module ex1010_qmap_map (sk, i_9_, i_2_, i_0_, i_1_, i_8_, i_6_, i_7_, i_5_, i_3_, i_4_, o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_);

	input i_9_;
	input i_2_;
	input i_0_;
	input i_1_;
	input i_8_;
	input i_6_;
	input i_7_;
	input i_5_;
	input i_3_;
	input i_4_;
	output o_0_;
	output o_1_;
	output o_2_;
	output o_3_;
	output o_4_;
	output o_5_;
	output o_6_;
	output o_7_;
	output o_8_;
	output o_9_;



	wire g217, g298, g364, g431, g486, g542, g585, g627, g662, g689, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11;
	wire g12, g13, g14, g15, g16, g17, g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29, g30, g31, g32;
	wire g33, g34, g35, g36, g37, g38, g39, g40, g41, g42, g43, g44, g45, g46, g47, g48, g49, g50, g51, g52, g53;
	wire g54, g55, g56, g57, g58, g59, g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g70, g71, g72, g73, g74;
	wire g75, g76, g77, g78, g79, g80, g81, g82, g83, g84, g85, g86, g765, g87, g88, g787, g774, g89, g90, g91, g92;
	wire g93, g94, g95, g96, g97, g98, g99, g100, g101, g102, g103, g104, g105, g106, g107, g108, g109, g110, g111, g112, g113;
	wire g114, g115, g116, g117, g118, g119, g120, g121, g122, g123, g124, g125, g126, g127, g128, g129, g130, g131, g132, g133, g134;
	wire g135, g136, g137, g138, g139, g140, g141, g142, g143, g144, g145, g146, g147, g148, g149, g150, g151, g152, g153, g154, g155;
	wire g156, g157, g158, g159, g160, g161, g162, g163, g164, g165, g166, g167, g168, g169, g170, g171, g172, g747, g173, g174, g175;
	wire g176, g177, g178, g179, g180, g181, g182, g183, g184, g185, g186, g187, g188, g189, g190, g191, g192, g193, g194, g195, g196;
	wire g197, g198, g199, g200, g201, g202, g203, g204, g205, g206, g207, g208, g209, g210, g211, g212, g213, g214, g215, g216, g758;
	wire g218, g219, g220, g221, g222, g223, g224, g225, g226, g227, g228, g229, g230, g231, g232, g233, g234, g235, g236, g237, g238;
	wire g239, g240, g241, g242, g243, g244, g245, g246, g247, g248, g249, g250, g251, g252, g253, g254, g255, g256, g257, g258, g259;
	wire g260, g261, g262, g263, g264, g265, g266, g267, g268, g269, g270, g271, g272, g273, g274, g275, g276, g277, g278, g279, g280;
	wire g281, g282, g283, g284, g285, g286, g287, g288, g289, g729, g290, g291, g292, g293, g294, g295, g296, g722, g297, g735, g299;
	wire g300, g301, g302, g303, g304, g305, g306, g307, g308, g309, g310, g311, g312, g313, g314, g315, g316, g317, g318, g319, g320;
	wire g321, g322, g323, g324, g325, g326, g327, g328, g329, g330, g331, g332, g333, g334, g335, g336, g337, g338, g339, g340, g341;
	wire g342, g343, g344, g345, g346, g347, g348, g349, g350, g351, g352, g353, g354, g355, g356, g357, g358, g359, g360, g711, g361;
	wire g362, g363, g365, g366, g367, g368, g369, g370, g371, g372, g373, g374, g375, g376, g377, g378, g379, g380, g381, g382, g383;
	wire g384, g385, g386, g387, g388, g389, g390, g391, g392, g393, g394, g395, g396, g397, g398, g399, g400, g401, g402, g403, g404;
	wire g405, g406, g407, g408, g409, g410, g411, g412, g413, g414, g415, g416, g417, g418, g419, g420, g421, g422, g423, g424, g425;
	wire g426, g427, g428, g429, g430, g432, g433, g434, g435, g436, g437, g438, g439, g440, g441, g442, g443, g444, g445, g446, g447;
	wire g448, g449, g450, g451, g452, g453, g454, g455, g456, g457, g458, g459, g460, g461, g462, g463, g464, g465, g466, g467, g468;
	wire g469, g470, g471, g472, g473, g474, g475, g476, g477, g478, g479, g480, g481, g482, g483, g704, g484, g485, g487, g488, g489;
	wire g490, g491, g492, g493, g494, g495, g496, g497, g498, g499, g500, g501, g502, g503, g504, g505, g506, g507, g508, g509, g510;
	wire g511, g512, g513, g514, g515, g516, g517, g518, g519, g520, g521, g522, g523, g524, g525, g526, g527, g528, g529, g530, g531;
	wire g532, g533, g534, g535, g536, g537, g538, g697, g539, g540, g541, g543, g544, g545, g546, g690, g547, g548, g549, g550, g551;
	wire g552, g553, g554, g555, g556, g557, g558, g559, g560, g561, g562, g563, g564, g565, g566, g567, g568, g569, g570, g571, g572;
	wire g573, g574, g575, g576, g577, g578, g579, g580, g581, g582, g583, g584, g586, g587, g588, g589, g590, g591, g592, g593, g594;
	wire g595, g596, g597, g598, g599, g600, g601, g602, g603, g604, g605, g606, g607, g608, g609, g610, g611, g612, g613, g614, g615;
	wire g616, g617, g618, g619, g620, g621, g622, g623, g624, g625, g626, g628, g629, g630, g631, g632, g633, g634, g635, g636, g637;
	wire g638, g639, g640, g641, g642, g643, g644, g645, g646, g647, g648, g649, g650, g651, g652, g653, g654, g655, g656, g657, g658;
	wire g659, g660, g661, g663, g664, g665, g666, g667, g668, g669, g670, g671, g672, g673, g674, g675, g676, g677, g678, g679, g680;
	wire g681, g682, g683, g684, g685, g686, g687, g688, g691, g692, g693, g694, g695, g696, g698, g699, g700, g701, g702, g703, g705;
	wire g706, g707, g708, g709, g710, g712, g713, g714, g717, g715, g716, g719, g720, g718, g721, g723, g724, g725, g726, g727, g728;
	wire g730, g731, g732, g733, g734, g736, g737, g738, g741, g739, g740, g744, g745, g742, g743, g746, g748, g749, g750, g753, g751;
	wire g752, g755, g756, g754, g757, g759, g760, g761, g762, g763, g764, g766, g767, g768, g770, g769, g772, g771, g773, g775, g776;
	wire g777, g780, g778, g779, g783, g784, g781, g782, g785, g786, g788, g789, g790, g793, g791, g792, g796, g797, g794, g795, g798;
	wire g799;

	lut_sub lut_5 ({g217}, o_0_);
	defparam lut_5.LUT_SIZE = 1;
	defparam lut_5.mask = 2'b10;

	lut_sub lut_9 ({g298}, o_1_);
	defparam lut_9.LUT_SIZE = 1;
	defparam lut_9.mask = 2'b10;

	lut_sub lut_13 ({g364}, o_2_);
	defparam lut_13.LUT_SIZE = 1;
	defparam lut_13.mask = 2'b10;

	lut_sub lut_17 ({g431}, o_3_);
	defparam lut_17.LUT_SIZE = 1;
	defparam lut_17.mask = 2'b10;

	lut_sub lut_21 ({g486}, o_4_);
	defparam lut_21.LUT_SIZE = 1;
	defparam lut_21.mask = 2'b10;

	lut_sub lut_25 ({g542}, o_5_);
	defparam lut_25.LUT_SIZE = 1;
	defparam lut_25.mask = 2'b10;

	lut_sub lut_29 ({g585}, o_6_);
	defparam lut_29.LUT_SIZE = 1;
	defparam lut_29.mask = 2'b10;

	lut_sub lut_33 ({g627}, o_7_);
	defparam lut_33.LUT_SIZE = 1;
	defparam lut_33.mask = 2'b10;

	lut_sub lut_37 ({g662}, o_8_);
	defparam lut_37.LUT_SIZE = 1;
	defparam lut_37.mask = 2'b10;

	lut_sub lut_41 ({g689}, o_9_);
	defparam lut_41.LUT_SIZE = 1;
	defparam lut_41.mask = 2'b10;

	lut_sub lut_45 ({i_2_, i_0_, i_1_}, g1);
	defparam lut_45.LUT_SIZE = 3;
	defparam lut_45.mask = 8'h7f;

	lut_sub lut_56 ({i_9_, g1}, g2);
	defparam lut_56.LUT_SIZE = 2;
	defparam lut_56.mask = 4'b1000;

	lut_sub lut_60 ({i_8_, i_6_, i_7_}, g3);
	defparam lut_60.LUT_SIZE = 3;
	defparam lut_60.mask = 8'hf7;

	lut_sub lut_70 ({i_5_, i_3_, i_4_}, g4);
	defparam lut_70.LUT_SIZE = 3;
	defparam lut_70.mask = 8'hef;

	lut_sub lut_82 ({g3, g4}, g5);
	defparam lut_82.LUT_SIZE = 2;
	defparam lut_82.mask = 4'b1000;

	lut_sub lut_86 ({i_2_, i_0_, i_1_}, g6);
	defparam lut_86.LUT_SIZE = 3;
	defparam lut_86.mask = 8'hf7;

	lut_sub lut_96 ({i_5_, i_3_, i_4_}, g7);
	defparam lut_96.LUT_SIZE = 3;
	defparam lut_96.mask = 8'h20;

	lut_sub lut_100 ({i_8_, i_6_, i_7_}, g8);
	defparam lut_100.LUT_SIZE = 3;
	defparam lut_100.mask = 8'h20;

	lut_sub lut_106 ({g7, g8}, g9);
	defparam lut_106.LUT_SIZE = 2;
	defparam lut_106.mask = 4'b0001;

	lut_sub lut_110 ({i_5_, i_3_, i_4_}, g10);
	defparam lut_110.LUT_SIZE = 3;
	defparam lut_110.mask = 8'h7f;

	lut_sub lut_120 ({i_2_, i_0_, i_1_}, g11);
	defparam lut_120.LUT_SIZE = 3;
	defparam lut_120.mask = 8'h04;

	lut_sub lut_126 ({g10, g11}, g12);
	defparam lut_126.LUT_SIZE = 2;
	defparam lut_126.mask = 4'b1011;

	lut_sub lut_132 ({i_2_, i_0_, i_1_, i_9_}, g13);
	defparam lut_132.LUT_SIZE = 4;
	defparam lut_132.mask = 16'hfdff;

	lut_sub lut_150 ({i_5_, i_3_, i_4_}, g14);
	defparam lut_150.LUT_SIZE = 3;
	defparam lut_150.mask = 8'hfe;

	lut_sub lut_162 ({g3, g14}, g15);
	defparam lut_162.LUT_SIZE = 2;
	defparam lut_162.mask = 4'b1000;

	lut_sub lut_166 ({i_8_, i_6_, i_7_}, g16);
	defparam lut_166.LUT_SIZE = 3;
	defparam lut_166.mask = 8'h40;

	lut_sub lut_172 ({g16, g4}, g17);
	defparam lut_172.LUT_SIZE = 2;
	defparam lut_172.mask = 4'b0010;

	lut_sub lut_176 ({i_8_, i_6_, i_7_}, g18);
	defparam lut_176.LUT_SIZE = 3;
	defparam lut_176.mask = 8'h80;

	lut_sub lut_182 ({g7, g18}, g19);
	defparam lut_182.LUT_SIZE = 2;
	defparam lut_182.mask = 4'b0001;

	lut_sub lut_186 ({i_9_, i_8_, i_6_, i_7_}, g20);
	defparam lut_186.LUT_SIZE = 4;
	defparam lut_186.mask = 16'h0004;

	lut_sub lut_190 ({i_2_, i_0_, i_1_, i_9_}, g21);
	defparam lut_190.LUT_SIZE = 4;
	defparam lut_190.mask = 16'hfff7;

	lut_sub lut_208 ({i_2_, i_0_, i_1_}, g22);
	defparam lut_208.LUT_SIZE = 3;
	defparam lut_208.mask = 8'h01;

	lut_sub lut_214 ({g22, g14}, g23);
	defparam lut_214.LUT_SIZE = 2;
	defparam lut_214.mask = 4'b0010;

	lut_sub lut_222 ({g20, g21, g19, g23}, g24);
	defparam lut_222.LUT_SIZE = 4;
	defparam lut_222.mask = 16'h3075;

	lut_sub lut_232 ({i_2_, i_0_, i_1_}, g25);
	defparam lut_232.LUT_SIZE = 3;
	defparam lut_232.mask = 8'h02;

	lut_sub lut_238 ({g25, g14}, g26);
	defparam lut_238.LUT_SIZE = 2;
	defparam lut_238.mask = 4'b0010;

	lut_sub lut_242 ({i_9_, i_8_, i_6_, i_7_}, g27);
	defparam lut_242.LUT_SIZE = 4;
	defparam lut_242.mask = 16'h0002;

	lut_sub lut_246 ({i_5_, i_3_, i_4_}, g28);
	defparam lut_246.LUT_SIZE = 3;
	defparam lut_246.mask = 8'hbf;

	lut_sub lut_258 ({g28, g6}, g29);
	defparam lut_258.LUT_SIZE = 2;
	defparam lut_258.mask = 4'b1000;

	lut_sub lut_262 ({i_5_, i_3_, i_4_}, g30);
	defparam lut_262.LUT_SIZE = 3;
	defparam lut_262.mask = 8'h08;

	lut_sub lut_268 ({g16, g30}, g31);
	defparam lut_268.LUT_SIZE = 2;
	defparam lut_268.mask = 4'b0001;

	lut_sub lut_274 ({g8, g10}, g32);
	defparam lut_274.LUT_SIZE = 2;
	defparam lut_274.mask = 4'b0010;

	lut_sub lut_280 ({i_2_, i_0_, i_1_, i_9_, g31, g32}, g33);
	defparam lut_280.LUT_SIZE = 6;
	defparam lut_280.mask = 64'h0000500000300000;

	lut_sub lut_292 ({g20, g26, g27, g29, g33}, g34);
	defparam lut_292.LUT_SIZE = 5;
	defparam lut_292.mask = 32'haaa08880;

	lut_sub lut_304 ({i_2_, i_0_, i_1_, i_9_}, g35);
	defparam lut_304.LUT_SIZE = 4;
	defparam lut_304.mask = 16'h2000;

	lut_sub lut_308 ({i_5_, i_3_, i_4_}, g36);
	defparam lut_308.LUT_SIZE = 3;
	defparam lut_308.mask = 8'h04;

	lut_sub lut_314 ({g36, g16}, g37);
	defparam lut_314.LUT_SIZE = 2;
	defparam lut_314.mask = 4'b1110;

	lut_sub lut_320 ({i_9_, i_8_, i_6_, i_7_}, g38);
	defparam lut_320.LUT_SIZE = 4;
	defparam lut_320.mask = 16'hffdf;

	lut_sub lut_338 ({i_2_, i_0_, i_1_}, g39);
	defparam lut_338.LUT_SIZE = 3;
	defparam lut_338.mask = 8'h40;

	lut_sub lut_342 ({i_9_, i_8_, i_6_, i_7_}, g40);
	defparam lut_342.LUT_SIZE = 4;
	defparam lut_342.mask = 16'h0080;

	lut_sub lut_351 ({g38, g39, g25, g10, g40}, g41);
	defparam lut_351.LUT_SIZE = 5;
	defparam lut_351.mask = 32'h0c4c0044;

	lut_sub lut_361 ({i_2_, i_0_, i_1_, i_9_}, g42);
	defparam lut_361.LUT_SIZE = 4;
	defparam lut_361.mask = 16'h0080;

	lut_sub lut_366 ({i_9_, g11}, g43);
	defparam lut_366.LUT_SIZE = 2;
	defparam lut_366.mask = 4'b1011;

	lut_sub lut_374 ({g28, g3}, g44);
	defparam lut_374.LUT_SIZE = 2;
	defparam lut_374.mask = 4'b1000;

	lut_sub lut_378 ({i_8_, i_6_, i_7_}, g45);
	defparam lut_378.LUT_SIZE = 3;
	defparam lut_378.mask = 8'hfd;

	lut_sub lut_390 ({g28, g45}, g46);
	defparam lut_390.LUT_SIZE = 2;
	defparam lut_390.mask = 4'b1000;

	lut_sub lut_398 ({g42, g43, g44, g46}, g47);
	defparam lut_398.LUT_SIZE = 4;
	defparam lut_398.mask = 16'h3075;

	lut_sub lut_412 ({g20, g28, g1, g47}, g48);
	defparam lut_412.LUT_SIZE = 4;
	defparam lut_412.mask = 16'haa2a;

	lut_sub lut_422 ({i_2_, i_0_, i_1_, i_9_}, g49);
	defparam lut_422.LUT_SIZE = 4;
	defparam lut_422.mask = 16'h0002;

	lut_sub lut_426 ({i_8_, i_6_, i_7_}, g50);
	defparam lut_426.LUT_SIZE = 3;
	defparam lut_426.mask = 8'hef;

	lut_sub lut_438 ({g50, g14}, g51);
	defparam lut_438.LUT_SIZE = 2;
	defparam lut_438.mask = 4'b1000;

	lut_sub lut_444 ({g39, g14}, g52);
	defparam lut_444.LUT_SIZE = 2;
	defparam lut_444.mask = 4'b0010;

	lut_sub lut_449 ({i_9_, g50}, g53);
	defparam lut_449.LUT_SIZE = 2;
	defparam lut_449.mask = 4'b0010;

	lut_sub lut_453 ({i_8_, i_6_, i_7_}, g54);
	defparam lut_453.LUT_SIZE = 3;
	defparam lut_453.mask = 8'hfb;

	lut_sub lut_465 ({g54, g30}, g55);
	defparam lut_465.LUT_SIZE = 2;
	defparam lut_465.mask = 4'b0100;

	lut_sub lut_473 ({g49, g52, g53, g55}, g56);
	defparam lut_473.LUT_SIZE = 4;
	defparam lut_473.mask = 16'h0357;

	lut_sub lut_485 ({g6, g4}, g57);
	defparam lut_485.LUT_SIZE = 2;
	defparam lut_485.mask = 4'b1000;

	lut_sub lut_489 ({i_9_, i_8_, i_6_, i_7_}, g58);
	defparam lut_489.LUT_SIZE = 4;
	defparam lut_489.mask = 16'hfffe;

	lut_sub lut_507 ({i_2_, i_0_, i_1_}, g59);
	defparam lut_507.LUT_SIZE = 3;
	defparam lut_507.mask = 8'h10;

	lut_sub lut_513 ({g7, g59}, g60);
	defparam lut_513.LUT_SIZE = 2;
	defparam lut_513.mask = 4'b0001;

	lut_sub lut_522 ({g39, g30, g57, g58, g60}, g61);
	defparam lut_522.LUT_SIZE = 5;
	defparam lut_522.mask = 32'h4c4c4ccc;

	lut_sub lut_540 ({g59, g4}, g62);
	defparam lut_540.LUT_SIZE = 2;
	defparam lut_540.mask = 4'b0010;

	lut_sub lut_544 ({i_2_, i_0_, i_1_}, g63);
	defparam lut_544.LUT_SIZE = 3;
	defparam lut_544.mask = 8'h20;

	lut_sub lut_550 ({g63, g14}, g64);
	defparam lut_550.LUT_SIZE = 2;
	defparam lut_550.mask = 4'b0010;

	lut_sub lut_557 ({g62, g53, g64}, g65);
	defparam lut_557.LUT_SIZE = 3;
	defparam lut_557.mask = 8'h13;

	lut_sub lut_568 ({g49, g51, g56, g61, g65}, g66);
	defparam lut_568.LUT_SIZE = 5;
	defparam lut_568.mask = 32'h80808000;

	lut_sub lut_579 ({g35, g37, g41, g48, g66}, g67);
	defparam lut_579.LUT_SIZE = 5;
	defparam lut_579.mask = 32'h10100010;

	lut_sub lut_585 ({i_6_, i_7_}, g68);
	defparam lut_585.LUT_SIZE = 2;
	defparam lut_585.mask = 4'b0100;

	lut_sub lut_590 ({i_9_, g68}, g69);
	defparam lut_590.LUT_SIZE = 2;
	defparam lut_590.mask = 4'b0001;

	lut_sub lut_599 ({g22, g36, g20, g58, g12}, g70);
	defparam lut_599.LUT_SIZE = 5;
	defparam lut_599.mask = 32'h8888888f;

	lut_sub lut_615 ({g6, g14}, g71);
	defparam lut_615.LUT_SIZE = 2;
	defparam lut_615.mask = 4'b1000;

	lut_sub lut_622 ({i_8_, g28, g59, g71}, g72);
	defparam lut_622.LUT_SIZE = 4;
	defparam lut_622.mask = 16'h5530;

	lut_sub lut_631 ({i_9_, i_8_, i_6_, i_7_}, g73);
	defparam lut_631.LUT_SIZE = 4;
	defparam lut_631.mask = 16'h0008;

	lut_sub lut_637 ({g4, g1}, g74);
	defparam lut_637.LUT_SIZE = 2;
	defparam lut_637.mask = 4'b0111;

	lut_sub lut_643 ({i_0_, i_1_}, g75);
	defparam lut_643.LUT_SIZE = 2;
	defparam lut_643.mask = 4'b0010;

	lut_sub lut_647 ({i_5_, i_3_, i_4_}, g76);
	defparam lut_647.LUT_SIZE = 3;
	defparam lut_647.mask = 8'hfd;

	lut_sub lut_659 ({g76, g45}, g77);
	defparam lut_659.LUT_SIZE = 2;
	defparam lut_659.mask = 4'b1000;

	lut_sub lut_663 ({i_0_, i_1_}, g78);
	defparam lut_663.LUT_SIZE = 2;
	defparam lut_663.mask = 4'b0001;

	lut_sub lut_668 ({i_2_, g78, i_9_}, g79);
	defparam lut_668.LUT_SIZE = 3;
	defparam lut_668.mask = 8'ha2;

	lut_sub lut_679 ({i_2_, g7, g75, g16, g77, g79}, g80);
	defparam lut_679.LUT_SIZE = 6;
	defparam lut_679.mask = 64'h0011001100000505;

	lut_sub lut_690 ({i_6_, i_7_}, g81);
	defparam lut_690.LUT_SIZE = 2;
	defparam lut_690.mask = 4'b0010;

	lut_sub lut_696 ({g63, g4}, g82);
	defparam lut_696.LUT_SIZE = 2;
	defparam lut_696.mask = 4'b0010;

	lut_sub lut_700 ({i_6_, i_7_}, g83);
	defparam lut_700.LUT_SIZE = 2;
	defparam lut_700.mask = 4'b0001;

	lut_sub lut_706 ({g76, g63}, g84);
	defparam lut_706.LUT_SIZE = 2;
	defparam lut_706.mask = 4'b0100;

	lut_sub lut_712 ({g54, g14}, g85);
	defparam lut_712.LUT_SIZE = 2;
	defparam lut_712.mask = 4'b1000;

	lut_sub lut_720 ({g35, g20, g84, g85}, g86);
	defparam lut_720.LUT_SIZE = 4;
	defparam lut_720.mask = 16'h0357;

	lut_sub lut_735 ({g73, g74, g80, g765, g86}, g87);
	defparam lut_735.LUT_SIZE = 5;
	defparam lut_735.mask = 32'h20200020;

	lut_sub lut_745 ({g69, g70, g72, g87}, g88);
	defparam lut_745.LUT_SIZE = 4;
	defparam lut_745.mask = 16'h5040;

	lut_sub lut_757 ({g787, g774, g24, g34, g67, g88}, g89);
	defparam lut_757.LUT_SIZE = 6;
	defparam lut_757.mask = 64'h0000000000000100;

	lut_sub lut_763 ({g36, g63}, g90);
	defparam lut_763.LUT_SIZE = 2;
	defparam lut_763.mask = 4'b0001;

	lut_sub lut_772 ({g22, g28, g73, g27, g90}, g91);
	defparam lut_772.LUT_SIZE = 5;
	defparam lut_772.mask = 32'h11111f11;

	lut_sub lut_786 ({i_3_, i_4_}, g92);
	defparam lut_786.LUT_SIZE = 2;
	defparam lut_786.mask = 4'b0001;

	lut_sub lut_794 ({g22, i_9_, g50, i_5_, g92, g18}, g93);
	defparam lut_794.LUT_SIZE = 6;
	defparam lut_794.mask = 64'h0000000030000101;

	lut_sub lut_803 ({g39, g4}, g94);
	defparam lut_803.LUT_SIZE = 2;
	defparam lut_803.mask = 4'b0010;

	lut_sub lut_809 ({i_6_, i_7_, g6, g10}, g95);
	defparam lut_809.LUT_SIZE = 4;
	defparam lut_809.mask = 16'h7fff;

	lut_sub lut_830 ({i_9_, i_8_, g83, g94, g95}, g96);
	defparam lut_830.LUT_SIZE = 5;
	defparam lut_830.mask = 32'h000003aa;

	lut_sub lut_841 ({g50, g10}, g97);
	defparam lut_841.LUT_SIZE = 2;
	defparam lut_841.mask = 4'b1000;

	lut_sub lut_849 ({g42, g13, g85, g97}, g98);
	defparam lut_849.LUT_SIZE = 4;
	defparam lut_849.mask = 16'h5073;

	lut_sub lut_861 ({g63, g30}, g99);
	defparam lut_861.LUT_SIZE = 2;
	defparam lut_861.mask = 4'b0001;

	lut_sub lut_868 ({g99, g40, g12}, g100);
	defparam lut_868.LUT_SIZE = 3;
	defparam lut_868.mask = 8'h23;

	lut_sub lut_876 ({g50, g36}, g101);
	defparam lut_876.LUT_SIZE = 2;
	defparam lut_876.mask = 4'b0100;

	lut_sub lut_884 ({i_2_, i_9_, g7, g101, g75, g3}, g102);
	defparam lut_884.LUT_SIZE = 6;
	defparam lut_884.mask = 64'h0303002203030000;

	lut_sub lut_900 ({g20, g25, g4}, g103);
	defparam lut_900.LUT_SIZE = 3;
	defparam lut_900.mask = 8'h02;

	lut_sub lut_909 ({g36, g20, g59, g53, g103}, g104);
	defparam lut_909.LUT_SIZE = 5;
	defparam lut_909.mask = 32'haaaaa8a0;

	lut_sub lut_930 ({g22, g50, g38, g35, g76}, g105);
	defparam lut_930.LUT_SIZE = 5;
	defparam lut_930.mask = 32'h2200a2a0;

	lut_sub lut_945 ({g7, g1, g14, g53, g27}, g106);
	defparam lut_945.LUT_SIZE = 5;
	defparam lut_945.mask = 32'h50007300;

	lut_sub lut_960 ({g100, g102, g104, g105, g106}, g107);
	defparam lut_960.LUT_SIZE = 5;
	defparam lut_960.mask = 32'h08000000;

	lut_sub lut_969 ({g91, g93, g96, g98, g107}, g108);
	defparam lut_969.LUT_SIZE = 5;
	defparam lut_969.mask = 32'h40000000;

	lut_sub lut_976 ({i_9_, g3, g63, g30}, g109);
	defparam lut_976.LUT_SIZE = 4;
	defparam lut_976.mask = 16'hef00;

	lut_sub lut_989 ({i_9_, g7, g39, g16}, g110);
	defparam lut_989.LUT_SIZE = 4;
	defparam lut_989.mask = 16'h00fe;

	lut_sub lut_1002 ({i_9_, i_8_, g81, g84, g62}, g111);
	defparam lut_1002.LUT_SIZE = 5;
	defparam lut_1002.mask = 32'h03000005;

	lut_sub lut_1011 ({g36, g1}, g112);
	defparam lut_1011.LUT_SIZE = 2;
	defparam lut_1011.mask = 4'b0010;

	lut_sub lut_1020 ({g20, g73, g30, g11, g112}, g113);
	defparam lut_1020.LUT_SIZE = 5;
	defparam lut_1020.mask = 32'h00550357;

	lut_sub lut_1038 ({g109, g110, g111, g113}, g114);
	defparam lut_1038.LUT_SIZE = 4;
	defparam lut_1038.mask = 16'h0888;

	lut_sub lut_1048 ({g38, g57, g53, g90}, g115);
	defparam lut_1048.LUT_SIZE = 4;
	defparam lut_1048.mask = 16'h5703;

	lut_sub lut_1060 ({g76, g16}, g116);
	defparam lut_1060.LUT_SIZE = 2;
	defparam lut_1060.mask = 4'b0100;

	lut_sub lut_1066 ({g10, g45}, g117);
	defparam lut_1066.LUT_SIZE = 2;
	defparam lut_1066.mask = 4'b1000;

	lut_sub lut_1074 ({g20, g13, g57, g117}, g118);
	defparam lut_1074.LUT_SIZE = 4;
	defparam lut_1074.mask = 16'h5073;

	lut_sub lut_1084 ({i_0_, i_1_}, g119);
	defparam lut_1084.LUT_SIZE = 2;
	defparam lut_1084.mask = 4'b0111;

	lut_sub lut_1092 ({g54, g76}, g120);
	defparam lut_1092.LUT_SIZE = 2;
	defparam lut_1092.mask = 4'b1000;

	lut_sub lut_1099 ({i_2_, i_9_, g119, g120, g9}, g121);
	defparam lut_1099.LUT_SIZE = 5;
	defparam lut_1099.mask = 32'h00503000;

	lut_sub lut_1108 ({g50, g28}, g122);
	defparam lut_1108.LUT_SIZE = 2;
	defparam lut_1108.mask = 4'b1000;

	lut_sub lut_1115 ({i_2_, g78, i_9_, g122, g17}, g123);
	defparam lut_1115.LUT_SIZE = 5;
	defparam lut_1115.mask = 32'h00300005;

	lut_sub lut_1124 ({g39, g76}, g124);
	defparam lut_1124.LUT_SIZE = 2;
	defparam lut_1124.mask = 4'b0010;

	lut_sub lut_1130 ({g50, g30}, g125);
	defparam lut_1130.LUT_SIZE = 2;
	defparam lut_1130.mask = 4'b0100;

	lut_sub lut_1140 ({g101, g35, g20, g124, g125, g13}, g126);
	defparam lut_1140.LUT_SIZE = 6;
	defparam lut_1140.mask = 64'hddd0ddd0ddd00000;

	lut_sub lut_1174 ({g20, g28, g25, g99}, g127);
	defparam lut_1174.LUT_SIZE = 4;
	defparam lut_1174.mask = 16'h0075;

	lut_sub lut_1187 ({g73, g84, g123, g126, g127}, g128);
	defparam lut_1187.LUT_SIZE = 5;
	defparam lut_1187.mask = 32'h20202000;

	lut_sub lut_1198 ({g42, g116, g118, g121, g128}, g129);
	defparam lut_1198.LUT_SIZE = 5;
	defparam lut_1198.mask = 32'h40404000;

	lut_sub lut_1208 ({i_9_, i_8_, g81, g36, g57, g11}, g130);
	defparam lut_1208.LUT_SIZE = 6;
	defparam lut_1208.mask = 64'h0005000000000033;

	lut_sub lut_1217 ({i_2_, i_0_, i_9_}, g131);
	defparam lut_1217.LUT_SIZE = 3;
	defparam lut_1217.mask = 8'h80;

	lut_sub lut_1227 ({g50, g35, g10, g2, g14, g131}, g132);
	defparam lut_1227.LUT_SIZE = 6;
	defparam lut_1227.mask = 64'h4404550400000000;

	lut_sub lut_1239 ({i_9_, g63}, g133);
	defparam lut_1239.LUT_SIZE = 2;
	defparam lut_1239.mask = 4'b1011;

	lut_sub lut_1247 ({g8, g28}, g134);
	defparam lut_1247.LUT_SIZE = 2;
	defparam lut_1247.mask = 4'b0010;

	lut_sub lut_1253 ({g8, g14}, g135);
	defparam lut_1253.LUT_SIZE = 2;
	defparam lut_1253.mask = 4'b0010;

	lut_sub lut_1263 ({g49, g13, g133, g134, g32, g135}, g136);
	defparam lut_1263.LUT_SIZE = 6;
	defparam lut_1263.mask = 64'h88ccaaff80c0a0f0;

	lut_sub lut_1294 ({i_9_, g16}, g137);
	defparam lut_1294.LUT_SIZE = 2;
	defparam lut_1294.mask = 4'b0001;

	lut_sub lut_1298 ({i_8_, i_6_, i_7_}, g138);
	defparam lut_1298.LUT_SIZE = 3;
	defparam lut_1298.mask = 8'h01;

	lut_sub lut_1304 ({g138, g14}, g139);
	defparam lut_1304.LUT_SIZE = 2;
	defparam lut_1304.mask = 4'b0010;

	lut_sub lut_1313 ({g7, g43, g137, g1, g139}, g140);
	defparam lut_1313.LUT_SIZE = 5;
	defparam lut_1313.mask = 32'h55005d0c;

	lut_sub lut_1329 ({g76, g138}, g141);
	defparam lut_1329.LUT_SIZE = 2;
	defparam lut_1329.mask = 4'b0100;

	lut_sub lut_1335 ({g36, g25}, g142);
	defparam lut_1335.LUT_SIZE = 2;
	defparam lut_1335.mask = 4'b1110;

	lut_sub lut_1345 ({g76, g11, g40, g142}, g143);
	defparam lut_1345.LUT_SIZE = 4;
	defparam lut_1345.mask = 16'h2322;

	lut_sub lut_1355 ({g25, g30}, g144);
	defparam lut_1355.LUT_SIZE = 2;
	defparam lut_1355.mask = 4'b0001;

	lut_sub lut_1365 ({g38, g42, g77, g27, g29, g144}, g145);
	defparam lut_1365.LUT_SIZE = 6;
	defparam lut_1365.mask = 64'h88888800fafafa00;

	lut_sub lut_1397 ({g21, g15, g141, g143, g145}, g146);
	defparam lut_1397.LUT_SIZE = 5;
	defparam lut_1397.mask = 32'h40004444;

	lut_sub lut_1410 ({g130, g132, g136, g140, g146}, g147);
	defparam lut_1410.LUT_SIZE = 5;
	defparam lut_1410.mask = 32'h04000000;

	lut_sub lut_1416 ({g54, g28}, g148);
	defparam lut_1416.LUT_SIZE = 2;
	defparam lut_1416.mask = 4'b1000;

	lut_sub lut_1425 ({i_9_, g36, g39, g45, g1, g148}, g149);
	defparam lut_1425.LUT_SIZE = 6;
	defparam lut_1425.mask = 64'h44444444000000f0;

	lut_sub lut_1445 ({g36, g20, g18, g21, g144}, g150);
	defparam lut_1445.LUT_SIZE = 5;
	defparam lut_1445.mask = 32'h00550c5d;

	lut_sub lut_1460 ({i_2_, i_9_, g75}, g151);
	defparam lut_1460.LUT_SIZE = 3;
	defparam lut_1460.mask = 8'hc4;

	lut_sub lut_1469 ({g78, g3, g30}, g152);
	defparam lut_1469.LUT_SIZE = 3;
	defparam lut_1469.mask = 8'h04;

	lut_sub lut_1477 ({i_2_, g76, g16, g151, g152}, g153);
	defparam lut_1477.LUT_SIZE = 5;
	defparam lut_1477.mask = 32'h11110300;

	lut_sub lut_1489 ({i_8_, i_6_, i_7_, g36, g133, g43}, g154);
	defparam lut_1489.LUT_SIZE = 6;
	defparam lut_1489.mask = 64'h0a00000000000c00;

	lut_sub lut_1500 ({g149, g150, g153, g154}, g155);
	defparam lut_1500.LUT_SIZE = 4;
	defparam lut_1500.mask = 16'h8000;

	lut_sub lut_1506 ({g54, g4}, g156);
	defparam lut_1506.LUT_SIZE = 2;
	defparam lut_1506.mask = 4'b1000;

	lut_sub lut_1512 ({g8, g4}, g157);
	defparam lut_1512.LUT_SIZE = 2;
	defparam lut_1512.mask = 4'b0010;

	lut_sub lut_1518 ({g8, g30}, g158);
	defparam lut_1518.LUT_SIZE = 2;
	defparam lut_1518.mask = 4'b0001;

	lut_sub lut_1526 ({g42, g156, g157, g158}, g159);
	defparam lut_1526.LUT_SIZE = 4;
	defparam lut_1526.mask = 16'h007f;

	lut_sub lut_1537 ({i_9_, i_8_, i_6_, g36}, g160);
	defparam lut_1537.LUT_SIZE = 4;
	defparam lut_1537.mask = 16'h1040;

	lut_sub lut_1544 ({g36, g54}, g161);
	defparam lut_1544.LUT_SIZE = 2;
	defparam lut_1544.mask = 4'b0010;

	lut_sub lut_1552 ({i_9_, g25, g3, g10, g161}, g162);
	defparam lut_1552.LUT_SIZE = 5;
	defparam lut_1552.mask = 32'h005500c0;

	lut_sub lut_1564 ({i_7_, g6, g160, g162}, g163);
	defparam lut_1564.LUT_SIZE = 4;
	defparam lut_1564.mask = 16'h8aaa;

	lut_sub lut_1578 ({g28, g25, g84, g53}, g164);
	defparam lut_1578.LUT_SIZE = 4;
	defparam lut_1578.mask = 16'h1511;

	lut_sub lut_1588 ({g18, g14}, g165);
	defparam lut_1588.LUT_SIZE = 2;
	defparam lut_1588.mask = 4'b0010;

	lut_sub lut_1596 ({g49, g50, g7, g165}, g166);
	defparam lut_1596.LUT_SIZE = 4;
	defparam lut_1596.mask = 16'h0075;

	lut_sub lut_1610 ({g38, g36, g39, g28, g137, g40}, g167);
	defparam lut_1610.LUT_SIZE = 6;
	defparam lut_1610.mask = 64'h003000ff00300075;

	lut_sub lut_1632 ({g7, g45}, g168);
	defparam lut_1632.LUT_SIZE = 2;
	defparam lut_1632.mask = 4'b0010;

	lut_sub lut_1638 ({g28, g16}, g169);
	defparam lut_1638.LUT_SIZE = 2;
	defparam lut_1638.mask = 4'b0100;

	lut_sub lut_1644 ({g7, g54}, g170);
	defparam lut_1644.LUT_SIZE = 2;
	defparam lut_1644.mask = 4'b0010;

	lut_sub lut_1650 ({g7, g138}, g171);
	defparam lut_1650.LUT_SIZE = 2;
	defparam lut_1650.mask = 4'b0001;

	lut_sub lut_1659 ({g99, g134, g43, g58, g171}, g172);
	defparam lut_1659.LUT_SIZE = 5;
	defparam lut_1659.mask = 32'haf0f2303;

	lut_sub lut_1682 ({g164, g166, g167, g747, g172}, g173);
	defparam lut_1682.LUT_SIZE = 5;
	defparam lut_1682.mask = 32'h10000000;

	lut_sub lut_1691 ({g2, g46, g159, g163, g173}, g174);
	defparam lut_1691.LUT_SIZE = 5;
	defparam lut_1691.mask = 32'h10101000;

	lut_sub lut_1700 ({g38, g6, g30}, g175);
	defparam lut_1700.LUT_SIZE = 3;
	defparam lut_1700.mask = 8'h40;

	lut_sub lut_1708 ({g39, g20, g10, g175}, g176);
	defparam lut_1708.LUT_SIZE = 4;
	defparam lut_1708.mask = 16'haaa2;

	lut_sub lut_1720 ({g3, g10}, g177);
	defparam lut_1720.LUT_SIZE = 2;
	defparam lut_1720.mask = 4'b1000;

	lut_sub lut_1728 ({g22, i_9_, g101, g16, g26}, g178);
	defparam lut_1728.LUT_SIZE = 5;
	defparam lut_1728.mask = 32'h00110f11;

	lut_sub lut_1741 ({g16, g10}, g179);
	defparam lut_1741.LUT_SIZE = 2;
	defparam lut_1741.mask = 4'b0010;

	lut_sub lut_1747 ({g36, g138}, g180);
	defparam lut_1747.LUT_SIZE = 2;
	defparam lut_1747.mask = 4'b0001;

	lut_sub lut_1755 ({g35, g179, g21, g180}, g181);
	defparam lut_1755.LUT_SIZE = 4;
	defparam lut_1755.mask = 16'h444f;

	lut_sub lut_1767 ({g30, g138}, g182);
	defparam lut_1767.LUT_SIZE = 2;
	defparam lut_1767.mask = 4'b0001;

	lut_sub lut_1773 ({g4, g18}, g183);
	defparam lut_1773.LUT_SIZE = 2;
	defparam lut_1773.mask = 4'b0100;

	lut_sub lut_1782 ({g42, g2, g182, g183, g44}, g184);
	defparam lut_1782.LUT_SIZE = 5;
	defparam lut_1782.mask = 32'hffc0aa80;

	lut_sub lut_1805 ({g49, g177, g178, g181, g184}, g185);
	defparam lut_1805.LUT_SIZE = 5;
	defparam lut_1805.mask = 32'h40404000;

	lut_sub lut_1813 ({g45, g14}, g186);
	defparam lut_1813.LUT_SIZE = 2;
	defparam lut_1813.mask = 4'b1000;

	lut_sub lut_1819 ({i_2_, i_0_, i_1_, i_9_, g179, g186}, g187);
	defparam lut_1819.LUT_SIZE = 6;
	defparam lut_1819.mask = 64'h0000300000500000;

	lut_sub lut_1831 ({g7, g36, g35, g42, g16}, g188);
	defparam lut_1831.LUT_SIZE = 5;
	defparam lut_1831.mask = 32'h00110515;

	lut_sub lut_1845 ({g38, g11, g14, g188}, g189);
	defparam lut_1845.LUT_SIZE = 4;
	defparam lut_1845.mask = 16'ha2aa;

	lut_sub lut_1859 ({g176, g185, g187, g189}, g190);
	defparam lut_1859.LUT_SIZE = 4;
	defparam lut_1859.mask = 16'h0004;

	lut_sub lut_1869 ({g115, g129, g147, g155, g174, g190}, g191);
	defparam lut_1869.LUT_SIZE = 6;
	defparam lut_1869.mask = 64'h0000000100000000;

	lut_sub lut_1873 ({i_9_, i_8_, i_6_}, g192);
	defparam lut_1873.LUT_SIZE = 3;
	defparam lut_1873.mask = 8'h04;

	lut_sub lut_1879 ({g36, g45}, g193);
	defparam lut_1879.LUT_SIZE = 2;
	defparam lut_1879.mask = 4'b0010;

	lut_sub lut_1887 ({i_9_, g7, g3, g11, g193}, g194);
	defparam lut_1887.LUT_SIZE = 5;
	defparam lut_1887.mask = 32'h00301111;

	lut_sub lut_1898 ({g36, g11}, g195);
	defparam lut_1898.LUT_SIZE = 2;
	defparam lut_1898.mask = 4'b0001;

	lut_sub lut_1907 ({g7, g38, g63, g53, g195}, g196);
	defparam lut_1907.LUT_SIZE = 5;
	defparam lut_1907.mask = 32'h11111f15;

	lut_sub lut_1923 ({i_9_, i_8_, i_6_, i_7_, g25}, g197);
	defparam lut_1923.LUT_SIZE = 5;
	defparam lut_1923.mask = 32'hc0c00040;

	lut_sub lut_1934 ({i_9_, i_8_, g30, g82, g197}, g198);
	defparam lut_1934.LUT_SIZE = 5;
	defparam lut_1934.mask = 32'h11000505;

	lut_sub lut_1947 ({i_2_, g78, g122, g139, g151}, g199);
	defparam lut_1947.LUT_SIZE = 5;
	defparam lut_1947.mask = 32'h00110505;

	lut_sub lut_1959 ({g50, g6, g30}, g200);
	defparam lut_1959.LUT_SIZE = 3;
	defparam lut_1959.mask = 8'h40;

	lut_sub lut_1965 ({g28, g138}, g201);
	defparam lut_1965.LUT_SIZE = 2;
	defparam lut_1965.mask = 4'b0100;

	lut_sub lut_1974 ({i_9_, g25, g59, g183, g141, g201}, g202);
	defparam lut_1974.LUT_SIZE = 6;
	defparam lut_1974.mask = 64'h003f003f00005555;

	lut_sub lut_2003 ({g21, g5, g198, g199, g200, g202}, g203);
	defparam lut_2003.LUT_SIZE = 6;
	defparam lut_2003.mask = 64'h8000000080008000;

	lut_sub lut_2011 ({i_9_, i_8_, i_7_, g59, g14}, g204);
	defparam lut_2011.LUT_SIZE = 5;
	defparam lut_2011.mask = 32'h00000200;

	lut_sub lut_2018 ({i_2_, i_9_, g50, g8, g119}, g205);
	defparam lut_2018.LUT_SIZE = 5;
	defparam lut_2018.mask = 32'ha0000022;

	lut_sub lut_2025 ({i_8_, i_7_}, g206);
	defparam lut_2025.LUT_SIZE = 2;
	defparam lut_2025.mask = 4'b0110;

	lut_sub lut_2031 ({i_9_, i_6_, g206}, g207);
	defparam lut_2031.LUT_SIZE = 3;
	defparam lut_2031.mask = 8'h08;

	lut_sub lut_2037 ({g28, g11}, g208);
	defparam lut_2037.LUT_SIZE = 2;
	defparam lut_2037.mask = 4'b0100;

	lut_sub lut_2043 ({g4, g138}, g209);
	defparam lut_2043.LUT_SIZE = 2;
	defparam lut_2043.mask = 4'b0100;

	lut_sub lut_2051 ({i_9_, g25, g18, g208, g209}, g210);
	defparam lut_2051.LUT_SIZE = 5;
	defparam lut_2051.mask = 32'h00550303;

	lut_sub lut_2064 ({g36, g3}, g211);
	defparam lut_2064.LUT_SIZE = 2;
	defparam lut_2064.mask = 4'b0010;

	lut_sub lut_2072 ({i_9_, g25, g45, g52, g211}, g212);
	defparam lut_2072.LUT_SIZE = 5;
	defparam lut_2072.mask = 32'h00553030;

	lut_sub lut_2087 ({i_5_, g39, g20, g92, g40}, g213);
	defparam lut_2087.LUT_SIZE = 5;
	defparam lut_2087.mask = 32'h00030011;

	lut_sub lut_2098 ({g207, g210, g212, g213}, g214);
	defparam lut_2098.LUT_SIZE = 4;
	defparam lut_2098.mask = 16'hc080;

	lut_sub lut_2108 ({g7, g204, g205, g214}, g215);
	defparam lut_2108.LUT_SIZE = 4;
	defparam lut_2108.mask = 16'h5040;

	lut_sub lut_2119 ({g192, g194, g196, g203, g215}, g216);
	defparam lut_2119.LUT_SIZE = 5;
	defparam lut_2119.mask = 32'h11001000;

	lut_sub lut_2131 ({g89, g108, g758, g114, g191, g216}, g217);
	defparam lut_2131.LUT_SIZE = 6;
	defparam lut_2131.mask = 64'h0000000000000001;

	lut_sub lut_2137 ({i_9_, i_8_, i_6_, i_7_, g29, g142}, g218);
	defparam lut_2137.LUT_SIZE = 6;
	defparam lut_2137.mask = 64'h000000000000300a;

	lut_sub lut_2148 ({g10, g1, g58, g218}, g219);
	defparam lut_2148.LUT_SIZE = 4;
	defparam lut_2148.mask = 16'h2aaa;

	lut_sub lut_2163 ({i_9_, g50, g124, g59, g134, g77}, g220);
	defparam lut_2163.LUT_SIZE = 6;
	defparam lut_2163.mask = 64'h0303030305ff0505;

	lut_sub lut_2190 ({g39, g28}, g221);
	defparam lut_2190.LUT_SIZE = 2;
	defparam lut_2190.mask = 4'b0010;

	lut_sub lut_2196 ({g76, g1}, g222);
	defparam lut_2196.LUT_SIZE = 2;
	defparam lut_2196.mask = 4'b1000;

	lut_sub lut_2205 ({g20, g42, g221, g135, g222}, g223);
	defparam lut_2205.LUT_SIZE = 5;
	defparam lut_2205.mask = 32'hffcca080;

	lut_sub lut_2225 ({g4, g11}, g224);
	defparam lut_2225.LUT_SIZE = 2;
	defparam lut_2225.mask = 4'b0100;

	lut_sub lut_2231 ({g50, g4}, g225);
	defparam lut_2231.LUT_SIZE = 2;
	defparam lut_2231.mask = 4'b1000;

	lut_sub lut_2239 ({g21, g27, g224, g225}, g226);
	defparam lut_2239.LUT_SIZE = 4;
	defparam lut_2239.mask = 16'h5703;

	lut_sub lut_2253 ({g219, g220, g223, g226}, g227);
	defparam lut_2253.LUT_SIZE = 4;
	defparam lut_2253.mask = 16'h0020;

	lut_sub lut_2259 ({g30, g45}, g228);
	defparam lut_2259.LUT_SIZE = 2;
	defparam lut_2259.mask = 4'b0010;

	lut_sub lut_2267 ({g35, g133, g165, g228}, g229);
	defparam lut_2267.LUT_SIZE = 4;
	defparam lut_2267.mask = 16'haf8c;

	lut_sub lut_2281 ({g8, g76}, g230);
	defparam lut_2281.LUT_SIZE = 2;
	defparam lut_2281.mask = 4'b0010;

	lut_sub lut_2290 ({g84, g1, g14, g40, g142}, g231);
	defparam lut_2290.LUT_SIZE = 5;
	defparam lut_2290.mask = 32'h32223333;

	lut_sub lut_2311 ({g42, g2, g186, g230, g231}, g232);
	defparam lut_2311.LUT_SIZE = 5;
	defparam lut_2311.mask = 32'haaa08880;

	lut_sub lut_2325 ({g30, g18}, g233);
	defparam lut_2325.LUT_SIZE = 2;
	defparam lut_2325.mask = 4'b0001;

	lut_sub lut_2334 ({g35, g28, g1, g40, g233}, g234);
	defparam lut_2334.LUT_SIZE = 5;
	defparam lut_2334.mask = 32'h30007555;

	lut_sub lut_2349 ({i_2_, i_0_, i_1_, g186}, g235);
	defparam lut_2349.LUT_SIZE = 4;
	defparam lut_2349.mask = 16'h3040;

	lut_sub lut_2361 ({g7, g6, g16, g4, g133, g53}, g236);
	defparam lut_2361.LUT_SIZE = 6;
	defparam lut_2361.mask = 64'h00c000c055d500c0;

	lut_sub lut_2383 ({i_2_, i_9_, g125, g234, g235, g236}, g237);
	defparam lut_2383.LUT_SIZE = 6;
	defparam lut_2383.mask = 64'ha080a0a08080a0a0;

	lut_sub lut_2403 ({i_9_, g50, g25, g60, g230}, g238);
	defparam lut_2403.LUT_SIZE = 5;
	defparam lut_2403.mask = 32'h05053300;

	lut_sub lut_2418 ({g49, g38, g182, g142}, g239);
	defparam lut_2418.LUT_SIZE = 4;
	defparam lut_2418.mask = 16'ha0b3;

	lut_sub lut_2430 ({g22, g30}, g240);
	defparam lut_2430.LUT_SIZE = 2;
	defparam lut_2430.mask = 4'b0001;

	lut_sub lut_2436 ({i_9_, i_8_, i_6_, i_7_, g26, g240}, g241);
	defparam lut_2436.LUT_SIZE = 6;
	defparam lut_2436.mask = 64'h0000000000050300;

	lut_sub lut_2446 ({g42, g233, g241}, g242);
	defparam lut_2446.LUT_SIZE = 3;
	defparam lut_2446.mask = 8'ha8;

	lut_sub lut_2457 ({g20, g28, g25, g137, g74}, g243);
	defparam lut_2457.LUT_SIZE = 5;
	defparam lut_2457.mask = 32'h0300abaa;

	lut_sub lut_2473 ({g10, g18}, g244);
	defparam lut_2473.LUT_SIZE = 2;
	defparam lut_2473.mask = 4'b0100;

	lut_sub lut_2482 ({g22, g38, g73, g4, g10}, g245);
	defparam lut_2482.LUT_SIZE = 5;
	defparam lut_2482.mask = 32'h0000ae0c;

	lut_sub lut_2495 ({g133, g244, g245}, g246);
	defparam lut_2495.LUT_SIZE = 3;
	defparam lut_2495.mask = 8'h8a;

	lut_sub lut_2507 ({g35, g42, g2, g161, g141, g244}, g247);
	defparam lut_2507.LUT_SIZE = 6;
	defparam lut_2507.mask = 64'hffaacc88f0a0c080;

	lut_sub lut_2542 ({g239, g242, g243, g246, g247}, g248);
	defparam lut_2542.LUT_SIZE = 5;
	defparam lut_2542.mask = 32'h00100000;

	lut_sub lut_2550 ({i_9_, g25, g3, g125, g62}, g249);
	defparam lut_2550.LUT_SIZE = 5;
	defparam lut_2550.mask = 32'h00335050;

	lut_sub lut_2565 ({g22, i_9_, g54, g122, g10}, g250);
	defparam lut_2565.LUT_SIZE = 5;
	defparam lut_2565.mask = 32'h0000a033;

	lut_sub lut_2576 ({g76, g18}, g251);
	defparam lut_2576.LUT_SIZE = 2;
	defparam lut_2576.mask = 4'b0100;

	lut_sub lut_2586 ({g42, g13, g43, g19, g165, g251}, g252);
	defparam lut_2586.LUT_SIZE = 6;
	defparam lut_2586.mask = 64'hc0ccf0ff8088a0aa;

	lut_sub lut_2621 ({g117, g133, g21, g161, g55}, g253);
	defparam lut_2621.LUT_SIZE = 5;
	defparam lut_2621.mask = 32'h8acf00cf;

	lut_sub lut_2644 ({g38, g73, g57, g1, g14}, g254);
	defparam lut_2644.LUT_SIZE = 5;
	defparam lut_2644.mask = 32'h888f000f;

	lut_sub lut_2663 ({g249, g250, g252, g253, g254}, g255);
	defparam lut_2663.LUT_SIZE = 5;
	defparam lut_2663.mask = 32'h02000000;

	lut_sub lut_2670 ({i_2_, i_0_, i_1_, g38, g30, g40}, g256);
	defparam lut_2670.LUT_SIZE = 6;
	defparam lut_2670.mask = 64'h1130001100000000;

	lut_sub lut_2682 ({i_2_, g119, g30, g10}, g257);
	defparam lut_2682.LUT_SIZE = 4;
	defparam lut_2682.mask = 16'h30a0;

	lut_sub lut_2694 ({g21, g58, g85, g141, g257}, g258);
	defparam lut_2694.LUT_SIZE = 5;
	defparam lut_2694.mask = 32'h80c0aaff;

	lut_sub lut_2714 ({g16, g14}, g259);
	defparam lut_2714.LUT_SIZE = 2;
	defparam lut_2714.mask = 4'b0010;

	lut_sub lut_2721 ({g49, g77, g259}, g260);
	defparam lut_2721.LUT_SIZE = 3;
	defparam lut_2721.mask = 8'h07;

	lut_sub lut_2732 ({g22, g38, g6, g76, g260}, g261);
	defparam lut_2732.LUT_SIZE = 5;
	defparam lut_2732.mask = 32'h2aaa22aa;

	lut_sub lut_2753 ({g133, g43, g169, g135, g211}, g262);
	defparam lut_2753.LUT_SIZE = 5;
	defparam lut_2753.mask = 32'h8088c0ff;

	lut_sub lut_2771 ({g10, g27}, g263);
	defparam lut_2771.LUT_SIZE = 2;
	defparam lut_2771.mask = 4'b0100;

	lut_sub lut_2779 ({i_9_, g25, g77, g209, g263}, g264);
	defparam lut_2779.LUT_SIZE = 5;
	defparam lut_2779.mask = 32'h005f0077;

	lut_sub lut_2799 ({i_9_, g39, g182, g44, g161, g251}, g265);
	defparam lut_2799.LUT_SIZE = 6;
	defparam lut_2799.mask = 64'h000055ff00003f3f;

	lut_sub lut_2831 ({g258, g261, g262, g264, g265}, g266);
	defparam lut_2831.LUT_SIZE = 5;
	defparam lut_2831.mask = 32'h00000008;

	lut_sub lut_2837 ({i_2_, g78, g180}, g267);
	defparam lut_2837.LUT_SIZE = 3;
	defparam lut_2837.mask = 8'he0;

	lut_sub lut_2848 ({g22, g42, g76, g27, g201}, g268);
	defparam lut_2848.LUT_SIZE = 5;
	defparam lut_2848.mask = 32'h00553075;

	lut_sub lut_2865 ({i_2_, i_9_, g8, g119, g10}, g269);
	defparam lut_2865.LUT_SIZE = 5;
	defparam lut_2865.mask = 32'hff000800;

	lut_sub lut_2881 ({g42, g124, g40, g15}, g270);
	defparam lut_2881.LUT_SIZE = 4;
	defparam lut_2881.mask = 16'h0357;

	lut_sub lut_2895 ({g22, i_9_, g36, g10, g18}, g271);
	defparam lut_2895.LUT_SIZE = 5;
	defparam lut_2895.mask = 32'h00004405;

	lut_sub lut_2902 ({i_0_, i_1_}, g272);
	defparam lut_2902.LUT_SIZE = 2;
	defparam lut_2902.mask = 4'b0100;

	lut_sub lut_2909 ({i_2_, i_9_, g272, g32, g141}, g273);
	defparam lut_2909.LUT_SIZE = 5;
	defparam lut_2909.mask = 32'h00030500;

	lut_sub lut_2919 ({i_2_, i_9_, g119, g31, g139}, g274);
	defparam lut_2919.LUT_SIZE = 5;
	defparam lut_2919.mask = 32'h50000030;

	lut_sub lut_2930 ({i_5_, g92, g11, g137, g1}, g275);
	defparam lut_2930.LUT_SIZE = 5;
	defparam lut_2930.mask = 32'h00030023;

	lut_sub lut_2942 ({g271, g273, g274, g275}, g276);
	defparam lut_2942.LUT_SIZE = 4;
	defparam lut_2942.mask = 16'h8000;

	lut_sub lut_2951 ({g267, g268, g269, g270, g276}, g277);
	defparam lut_2951.LUT_SIZE = 5;
	defparam lut_2951.mask = 32'h40004400;

	lut_sub lut_2963 ({g238, g248, g255, g256, g266, g277}, g278);
	defparam lut_2963.LUT_SIZE = 6;
	defparam lut_2963.mask = 64'h0000001000000000;

	lut_sub lut_2971 ({g43, g21, g51, g157}, g279);
	defparam lut_2971.LUT_SIZE = 4;
	defparam lut_2971.mask = 16'h7530;

	lut_sub lut_2986 ({g20, g122, g43, g179, g60}, g280);
	defparam lut_2986.LUT_SIZE = 5;
	defparam lut_2986.mask = 32'hcf0f8a0a;

	lut_sub lut_3008 ({g57, g137, g2, g201}, g281);
	defparam lut_3008.LUT_SIZE = 4;
	defparam lut_3008.mask = 16'h111f;

	lut_sub lut_3021 ({g38, g175, g26}, g282);
	defparam lut_3021.LUT_SIZE = 3;
	defparam lut_3021.mask = 8'h8c;

	lut_sub lut_3032 ({g73, g43, g64, g85, g240}, g283);
	defparam lut_3032.LUT_SIZE = 5;
	defparam lut_3032.mask = 32'hccff80a0;

	lut_sub lut_3054 ({i_9_, g50, g28, g63, g45}, g284);
	defparam lut_3054.LUT_SIZE = 5;
	defparam lut_3054.mask = 32'h20203000;

	lut_sub lut_3064 ({i_2_, i_0_, i_1_, g7, g36, g40}, g285);
	defparam lut_3064.LUT_SIZE = 6;
	defparam lut_3064.mask = 64'h0000001105000005;

	lut_sub lut_3078 ({g54, g10, g133, g284, g285}, g286);
	defparam lut_3078.LUT_SIZE = 5;
	defparam lut_3078.mask = 32'h08888888;

	lut_sub lut_3093 ({g21, g158, g282, g283, g286}, g287);
	defparam lut_3093.LUT_SIZE = 5;
	defparam lut_3093.mask = 32'h01000101;

	lut_sub lut_3102 ({i_2_, g78, i_9_, g117, g230}, g288);
	defparam lut_3102.LUT_SIZE = 5;
	defparam lut_3102.mask = 32'h00500030;

	lut_sub lut_3114 ({g76, g1, g40, g150, g288}, g289);
	defparam lut_3114.LUT_SIZE = 5;
	defparam lut_3114.mask = 32'h80888888;

	lut_sub lut_3129 ({g279, g729, g281, g287, g289}, g290);
	defparam lut_3129.LUT_SIZE = 5;
	defparam lut_3129.mask = 32'h00100000;

	lut_sub lut_3135 ({i_9_, i_5_, i_3_, i_4_, g3, g45}, g291);
	defparam lut_3135.LUT_SIZE = 6;
	defparam lut_3135.mask = 64'h000000a000c00000;

	lut_sub lut_3144 ({i_0_, i_1_, g9, g46}, g292);
	defparam lut_3144.LUT_SIZE = 4;
	defparam lut_3144.mask = 16'h0250;

	lut_sub lut_3154 ({i_2_, i_9_, g119, g125, g117, g292}, g293);
	defparam lut_3154.LUT_SIZE = 6;
	defparam lut_3154.mask = 64'h0f00000077550000;

	lut_sub lut_3174 ({g73, g23, g293}, g294);
	defparam lut_3174.LUT_SIZE = 3;
	defparam lut_3174.mask = 8'ha8;

	lut_sub lut_3185 ({g35, g28, g2, g18, g225}, g295);
	defparam lut_3185.LUT_SIZE = 5;
	defparam lut_3185.mask = 32'h05053705;

	lut_sub lut_3203 ({g181, g70, g295, g189}, g296);
	defparam lut_3203.LUT_SIZE = 4;
	defparam lut_3203.mask = 16'h4000;

	lut_sub lut_3213 ({g59, g290, g722, g291, g294, g296}, g297);
	defparam lut_3213.LUT_SIZE = 6;
	defparam lut_3213.mask = 64'h0000001100000010;

	lut_sub lut_3225 ({g227, g735, g232, g237, g278, g297}, g298);
	defparam lut_3225.LUT_SIZE = 6;
	defparam lut_3225.mask = 64'h0000000000000001;

	lut_sub lut_3233 ({g22, i_9_, g25, g134, g171}, g299);
	defparam lut_3233.LUT_SIZE = 5;
	defparam lut_3233.mask = 32'h03000355;

	lut_sub lut_3249 ({g22, g73, g30, g11, g137}, g300);
	defparam lut_3249.LUT_SIZE = 5;
	defparam lut_3249.mask = 32'h0101010f;

	lut_sub lut_3263 ({g20, g6, g10, g300}, g301);
	defparam lut_3263.LUT_SIZE = 4;
	defparam lut_3263.mask = 16'haa2a;

	lut_sub lut_3275 ({g6, g76}, g302);
	defparam lut_3275.LUT_SIZE = 2;
	defparam lut_3275.mask = 4'b1000;

	lut_sub lut_3284 ({g28, g42, g63, g40, g139}, g303);
	defparam lut_3284.LUT_SIZE = 5;
	defparam lut_3284.mask = 32'h03570055;

	lut_sub lut_3301 ({g27, g302, g303}, g304);
	defparam lut_3301.LUT_SIZE = 3;
	defparam lut_3301.mask = 8'ha8;

	lut_sub lut_3311 ({i_9_, g50, g7, g6, g62}, g305);
	defparam lut_3311.LUT_SIZE = 5;
	defparam lut_3311.mask = 32'h0c005500;

	lut_sub lut_3323 ({g49, g28, g18}, g306);
	defparam lut_3323.LUT_SIZE = 3;
	defparam lut_3323.mask = 8'h04;

	lut_sub lut_3329 ({g76, g59}, g307);
	defparam lut_3329.LUT_SIZE = 2;
	defparam lut_3329.mask = 4'b0100;

	lut_sub lut_3338 ({g22, g10, g53, g306, g307}, g308);
	defparam lut_3338.LUT_SIZE = 5;
	defparam lut_3338.mask = 32'hc8c8c0c8;

	lut_sub lut_3357 ({g49, g1, g183, g14, g40}, g309);
	defparam lut_3357.LUT_SIZE = 5;
	defparam lut_3357.mask = 32'h44004f0f;

	lut_sub lut_3376 ({g22, g38, g36, g39, g58}, g310);
	defparam lut_3376.LUT_SIZE = 5;
	defparam lut_3376.mask = 32'h03000b0a;

	lut_sub lut_3389 ({g35, g170, g310}, g311);
	defparam lut_3389.LUT_SIZE = 3;
	defparam lut_3389.mask = 8'ha8;

	lut_sub lut_3400 ({g49, g141, g308, g309, g311}, g312);
	defparam lut_3400.LUT_SIZE = 5;
	defparam lut_3400.mask = 32'h04040400;

	lut_sub lut_3411 ({g76, g3, g13, g305, g312}, g313);
	defparam lut_3411.LUT_SIZE = 5;
	defparam lut_3411.mask = 32'h04444444;

	lut_sub lut_3426 ({g234, g299, g301, g304, g313}, g314);
	defparam lut_3426.LUT_SIZE = 5;
	defparam lut_3426.mask = 32'h01000000;

	lut_sub lut_3434 ({i_9_, g39, g3, g55, g302}, g315);
	defparam lut_3434.LUT_SIZE = 5;
	defparam lut_3434.mask = 32'h00335050;

	lut_sub lut_3450 ({g73, g133, g64, g19, g208}, g316);
	defparam lut_3450.LUT_SIZE = 5;
	defparam lut_3450.mask = 32'hccff80a0;

	lut_sub lut_3472 ({g2, g251, g315, g316}, g317);
	defparam lut_3472.LUT_SIZE = 4;
	defparam lut_3472.mask = 16'h4440;

	lut_sub lut_3482 ({g38, g94, g58, g23}, g318);
	defparam lut_3482.LUT_SIZE = 4;
	defparam lut_3482.mask = 16'h4f44;

	lut_sub lut_3497 ({g28, g73, g63, g13, g18}, g319);
	defparam lut_3497.LUT_SIZE = 5;
	defparam lut_3497.mask = 32'h444f0000;

	lut_sub lut_3511 ({g73, g26, g318, g319}, g320);
	defparam lut_3511.LUT_SIZE = 4;
	defparam lut_3511.mask = 16'h8880;

	lut_sub lut_3521 ({g7, g20, g6, g320}, g321);
	defparam lut_3521.LUT_SIZE = 4;
	defparam lut_3521.mask = 16'h5551;

	lut_sub lut_3535 ({i_9_, g6, g45, g94, g171}, g322);
	defparam lut_3535.LUT_SIZE = 5;
	defparam lut_3535.mask = 32'h55003030;

	lut_sub lut_3552 ({g73, g57, g94, g58, g82, g195}, g323);
	defparam lut_3552.LUT_SIZE = 6;
	defparam lut_3552.mask = 64'hffff0f0f88000800;

	lut_sub lut_3586 ({g49, g35, g170, g228}, g324);
	defparam lut_3586.LUT_SIZE = 4;
	defparam lut_3586.mask = 16'h0537;

	lut_sub lut_3601 ({g53, g112, g322, g323, g324}, g325);
	defparam lut_3601.LUT_SIZE = 5;
	defparam lut_3601.mask = 32'h20202000;

	lut_sub lut_3612 ({g7, g35, g16, g2, g225}, g326);
	defparam lut_3612.LUT_SIZE = 5;
	defparam lut_3612.mask = 32'h00550757;

	lut_sub lut_3630 ({i_9_, g50, g7, g31}, g327);
	defparam lut_3630.LUT_SIZE = 4;
	defparam lut_3630.mask = 16'h3055;

	lut_sub lut_3644 ({g59, g131, g325, g326, g327}, g328);
	defparam lut_3644.LUT_SIZE = 5;
	defparam lut_3644.mask = 32'h0f0c0a08;

	lut_sub lut_3659 ({g22, i_5_, i_3_, i_4_, g20, g207}, g329);
	defparam lut_3659.LUT_SIZE = 6;
	defparam lut_3659.mask = 64'h0000000051000000;

	lut_sub lut_3669 ({i_2_, g272, g168, g79, g97}, g330);
	defparam lut_3669.LUT_SIZE = 5;
	defparam lut_3669.mask = 32'h00031111;

	lut_sub lut_3678 ({i_9_, i_8_, i_6_, i_7_}, g331);
	defparam lut_3678.LUT_SIZE = 4;
	defparam lut_3678.mask = 16'h0060;

	lut_sub lut_3688 ({g38, g137, g64, g195, g331}, g332);
	defparam lut_3688.LUT_SIZE = 5;
	defparam lut_3688.mask = 32'h11150105;

	lut_sub lut_3703 ({i_9_, g50, g36, g6, g170}, g333);
	defparam lut_3703.LUT_SIZE = 5;
	defparam lut_3703.mask = 32'h44440c00;

	lut_sub lut_3716 ({g21, g60, g27, g171}, g334);
	defparam lut_3716.LUT_SIZE = 4;
	defparam lut_3716.mask = 16'h5703;

	lut_sub lut_3731 ({g40, g195, g332, g333, g334}, g335);
	defparam lut_3731.LUT_SIZE = 5;
	defparam lut_3731.mask = 32'h80808000;

	lut_sub lut_3742 ({g28, g40, g329, g330, g335}, g336);
	defparam lut_3742.LUT_SIZE = 5;
	defparam lut_3742.mask = 32'h40404440;

	lut_sub lut_3754 ({i_9_, g39, g30, g44, g58}, g337);
	defparam lut_3754.LUT_SIZE = 5;
	defparam lut_3754.mask = 32'h003b000a;

	lut_sub lut_3770 ({g49, g53, g82, g19, g230, g337}, g338);
	defparam lut_3770.LUT_SIZE = 6;
	defparam lut_3770.mask = 64'haaaaaa0080808000;

	lut_sub lut_3793 ({g22, i_9_, g28, g84, g45, g177}, g339);
	defparam lut_3793.LUT_SIZE = 6;
	defparam lut_3793.mask = 64'h00000c0ccc005d5d;

	lut_sub lut_3817 ({g30, g11, g58}, g340);
	defparam lut_3817.LUT_SIZE = 3;
	defparam lut_3817.mask = 8'h02;

	lut_sub lut_3826 ({g39, g10, g53, g144, g340}, g341);
	defparam lut_3826.LUT_SIZE = 5;
	defparam lut_3826.mask = 32'ha8a8a0a8;

	lut_sub lut_3846 ({g116, g59, g10, g43, g137, g259}, g342);
	defparam lut_3846.LUT_SIZE = 6;
	defparam lut_3846.mask = 64'h505073505050ffff;

	lut_sub lut_3885 ({g49, i_6_, g36, g39, g73, g206}, g343);
	defparam lut_3885.LUT_SIZE = 6;
	defparam lut_3885.mask = 64'h00030003000300ab;

	lut_sub lut_3899 ({i_9_, i_8_, i_6_, i_7_, i_5_}, g344);
	defparam lut_3899.LUT_SIZE = 5;
	defparam lut_3899.mask = 32'h00008004;

	lut_sub lut_3906 ({i_3_, i_4_, g63, g344}, g345);
	defparam lut_3906.LUT_SIZE = 4;
	defparam lut_3906.mask = 16'h1000;

	lut_sub lut_3914 ({i_6_, g76, g9, g133, g206}, g346);
	defparam lut_3914.LUT_SIZE = 5;
	defparam lut_3914.mask = 32'h8c0c0c0c;

	lut_sub lut_3930 ({g38, g28, g10, g1}, g347);
	defparam lut_3930.LUT_SIZE = 4;
	defparam lut_3930.mask = 16'ha800;

	lut_sub lut_3941 ({g35, g169, g345, g346, g347}, g348);
	defparam lut_3941.LUT_SIZE = 5;
	defparam lut_3941.mask = 32'h80808000;

	lut_sub lut_3952 ({g339, g341, g342, g343, g348}, g349);
	defparam lut_3952.LUT_SIZE = 5;
	defparam lut_3952.mask = 32'h00400000;

	lut_sub lut_3956 ({i_6_, i_7_, i_5_, i_3_}, g350);
	defparam lut_3956.LUT_SIZE = 4;
	defparam lut_3956.mask = 16'h4000;

	lut_sub lut_3962 ({g22, i_9_, i_8_, i_4_, g350}, g351);
	defparam lut_3962.LUT_SIZE = 5;
	defparam lut_3962.mask = 32'h00000014;

	lut_sub lut_3968 ({i_2_, i_9_, i_7_, g272}, g352);
	defparam lut_3968.LUT_SIZE = 4;
	defparam lut_3968.mask = 16'h1040;

	lut_sub lut_3975 ({i_8_, i_6_, g4, g352}, g353);
	defparam lut_3975.LUT_SIZE = 4;
	defparam lut_3975.mask = 16'h0004;

	lut_sub lut_3981 ({g7, g25}, g354);
	defparam lut_3981.LUT_SIZE = 2;
	defparam lut_3981.mask = 4'b0001;

	lut_sub lut_3988 ({i_9_, i_8_, g83, g82, g354}, g355);
	defparam lut_3988.LUT_SIZE = 5;
	defparam lut_3988.mask = 32'h00000503;

	lut_sub lut_3997 ({g10, g138}, g356);
	defparam lut_3997.LUT_SIZE = 2;
	defparam lut_3997.mask = 4'b0100;

	lut_sub lut_4005 ({i_2_, g119, g157, g151, g356}, g357);
	defparam lut_4005.LUT_SIZE = 5;
	defparam lut_4005.mask = 32'h11000303;

	lut_sub lut_4014 ({i_2_, i_9_, i_8_, i_6_, i_7_}, g358);
	defparam lut_4014.LUT_SIZE = 5;
	defparam lut_4014.mask = 32'hfffdffef;

	lut_sub lut_4050 ({g38, g28, g59}, g359);
	defparam lut_4050.LUT_SIZE = 3;
	defparam lut_4050.mask = 8'h40;

	lut_sub lut_4059 ({g40, g27, g142, g90, g359}, g360);
	defparam lut_4059.LUT_SIZE = 5;
	defparam lut_4059.mask = 32'haa0a8808;

	lut_sub lut_4076 ({g20, g307, g357, g711, g360}, g361);
	defparam lut_4076.LUT_SIZE = 5;
	defparam lut_4076.mask = 32'h10101000;

	lut_sub lut_4087 ({g56, g351, g353, g355, g361}, g362);
	defparam lut_4087.LUT_SIZE = 5;
	defparam lut_4087.mask = 32'h40000000;

	lut_sub lut_4097 ({g729, g248, g336, g338, g349, g362}, g363);
	defparam lut_4097.LUT_SIZE = 6;
	defparam lut_4097.mask = 64'h0000000000000001;

	lut_sub lut_4107 ({g108, g314, g317, g321, g328, g363}, g364);
	defparam lut_4107.LUT_SIZE = 6;
	defparam lut_4107.mask = 64'h0000000000000001;

	lut_sub lut_4116 ({g35, g76, g1, g40, g201}, g365);
	defparam lut_4116.LUT_SIZE = 5;
	defparam lut_4116.mask = 32'h30007555;

	lut_sub lut_4133 ({i_9_, g116, g63, g161}, g366);
	defparam lut_4133.LUT_SIZE = 4;
	defparam lut_4133.mask = 16'h1103;

	lut_sub lut_4144 ({g133, g64, g27, g165}, g367);
	defparam lut_4144.LUT_SIZE = 4;
	defparam lut_4144.mask = 16'h5703;

	lut_sub lut_4158 ({g38, g307, g354, g367}, g368);
	defparam lut_4158.LUT_SIZE = 4;
	defparam lut_4158.mask = 16'h80aa;

	lut_sub lut_4172 ({g35, g43, g169, g58, g71, g171}, g369);
	defparam lut_4172.LUT_SIZE = 6;
	defparam lut_4172.mask = 64'hcf00cfcf8a008a8a;

	lut_sub lut_4207 ({g8, g36, g42, g13, g183}, g370);
	defparam lut_4207.LUT_SIZE = 5;
	defparam lut_4207.mask = 32'h050505cd;

	lut_sub lut_4226 ({g365, g366, g368, g369, g370}, g371);
	defparam lut_4226.LUT_SIZE = 5;
	defparam lut_4226.mask = 32'h02000000;

	lut_sub lut_4234 ({g59, g10, g58, g371}, g372);
	defparam lut_4234.LUT_SIZE = 4;
	defparam lut_4234.mask = 16'h5515;

	lut_sub lut_4249 ({g49, g7, g3, g21, g156}, g373);
	defparam lut_4249.LUT_SIZE = 5;
	defparam lut_4249.mask = 32'h445444f4;

	lut_sub lut_4267 ({i_9_, g39, g101, g31}, g374);
	defparam lut_4267.LUT_SIZE = 4;
	defparam lut_4267.mask = 16'h0503;

	lut_sub lut_4277 ({g43, g37, g55}, g375);
	defparam lut_4277.LUT_SIZE = 3;
	defparam lut_4277.mask = 8'hd0;

	lut_sub lut_4288 ({g76, g73, g11, g90, g375}, g376);
	defparam lut_4288.LUT_SIZE = 5;
	defparam lut_4288.mask = 32'haa80aa88;

	lut_sub lut_4307 ({g20, g28, g25, g10, g137}, g377);
	defparam lut_4307.LUT_SIZE = 5;
	defparam lut_4307.mask = 32'h04040f04;

	lut_sub lut_4320 ({g35, g165, g377}, g378);
	defparam lut_4320.LUT_SIZE = 3;
	defparam lut_4320.mask = 8'ha8;

	lut_sub lut_4329 ({g2, g77, g115}, g379);
	defparam lut_4329.LUT_SIZE = 3;
	defparam lut_4329.mask = 8'ha8;

	lut_sub lut_4340 ({g24, g374, g376, g378, g379}, g380);
	defparam lut_4340.LUT_SIZE = 5;
	defparam lut_4340.mask = 32'h01000000;

	lut_sub lut_4346 ({i_2_, i_0_, i_9_, g373, g380}, g381);
	defparam lut_4346.LUT_SIZE = 5;
	defparam lut_4346.mask = 32'h55555545;

	lut_sub lut_4368 ({i_9_, g7, g25, g16, g157}, g382);
	defparam lut_4368.LUT_SIZE = 5;
	defparam lut_4368.mask = 32'h00030505;

	lut_sub lut_4382 ({g42, g21, g32, g135, g244}, g383);
	defparam lut_4382.LUT_SIZE = 5;
	defparam lut_4382.mask = 32'hf0ff8088;

	lut_sub lut_4405 ({i_9_, g16, g124, g59, g1, g14}, g384);
	defparam lut_4405.LUT_SIZE = 6;
	defparam lut_4405.mask = 64'h00000a0a000088ff;

	lut_sub lut_4427 ({g22, g7, g221, g14, g53}, g385);
	defparam lut_4427.LUT_SIZE = 5;
	defparam lut_4427.mask = 32'h05054555;

	lut_sub lut_4444 ({i_9_, i_8_, g68, g28, g63}, g386);
	defparam lut_4444.LUT_SIZE = 5;
	defparam lut_4444.mask = 32'h04000004;

	lut_sub lut_4453 ({g20, g84, g62, g386}, g387);
	defparam lut_4453.LUT_SIZE = 4;
	defparam lut_4453.mask = 16'haa80;

	lut_sub lut_4467 ({g49, g117, g134, g2, g179, g171}, g388);
	defparam lut_4467.LUT_SIZE = 6;
	defparam lut_4467.mask = 64'hfaf0f0f0c8c0c0c0;

	lut_sub lut_4502 ({g22, g20, g10, g40, g307}, g389);
	defparam lut_4502.LUT_SIZE = 5;
	defparam lut_4502.mask = 32'h111111f1;

	lut_sub lut_4519 ({g40, g144, g389}, g390);
	defparam lut_4519.LUT_SIZE = 3;
	defparam lut_4519.mask = 8'ha8;

	lut_sub lut_4531 ({g383, g384, g385, g387, g388, g390}, g391);
	defparam lut_4531.LUT_SIZE = 6;
	defparam lut_4531.mask = 64'h0000000001000000;

	lut_sub lut_4538 ({g133, g5, g80}, g392);
	defparam lut_4538.LUT_SIZE = 3;
	defparam lut_4538.mask = 8'h8a;

	lut_sub lut_4546 ({i_2_, i_0_, i_1_, g4, g137}, g393);
	defparam lut_4546.LUT_SIZE = 5;
	defparam lut_4546.mask = 32'hc0000040;

	lut_sub lut_4553 ({i_9_, i_8_, i_6_, g393}, g394);
	defparam lut_4553.LUT_SIZE = 4;
	defparam lut_4553.mask = 16'h0040;

	lut_sub lut_4562 ({g7, g38, g39, g43, g156}, g395);
	defparam lut_4562.LUT_SIZE = 5;
	defparam lut_4562.mask = 32'h44444f44;

	lut_sub lut_4580 ({g28, g2, g18, g395}, g396);
	defparam lut_4580.LUT_SIZE = 4;
	defparam lut_4580.mask = 16'ha8aa;

	lut_sub lut_4594 ({g25, g40, g394, g396}, g397);
	defparam lut_4594.LUT_SIZE = 4;
	defparam lut_4594.mask = 16'h5444;

	lut_sub lut_4606 ({i_9_, g54, g45, g60, g240}, g398);
	defparam lut_4606.LUT_SIZE = 5;
	defparam lut_4606.mask = 32'h33005050;

	lut_sub lut_4621 ({g22, i_9_, g50, g76, g156}, g399);
	defparam lut_4621.LUT_SIZE = 5;
	defparam lut_4621.mask = 32'h000055c0;

	lut_sub lut_4634 ({i_9_, g6, g3, g30, g179}, g400);
	defparam lut_4634.LUT_SIZE = 5;
	defparam lut_4634.mask = 32'h55003000;

	lut_sub lut_4645 ({i_2_, i_9_, g7, g16}, g401);
	defparam lut_4645.LUT_SIZE = 4;
	defparam lut_4645.mask = 16'h5051;

	lut_sub lut_4656 ({i_2_, i_9_, g119, g10, g401}, g402);
	defparam lut_4656.LUT_SIZE = 5;
	defparam lut_4656.mask = 32'h40500050;

	lut_sub lut_4667 ({g28, g18, g21}, g403);
	defparam lut_4667.LUT_SIZE = 3;
	defparam lut_4667.mask = 8'h20;

	lut_sub lut_4676 ({g133, g53, g46, g224, g403}, g404);
	defparam lut_4676.LUT_SIZE = 5;
	defparam lut_4676.mask = 32'ha080aa88;

	lut_sub lut_4693 ({g398, g399, g400, g402, g404}, g405);
	defparam lut_4693.LUT_SIZE = 5;
	defparam lut_4693.mask = 32'h40000000;

	lut_sub lut_4701 ({i_9_, g25, g5, g148, g405}, g406);
	defparam lut_4701.LUT_SIZE = 5;
	defparam lut_4701.mask = 32'h55445550;

	lut_sub lut_4719 ({i_9_, g59, g37, g19}, g407);
	defparam lut_4719.LUT_SIZE = 4;
	defparam lut_4719.mask = 16'h0c05;

	lut_sub lut_4730 ({i_9_, g39, g76, g3, g209}, g408);
	defparam lut_4730.LUT_SIZE = 5;
	defparam lut_4730.mask = 32'h00c00055;

	lut_sub lut_4742 ({i_9_, i_5_, g6, g45, g11}, g409);
	defparam lut_4742.LUT_SIZE = 5;
	defparam lut_4742.mask = 32'hc0000044;

	lut_sub lut_4752 ({i_3_, i_4_, g407, g408, g409}, g410);
	defparam lut_4752.LUT_SIZE = 5;
	defparam lut_4752.mask = 32'hc0c080c0;

	lut_sub lut_4765 ({i_2_, i_9_, g119, g233, g259}, g411);
	defparam lut_4765.LUT_SIZE = 5;
	defparam lut_4765.mask = 32'h50000030;

	lut_sub lut_4777 ({g7, g63, g13, g27, g193}, g412);
	defparam lut_4777.LUT_SIZE = 5;
	defparam lut_4777.mask = 32'h50505073;

	lut_sub lut_4796 ({g22, g28, g2, g177, g58}, g413);
	defparam lut_4796.LUT_SIZE = 5;
	defparam lut_4796.mask = 32'h0303ab03;

	lut_sub lut_4815 ({g35, g85, g411, g412, g413}, g414);
	defparam lut_4815.LUT_SIZE = 5;
	defparam lut_4815.mask = 32'h80808000;

	lut_sub lut_4825 ({i_8_, g7, g36, g63, g69}, g415);
	defparam lut_4825.LUT_SIZE = 5;
	defparam lut_4825.mask = 32'h00110101;

	lut_sub lut_4836 ({i_9_, g39, g76, g16, g4}, g416);
	defparam lut_4836.LUT_SIZE = 5;
	defparam lut_4836.mask = 32'h00300022;

	lut_sub lut_4847 ({g42, g193, g415, g416}, g417);
	defparam lut_4847.LUT_SIZE = 4;
	defparam lut_4847.mask = 16'h8880;

	lut_sub lut_4858 ({g22, i_9_, g3, g63, g10, g31}, g418);
	defparam lut_4858.LUT_SIZE = 6;
	defparam lut_4858.mask = 64'h0c000c005d550c00;

	lut_sub lut_4879 ({i_9_, i_6_, g39, g30, g206}, g419);
	defparam lut_4879.LUT_SIZE = 5;
	defparam lut_4879.mask = 32'h00000001;

	lut_sub lut_4888 ({g20, g13, g161, g112, g208}, g420);
	defparam lut_4888.LUT_SIZE = 5;
	defparam lut_4888.mask = 32'hf0ff8088;

	lut_sub lut_4911 ({g38, g35, g120, g9, g57}, g421);
	defparam lut_4911.LUT_SIZE = 5;
	defparam lut_4911.mask = 32'haa80ffc0;

	lut_sub lut_4933 ({g76, g3, g4, g45}, g422);
	defparam lut_4933.LUT_SIZE = 4;
	defparam lut_4933.mask = 16'hf888;

	lut_sub lut_4947 ({g122, g2, g15, g422}, g423);
	defparam lut_4947.LUT_SIZE = 4;
	defparam lut_4947.mask = 16'h070f;

	lut_sub lut_4957 ({i_9_, i_8_, i_7_}, g424);
	defparam lut_4957.LUT_SIZE = 3;
	defparam lut_4957.mask = 8'h01;

	lut_sub lut_4963 ({i_6_, i_5_, i_3_, i_4_, g25, g424}, g425);
	defparam lut_4963.LUT_SIZE = 6;
	defparam lut_4963.mask = 64'h1000000000001000;

	lut_sub lut_4971 ({i_5_, i_3_, i_4_, g39, g59, g40}, g426);
	defparam lut_4971.LUT_SIZE = 6;
	defparam lut_4971.mask = 64'h0505000000110000;

	lut_sub lut_4985 ({g26, g27, g354, g425, g426}, g427);
	defparam lut_4985.LUT_SIZE = 5;
	defparam lut_4985.mask = 32'h88808800;

	lut_sub lut_4998 ({g419, g420, g421, g423, g427}, g428);
	defparam lut_4998.LUT_SIZE = 5;
	defparam lut_4998.mask = 32'h00040000;

	lut_sub lut_5007 ({g255, g414, g417, g418, g428}, g429);
	defparam lut_5007.LUT_SIZE = 5;
	defparam lut_5007.mask = 32'h00000004;

	lut_sub lut_5017 ({g392, g203, g397, g406, g410, g429}, g430);
	defparam lut_5017.LUT_SIZE = 6;
	defparam lut_5017.mask = 64'h0000000000000001;

	lut_sub lut_5027 ({g314, g372, g381, g382, g391, g430}, g431);
	defparam lut_5027.LUT_SIZE = 6;
	defparam lut_5027.mask = 64'h0000000000000010;

	lut_sub lut_5034 ({i_2_, i_9_, g272, g157, g233}, g432);
	defparam lut_5034.LUT_SIZE = 5;
	defparam lut_5034.mask = 32'h03000005;

	lut_sub lut_5045 ({i_9_, g50, g7, g6, g221}, g433);
	defparam lut_5045.LUT_SIZE = 5;
	defparam lut_5045.mask = 32'h0c005500;

	lut_sub lut_5058 ({g20, g240, g432, g433}, g434);
	defparam lut_5058.LUT_SIZE = 4;
	defparam lut_5058.mask = 16'h8880;

	lut_sub lut_5069 ({i_9_, g8, g28, g63, g11, g138}, g435);
	defparam lut_5069.LUT_SIZE = 6;
	defparam lut_5069.mask = 64'h0500050000003300;

	lut_sub lut_5084 ({i_2_, g78, g156, g31, g151}, g436);
	defparam lut_5084.LUT_SIZE = 5;
	defparam lut_5084.mask = 32'h00051111;

	lut_sub lut_5098 ({g22, i_9_, g9, g11, g165, g193}, g437);
	defparam lut_5098.LUT_SIZE = 6;
	defparam lut_5098.mask = 64'h0505030305ff5757;

	lut_sub lut_5132 ({i_9_, g25, g44, g31}, g438);
	defparam lut_5132.LUT_SIZE = 4;
	defparam lut_5132.mask = 16'h0305;

	lut_sub lut_5143 ({i_9_, g54, g59, g10, g31}, g439);
	defparam lut_5143.LUT_SIZE = 5;
	defparam lut_5143.mask = 32'h05050c00;

	lut_sub lut_5154 ({g25, g76}, g440);
	defparam lut_5154.LUT_SIZE = 2;
	defparam lut_5154.mask = 4'b0010;

	lut_sub lut_5164 ({g20, g53, g27, g12, g208, g440}, g441);
	defparam lut_5164.LUT_SIZE = 6;
	defparam lut_5164.mask = 64'hff0a88080f0a0808;

	lut_sub lut_5192 ({g7, g42, g3, g356}, g442);
	defparam lut_5192.LUT_SIZE = 4;
	defparam lut_5192.mask = 16'h050d;

	lut_sub lut_5203 ({g120, g4, g45}, g443);
	defparam lut_5203.LUT_SIZE = 3;
	defparam lut_5203.mask = 8'h70;

	lut_sub lut_5214 ({g13, g161, g51, g442, g443}, g444);
	defparam lut_5214.LUT_SIZE = 5;
	defparam lut_5214.mask = 32'h4000cccc;

	lut_sub lut_5228 ({g49, i_5_, i_3_, i_4_, g3}, g445);
	defparam lut_5228.LUT_SIZE = 5;
	defparam lut_5228.mask = 32'h00002280;

	lut_sub lut_5238 ({g35, g5, g230, g445}, g446);
	defparam lut_5238.LUT_SIZE = 4;
	defparam lut_5238.mask = 16'haa80;

	lut_sub lut_5249 ({i_5_, i_4_, g8, g117, g133}, g447);
	defparam lut_5249.LUT_SIZE = 5;
	defparam lut_5249.mask = 32'h222a2222;

	lut_sub lut_5266 ({g22, g28, g73, g27, g90}, g448);
	defparam lut_5266.LUT_SIZE = 5;
	defparam lut_5266.mask = 32'h15151f15;

	lut_sub lut_5288 ({g63, g263, g446, g447, g448}, g449);
	defparam lut_5288.LUT_SIZE = 5;
	defparam lut_5288.mask = 32'h08080800;

	lut_sub lut_5299 ({g438, g439, g441, g444, g449}, g450);
	defparam lut_5299.LUT_SIZE = 5;
	defparam lut_5299.mask = 32'h01000000;

	lut_sub lut_5304 ({i_9_, i_3_, i_4_, g1}, g451);
	defparam lut_5304.LUT_SIZE = 4;
	defparam lut_5304.mask = 16'h0280;

	lut_sub lut_5313 ({i_9_, g63, g11, g51, g32}, g452);
	defparam lut_5313.LUT_SIZE = 5;
	defparam lut_5313.mask = 32'h03030055;

	lut_sub lut_5330 ({g2, g21, g40, g64, g15, g165}, g453);
	defparam lut_5330.LUT_SIZE = 6;
	defparam lut_5330.mask = 64'hccc0fff08880aaa0;

	lut_sub lut_5365 ({g7, g39, g42, g58, g209}, g454);
	defparam lut_5365.LUT_SIZE = 5;
	defparam lut_5365.mask = 32'h050505cd;

	lut_sub lut_5384 ({g137, g302, g452, g453, g454}, g455);
	defparam lut_5384.LUT_SIZE = 5;
	defparam lut_5384.mask = 32'h20202000;

	lut_sub lut_5395 ({i_5_, g54, g308, g389, g451, g455}, g456);
	defparam lut_5395.LUT_SIZE = 6;
	defparam lut_5395.mask = 64'h0040005000500050;

	lut_sub lut_5409 ({g73, g124, g133, g97}, g457);
	defparam lut_5409.LUT_SIZE = 4;
	defparam lut_5409.mask = 16'h444f;

	lut_sub lut_5419 ({i_9_, i_8_, i_6_, i_7_}, g458);
	defparam lut_5419.LUT_SIZE = 4;
	defparam lut_5419.mask = 16'h0090;

	lut_sub lut_5426 ({i_5_, i_3_, i_4_, g11, g40}, g459);
	defparam lut_5426.LUT_SIZE = 5;
	defparam lut_5426.mask = 32'h30010000;

	lut_sub lut_5436 ({g4, g53, g458, g459}, g460);
	defparam lut_5436.LUT_SIZE = 4;
	defparam lut_5436.mask = 16'h1101;

	lut_sub lut_5446 ({g9, g21, g169, g32}, g461);
	defparam lut_5446.LUT_SIZE = 4;
	defparam lut_5446.mask = 16'h70f0;

	lut_sub lut_5462 ({g35, g120, g43, g2, g85, g186}, g462);
	defparam lut_5462.LUT_SIZE = 6;
	defparam lut_5462.mask = 64'hfcfc00fca8a800a8;

	lut_sub lut_5498 ({g49, g38, g76, g3, g138, g112}, g463);
	defparam lut_5498.LUT_SIZE = 6;
	defparam lut_5498.mask = 64'h55550000f755f300;

	lut_sub lut_5531 ({g73, g440, g461, g462, g463}, g464);
	defparam lut_5531.LUT_SIZE = 5;
	defparam lut_5531.mask = 32'h20202000;

	lut_sub lut_5538 ({i_9_, i_8_, i_6_, i_7_, g76}, g465);
	defparam lut_5538.LUT_SIZE = 5;
	defparam lut_5538.mask = 32'h000000c2;

	lut_sub lut_5546 ({i_5_, i_4_, g11, g465}, g466);
	defparam lut_5546.LUT_SIZE = 4;
	defparam lut_5546.mask = 16'h0010;

	lut_sub lut_5556 ({g30, g58, g457, g460, g464, g466}, g467);
	defparam lut_5556.LUT_SIZE = 6;
	defparam lut_5556.mask = 64'h2000300020002000;

	lut_sub lut_5570 ({g129, g436, g437, g450, g456, g467}, g468);
	defparam lut_5570.LUT_SIZE = 6;
	defparam lut_5570.mask = 64'h0000000001000000;

	lut_sub lut_5579 ({g20, g73, g63, g10, g307}, g469);
	defparam lut_5579.LUT_SIZE = 5;
	defparam lut_5579.mask = 32'h04550c5d;

	lut_sub lut_5598 ({i_2_, i_9_, g36, g54, g75, g51}, g470);
	defparam lut_5598.LUT_SIZE = 6;
	defparam lut_5598.mask = 64'h1111000000000030;

	lut_sub lut_5611 ({g117, g133, g21, g31}, g471);
	defparam lut_5611.LUT_SIZE = 4;
	defparam lut_5611.mask = 16'h50dc;

	lut_sub lut_5625 ({g49, g42, g211, g225}, g472);
	defparam lut_5625.LUT_SIZE = 4;
	defparam lut_5625.mask = 16'h0537;

	lut_sub lut_5640 ({g20, g208, g470, g471, g472}, g473);
	defparam lut_5640.LUT_SIZE = 5;
	defparam lut_5640.mask = 32'h80808000;

	lut_sub lut_5648 ({i_9_, i_8_, i_6_, g469, g473}, g474);
	defparam lut_5648.LUT_SIZE = 5;
	defparam lut_5648.mask = 32'h55555545;

	lut_sub lut_5669 ({g28, g1, g40}, g475);
	defparam lut_5669.LUT_SIZE = 3;
	defparam lut_5669.mask = 8'hd0;

	lut_sub lut_5679 ({g22, g1, g53, g458}, g476);
	defparam lut_5679.LUT_SIZE = 4;
	defparam lut_5679.mask = 16'h1055;

	lut_sub lut_5691 ({i_9_, g28, g63, g45, g94}, g477);
	defparam lut_5691.LUT_SIZE = 5;
	defparam lut_5691.mask = 32'h44440c00;

	lut_sub lut_5705 ({g20, g30, g59, g120, g2}, g478);
	defparam lut_5705.LUT_SIZE = 5;
	defparam lut_5705.mask = 32'h1111111f;

	lut_sub lut_5723 ({g475, g476, g477, g478}, g479);
	defparam lut_5723.LUT_SIZE = 4;
	defparam lut_5723.mask = 16'h8880;

	lut_sub lut_5729 ({i_2_, i_0_, i_1_, i_9_}, g480);
	defparam lut_5729.LUT_SIZE = 4;
	defparam lut_5729.mask = 16'hfddf;

	lut_sub lut_5749 ({i_2_, g78, i_9_, g201, g228}, g481);
	defparam lut_5749.LUT_SIZE = 5;
	defparam lut_5749.mask = 32'h00300050;

	lut_sub lut_5759 ({g22, i_9_, g15, g251}, g482);
	defparam lut_5759.LUT_SIZE = 4;
	defparam lut_5759.mask = 16'h0035;

	lut_sub lut_5770 ({g42, g73, g74, g77}, g483);
	defparam lut_5770.LUT_SIZE = 4;
	defparam lut_5770.mask = 16'h0c5d;

	lut_sub lut_5784 ({g704, g481, g482, g483}, g484);
	defparam lut_5784.LUT_SIZE = 4;
	defparam lut_5784.mask = 16'h0080;

	lut_sub lut_5792 ({g290, g474, g479, g484}, g485);
	defparam lut_5792.LUT_SIZE = 4;
	defparam lut_5792.mask = 16'h0001;

	lut_sub lut_5802 ({g34, g336, g434, g435, g468, g485}, g486);
	defparam lut_5802.LUT_SIZE = 6;
	defparam lut_5802.mask = 64'h0000000000000010;

	lut_sub lut_5809 ({i_2_, g36, g18, g209}, g487);
	defparam lut_5809.LUT_SIZE = 4;
	defparam lut_5809.mask = 16'h5503;

	lut_sub lut_5822 ({g78, i_9_, g16, g29, g487}, g488);
	defparam lut_5822.LUT_SIZE = 5;
	defparam lut_5822.mask = 32'h00035503;

	lut_sub lut_5838 ({g22, g7, g35, g18, g53}, g489);
	defparam lut_5838.LUT_SIZE = 5;
	defparam lut_5838.mask = 32'h00030057;

	lut_sub lut_5852 ({g49, g134, g5, g306}, g490);
	defparam lut_5852.LUT_SIZE = 4;
	defparam lut_5852.mask = 16'haa80;

	lut_sub lut_5865 ({g38, g36, g59, g1, g58}, g491);
	defparam lut_5865.LUT_SIZE = 5;
	defparam lut_5865.mask = 32'h00ce000a;

	lut_sub lut_5881 ({g25, g73, g10, g43, g82, g211}, g492);
	defparam lut_5881.LUT_SIZE = 6;
	defparam lut_5881.mask = 64'h505073735050ff73;

	lut_sub lut_5920 ({g73, g240, g490, g491, g492}, g493);
	defparam lut_5920.LUT_SIZE = 5;
	defparam lut_5920.mask = 32'h08080800;

	lut_sub lut_5931 ({i_9_, g25, g30, g120, g138, g208}, g494);
	defparam lut_5931.LUT_SIZE = 6;
	defparam lut_5931.mask = 64'h0000003311111f1f;

	lut_sub lut_5956 ({g43, g58, g148, g222}, g495);
	defparam lut_5956.LUT_SIZE = 4;
	defparam lut_5956.mask = 16'h7350;

	lut_sub lut_5971 ({g20, g28, g1, g40, g62}, g496);
	defparam lut_5971.LUT_SIZE = 5;
	defparam lut_5971.mask = 32'h1111f111;

	lut_sub lut_5990 ({g118, g392, g494, g495, g496}, g497);
	defparam lut_5990.LUT_SIZE = 5;
	defparam lut_5990.mask = 32'h00800000;

	lut_sub lut_5999 ({g295, g488, g489, g493, g497}, g498);
	defparam lut_5999.LUT_SIZE = 5;
	defparam lut_5999.mask = 32'h10000000;

	lut_sub lut_6008 ({i_9_, g59, g45, g11, g44, g14}, g499);
	defparam lut_6008.LUT_SIZE = 6;
	defparam lut_6008.mask = 64'h000033330a000a00;

	lut_sub lut_6026 ({g36, g119, g18}, g500);
	defparam lut_6026.LUT_SIZE = 3;
	defparam lut_6026.mask = 8'h04;

	lut_sub lut_6034 ({i_2_, g7, g3, g151, g500}, g501);
	defparam lut_6034.LUT_SIZE = 5;
	defparam lut_6034.mask = 32'h11110030;

	lut_sub lut_6048 ({g30, g168, g11, g2, g53}, g502);
	defparam lut_6048.LUT_SIZE = 5;
	defparam lut_6048.mask = 32'h00330537;

	lut_sub lut_6066 ({g279, g499, g501, g502}, g503);
	defparam lut_6066.LUT_SIZE = 4;
	defparam lut_6066.mask = 16'h8000;

	lut_sub lut_6073 ({i_9_, i_8_, g81, g23, g440}, g504);
	defparam lut_6073.LUT_SIZE = 5;
	defparam lut_6073.mask = 32'h00000503;

	lut_sub lut_6084 ({g42, g133, g141, g171}, g505);
	defparam lut_6084.LUT_SIZE = 4;
	defparam lut_6084.mask = 16'h5073;

	lut_sub lut_6098 ({i_9_, g50, g28, g11, g14}, g506);
	defparam lut_6098.LUT_SIZE = 5;
	defparam lut_6098.mask = 32'h30002200;

	lut_sub lut_6110 ({g58, g90, g504, g505, g506}, g507);
	defparam lut_6110.LUT_SIZE = 5;
	defparam lut_6110.mask = 32'h80008080;

	lut_sub lut_6120 ({i_9_, g50, g7, g75, g74}, g508);
	defparam lut_6120.LUT_SIZE = 5;
	defparam lut_6120.mask = 32'h0300aa00;

	lut_sub lut_6133 ({g1, g14, g27, g508}, g509);
	defparam lut_6133.LUT_SIZE = 4;
	defparam lut_6133.mask = 16'h8aaa;

	lut_sub lut_6147 ({g28, g25, g73, g509}, g510);
	defparam lut_6147.LUT_SIZE = 4;
	defparam lut_6147.mask = 16'h5455;

	lut_sub lut_6158 ({i_9_, i_6_, g206}, g511);
	defparam lut_6158.LUT_SIZE = 3;
	defparam lut_6158.mask = 8'h02;

	lut_sub lut_6165 ({i_2_, i_0_, i_1_, g7, g38, g511}, g512);
	defparam lut_6165.LUT_SIZE = 6;
	defparam lut_6165.mask = 64'h0000000400000500;

	lut_sub lut_6174 ({i_2_, i_9_, g272, g141, g244}, g513);
	defparam lut_6174.LUT_SIZE = 5;
	defparam lut_6174.mask = 32'h03000500;

	lut_sub lut_6185 ({i_9_, g39, g6, g122, g55}, g514);
	defparam lut_6185.LUT_SIZE = 5;
	defparam lut_6185.mask = 32'h00335050;

	lut_sub lut_6199 ({g25, g4, g45}, g515);
	defparam lut_6199.LUT_SIZE = 3;
	defparam lut_6199.mask = 8'h08;

	lut_sub lut_6207 ({i_9_, g54, g59, g14, g515}, g516);
	defparam lut_6207.LUT_SIZE = 5;
	defparam lut_6207.mask = 32'h55550c00;

	lut_sub lut_6222 ({i_5_, i_3_, i_4_, g8, g54}, g517);
	defparam lut_6222.LUT_SIZE = 5;
	defparam lut_6222.mask = 32'h00000bb0;

	lut_sub lut_6235 ({g22, i_9_, g36, g20, g517}, g518);
	defparam lut_6235.LUT_SIZE = 5;
	defparam lut_6235.mask = 32'h00000015;

	lut_sub lut_6246 ({g38, g76, g514, g516, g518}, g519);
	defparam lut_6246.LUT_SIZE = 5;
	defparam lut_6246.mask = 32'h808080c0;

	lut_sub lut_6259 ({g59, g58, g512, g513, g519}, g520);
	defparam lut_6259.LUT_SIZE = 5;
	defparam lut_6259.mask = 32'h40444040;

	lut_sub lut_6269 ({g49, i_3_, i_4_, g13}, g521);
	defparam lut_6269.LUT_SIZE = 4;
	defparam lut_6269.mask = 16'h02c0;

	lut_sub lut_6280 ({g50, g76, g13, g46, g157}, g522);
	defparam lut_6280.LUT_SIZE = 5;
	defparam lut_6280.mask = 32'hf0707070;

	lut_sub lut_6299 ({i_5_, g8, g521, g522}, g523);
	defparam lut_6299.LUT_SIZE = 4;
	defparam lut_6299.mask = 16'haaa8;

	lut_sub lut_6311 ({g22, i_9_, i_5_, i_3_, i_4_, g138}, g524);
	defparam lut_6311.LUT_SIZE = 6;
	defparam lut_6311.mask = 64'h0000000000010004;

	lut_sub lut_6320 ({g35, g183, g148, g524}, g525);
	defparam lut_6320.LUT_SIZE = 4;
	defparam lut_6320.mask = 16'haa80;

	lut_sub lut_6332 ({g22, i_9_, g28, g16, g45}, g526);
	defparam lut_6332.LUT_SIZE = 5;
	defparam lut_6332.mask = 32'h000030a0;

	lut_sub lut_6345 ({g120, g43, g161, g251, g228, g526}, g527);
	defparam lut_6345.LUT_SIZE = 6;
	defparam lut_6345.mask = 64'h8000aaaa0000aaaa;

	lut_sub lut_6370 ({g168, g21, g55, g356, g103}, g528);
	defparam lut_6370.LUT_SIZE = 5;
	defparam lut_6370.mask = 32'h80aa00aa;

	lut_sub lut_6386 ({i_9_, g59, g1, g244, g263}, g529);
	defparam lut_6386.LUT_SIZE = 5;
	defparam lut_6386.mask = 32'h70755055;

	lut_sub lut_6408 ({g16, g30, g133, g139, g90}, g530);
	defparam lut_6408.LUT_SIZE = 5;
	defparam lut_6408.mask = 32'h303075f5;

	lut_sub lut_6432 ({g20, g99, g527, g528, g529, g530}, g531);
	defparam lut_6432.LUT_SIZE = 6;
	defparam lut_6432.mask = 64'h0008000800080000;

	lut_sub lut_6440 ({i_9_, i_8_, i_6_, g59, g14}, g532);
	defparam lut_6440.LUT_SIZE = 5;
	defparam lut_6440.mask = 32'h00000002;

	lut_sub lut_6449 ({g20, g137, g52, g71, g532}, g533);
	defparam lut_6449.LUT_SIZE = 5;
	defparam lut_6449.mask = 32'haaa08880;

	lut_sub lut_6464 ({g22, i_7_, i_5_, g92, g192}, g534);
	defparam lut_6464.LUT_SIZE = 5;
	defparam lut_6464.mask = 32'h00000110;

	lut_sub lut_6473 ({i_9_, g6, g165, g193, g534}, g535);
	defparam lut_6473.LUT_SIZE = 5;
	defparam lut_6473.mask = 32'ha0aa88aa;

	lut_sub lut_6489 ({i_9_, i_8_, i_6_, i_7_, g119}, g536);
	defparam lut_6489.LUT_SIZE = 5;
	defparam lut_6489.mask = 32'h00008008;

	lut_sub lut_6499 ({i_2_, g7, g75, g73, g14, g40}, g537);
	defparam lut_6499.LUT_SIZE = 6;
	defparam lut_6499.mask = 64'h000c005d0000000f;

	lut_sub lut_6518 ({g27, g29, g475, g536, g537}, g538);
	defparam lut_6518.LUT_SIZE = 5;
	defparam lut_6518.mask = 32'haaa8a8a8;

	lut_sub lut_6539 ({g303, g697, g533, g535, g538}, g539);
	defparam lut_6539.LUT_SIZE = 5;
	defparam lut_6539.mask = 32'h00010000;

	lut_sub lut_6549 ({g774, g114, g523, g525, g531, g539}, g540);
	defparam lut_6549.LUT_SIZE = 6;
	defparam lut_6549.mask = 64'h0000000000000001;

	lut_sub lut_6559 ({g227, g338, g434, g510, g520, g540}, g541);
	defparam lut_6559.LUT_SIZE = 6;
	defparam lut_6559.mask = 64'h0000000000000001;

	lut_sub lut_6568 ({g381, g498, g503, g507, g541}, g542);
	defparam lut_6568.LUT_SIZE = 5;
	defparam lut_6568.mask = 32'h00000001;

	lut_sub lut_6576 ({g20, g52, g58, g302}, g543);
	defparam lut_6576.LUT_SIZE = 4;
	defparam lut_6576.mask = 16'hf2a2;

	lut_sub lut_6591 ({i_9_, g6, g46, g19, g488}, g544);
	defparam lut_6591.LUT_SIZE = 5;
	defparam lut_6591.mask = 32'h88aaa0aa;

	lut_sub lut_6611 ({g220, g339, g424, g543, g544}, g545);
	defparam lut_6611.LUT_SIZE = 5;
	defparam lut_6611.mask = 32'h51000000;

	lut_sub lut_6619 ({i_0_, i_1_, g135, g251}, g546);
	defparam lut_6619.LUT_SIZE = 4;
	defparam lut_6619.mask = 16'h0305;

	lut_sub lut_6628 ({i_2_, i_9_, g546, g690}, g547);
	defparam lut_6628.LUT_SIZE = 4;
	defparam lut_6628.mask = 16'h4555;

	lut_sub lut_6641 ({i_8_, g36, g68, g59}, g548);
	defparam lut_6641.LUT_SIZE = 4;
	defparam lut_6641.mask = 16'hfe00;

	lut_sub lut_6654 ({g22, i_9_, i_8_, g83, g10}, g549);
	defparam lut_6654.LUT_SIZE = 5;
	defparam lut_6654.mask = 32'h00f000f2;

	lut_sub lut_6666 ({i_9_, i_6_, i_7_}, g550);
	defparam lut_6666.LUT_SIZE = 3;
	defparam lut_6666.mask = 8'h08;

	lut_sub lut_6674 ({i_8_, g39, g30, g71, g550}, g551);
	defparam lut_6674.LUT_SIZE = 5;
	defparam lut_6674.mask = 32'h00051111;

	lut_sub lut_6688 ({i_9_, g38, g30, g59, g94, g46}, g552);
	defparam lut_6688.LUT_SIZE = 6;
	defparam lut_6688.mask = 64'h373f0505333f0000;

	lut_sub lut_6721 ({g49, g35, g116, g135, g259}, g553);
	defparam lut_6721.LUT_SIZE = 5;
	defparam lut_6721.mask = 32'hffaac080;

	lut_sub lut_6744 ({i_9_, g50, g28, g63, g11, g182}, g554);
	defparam lut_6744.LUT_SIZE = 6;
	defparam lut_6744.mask = 64'h111111113f000000;

	lut_sub lut_6765 ({g101, g42, g209, g148}, g555);
	defparam lut_6765.LUT_SIZE = 4;
	defparam lut_6765.mask = 16'h070f;

	lut_sub lut_6779 ({g268, g553, g554, g555}, g556);
	defparam lut_6779.LUT_SIZE = 4;
	defparam lut_6779.mask = 16'h0800;

	lut_sub lut_6788 ({g548, g549, g551, g552, g556}, g557);
	defparam lut_6788.LUT_SIZE = 5;
	defparam lut_6788.mask = 32'h40004040;

	lut_sub lut_6798 ({i_9_, g50, g7, g45, g11}, g558);
	defparam lut_6798.LUT_SIZE = 5;
	defparam lut_6798.mask = 32'h04040500;

	lut_sub lut_6810 ({g43, g37, g230, g225, g558}, g559);
	defparam lut_6810.LUT_SIZE = 5;
	defparam lut_6810.mask = 32'h0080aaaa;

	lut_sub lut_6825 ({i_9_, g16, g138, g112}, g560);
	defparam lut_6825.LUT_SIZE = 4;
	defparam lut_6825.mask = 16'h1105;

	lut_sub lut_6836 ({g13, g158, g259, g560}, g561);
	defparam lut_6836.LUT_SIZE = 4;
	defparam lut_6836.mask = 16'h80aa;

	lut_sub lut_6846 ({i_2_, i_9_, g36, g76}, g562);
	defparam lut_6846.LUT_SIZE = 4;
	defparam lut_6846.mask = 16'ha003;

	lut_sub lut_6858 ({g54, g10, g133, g18, g141}, g563);
	defparam lut_6858.LUT_SIZE = 5;
	defparam lut_6858.mask = 32'hf0507050;

	lut_sub lut_6876 ({g50, g75, g562, g563}, g564);
	defparam lut_6876.LUT_SIZE = 4;
	defparam lut_6876.mask = 16'ha8aa;

	lut_sub lut_6892 ({g81, g35, g10, g2, g233, g228}, g565);
	defparam lut_6892.LUT_SIZE = 6;
	defparam lut_6892.mask = 64'h030357570f035f57;

	lut_sub lut_6926 ({i_9_, i_8_, i_5_, i_3_, i_4_}, g566);
	defparam lut_6926.LUT_SIZE = 5;
	defparam lut_6926.mask = 32'h00000021;

	lut_sub lut_6935 ({i_7_, g6, g73, g14, g566}, g567);
	defparam lut_6935.LUT_SIZE = 5;
	defparam lut_6935.mask = 32'h45000000;

	lut_sub lut_6944 ({i_2_, i_0_, i_1_, g28, g73, g40}, g568);
	defparam lut_6944.LUT_SIZE = 6;
	defparam lut_6944.mask = 64'h5000305000000000;

	lut_sub lut_6957 ({g7, g27, g567, g568}, g569);
	defparam lut_6957.LUT_SIZE = 4;
	defparam lut_6957.mask = 16'ha888;

	lut_sub lut_6970 ({g559, g561, g564, g565, g569}, g570);
	defparam lut_6970.LUT_SIZE = 5;
	defparam lut_6970.mask = 32'h00000004;

	lut_sub lut_6976 ({i_9_, i_8_, g81, g124}, g571);
	defparam lut_6976.LUT_SIZE = 4;
	defparam lut_6976.mask = 16'h0110;

	lut_sub lut_6987 ({g39, g20, g10, g14, g58, g424}, g572);
	defparam lut_6987.LUT_SIZE = 6;
	defparam lut_6987.mask = 64'h0000000054005450;

	lut_sub lut_7002 ({g49, g32, g157, g251}, g573);
	defparam lut_7002.LUT_SIZE = 4;
	defparam lut_7002.mask = 16'h007f;

	lut_sub lut_7017 ({g460, g464, g571, g572, g573}, g574);
	defparam lut_7017.LUT_SIZE = 5;
	defparam lut_7017.mask = 32'h00800000;

	lut_sub lut_7025 ({i_2_, i_9_, g28, g119, g16, g180}, g575);
	defparam lut_7025.LUT_SIZE = 6;
	defparam lut_7025.mask = 64'h0000300030005050;

	lut_sub lut_7041 ({i_9_, g7, g36, g16, g45, g11}, g576);
	defparam lut_7041.LUT_SIZE = 6;
	defparam lut_7041.mask = 64'h0000000000054445;

	lut_sub lut_7054 ({i_9_, g7, g3, g125}, g577);
	defparam lut_7054.LUT_SIZE = 4;
	defparam lut_7054.mask = 16'h0c55;

	lut_sub lut_7064 ({i_9_, i_3_, i_4_, g25}, g578);
	defparam lut_7064.LUT_SIZE = 4;
	defparam lut_7064.mask = 16'h4004;

	lut_sub lut_7073 ({i_5_, g54, g63, g577, g578}, g579);
	defparam lut_7073.LUT_SIZE = 5;
	defparam lut_7073.mask = 32'h57030303;

	lut_sub lut_7092 ({i_9_, g39, g3, g92, g117, g224}, g580);
	defparam lut_7092.LUT_SIZE = 6;
	defparam lut_7092.mask = 64'h0000333355005f00;

	lut_sub lut_7117 ({g26, g58, g53, g440}, g581);
	defparam lut_7117.LUT_SIZE = 4;
	defparam lut_7117.mask = 16'h5073;

	lut_sub lut_7132 ({i_9_, g25, g120, g183, g179, g581}, g582);
	defparam lut_7132.LUT_SIZE = 6;
	defparam lut_7132.mask = 64'haaaa8800aaaaa0a0;

	lut_sub lut_7162 ({g575, g576, g579, g580, g582}, g583);
	defparam lut_7162.LUT_SIZE = 5;
	defparam lut_7162.mask = 32'h40000000;

	lut_sub lut_7172 ({g547, g735, g557, g570, g574, g583}, g584);
	defparam lut_7172.LUT_SIZE = 6;
	defparam lut_7172.mask = 64'h0000000000000001;

	lut_sub lut_7181 ({g89, g372, g507, g545, g584}, g585);
	defparam lut_7181.LUT_SIZE = 5;
	defparam lut_7181.mask = 32'h00000001;

	lut_sub lut_7188 ({i_9_, g101, g59, g141}, g586);
	defparam lut_7188.LUT_SIZE = 4;
	defparam lut_7188.mask = 16'h0311;

	lut_sub lut_7199 ({g22, g36, g26, g53}, g587);
	defparam lut_7199.LUT_SIZE = 4;
	defparam lut_7199.mask = 16'h1115;

	lut_sub lut_7211 ({g50, g35, g76, g587}, g588);
	defparam lut_7211.LUT_SIZE = 4;
	defparam lut_7211.mask = 16'ha2aa;

	lut_sub lut_7225 ({g124, g137, g2, g46}, g589);
	defparam lut_7225.LUT_SIZE = 4;
	defparam lut_7225.mask = 16'h111f;

	lut_sub lut_7240 ({g22, g36, g6, g73, g4}, g590);
	defparam lut_7240.LUT_SIZE = 5;
	defparam lut_7240.mask = 32'h00302232;

	lut_sub lut_7254 ({g39, g20, g30, g59}, g591);
	defparam lut_7254.LUT_SIZE = 4;
	defparam lut_7254.mask = 16'h0103;

	lut_sub lut_7265 ({g42, g116, g340, g590, g591}, g592);
	defparam lut_7265.LUT_SIZE = 5;
	defparam lut_7265.mask = 32'h80808000;

	lut_sub lut_7276 ({g404, g586, g588, g589, g592}, g593);
	defparam lut_7276.LUT_SIZE = 5;
	defparam lut_7276.mask = 32'h00000400;

	lut_sub lut_7284 ({g62, g27, g192, g224}, g594);
	defparam lut_7284.LUT_SIZE = 4;
	defparam lut_7284.mask = 16'h0537;

	lut_sub lut_7298 ({g49, g17, g193, g594}, g595);
	defparam lut_7298.LUT_SIZE = 4;
	defparam lut_7298.mask = 16'haa80;

	lut_sub lut_7310 ({g125, g13, g2, g161}, g596);
	defparam lut_7310.LUT_SIZE = 4;
	defparam lut_7310.mask = 16'h11f1;

	lut_sub lut_7324 ({g495, g325, g595, g596}, g597);
	defparam lut_7324.LUT_SIZE = 4;
	defparam lut_7324.mask = 16'h0200;

	lut_sub lut_7332 ({i_9_, g39, g45, g139, g208}, g598);
	defparam lut_7332.LUT_SIZE = 5;
	defparam lut_7332.mask = 32'h00335050;

	lut_sub lut_7346 ({i_9_, g120, g11, g5}, g599);
	defparam lut_7346.LUT_SIZE = 4;
	defparam lut_7346.mask = 16'h1103;

	lut_sub lut_7356 ({i_9_, g63, g179, g158}, g600);
	defparam lut_7356.LUT_SIZE = 4;
	defparam lut_7356.mask = 16'h0503;

	lut_sub lut_7367 ({g22, i_9_, g10, g45, g148}, g601);
	defparam lut_7367.LUT_SIZE = 5;
	defparam lut_7367.mask = 32'h000055c0;

	lut_sub lut_7381 ({g365, g598, g599, g600, g601}, g602);
	defparam lut_7381.LUT_SIZE = 5;
	defparam lut_7381.mask = 32'h80000000;

	lut_sub lut_7389 ({i_9_, g59, g177, g55, g602}, g603);
	defparam lut_7389.LUT_SIZE = 5;
	defparam lut_7389.mask = 32'h55445550;

	lut_sub lut_7407 ({i_2_, i_9_, g272, g156, g169}, g604);
	defparam lut_7407.LUT_SIZE = 5;
	defparam lut_7407.mask = 32'h03000005;

	lut_sub lut_7417 ({g28, g3, g1}, g605);
	defparam lut_7417.LUT_SIZE = 3;
	defparam lut_7417.mask = 8'h80;

	lut_sub lut_7426 ({g7, g20, g16, g63, g13}, g606);
	defparam lut_7426.LUT_SIZE = 5;
	defparam lut_7426.mask = 32'h00000a3b;

	lut_sub lut_7439 ({g133, g139, g606}, g607);
	defparam lut_7439.LUT_SIZE = 3;
	defparam lut_7439.mask = 8'h8a;

	lut_sub lut_7449 ({g101, g42, g43, g180}, g608);
	defparam lut_7449.LUT_SIZE = 4;
	defparam lut_7449.mask = 16'h05cd;

	lut_sub lut_7464 ({g57, g40, g457, g607, g608}, g609);
	defparam lut_7464.LUT_SIZE = 5;
	defparam lut_7464.mask = 32'h20202000;

	lut_sub lut_7475 ({i_9_, g39, g239, g356, g605, g609}, g610);
	defparam lut_7475.LUT_SIZE = 6;
	defparam lut_7475.mask = 64'h5500500044004400;

	lut_sub lut_7491 ({i_5_, i_3_, i_4_, g63, g137, g58}, g611);
	defparam lut_7491.LUT_SIZE = 6;
	defparam lut_7491.mask = 64'h000300000000000a;

	lut_sub lut_7503 ({g7, g28, g73, g59, g1}, g612);
	defparam lut_7503.LUT_SIZE = 5;
	defparam lut_7503.mask = 32'h03000b0a;

	lut_sub lut_7517 ({i_9_, g50, i_5_, g6, g92, g45}, g613);
	defparam lut_7517.LUT_SIZE = 6;
	defparam lut_7517.mask = 64'h2000200000300000;

	lut_sub lut_7528 ({g38, g1, g14, g613}, g614);
	defparam lut_7528.LUT_SIZE = 4;
	defparam lut_7528.mask = 16'h2aaa;

	lut_sub lut_7543 ({g7, g28, g25, g6, g40}, g615);
	defparam lut_7543.LUT_SIZE = 5;
	defparam lut_7543.mask = 32'h05004545;

	lut_sub lut_7560 ({g38, g42, g122, g17, g46, g29}, g616);
	defparam lut_7560.LUT_SIZE = 6;
	defparam lut_7560.mask = 64'haaaa8000ffffc000;

	lut_sub lut_7595 ({g101, g21, g53, g23, g97}, g617);
	defparam lut_7595.LUT_SIZE = 5;
	defparam lut_7595.mask = 32'ha8fc00fc;

	lut_sub lut_7618 ({g21, g165, g615, g616, g617}, g618);
	defparam lut_7618.LUT_SIZE = 5;
	defparam lut_7618.mask = 32'h10001010;

	lut_sub lut_7629 ({g13, g177, g612, g614, g618}, g619);
	defparam lut_7629.LUT_SIZE = 5;
	defparam lut_7629.mask = 32'h10001010;

	lut_sub lut_7639 ({g8, g36, g122, g133}, g620);
	defparam lut_7639.LUT_SIZE = 4;
	defparam lut_7639.mask = 16'h222a;

	lut_sub lut_7651 ({g35, g43, g165, g244}, g621);
	defparam lut_7651.LUT_SIZE = 4;
	defparam lut_7651.mask = 16'h3075;

	lut_sub lut_7666 ({g7, g39, g16, g133, g53}, g622);
	defparam lut_7666.LUT_SIZE = 5;
	defparam lut_7666.mask = 32'h00000c5d;

	lut_sub lut_7681 ({g620, g176, g185, g621, g622}, g623);
	defparam lut_7681.LUT_SIZE = 5;
	defparam lut_7681.mask = 32'h00080000;

	lut_sub lut_7690 ({g604, g610, g611, g619, g623}, g624);
	defparam lut_7690.LUT_SIZE = 5;
	defparam lut_7690.mask = 32'h00100000;

	lut_sub lut_7696 ({i_9_, i_8_, i_6_, i_7_, g99, g195}, g625);
	defparam lut_7696.LUT_SIZE = 6;
	defparam lut_7696.mask = 64'h0000000000003500;

	lut_sub lut_7708 ({g547, g397, g474, g503, g625}, g626);
	defparam lut_7708.LUT_SIZE = 5;
	defparam lut_7708.mask = 32'h00000002;

	lut_sub lut_7718 ({g237, g593, g597, g603, g624, g626}, g627);
	defparam lut_7718.LUT_SIZE = 6;
	defparam lut_7718.mask = 64'h0000000000000001;

	lut_sub lut_7725 ({g22, i_9_, g182, g186}, g628);
	defparam lut_7725.LUT_SIZE = 4;
	defparam lut_7725.mask = 16'h0053;

	lut_sub lut_7736 ({g20, g137, g60, g307}, g629);
	defparam lut_7736.LUT_SIZE = 4;
	defparam lut_7736.mask = 16'h0357;

	lut_sub lut_7751 ({g38, g137, g52, g222, g331}, g630);
	defparam lut_7751.LUT_SIZE = 5;
	defparam lut_7751.mask = 32'h05150111;

	lut_sub lut_7767 ({g76, g3, g21, g171, g193}, g631);
	defparam lut_7767.LUT_SIZE = 5;
	defparam lut_7767.mask = 32'hf0707070;

	lut_sub lut_7787 ({g53, g440, g630, g631}, g632);
	defparam lut_7787.LUT_SIZE = 4;
	defparam lut_7787.mask = 16'h8880;

	lut_sub lut_7798 ({g43, g209, g628, g629, g632}, g633);
	defparam lut_7798.LUT_SIZE = 5;
	defparam lut_7798.mask = 32'h40004040;

	lut_sub lut_7806 ({i_5_, i_3_, i_4_, g25, g137}, g634);
	defparam lut_7806.LUT_SIZE = 5;
	defparam lut_7806.mask = 32'h00000013;

	lut_sub lut_7813 ({i_9_, i_8_, i_6_, g634}, g635);
	defparam lut_7813.LUT_SIZE = 4;
	defparam lut_7813.mask = 16'h0040;

	lut_sub lut_7822 ({g40, g243, g440, g633, g635}, g636);
	defparam lut_7822.LUT_SIZE = 5;
	defparam lut_7822.mask = 32'h32002200;

	lut_sub lut_7834 ({i_9_, g6, g30, g134, g138}, g637);
	defparam lut_7834.LUT_SIZE = 5;
	defparam lut_7834.mask = 32'h33000500;

	lut_sub lut_7847 ({i_9_, g7, g63, g30, g138}, g638);
	defparam lut_7847.LUT_SIZE = 5;
	defparam lut_7847.mask = 32'h01010005;

	lut_sub lut_7854 ({i_9_, i_8_, i_6_, i_7_, i_5_}, g639);
	defparam lut_7854.LUT_SIZE = 5;
	defparam lut_7854.mask = 32'h00000042;

	lut_sub lut_7861 ({i_3_, i_4_, g1, g639}, g640);
	defparam lut_7861.LUT_SIZE = 4;
	defparam lut_7861.mask = 16'h0040;

	lut_sub lut_7869 ({g13, g85, g638, g640}, g641);
	defparam lut_7869.LUT_SIZE = 4;
	defparam lut_7869.mask = 16'h8088;

	lut_sub lut_7880 ({g36, g54, g28, g6, g58}, g642);
	defparam lut_7880.LUT_SIZE = 5;
	defparam lut_7880.mask = 32'h8080cc80;

	lut_sub lut_7894 ({i_2_, g78, i_9_, g122, g168, g85}, g643);
	defparam lut_7894.LUT_SIZE = 6;
	defparam lut_7894.mask = 64'h0000330f00005533;

	lut_sub lut_7918 ({i_9_, g39, g1, g37, g32, g228}, g644);
	defparam lut_7918.LUT_SIZE = 6;
	defparam lut_7918.mask = 64'hf000f3335500f5f0;

	lut_sub lut_7951 ({i_9_, i_5_, i_3_, i_4_, g3, g11}, g645);
	defparam lut_7951.LUT_SIZE = 6;
	defparam lut_7951.mask = 64'h0000404000000004;

	lut_sub lut_7963 ({g35, g42, g3, g10, g18, g21}, g646);
	defparam lut_7963.LUT_SIZE = 6;
	defparam lut_7963.mask = 64'h2020f020f020f020;

	lut_sub lut_7988 ({g7, g16, g43, g645, g646}, g647);
	defparam lut_7988.LUT_SIZE = 5;
	defparam lut_7988.mask = 32'h88888808;

	lut_sub lut_8003 ({g641, g642, g643, g644, g647}, g648);
	defparam lut_8003.LUT_SIZE = 5;
	defparam lut_8003.mask = 32'h00004000;

	lut_sub lut_8010 ({g78, g54, g10}, g649);
	defparam lut_8010.LUT_SIZE = 3;
	defparam lut_8010.mask = 8'h08;

	lut_sub lut_8018 ({i_2_, g16, g14, g151, g649}, g650);
	defparam lut_8018.LUT_SIZE = 5;
	defparam lut_8018.mask = 32'h11110030;

	lut_sub lut_8031 ({g22, i_9_, g1, g44, g156}, g651);
	defparam lut_8031.LUT_SIZE = 5;
	defparam lut_8031.mask = 32'h30003055;

	lut_sub lut_8046 ({i_9_, g16, g63, g156, g354}, g652);
	defparam lut_8046.LUT_SIZE = 5;
	defparam lut_8046.mask = 32'h03030055;

	lut_sub lut_8061 ({g22, i_9_, g7, g40, g356}, g653);
	defparam lut_8061.LUT_SIZE = 5;
	defparam lut_8061.mask = 32'h00005703;

	lut_sub lut_8076 ({g133, g422, g651, g652, g653}, g654);
	defparam lut_8076.LUT_SIZE = 5;
	defparam lut_8076.mask = 32'h80008080;

	lut_sub lut_8086 ({g219, g494, g650, g654}, g655);
	defparam lut_8086.LUT_SIZE = 4;
	defparam lut_8086.mask = 16'h0040;

	lut_sub lut_8095 ({g147, g610, g637, g648, g655}, g656);
	defparam lut_8095.LUT_SIZE = 5;
	defparam lut_8095.mask = 32'h00000010;

	lut_sub lut_8103 ({i_9_, g39, g3, g30, g77}, g657);
	defparam lut_8103.LUT_SIZE = 5;
	defparam lut_8103.mask = 32'h00300055;

	lut_sub lut_8115 ({i_9_, g25, g17, g139}, g658);
	defparam lut_8115.LUT_SIZE = 4;
	defparam lut_8115.mask = 16'h0305;

	lut_sub lut_8124 ({i_2_, g78, i_9_, g4}, g659);
	defparam lut_8124.LUT_SIZE = 4;
	defparam lut_8124.mask = 16'h0b03;

	lut_sub lut_8137 ({g787, g401, g657, g658, g659}, g660);
	defparam lut_8137.LUT_SIZE = 5;
	defparam lut_8137.mask = 32'h0000c080;

	lut_sub lut_8148 ({g294, g382, g391, g510, g660}, g661);
	defparam lut_8148.LUT_SIZE = 5;
	defparam lut_8148.mask = 32'h00000100;

	lut_sub lut_8158 ({g317, g479, g557, g636, g656, g661}, g662);
	defparam lut_8158.LUT_SIZE = 6;
	defparam lut_8158.mask = 64'h0000000000000001;

	lut_sub lut_8166 ({i_9_, g45, g221, g138, g302}, g663);
	defparam lut_8166.LUT_SIZE = 5;
	defparam lut_8166.mask = 32'h0f001111;

	lut_sub lut_8177 ({i_9_, i_8_, i_6_, i_7_, i_5_}, g664);
	defparam lut_8177.LUT_SIZE = 5;
	defparam lut_8177.mask = 32'h00002040;

	lut_sub lut_8185 ({g22, i_3_, i_4_, g206, g664}, g665);
	defparam lut_8185.LUT_SIZE = 5;
	defparam lut_8185.mask = 32'h00000100;

	lut_sub lut_8193 ({i_9_, g8, g59, g10, g142}, g666);
	defparam lut_8193.LUT_SIZE = 5;
	defparam lut_8193.mask = 32'h00aa000c;

	lut_sub lut_8207 ({g35, g116, g43, g158, g193}, g667);
	defparam lut_8207.LUT_SIZE = 5;
	defparam lut_8207.mask = 32'hcf0f8a0a;

	lut_sub lut_8229 ({g13, g141, g225, g667}, g668);
	defparam lut_8229.LUT_SIZE = 4;
	defparam lut_8229.mask = 16'h4055;

	lut_sub lut_8238 ({i_9_, i_8_, i_6_, g221}, g669);
	defparam lut_8238.LUT_SIZE = 4;
	defparam lut_8238.mask = 16'h0001;

	lut_sub lut_8244 ({i_9_, i_5_, g16, g138}, g670);
	defparam lut_8244.LUT_SIZE = 4;
	defparam lut_8244.mask = 16'h0053;

	lut_sub lut_8254 ({i_3_, i_4_, g63, g669, g670}, g671);
	defparam lut_8254.LUT_SIZE = 5;
	defparam lut_8254.mask = 32'hc8cccccc;

	lut_sub lut_8277 ({g663, g665, g666, g668, g671}, g672);
	defparam lut_8277.LUT_SIZE = 5;
	defparam lut_8277.mask = 32'h10000000;

	lut_sub lut_8283 ({g22, i_9_, i_3_, i_4_, g68}, g673);
	defparam lut_8283.LUT_SIZE = 5;
	defparam lut_8283.mask = 32'h00000004;

	lut_sub lut_8292 ({g7, g20, g76, g137, g673}, g674);
	defparam lut_8292.LUT_SIZE = 5;
	defparam lut_8292.mask = 32'h10115055;

	lut_sub lut_8306 ({g242, g232}, g675);
	defparam lut_8306.LUT_SIZE = 2;
	defparam lut_8306.mask = 4'b0001;

	lut_sub lut_8314 ({g16, g45, g133, g14}, g676);
	defparam lut_8314.LUT_SIZE = 4;
	defparam lut_8314.mask = 16'h8088;

	lut_sub lut_8324 ({g7, g1, g27, g676}, g677);
	defparam lut_8324.LUT_SIZE = 4;
	defparam lut_8324.mask = 16'haa8a;

	lut_sub lut_8338 ({i_2_, i_9_, g119, g182, g55, g97}, g678);
	defparam lut_8338.LUT_SIZE = 6;
	defparam lut_8338.mask = 64'h550033000f005500;

	lut_sub lut_8361 ({i_9_, g30, g59, g45, g18}, g679);
	defparam lut_8361.LUT_SIZE = 5;
	defparam lut_8361.mask = 32'h0005000c;

	lut_sub lut_8373 ({g21, g40, g112, g233, g679}, g680);
	defparam lut_8373.LUT_SIZE = 5;
	defparam lut_8373.mask = 32'h8880aaa0;

	lut_sub lut_8390 ({g38, g25, g4, g10, g11}, g681);
	defparam lut_8390.LUT_SIZE = 5;
	defparam lut_8390.mask = 32'h50dc0000;

	lut_sub lut_8404 ({g2, g158, g201, g681}, g682);
	defparam lut_8404.LUT_SIZE = 4;
	defparam lut_8404.mask = 16'haa80;

	lut_sub lut_8418 ({g28, g42, g59, g10, g18, g58}, g683);
	defparam lut_8418.LUT_SIZE = 6;
	defparam lut_8418.mask = 64'h00aa33bb00a000a0;

	lut_sub lut_8443 ({i_8_, g7, g35, g68, g42}, g684);
	defparam lut_8443.LUT_SIZE = 5;
	defparam lut_8443.mask = 32'h00110013;

	lut_sub lut_8455 ({g35, g180, g259, g684}, g685);
	defparam lut_8455.LUT_SIZE = 4;
	defparam lut_8455.mask = 16'haa80;

	lut_sub lut_8467 ({g680, g682, g683, g685}, g686);
	defparam lut_8467.LUT_SIZE = 4;
	defparam lut_8467.mask = 16'h0004;

	lut_sub lut_8475 ({g155, g677, g678, g686}, g687);
	defparam lut_8475.LUT_SIZE = 4;
	defparam lut_8475.mask = 16'h0004;

	lut_sub lut_8485 ({g575, g593, g633, g674, g675, g687}, g688);
	defparam lut_8485.LUT_SIZE = 6;
	defparam lut_8485.mask = 64'h0000001000000000;

	lut_sub lut_8495 ({g321, g414, g484, g498, g672, g688}, g689);
	defparam lut_8495.LUT_SIZE = 6;
	defparam lut_8495.mask = 64'h0000000000000001;

	lut_sub lut_8501 ({g4, g691}, g690);
	defparam lut_8501.LUT_SIZE = 2;
	defparam lut_8501.mask = 4'b1000;

	lut_sub lut_8507 ({g4, g692}, g691);
	defparam lut_8507.LUT_SIZE = 2;
	defparam lut_8507.mask = 4'b0100;

	lut_sub lut_8513 ({g693, g694}, g692);
	defparam lut_8513.LUT_SIZE = 2;
	defparam lut_8513.mask = 4'b1000;

	lut_sub lut_8518 ({i_1_, g695}, g693);
	defparam lut_8518.LUT_SIZE = 2;
	defparam lut_8518.mask = 4'b0100;

	lut_sub lut_8523 ({i_1_, g696}, g694);
	defparam lut_8523.LUT_SIZE = 2;
	defparam lut_8523.mask = 4'b0001;

	lut_sub lut_8529 ({g511, i_0_, g38, i_2_}, g695);
	defparam lut_8529.LUT_SIZE = 4;
	defparam lut_8529.mask = 16'hff7f;

	lut_sub lut_8549 ({g511, i_0_, g58, i_2_}, g696);
	defparam lut_8549.LUT_SIZE = 4;
	defparam lut_8549.mask = 16'hfff7;

	lut_sub lut_8568 ({i_9_, g698}, g697);
	defparam lut_8568.LUT_SIZE = 2;
	defparam lut_8568.mask = 4'b0010;

	lut_sub lut_8573 ({i_9_, g699}, g698);
	defparam lut_8573.LUT_SIZE = 2;
	defparam lut_8573.mask = 4'b0001;

	lut_sub lut_8579 ({g700, g701}, g699);
	defparam lut_8579.LUT_SIZE = 2;
	defparam lut_8579.mask = 4'b1000;

	lut_sub lut_8584 ({i_7_, g702}, g700);
	defparam lut_8584.LUT_SIZE = 2;
	defparam lut_8584.mask = 4'b0100;

	lut_sub lut_8589 ({i_7_, g703}, g701);
	defparam lut_8589.LUT_SIZE = 2;
	defparam lut_8589.mask = 4'b0001;

	lut_sub lut_8595 ({g6, i_6_, g7, i_8_}, g702);
	defparam lut_8595.LUT_SIZE = 4;
	defparam lut_8595.mask = 16'hfeff;

	lut_sub lut_8614 ({i_6_, g74, i_8_}, g703);
	defparam lut_8614.LUT_SIZE = 3;
	defparam lut_8614.mask = 8'h7f;

	lut_sub lut_8625 ({i_5_, g705}, g704);
	defparam lut_8625.LUT_SIZE = 2;
	defparam lut_8625.mask = 4'b1000;

	lut_sub lut_8630 ({i_5_, g706}, g705);
	defparam lut_8630.LUT_SIZE = 2;
	defparam lut_8630.mask = 4'b0100;

	lut_sub lut_8636 ({g707, g708}, g706);
	defparam lut_8636.LUT_SIZE = 2;
	defparam lut_8636.mask = 4'b1000;

	lut_sub lut_8641 ({i_4_, g709}, g707);
	defparam lut_8641.LUT_SIZE = 2;
	defparam lut_8641.mask = 4'b0100;

	lut_sub lut_8646 ({i_4_, g710}, g708);
	defparam lut_8646.LUT_SIZE = 2;
	defparam lut_8646.mask = 4'b0001;

	lut_sub lut_8653 ({g480, g138, g13, i_3_}, g709);
	defparam lut_8653.LUT_SIZE = 4;
	defparam lut_8653.mask = 16'hf7ff;

	lut_sub lut_8674 ({g480, g138, g43, i_3_}, g710);
	defparam lut_8674.LUT_SIZE = 4;
	defparam lut_8674.mask = 16'hf7ff;

	lut_sub lut_8694 ({g712, g713}, g711);
	defparam lut_8694.LUT_SIZE = 2;
	defparam lut_8694.mask = 4'b1000;

	lut_sub lut_8700 ({g358, g714}, g712);
	defparam lut_8700.LUT_SIZE = 2;
	defparam lut_8700.mask = 4'b0100;

	lut_sub lut_8706 ({g358, g717}, g713);
	defparam lut_8706.LUT_SIZE = 2;
	defparam lut_8706.mask = 4'b0001;

	lut_sub lut_8712 ({g715, g716}, g714);
	defparam lut_8712.LUT_SIZE = 2;
	defparam lut_8712.mask = 4'b1000;

	lut_sub lut_8717 ({i_4_, g719}, g715);
	defparam lut_8717.LUT_SIZE = 2;
	defparam lut_8717.mask = 4'b0100;

	lut_sub lut_8722 ({i_4_, g720}, g716);
	defparam lut_8722.LUT_SIZE = 2;
	defparam lut_8722.mask = 4'b0001;

	lut_sub lut_8727 ({i_4_, g718}, g717);
	defparam lut_8727.LUT_SIZE = 2;
	defparam lut_8727.mask = 4'b0010;

	lut_sub lut_8732 ({i_4_, g721}, g718);
	defparam lut_8732.LUT_SIZE = 2;
	defparam lut_8732.mask = 4'b0001;

	lut_sub lut_8737 ({i_3_, g119, i_5_}, g719);
	defparam lut_8737.LUT_SIZE = 3;
	defparam lut_8737.mask = 8'hfb;

	lut_sub lut_8749 ({g21, i_3_, g138, i_5_}, g720);
	defparam lut_8749.LUT_SIZE = 4;
	defparam lut_8749.mask = 16'hdeff;

	lut_sub lut_8768 ({g21, i_3_, g138, i_5_}, g721);
	defparam lut_8768.LUT_SIZE = 4;
	defparam lut_8768.mask = 16'hdeff;

	lut_sub lut_8786 ({i_9_, g723}, g722);
	defparam lut_8786.LUT_SIZE = 2;
	defparam lut_8786.mask = 4'b0010;

	lut_sub lut_8791 ({i_9_, g724}, g723);
	defparam lut_8791.LUT_SIZE = 2;
	defparam lut_8791.mask = 4'b0001;

	lut_sub lut_8797 ({g725, g726}, g724);
	defparam lut_8797.LUT_SIZE = 2;
	defparam lut_8797.mask = 4'b1000;

	lut_sub lut_8802 ({i_7_, g727}, g725);
	defparam lut_8802.LUT_SIZE = 2;
	defparam lut_8802.mask = 4'b0100;

	lut_sub lut_8807 ({i_7_, g728}, g726);
	defparam lut_8807.LUT_SIZE = 2;
	defparam lut_8807.mask = 4'b0001;

	lut_sub lut_8812 ({i_6_, g142, i_8_}, g727);
	defparam lut_8812.LUT_SIZE = 3;
	defparam lut_8812.mask = 8'hbf;

	lut_sub lut_8824 ({g11, i_6_, g14, i_8_}, g728);
	defparam lut_8824.LUT_SIZE = 4;
	defparam lut_8824.mask = 16'hffbf;

	lut_sub lut_8844 ({g280, g730}, g729);
	defparam lut_8844.LUT_SIZE = 2;
	defparam lut_8844.mask = 4'b0001;

	lut_sub lut_8850 ({g731, g732}, g730);
	defparam lut_8850.LUT_SIZE = 2;
	defparam lut_8850.mask = 4'b1000;

	lut_sub lut_8855 ({i_8_, g733}, g731);
	defparam lut_8855.LUT_SIZE = 2;
	defparam lut_8855.mask = 4'b0100;

	lut_sub lut_8860 ({i_8_, g734}, g732);
	defparam lut_8860.LUT_SIZE = 2;
	defparam lut_8860.mask = 4'b0001;

	lut_sub lut_8865 ({g95, i_9_}, g733);
	defparam lut_8865.LUT_SIZE = 2;
	defparam lut_8865.mask = 4'b1011;

	lut_sub lut_8874 ({g1, g68, g14, i_9_}, g734);
	defparam lut_8874.LUT_SIZE = 4;
	defparam lut_8874.mask = 16'hfbff;

	lut_sub lut_8894 ({g736, g737}, g735);
	defparam lut_8894.LUT_SIZE = 2;
	defparam lut_8894.mask = 4'b1000;

	lut_sub lut_8900 ({g45, g738}, g736);
	defparam lut_8900.LUT_SIZE = 2;
	defparam lut_8900.mask = 4'b0100;

	lut_sub lut_8906 ({g45, g741}, g737);
	defparam lut_8906.LUT_SIZE = 2;
	defparam lut_8906.mask = 4'b0001;

	lut_sub lut_8912 ({g739, g740}, g738);
	defparam lut_8912.LUT_SIZE = 2;
	defparam lut_8912.mask = 4'b1000;

	lut_sub lut_8917 ({i_9_, g744}, g739);
	defparam lut_8917.LUT_SIZE = 2;
	defparam lut_8917.mask = 4'b0100;

	lut_sub lut_8922 ({i_9_, g745}, g740);
	defparam lut_8922.LUT_SIZE = 2;
	defparam lut_8922.mask = 4'b0001;

	lut_sub lut_8928 ({g742, g743}, g741);
	defparam lut_8928.LUT_SIZE = 2;
	defparam lut_8928.mask = 4'b1000;

	lut_sub lut_8933 ({i_9_, g746}, g742);
	defparam lut_8933.LUT_SIZE = 2;
	defparam lut_8933.mask = 4'b0100;

	lut_sub lut_8938 ({i_9_, g229}, g743);
	defparam lut_8938.LUT_SIZE = 2;
	defparam lut_8938.mask = 4'b0001;

	lut_sub lut_8946 ({g10, g54, g1, g229}, g744);
	defparam lut_8946.LUT_SIZE = 4;
	defparam lut_8946.mask = 16'h1555;

	lut_sub lut_8959 ({g10, g39, g229}, g745);
	defparam lut_8959.LUT_SIZE = 3;
	defparam lut_8959.mask = 8'h45;

	lut_sub lut_8969 ({g10, g54, g1, g229}, g746);
	defparam lut_8969.LUT_SIZE = 4;
	defparam lut_8969.mask = 16'h1555;

	lut_sub lut_8981 ({g748, g749}, g747);
	defparam lut_8981.LUT_SIZE = 2;
	defparam lut_8981.mask = 4'b1000;

	lut_sub lut_8987 ({g133, g750}, g748);
	defparam lut_8987.LUT_SIZE = 2;
	defparam lut_8987.mask = 4'b0100;

	lut_sub lut_8993 ({g133, g753}, g749);
	defparam lut_8993.LUT_SIZE = 2;
	defparam lut_8993.mask = 4'b0001;

	lut_sub lut_8999 ({g751, g752}, g750);
	defparam lut_8999.LUT_SIZE = 2;
	defparam lut_8999.mask = 4'b1000;

	lut_sub lut_9004 ({i_8_, g755}, g751);
	defparam lut_9004.LUT_SIZE = 2;
	defparam lut_9004.mask = 4'b0100;

	lut_sub lut_9009 ({i_8_, g756}, g752);
	defparam lut_9009.LUT_SIZE = 2;
	defparam lut_9009.mask = 4'b0001;

	lut_sub lut_9014 ({i_8_, g754}, g753);
	defparam lut_9014.LUT_SIZE = 2;
	defparam lut_9014.mask = 4'b1000;

	lut_sub lut_9019 ({i_8_, g757}, g754);
	defparam lut_9019.LUT_SIZE = 2;
	defparam lut_9019.mask = 4'b0100;

	lut_sub lut_9024 ({i_7_, i_6_, g28}, g755);
	defparam lut_9024.LUT_SIZE = 3;
	defparam lut_9024.mask = 8'hf7;

	lut_sub lut_9036 ({i_7_, i_6_, g7, g28}, g756);
	defparam lut_9036.LUT_SIZE = 4;
	defparam lut_9036.mask = 16'hfc4f;

	lut_sub lut_9052 ({i_7_, i_6_, g13, g28}, g757);
	defparam lut_9052.LUT_SIZE = 4;
	defparam lut_9052.mask = 16'hff7f;

	lut_sub lut_9071 ({i_2_, g759}, g758);
	defparam lut_9071.LUT_SIZE = 2;
	defparam lut_9071.mask = 4'b0010;

	lut_sub lut_9076 ({i_2_, g760}, g759);
	defparam lut_9076.LUT_SIZE = 2;
	defparam lut_9076.mask = 4'b0001;

	lut_sub lut_9082 ({g761, g762}, g760);
	defparam lut_9082.LUT_SIZE = 2;
	defparam lut_9082.mask = 4'b1000;

	lut_sub lut_9087 ({i_1_, g763}, g761);
	defparam lut_9087.LUT_SIZE = 2;
	defparam lut_9087.mask = 4'b0100;

	lut_sub lut_9092 ({i_1_, g764}, g762);
	defparam lut_9092.LUT_SIZE = 2;
	defparam lut_9092.mask = 4'b0001;

	lut_sub lut_9097 ({i_9_, g37, i_0_}, g763);
	defparam lut_9097.LUT_SIZE = 3;
	defparam lut_9097.mask = 8'hbf;

	lut_sub lut_9109 ({g50, i_9_, g76, i_0_}, g764);
	defparam lut_9109.LUT_SIZE = 4;
	defparam lut_9109.mask = 16'hbfff;

	lut_sub lut_9129 ({g766, g767}, g765);
	defparam lut_9129.LUT_SIZE = 2;
	defparam lut_9129.mask = 4'b1000;

	lut_sub lut_9134 ({i_8_, g768}, g766);
	defparam lut_9134.LUT_SIZE = 2;
	defparam lut_9134.mask = 4'b0100;

	lut_sub lut_9139 ({i_8_, g770}, g767);
	defparam lut_9139.LUT_SIZE = 2;
	defparam lut_9139.mask = 4'b0001;

	lut_sub lut_9144 ({i_7_, g769}, g768);
	defparam lut_9144.LUT_SIZE = 2;
	defparam lut_9144.mask = 4'b1000;

	lut_sub lut_9149 ({i_7_, g772}, g769);
	defparam lut_9149.LUT_SIZE = 2;
	defparam lut_9149.mask = 4'b0100;

	lut_sub lut_9154 ({i_7_, g771}, g770);
	defparam lut_9154.LUT_SIZE = 2;
	defparam lut_9154.mask = 4'b0010;

	lut_sub lut_9159 ({i_7_, g773}, g771);
	defparam lut_9159.LUT_SIZE = 2;
	defparam lut_9159.mask = 4'b0001;

	lut_sub lut_9164 ({i_9_, g82, i_6_}, g772);
	defparam lut_9164.LUT_SIZE = 3;
	defparam lut_9164.mask = 8'hfe;

	lut_sub lut_9176 ({g11, i_9_, g7, i_6_}, g773);
	defparam lut_9176.LUT_SIZE = 4;
	defparam lut_9176.mask = 16'hfffe;

	lut_sub lut_9196 ({g775, g776}, g774);
	defparam lut_9196.LUT_SIZE = 2;
	defparam lut_9196.mask = 4'b1000;

	lut_sub lut_9202 ({g15, g777}, g775);
	defparam lut_9202.LUT_SIZE = 2;
	defparam lut_9202.mask = 4'b0100;

	lut_sub lut_9208 ({g15, g780}, g776);
	defparam lut_9208.LUT_SIZE = 2;
	defparam lut_9208.mask = 4'b0001;

	lut_sub lut_9214 ({g778, g779}, g777);
	defparam lut_9214.LUT_SIZE = 2;
	defparam lut_9214.mask = 4'b1000;

	lut_sub lut_9219 ({i_9_, g783}, g778);
	defparam lut_9219.LUT_SIZE = 2;
	defparam lut_9219.mask = 4'b0100;

	lut_sub lut_9224 ({i_9_, g784}, g779);
	defparam lut_9224.LUT_SIZE = 2;
	defparam lut_9224.mask = 4'b0001;

	lut_sub lut_9230 ({g781, g782}, g780);
	defparam lut_9230.LUT_SIZE = 2;
	defparam lut_9230.mask = 4'b1000;

	lut_sub lut_9235 ({i_9_, g785}, g781);
	defparam lut_9235.LUT_SIZE = 2;
	defparam lut_9235.mask = 4'b0100;

	lut_sub lut_9240 ({i_9_, g786}, g782);
	defparam lut_9240.LUT_SIZE = 2;
	defparam lut_9240.mask = 4'b0001;

	lut_sub lut_9245 ({i_1_, i_0_, g17, i_2_}, g783);
	defparam lut_9245.LUT_SIZE = 4;
	defparam lut_9245.mask = 16'hdfff;

	lut_sub lut_9264 ({i_1_, i_0_, g19, i_2_}, g784);
	defparam lut_9264.LUT_SIZE = 4;
	defparam lut_9264.mask = 16'hffef;

	lut_sub lut_9283 ({i_1_, i_0_, g17, i_2_}, g785);
	defparam lut_9283.LUT_SIZE = 4;
	defparam lut_9283.mask = 16'hdff5;

	lut_sub lut_9300 ({i_1_, i_0_, g19, i_2_}, g786);
	defparam lut_9300.LUT_SIZE = 4;
	defparam lut_9300.mask = 16'hffef;

	lut_sub lut_9320 ({g788, g789}, g787);
	defparam lut_9320.LUT_SIZE = 2;
	defparam lut_9320.mask = 4'b1000;

	lut_sub lut_9326 ({g1, g790}, g788);
	defparam lut_9326.LUT_SIZE = 2;
	defparam lut_9326.mask = 4'b0100;

	lut_sub lut_9332 ({g1, g793}, g789);
	defparam lut_9332.LUT_SIZE = 2;
	defparam lut_9332.mask = 4'b0001;

	lut_sub lut_9338 ({g791, g792}, g790);
	defparam lut_9338.LUT_SIZE = 2;
	defparam lut_9338.mask = 4'b1000;

	lut_sub lut_9343 ({i_9_, g796}, g791);
	defparam lut_9343.LUT_SIZE = 2;
	defparam lut_9343.mask = 4'b0100;

	lut_sub lut_9348 ({i_9_, g797}, g792);
	defparam lut_9348.LUT_SIZE = 2;
	defparam lut_9348.mask = 4'b0001;

	lut_sub lut_9354 ({g794, g795}, g793);
	defparam lut_9354.LUT_SIZE = 2;
	defparam lut_9354.mask = 4'b1000;

	lut_sub lut_9359 ({i_9_, g798}, g794);
	defparam lut_9359.LUT_SIZE = 2;
	defparam lut_9359.mask = 4'b0100;

	lut_sub lut_9364 ({i_9_, g799}, g795);
	defparam lut_9364.LUT_SIZE = 2;
	defparam lut_9364.mask = 4'b0001;

	lut_sub lut_9372 ({g6, g4, g9, g3}, g796);
	defparam lut_9372.LUT_SIZE = 4;
	defparam lut_9372.mask = 16'h4c5f;

	lut_sub lut_9386 ({g12, g3}, g797);
	defparam lut_9386.LUT_SIZE = 2;
	defparam lut_9386.mask = 4'b0111;

	lut_sub lut_9394 ({g6, g9}, g798);
	defparam lut_9394.LUT_SIZE = 2;
	defparam lut_9394.mask = 4'b1011;

	lut_sub lut_9402 ({g12, g3}, g799);
	defparam lut_9402.LUT_SIZE = 2;
	defparam lut_9402.mask = 4'b0111;


endmodule