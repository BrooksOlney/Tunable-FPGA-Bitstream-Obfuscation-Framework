module ks_spla_qmap_map (sk, i_0_, i_1_, i_8_, i_6_, i_7_, i_9_, i_10_, i_11_, i_15_, i_12_, i_13_, i_14_, i_4_, i_3_, i_5_, i_2_, o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_, o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_, o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_, o_41_, o_42_, o_43_, o_44_, o_45_);

	input i_0_;
	input i_1_;
	input i_8_;
	input i_6_;
	input i_7_;
	input i_9_;
	input i_10_;
	input i_11_;
	input i_15_;
	input i_12_;
	input i_13_;
	input i_14_;
	input i_4_;
	input i_3_;
	input i_5_;
	input i_2_;
	output o_0_;
	output o_1_;
	output o_2_;
	output o_3_;
	output o_4_;
	output o_5_;
	output o_6_;
	output o_7_;
	output o_8_;
	output o_9_;
	output o_10_;
	output o_11_;
	output o_12_;
	output o_13_;
	output o_14_;
	output o_15_;
	output o_16_;
	output o_17_;
	output o_18_;
	output o_19_;
	output o_20_;
	output o_21_;
	output o_22_;
	output o_23_;
	output o_24_;
	output o_25_;
	output o_26_;
	output o_27_;
	output o_28_;
	output o_29_;
	output o_30_;
	output o_31_;
	output o_32_;
	output o_33_;
	output o_34_;
	output o_35_;
	output o_36_;
	output o_37_;
	output o_38_;
	output o_39_;
	output o_40_;
	output o_41_;
	output o_42_;
	output o_43_;
	output o_44_;
	output o_45_;

	input [127 : 0] sk /* synthesis noprune */;


	wire g9, g11, g52, g456, g458, g621, g812, g845, g846, g923, g963, g989, g1003, g1456, g1018, g1057, g1454, g1077, g1125, g1128, g1129;
	wire g1253, g1346, g1393, g1417, g1422, g1424, g1426, g1437, g1449, g1451, g1, g2, g3, g4, g5, g6, g7, g8, g10, g12, g14;
	wire g15, g16, g17, g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29, g30, g31, g32, g33, g34, g35;
	wire g36, g37, g38, g39, g40, g41, g42, g43, g44, g45, g46, g47, g48, g49, g50, g51, g53, g54, g55, g56, g57;
	wire g58, g59, g60, g61, g62, g63, g64, g65, g66, g68, g69, g70, g71, g72, g73, g74, g75, g76, g77, g78, g79;
	wire g80, g81, g82, g83, g84, g85, g86, g87, g88, g89, g90, g91, g92, g93, g94, g95, g96, g97, g98, g99, g100;
	wire g101, g102, g103, g104, g105, g106, g107, g108, g109, g110, g111, g112, g113, g114, g115, g116, g117, g118, g119, g120, g121;
	wire g122, g123, g124, g125, g126, g127, g128, g129, g130, g131, g1639, g132, g133, g134, g135, g136, g137, g138, g139, g140, g141;
	wire g142, g143, g144, g145, g146, g147, g148, g149, g150, g151, g152, g153, g154, g155, g156, g157, g158, g159, g160, g161, g162;
	wire g163, g164, g165, g166, g167, g168, g169, g170, g171, g172, g173, g174, g175, g176, g177, g178, g179, g180, g181, g182, g183;
	wire g184, g185, g186, g187, g188, g189, g190, g191, g192, g193, g194, g195, g196, g197, g198, g199, g200, g201, g202, g203, g204;
	wire g205, g206, g207, g208, g209, g210, g211, g212, g213, g214, g215, g216, g217, g218, g219, g220, g221, g222, g223, g224, g225;
	wire g226, g227, g228, g229, g230, g231, g232, g233, g234, g235, g236, g237, g238, g239, g240, g241, g242, g243, g244, g245, g246;
	wire g247, g248, g249, g250, g251, g252, g253, g254, g255, g256, g257, g258, g259, g260, g261, g262, g263, g264, g265, g266, g267;
	wire g268, g269, g270, g271, g272, g273, g274, g275, g276, g277, g278, g279, g280, g281, g282, g283, g284, g285, g286, g287, g288;
	wire g289, g290, g291, g292, g293, g294, g295, g296, g297, g298, g299, g300, g301, g302, g303, g304, g305, g306, g307, g308, g309;
	wire g310, g311, g312, g313, g314, g315, g1632, g316, g317, g318, g319, g320, g1625, g321, g322, g323, g324, g325, g326, g327, g328;
	wire g329, g330, g1606, g331, g1613, g332, g333, g334, g335, g336, g337, g338, g339, g340, g341, g342, g343, g344, g345, g346, g347;
	wire g348, g349, g350, g351, g352, g353, g354, g355, g356, g357, g358, g359, g360, g361, g362, g363, g364, g365, g366, g367, g368;
	wire g369, g370, g371, g372, g373, g374, g375, g376, g377, g378, g379, g380, g381, g382, g383, g384, g385, g386, g387, g388, g389;
	wire g390, g391, g392, g393, g394, g395, g396, g397, g398, g399, g400, g401, g402, g403, g404, g405, g406, g407, g408, g409, g410;
	wire g411, g412, g413, g414, g415, g416, g417, g418, g419, g420, g421, g422, g423, g424, g425, g426, g427, g428, g429, g430, g431;
	wire g432, g433, g434, g435, g436, g437, g438, g439, g440, g441, g1593, g442, g443, g444, g445, g446, g447, g448, g449, g450, g451;
	wire g452, g453, g454, g1584, g455, g457, g459, g460, g461, g462, g463, g464, g465, g466, g467, g468, g469, g470, g471, g472, g473;
	wire g474, g475, g476, g477, g478, g479, g480, g481, g482, g483, g484, g485, g486, g487, g488, g489, g490, g491, g492, g493, g494;
	wire g495, g496, g497, g498, g499, g500, g501, g502, g503, g504, g505, g506, g507, g508, g509, g510, g511, g512, g513, g514, g515;
	wire g516, g517, g518, g1577, g519, g520, g521, g522, g523, g524, g1564, g525, g526, g527, g528, g529, g530, g531, g532, g533, g534;
	wire g535, g536, g1459, g537, g538, g539, g540, g541, g542, g543, g544, g545, g546, g547, g548, g549, g550, g551, g552, g553, g554;
	wire g555, g556, g557, g558, g559, g560, g561, g562, g563, g564, g565, g566, g567, g568, g569, g570, g571, g572, g573, g574, g575;
	wire g576, g577, g578, g579, g580, g1554, g1543, g581, g582, g583, g584, g585, g586, g587, g588, g589, g590, g591, g592, g593, g594;
	wire g595, g596, g597, g598, g599, g600, g601, g602, g603, g604, g605, g606, g607, g608, g609, g610, g611, g612, g613, g614, g615;
	wire g616, g617, g618, g1458, g619, g620, g623, g624, g625, g626, g627, g628, g629, g630, g631, g632, g633, g634, g635, g636, g637;
	wire g638, g639, g640, g641, g642, g643, g644, g645, g646, g647, g648, g649, g650, g651, g652, g653, g654, g655, g656, g657, g658;
	wire g659, g660, g661, g662, g663, g664, g665, g666, g667, g668, g669, g670, g671, g672, g673, g674, g675, g676, g677, g678, g679;
	wire g680, g681, g682, g683, g684, g685, g686, g687, g688, g689, g690, g1457, g691, g692, g693, g694, g695, g696, g697, g698, g699;
	wire g700, g701, g702, g703, g704, g705, g706, g1531, g707, g708, g709, g710, g711, g712, g713, g714, g715, g716, g717, g718, g719;
	wire g720, g721, g722, g723, g724, g725, g726, g727, g728, g729, g730, g731, g732, g733, g734, g735, g736, g737, g738, g739, g740;
	wire g741, g742, g743, g744, g745, g746, g747, g1518, g748, g749, g750, g751, g752, g753, g754, g755, g756, g757, g758, g759, g760;
	wire g761, g762, g763, g764, g765, g766, g767, g768, g769, g770, g771, g772, g773, g774, g775, g776, g777, g778, g779, g780, g781;
	wire g782, g783, g784, g785, g786, g787, g788, g789, g790, g791, g792, g793, g794, g795, g796, g797, g798, g799, g800, g801, g802;
	wire g803, g804, g805, g806, g807, g808, g809, g810, g811, g813, g814, g815, g816, g817, g818, g819, g820, g821, g822, g823, g824;
	wire g825, g826, g827, g828, g829, g830, g831, g832, g833, g834, g835, g836, g837, g838, g839, g840, g841, g842, g843, g1511, g844;
	wire g847, g848, g849, g850, g851, g852, g853, g854, g855, g856, g857, g858, g859, g860, g861, g862, g863, g864, g865, g866, g867;
	wire g868, g869, g870, g871, g872, g1501, g1488, g873, g874, g875, g876, g877, g878, g879, g880, g881, g882, g883, g884, g885, g886;
	wire g887, g888, g889, g890, g891, g892, g893, g894, g895, g896, g1478, g897, g898, g899, g900, g901, g902, g903, g904, g905, g906;
	wire g907, g908, g909, g910, g911, g912, g913, g914, g915, g916, g917, g918, g919, g920, g921, g922, g924, g925, g926, g927, g928;
	wire g929, g930, g931, g932, g933, g934, g935, g936, g937, g938, g939, g940, g941, g942, g943, g944, g945, g946, g947, g948, g949;
	wire g950, g1467, g951, g952, g953, g954, g955, g956, g957, g958, g959, g960, g961, g962, g964, g965, g966, g967, g968, g969, g970;
	wire g971, g972, g973, g974, g975, g976, g977, g978, g979, g980, g981, g982, g983, g984, g985, g986, g987, g988, g990, g991, g992;
	wire g993, g994, g995, g996, g997, g998, g999, g1000, g1001, g1002, g1004, g1005, g1006, g1007, g1008, g1009, g1010, g1011, g1012, g1013, g1455;
	wire g1014, g1015, g1016, g1017, g1019, g1020, g1021, g1022, g1023, g1024, g1025, g1026, g1027, g1028, g1029, g1030, g1031, g1032, g1033, g1034, g1035;
	wire g1036, g1037, g1038, g1039, g1040, g1041, g1042, g1043, g1044, g1045, g1046, g1047, g1048, g1049, g1050, g1051, g1052, g1053, g1054, g1055, g1056;
	wire g1058, g1060, g1062, g1063, g1064, g1065, g1067, g1068, g1069, g1070, g1071, g1072, g1073, g1074, g1075, g1076, g1080, g1081, g1082, g1084, g1085;
	wire g1086, g1087, g1088, g1090, g1091, g1094, g1095, g1096, g1097, g1098, g1099, g1100, g1101, g1102, g1103, g1104, g1105, g1106, g1107, g1108, g1109;
	wire g1110, g1111, g1112, g1460, g1113, g1114, g1115, g1116, g1117, g1118, g1119, g1122, g1123, g1124, g1126, g1127, g1130, g1131, g1132, g1133, g1134;
	wire g1135, g1136, g1137, g1138, g1139, g1140, g1141, g1142, g1143, g1144, g1145, g1146, g1147, g1148, g1149, g1150, g1151, g1152, g1153, g1154, g1155;
	wire g1156, g1157, g1158, g1159, g1160, g1161, g1162, g1163, g1164, g1165, g1166, g1167, g1168, g1169, g1170, g1171, g1172, g1173, g1174, g1175, g1176;
	wire g1177, g1178, g1179, g1180, g1181, g1182, g1453, g1183, g1184, g1185, g1186, g1452, g1187, g1188, g1189, g1190, g1191, g1192, g1193, g1194, g1195;
	wire g1196, g1197, g1198, g1199, g1200, g1201, g1202, g1203, g1204, g1205, g1206, g1207, g1208, g1209, g1210, g1211, g1212, g1213, g1214, g1215, g1216;
	wire g1217, g1218, g1219, g1220, g1221, g1222, g1223, g1224, g1225, g1226, g1227, g1228, g1229, g1230, g1231, g1232, g1233, g1234, g1235, g1236, g1237;
	wire g1238, g1239, g1240, g1241, g1242, g1243, g1244, g1245, g1246, g1247, g1248, g1249, g1250, g1251, g1252, g1254, g1255, g1256, g1257, g1258, g1259;
	wire g1260, g1261, g1262, g1263, g1264, g1265, g1266, g1267, g1268, g1269, g1270, g1271, g1272, g1273, g1274, g1275, g1276, g1277, g1278, g1279, g1280;
	wire g1281, g1282, g1283, g1284, g1285, g1286, g1287, g1288, g1289, g1290, g1291, g1292, g1293, g1294, g1295, g1296, g1297, g1298, g1299, g1300, g1301;
	wire g1302, g1303, g1304, g1305, g1306, g1307, g1308, g1309, g1310, g1311, g1312, g1313, g1314, g1315, g1316, g1317, g1318, g1319, g1320, g1321, g1322;
	wire g1323, g1324, g1325, g1326, g1327, g1328, g1329, g1330, g1331, g1332, g1333, g1334, g1335, g1336, g1337, g1338, g1339, g1340, g1341, g1342, g1343;
	wire g1344, g1345, g1347, g1348, g1349, g1350, g1351, g1352, g1353, g1354, g1355, g1356, g1357, g1358, g1359, g1360, g1361, g1362, g1363, g1364, g1365;
	wire g1366, g1367, g1368, g1369, g1370, g1371, g1372, g1373, g1374, g1375, g1376, g1377, g1378, g1379, g1380, g1381, g1382, g1383, g1384, g1385, g1386;
	wire g1387, g1388, g1389, g1390, g1391, g1392, g1394, g1395, g1396, g1397, g1398, g1399, g1400, g1401, g1402, g1403, g1404, g1405, g1406, g1407, g1408;
	wire g1409, g1410, g1411, g1412, g1413, g1414, g1415, g1416, g1418, g1419, g1420, g1421, g1423, g1427, g1428, g1429, g1430, g1431, g1432, g1433, g1434;
	wire g1435, g1436, g1438, g1439, g1440, g1441, g1442, g1443, g1444, g1445, g1446, g1447, g1448, g1450, g1461, g1462, g1463, g1464, g1465, g1466, g1468;
	wire g1469, g1470, g1472, g1471, g1475, g1473, g1474, g1476, g1477, g1479, g1480, g1481, g1482, g1485, g1483, g1484, g1486, g1487, g1489, g1490, g1491;
	wire g1494, g1492, g1493, g1497, g1498, g1495, g1496, g1499, g1500, g1502, g1503, g1504, g1505, g1508, g1506, g1507, g1509, g1510, g1512, g1513, g1514;
	wire g1515, g1516, g1517, g1519, g1520, g1521, g1524, g1522, g1523, g1527, g1528, g1525, g1526, g1529, g1530, g1532, g1533, g1534, g1537, g1535, g1536;
	wire g1540, g1538, g1539, g1541, g1542, g1544, g1545, g1546, g1549, g1547, g1548, g1550, g1551, g1552, g1553, g1555, g1556, g1557, g1558, g1561, g1559;
	wire g1560, g1562, g1563, g1565, g1566, g1567, g1570, g1568, g1569, g1573, g1574, g1571, g1572, g1575, g1576, g1578, g1579, g1580, g1581, g1582, g1583;
	wire g1585, g1586, g1587, g1589, g1588, g1591, g1590, g1592, g1594, g1595, g1596, g1599, g1597, g1598, g1602, g1603, g1600, g1601, g1604, g1605, g1607;
	wire g1608, g1609, g1610, g1611, g1612, g1614, g1615, g1616, g1619, g1617, g1618, g1622, g1623, g1620, g1621, g1624, g1626, g1627, g1628, g1629, g1630;
	wire g1631, g1633, g1634, g1635, g1636, g1637, g1638, g1640, g1641, g1642, g1643, g1646, g1644, g1645, g1647, g1648;

	assign o_0_ = (((sk[0]) & (!g9)));
	assign o_1_ = (((sk[1]) & (!g11)));
	assign o_3_ = (((sk[2]) & (!g52)));
	assign o_5_ = (((sk[3]) & (!g456)));
	assign o_6_ = (((sk[4]) & (!g458)));
	assign o_7_ = (((sk[5]) & (!g621)));
	assign o_9_ = (((sk[6]) & (!g812)));
	assign o_10_ = (((sk[7]) & (!g845)));
	assign o_11_ = (((sk[8]) & (!g846)));
	assign o_12_ = (((sk[9]) & (!g923)));
	assign o_13_ = (((sk[10]) & (!g963)));
	assign o_14_ = (((sk[11]) & (!g989)));
	assign o_15_ = (((sk[12]) & (!g1003)));
	assign o_16_ = (((sk[13]) & (!g1456)));
	assign o_17_ = (((sk[14]) & (!g1018)));
	assign o_18_ = (((sk[15]) & (!g1057)));
	assign o_22_ = (((sk[16]) & (!g1454)));
	assign o_23_ = (((sk[17]) & (!g1077)));
	assign o_32_ = (((sk[18]) & (!g1125)));
	assign o_33_ = (((sk[19]) & (!g1128)));
	assign o_34_ = (((sk[20]) & (!g1129)));
	assign o_35_ = (((sk[21]) & (!g1253)));
	assign o_36_ = (((sk[22]) & (!g1346)));
	assign o_37_ = (((sk[23]) & (!g1393)));
	assign o_38_ = (((sk[24]) & (!g1417)));
	assign o_39_ = (((sk[25]) & (!g1422)));
	assign o_40_ = (((sk[26]) & (!g1424)));
	assign o_42_ = (((sk[27]) & (!g1426)));
	assign o_43_ = (((sk[28]) & (!g1437)));
	assign o_44_ = (((sk[29]) & (!g1449)));
	assign o_45_ = (((sk[30]) & (!g1451)));
	assign g1 = (((!sk[31]) & (i_6_) & (!i_7_)) + ((!sk[31]) & (i_6_) & (i_7_)) + ((sk[31]) & (!i_6_) & (!i_7_)));
	assign g2 = (((!i_8_) & (sk[32]) & (g1)) + ((i_8_) & (!sk[32]) & (!g1)) + ((i_8_) & (!sk[32]) & (g1)));
	assign g3 = (((!i_9_) & (!sk[33]) & (!i_10_) & (i_11_) & (!i_15_)) + ((!i_9_) & (!sk[33]) & (!i_10_) & (i_11_) & (i_15_)) + ((!i_9_) & (!sk[33]) & (i_10_) & (!i_11_) & (i_15_)) + ((!i_9_) & (!sk[33]) & (i_10_) & (i_11_) & (!i_15_)) + ((!i_9_) & (!sk[33]) & (i_10_) & (i_11_) & (i_15_)) + ((!i_9_) & (sk[33]) & (!i_10_) & (!i_11_) & (!i_15_)) + ((i_9_) & (!sk[33]) & (!i_10_) & (!i_11_) & (!i_15_)) + ((i_9_) & (!sk[33]) & (!i_10_) & (!i_11_) & (i_15_)) + ((i_9_) & (!sk[33]) & (!i_10_) & (i_11_) & (!i_15_)) + ((i_9_) & (!sk[33]) & (!i_10_) & (i_11_) & (i_15_)) + ((i_9_) & (!sk[33]) & (i_10_) & (!i_11_) & (!i_15_)) + ((i_9_) & (!sk[33]) & (i_10_) & (!i_11_) & (i_15_)) + ((i_9_) & (!sk[33]) & (i_10_) & (i_11_) & (!i_15_)) + ((i_9_) & (!sk[33]) & (i_10_) & (i_11_) & (i_15_)));
	assign g4 = (((!i_12_) & (sk[34]) & (!i_13_) & (!i_14_)) + ((i_12_) & (!sk[34]) & (!i_13_) & (!i_14_)) + ((i_12_) & (!sk[34]) & (!i_13_) & (i_14_)) + ((i_12_) & (!sk[34]) & (i_13_) & (!i_14_)) + ((i_12_) & (!sk[34]) & (i_13_) & (i_14_)));
	assign g5 = (((!sk[35]) & (g3) & (!g4)) + ((!sk[35]) & (g3) & (g4)) + ((sk[35]) & (g3) & (g4)));
	assign g6 = (((!i_4_) & (sk[36]) & (!i_3_) & (i_5_)) + ((i_4_) & (!sk[36]) & (!i_3_) & (!i_5_)) + ((i_4_) & (!sk[36]) & (!i_3_) & (i_5_)) + ((i_4_) & (!sk[36]) & (i_3_) & (!i_5_)) + ((i_4_) & (!sk[36]) & (i_3_) & (i_5_)));
	assign g7 = (((!i_0_) & (!i_1_) & (g6) & (!sk[37]) & (!i_2_)) + ((!i_0_) & (!i_1_) & (g6) & (!sk[37]) & (i_2_)) + ((!i_0_) & (i_1_) & (!g6) & (!sk[37]) & (i_2_)) + ((!i_0_) & (i_1_) & (g6) & (!sk[37]) & (!i_2_)) + ((!i_0_) & (i_1_) & (g6) & (!sk[37]) & (i_2_)) + ((i_0_) & (!i_1_) & (!g6) & (!sk[37]) & (!i_2_)) + ((i_0_) & (!i_1_) & (!g6) & (!sk[37]) & (i_2_)) + ((i_0_) & (!i_1_) & (g6) & (!sk[37]) & (!i_2_)) + ((i_0_) & (!i_1_) & (g6) & (!sk[37]) & (i_2_)) + ((i_0_) & (i_1_) & (!g6) & (!sk[37]) & (!i_2_)) + ((i_0_) & (i_1_) & (!g6) & (!sk[37]) & (i_2_)) + ((i_0_) & (i_1_) & (g6) & (!sk[37]) & (!i_2_)) + ((i_0_) & (i_1_) & (g6) & (!sk[37]) & (i_2_)) + ((i_0_) & (i_1_) & (g6) & (sk[37]) & (!i_2_)));
	assign g8 = (((!sk[38]) & (g5) & (!g7)) + ((!sk[38]) & (g5) & (g7)) + ((sk[38]) & (g5) & (g7)));
	assign g9 = (((!i_0_) & (!i_1_) & (!sk[39]) & (g2) & (!g8)) + ((!i_0_) & (!i_1_) & (!sk[39]) & (g2) & (g8)) + ((!i_0_) & (!i_1_) & (sk[39]) & (!g2) & (!g8)) + ((!i_0_) & (!i_1_) & (sk[39]) & (!g2) & (g8)) + ((!i_0_) & (!i_1_) & (sk[39]) & (g2) & (!g8)) + ((!i_0_) & (i_1_) & (!sk[39]) & (!g2) & (g8)) + ((!i_0_) & (i_1_) & (!sk[39]) & (g2) & (!g8)) + ((!i_0_) & (i_1_) & (!sk[39]) & (g2) & (g8)) + ((!i_0_) & (i_1_) & (sk[39]) & (!g2) & (!g8)) + ((!i_0_) & (i_1_) & (sk[39]) & (!g2) & (g8)) + ((!i_0_) & (i_1_) & (sk[39]) & (g2) & (!g8)) + ((i_0_) & (!i_1_) & (!sk[39]) & (!g2) & (!g8)) + ((i_0_) & (!i_1_) & (!sk[39]) & (!g2) & (g8)) + ((i_0_) & (!i_1_) & (!sk[39]) & (g2) & (!g8)) + ((i_0_) & (!i_1_) & (!sk[39]) & (g2) & (g8)) + ((i_0_) & (i_1_) & (!sk[39]) & (!g2) & (!g8)) + ((i_0_) & (i_1_) & (!sk[39]) & (!g2) & (g8)) + ((i_0_) & (i_1_) & (!sk[39]) & (g2) & (!g8)) + ((i_0_) & (i_1_) & (!sk[39]) & (g2) & (g8)) + ((i_0_) & (i_1_) & (sk[39]) & (!g2) & (!g8)) + ((i_0_) & (i_1_) & (sk[39]) & (!g2) & (g8)) + ((i_0_) & (i_1_) & (sk[39]) & (g2) & (!g8)));
	assign g10 = (((!sk[40]) & (i_6_) & (!i_7_)) + ((!sk[40]) & (i_6_) & (i_7_)) + ((sk[40]) & (!i_6_) & (i_7_)));
	assign g11 = (((!i_0_) & (!i_1_) & (!i_8_) & (!i_2_) & (!g8) & (!g10)) + ((!i_0_) & (!i_1_) & (!i_8_) & (!i_2_) & (!g8) & (g10)) + ((!i_0_) & (!i_1_) & (!i_8_) & (!i_2_) & (g8) & (!g10)) + ((!i_0_) & (!i_1_) & (i_8_) & (!i_2_) & (!g8) & (!g10)) + ((!i_0_) & (!i_1_) & (i_8_) & (!i_2_) & (!g8) & (g10)) + ((!i_0_) & (!i_1_) & (i_8_) & (!i_2_) & (g8) & (!g10)) + ((!i_0_) & (!i_1_) & (i_8_) & (!i_2_) & (g8) & (g10)) + ((!i_0_) & (i_1_) & (!i_8_) & (!i_2_) & (!g8) & (!g10)) + ((!i_0_) & (i_1_) & (!i_8_) & (!i_2_) & (!g8) & (g10)) + ((!i_0_) & (i_1_) & (!i_8_) & (!i_2_) & (g8) & (!g10)) + ((!i_0_) & (i_1_) & (i_8_) & (!i_2_) & (!g8) & (!g10)) + ((!i_0_) & (i_1_) & (i_8_) & (!i_2_) & (!g8) & (g10)) + ((!i_0_) & (i_1_) & (i_8_) & (!i_2_) & (g8) & (!g10)) + ((!i_0_) & (i_1_) & (i_8_) & (!i_2_) & (g8) & (g10)) + ((i_0_) & (!i_1_) & (!i_8_) & (i_2_) & (!g8) & (!g10)) + ((i_0_) & (!i_1_) & (!i_8_) & (i_2_) & (!g8) & (g10)) + ((i_0_) & (!i_1_) & (!i_8_) & (i_2_) & (g8) & (!g10)) + ((i_0_) & (!i_1_) & (i_8_) & (i_2_) & (!g8) & (!g10)) + ((i_0_) & (!i_1_) & (i_8_) & (i_2_) & (!g8) & (g10)) + ((i_0_) & (!i_1_) & (i_8_) & (i_2_) & (g8) & (!g10)) + ((i_0_) & (!i_1_) & (i_8_) & (i_2_) & (g8) & (g10)) + ((i_0_) & (i_1_) & (!i_8_) & (!i_2_) & (!g8) & (!g10)) + ((i_0_) & (i_1_) & (!i_8_) & (!i_2_) & (!g8) & (g10)) + ((i_0_) & (i_1_) & (!i_8_) & (!i_2_) & (g8) & (!g10)) + ((i_0_) & (i_1_) & (!i_8_) & (i_2_) & (!g8) & (!g10)) + ((i_0_) & (i_1_) & (!i_8_) & (i_2_) & (!g8) & (g10)) + ((i_0_) & (i_1_) & (!i_8_) & (i_2_) & (g8) & (!g10)) + ((i_0_) & (i_1_) & (i_8_) & (!i_2_) & (!g8) & (!g10)) + ((i_0_) & (i_1_) & (i_8_) & (!i_2_) & (!g8) & (g10)) + ((i_0_) & (i_1_) & (i_8_) & (!i_2_) & (g8) & (!g10)) + ((i_0_) & (i_1_) & (i_8_) & (!i_2_) & (g8) & (g10)) + ((i_0_) & (i_1_) & (i_8_) & (i_2_) & (!g8) & (!g10)) + ((i_0_) & (i_1_) & (i_8_) & (i_2_) & (!g8) & (g10)) + ((i_0_) & (i_1_) & (i_8_) & (i_2_) & (g8) & (!g10)) + ((i_0_) & (i_1_) & (i_8_) & (i_2_) & (g8) & (g10)));
	assign g12 = (((!i_0_) & (!i_1_) & (!sk[42]) & (g5) & (!i_2_)) + ((!i_0_) & (!i_1_) & (!sk[42]) & (g5) & (i_2_)) + ((!i_0_) & (i_1_) & (!sk[42]) & (!g5) & (i_2_)) + ((!i_0_) & (i_1_) & (!sk[42]) & (g5) & (!i_2_)) + ((!i_0_) & (i_1_) & (!sk[42]) & (g5) & (i_2_)) + ((i_0_) & (!i_1_) & (!sk[42]) & (!g5) & (!i_2_)) + ((i_0_) & (!i_1_) & (!sk[42]) & (!g5) & (i_2_)) + ((i_0_) & (!i_1_) & (!sk[42]) & (g5) & (!i_2_)) + ((i_0_) & (!i_1_) & (!sk[42]) & (g5) & (i_2_)) + ((i_0_) & (i_1_) & (!sk[42]) & (!g5) & (!i_2_)) + ((i_0_) & (i_1_) & (!sk[42]) & (!g5) & (i_2_)) + ((i_0_) & (i_1_) & (!sk[42]) & (g5) & (!i_2_)) + ((i_0_) & (i_1_) & (!sk[42]) & (g5) & (i_2_)) + ((i_0_) & (i_1_) & (sk[42]) & (g5) & (!i_2_)));
	assign o_2_ = (((!i_8_) & (!i_6_) & (!sk[43]) & (g6) & (!g12)) + ((!i_8_) & (!i_6_) & (!sk[43]) & (g6) & (g12)) + ((!i_8_) & (!i_6_) & (sk[43]) & (g6) & (g12)) + ((!i_8_) & (i_6_) & (!sk[43]) & (!g6) & (g12)) + ((!i_8_) & (i_6_) & (!sk[43]) & (g6) & (!g12)) + ((!i_8_) & (i_6_) & (!sk[43]) & (g6) & (g12)) + ((i_8_) & (!i_6_) & (!sk[43]) & (!g6) & (!g12)) + ((i_8_) & (!i_6_) & (!sk[43]) & (!g6) & (g12)) + ((i_8_) & (!i_6_) & (!sk[43]) & (g6) & (!g12)) + ((i_8_) & (!i_6_) & (!sk[43]) & (g6) & (g12)) + ((i_8_) & (i_6_) & (!sk[43]) & (!g6) & (!g12)) + ((i_8_) & (i_6_) & (!sk[43]) & (!g6) & (g12)) + ((i_8_) & (i_6_) & (!sk[43]) & (g6) & (!g12)) + ((i_8_) & (i_6_) & (!sk[43]) & (g6) & (g12)));
	assign g14 = (((!i_0_) & (i_1_) & (sk[44]) & (!i_2_)) + ((i_0_) & (!i_1_) & (!sk[44]) & (!i_2_)) + ((i_0_) & (!i_1_) & (!sk[44]) & (i_2_)) + ((i_0_) & (i_1_) & (!sk[44]) & (!i_2_)) + ((i_0_) & (i_1_) & (!sk[44]) & (i_2_)));
	assign g15 = (((!i_4_) & (sk[45]) & (!i_3_) & (!i_5_)) + ((i_4_) & (!sk[45]) & (!i_3_) & (!i_5_)) + ((i_4_) & (!sk[45]) & (!i_3_) & (i_5_)) + ((i_4_) & (!sk[45]) & (i_3_) & (!i_5_)) + ((i_4_) & (!sk[45]) & (i_3_) & (i_5_)));
	assign g16 = (((g14) & (!sk[46]) & (!g15)) + ((g14) & (!sk[46]) & (g15)) + ((g14) & (sk[46]) & (g15)));
	assign g17 = (((!i_9_) & (!i_10_) & (!sk[47]) & (i_11_) & (!i_15_)) + ((!i_9_) & (!i_10_) & (!sk[47]) & (i_11_) & (i_15_)) + ((!i_9_) & (i_10_) & (!sk[47]) & (!i_11_) & (i_15_)) + ((!i_9_) & (i_10_) & (!sk[47]) & (i_11_) & (!i_15_)) + ((!i_9_) & (i_10_) & (!sk[47]) & (i_11_) & (i_15_)) + ((i_9_) & (!i_10_) & (!sk[47]) & (!i_11_) & (!i_15_)) + ((i_9_) & (!i_10_) & (!sk[47]) & (!i_11_) & (i_15_)) + ((i_9_) & (!i_10_) & (!sk[47]) & (i_11_) & (!i_15_)) + ((i_9_) & (!i_10_) & (!sk[47]) & (i_11_) & (i_15_)) + ((i_9_) & (!i_10_) & (sk[47]) & (!i_11_) & (i_15_)) + ((i_9_) & (i_10_) & (!sk[47]) & (!i_11_) & (!i_15_)) + ((i_9_) & (i_10_) & (!sk[47]) & (!i_11_) & (i_15_)) + ((i_9_) & (i_10_) & (!sk[47]) & (i_11_) & (!i_15_)) + ((i_9_) & (i_10_) & (!sk[47]) & (i_11_) & (i_15_)));
	assign g18 = (((!sk[48]) & (g4) & (!g17)) + ((!sk[48]) & (g4) & (g17)) + ((sk[48]) & (g4) & (g17)));
	assign g19 = (((!i_12_) & (sk[49]) & (i_13_) & (!i_14_)) + ((i_12_) & (!sk[49]) & (!i_13_) & (!i_14_)) + ((i_12_) & (!sk[49]) & (!i_13_) & (i_14_)) + ((i_12_) & (!sk[49]) & (i_13_) & (!i_14_)) + ((i_12_) & (!sk[49]) & (i_13_) & (i_14_)));
	assign g20 = (((!sk[50]) & (!i_9_) & (!i_10_) & (i_11_) & (!i_15_)) + ((!sk[50]) & (!i_9_) & (!i_10_) & (i_11_) & (i_15_)) + ((!sk[50]) & (!i_9_) & (i_10_) & (!i_11_) & (i_15_)) + ((!sk[50]) & (!i_9_) & (i_10_) & (i_11_) & (!i_15_)) + ((!sk[50]) & (!i_9_) & (i_10_) & (i_11_) & (i_15_)) + ((!sk[50]) & (i_9_) & (!i_10_) & (!i_11_) & (!i_15_)) + ((!sk[50]) & (i_9_) & (!i_10_) & (!i_11_) & (i_15_)) + ((!sk[50]) & (i_9_) & (!i_10_) & (i_11_) & (!i_15_)) + ((!sk[50]) & (i_9_) & (!i_10_) & (i_11_) & (i_15_)) + ((!sk[50]) & (i_9_) & (i_10_) & (!i_11_) & (!i_15_)) + ((!sk[50]) & (i_9_) & (i_10_) & (!i_11_) & (i_15_)) + ((!sk[50]) & (i_9_) & (i_10_) & (i_11_) & (!i_15_)) + ((!sk[50]) & (i_9_) & (i_10_) & (i_11_) & (i_15_)) + ((sk[50]) & (!i_9_) & (i_10_) & (!i_11_) & (!i_15_)));
	assign g21 = (((!sk[51]) & (g19) & (!g20)) + ((!sk[51]) & (g19) & (g20)) + ((sk[51]) & (g19) & (g20)));
	assign g22 = (((!i_9_) & (!i_10_) & (!sk[52]) & (i_11_) & (!i_15_)) + ((!i_9_) & (!i_10_) & (!sk[52]) & (i_11_) & (i_15_)) + ((!i_9_) & (!i_10_) & (sk[52]) & (!i_11_) & (!i_15_)) + ((!i_9_) & (!i_10_) & (sk[52]) & (!i_11_) & (i_15_)) + ((!i_9_) & (!i_10_) & (sk[52]) & (i_11_) & (!i_15_)) + ((!i_9_) & (!i_10_) & (sk[52]) & (i_11_) & (i_15_)) + ((!i_9_) & (i_10_) & (!sk[52]) & (!i_11_) & (i_15_)) + ((!i_9_) & (i_10_) & (!sk[52]) & (i_11_) & (!i_15_)) + ((!i_9_) & (i_10_) & (!sk[52]) & (i_11_) & (i_15_)) + ((!i_9_) & (i_10_) & (sk[52]) & (!i_11_) & (!i_15_)) + ((!i_9_) & (i_10_) & (sk[52]) & (i_11_) & (!i_15_)) + ((!i_9_) & (i_10_) & (sk[52]) & (i_11_) & (i_15_)) + ((i_9_) & (!i_10_) & (!sk[52]) & (!i_11_) & (!i_15_)) + ((i_9_) & (!i_10_) & (!sk[52]) & (!i_11_) & (i_15_)) + ((i_9_) & (!i_10_) & (!sk[52]) & (i_11_) & (!i_15_)) + ((i_9_) & (!i_10_) & (!sk[52]) & (i_11_) & (i_15_)) + ((i_9_) & (!i_10_) & (sk[52]) & (!i_11_) & (!i_15_)) + ((i_9_) & (!i_10_) & (sk[52]) & (!i_11_) & (i_15_)) + ((i_9_) & (!i_10_) & (sk[52]) & (i_11_) & (!i_15_)) + ((i_9_) & (!i_10_) & (sk[52]) & (i_11_) & (i_15_)) + ((i_9_) & (i_10_) & (!sk[52]) & (!i_11_) & (!i_15_)) + ((i_9_) & (i_10_) & (!sk[52]) & (!i_11_) & (i_15_)) + ((i_9_) & (i_10_) & (!sk[52]) & (i_11_) & (!i_15_)) + ((i_9_) & (i_10_) & (!sk[52]) & (i_11_) & (i_15_)) + ((i_9_) & (i_10_) & (sk[52]) & (!i_11_) & (!i_15_)) + ((i_9_) & (i_10_) & (sk[52]) & (!i_11_) & (i_15_)) + ((i_9_) & (i_10_) & (sk[52]) & (i_11_) & (!i_15_)) + ((i_9_) & (i_10_) & (sk[52]) & (i_11_) & (i_15_)));
	assign g23 = (((!g4) & (sk[53]) & (!g22)) + ((!g4) & (sk[53]) & (g22)) + ((g4) & (!sk[53]) & (!g22)) + ((g4) & (!sk[53]) & (g22)) + ((g4) & (sk[53]) & (g22)));
	assign g24 = (((!sk[54]) & (i_12_) & (!i_13_) & (!i_14_)) + ((!sk[54]) & (i_12_) & (!i_13_) & (i_14_)) + ((!sk[54]) & (i_12_) & (i_13_) & (!i_14_)) + ((!sk[54]) & (i_12_) & (i_13_) & (i_14_)) + ((sk[54]) & (!i_12_) & (!i_13_) & (!i_14_)) + ((sk[54]) & (!i_12_) & (i_13_) & (!i_14_)) + ((sk[54]) & (!i_12_) & (i_13_) & (i_14_)) + ((sk[54]) & (i_12_) & (!i_13_) & (!i_14_)) + ((sk[54]) & (i_12_) & (!i_13_) & (i_14_)) + ((sk[54]) & (i_12_) & (i_13_) & (!i_14_)) + ((sk[54]) & (i_12_) & (i_13_) & (i_14_)));
	assign g25 = (((!sk[55]) & (g20) & (!g24)) + ((!sk[55]) & (g20) & (g24)) + ((sk[55]) & (!g20) & (!g24)) + ((sk[55]) & (!g20) & (g24)) + ((sk[55]) & (g20) & (g24)));
	assign g26 = (((!g18) & (!g21) & (g23) & (!sk[56]) & (!g25)) + ((!g18) & (!g21) & (g23) & (!sk[56]) & (g25)) + ((!g18) & (!g21) & (g23) & (sk[56]) & (g25)) + ((!g18) & (g21) & (!g23) & (!sk[56]) & (g25)) + ((!g18) & (g21) & (g23) & (!sk[56]) & (!g25)) + ((!g18) & (g21) & (g23) & (!sk[56]) & (g25)) + ((g18) & (!g21) & (!g23) & (!sk[56]) & (!g25)) + ((g18) & (!g21) & (!g23) & (!sk[56]) & (g25)) + ((g18) & (!g21) & (g23) & (!sk[56]) & (!g25)) + ((g18) & (!g21) & (g23) & (!sk[56]) & (g25)) + ((g18) & (g21) & (!g23) & (!sk[56]) & (!g25)) + ((g18) & (g21) & (!g23) & (!sk[56]) & (g25)) + ((g18) & (g21) & (g23) & (!sk[56]) & (!g25)) + ((g18) & (g21) & (g23) & (!sk[56]) & (g25)));
	assign g27 = (((!i_9_) & (!sk[57]) & (!i_10_) & (i_11_) & (!i_15_)) + ((!i_9_) & (!sk[57]) & (!i_10_) & (i_11_) & (i_15_)) + ((!i_9_) & (!sk[57]) & (i_10_) & (!i_11_) & (i_15_)) + ((!i_9_) & (!sk[57]) & (i_10_) & (i_11_) & (!i_15_)) + ((!i_9_) & (!sk[57]) & (i_10_) & (i_11_) & (i_15_)) + ((i_9_) & (!sk[57]) & (!i_10_) & (!i_11_) & (!i_15_)) + ((i_9_) & (!sk[57]) & (!i_10_) & (!i_11_) & (i_15_)) + ((i_9_) & (!sk[57]) & (!i_10_) & (i_11_) & (!i_15_)) + ((i_9_) & (!sk[57]) & (!i_10_) & (i_11_) & (i_15_)) + ((i_9_) & (!sk[57]) & (i_10_) & (!i_11_) & (!i_15_)) + ((i_9_) & (!sk[57]) & (i_10_) & (!i_11_) & (i_15_)) + ((i_9_) & (!sk[57]) & (i_10_) & (i_11_) & (!i_15_)) + ((i_9_) & (!sk[57]) & (i_10_) & (i_11_) & (i_15_)) + ((i_9_) & (sk[57]) & (!i_10_) & (!i_11_) & (!i_15_)));
	assign g28 = (((!sk[58]) & (g24) & (!g27)) + ((!sk[58]) & (g24) & (g27)) + ((sk[58]) & (!g24) & (g27)));
	assign g29 = (((!g2) & (!g10) & (!g26) & (sk[59]) & (!g28)) + ((!g2) & (!g10) & (!g26) & (sk[59]) & (g28)) + ((!g2) & (!g10) & (g26) & (!sk[59]) & (!g28)) + ((!g2) & (!g10) & (g26) & (!sk[59]) & (g28)) + ((!g2) & (!g10) & (g26) & (sk[59]) & (!g28)) + ((!g2) & (!g10) & (g26) & (sk[59]) & (g28)) + ((!g2) & (g10) & (!g26) & (!sk[59]) & (g28)) + ((!g2) & (g10) & (g26) & (!sk[59]) & (!g28)) + ((!g2) & (g10) & (g26) & (!sk[59]) & (g28)) + ((g2) & (!g10) & (!g26) & (!sk[59]) & (!g28)) + ((g2) & (!g10) & (!g26) & (!sk[59]) & (g28)) + ((g2) & (!g10) & (g26) & (!sk[59]) & (!g28)) + ((g2) & (!g10) & (g26) & (!sk[59]) & (g28)) + ((g2) & (!g10) & (g26) & (sk[59]) & (!g28)) + ((g2) & (g10) & (!g26) & (!sk[59]) & (!g28)) + ((g2) & (g10) & (!g26) & (!sk[59]) & (g28)) + ((g2) & (g10) & (g26) & (!sk[59]) & (!g28)) + ((g2) & (g10) & (g26) & (!sk[59]) & (g28)));
	assign g30 = (((i_8_) & (!sk[60]) & (!g1)) + ((i_8_) & (!sk[60]) & (g1)) + ((i_8_) & (sk[60]) & (g1)));
	assign g31 = (((g4) & (!g20) & (!sk[61]) & (!g27)) + ((g4) & (!g20) & (!sk[61]) & (g27)) + ((g4) & (!g20) & (sk[61]) & (g27)) + ((g4) & (g20) & (!sk[61]) & (!g27)) + ((g4) & (g20) & (!sk[61]) & (g27)) + ((g4) & (g20) & (sk[61]) & (!g27)) + ((g4) & (g20) & (sk[61]) & (g27)));
	assign g32 = (((!sk[62]) & (!g5) & (!g16) & (!g29) & (!g30) & (g31)) + ((!sk[62]) & (!g5) & (!g16) & (!g29) & (g30) & (g31)) + ((!sk[62]) & (!g5) & (!g16) & (g29) & (!g30) & (g31)) + ((!sk[62]) & (!g5) & (!g16) & (g29) & (g30) & (g31)) + ((!sk[62]) & (!g5) & (g16) & (!g29) & (!g30) & (g31)) + ((!sk[62]) & (!g5) & (g16) & (!g29) & (g30) & (g31)) + ((!sk[62]) & (!g5) & (g16) & (g29) & (!g30) & (g31)) + ((!sk[62]) & (!g5) & (g16) & (g29) & (g30) & (g31)) + ((!sk[62]) & (g5) & (!g16) & (!g29) & (!g30) & (!g31)) + ((!sk[62]) & (g5) & (!g16) & (!g29) & (!g30) & (g31)) + ((!sk[62]) & (g5) & (!g16) & (!g29) & (g30) & (!g31)) + ((!sk[62]) & (g5) & (!g16) & (!g29) & (g30) & (g31)) + ((!sk[62]) & (g5) & (!g16) & (g29) & (!g30) & (!g31)) + ((!sk[62]) & (g5) & (!g16) & (g29) & (!g30) & (g31)) + ((!sk[62]) & (g5) & (!g16) & (g29) & (g30) & (!g31)) + ((!sk[62]) & (g5) & (!g16) & (g29) & (g30) & (g31)) + ((!sk[62]) & (g5) & (g16) & (!g29) & (!g30) & (!g31)) + ((!sk[62]) & (g5) & (g16) & (!g29) & (!g30) & (g31)) + ((!sk[62]) & (g5) & (g16) & (!g29) & (g30) & (!g31)) + ((!sk[62]) & (g5) & (g16) & (!g29) & (g30) & (g31)) + ((!sk[62]) & (g5) & (g16) & (g29) & (!g30) & (!g31)) + ((!sk[62]) & (g5) & (g16) & (g29) & (!g30) & (g31)) + ((!sk[62]) & (g5) & (g16) & (g29) & (g30) & (!g31)) + ((!sk[62]) & (g5) & (g16) & (g29) & (g30) & (g31)) + ((sk[62]) & (!g5) & (g16) & (!g29) & (!g30) & (!g31)) + ((sk[62]) & (!g5) & (g16) & (!g29) & (!g30) & (g31)) + ((sk[62]) & (!g5) & (g16) & (!g29) & (g30) & (!g31)) + ((sk[62]) & (!g5) & (g16) & (!g29) & (g30) & (g31)) + ((sk[62]) & (!g5) & (g16) & (g29) & (g30) & (g31)) + ((sk[62]) & (g5) & (g16) & (!g29) & (!g30) & (!g31)) + ((sk[62]) & (g5) & (g16) & (!g29) & (!g30) & (g31)) + ((sk[62]) & (g5) & (g16) & (!g29) & (g30) & (!g31)) + ((sk[62]) & (g5) & (g16) & (!g29) & (g30) & (g31)) + ((sk[62]) & (g5) & (g16) & (g29) & (g30) & (!g31)) + ((sk[62]) & (g5) & (g16) & (g29) & (g30) & (g31)));
	assign g33 = (((g19) & (!sk[63]) & (!g27)) + ((g19) & (!sk[63]) & (g27)) + ((g19) & (sk[63]) & (g27)));
	assign g34 = (((i_9_) & (!sk[64]) & (!i_10_)) + ((i_9_) & (!sk[64]) & (i_10_)) + ((i_9_) & (sk[64]) & (i_10_)));
	assign g35 = (((!i_11_) & (!i_15_) & (sk[65]) & (g34)) + ((i_11_) & (!i_15_) & (!sk[65]) & (!g34)) + ((i_11_) & (!i_15_) & (!sk[65]) & (g34)) + ((i_11_) & (i_15_) & (!sk[65]) & (!g34)) + ((i_11_) & (i_15_) & (!sk[65]) & (g34)));
	assign g36 = (((!i_9_) & (!i_10_) & (!sk[66]) & (i_11_) & (!i_15_)) + ((!i_9_) & (!i_10_) & (!sk[66]) & (i_11_) & (i_15_)) + ((!i_9_) & (i_10_) & (!sk[66]) & (!i_11_) & (i_15_)) + ((!i_9_) & (i_10_) & (!sk[66]) & (i_11_) & (!i_15_)) + ((!i_9_) & (i_10_) & (!sk[66]) & (i_11_) & (i_15_)) + ((i_9_) & (!i_10_) & (!sk[66]) & (!i_11_) & (!i_15_)) + ((i_9_) & (!i_10_) & (!sk[66]) & (!i_11_) & (i_15_)) + ((i_9_) & (!i_10_) & (!sk[66]) & (i_11_) & (!i_15_)) + ((i_9_) & (!i_10_) & (!sk[66]) & (i_11_) & (i_15_)) + ((i_9_) & (i_10_) & (!sk[66]) & (!i_11_) & (!i_15_)) + ((i_9_) & (i_10_) & (!sk[66]) & (!i_11_) & (i_15_)) + ((i_9_) & (i_10_) & (!sk[66]) & (i_11_) & (!i_15_)) + ((i_9_) & (i_10_) & (!sk[66]) & (i_11_) & (i_15_)) + ((i_9_) & (i_10_) & (sk[66]) & (!i_11_) & (i_15_)));
	assign g37 = (((!g4) & (sk[67]) & (!g36)) + ((!g4) & (sk[67]) & (g36)) + ((g4) & (!sk[67]) & (!g36)) + ((g4) & (!sk[67]) & (g36)) + ((g4) & (sk[67]) & (!g36)));
	assign g38 = (((!g19) & (!g24) & (!g35) & (sk[68]) & (g37)) + ((!g19) & (!g24) & (g35) & (!sk[68]) & (!g37)) + ((!g19) & (!g24) & (g35) & (!sk[68]) & (g37)) + ((!g19) & (g24) & (!g35) & (!sk[68]) & (g37)) + ((!g19) & (g24) & (!g35) & (sk[68]) & (g37)) + ((!g19) & (g24) & (g35) & (!sk[68]) & (!g37)) + ((!g19) & (g24) & (g35) & (!sk[68]) & (g37)) + ((!g19) & (g24) & (g35) & (sk[68]) & (g37)) + ((g19) & (!g24) & (!g35) & (!sk[68]) & (!g37)) + ((g19) & (!g24) & (!g35) & (!sk[68]) & (g37)) + ((g19) & (!g24) & (!g35) & (sk[68]) & (g37)) + ((g19) & (!g24) & (g35) & (!sk[68]) & (!g37)) + ((g19) & (!g24) & (g35) & (!sk[68]) & (g37)) + ((g19) & (g24) & (!g35) & (!sk[68]) & (!g37)) + ((g19) & (g24) & (!g35) & (!sk[68]) & (g37)) + ((g19) & (g24) & (!g35) & (sk[68]) & (g37)) + ((g19) & (g24) & (g35) & (!sk[68]) & (!g37)) + ((g19) & (g24) & (g35) & (!sk[68]) & (g37)));
	assign g39 = (((!sk[69]) & (!g2) & (!g16) & (g33) & (!g38)) + ((!sk[69]) & (!g2) & (!g16) & (g33) & (g38)) + ((!sk[69]) & (!g2) & (g16) & (!g33) & (g38)) + ((!sk[69]) & (!g2) & (g16) & (g33) & (!g38)) + ((!sk[69]) & (!g2) & (g16) & (g33) & (g38)) + ((!sk[69]) & (g2) & (!g16) & (!g33) & (!g38)) + ((!sk[69]) & (g2) & (!g16) & (!g33) & (g38)) + ((!sk[69]) & (g2) & (!g16) & (g33) & (!g38)) + ((!sk[69]) & (g2) & (!g16) & (g33) & (g38)) + ((!sk[69]) & (g2) & (g16) & (!g33) & (!g38)) + ((!sk[69]) & (g2) & (g16) & (!g33) & (g38)) + ((!sk[69]) & (g2) & (g16) & (g33) & (!g38)) + ((!sk[69]) & (g2) & (g16) & (g33) & (g38)) + ((sk[69]) & (g2) & (g16) & (!g33) & (!g38)) + ((sk[69]) & (g2) & (g16) & (g33) & (!g38)) + ((sk[69]) & (g2) & (g16) & (g33) & (g38)));
	assign g40 = (((!sk[70]) & (i_0_) & (!i_1_) & (!i_3_)) + ((!sk[70]) & (i_0_) & (!i_1_) & (i_3_)) + ((!sk[70]) & (i_0_) & (i_1_) & (!i_3_)) + ((!sk[70]) & (i_0_) & (i_1_) & (i_3_)) + ((sk[70]) & (i_0_) & (!i_1_) & (!i_3_)));
	assign g41 = (((!i_4_) & (sk[71]) & (!g39) & (!g40)) + ((i_4_) & (!sk[71]) & (!g39) & (!g40)) + ((i_4_) & (!sk[71]) & (!g39) & (g40)) + ((i_4_) & (!sk[71]) & (g39) & (!g40)) + ((i_4_) & (!sk[71]) & (g39) & (g40)) + ((i_4_) & (sk[71]) & (!g39) & (!g40)) + ((i_4_) & (sk[71]) & (!g39) & (g40)));
	assign g42 = (((!sk[72]) & (i_6_) & (!i_7_)) + ((!sk[72]) & (i_6_) & (i_7_)) + ((sk[72]) & (i_6_) & (!i_7_)));
	assign g43 = (((!sk[73]) & (i_8_) & (!g42)) + ((!sk[73]) & (i_8_) & (g42)) + ((sk[73]) & (!i_8_) & (g42)));
	assign g44 = (((!g16) & (!g43) & (g33) & (!sk[74]) & (!g38)) + ((!g16) & (!g43) & (g33) & (!sk[74]) & (g38)) + ((!g16) & (g43) & (!g33) & (!sk[74]) & (g38)) + ((!g16) & (g43) & (g33) & (!sk[74]) & (!g38)) + ((!g16) & (g43) & (g33) & (!sk[74]) & (g38)) + ((g16) & (!g43) & (!g33) & (!sk[74]) & (!g38)) + ((g16) & (!g43) & (!g33) & (!sk[74]) & (g38)) + ((g16) & (!g43) & (g33) & (!sk[74]) & (!g38)) + ((g16) & (!g43) & (g33) & (!sk[74]) & (g38)) + ((g16) & (g43) & (!g33) & (!sk[74]) & (!g38)) + ((g16) & (g43) & (!g33) & (!sk[74]) & (g38)) + ((g16) & (g43) & (!g33) & (sk[74]) & (!g38)) + ((g16) & (g43) & (g33) & (!sk[74]) & (!g38)) + ((g16) & (g43) & (g33) & (!sk[74]) & (g38)) + ((g16) & (g43) & (g33) & (sk[74]) & (!g38)) + ((g16) & (g43) & (g33) & (sk[74]) & (g38)));
	assign g45 = (((i_6_) & (!sk[75]) & (!i_7_)) + ((i_6_) & (!sk[75]) & (i_7_)) + ((i_6_) & (sk[75]) & (i_7_)));
	assign g46 = (((!g16) & (!sk[76]) & (!g26) & (g43) & (!g45)) + ((!g16) & (!sk[76]) & (!g26) & (g43) & (g45)) + ((!g16) & (!sk[76]) & (g26) & (!g43) & (g45)) + ((!g16) & (!sk[76]) & (g26) & (g43) & (!g45)) + ((!g16) & (!sk[76]) & (g26) & (g43) & (g45)) + ((g16) & (!sk[76]) & (!g26) & (!g43) & (!g45)) + ((g16) & (!sk[76]) & (!g26) & (!g43) & (g45)) + ((g16) & (!sk[76]) & (!g26) & (g43) & (!g45)) + ((g16) & (!sk[76]) & (!g26) & (g43) & (g45)) + ((g16) & (!sk[76]) & (g26) & (!g43) & (!g45)) + ((g16) & (!sk[76]) & (g26) & (!g43) & (g45)) + ((g16) & (!sk[76]) & (g26) & (g43) & (!g45)) + ((g16) & (!sk[76]) & (g26) & (g43) & (g45)) + ((g16) & (sk[76]) & (!g26) & (!g43) & (g45)) + ((g16) & (sk[76]) & (!g26) & (g43) & (!g45)) + ((g16) & (sk[76]) & (!g26) & (g43) & (g45)) + ((g16) & (sk[76]) & (g26) & (!g43) & (g45)) + ((g16) & (sk[76]) & (g26) & (g43) & (g45)));
	assign g47 = (((!i_8_) & (!g4) & (!sk[77]) & (g16) & (!g24)) + ((!i_8_) & (!g4) & (!sk[77]) & (g16) & (g24)) + ((!i_8_) & (!g4) & (sk[77]) & (g16) & (!g24)) + ((!i_8_) & (g4) & (!sk[77]) & (!g16) & (g24)) + ((!i_8_) & (g4) & (!sk[77]) & (g16) & (!g24)) + ((!i_8_) & (g4) & (!sk[77]) & (g16) & (g24)) + ((!i_8_) & (g4) & (sk[77]) & (g16) & (!g24)) + ((i_8_) & (!g4) & (!sk[77]) & (!g16) & (!g24)) + ((i_8_) & (!g4) & (!sk[77]) & (!g16) & (g24)) + ((i_8_) & (!g4) & (!sk[77]) & (g16) & (!g24)) + ((i_8_) & (!g4) & (!sk[77]) & (g16) & (g24)) + ((i_8_) & (g4) & (!sk[77]) & (!g16) & (!g24)) + ((i_8_) & (g4) & (!sk[77]) & (!g16) & (g24)) + ((i_8_) & (g4) & (!sk[77]) & (g16) & (!g24)) + ((i_8_) & (g4) & (!sk[77]) & (g16) & (g24)) + ((i_8_) & (g4) & (sk[77]) & (g16) & (!g24)) + ((i_8_) & (g4) & (sk[77]) & (g16) & (g24)));
	assign g48 = (((!sk[78]) & (g4) & (!g20)) + ((!sk[78]) & (g4) & (g20)) + ((sk[78]) & (g4) & (g20)));
	assign g49 = (((i_8_) & (!sk[79]) & (!g42)) + ((i_8_) & (!sk[79]) & (g42)) + ((i_8_) & (sk[79]) & (g42)));
	assign g50 = (((!g5) & (!sk[80]) & (!g16) & (g48) & (!g49)) + ((!g5) & (!sk[80]) & (!g16) & (g48) & (g49)) + ((!g5) & (!sk[80]) & (g16) & (!g48) & (g49)) + ((!g5) & (!sk[80]) & (g16) & (g48) & (!g49)) + ((!g5) & (!sk[80]) & (g16) & (g48) & (g49)) + ((!g5) & (sk[80]) & (g16) & (g48) & (g49)) + ((g5) & (!sk[80]) & (!g16) & (!g48) & (!g49)) + ((g5) & (!sk[80]) & (!g16) & (!g48) & (g49)) + ((g5) & (!sk[80]) & (!g16) & (g48) & (!g49)) + ((g5) & (!sk[80]) & (!g16) & (g48) & (g49)) + ((g5) & (!sk[80]) & (g16) & (!g48) & (!g49)) + ((g5) & (!sk[80]) & (g16) & (!g48) & (g49)) + ((g5) & (!sk[80]) & (g16) & (g48) & (!g49)) + ((g5) & (!sk[80]) & (g16) & (g48) & (g49)) + ((g5) & (sk[80]) & (g16) & (!g48) & (g49)) + ((g5) & (sk[80]) & (g16) & (g48) & (g49)));
	assign g51 = (((!g27) & (!g42) & (!g44) & (!g46) & (!g47) & (!g50)) + ((!g27) & (!g42) & (!g44) & (!g46) & (g47) & (!g50)) + ((!g27) & (g42) & (!g44) & (!g46) & (!g47) & (!g50)) + ((!g27) & (g42) & (!g44) & (!g46) & (g47) & (!g50)) + ((g27) & (!g42) & (!g44) & (!g46) & (!g47) & (!g50)) + ((g27) & (!g42) & (!g44) & (!g46) & (g47) & (!g50)) + ((g27) & (g42) & (!g44) & (!g46) & (!g47) & (!g50)));
	assign g52 = (((!sk[82]) & (g32) & (!g41) & (!g51)) + ((!sk[82]) & (g32) & (!g41) & (g51)) + ((!sk[82]) & (g32) & (g41) & (!g51)) + ((!sk[82]) & (g32) & (g41) & (g51)) + ((sk[82]) & (!g32) & (g41) & (g51)));
	assign g53 = (((!i_9_) & (sk[83]) & (i_10_)) + ((i_9_) & (!sk[83]) & (!i_10_)) + ((i_9_) & (!sk[83]) & (i_10_)) + ((i_9_) & (sk[83]) & (!i_10_)));
	assign g54 = (((i_4_) & (!i_3_) & (!sk[84]) & (!i_5_)) + ((i_4_) & (!i_3_) & (!sk[84]) & (i_5_)) + ((i_4_) & (!i_3_) & (sk[84]) & (!i_5_)) + ((i_4_) & (i_3_) & (!sk[84]) & (!i_5_)) + ((i_4_) & (i_3_) & (!sk[84]) & (i_5_)));
	assign g55 = (((g14) & (!sk[85]) & (!g54)) + ((g14) & (!sk[85]) & (g54)) + ((g14) & (sk[85]) & (g54)));
	assign g56 = (((!i_12_) & (!i_13_) & (sk[86]) & (i_14_)) + ((!i_12_) & (i_13_) & (sk[86]) & (!i_14_)) + ((i_12_) & (!i_13_) & (!sk[86]) & (!i_14_)) + ((i_12_) & (!i_13_) & (!sk[86]) & (i_14_)) + ((i_12_) & (i_13_) & (!sk[86]) & (!i_14_)) + ((i_12_) & (i_13_) & (!sk[86]) & (i_14_)));
	assign g57 = (((!g2) & (!g35) & (!sk[87]) & (!g37) & (!g55) & (g56)) + ((!g2) & (!g35) & (!sk[87]) & (!g37) & (g55) & (g56)) + ((!g2) & (!g35) & (!sk[87]) & (g37) & (!g55) & (g56)) + ((!g2) & (!g35) & (!sk[87]) & (g37) & (g55) & (g56)) + ((!g2) & (g35) & (!sk[87]) & (!g37) & (!g55) & (g56)) + ((!g2) & (g35) & (!sk[87]) & (!g37) & (g55) & (g56)) + ((!g2) & (g35) & (!sk[87]) & (g37) & (!g55) & (g56)) + ((!g2) & (g35) & (!sk[87]) & (g37) & (g55) & (g56)) + ((g2) & (!g35) & (!sk[87]) & (!g37) & (!g55) & (!g56)) + ((g2) & (!g35) & (!sk[87]) & (!g37) & (!g55) & (g56)) + ((g2) & (!g35) & (!sk[87]) & (!g37) & (g55) & (!g56)) + ((g2) & (!g35) & (!sk[87]) & (!g37) & (g55) & (g56)) + ((g2) & (!g35) & (!sk[87]) & (g37) & (!g55) & (!g56)) + ((g2) & (!g35) & (!sk[87]) & (g37) & (!g55) & (g56)) + ((g2) & (!g35) & (!sk[87]) & (g37) & (g55) & (!g56)) + ((g2) & (!g35) & (!sk[87]) & (g37) & (g55) & (g56)) + ((g2) & (!g35) & (sk[87]) & (!g37) & (g55) & (!g56)) + ((g2) & (!g35) & (sk[87]) & (!g37) & (g55) & (g56)) + ((g2) & (g35) & (!sk[87]) & (!g37) & (!g55) & (!g56)) + ((g2) & (g35) & (!sk[87]) & (!g37) & (!g55) & (g56)) + ((g2) & (g35) & (!sk[87]) & (!g37) & (g55) & (!g56)) + ((g2) & (g35) & (!sk[87]) & (!g37) & (g55) & (g56)) + ((g2) & (g35) & (!sk[87]) & (g37) & (!g55) & (!g56)) + ((g2) & (g35) & (!sk[87]) & (g37) & (!g55) & (g56)) + ((g2) & (g35) & (!sk[87]) & (g37) & (g55) & (!g56)) + ((g2) & (g35) & (!sk[87]) & (g37) & (g55) & (g56)) + ((g2) & (g35) & (sk[87]) & (!g37) & (g55) & (!g56)) + ((g2) & (g35) & (sk[87]) & (!g37) & (g55) & (g56)) + ((g2) & (g35) & (sk[87]) & (g37) & (g55) & (g56)));
	assign g58 = (((!i_0_) & (!i_1_) & (!sk[88]) & (!i_2_) & (!g10) & (g54)) + ((!i_0_) & (!i_1_) & (!sk[88]) & (!i_2_) & (g10) & (g54)) + ((!i_0_) & (!i_1_) & (!sk[88]) & (i_2_) & (!g10) & (g54)) + ((!i_0_) & (!i_1_) & (!sk[88]) & (i_2_) & (g10) & (g54)) + ((!i_0_) & (i_1_) & (!sk[88]) & (!i_2_) & (!g10) & (g54)) + ((!i_0_) & (i_1_) & (!sk[88]) & (!i_2_) & (g10) & (g54)) + ((!i_0_) & (i_1_) & (!sk[88]) & (i_2_) & (!g10) & (g54)) + ((!i_0_) & (i_1_) & (!sk[88]) & (i_2_) & (g10) & (g54)) + ((!i_0_) & (i_1_) & (sk[88]) & (!i_2_) & (g10) & (g54)) + ((i_0_) & (!i_1_) & (!sk[88]) & (!i_2_) & (!g10) & (!g54)) + ((i_0_) & (!i_1_) & (!sk[88]) & (!i_2_) & (!g10) & (g54)) + ((i_0_) & (!i_1_) & (!sk[88]) & (!i_2_) & (g10) & (!g54)) + ((i_0_) & (!i_1_) & (!sk[88]) & (!i_2_) & (g10) & (g54)) + ((i_0_) & (!i_1_) & (!sk[88]) & (i_2_) & (!g10) & (!g54)) + ((i_0_) & (!i_1_) & (!sk[88]) & (i_2_) & (!g10) & (g54)) + ((i_0_) & (!i_1_) & (!sk[88]) & (i_2_) & (g10) & (!g54)) + ((i_0_) & (!i_1_) & (!sk[88]) & (i_2_) & (g10) & (g54)) + ((i_0_) & (!i_1_) & (sk[88]) & (!i_2_) & (!g10) & (g54)) + ((i_0_) & (!i_1_) & (sk[88]) & (!i_2_) & (g10) & (g54)) + ((i_0_) & (!i_1_) & (sk[88]) & (i_2_) & (!g10) & (g54)) + ((i_0_) & (!i_1_) & (sk[88]) & (i_2_) & (g10) & (g54)) + ((i_0_) & (i_1_) & (!sk[88]) & (!i_2_) & (!g10) & (!g54)) + ((i_0_) & (i_1_) & (!sk[88]) & (!i_2_) & (!g10) & (g54)) + ((i_0_) & (i_1_) & (!sk[88]) & (!i_2_) & (g10) & (!g54)) + ((i_0_) & (i_1_) & (!sk[88]) & (!i_2_) & (g10) & (g54)) + ((i_0_) & (i_1_) & (!sk[88]) & (i_2_) & (!g10) & (!g54)) + ((i_0_) & (i_1_) & (!sk[88]) & (i_2_) & (!g10) & (g54)) + ((i_0_) & (i_1_) & (!sk[88]) & (i_2_) & (g10) & (!g54)) + ((i_0_) & (i_1_) & (!sk[88]) & (i_2_) & (g10) & (g54)));
	assign g59 = (((!g2) & (!g26) & (!g28) & (!g33) & (!g55) & (!g58)) + ((!g2) & (!g26) & (!g28) & (!g33) & (g55) & (!g58)) + ((!g2) & (!g26) & (!g28) & (g33) & (!g55) & (!g58)) + ((!g2) & (!g26) & (!g28) & (g33) & (g55) & (!g58)) + ((!g2) & (!g26) & (g28) & (!g33) & (!g55) & (!g58)) + ((!g2) & (!g26) & (g28) & (!g33) & (g55) & (!g58)) + ((!g2) & (!g26) & (g28) & (g33) & (!g55) & (!g58)) + ((!g2) & (!g26) & (g28) & (g33) & (g55) & (!g58)) + ((!g2) & (g26) & (!g28) & (!g33) & (!g55) & (!g58)) + ((!g2) & (g26) & (!g28) & (!g33) & (g55) & (!g58)) + ((!g2) & (g26) & (!g28) & (g33) & (!g55) & (!g58)) + ((!g2) & (g26) & (!g28) & (g33) & (g55) & (!g58)) + ((!g2) & (g26) & (g28) & (!g33) & (!g55) & (!g58)) + ((!g2) & (g26) & (g28) & (!g33) & (g55) & (!g58)) + ((!g2) & (g26) & (g28) & (g33) & (!g55) & (!g58)) + ((!g2) & (g26) & (g28) & (g33) & (g55) & (!g58)) + ((g2) & (!g26) & (!g28) & (!g33) & (!g55) & (!g58)) + ((g2) & (!g26) & (!g28) & (g33) & (!g55) & (!g58)) + ((g2) & (!g26) & (g28) & (!g33) & (!g55) & (!g58)) + ((g2) & (!g26) & (g28) & (g33) & (!g55) & (!g58)) + ((g2) & (g26) & (!g28) & (!g33) & (!g55) & (!g58)) + ((g2) & (g26) & (!g28) & (!g33) & (g55) & (!g58)) + ((g2) & (g26) & (!g28) & (g33) & (!g55) & (!g58)) + ((g2) & (g26) & (g28) & (!g33) & (!g55) & (!g58)) + ((g2) & (g26) & (g28) & (g33) & (!g55) & (!g58)));
	assign g60 = (((!sk[90]) & (i_11_) & (!i_15_) & (!g4)) + ((!sk[90]) & (i_11_) & (!i_15_) & (g4)) + ((!sk[90]) & (i_11_) & (i_15_) & (!g4)) + ((!sk[90]) & (i_11_) & (i_15_) & (g4)) + ((sk[90]) & (!i_11_) & (!i_15_) & (g4)));
	assign g61 = (((!g30) & (!g53) & (!g55) & (!g57) & (g59) & (!g60)) + ((!g30) & (!g53) & (!g55) & (!g57) & (g59) & (g60)) + ((!g30) & (!g53) & (g55) & (!g57) & (g59) & (!g60)) + ((!g30) & (!g53) & (g55) & (!g57) & (g59) & (g60)) + ((!g30) & (g53) & (!g55) & (!g57) & (g59) & (!g60)) + ((!g30) & (g53) & (!g55) & (!g57) & (g59) & (g60)) + ((!g30) & (g53) & (g55) & (!g57) & (g59) & (!g60)) + ((!g30) & (g53) & (g55) & (!g57) & (g59) & (g60)) + ((g30) & (!g53) & (!g55) & (!g57) & (g59) & (!g60)) + ((g30) & (!g53) & (!g55) & (!g57) & (g59) & (g60)) + ((g30) & (!g53) & (g55) & (!g57) & (g59) & (!g60)) + ((g30) & (!g53) & (g55) & (!g57) & (g59) & (g60)) + ((g30) & (g53) & (!g55) & (!g57) & (g59) & (!g60)) + ((g30) & (g53) & (!g55) & (!g57) & (g59) & (g60)) + ((g30) & (g53) & (g55) & (!g57) & (g59) & (!g60)));
	assign g62 = (((!sk[92]) & (!i_4_) & (!i_3_) & (i_5_)) + ((!sk[92]) & (!i_4_) & (i_3_) & (i_5_)) + ((!sk[92]) & (i_4_) & (!i_3_) & (i_5_)) + ((!sk[92]) & (i_4_) & (i_3_) & (!i_5_)) + ((!sk[92]) & (i_4_) & (i_3_) & (i_5_)) + ((sk[92]) & (i_4_) & (!i_3_) & (i_5_)));
	assign g63 = (((!i_0_) & (!i_1_) & (!sk[93]) & (g62)) + ((!i_0_) & (i_1_) & (!sk[93]) & (g62)) + ((i_0_) & (!i_1_) & (!sk[93]) & (g62)) + ((i_0_) & (!i_1_) & (sk[93]) & (g62)) + ((i_0_) & (i_1_) & (!sk[93]) & (!g62)) + ((i_0_) & (i_1_) & (!sk[93]) & (g62)));
	assign g64 = (((!g26) & (!g28) & (!g43) & (!sk[94]) & (g33) & (g55)) + ((!g26) & (!g28) & (g43) & (!sk[94]) & (g33) & (g55)) + ((!g26) & (!g28) & (g43) & (sk[94]) & (!g33) & (g55)) + ((!g26) & (!g28) & (g43) & (sk[94]) & (g33) & (g55)) + ((!g26) & (g28) & (!g43) & (!sk[94]) & (!g33) & (!g55)) + ((!g26) & (g28) & (!g43) & (!sk[94]) & (!g33) & (g55)) + ((!g26) & (g28) & (!g43) & (!sk[94]) & (g33) & (!g55)) + ((!g26) & (g28) & (!g43) & (!sk[94]) & (g33) & (g55)) + ((!g26) & (g28) & (g43) & (!sk[94]) & (!g33) & (!g55)) + ((!g26) & (g28) & (g43) & (!sk[94]) & (!g33) & (g55)) + ((!g26) & (g28) & (g43) & (!sk[94]) & (g33) & (!g55)) + ((!g26) & (g28) & (g43) & (!sk[94]) & (g33) & (g55)) + ((!g26) & (g28) & (g43) & (sk[94]) & (!g33) & (g55)) + ((!g26) & (g28) & (g43) & (sk[94]) & (g33) & (g55)) + ((g26) & (!g28) & (!g43) & (!sk[94]) & (g33) & (g55)) + ((g26) & (!g28) & (g43) & (!sk[94]) & (g33) & (g55)) + ((g26) & (!g28) & (g43) & (sk[94]) & (g33) & (g55)) + ((g26) & (g28) & (!g43) & (!sk[94]) & (!g33) & (!g55)) + ((g26) & (g28) & (!g43) & (!sk[94]) & (!g33) & (g55)) + ((g26) & (g28) & (!g43) & (!sk[94]) & (g33) & (!g55)) + ((g26) & (g28) & (!g43) & (!sk[94]) & (g33) & (g55)) + ((g26) & (g28) & (g43) & (!sk[94]) & (!g33) & (!g55)) + ((g26) & (g28) & (g43) & (!sk[94]) & (!g33) & (g55)) + ((g26) & (g28) & (g43) & (!sk[94]) & (g33) & (!g55)) + ((g26) & (g28) & (g43) & (!sk[94]) & (g33) & (g55)) + ((g26) & (g28) & (g43) & (sk[94]) & (!g33) & (g55)) + ((g26) & (g28) & (g43) & (sk[94]) & (g33) & (g55)));
	assign g65 = (((!sk[95]) & (!i_6_) & (!i_7_) & (!g55) & (g63) & (g64)) + ((!sk[95]) & (!i_6_) & (!i_7_) & (g55) & (g63) & (g64)) + ((!sk[95]) & (!i_6_) & (i_7_) & (!g55) & (!g63) & (!g64)) + ((!sk[95]) & (!i_6_) & (i_7_) & (!g55) & (!g63) & (g64)) + ((!sk[95]) & (!i_6_) & (i_7_) & (!g55) & (g63) & (!g64)) + ((!sk[95]) & (!i_6_) & (i_7_) & (!g55) & (g63) & (g64)) + ((!sk[95]) & (!i_6_) & (i_7_) & (g55) & (!g63) & (!g64)) + ((!sk[95]) & (!i_6_) & (i_7_) & (g55) & (!g63) & (g64)) + ((!sk[95]) & (!i_6_) & (i_7_) & (g55) & (g63) & (!g64)) + ((!sk[95]) & (!i_6_) & (i_7_) & (g55) & (g63) & (g64)) + ((!sk[95]) & (i_6_) & (!i_7_) & (!g55) & (g63) & (g64)) + ((!sk[95]) & (i_6_) & (!i_7_) & (g55) & (g63) & (g64)) + ((!sk[95]) & (i_6_) & (i_7_) & (!g55) & (!g63) & (!g64)) + ((!sk[95]) & (i_6_) & (i_7_) & (!g55) & (!g63) & (g64)) + ((!sk[95]) & (i_6_) & (i_7_) & (!g55) & (g63) & (!g64)) + ((!sk[95]) & (i_6_) & (i_7_) & (!g55) & (g63) & (g64)) + ((!sk[95]) & (i_6_) & (i_7_) & (g55) & (!g63) & (!g64)) + ((!sk[95]) & (i_6_) & (i_7_) & (g55) & (!g63) & (g64)) + ((!sk[95]) & (i_6_) & (i_7_) & (g55) & (g63) & (!g64)) + ((!sk[95]) & (i_6_) & (i_7_) & (g55) & (g63) & (g64)) + ((sk[95]) & (!i_6_) & (!i_7_) & (!g55) & (!g63) & (!g64)) + ((sk[95]) & (!i_6_) & (!i_7_) & (g55) & (!g63) & (!g64)) + ((sk[95]) & (!i_6_) & (i_7_) & (!g55) & (!g63) & (!g64)) + ((sk[95]) & (!i_6_) & (i_7_) & (g55) & (!g63) & (!g64)) + ((sk[95]) & (i_6_) & (!i_7_) & (!g55) & (!g63) & (!g64)) + ((sk[95]) & (i_6_) & (!i_7_) & (g55) & (!g63) & (!g64)) + ((sk[95]) & (i_6_) & (i_7_) & (!g55) & (!g63) & (!g64)));
	assign g66 = (((!i_8_) & (!g31) & (!g42) & (!g38) & (!g55) & (g65)) + ((!i_8_) & (!g31) & (!g42) & (!g38) & (g55) & (g65)) + ((!i_8_) & (!g31) & (!g42) & (g38) & (!g55) & (g65)) + ((!i_8_) & (!g31) & (!g42) & (g38) & (g55) & (g65)) + ((!i_8_) & (!g31) & (g42) & (!g38) & (!g55) & (g65)) + ((!i_8_) & (!g31) & (g42) & (g38) & (!g55) & (g65)) + ((!i_8_) & (!g31) & (g42) & (g38) & (g55) & (g65)) + ((!i_8_) & (g31) & (!g42) & (!g38) & (!g55) & (g65)) + ((!i_8_) & (g31) & (!g42) & (!g38) & (g55) & (g65)) + ((!i_8_) & (g31) & (!g42) & (g38) & (!g55) & (g65)) + ((!i_8_) & (g31) & (!g42) & (g38) & (g55) & (g65)) + ((!i_8_) & (g31) & (g42) & (!g38) & (!g55) & (g65)) + ((!i_8_) & (g31) & (g42) & (g38) & (!g55) & (g65)) + ((!i_8_) & (g31) & (g42) & (g38) & (g55) & (g65)) + ((i_8_) & (!g31) & (!g42) & (!g38) & (!g55) & (g65)) + ((i_8_) & (!g31) & (!g42) & (!g38) & (g55) & (g65)) + ((i_8_) & (!g31) & (!g42) & (g38) & (!g55) & (g65)) + ((i_8_) & (!g31) & (!g42) & (g38) & (g55) & (g65)) + ((i_8_) & (!g31) & (g42) & (!g38) & (!g55) & (g65)) + ((i_8_) & (!g31) & (g42) & (!g38) & (g55) & (g65)) + ((i_8_) & (!g31) & (g42) & (g38) & (!g55) & (g65)) + ((i_8_) & (!g31) & (g42) & (g38) & (g55) & (g65)) + ((i_8_) & (g31) & (!g42) & (!g38) & (!g55) & (g65)) + ((i_8_) & (g31) & (!g42) & (!g38) & (g55) & (g65)) + ((i_8_) & (g31) & (!g42) & (g38) & (!g55) & (g65)) + ((i_8_) & (g31) & (!g42) & (g38) & (g55) & (g65)) + ((i_8_) & (g31) & (g42) & (!g38) & (!g55) & (g65)) + ((i_8_) & (g31) & (g42) & (g38) & (!g55) & (g65)));
	assign o_4_ = (((!g61) & (!sk[97]) & (g66)) + ((!g61) & (sk[97]) & (!g66)) + ((!g61) & (sk[97]) & (g66)) + ((g61) & (!sk[97]) & (g66)) + ((g61) & (sk[97]) & (!g66)));
	assign g68 = (((!i_12_) & (!sk[98]) & (!i_13_) & (i_14_)) + ((!i_12_) & (!sk[98]) & (i_13_) & (i_14_)) + ((!i_12_) & (sk[98]) & (!i_13_) & (!i_14_)) + ((!i_12_) & (sk[98]) & (!i_13_) & (i_14_)) + ((!i_12_) & (sk[98]) & (i_13_) & (!i_14_)) + ((!i_12_) & (sk[98]) & (i_13_) & (i_14_)) + ((i_12_) & (!sk[98]) & (!i_13_) & (i_14_)) + ((i_12_) & (!sk[98]) & (i_13_) & (!i_14_)) + ((i_12_) & (!sk[98]) & (i_13_) & (i_14_)) + ((i_12_) & (sk[98]) & (!i_13_) & (i_14_)) + ((i_12_) & (sk[98]) & (i_13_) & (!i_14_)) + ((i_12_) & (sk[98]) & (i_13_) & (i_14_)));
	assign g69 = (((!i_9_) & (!i_10_) & (!i_11_) & (!sk[99]) & (i_15_)) + ((!i_9_) & (!i_10_) & (!i_11_) & (sk[99]) & (i_15_)) + ((!i_9_) & (!i_10_) & (i_11_) & (!sk[99]) & (i_15_)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[99]) & (i_15_)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[99]) & (i_15_)) + ((i_9_) & (!i_10_) & (!i_11_) & (!sk[99]) & (!i_15_)) + ((i_9_) & (!i_10_) & (!i_11_) & (!sk[99]) & (i_15_)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[99]) & (!i_15_)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[99]) & (i_15_)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[99]) & (!i_15_)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[99]) & (i_15_)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[99]) & (!i_15_)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[99]) & (i_15_)));
	assign g70 = (((!sk[100]) & (g68) & (g69)) + ((sk[100]) & (!g68) & (g69)));
	assign g71 = (((!sk[101]) & (i_0_) & (i_1_) & (!i_2_)) + ((!sk[101]) & (i_0_) & (i_1_) & (i_2_)) + ((sk[101]) & (!i_0_) & (!i_1_) & (!i_2_)));
	assign g72 = (((!sk[102]) & (g62) & (g71)) + ((sk[102]) & (g62) & (g71)));
	assign g73 = (((g10) & (!sk[103]) & (g72)) + ((g10) & (sk[103]) & (g72)));
	assign g74 = (((!i_8_) & (sk[104]) & (g73)) + ((i_8_) & (!sk[104]) & (g73)));
	assign g75 = (((!sk[105]) & (i_8_) & (g73)) + ((sk[105]) & (!i_8_) & (!g73)) + ((sk[105]) & (!i_8_) & (g73)) + ((sk[105]) & (i_8_) & (!g73)));
	assign g76 = (((!i_12_) & (sk[106]) & (!i_13_) & (!i_14_)) + ((!i_12_) & (sk[106]) & (!i_13_) & (i_14_)) + ((!i_12_) & (sk[106]) & (i_13_) & (!i_14_)) + ((i_12_) & (!sk[106]) & (i_13_) & (!i_14_)) + ((i_12_) & (!sk[106]) & (i_13_) & (i_14_)) + ((i_12_) & (sk[106]) & (!i_13_) & (!i_14_)) + ((i_12_) & (sk[106]) & (!i_13_) & (i_14_)) + ((i_12_) & (sk[106]) & (i_13_) & (!i_14_)) + ((i_12_) & (sk[106]) & (i_13_) & (i_14_)));
	assign g77 = (((!sk[107]) & (g3) & (g76)) + ((sk[107]) & (g3) & (!g76)));
	assign g78 = (((!sk[108]) & (g22) & (g68)) + ((sk[108]) & (!g22) & (g68)) + ((sk[108]) & (g22) & (!g68)) + ((sk[108]) & (g22) & (g68)));
	assign g79 = (((!g20) & (sk[109]) & (!g76)) + ((!g20) & (sk[109]) & (g76)) + ((g20) & (!sk[109]) & (g76)) + ((g20) & (sk[109]) & (g76)));
	assign g80 = (((!i_9_) & (sk[110]) & (!i_10_)) + ((i_9_) & (!sk[110]) & (i_10_)));
	assign g81 = (((!sk[111]) & (g80) & (i_11_) & (!i_15_)) + ((!sk[111]) & (g80) & (i_11_) & (i_15_)) + ((sk[111]) & (g80) & (i_11_) & (i_15_)));
	assign g82 = (((!sk[112]) & (g68) & (g81)) + ((sk[112]) & (!g68) & (g81)));
	assign g83 = (((g80) & (!sk[113]) & (i_11_) & (!i_15_)) + ((g80) & (!sk[113]) & (i_11_) & (i_15_)) + ((g80) & (sk[113]) & (i_11_) & (!i_15_)));
	assign g84 = (((!i_8_) & (!g73) & (!g76) & (g82) & (!sk[114]) & (!g83)) + ((!i_8_) & (!g73) & (!g76) & (g82) & (!sk[114]) & (g83)) + ((!i_8_) & (!g73) & (g76) & (!g82) & (!sk[114]) & (!g83)) + ((!i_8_) & (!g73) & (g76) & (!g82) & (!sk[114]) & (g83)) + ((!i_8_) & (!g73) & (g76) & (g82) & (!sk[114]) & (!g83)) + ((!i_8_) & (!g73) & (g76) & (g82) & (!sk[114]) & (g83)) + ((!i_8_) & (g73) & (!g76) & (g82) & (!sk[114]) & (!g83)) + ((!i_8_) & (g73) & (!g76) & (g82) & (!sk[114]) & (g83)) + ((!i_8_) & (g73) & (g76) & (!g82) & (!sk[114]) & (!g83)) + ((!i_8_) & (g73) & (g76) & (!g82) & (!sk[114]) & (g83)) + ((!i_8_) & (g73) & (g76) & (g82) & (!sk[114]) & (!g83)) + ((!i_8_) & (g73) & (g76) & (g82) & (!sk[114]) & (g83)) + ((i_8_) & (!g73) & (!g76) & (g82) & (!sk[114]) & (!g83)) + ((i_8_) & (!g73) & (!g76) & (g82) & (!sk[114]) & (g83)) + ((i_8_) & (!g73) & (g76) & (!g82) & (!sk[114]) & (!g83)) + ((i_8_) & (!g73) & (g76) & (!g82) & (!sk[114]) & (g83)) + ((i_8_) & (!g73) & (g76) & (g82) & (!sk[114]) & (!g83)) + ((i_8_) & (!g73) & (g76) & (g82) & (!sk[114]) & (g83)) + ((i_8_) & (g73) & (!g76) & (!g82) & (sk[114]) & (g83)) + ((i_8_) & (g73) & (!g76) & (g82) & (!sk[114]) & (!g83)) + ((i_8_) & (g73) & (!g76) & (g82) & (!sk[114]) & (g83)) + ((i_8_) & (g73) & (!g76) & (g82) & (sk[114]) & (!g83)) + ((i_8_) & (g73) & (!g76) & (g82) & (sk[114]) & (g83)) + ((i_8_) & (g73) & (g76) & (!g82) & (!sk[114]) & (!g83)) + ((i_8_) & (g73) & (g76) & (!g82) & (!sk[114]) & (g83)) + ((i_8_) & (g73) & (g76) & (g82) & (!sk[114]) & (!g83)) + ((i_8_) & (g73) & (g76) & (g82) & (!sk[114]) & (g83)) + ((i_8_) & (g73) & (g76) & (g82) & (sk[114]) & (!g83)) + ((i_8_) & (g73) & (g76) & (g82) & (sk[114]) & (g83)));
	assign g85 = (((!g75) & (!g77) & (!g70) & (g78) & (g79) & (!g84)) + ((g75) & (!g77) & (!g70) & (!g78) & (!g79) & (!g84)) + ((g75) & (!g77) & (!g70) & (!g78) & (g79) & (!g84)) + ((g75) & (!g77) & (!g70) & (g78) & (!g79) & (!g84)) + ((g75) & (!g77) & (!g70) & (g78) & (g79) & (!g84)) + ((g75) & (!g77) & (g70) & (!g78) & (!g79) & (!g84)) + ((g75) & (!g77) & (g70) & (!g78) & (g79) & (!g84)) + ((g75) & (!g77) & (g70) & (g78) & (!g79) & (!g84)) + ((g75) & (!g77) & (g70) & (g78) & (g79) & (!g84)) + ((g75) & (g77) & (!g70) & (!g78) & (!g79) & (!g84)) + ((g75) & (g77) & (!g70) & (!g78) & (g79) & (!g84)) + ((g75) & (g77) & (!g70) & (g78) & (!g79) & (!g84)) + ((g75) & (g77) & (!g70) & (g78) & (g79) & (!g84)) + ((g75) & (g77) & (g70) & (!g78) & (!g79) & (!g84)) + ((g75) & (g77) & (g70) & (!g78) & (g79) & (!g84)) + ((g75) & (g77) & (g70) & (g78) & (!g79) & (!g84)) + ((g75) & (g77) & (g70) & (g78) & (g79) & (!g84)));
	assign g86 = (((!i_9_) & (!sk[116]) & (!i_10_) & (!i_11_) & (i_15_)) + ((!i_9_) & (!sk[116]) & (!i_10_) & (i_11_) & (i_15_)) + ((!i_9_) & (!sk[116]) & (i_10_) & (!i_11_) & (i_15_)) + ((!i_9_) & (!sk[116]) & (i_10_) & (i_11_) & (i_15_)) + ((i_9_) & (!sk[116]) & (!i_10_) & (!i_11_) & (i_15_)) + ((i_9_) & (!sk[116]) & (!i_10_) & (i_11_) & (i_15_)) + ((i_9_) & (!sk[116]) & (i_10_) & (!i_11_) & (!i_15_)) + ((i_9_) & (!sk[116]) & (i_10_) & (!i_11_) & (i_15_)) + ((i_9_) & (!sk[116]) & (i_10_) & (i_11_) & (!i_15_)) + ((i_9_) & (!sk[116]) & (i_10_) & (i_11_) & (i_15_)) + ((i_9_) & (sk[116]) & (!i_10_) & (i_11_) & (!i_15_)));
	assign g87 = (((!sk[117]) & (g76) & (g86)) + ((sk[117]) & (!g76) & (!g86)) + ((sk[117]) & (g76) & (!g86)) + ((sk[117]) & (g76) & (g86)));
	assign g88 = (((!i_9_) & (!sk[118]) & (!i_10_) & (!i_11_) & (i_15_)) + ((!i_9_) & (!sk[118]) & (!i_10_) & (i_11_) & (i_15_)) + ((!i_9_) & (!sk[118]) & (i_10_) & (!i_11_) & (i_15_)) + ((!i_9_) & (!sk[118]) & (i_10_) & (i_11_) & (i_15_)) + ((i_9_) & (!sk[118]) & (!i_10_) & (!i_11_) & (i_15_)) + ((i_9_) & (!sk[118]) & (!i_10_) & (i_11_) & (i_15_)) + ((i_9_) & (!sk[118]) & (i_10_) & (!i_11_) & (!i_15_)) + ((i_9_) & (!sk[118]) & (i_10_) & (!i_11_) & (i_15_)) + ((i_9_) & (!sk[118]) & (i_10_) & (i_11_) & (!i_15_)) + ((i_9_) & (!sk[118]) & (i_10_) & (i_11_) & (i_15_)) + ((i_9_) & (sk[118]) & (!i_10_) & (i_11_) & (i_15_)));
	assign g89 = (((!sk[119]) & (g68) & (g88)) + ((sk[119]) & (!g68) & (!g88)) + ((sk[119]) & (g68) & (!g88)) + ((sk[119]) & (g68) & (g88)));
	assign g90 = (((!sk[120]) & (g36) & (g68)) + ((sk[120]) & (g36) & (!g68)));
	assign g91 = (((!i_9_) & (!sk[121]) & (!i_10_) & (!i_11_) & (i_15_)) + ((!i_9_) & (!sk[121]) & (!i_10_) & (i_11_) & (i_15_)) + ((!i_9_) & (!sk[121]) & (i_10_) & (!i_11_) & (i_15_)) + ((!i_9_) & (!sk[121]) & (i_10_) & (i_11_) & (i_15_)) + ((!i_9_) & (sk[121]) & (!i_10_) & (!i_11_) & (!i_15_)) + ((!i_9_) & (sk[121]) & (!i_10_) & (!i_11_) & (i_15_)) + ((!i_9_) & (sk[121]) & (!i_10_) & (i_11_) & (!i_15_)) + ((!i_9_) & (sk[121]) & (!i_10_) & (i_11_) & (i_15_)) + ((!i_9_) & (sk[121]) & (i_10_) & (!i_11_) & (!i_15_)) + ((!i_9_) & (sk[121]) & (i_10_) & (!i_11_) & (i_15_)) + ((!i_9_) & (sk[121]) & (i_10_) & (i_11_) & (!i_15_)) + ((!i_9_) & (sk[121]) & (i_10_) & (i_11_) & (i_15_)) + ((i_9_) & (!sk[121]) & (!i_10_) & (!i_11_) & (i_15_)) + ((i_9_) & (!sk[121]) & (!i_10_) & (i_11_) & (i_15_)) + ((i_9_) & (!sk[121]) & (i_10_) & (!i_11_) & (!i_15_)) + ((i_9_) & (!sk[121]) & (i_10_) & (!i_11_) & (i_15_)) + ((i_9_) & (!sk[121]) & (i_10_) & (i_11_) & (!i_15_)) + ((i_9_) & (!sk[121]) & (i_10_) & (i_11_) & (i_15_)) + ((i_9_) & (sk[121]) & (!i_10_) & (!i_11_) & (!i_15_)) + ((i_9_) & (sk[121]) & (!i_10_) & (!i_11_) & (i_15_)) + ((i_9_) & (sk[121]) & (!i_10_) & (i_11_) & (!i_15_)) + ((i_9_) & (sk[121]) & (!i_10_) & (i_11_) & (i_15_)) + ((i_9_) & (sk[121]) & (i_10_) & (!i_11_) & (!i_15_)) + ((i_9_) & (sk[121]) & (i_10_) & (!i_11_) & (i_15_)) + ((i_9_) & (sk[121]) & (i_10_) & (i_11_) & (!i_15_)));
	assign g92 = (((!sk[122]) & (g68) & (g91)) + ((sk[122]) & (!g68) & (!g91)));
	assign g93 = (((!i_15_) & (sk[123]) & (!g76)) + ((i_15_) & (!sk[123]) & (g76)));
	assign g94 = (((g80) & (!sk[124]) & (g93)) + ((g80) & (sk[124]) & (g93)));
	assign g95 = (((!i_8_) & (g73) & (!g90) & (!g82) & (!g92) & (g94)) + ((!i_8_) & (g73) & (!g90) & (!g82) & (g92) & (!g94)) + ((!i_8_) & (g73) & (!g90) & (!g82) & (g92) & (g94)) + ((!i_8_) & (g73) & (!g90) & (g82) & (!g92) & (!g94)) + ((!i_8_) & (g73) & (!g90) & (g82) & (!g92) & (g94)) + ((!i_8_) & (g73) & (!g90) & (g82) & (g92) & (!g94)) + ((!i_8_) & (g73) & (!g90) & (g82) & (g92) & (g94)) + ((!i_8_) & (g73) & (g90) & (!g82) & (!g92) & (!g94)) + ((!i_8_) & (g73) & (g90) & (!g82) & (!g92) & (g94)) + ((!i_8_) & (g73) & (g90) & (!g82) & (g92) & (!g94)) + ((!i_8_) & (g73) & (g90) & (!g82) & (g92) & (g94)) + ((!i_8_) & (g73) & (g90) & (g82) & (!g92) & (!g94)) + ((!i_8_) & (g73) & (g90) & (g82) & (!g92) & (g94)) + ((!i_8_) & (g73) & (g90) & (g82) & (g92) & (!g94)) + ((!i_8_) & (g73) & (g90) & (g82) & (g92) & (g94)) + ((i_8_) & (g73) & (g90) & (!g82) & (!g92) & (!g94)) + ((i_8_) & (g73) & (g90) & (!g82) & (!g92) & (g94)) + ((i_8_) & (g73) & (g90) & (!g82) & (g92) & (!g94)) + ((i_8_) & (g73) & (g90) & (!g82) & (g92) & (g94)) + ((i_8_) & (g73) & (g90) & (g82) & (!g92) & (!g94)) + ((i_8_) & (g73) & (g90) & (g82) & (!g92) & (g94)) + ((i_8_) & (g73) & (g90) & (g82) & (g92) & (!g94)) + ((i_8_) & (g73) & (g90) & (g82) & (g92) & (g94)));
	assign g96 = (((!g87) & (!g78) & (!g74) & (!g79) & (!g89) & (!g95)) + ((!g87) & (!g78) & (!g74) & (!g79) & (g89) & (!g95)) + ((!g87) & (!g78) & (!g74) & (g79) & (!g89) & (!g95)) + ((!g87) & (!g78) & (!g74) & (g79) & (g89) & (!g95)) + ((!g87) & (g78) & (!g74) & (!g79) & (!g89) & (!g95)) + ((!g87) & (g78) & (!g74) & (!g79) & (g89) & (!g95)) + ((!g87) & (g78) & (!g74) & (g79) & (!g89) & (!g95)) + ((!g87) & (g78) & (!g74) & (g79) & (g89) & (!g95)) + ((g87) & (!g78) & (!g74) & (!g79) & (!g89) & (!g95)) + ((g87) & (!g78) & (!g74) & (!g79) & (g89) & (!g95)) + ((g87) & (!g78) & (!g74) & (g79) & (!g89) & (!g95)) + ((g87) & (!g78) & (!g74) & (g79) & (g89) & (!g95)) + ((g87) & (g78) & (!g74) & (!g79) & (!g89) & (!g95)) + ((g87) & (g78) & (!g74) & (!g79) & (g89) & (!g95)) + ((g87) & (g78) & (!g74) & (g79) & (!g89) & (!g95)) + ((g87) & (g78) & (!g74) & (g79) & (g89) & (!g95)) + ((g87) & (g78) & (g74) & (g79) & (g89) & (!g95)));
	assign g97 = (((!sk[127]) & (g17) & (g68)) + ((sk[127]) & (!g17) & (!g68)) + ((sk[127]) & (!g17) & (g68)) + ((sk[127]) & (g17) & (g68)));
	assign g98 = (((!sk[0]) & (g27) & (g76)) + ((sk[0]) & (g27) & (!g76)));
	assign g99 = (((!sk[1]) & (g73) & (g97) & (!g98)) + ((!sk[1]) & (g73) & (g97) & (g98)) + ((sk[1]) & (g73) & (!g97) & (!g98)) + ((sk[1]) & (g73) & (!g97) & (g98)) + ((sk[1]) & (g73) & (g97) & (g98)));
	assign g100 = (((!g70) & (!g74) & (!g85) & (g96) & (!sk[2]) & (!g99)) + ((!g70) & (!g74) & (!g85) & (g96) & (!sk[2]) & (g99)) + ((!g70) & (!g74) & (g85) & (!g96) & (!sk[2]) & (!g99)) + ((!g70) & (!g74) & (g85) & (!g96) & (!sk[2]) & (g99)) + ((!g70) & (!g74) & (g85) & (g96) & (!sk[2]) & (!g99)) + ((!g70) & (!g74) & (g85) & (g96) & (!sk[2]) & (g99)) + ((!g70) & (!g74) & (g85) & (g96) & (sk[2]) & (!g99)) + ((!g70) & (g74) & (!g85) & (g96) & (!sk[2]) & (!g99)) + ((!g70) & (g74) & (!g85) & (g96) & (!sk[2]) & (g99)) + ((!g70) & (g74) & (g85) & (!g96) & (!sk[2]) & (!g99)) + ((!g70) & (g74) & (g85) & (!g96) & (!sk[2]) & (g99)) + ((!g70) & (g74) & (g85) & (g96) & (!sk[2]) & (!g99)) + ((!g70) & (g74) & (g85) & (g96) & (!sk[2]) & (g99)) + ((!g70) & (g74) & (g85) & (g96) & (sk[2]) & (!g99)) + ((g70) & (!g74) & (!g85) & (g96) & (!sk[2]) & (!g99)) + ((g70) & (!g74) & (!g85) & (g96) & (!sk[2]) & (g99)) + ((g70) & (!g74) & (g85) & (!g96) & (!sk[2]) & (!g99)) + ((g70) & (!g74) & (g85) & (!g96) & (!sk[2]) & (g99)) + ((g70) & (!g74) & (g85) & (g96) & (!sk[2]) & (!g99)) + ((g70) & (!g74) & (g85) & (g96) & (!sk[2]) & (g99)) + ((g70) & (!g74) & (g85) & (g96) & (sk[2]) & (!g99)) + ((g70) & (g74) & (!g85) & (g96) & (!sk[2]) & (!g99)) + ((g70) & (g74) & (!g85) & (g96) & (!sk[2]) & (g99)) + ((g70) & (g74) & (g85) & (!g96) & (!sk[2]) & (!g99)) + ((g70) & (g74) & (g85) & (!g96) & (!sk[2]) & (g99)) + ((g70) & (g74) & (g85) & (g96) & (!sk[2]) & (!g99)) + ((g70) & (g74) & (g85) & (g96) & (!sk[2]) & (g99)));
	assign g101 = (((!sk[3]) & (i_8_) & (i_6_) & (!i_7_)) + ((!sk[3]) & (i_8_) & (i_6_) & (i_7_)) + ((sk[3]) & (!i_8_) & (i_6_) & (i_7_)));
	assign g102 = (((!sk[4]) & (g72) & (g101)) + ((sk[4]) & (g72) & (g101)));
	assign g103 = (((!g76) & (!sk[5]) & (!g102) & (!g82) & (g83)) + ((!g76) & (!sk[5]) & (!g102) & (g82) & (g83)) + ((!g76) & (!sk[5]) & (g102) & (!g82) & (g83)) + ((!g76) & (!sk[5]) & (g102) & (g82) & (g83)) + ((!g76) & (sk[5]) & (g102) & (!g82) & (g83)) + ((!g76) & (sk[5]) & (g102) & (g82) & (!g83)) + ((!g76) & (sk[5]) & (g102) & (g82) & (g83)) + ((g76) & (!sk[5]) & (!g102) & (!g82) & (g83)) + ((g76) & (!sk[5]) & (!g102) & (g82) & (g83)) + ((g76) & (!sk[5]) & (g102) & (!g82) & (!g83)) + ((g76) & (!sk[5]) & (g102) & (!g82) & (g83)) + ((g76) & (!sk[5]) & (g102) & (g82) & (!g83)) + ((g76) & (!sk[5]) & (g102) & (g82) & (g83)) + ((g76) & (sk[5]) & (g102) & (g82) & (!g83)) + ((g76) & (sk[5]) & (g102) & (g82) & (g83)));
	assign g104 = (((!sk[6]) & (g87) & (g102) & (!g89)) + ((!sk[6]) & (g87) & (g102) & (g89)) + ((sk[6]) & (!g87) & (g102) & (!g89)) + ((sk[6]) & (!g87) & (g102) & (g89)) + ((sk[6]) & (g87) & (g102) & (!g89)));
	assign g105 = (((!i_8_) & (!g45) & (sk[7]) & (!g72)) + ((!i_8_) & (!g45) & (sk[7]) & (g72)) + ((!i_8_) & (g45) & (!sk[7]) & (!g72)) + ((!i_8_) & (g45) & (!sk[7]) & (g72)) + ((!i_8_) & (g45) & (sk[7]) & (!g72)) + ((!i_8_) & (g45) & (sk[7]) & (g72)) + ((i_8_) & (!g45) & (!sk[7]) & (!g72)) + ((i_8_) & (!g45) & (!sk[7]) & (g72)) + ((i_8_) & (!g45) & (sk[7]) & (!g72)) + ((i_8_) & (!g45) & (sk[7]) & (g72)) + ((i_8_) & (g45) & (!sk[7]) & (!g72)) + ((i_8_) & (g45) & (!sk[7]) & (g72)) + ((i_8_) & (g45) & (sk[7]) & (!g72)));
	assign g106 = (((!sk[8]) & (g76) & (!g82) & (!g83) & (!g105)) + ((!sk[8]) & (g76) & (!g82) & (!g83) & (g105)) + ((!sk[8]) & (g76) & (!g82) & (g83) & (!g105)) + ((!sk[8]) & (g76) & (!g82) & (g83) & (g105)) + ((!sk[8]) & (g76) & (g82) & (!g83) & (!g105)) + ((!sk[8]) & (g76) & (g82) & (!g83) & (g105)) + ((!sk[8]) & (g76) & (g82) & (g83) & (!g105)) + ((!sk[8]) & (g76) & (g82) & (g83) & (g105)) + ((sk[8]) & (!g76) & (!g82) & (g83) & (!g105)) + ((sk[8]) & (!g76) & (g82) & (!g83) & (!g105)) + ((sk[8]) & (!g76) & (g82) & (g83) & (!g105)) + ((sk[8]) & (g76) & (g82) & (!g83) & (!g105)) + ((sk[8]) & (g76) & (g82) & (g83) & (!g105)));
	assign g107 = (((!i_11_) & (!sk[9]) & (i_15_) & (!g34)) + ((!i_11_) & (!sk[9]) & (i_15_) & (g34)) + ((!i_11_) & (sk[9]) & (!i_15_) & (!g34)) + ((!i_11_) & (sk[9]) & (!i_15_) & (g34)) + ((!i_11_) & (sk[9]) & (i_15_) & (!g34)) + ((!i_11_) & (sk[9]) & (i_15_) & (g34)) + ((i_11_) & (!sk[9]) & (!i_15_) & (!g34)) + ((i_11_) & (!sk[9]) & (!i_15_) & (g34)) + ((i_11_) & (!sk[9]) & (i_15_) & (!g34)) + ((i_11_) & (!sk[9]) & (i_15_) & (g34)) + ((i_11_) & (sk[9]) & (!i_15_) & (!g34)) + ((i_11_) & (sk[9]) & (i_15_) & (!g34)) + ((i_11_) & (sk[9]) & (i_15_) & (g34)));
	assign g108 = (((!sk[10]) & (g76) & (!g107)) + ((!sk[10]) & (g76) & (g107)) + ((sk[10]) & (!g76) & (!g107)));
	assign g109 = (((g35) & (!sk[11]) & (!g76)) + ((g35) & (!sk[11]) & (g76)) + ((g35) & (sk[11]) & (!g76)));
	assign g110 = (((!g108) & (!g109) & (!g90) & (!g98) & (g102) & (!g78)) + ((!g108) & (!g109) & (!g90) & (g98) & (g102) & (!g78)) + ((!g108) & (!g109) & (!g90) & (g98) & (g102) & (g78)) + ((!g108) & (!g109) & (g90) & (!g98) & (g102) & (!g78)) + ((!g108) & (!g109) & (g90) & (!g98) & (g102) & (g78)) + ((!g108) & (!g109) & (g90) & (g98) & (g102) & (!g78)) + ((!g108) & (!g109) & (g90) & (g98) & (g102) & (g78)) + ((!g108) & (g109) & (!g90) & (!g98) & (g102) & (!g78)) + ((!g108) & (g109) & (!g90) & (!g98) & (g102) & (g78)) + ((!g108) & (g109) & (!g90) & (g98) & (g102) & (!g78)) + ((!g108) & (g109) & (!g90) & (g98) & (g102) & (g78)) + ((!g108) & (g109) & (g90) & (!g98) & (g102) & (!g78)) + ((!g108) & (g109) & (g90) & (!g98) & (g102) & (g78)) + ((!g108) & (g109) & (g90) & (g98) & (g102) & (!g78)) + ((!g108) & (g109) & (g90) & (g98) & (g102) & (g78)) + ((g108) & (!g109) & (!g90) & (!g98) & (g102) & (!g78)) + ((g108) & (!g109) & (!g90) & (!g98) & (g102) & (g78)) + ((g108) & (!g109) & (!g90) & (g98) & (g102) & (!g78)) + ((g108) & (!g109) & (!g90) & (g98) & (g102) & (g78)) + ((g108) & (!g109) & (g90) & (!g98) & (g102) & (!g78)) + ((g108) & (!g109) & (g90) & (!g98) & (g102) & (g78)) + ((g108) & (!g109) & (g90) & (g98) & (g102) & (!g78)) + ((g108) & (!g109) & (g90) & (g98) & (g102) & (g78)) + ((g108) & (g109) & (!g90) & (!g98) & (g102) & (!g78)) + ((g108) & (g109) & (!g90) & (!g98) & (g102) & (g78)) + ((g108) & (g109) & (!g90) & (g98) & (g102) & (!g78)) + ((g108) & (g109) & (!g90) & (g98) & (g102) & (g78)) + ((g108) & (g109) & (g90) & (!g98) & (g102) & (!g78)) + ((g108) & (g109) & (g90) & (!g98) & (g102) & (g78)) + ((g108) & (g109) & (g90) & (g98) & (g102) & (!g78)) + ((g108) & (g109) & (g90) & (g98) & (g102) & (g78)));
	assign g111 = (((!sk[13]) & (g103) & (!g104) & (!g106) & (!g110)) + ((!sk[13]) & (g103) & (!g104) & (!g106) & (g110)) + ((!sk[13]) & (g103) & (!g104) & (g106) & (!g110)) + ((!sk[13]) & (g103) & (!g104) & (g106) & (g110)) + ((!sk[13]) & (g103) & (g104) & (!g106) & (!g110)) + ((!sk[13]) & (g103) & (g104) & (!g106) & (g110)) + ((!sk[13]) & (g103) & (g104) & (g106) & (!g110)) + ((!sk[13]) & (g103) & (g104) & (g106) & (g110)) + ((sk[13]) & (!g103) & (!g104) & (!g106) & (!g110)));
	assign g112 = (((!sk[14]) & (!i_9_) & (i_10_) & (!i_11_)) + ((!sk[14]) & (!i_9_) & (i_10_) & (i_11_)) + ((!sk[14]) & (i_9_) & (!i_10_) & (!i_11_)) + ((!sk[14]) & (i_9_) & (!i_10_) & (i_11_)) + ((!sk[14]) & (i_9_) & (i_10_) & (!i_11_)) + ((!sk[14]) & (i_9_) & (i_10_) & (i_11_)) + ((sk[14]) & (!i_9_) & (i_10_) & (i_11_)));
	assign g113 = (((!sk[15]) & (i_15_) & (!g112)) + ((!sk[15]) & (i_15_) & (g112)) + ((sk[15]) & (!i_15_) & (!g112)) + ((sk[15]) & (!i_15_) & (g112)) + ((sk[15]) & (i_15_) & (!g112)));
	assign g114 = (((!g68) & (sk[16]) & (g113)) + ((g68) & (!sk[16]) & (!g113)) + ((g68) & (!sk[16]) & (g113)) + ((g68) & (sk[16]) & (!g113)) + ((g68) & (sk[16]) & (g113)));
	assign g115 = (((!g109) & (!g90) & (sk[17]) & (g77) & (!g105)) + ((!g109) & (g90) & (sk[17]) & (!g77) & (!g105)) + ((!g109) & (g90) & (sk[17]) & (g77) & (!g105)) + ((g109) & (!g90) & (!sk[17]) & (!g77) & (!g105)) + ((g109) & (!g90) & (!sk[17]) & (!g77) & (g105)) + ((g109) & (!g90) & (!sk[17]) & (g77) & (!g105)) + ((g109) & (!g90) & (!sk[17]) & (g77) & (g105)) + ((g109) & (!g90) & (sk[17]) & (!g77) & (!g105)) + ((g109) & (!g90) & (sk[17]) & (g77) & (!g105)) + ((g109) & (g90) & (!sk[17]) & (!g77) & (!g105)) + ((g109) & (g90) & (!sk[17]) & (!g77) & (g105)) + ((g109) & (g90) & (!sk[17]) & (g77) & (!g105)) + ((g109) & (g90) & (!sk[17]) & (g77) & (g105)) + ((g109) & (g90) & (sk[17]) & (!g77) & (!g105)) + ((g109) & (g90) & (sk[17]) & (g77) & (!g105)));
	assign g116 = (((!g102) & (!sk[18]) & (!g92) & (g79) & (!g114) & (!g115)) + ((!g102) & (!sk[18]) & (!g92) & (g79) & (!g114) & (g115)) + ((!g102) & (!sk[18]) & (!g92) & (g79) & (g114) & (!g115)) + ((!g102) & (!sk[18]) & (!g92) & (g79) & (g114) & (g115)) + ((!g102) & (!sk[18]) & (g92) & (g79) & (!g114) & (!g115)) + ((!g102) & (!sk[18]) & (g92) & (g79) & (!g114) & (g115)) + ((!g102) & (!sk[18]) & (g92) & (g79) & (g114) & (!g115)) + ((!g102) & (!sk[18]) & (g92) & (g79) & (g114) & (g115)) + ((!g102) & (sk[18]) & (!g92) & (!g79) & (!g114) & (!g115)) + ((!g102) & (sk[18]) & (!g92) & (!g79) & (g114) & (!g115)) + ((!g102) & (sk[18]) & (!g92) & (g79) & (!g114) & (!g115)) + ((!g102) & (sk[18]) & (!g92) & (g79) & (g114) & (!g115)) + ((!g102) & (sk[18]) & (g92) & (!g79) & (!g114) & (!g115)) + ((!g102) & (sk[18]) & (g92) & (!g79) & (g114) & (!g115)) + ((!g102) & (sk[18]) & (g92) & (g79) & (!g114) & (!g115)) + ((!g102) & (sk[18]) & (g92) & (g79) & (g114) & (!g115)) + ((g102) & (!sk[18]) & (!g92) & (!g79) & (!g114) & (g115)) + ((g102) & (!sk[18]) & (!g92) & (!g79) & (g114) & (g115)) + ((g102) & (!sk[18]) & (!g92) & (g79) & (!g114) & (!g115)) + ((g102) & (!sk[18]) & (!g92) & (g79) & (!g114) & (g115)) + ((g102) & (!sk[18]) & (!g92) & (g79) & (g114) & (!g115)) + ((g102) & (!sk[18]) & (!g92) & (g79) & (g114) & (g115)) + ((g102) & (!sk[18]) & (g92) & (!g79) & (!g114) & (g115)) + ((g102) & (!sk[18]) & (g92) & (!g79) & (g114) & (g115)) + ((g102) & (!sk[18]) & (g92) & (g79) & (!g114) & (!g115)) + ((g102) & (!sk[18]) & (g92) & (g79) & (!g114) & (g115)) + ((g102) & (!sk[18]) & (g92) & (g79) & (g114) & (!g115)) + ((g102) & (!sk[18]) & (g92) & (g79) & (g114) & (g115)) + ((g102) & (sk[18]) & (!g92) & (g79) & (g114) & (!g115)));
	assign g117 = (((!sk[19]) & (g111) & (!g116)) + ((!sk[19]) & (g111) & (g116)) + ((sk[19]) & (g111) & (g116)));
	assign g118 = (((g6) & (!sk[20]) & (!g71)) + ((g6) & (!sk[20]) & (g71)) + ((g6) & (sk[20]) & (g71)));
	assign g119 = (((!sk[21]) & (!i_8_) & (g10) & (!g118)) + ((!sk[21]) & (!i_8_) & (g10) & (g118)) + ((!sk[21]) & (i_8_) & (!g10) & (!g118)) + ((!sk[21]) & (i_8_) & (!g10) & (g118)) + ((!sk[21]) & (i_8_) & (g10) & (!g118)) + ((!sk[21]) & (i_8_) & (g10) & (g118)) + ((sk[21]) & (i_8_) & (g10) & (g118)));
	assign g120 = (((!sk[22]) & (g54) & (!g71)) + ((!sk[22]) & (g54) & (g71)) + ((sk[22]) & (g54) & (g71)));
	assign g121 = (((!i_8_) & (g45) & (!sk[23]) & (!g120)) + ((!i_8_) & (g45) & (!sk[23]) & (g120)) + ((i_8_) & (!g45) & (!sk[23]) & (!g120)) + ((i_8_) & (!g45) & (!sk[23]) & (g120)) + ((i_8_) & (g45) & (!sk[23]) & (!g120)) + ((i_8_) & (g45) & (!sk[23]) & (g120)) + ((i_8_) & (g45) & (sk[23]) & (g120)));
	assign g122 = (((!sk[24]) & (g49) & (!g118)) + ((!sk[24]) & (g49) & (g118)) + ((sk[24]) & (g49) & (g118)));
	assign g123 = (((!sk[25]) & (g30) & (!g118)) + ((!sk[25]) & (g30) & (g118)) + ((sk[25]) & (!g30) & (!g118)) + ((sk[25]) & (!g30) & (g118)) + ((sk[25]) & (g30) & (!g118)));
	assign g124 = (((!g70) & (g122) & (sk[26]) & (!g123) & (!g114)) + ((!g70) & (g122) & (sk[26]) & (g123) & (!g114)) + ((g70) & (!g122) & (!sk[26]) & (!g123) & (!g114)) + ((g70) & (!g122) & (!sk[26]) & (!g123) & (g114)) + ((g70) & (!g122) & (!sk[26]) & (g123) & (!g114)) + ((g70) & (!g122) & (!sk[26]) & (g123) & (g114)) + ((g70) & (!g122) & (sk[26]) & (!g123) & (!g114)) + ((g70) & (!g122) & (sk[26]) & (!g123) & (g114)) + ((g70) & (g122) & (!sk[26]) & (!g123) & (!g114)) + ((g70) & (g122) & (!sk[26]) & (!g123) & (g114)) + ((g70) & (g122) & (!sk[26]) & (g123) & (!g114)) + ((g70) & (g122) & (!sk[26]) & (g123) & (g114)) + ((g70) & (g122) & (sk[26]) & (!g123) & (!g114)) + ((g70) & (g122) & (sk[26]) & (!g123) & (g114)) + ((g70) & (g122) & (sk[26]) & (g123) & (!g114)));
	assign g125 = (((g49) & (!sk[27]) & (!g120)) + ((g49) & (!sk[27]) & (g120)) + ((g49) & (sk[27]) & (g120)));
	assign g126 = (((!i_15_) & (sk[28]) & (!g112)) + ((i_15_) & (!sk[28]) & (!g112)) + ((i_15_) & (!sk[28]) & (g112)) + ((i_15_) & (sk[28]) & (!g112)) + ((i_15_) & (sk[28]) & (g112)));
	assign g127 = (((!sk[29]) & (g76) & (!g126)) + ((!sk[29]) & (g76) & (g126)) + ((sk[29]) & (!g76) & (!g126)));
	assign g128 = (((!g125) & (!g77) & (!sk[30]) & (g127) & (!g123) & (!g119)) + ((!g125) & (!g77) & (!sk[30]) & (g127) & (!g123) & (g119)) + ((!g125) & (!g77) & (!sk[30]) & (g127) & (g123) & (!g119)) + ((!g125) & (!g77) & (!sk[30]) & (g127) & (g123) & (g119)) + ((!g125) & (!g77) & (sk[30]) & (!g127) & (!g123) & (!g119)) + ((!g125) & (!g77) & (sk[30]) & (!g127) & (!g123) & (g119)) + ((!g125) & (!g77) & (sk[30]) & (!g127) & (g123) & (!g119)) + ((!g125) & (!g77) & (sk[30]) & (!g127) & (g123) & (g119)) + ((!g125) & (!g77) & (sk[30]) & (g127) & (!g123) & (!g119)) + ((!g125) & (!g77) & (sk[30]) & (g127) & (!g123) & (g119)) + ((!g125) & (!g77) & (sk[30]) & (g127) & (g123) & (!g119)) + ((!g125) & (!g77) & (sk[30]) & (g127) & (g123) & (g119)) + ((!g125) & (g77) & (!sk[30]) & (g127) & (!g123) & (!g119)) + ((!g125) & (g77) & (!sk[30]) & (g127) & (!g123) & (g119)) + ((!g125) & (g77) & (!sk[30]) & (g127) & (g123) & (!g119)) + ((!g125) & (g77) & (!sk[30]) & (g127) & (g123) & (g119)) + ((!g125) & (g77) & (sk[30]) & (!g127) & (g123) & (!g119)) + ((!g125) & (g77) & (sk[30]) & (g127) & (g123) & (!g119)) + ((g125) & (!g77) & (!sk[30]) & (!g127) & (!g123) & (g119)) + ((g125) & (!g77) & (!sk[30]) & (!g127) & (g123) & (g119)) + ((g125) & (!g77) & (!sk[30]) & (g127) & (!g123) & (!g119)) + ((g125) & (!g77) & (!sk[30]) & (g127) & (!g123) & (g119)) + ((g125) & (!g77) & (!sk[30]) & (g127) & (g123) & (!g119)) + ((g125) & (!g77) & (!sk[30]) & (g127) & (g123) & (g119)) + ((g125) & (!g77) & (sk[30]) & (!g127) & (!g123) & (!g119)) + ((g125) & (!g77) & (sk[30]) & (!g127) & (!g123) & (g119)) + ((g125) & (!g77) & (sk[30]) & (!g127) & (g123) & (!g119)) + ((g125) & (!g77) & (sk[30]) & (!g127) & (g123) & (g119)) + ((g125) & (g77) & (!sk[30]) & (!g127) & (!g123) & (g119)) + ((g125) & (g77) & (!sk[30]) & (!g127) & (g123) & (g119)) + ((g125) & (g77) & (!sk[30]) & (g127) & (!g123) & (!g119)) + ((g125) & (g77) & (!sk[30]) & (g127) & (!g123) & (g119)) + ((g125) & (g77) & (!sk[30]) & (g127) & (g123) & (!g119)) + ((g125) & (g77) & (!sk[30]) & (g127) & (g123) & (g119)) + ((g125) & (g77) & (sk[30]) & (!g127) & (g123) & (!g119)));
	assign g129 = (((!g70) & (!g119) & (!g121) & (!g124) & (sk[31]) & (g128)) + ((!g70) & (!g119) & (g121) & (!g124) & (!sk[31]) & (!g128)) + ((!g70) & (!g119) & (g121) & (!g124) & (!sk[31]) & (g128)) + ((!g70) & (!g119) & (g121) & (!g124) & (sk[31]) & (g128)) + ((!g70) & (!g119) & (g121) & (g124) & (!sk[31]) & (!g128)) + ((!g70) & (!g119) & (g121) & (g124) & (!sk[31]) & (g128)) + ((!g70) & (g119) & (!g121) & (!g124) & (sk[31]) & (g128)) + ((!g70) & (g119) & (g121) & (!g124) & (!sk[31]) & (!g128)) + ((!g70) & (g119) & (g121) & (!g124) & (!sk[31]) & (g128)) + ((!g70) & (g119) & (g121) & (!g124) & (sk[31]) & (g128)) + ((!g70) & (g119) & (g121) & (g124) & (!sk[31]) & (!g128)) + ((!g70) & (g119) & (g121) & (g124) & (!sk[31]) & (g128)) + ((g70) & (!g119) & (!g121) & (!g124) & (!sk[31]) & (g128)) + ((g70) & (!g119) & (!g121) & (!g124) & (sk[31]) & (g128)) + ((g70) & (!g119) & (!g121) & (g124) & (!sk[31]) & (g128)) + ((g70) & (!g119) & (g121) & (!g124) & (!sk[31]) & (!g128)) + ((g70) & (!g119) & (g121) & (!g124) & (!sk[31]) & (g128)) + ((g70) & (!g119) & (g121) & (g124) & (!sk[31]) & (!g128)) + ((g70) & (!g119) & (g121) & (g124) & (!sk[31]) & (g128)) + ((g70) & (g119) & (!g121) & (!g124) & (!sk[31]) & (g128)) + ((g70) & (g119) & (!g121) & (g124) & (!sk[31]) & (g128)) + ((g70) & (g119) & (g121) & (!g124) & (!sk[31]) & (!g128)) + ((g70) & (g119) & (g121) & (!g124) & (!sk[31]) & (g128)) + ((g70) & (g119) & (g121) & (g124) & (!sk[31]) & (!g128)) + ((g70) & (g119) & (g121) & (g124) & (!sk[31]) & (g128)));
	assign g130 = (((!sk[32]) & (g2) & (!g118)) + ((!sk[32]) & (g2) & (g118)) + ((sk[32]) & (!g2) & (!g118)) + ((sk[32]) & (!g2) & (g118)) + ((sk[32]) & (g2) & (!g118)));
	assign g131 = (((!sk[33]) & (g43) & (!g120)) + ((!sk[33]) & (g43) & (g120)) + ((sk[33]) & (!g43) & (!g120)) + ((sk[33]) & (!g43) & (g120)) + ((sk[33]) & (g43) & (!g120)));
	assign g132 = (((!i_8_) & (!g73) & (!g108) & (sk[34]) & (!g92) & (g1639)) + ((!i_8_) & (!g73) & (!g108) & (sk[34]) & (g92) & (g1639)) + ((!i_8_) & (!g73) & (g108) & (!sk[34]) & (!g92) & (!g1639)) + ((!i_8_) & (!g73) & (g108) & (!sk[34]) & (!g92) & (g1639)) + ((!i_8_) & (!g73) & (g108) & (!sk[34]) & (g92) & (!g1639)) + ((!i_8_) & (!g73) & (g108) & (!sk[34]) & (g92) & (g1639)) + ((!i_8_) & (!g73) & (g108) & (sk[34]) & (!g92) & (g1639)) + ((!i_8_) & (!g73) & (g108) & (sk[34]) & (g92) & (g1639)) + ((!i_8_) & (g73) & (!g108) & (sk[34]) & (!g92) & (g1639)) + ((!i_8_) & (g73) & (!g108) & (sk[34]) & (g92) & (g1639)) + ((!i_8_) & (g73) & (g108) & (!sk[34]) & (!g92) & (!g1639)) + ((!i_8_) & (g73) & (g108) & (!sk[34]) & (!g92) & (g1639)) + ((!i_8_) & (g73) & (g108) & (!sk[34]) & (g92) & (!g1639)) + ((!i_8_) & (g73) & (g108) & (!sk[34]) & (g92) & (g1639)) + ((i_8_) & (!g73) & (!g108) & (!sk[34]) & (!g92) & (g1639)) + ((i_8_) & (!g73) & (!g108) & (!sk[34]) & (g92) & (g1639)) + ((i_8_) & (!g73) & (!g108) & (sk[34]) & (!g92) & (g1639)) + ((i_8_) & (!g73) & (!g108) & (sk[34]) & (g92) & (g1639)) + ((i_8_) & (!g73) & (g108) & (!sk[34]) & (!g92) & (!g1639)) + ((i_8_) & (!g73) & (g108) & (!sk[34]) & (!g92) & (g1639)) + ((i_8_) & (!g73) & (g108) & (!sk[34]) & (g92) & (!g1639)) + ((i_8_) & (!g73) & (g108) & (!sk[34]) & (g92) & (g1639)) + ((i_8_) & (!g73) & (g108) & (sk[34]) & (!g92) & (g1639)) + ((i_8_) & (!g73) & (g108) & (sk[34]) & (g92) & (g1639)) + ((i_8_) & (g73) & (!g108) & (!sk[34]) & (!g92) & (g1639)) + ((i_8_) & (g73) & (!g108) & (!sk[34]) & (g92) & (g1639)) + ((i_8_) & (g73) & (!g108) & (sk[34]) & (!g92) & (g1639)) + ((i_8_) & (g73) & (g108) & (!sk[34]) & (!g92) & (!g1639)) + ((i_8_) & (g73) & (g108) & (!sk[34]) & (!g92) & (g1639)) + ((i_8_) & (g73) & (g108) & (!sk[34]) & (g92) & (!g1639)) + ((i_8_) & (g73) & (g108) & (!sk[34]) & (g92) & (g1639)) + ((i_8_) & (g73) & (g108) & (sk[34]) & (!g92) & (g1639)));
	assign g133 = (((!g108) & (!sk[35]) & (g92) & (!g123)) + ((!g108) & (!sk[35]) & (g92) & (g123)) + ((!g108) & (sk[35]) & (g92) & (!g123)) + ((g108) & (!sk[35]) & (!g92) & (!g123)) + ((g108) & (!sk[35]) & (!g92) & (g123)) + ((g108) & (!sk[35]) & (g92) & (!g123)) + ((g108) & (!sk[35]) & (g92) & (g123)) + ((g108) & (sk[35]) & (!g92) & (!g123)) + ((g108) & (sk[35]) & (g92) & (!g123)));
	assign g134 = (((!g108) & (g92) & (!sk[36]) & (!g130)) + ((!g108) & (g92) & (!sk[36]) & (g130)) + ((!g108) & (g92) & (sk[36]) & (!g130)) + ((g108) & (!g92) & (!sk[36]) & (!g130)) + ((g108) & (!g92) & (!sk[36]) & (g130)) + ((g108) & (!g92) & (sk[36]) & (!g130)) + ((g108) & (g92) & (!sk[36]) & (!g130)) + ((g108) & (g92) & (!sk[36]) & (g130)) + ((g108) & (g92) & (sk[36]) & (!g130)));
	assign g135 = (((!g43) & (sk[37]) & (!g118)) + ((!g43) & (sk[37]) & (g118)) + ((g43) & (!sk[37]) & (!g118)) + ((g43) & (!sk[37]) & (g118)) + ((g43) & (sk[37]) & (!g118)));
	assign g136 = (((!g76) & (g122) & (sk[38]) & (!g82) & (g83)) + ((!g76) & (g122) & (sk[38]) & (g82) & (!g83)) + ((!g76) & (g122) & (sk[38]) & (g82) & (g83)) + ((g76) & (!g122) & (!sk[38]) & (!g82) & (!g83)) + ((g76) & (!g122) & (!sk[38]) & (!g82) & (g83)) + ((g76) & (!g122) & (!sk[38]) & (g82) & (!g83)) + ((g76) & (!g122) & (!sk[38]) & (g82) & (g83)) + ((g76) & (g122) & (!sk[38]) & (!g82) & (!g83)) + ((g76) & (g122) & (!sk[38]) & (!g82) & (g83)) + ((g76) & (g122) & (!sk[38]) & (g82) & (!g83)) + ((g76) & (g122) & (!sk[38]) & (g82) & (g83)) + ((g76) & (g122) & (sk[38]) & (g82) & (!g83)) + ((g76) & (g122) & (sk[38]) & (g82) & (g83)));
	assign g137 = (((!sk[39]) & (g78) & (!g135) & (!g122) & (!g89)) + ((!sk[39]) & (g78) & (!g135) & (!g122) & (g89)) + ((!sk[39]) & (g78) & (!g135) & (g122) & (!g89)) + ((!sk[39]) & (g78) & (!g135) & (g122) & (g89)) + ((!sk[39]) & (g78) & (g135) & (!g122) & (!g89)) + ((!sk[39]) & (g78) & (g135) & (!g122) & (g89)) + ((!sk[39]) & (g78) & (g135) & (g122) & (!g89)) + ((!sk[39]) & (g78) & (g135) & (g122) & (g89)) + ((sk[39]) & (!g78) & (!g135) & (!g122) & (!g89)) + ((sk[39]) & (!g78) & (!g135) & (g122) & (!g89)) + ((sk[39]) & (!g78) & (!g135) & (g122) & (g89)) + ((sk[39]) & (!g78) & (g135) & (g122) & (!g89)) + ((sk[39]) & (!g78) & (g135) & (g122) & (g89)) + ((sk[39]) & (g78) & (!g135) & (!g122) & (!g89)) + ((sk[39]) & (g78) & (!g135) & (g122) & (!g89)));
	assign g138 = (((!g97) & (!g98) & (g135) & (!g122) & (!g136) & (!g137)) + ((!g97) & (g98) & (g135) & (!g122) & (!g136) & (!g137)) + ((g97) & (!g98) & (!g135) & (!g122) & (!g136) & (!g137)) + ((g97) & (!g98) & (!g135) & (g122) & (!g136) & (!g137)) + ((g97) & (!g98) & (g135) & (!g122) & (!g136) & (!g137)) + ((g97) & (!g98) & (g135) & (g122) & (!g136) & (!g137)) + ((g97) & (g98) & (g135) & (!g122) & (!g136) & (!g137)));
	assign g139 = (((!sk[41]) & (g76) & (!g82) & (!g83) & (!g130)) + ((!sk[41]) & (g76) & (!g82) & (!g83) & (g130)) + ((!sk[41]) & (g76) & (!g82) & (g83) & (!g130)) + ((!sk[41]) & (g76) & (!g82) & (g83) & (g130)) + ((!sk[41]) & (g76) & (g82) & (!g83) & (!g130)) + ((!sk[41]) & (g76) & (g82) & (!g83) & (g130)) + ((!sk[41]) & (g76) & (g82) & (g83) & (!g130)) + ((!sk[41]) & (g76) & (g82) & (g83) & (g130)) + ((sk[41]) & (!g76) & (!g82) & (g83) & (!g130)) + ((sk[41]) & (!g76) & (g82) & (!g83) & (!g130)) + ((sk[41]) & (!g76) & (g82) & (g83) & (!g130)) + ((sk[41]) & (g76) & (g82) & (!g83) & (!g130)) + ((sk[41]) & (g76) & (g82) & (g83) & (!g130)));
	assign g140 = (((!g109) & (g90) & (!sk[42]) & (!g130)) + ((!g109) & (g90) & (!sk[42]) & (g130)) + ((!g109) & (g90) & (sk[42]) & (!g130)) + ((g109) & (!g90) & (!sk[42]) & (!g130)) + ((g109) & (!g90) & (!sk[42]) & (g130)) + ((g109) & (!g90) & (sk[42]) & (!g130)) + ((g109) & (g90) & (!sk[42]) & (!g130)) + ((g109) & (g90) & (!sk[42]) & (g130)) + ((g109) & (g90) & (sk[42]) & (!g130)));
	assign g141 = (((!sk[43]) & (g87) & (!g127) & (!g79) & (!g123)) + ((!sk[43]) & (g87) & (!g127) & (!g79) & (g123)) + ((!sk[43]) & (g87) & (!g127) & (g79) & (!g123)) + ((!sk[43]) & (g87) & (!g127) & (g79) & (g123)) + ((!sk[43]) & (g87) & (g127) & (!g79) & (!g123)) + ((!sk[43]) & (g87) & (g127) & (!g79) & (g123)) + ((!sk[43]) & (g87) & (g127) & (g79) & (!g123)) + ((!sk[43]) & (g87) & (g127) & (g79) & (g123)) + ((sk[43]) & (!g87) & (!g127) & (!g79) & (!g123)) + ((sk[43]) & (!g87) & (!g127) & (g79) & (!g123)) + ((sk[43]) & (!g87) & (g127) & (!g79) & (!g123)) + ((sk[43]) & (!g87) & (g127) & (g79) & (!g123)) + ((sk[43]) & (g87) & (!g127) & (!g79) & (!g123)) + ((sk[43]) & (g87) & (g127) & (!g79) & (!g123)) + ((sk[43]) & (g87) & (g127) & (g79) & (!g123)));
	assign g142 = (((!sk[44]) & (!i_8_) & (g10) & (!g118)) + ((!sk[44]) & (!i_8_) & (g10) & (g118)) + ((!sk[44]) & (i_8_) & (!g10) & (!g118)) + ((!sk[44]) & (i_8_) & (!g10) & (g118)) + ((!sk[44]) & (i_8_) & (g10) & (!g118)) + ((!sk[44]) & (i_8_) & (g10) & (g118)) + ((sk[44]) & (!i_8_) & (!g10) & (!g118)) + ((sk[44]) & (!i_8_) & (!g10) & (g118)) + ((sk[44]) & (!i_8_) & (g10) & (!g118)) + ((sk[44]) & (i_8_) & (!g10) & (!g118)) + ((sk[44]) & (i_8_) & (!g10) & (g118)) + ((sk[44]) & (i_8_) & (g10) & (!g118)) + ((sk[44]) & (i_8_) & (g10) & (g118)));
	assign g143 = (((!g97) & (!g82) & (sk[45]) & (!g142)) + ((!g97) & (g82) & (!sk[45]) & (!g142)) + ((!g97) & (g82) & (!sk[45]) & (g142)) + ((!g97) & (g82) & (sk[45]) & (!g142)) + ((g97) & (!g82) & (!sk[45]) & (!g142)) + ((g97) & (!g82) & (!sk[45]) & (g142)) + ((g97) & (g82) & (!sk[45]) & (!g142)) + ((g97) & (g82) & (!sk[45]) & (g142)) + ((g97) & (g82) & (sk[45]) & (!g142)));
	assign g144 = (((!sk[46]) & (g42) & (!g120)) + ((!sk[46]) & (g42) & (g120)) + ((sk[46]) & (g42) & (g120)));
	assign g145 = (((!g87) & (!g144) & (!g122) & (!g89) & (sk[47]) & (g105)) + ((!g87) & (!g144) & (!g122) & (g89) & (sk[47]) & (g105)) + ((!g87) & (!g144) & (g122) & (!g89) & (!sk[47]) & (!g105)) + ((!g87) & (!g144) & (g122) & (!g89) & (!sk[47]) & (g105)) + ((!g87) & (!g144) & (g122) & (g89) & (!sk[47]) & (!g105)) + ((!g87) & (!g144) & (g122) & (g89) & (!sk[47]) & (g105)) + ((!g87) & (!g144) & (g122) & (g89) & (sk[47]) & (g105)) + ((!g87) & (g144) & (!g122) & (g89) & (sk[47]) & (g105)) + ((!g87) & (g144) & (g122) & (!g89) & (!sk[47]) & (!g105)) + ((!g87) & (g144) & (g122) & (!g89) & (!sk[47]) & (g105)) + ((!g87) & (g144) & (g122) & (g89) & (!sk[47]) & (!g105)) + ((!g87) & (g144) & (g122) & (g89) & (!sk[47]) & (g105)) + ((!g87) & (g144) & (g122) & (g89) & (sk[47]) & (g105)) + ((g87) & (!g144) & (!g122) & (!g89) & (!sk[47]) & (g105)) + ((g87) & (!g144) & (!g122) & (!g89) & (sk[47]) & (g105)) + ((g87) & (!g144) & (!g122) & (g89) & (!sk[47]) & (g105)) + ((g87) & (!g144) & (!g122) & (g89) & (sk[47]) & (!g105)) + ((g87) & (!g144) & (!g122) & (g89) & (sk[47]) & (g105)) + ((g87) & (!g144) & (g122) & (!g89) & (!sk[47]) & (!g105)) + ((g87) & (!g144) & (g122) & (!g89) & (!sk[47]) & (g105)) + ((g87) & (!g144) & (g122) & (g89) & (!sk[47]) & (!g105)) + ((g87) & (!g144) & (g122) & (g89) & (!sk[47]) & (g105)) + ((g87) & (!g144) & (g122) & (g89) & (sk[47]) & (!g105)) + ((g87) & (!g144) & (g122) & (g89) & (sk[47]) & (g105)) + ((g87) & (g144) & (!g122) & (!g89) & (!sk[47]) & (g105)) + ((g87) & (g144) & (!g122) & (g89) & (!sk[47]) & (g105)) + ((g87) & (g144) & (!g122) & (g89) & (sk[47]) & (!g105)) + ((g87) & (g144) & (!g122) & (g89) & (sk[47]) & (g105)) + ((g87) & (g144) & (g122) & (!g89) & (!sk[47]) & (!g105)) + ((g87) & (g144) & (g122) & (!g89) & (!sk[47]) & (g105)) + ((g87) & (g144) & (g122) & (g89) & (!sk[47]) & (!g105)) + ((g87) & (g144) & (g122) & (g89) & (!sk[47]) & (g105)) + ((g87) & (g144) & (g122) & (g89) & (sk[47]) & (!g105)) + ((g87) & (g144) & (g122) & (g89) & (sk[47]) & (g105)));
	assign g146 = (((!sk[48]) & (!g139) & (!g140) & (g141) & (!g143) & (!g145)) + ((!sk[48]) & (!g139) & (!g140) & (g141) & (!g143) & (g145)) + ((!sk[48]) & (!g139) & (!g140) & (g141) & (g143) & (!g145)) + ((!sk[48]) & (!g139) & (!g140) & (g141) & (g143) & (g145)) + ((!sk[48]) & (!g139) & (g140) & (g141) & (!g143) & (!g145)) + ((!sk[48]) & (!g139) & (g140) & (g141) & (!g143) & (g145)) + ((!sk[48]) & (!g139) & (g140) & (g141) & (g143) & (!g145)) + ((!sk[48]) & (!g139) & (g140) & (g141) & (g143) & (g145)) + ((!sk[48]) & (g139) & (!g140) & (!g141) & (!g143) & (g145)) + ((!sk[48]) & (g139) & (!g140) & (!g141) & (g143) & (g145)) + ((!sk[48]) & (g139) & (!g140) & (g141) & (!g143) & (!g145)) + ((!sk[48]) & (g139) & (!g140) & (g141) & (!g143) & (g145)) + ((!sk[48]) & (g139) & (!g140) & (g141) & (g143) & (!g145)) + ((!sk[48]) & (g139) & (!g140) & (g141) & (g143) & (g145)) + ((!sk[48]) & (g139) & (g140) & (!g141) & (!g143) & (g145)) + ((!sk[48]) & (g139) & (g140) & (!g141) & (g143) & (g145)) + ((!sk[48]) & (g139) & (g140) & (g141) & (!g143) & (!g145)) + ((!sk[48]) & (g139) & (g140) & (g141) & (!g143) & (g145)) + ((!sk[48]) & (g139) & (g140) & (g141) & (g143) & (!g145)) + ((!sk[48]) & (g139) & (g140) & (g141) & (g143) & (g145)) + ((sk[48]) & (!g139) & (!g140) & (!g141) & (!g143) & (g145)));
	assign g147 = (((!sk[49]) & (!g109) & (g90) & (!g123)) + ((!sk[49]) & (!g109) & (g90) & (g123)) + ((!sk[49]) & (g109) & (!g90) & (!g123)) + ((!sk[49]) & (g109) & (!g90) & (g123)) + ((!sk[49]) & (g109) & (g90) & (!g123)) + ((!sk[49]) & (g109) & (g90) & (g123)) + ((sk[49]) & (!g109) & (g90) & (!g123)) + ((sk[49]) & (g109) & (!g90) & (!g123)) + ((sk[49]) & (g109) & (g90) & (!g123)));
	assign g148 = (((!g97) & (!g98) & (sk[50]) & (!g105)) + ((!g97) & (g98) & (!sk[50]) & (!g105)) + ((!g97) & (g98) & (!sk[50]) & (g105)) + ((!g97) & (g98) & (sk[50]) & (!g105)) + ((g97) & (!g98) & (!sk[50]) & (!g105)) + ((g97) & (!g98) & (!sk[50]) & (g105)) + ((g97) & (g98) & (!sk[50]) & (!g105)) + ((g97) & (g98) & (!sk[50]) & (g105)) + ((g97) & (g98) & (sk[50]) & (!g105)));
	assign g149 = (((!g127) & (!g78) & (!g135) & (!g79) & (g114) & (g105)) + ((!g127) & (!g78) & (!g135) & (g79) & (g114) & (g105)) + ((!g127) & (!g78) & (g135) & (!g79) & (!g114) & (g105)) + ((!g127) & (!g78) & (g135) & (!g79) & (g114) & (g105)) + ((!g127) & (!g78) & (g135) & (g79) & (!g114) & (g105)) + ((!g127) & (!g78) & (g135) & (g79) & (g114) & (g105)) + ((!g127) & (g78) & (!g135) & (!g79) & (g114) & (g105)) + ((!g127) & (g78) & (!g135) & (g79) & (g114) & (!g105)) + ((!g127) & (g78) & (!g135) & (g79) & (g114) & (g105)) + ((!g127) & (g78) & (g135) & (!g79) & (!g114) & (g105)) + ((!g127) & (g78) & (g135) & (!g79) & (g114) & (g105)) + ((!g127) & (g78) & (g135) & (g79) & (!g114) & (g105)) + ((!g127) & (g78) & (g135) & (g79) & (g114) & (!g105)) + ((!g127) & (g78) & (g135) & (g79) & (g114) & (g105)) + ((g127) & (!g78) & (!g135) & (!g79) & (g114) & (g105)) + ((g127) & (!g78) & (!g135) & (g79) & (g114) & (g105)) + ((g127) & (!g78) & (g135) & (!g79) & (!g114) & (g105)) + ((g127) & (!g78) & (g135) & (!g79) & (g114) & (g105)) + ((g127) & (!g78) & (g135) & (g79) & (!g114) & (g105)) + ((g127) & (!g78) & (g135) & (g79) & (g114) & (g105)) + ((g127) & (g78) & (!g135) & (!g79) & (g114) & (g105)) + ((g127) & (g78) & (!g135) & (g79) & (g114) & (g105)) + ((g127) & (g78) & (g135) & (!g79) & (!g114) & (g105)) + ((g127) & (g78) & (g135) & (!g79) & (g114) & (g105)) + ((g127) & (g78) & (g135) & (g79) & (!g114) & (g105)) + ((g127) & (g78) & (g135) & (g79) & (g114) & (g105)));
	assign g150 = (((!g77) & (!g97) & (!g102) & (!g147) & (!g148) & (g149)) + ((!g77) & (g97) & (!g102) & (!g147) & (!g148) & (g149)) + ((!g77) & (g97) & (g102) & (!g147) & (!g148) & (g149)) + ((g77) & (!g97) & (!g102) & (!g147) & (!g148) & (g149)) + ((g77) & (g97) & (!g102) & (!g147) & (!g148) & (g149)));
	assign g151 = (((!i_9_) & (!i_10_) & (sk[53]) & (i_11_) & (!g142)) + ((i_9_) & (!i_10_) & (!sk[53]) & (!i_11_) & (!g142)) + ((i_9_) & (!i_10_) & (!sk[53]) & (!i_11_) & (g142)) + ((i_9_) & (!i_10_) & (!sk[53]) & (i_11_) & (!g142)) + ((i_9_) & (!i_10_) & (!sk[53]) & (i_11_) & (g142)) + ((i_9_) & (!i_10_) & (sk[53]) & (!i_11_) & (!g142)) + ((i_9_) & (i_10_) & (!sk[53]) & (!i_11_) & (!g142)) + ((i_9_) & (i_10_) & (!sk[53]) & (!i_11_) & (g142)) + ((i_9_) & (i_10_) & (!sk[53]) & (i_11_) & (!g142)) + ((i_9_) & (i_10_) & (!sk[53]) & (i_11_) & (g142)));
	assign g152 = (((!g73) & (!g127) & (!g93) & (sk[54]) & (!g114) & (!g151)) + ((!g73) & (!g127) & (!g93) & (sk[54]) & (!g114) & (g151)) + ((!g73) & (!g127) & (!g93) & (sk[54]) & (g114) & (!g151)) + ((!g73) & (!g127) & (!g93) & (sk[54]) & (g114) & (g151)) + ((!g73) & (!g127) & (g93) & (!sk[54]) & (!g114) & (!g151)) + ((!g73) & (!g127) & (g93) & (!sk[54]) & (!g114) & (g151)) + ((!g73) & (!g127) & (g93) & (!sk[54]) & (g114) & (!g151)) + ((!g73) & (!g127) & (g93) & (!sk[54]) & (g114) & (g151)) + ((!g73) & (!g127) & (g93) & (sk[54]) & (!g114) & (!g151)) + ((!g73) & (!g127) & (g93) & (sk[54]) & (g114) & (!g151)) + ((!g73) & (g127) & (!g93) & (sk[54]) & (!g114) & (!g151)) + ((!g73) & (g127) & (!g93) & (sk[54]) & (!g114) & (g151)) + ((!g73) & (g127) & (!g93) & (sk[54]) & (g114) & (!g151)) + ((!g73) & (g127) & (!g93) & (sk[54]) & (g114) & (g151)) + ((!g73) & (g127) & (g93) & (!sk[54]) & (!g114) & (!g151)) + ((!g73) & (g127) & (g93) & (!sk[54]) & (!g114) & (g151)) + ((!g73) & (g127) & (g93) & (!sk[54]) & (g114) & (!g151)) + ((!g73) & (g127) & (g93) & (!sk[54]) & (g114) & (g151)) + ((!g73) & (g127) & (g93) & (sk[54]) & (!g114) & (!g151)) + ((!g73) & (g127) & (g93) & (sk[54]) & (g114) & (!g151)) + ((g73) & (!g127) & (!g93) & (!sk[54]) & (!g114) & (g151)) + ((g73) & (!g127) & (!g93) & (!sk[54]) & (g114) & (g151)) + ((g73) & (!g127) & (!g93) & (sk[54]) & (g114) & (!g151)) + ((g73) & (!g127) & (!g93) & (sk[54]) & (g114) & (g151)) + ((g73) & (!g127) & (g93) & (!sk[54]) & (!g114) & (!g151)) + ((g73) & (!g127) & (g93) & (!sk[54]) & (!g114) & (g151)) + ((g73) & (!g127) & (g93) & (!sk[54]) & (g114) & (!g151)) + ((g73) & (!g127) & (g93) & (!sk[54]) & (g114) & (g151)) + ((g73) & (!g127) & (g93) & (sk[54]) & (g114) & (!g151)) + ((g73) & (g127) & (!g93) & (!sk[54]) & (!g114) & (g151)) + ((g73) & (g127) & (!g93) & (!sk[54]) & (g114) & (g151)) + ((g73) & (g127) & (g93) & (!sk[54]) & (!g114) & (!g151)) + ((g73) & (g127) & (g93) & (!sk[54]) & (!g114) & (g151)) + ((g73) & (g127) & (g93) & (!sk[54]) & (g114) & (!g151)) + ((g73) & (g127) & (g93) & (!sk[54]) & (g114) & (g151)));
	assign g153 = (((!g133) & (!g134) & (g138) & (g146) & (g150) & (g152)));
	assign g154 = (((!i_8_) & (!g10) & (sk[56]) & (!g120)) + ((!i_8_) & (!g10) & (sk[56]) & (g120)) + ((!i_8_) & (g10) & (!sk[56]) & (!g120)) + ((!i_8_) & (g10) & (!sk[56]) & (g120)) + ((!i_8_) & (g10) & (sk[56]) & (!g120)) + ((!i_8_) & (g10) & (sk[56]) & (g120)) + ((i_8_) & (!g10) & (!sk[56]) & (g120)) + ((i_8_) & (!g10) & (sk[56]) & (!g120)) + ((i_8_) & (!g10) & (sk[56]) & (g120)) + ((i_8_) & (g10) & (!sk[56]) & (!g120)) + ((i_8_) & (g10) & (!sk[56]) & (g120)) + ((i_8_) & (g10) & (sk[56]) & (!g120)));
	assign g155 = (((!g125) & (g154) & (!sk[57]) & (!g122)) + ((!g125) & (g154) & (!sk[57]) & (g122)) + ((!g125) & (g154) & (sk[57]) & (!g122)) + ((g125) & (!g154) & (!sk[57]) & (g122)) + ((g125) & (g154) & (!sk[57]) & (!g122)) + ((g125) & (g154) & (!sk[57]) & (g122)));
	assign g156 = (((!sk[58]) & (!i_15_) & (!g34) & (!g108) & (g68) & (!g155)) + ((!sk[58]) & (!i_15_) & (!g34) & (!g108) & (g68) & (g155)) + ((!sk[58]) & (!i_15_) & (!g34) & (g108) & (!g68) & (!g155)) + ((!sk[58]) & (!i_15_) & (!g34) & (g108) & (!g68) & (g155)) + ((!sk[58]) & (!i_15_) & (!g34) & (g108) & (g68) & (!g155)) + ((!sk[58]) & (!i_15_) & (!g34) & (g108) & (g68) & (g155)) + ((!sk[58]) & (!i_15_) & (g34) & (!g108) & (!g68) & (!g155)) + ((!sk[58]) & (!i_15_) & (g34) & (!g108) & (!g68) & (g155)) + ((!sk[58]) & (!i_15_) & (g34) & (!g108) & (g68) & (!g155)) + ((!sk[58]) & (!i_15_) & (g34) & (!g108) & (g68) & (g155)) + ((!sk[58]) & (!i_15_) & (g34) & (g108) & (!g68) & (!g155)) + ((!sk[58]) & (!i_15_) & (g34) & (g108) & (!g68) & (g155)) + ((!sk[58]) & (!i_15_) & (g34) & (g108) & (g68) & (!g155)) + ((!sk[58]) & (!i_15_) & (g34) & (g108) & (g68) & (g155)) + ((!sk[58]) & (i_15_) & (!g34) & (!g108) & (g68) & (!g155)) + ((!sk[58]) & (i_15_) & (!g34) & (!g108) & (g68) & (g155)) + ((!sk[58]) & (i_15_) & (!g34) & (g108) & (!g68) & (!g155)) + ((!sk[58]) & (i_15_) & (!g34) & (g108) & (!g68) & (g155)) + ((!sk[58]) & (i_15_) & (!g34) & (g108) & (g68) & (!g155)) + ((!sk[58]) & (i_15_) & (!g34) & (g108) & (g68) & (g155)) + ((!sk[58]) & (i_15_) & (g34) & (!g108) & (!g68) & (!g155)) + ((!sk[58]) & (i_15_) & (g34) & (!g108) & (!g68) & (g155)) + ((!sk[58]) & (i_15_) & (g34) & (!g108) & (g68) & (!g155)) + ((!sk[58]) & (i_15_) & (g34) & (!g108) & (g68) & (g155)) + ((!sk[58]) & (i_15_) & (g34) & (g108) & (!g68) & (!g155)) + ((!sk[58]) & (i_15_) & (g34) & (g108) & (!g68) & (g155)) + ((!sk[58]) & (i_15_) & (g34) & (g108) & (g68) & (!g155)) + ((!sk[58]) & (i_15_) & (g34) & (g108) & (g68) & (g155)) + ((sk[58]) & (!i_15_) & (!g34) & (g108) & (!g68) & (!g155)) + ((sk[58]) & (!i_15_) & (!g34) & (g108) & (g68) & (!g155)) + ((sk[58]) & (!i_15_) & (g34) & (g108) & (!g68) & (!g155)) + ((sk[58]) & (!i_15_) & (g34) & (g108) & (g68) & (!g155)) + ((sk[58]) & (i_15_) & (!g34) & (g108) & (!g68) & (!g155)) + ((sk[58]) & (i_15_) & (!g34) & (g108) & (g68) & (!g155)) + ((sk[58]) & (i_15_) & (g34) & (!g108) & (!g68) & (!g155)) + ((sk[58]) & (i_15_) & (g34) & (g108) & (!g68) & (!g155)) + ((sk[58]) & (i_15_) & (g34) & (g108) & (g68) & (!g155)));
	assign g157 = (((!g43) & (!sk[59]) & (g72)) + ((g43) & (!sk[59]) & (g72)) + ((g43) & (sk[59]) & (g72)));
	assign g158 = (((!g157) & (!g90) & (!g78) & (sk[60]) & (!g135)) + ((!g157) & (g90) & (!g78) & (!sk[60]) & (!g135)) + ((!g157) & (g90) & (!g78) & (!sk[60]) & (g135)) + ((!g157) & (g90) & (!g78) & (sk[60]) & (!g135)) + ((!g157) & (g90) & (g78) & (!sk[60]) & (!g135)) + ((!g157) & (g90) & (g78) & (!sk[60]) & (g135)) + ((g157) & (!g90) & (!g78) & (sk[60]) & (!g135)) + ((g157) & (g90) & (!g78) & (!sk[60]) & (!g135)) + ((g157) & (g90) & (!g78) & (!sk[60]) & (g135)) + ((g157) & (g90) & (!g78) & (sk[60]) & (!g135)) + ((g157) & (g90) & (!g78) & (sk[60]) & (g135)) + ((g157) & (g90) & (g78) & (!sk[60]) & (!g135)) + ((g157) & (g90) & (g78) & (!sk[60]) & (g135)) + ((g157) & (g90) & (g78) & (sk[60]) & (!g135)) + ((g157) & (g90) & (g78) & (sk[60]) & (g135)));
	assign g159 = (((!i_8_) & (!sk[61]) & (g10) & (!g120)) + ((!i_8_) & (!sk[61]) & (g10) & (g120)) + ((!i_8_) & (sk[61]) & (!g10) & (!g120)) + ((!i_8_) & (sk[61]) & (!g10) & (g120)) + ((!i_8_) & (sk[61]) & (g10) & (!g120)) + ((i_8_) & (!sk[61]) & (!g10) & (g120)) + ((i_8_) & (!sk[61]) & (g10) & (!g120)) + ((i_8_) & (!sk[61]) & (g10) & (g120)) + ((i_8_) & (sk[61]) & (!g10) & (!g120)) + ((i_8_) & (sk[61]) & (!g10) & (g120)) + ((i_8_) & (sk[61]) & (g10) & (!g120)) + ((i_8_) & (sk[61]) & (g10) & (g120)));
	assign g160 = (((!g87) & (!g98) & (sk[62]) & (!g144) & (!g159)) + ((!g87) & (!g98) & (sk[62]) & (g144) & (!g159)) + ((!g87) & (g98) & (!sk[62]) & (!g144) & (!g159)) + ((!g87) & (g98) & (!sk[62]) & (!g144) & (g159)) + ((!g87) & (g98) & (!sk[62]) & (g144) & (!g159)) + ((!g87) & (g98) & (!sk[62]) & (g144) & (g159)) + ((!g87) & (g98) & (sk[62]) & (!g144) & (!g159)) + ((!g87) & (g98) & (sk[62]) & (g144) & (!g159)) + ((!g87) & (g98) & (sk[62]) & (g144) & (g159)) + ((g87) & (g98) & (!sk[62]) & (!g144) & (!g159)) + ((g87) & (g98) & (!sk[62]) & (!g144) & (g159)) + ((g87) & (g98) & (!sk[62]) & (g144) & (!g159)) + ((g87) & (g98) & (!sk[62]) & (g144) & (g159)) + ((g87) & (g98) & (sk[62]) & (g144) & (!g159)) + ((g87) & (g98) & (sk[62]) & (g144) & (g159)));
	assign g161 = (((!g49) & (!sk[63]) & (g72)) + ((g49) & (!sk[63]) & (g72)) + ((g49) & (sk[63]) & (g72)));
	assign g162 = (((!i_8_) & (!g73) & (!g108) & (!g109) & (!g154) & (!g122)) + ((!i_8_) & (!g73) & (!g108) & (!g109) & (!g154) & (g122)) + ((!i_8_) & (!g73) & (!g108) & (!g109) & (g154) & (!g122)) + ((!i_8_) & (!g73) & (!g108) & (!g109) & (g154) & (g122)) + ((!i_8_) & (!g73) & (!g108) & (g109) & (g154) & (!g122)) + ((!i_8_) & (!g73) & (g108) & (!g109) & (!g154) & (!g122)) + ((!i_8_) & (!g73) & (g108) & (!g109) & (!g154) & (g122)) + ((!i_8_) & (!g73) & (g108) & (!g109) & (g154) & (!g122)) + ((!i_8_) & (!g73) & (g108) & (!g109) & (g154) & (g122)) + ((!i_8_) & (!g73) & (g108) & (g109) & (g154) & (!g122)) + ((!i_8_) & (g73) & (!g108) & (!g109) & (!g154) & (!g122)) + ((!i_8_) & (g73) & (!g108) & (!g109) & (!g154) & (g122)) + ((!i_8_) & (g73) & (!g108) & (!g109) & (g154) & (!g122)) + ((!i_8_) & (g73) & (!g108) & (!g109) & (g154) & (g122)) + ((!i_8_) & (g73) & (g108) & (!g109) & (!g154) & (!g122)) + ((!i_8_) & (g73) & (g108) & (!g109) & (!g154) & (g122)) + ((!i_8_) & (g73) & (g108) & (!g109) & (g154) & (!g122)) + ((!i_8_) & (g73) & (g108) & (!g109) & (g154) & (g122)) + ((i_8_) & (!g73) & (!g108) & (!g109) & (!g154) & (!g122)) + ((i_8_) & (!g73) & (!g108) & (!g109) & (!g154) & (g122)) + ((i_8_) & (!g73) & (!g108) & (!g109) & (g154) & (!g122)) + ((i_8_) & (!g73) & (!g108) & (!g109) & (g154) & (g122)) + ((i_8_) & (!g73) & (!g108) & (g109) & (g154) & (!g122)) + ((i_8_) & (!g73) & (g108) & (!g109) & (!g154) & (!g122)) + ((i_8_) & (!g73) & (g108) & (!g109) & (!g154) & (g122)) + ((i_8_) & (!g73) & (g108) & (!g109) & (g154) & (!g122)) + ((i_8_) & (!g73) & (g108) & (!g109) & (g154) & (g122)) + ((i_8_) & (!g73) & (g108) & (g109) & (g154) & (!g122)) + ((i_8_) & (g73) & (!g108) & (!g109) & (!g154) & (!g122)) + ((i_8_) & (g73) & (!g108) & (!g109) & (!g154) & (g122)) + ((i_8_) & (g73) & (!g108) & (!g109) & (g154) & (!g122)) + ((i_8_) & (g73) & (!g108) & (!g109) & (g154) & (g122)));
	assign g163 = (((!g109) & (!g161) & (!g87) & (!g125) & (!g78) & (g162)) + ((!g109) & (!g161) & (!g87) & (!g125) & (g78) & (g162)) + ((!g109) & (!g161) & (g87) & (!g125) & (!g78) & (g162)) + ((!g109) & (!g161) & (g87) & (!g125) & (g78) & (g162)) + ((!g109) & (!g161) & (g87) & (g125) & (g78) & (g162)) + ((!g109) & (g161) & (!g87) & (!g125) & (!g78) & (g162)) + ((!g109) & (g161) & (!g87) & (!g125) & (g78) & (g162)) + ((!g109) & (g161) & (g87) & (!g125) & (!g78) & (g162)) + ((!g109) & (g161) & (g87) & (!g125) & (g78) & (g162)) + ((!g109) & (g161) & (g87) & (g125) & (g78) & (g162)) + ((g109) & (!g161) & (!g87) & (!g125) & (!g78) & (g162)) + ((g109) & (!g161) & (!g87) & (!g125) & (g78) & (g162)) + ((g109) & (!g161) & (g87) & (!g125) & (!g78) & (g162)) + ((g109) & (!g161) & (g87) & (!g125) & (g78) & (g162)));
	assign g164 = (((!g30) & (!sk[66]) & (g120)) + ((g30) & (!sk[66]) & (g120)) + ((g30) & (sk[66]) & (g120)));
	assign g165 = (((!g42) & (!sk[67]) & (g118)) + ((g42) & (!sk[67]) & (g118)) + ((g42) & (sk[67]) & (g118)));
	assign g166 = (((!i_4_) & (!i_3_) & (sk[68]) & (i_5_) & (g71)) + ((!i_4_) & (i_3_) & (!sk[68]) & (!i_5_) & (!g71)) + ((!i_4_) & (i_3_) & (!sk[68]) & (!i_5_) & (g71)) + ((!i_4_) & (i_3_) & (!sk[68]) & (i_5_) & (!g71)) + ((!i_4_) & (i_3_) & (!sk[68]) & (i_5_) & (g71)) + ((i_4_) & (!i_3_) & (sk[68]) & (!i_5_) & (g71)) + ((i_4_) & (i_3_) & (!sk[68]) & (!i_5_) & (!g71)) + ((i_4_) & (i_3_) & (!sk[68]) & (!i_5_) & (g71)) + ((i_4_) & (i_3_) & (!sk[68]) & (i_5_) & (!g71)) + ((i_4_) & (i_3_) & (!sk[68]) & (i_5_) & (g71)));
	assign g167 = (((!g101) & (!sk[69]) & (g166)) + ((g101) & (!sk[69]) & (g166)) + ((g101) & (sk[69]) & (g166)));
	assign g168 = (((!g45) & (!sk[70]) & (g72)) + ((g45) & (!sk[70]) & (g72)) + ((g45) & (sk[70]) & (g72)));
	assign g169 = (((!i_8_) & (i_6_) & (!sk[71]) & (!g120) & (!g77)) + ((!i_8_) & (i_6_) & (!sk[71]) & (!g120) & (g77)) + ((!i_8_) & (i_6_) & (!sk[71]) & (g120) & (!g77)) + ((!i_8_) & (i_6_) & (!sk[71]) & (g120) & (g77)) + ((i_8_) & (i_6_) & (!sk[71]) & (!g120) & (!g77)) + ((i_8_) & (i_6_) & (!sk[71]) & (!g120) & (g77)) + ((i_8_) & (i_6_) & (!sk[71]) & (g120) & (!g77)) + ((i_8_) & (i_6_) & (!sk[71]) & (g120) & (g77)) + ((i_8_) & (i_6_) & (sk[71]) & (g120) & (g77)));
	assign g170 = (((!g125) & (!g167) & (!g97) & (!g70) & (!g168) & (!g169)) + ((!g125) & (!g167) & (!g97) & (!g70) & (g168) & (!g169)) + ((!g125) & (!g167) & (!g97) & (g70) & (!g168) & (!g169)) + ((!g125) & (!g167) & (g97) & (!g70) & (!g168) & (!g169)) + ((!g125) & (!g167) & (g97) & (!g70) & (g168) & (!g169)) + ((!g125) & (!g167) & (g97) & (g70) & (!g168) & (!g169)) + ((!g125) & (g167) & (g97) & (!g70) & (!g168) & (!g169)) + ((!g125) & (g167) & (g97) & (!g70) & (g168) & (!g169)) + ((!g125) & (g167) & (g97) & (g70) & (!g168) & (!g169)) + ((g125) & (!g167) & (!g97) & (!g70) & (!g168) & (!g169)) + ((g125) & (!g167) & (!g97) & (!g70) & (g168) & (!g169)) + ((g125) & (!g167) & (g97) & (!g70) & (!g168) & (!g169)) + ((g125) & (!g167) & (g97) & (!g70) & (g168) & (!g169)) + ((g125) & (g167) & (g97) & (!g70) & (!g168) & (!g169)) + ((g125) & (g167) & (g97) & (!g70) & (g168) & (!g169)));
	assign g171 = (((!g87) & (!g127) & (!g164) & (!g102) & (!g165) & (g170)) + ((!g87) & (!g127) & (!g164) & (g102) & (!g165) & (g170)) + ((!g87) & (!g127) & (g164) & (!g102) & (!g165) & (g170)) + ((!g87) & (!g127) & (g164) & (g102) & (!g165) & (g170)) + ((!g87) & (g127) & (!g164) & (!g102) & (!g165) & (g170)) + ((g87) & (!g127) & (!g164) & (!g102) & (!g165) & (g170)) + ((g87) & (!g127) & (!g164) & (!g102) & (g165) & (g170)) + ((g87) & (!g127) & (!g164) & (g102) & (!g165) & (g170)) + ((g87) & (!g127) & (!g164) & (g102) & (g165) & (g170)) + ((g87) & (!g127) & (g164) & (!g102) & (!g165) & (g170)) + ((g87) & (!g127) & (g164) & (!g102) & (g165) & (g170)) + ((g87) & (!g127) & (g164) & (g102) & (!g165) & (g170)) + ((g87) & (!g127) & (g164) & (g102) & (g165) & (g170)) + ((g87) & (g127) & (!g164) & (!g102) & (!g165) & (g170)) + ((g87) & (g127) & (!g164) & (!g102) & (g165) & (g170)));
	assign g172 = (((!g156) & (!sk[74]) & (!g158) & (!g160) & (g163) & (!g171)) + ((!g156) & (!sk[74]) & (!g158) & (!g160) & (g163) & (g171)) + ((!g156) & (!sk[74]) & (!g158) & (g160) & (!g163) & (!g171)) + ((!g156) & (!sk[74]) & (!g158) & (g160) & (!g163) & (g171)) + ((!g156) & (!sk[74]) & (!g158) & (g160) & (g163) & (!g171)) + ((!g156) & (!sk[74]) & (!g158) & (g160) & (g163) & (g171)) + ((!g156) & (!sk[74]) & (g158) & (!g160) & (!g163) & (!g171)) + ((!g156) & (!sk[74]) & (g158) & (!g160) & (!g163) & (g171)) + ((!g156) & (!sk[74]) & (g158) & (!g160) & (g163) & (!g171)) + ((!g156) & (!sk[74]) & (g158) & (!g160) & (g163) & (g171)) + ((!g156) & (!sk[74]) & (g158) & (g160) & (!g163) & (!g171)) + ((!g156) & (!sk[74]) & (g158) & (g160) & (!g163) & (g171)) + ((!g156) & (!sk[74]) & (g158) & (g160) & (g163) & (!g171)) + ((!g156) & (!sk[74]) & (g158) & (g160) & (g163) & (g171)) + ((!g156) & (sk[74]) & (!g158) & (!g160) & (g163) & (g171)) + ((g156) & (!sk[74]) & (!g158) & (!g160) & (g163) & (!g171)) + ((g156) & (!sk[74]) & (!g158) & (!g160) & (g163) & (g171)) + ((g156) & (!sk[74]) & (!g158) & (g160) & (!g163) & (!g171)) + ((g156) & (!sk[74]) & (!g158) & (g160) & (!g163) & (g171)) + ((g156) & (!sk[74]) & (!g158) & (g160) & (g163) & (!g171)) + ((g156) & (!sk[74]) & (!g158) & (g160) & (g163) & (g171)) + ((g156) & (!sk[74]) & (g158) & (!g160) & (!g163) & (!g171)) + ((g156) & (!sk[74]) & (g158) & (!g160) & (!g163) & (g171)) + ((g156) & (!sk[74]) & (g158) & (!g160) & (g163) & (!g171)) + ((g156) & (!sk[74]) & (g158) & (!g160) & (g163) & (g171)) + ((g156) & (!sk[74]) & (g158) & (g160) & (!g163) & (!g171)) + ((g156) & (!sk[74]) & (g158) & (g160) & (!g163) & (g171)) + ((g156) & (!sk[74]) & (g158) & (g160) & (g163) & (!g171)) + ((g156) & (!sk[74]) & (g158) & (g160) & (g163) & (g171)));
	assign g173 = (((g100) & (g117) & (g129) & (g132) & (g153) & (g172)));
	assign g174 = (((!i_12_) & (!sk[76]) & (i_13_) & (!i_14_)) + ((!i_12_) & (!sk[76]) & (i_13_) & (i_14_)) + ((!i_12_) & (sk[76]) & (!i_13_) & (!i_14_)) + ((!i_12_) & (sk[76]) & (!i_13_) & (i_14_)) + ((!i_12_) & (sk[76]) & (i_13_) & (!i_14_)) + ((!i_12_) & (sk[76]) & (i_13_) & (i_14_)) + ((i_12_) & (!sk[76]) & (!i_13_) & (i_14_)) + ((i_12_) & (!sk[76]) & (i_13_) & (!i_14_)) + ((i_12_) & (!sk[76]) & (i_13_) & (i_14_)) + ((i_12_) & (sk[76]) & (!i_13_) & (!i_14_)) + ((i_12_) & (sk[76]) & (!i_13_) & (i_14_)) + ((i_12_) & (sk[76]) & (i_13_) & (!i_14_)));
	assign g175 = (((!g20) & (!sk[77]) & (g174)) + ((g20) & (!sk[77]) & (g174)) + ((g20) & (sk[77]) & (!g174)));
	assign g176 = (((!i_12_) & (!sk[78]) & (i_13_) & (!i_14_)) + ((!i_12_) & (!sk[78]) & (i_13_) & (i_14_)) + ((!i_12_) & (sk[78]) & (!i_13_) & (!i_14_)) + ((!i_12_) & (sk[78]) & (!i_13_) & (i_14_)) + ((!i_12_) & (sk[78]) & (i_13_) & (!i_14_)) + ((!i_12_) & (sk[78]) & (i_13_) & (i_14_)) + ((i_12_) & (!sk[78]) & (!i_13_) & (i_14_)) + ((i_12_) & (!sk[78]) & (i_13_) & (!i_14_)) + ((i_12_) & (!sk[78]) & (i_13_) & (i_14_)) + ((i_12_) & (sk[78]) & (!i_13_) & (!i_14_)) + ((i_12_) & (sk[78]) & (i_13_) & (!i_14_)) + ((i_12_) & (sk[78]) & (i_13_) & (i_14_)));
	assign g177 = (((!g22) & (!sk[79]) & (g176)) + ((!g22) & (sk[79]) & (!g176)) + ((g22) & (!sk[79]) & (g176)));
	assign g178 = (((!sk[80]) & (!g75) & (g175) & (!g177)) + ((!sk[80]) & (!g75) & (g175) & (g177)) + ((!sk[80]) & (g75) & (!g175) & (g177)) + ((!sk[80]) & (g75) & (g175) & (!g177)) + ((!sk[80]) & (g75) & (g175) & (g177)) + ((sk[80]) & (!g75) & (!g175) & (g177)) + ((sk[80]) & (!g75) & (g175) & (!g177)) + ((sk[80]) & (!g75) & (g175) & (g177)));
	assign g179 = (((!g17) & (!sk[81]) & (g176)) + ((g17) & (!sk[81]) & (g176)) + ((g17) & (sk[81]) & (!g176)));
	assign g180 = (((!sk[82]) & (!g27) & (g174)) + ((!sk[82]) & (g27) & (g174)) + ((sk[82]) & (g27) & (!g174)));
	assign g181 = (((!g75) & (!g179) & (sk[83]) & (g180)) + ((!g75) & (g179) & (!sk[83]) & (!g180)) + ((!g75) & (g179) & (!sk[83]) & (g180)) + ((!g75) & (g179) & (sk[83]) & (!g180)) + ((!g75) & (g179) & (sk[83]) & (g180)) + ((g75) & (!g179) & (!sk[83]) & (g180)) + ((g75) & (g179) & (!sk[83]) & (!g180)) + ((g75) & (g179) & (!sk[83]) & (g180)));
	assign g182 = (((!sk[84]) & (!g81) & (g176)) + ((!sk[84]) & (g81) & (g176)) + ((sk[84]) & (g81) & (!g176)));
	assign g183 = (((!sk[85]) & (!g83) & (g174)) + ((!sk[85]) & (g83) & (g174)) + ((sk[85]) & (g83) & (!g174)));
	assign g184 = (((!g74) & (!sk[86]) & (g182) & (!g183)) + ((!g74) & (!sk[86]) & (g182) & (g183)) + ((g74) & (!sk[86]) & (!g182) & (g183)) + ((g74) & (!sk[86]) & (g182) & (!g183)) + ((g74) & (!sk[86]) & (g182) & (g183)) + ((g74) & (sk[86]) & (!g182) & (g183)) + ((g74) & (sk[86]) & (g182) & (!g183)) + ((g74) & (sk[86]) & (g182) & (g183)));
	assign g185 = (((!sk[87]) & (!g91) & (g176)) + ((!sk[87]) & (g91) & (g176)) + ((sk[87]) & (!g91) & (!g176)));
	assign g186 = (((!g36) & (!sk[88]) & (g176)) + ((g36) & (!sk[88]) & (g176)) + ((g36) & (sk[88]) & (!g176)));
	assign g187 = (((!g88) & (!sk[89]) & (g176)) + ((g88) & (!sk[89]) & (g176)) + ((g88) & (sk[89]) & (!g176)));
	assign g188 = (((!g3) & (!sk[90]) & (g174)) + ((g3) & (!sk[90]) & (g174)) + ((g3) & (sk[90]) & (!g174)));
	assign g189 = (((!i_8_) & (g73) & (!g179) & (!g188) & (!g175) & (g180)) + ((!i_8_) & (g73) & (!g179) & (!g188) & (g175) & (!g180)) + ((!i_8_) & (g73) & (!g179) & (!g188) & (g175) & (g180)) + ((!i_8_) & (g73) & (!g179) & (g188) & (!g175) & (!g180)) + ((!i_8_) & (g73) & (!g179) & (g188) & (!g175) & (g180)) + ((!i_8_) & (g73) & (!g179) & (g188) & (g175) & (!g180)) + ((!i_8_) & (g73) & (!g179) & (g188) & (g175) & (g180)) + ((!i_8_) & (g73) & (g179) & (!g188) & (!g175) & (!g180)) + ((!i_8_) & (g73) & (g179) & (!g188) & (!g175) & (g180)) + ((!i_8_) & (g73) & (g179) & (!g188) & (g175) & (!g180)) + ((!i_8_) & (g73) & (g179) & (!g188) & (g175) & (g180)) + ((!i_8_) & (g73) & (g179) & (g188) & (!g175) & (!g180)) + ((!i_8_) & (g73) & (g179) & (g188) & (!g175) & (g180)) + ((!i_8_) & (g73) & (g179) & (g188) & (g175) & (!g180)) + ((!i_8_) & (g73) & (g179) & (g188) & (g175) & (g180)));
	assign g190 = (((!g75) & (!g185) & (!g186) & (!sk[92]) & (g187) & (!g189)) + ((!g75) & (!g185) & (!g186) & (!sk[92]) & (g187) & (g189)) + ((!g75) & (!g185) & (!g186) & (sk[92]) & (!g187) & (!g189)) + ((!g75) & (!g185) & (g186) & (!sk[92]) & (!g187) & (!g189)) + ((!g75) & (!g185) & (g186) & (!sk[92]) & (!g187) & (g189)) + ((!g75) & (!g185) & (g186) & (!sk[92]) & (g187) & (!g189)) + ((!g75) & (!g185) & (g186) & (!sk[92]) & (g187) & (g189)) + ((!g75) & (g185) & (!g186) & (!sk[92]) & (!g187) & (!g189)) + ((!g75) & (g185) & (!g186) & (!sk[92]) & (!g187) & (g189)) + ((!g75) & (g185) & (!g186) & (!sk[92]) & (g187) & (!g189)) + ((!g75) & (g185) & (!g186) & (!sk[92]) & (g187) & (g189)) + ((!g75) & (g185) & (g186) & (!sk[92]) & (!g187) & (!g189)) + ((!g75) & (g185) & (g186) & (!sk[92]) & (!g187) & (g189)) + ((!g75) & (g185) & (g186) & (!sk[92]) & (g187) & (!g189)) + ((!g75) & (g185) & (g186) & (!sk[92]) & (g187) & (g189)) + ((g75) & (!g185) & (!g186) & (!sk[92]) & (g187) & (!g189)) + ((g75) & (!g185) & (!g186) & (!sk[92]) & (g187) & (g189)) + ((g75) & (!g185) & (!g186) & (sk[92]) & (!g187) & (!g189)) + ((g75) & (!g185) & (!g186) & (sk[92]) & (g187) & (!g189)) + ((g75) & (!g185) & (g186) & (!sk[92]) & (!g187) & (!g189)) + ((g75) & (!g185) & (g186) & (!sk[92]) & (!g187) & (g189)) + ((g75) & (!g185) & (g186) & (!sk[92]) & (g187) & (!g189)) + ((g75) & (!g185) & (g186) & (!sk[92]) & (g187) & (g189)) + ((g75) & (!g185) & (g186) & (sk[92]) & (!g187) & (!g189)) + ((g75) & (!g185) & (g186) & (sk[92]) & (g187) & (!g189)) + ((g75) & (g185) & (!g186) & (!sk[92]) & (!g187) & (!g189)) + ((g75) & (g185) & (!g186) & (!sk[92]) & (!g187) & (g189)) + ((g75) & (g185) & (!g186) & (!sk[92]) & (g187) & (!g189)) + ((g75) & (g185) & (!g186) & (!sk[92]) & (g187) & (g189)) + ((g75) & (g185) & (!g186) & (sk[92]) & (!g187) & (!g189)) + ((g75) & (g185) & (!g186) & (sk[92]) & (g187) & (!g189)) + ((g75) & (g185) & (g186) & (!sk[92]) & (!g187) & (!g189)) + ((g75) & (g185) & (g186) & (!sk[92]) & (!g187) & (g189)) + ((g75) & (g185) & (g186) & (!sk[92]) & (g187) & (!g189)) + ((g75) & (g185) & (g186) & (!sk[92]) & (g187) & (g189)) + ((g75) & (g185) & (g186) & (sk[92]) & (!g187) & (!g189)) + ((g75) & (g185) & (g186) & (sk[92]) & (g187) & (!g189)));
	assign g191 = (((!g86) & (!sk[93]) & (g174)) + ((g86) & (!sk[93]) & (g174)) + ((g86) & (sk[93]) & (!g174)));
	assign g192 = (((!g35) & (!sk[94]) & (g174)) + ((g35) & (!sk[94]) & (g174)) + ((g35) & (sk[94]) & (!g174)));
	assign g193 = (((!g74) & (!g191) & (!g186) & (!sk[95]) & (g187) & (!g192)) + ((!g74) & (!g191) & (!g186) & (!sk[95]) & (g187) & (g192)) + ((!g74) & (!g191) & (g186) & (!sk[95]) & (!g187) & (!g192)) + ((!g74) & (!g191) & (g186) & (!sk[95]) & (!g187) & (g192)) + ((!g74) & (!g191) & (g186) & (!sk[95]) & (g187) & (!g192)) + ((!g74) & (!g191) & (g186) & (!sk[95]) & (g187) & (g192)) + ((!g74) & (g191) & (!g186) & (!sk[95]) & (!g187) & (!g192)) + ((!g74) & (g191) & (!g186) & (!sk[95]) & (!g187) & (g192)) + ((!g74) & (g191) & (!g186) & (!sk[95]) & (g187) & (!g192)) + ((!g74) & (g191) & (!g186) & (!sk[95]) & (g187) & (g192)) + ((!g74) & (g191) & (g186) & (!sk[95]) & (!g187) & (!g192)) + ((!g74) & (g191) & (g186) & (!sk[95]) & (!g187) & (g192)) + ((!g74) & (g191) & (g186) & (!sk[95]) & (g187) & (!g192)) + ((!g74) & (g191) & (g186) & (!sk[95]) & (g187) & (g192)) + ((g74) & (!g191) & (!g186) & (!sk[95]) & (g187) & (!g192)) + ((g74) & (!g191) & (!g186) & (!sk[95]) & (g187) & (g192)) + ((g74) & (!g191) & (!g186) & (sk[95]) & (!g187) & (g192)) + ((g74) & (!g191) & (!g186) & (sk[95]) & (g187) & (!g192)) + ((g74) & (!g191) & (!g186) & (sk[95]) & (g187) & (g192)) + ((g74) & (!g191) & (g186) & (!sk[95]) & (!g187) & (!g192)) + ((g74) & (!g191) & (g186) & (!sk[95]) & (!g187) & (g192)) + ((g74) & (!g191) & (g186) & (!sk[95]) & (g187) & (!g192)) + ((g74) & (!g191) & (g186) & (!sk[95]) & (g187) & (g192)) + ((g74) & (!g191) & (g186) & (sk[95]) & (!g187) & (!g192)) + ((g74) & (!g191) & (g186) & (sk[95]) & (!g187) & (g192)) + ((g74) & (!g191) & (g186) & (sk[95]) & (g187) & (!g192)) + ((g74) & (!g191) & (g186) & (sk[95]) & (g187) & (g192)) + ((g74) & (g191) & (!g186) & (!sk[95]) & (!g187) & (!g192)) + ((g74) & (g191) & (!g186) & (!sk[95]) & (!g187) & (g192)) + ((g74) & (g191) & (!g186) & (!sk[95]) & (g187) & (!g192)) + ((g74) & (g191) & (!g186) & (!sk[95]) & (g187) & (g192)) + ((g74) & (g191) & (!g186) & (sk[95]) & (!g187) & (!g192)) + ((g74) & (g191) & (!g186) & (sk[95]) & (!g187) & (g192)) + ((g74) & (g191) & (!g186) & (sk[95]) & (g187) & (!g192)) + ((g74) & (g191) & (!g186) & (sk[95]) & (g187) & (g192)) + ((g74) & (g191) & (g186) & (!sk[95]) & (!g187) & (!g192)) + ((g74) & (g191) & (g186) & (!sk[95]) & (!g187) & (g192)) + ((g74) & (g191) & (g186) & (!sk[95]) & (g187) & (!g192)) + ((g74) & (g191) & (g186) & (!sk[95]) & (g187) & (g192)) + ((g74) & (g191) & (g186) & (sk[95]) & (!g187) & (!g192)) + ((g74) & (g191) & (g186) & (sk[95]) & (!g187) & (g192)) + ((g74) & (g191) & (g186) & (sk[95]) & (g187) & (!g192)) + ((g74) & (g191) & (g186) & (sk[95]) & (g187) & (g192)));
	assign g194 = (((!g69) & (!sk[96]) & (g176)) + ((g69) & (!sk[96]) & (g176)) + ((g69) & (sk[96]) & (!g176)));
	assign g195 = (((!g75) & (!sk[97]) & (!g194) & (!g188) & (g182) & (!g183)) + ((!g75) & (!sk[97]) & (!g194) & (!g188) & (g182) & (g183)) + ((!g75) & (!sk[97]) & (!g194) & (g188) & (!g182) & (!g183)) + ((!g75) & (!sk[97]) & (!g194) & (g188) & (!g182) & (g183)) + ((!g75) & (!sk[97]) & (!g194) & (g188) & (g182) & (!g183)) + ((!g75) & (!sk[97]) & (!g194) & (g188) & (g182) & (g183)) + ((!g75) & (!sk[97]) & (g194) & (!g188) & (!g182) & (!g183)) + ((!g75) & (!sk[97]) & (g194) & (!g188) & (!g182) & (g183)) + ((!g75) & (!sk[97]) & (g194) & (!g188) & (g182) & (!g183)) + ((!g75) & (!sk[97]) & (g194) & (!g188) & (g182) & (g183)) + ((!g75) & (!sk[97]) & (g194) & (g188) & (!g182) & (!g183)) + ((!g75) & (!sk[97]) & (g194) & (g188) & (!g182) & (g183)) + ((!g75) & (!sk[97]) & (g194) & (g188) & (g182) & (!g183)) + ((!g75) & (!sk[97]) & (g194) & (g188) & (g182) & (g183)) + ((!g75) & (sk[97]) & (!g194) & (!g188) & (!g182) & (g183)) + ((!g75) & (sk[97]) & (!g194) & (!g188) & (g182) & (!g183)) + ((!g75) & (sk[97]) & (!g194) & (!g188) & (g182) & (g183)) + ((!g75) & (sk[97]) & (!g194) & (g188) & (!g182) & (!g183)) + ((!g75) & (sk[97]) & (!g194) & (g188) & (!g182) & (g183)) + ((!g75) & (sk[97]) & (!g194) & (g188) & (g182) & (!g183)) + ((!g75) & (sk[97]) & (!g194) & (g188) & (g182) & (g183)) + ((!g75) & (sk[97]) & (g194) & (!g188) & (!g182) & (!g183)) + ((!g75) & (sk[97]) & (g194) & (!g188) & (!g182) & (g183)) + ((!g75) & (sk[97]) & (g194) & (!g188) & (g182) & (!g183)) + ((!g75) & (sk[97]) & (g194) & (!g188) & (g182) & (g183)) + ((!g75) & (sk[97]) & (g194) & (g188) & (!g182) & (!g183)) + ((!g75) & (sk[97]) & (g194) & (g188) & (!g182) & (g183)) + ((!g75) & (sk[97]) & (g194) & (g188) & (g182) & (!g183)) + ((!g75) & (sk[97]) & (g194) & (g188) & (g182) & (g183)) + ((g75) & (!sk[97]) & (!g194) & (!g188) & (g182) & (!g183)) + ((g75) & (!sk[97]) & (!g194) & (!g188) & (g182) & (g183)) + ((g75) & (!sk[97]) & (!g194) & (g188) & (!g182) & (!g183)) + ((g75) & (!sk[97]) & (!g194) & (g188) & (!g182) & (g183)) + ((g75) & (!sk[97]) & (!g194) & (g188) & (g182) & (!g183)) + ((g75) & (!sk[97]) & (!g194) & (g188) & (g182) & (g183)) + ((g75) & (!sk[97]) & (g194) & (!g188) & (!g182) & (!g183)) + ((g75) & (!sk[97]) & (g194) & (!g188) & (!g182) & (g183)) + ((g75) & (!sk[97]) & (g194) & (!g188) & (g182) & (!g183)) + ((g75) & (!sk[97]) & (g194) & (!g188) & (g182) & (g183)) + ((g75) & (!sk[97]) & (g194) & (g188) & (!g182) & (!g183)) + ((g75) & (!sk[97]) & (g194) & (g188) & (!g182) & (g183)) + ((g75) & (!sk[97]) & (g194) & (g188) & (g182) & (!g183)) + ((g75) & (!sk[97]) & (g194) & (g188) & (g182) & (g183)));
	assign g196 = (((!g178) & (!g181) & (!g184) & (g190) & (!g193) & (!g195)));
	assign g197 = (((!g113) & (!sk[99]) & (g176)) + ((!g113) & (sk[99]) & (!g176)) + ((g113) & (!sk[99]) & (g176)));
	assign g198 = (((!g123) & (!sk[100]) & (g194) & (!g188)) + ((!g123) & (!sk[100]) & (g194) & (g188)) + ((!g123) & (sk[100]) & (!g194) & (g188)) + ((!g123) & (sk[100]) & (g194) & (!g188)) + ((!g123) & (sk[100]) & (g194) & (g188)) + ((g123) & (!sk[100]) & (!g194) & (g188)) + ((g123) & (!sk[100]) & (g194) & (!g188)) + ((g123) & (!sk[100]) & (g194) & (g188)));
	assign g199 = (((!g105) & (!g119) & (sk[101]) & (g188)) + ((!g105) & (g119) & (!sk[101]) & (!g188)) + ((!g105) & (g119) & (!sk[101]) & (g188)) + ((!g105) & (g119) & (sk[101]) & (g188)) + ((g105) & (!g119) & (!sk[101]) & (g188)) + ((g105) & (g119) & (!sk[101]) & (!g188)) + ((g105) & (g119) & (!sk[101]) & (g188)) + ((g105) & (g119) & (sk[101]) & (g188)));
	assign g200 = (((!sk[102]) & (!g126) & (g174)) + ((!sk[102]) & (g126) & (g174)) + ((sk[102]) & (!g126) & (!g174)));
	assign g201 = (((!g125) & (!g122) & (!g123) & (!g197) & (sk[103]) & (!g200)) + ((!g125) & (!g122) & (!g123) & (!g197) & (sk[103]) & (g200)) + ((!g125) & (!g122) & (!g123) & (g197) & (!sk[103]) & (!g200)) + ((!g125) & (!g122) & (!g123) & (g197) & (!sk[103]) & (g200)) + ((!g125) & (!g122) & (g123) & (!g197) & (!sk[103]) & (!g200)) + ((!g125) & (!g122) & (g123) & (!g197) & (!sk[103]) & (g200)) + ((!g125) & (!g122) & (g123) & (!g197) & (sk[103]) & (!g200)) + ((!g125) & (!g122) & (g123) & (!g197) & (sk[103]) & (g200)) + ((!g125) & (!g122) & (g123) & (g197) & (!sk[103]) & (!g200)) + ((!g125) & (!g122) & (g123) & (g197) & (!sk[103]) & (g200)) + ((!g125) & (!g122) & (g123) & (g197) & (sk[103]) & (!g200)) + ((!g125) & (!g122) & (g123) & (g197) & (sk[103]) & (g200)) + ((!g125) & (g122) & (!g123) & (!g197) & (!sk[103]) & (!g200)) + ((!g125) & (g122) & (!g123) & (!g197) & (!sk[103]) & (g200)) + ((!g125) & (g122) & (!g123) & (!g197) & (sk[103]) & (!g200)) + ((!g125) & (g122) & (!g123) & (g197) & (!sk[103]) & (!g200)) + ((!g125) & (g122) & (!g123) & (g197) & (!sk[103]) & (g200)) + ((!g125) & (g122) & (g123) & (!g197) & (!sk[103]) & (!g200)) + ((!g125) & (g122) & (g123) & (!g197) & (!sk[103]) & (g200)) + ((!g125) & (g122) & (g123) & (!g197) & (sk[103]) & (!g200)) + ((!g125) & (g122) & (g123) & (g197) & (!sk[103]) & (!g200)) + ((!g125) & (g122) & (g123) & (g197) & (!sk[103]) & (g200)) + ((g125) & (!g122) & (!g123) & (!g197) & (sk[103]) & (!g200)) + ((g125) & (!g122) & (!g123) & (g197) & (!sk[103]) & (!g200)) + ((g125) & (!g122) & (!g123) & (g197) & (!sk[103]) & (g200)) + ((g125) & (!g122) & (g123) & (!g197) & (!sk[103]) & (!g200)) + ((g125) & (!g122) & (g123) & (!g197) & (!sk[103]) & (g200)) + ((g125) & (!g122) & (g123) & (!g197) & (sk[103]) & (!g200)) + ((g125) & (!g122) & (g123) & (g197) & (!sk[103]) & (!g200)) + ((g125) & (!g122) & (g123) & (g197) & (!sk[103]) & (g200)) + ((g125) & (g122) & (!g123) & (!g197) & (!sk[103]) & (!g200)) + ((g125) & (g122) & (!g123) & (!g197) & (!sk[103]) & (g200)) + ((g125) & (g122) & (!g123) & (!g197) & (sk[103]) & (!g200)) + ((g125) & (g122) & (!g123) & (g197) & (!sk[103]) & (!g200)) + ((g125) & (g122) & (!g123) & (g197) & (!sk[103]) & (g200)) + ((g125) & (g122) & (g123) & (!g197) & (!sk[103]) & (!g200)) + ((g125) & (g122) & (g123) & (!g197) & (!sk[103]) & (g200)) + ((g125) & (g122) & (g123) & (!g197) & (sk[103]) & (!g200)) + ((g125) & (g122) & (g123) & (g197) & (!sk[103]) & (!g200)) + ((g125) & (g122) & (g123) & (g197) & (!sk[103]) & (g200)));
	assign g202 = (((!g121) & (!g194) & (!g198) & (!sk[104]) & (g199) & (!g201)) + ((!g121) & (!g194) & (!g198) & (!sk[104]) & (g199) & (g201)) + ((!g121) & (!g194) & (!g198) & (sk[104]) & (!g199) & (g201)) + ((!g121) & (!g194) & (g198) & (!sk[104]) & (!g199) & (!g201)) + ((!g121) & (!g194) & (g198) & (!sk[104]) & (!g199) & (g201)) + ((!g121) & (!g194) & (g198) & (!sk[104]) & (g199) & (!g201)) + ((!g121) & (!g194) & (g198) & (!sk[104]) & (g199) & (g201)) + ((!g121) & (g194) & (!g198) & (!sk[104]) & (!g199) & (!g201)) + ((!g121) & (g194) & (!g198) & (!sk[104]) & (!g199) & (g201)) + ((!g121) & (g194) & (!g198) & (!sk[104]) & (g199) & (!g201)) + ((!g121) & (g194) & (!g198) & (!sk[104]) & (g199) & (g201)) + ((!g121) & (g194) & (!g198) & (sk[104]) & (!g199) & (g201)) + ((!g121) & (g194) & (g198) & (!sk[104]) & (!g199) & (!g201)) + ((!g121) & (g194) & (g198) & (!sk[104]) & (!g199) & (g201)) + ((!g121) & (g194) & (g198) & (!sk[104]) & (g199) & (!g201)) + ((!g121) & (g194) & (g198) & (!sk[104]) & (g199) & (g201)) + ((g121) & (!g194) & (!g198) & (!sk[104]) & (g199) & (!g201)) + ((g121) & (!g194) & (!g198) & (!sk[104]) & (g199) & (g201)) + ((g121) & (!g194) & (!g198) & (sk[104]) & (!g199) & (g201)) + ((g121) & (!g194) & (g198) & (!sk[104]) & (!g199) & (!g201)) + ((g121) & (!g194) & (g198) & (!sk[104]) & (!g199) & (g201)) + ((g121) & (!g194) & (g198) & (!sk[104]) & (g199) & (!g201)) + ((g121) & (!g194) & (g198) & (!sk[104]) & (g199) & (g201)) + ((g121) & (g194) & (!g198) & (!sk[104]) & (!g199) & (!g201)) + ((g121) & (g194) & (!g198) & (!sk[104]) & (!g199) & (g201)) + ((g121) & (g194) & (!g198) & (!sk[104]) & (g199) & (!g201)) + ((g121) & (g194) & (!g198) & (!sk[104]) & (g199) & (g201)) + ((g121) & (g194) & (g198) & (!sk[104]) & (!g199) & (!g201)) + ((g121) & (g194) & (g198) & (!sk[104]) & (!g199) & (g201)) + ((g121) & (g194) & (g198) & (!sk[104]) & (g199) & (!g201)) + ((g121) & (g194) & (g198) & (!sk[104]) & (g199) & (g201)));
	assign g203 = (((!g75) & (!g164) & (!g122) & (!g194) & (!g197) & (g202)) + ((!g75) & (!g164) & (!g122) & (g194) & (!g197) & (g202)) + ((!g75) & (!g164) & (g122) & (!g194) & (!g197) & (g202)) + ((!g75) & (g164) & (!g122) & (!g194) & (!g197) & (g202)) + ((!g75) & (g164) & (!g122) & (g194) & (!g197) & (g202)) + ((!g75) & (g164) & (g122) & (!g194) & (!g197) & (g202)) + ((g75) & (!g164) & (!g122) & (!g194) & (!g197) & (g202)) + ((g75) & (!g164) & (!g122) & (!g194) & (g197) & (g202)) + ((g75) & (!g164) & (!g122) & (g194) & (!g197) & (g202)) + ((g75) & (!g164) & (!g122) & (g194) & (g197) & (g202)) + ((g75) & (!g164) & (g122) & (!g194) & (!g197) & (g202)) + ((g75) & (!g164) & (g122) & (!g194) & (g197) & (g202)) + ((g75) & (g164) & (!g122) & (!g194) & (!g197) & (g202)) + ((g75) & (g164) & (!g122) & (g194) & (!g197) & (g202)) + ((g75) & (g164) & (g122) & (!g194) & (!g197) & (g202)));
	assign g204 = (((!g125) & (!sk[106]) & (!g131) & (!g185) & (g186) & (!g192)) + ((!g125) & (!sk[106]) & (!g131) & (!g185) & (g186) & (g192)) + ((!g125) & (!sk[106]) & (!g131) & (g185) & (!g186) & (!g192)) + ((!g125) & (!sk[106]) & (!g131) & (g185) & (!g186) & (g192)) + ((!g125) & (!sk[106]) & (!g131) & (g185) & (g186) & (!g192)) + ((!g125) & (!sk[106]) & (!g131) & (g185) & (g186) & (g192)) + ((!g125) & (!sk[106]) & (g131) & (!g185) & (!g186) & (!g192)) + ((!g125) & (!sk[106]) & (g131) & (!g185) & (!g186) & (g192)) + ((!g125) & (!sk[106]) & (g131) & (!g185) & (g186) & (!g192)) + ((!g125) & (!sk[106]) & (g131) & (!g185) & (g186) & (g192)) + ((!g125) & (!sk[106]) & (g131) & (g185) & (!g186) & (!g192)) + ((!g125) & (!sk[106]) & (g131) & (g185) & (!g186) & (g192)) + ((!g125) & (!sk[106]) & (g131) & (g185) & (g186) & (!g192)) + ((!g125) & (!sk[106]) & (g131) & (g185) & (g186) & (g192)) + ((!g125) & (sk[106]) & (!g131) & (!g185) & (!g186) & (!g192)) + ((!g125) & (sk[106]) & (!g131) & (g185) & (!g186) & (!g192)) + ((!g125) & (sk[106]) & (g131) & (!g185) & (!g186) & (!g192)) + ((!g125) & (sk[106]) & (g131) & (!g185) & (!g186) & (g192)) + ((!g125) & (sk[106]) & (g131) & (!g185) & (g186) & (!g192)) + ((!g125) & (sk[106]) & (g131) & (!g185) & (g186) & (g192)) + ((!g125) & (sk[106]) & (g131) & (g185) & (!g186) & (!g192)) + ((!g125) & (sk[106]) & (g131) & (g185) & (!g186) & (g192)) + ((!g125) & (sk[106]) & (g131) & (g185) & (g186) & (!g192)) + ((!g125) & (sk[106]) & (g131) & (g185) & (g186) & (g192)) + ((g125) & (!sk[106]) & (!g131) & (!g185) & (g186) & (!g192)) + ((g125) & (!sk[106]) & (!g131) & (!g185) & (g186) & (g192)) + ((g125) & (!sk[106]) & (!g131) & (g185) & (!g186) & (!g192)) + ((g125) & (!sk[106]) & (!g131) & (g185) & (!g186) & (g192)) + ((g125) & (!sk[106]) & (!g131) & (g185) & (g186) & (!g192)) + ((g125) & (!sk[106]) & (!g131) & (g185) & (g186) & (g192)) + ((g125) & (!sk[106]) & (g131) & (!g185) & (!g186) & (!g192)) + ((g125) & (!sk[106]) & (g131) & (!g185) & (!g186) & (g192)) + ((g125) & (!sk[106]) & (g131) & (!g185) & (g186) & (!g192)) + ((g125) & (!sk[106]) & (g131) & (!g185) & (g186) & (g192)) + ((g125) & (!sk[106]) & (g131) & (g185) & (!g186) & (!g192)) + ((g125) & (!sk[106]) & (g131) & (g185) & (!g186) & (g192)) + ((g125) & (!sk[106]) & (g131) & (g185) & (g186) & (!g192)) + ((g125) & (!sk[106]) & (g131) & (g185) & (g186) & (g192)) + ((g125) & (sk[106]) & (!g131) & (!g185) & (!g186) & (!g192)) + ((g125) & (sk[106]) & (g131) & (!g185) & (!g186) & (!g192)) + ((g125) & (sk[106]) & (g131) & (!g185) & (!g186) & (g192)) + ((g125) & (sk[106]) & (g131) & (!g185) & (g186) & (!g192)) + ((g125) & (sk[106]) & (g131) & (!g185) & (g186) & (g192)));
	assign g205 = (((!g125) & (!sk[107]) & (g194) & (!g188)) + ((!g125) & (!sk[107]) & (g194) & (g188)) + ((g125) & (!sk[107]) & (!g194) & (g188)) + ((g125) & (!sk[107]) & (g194) & (!g188)) + ((g125) & (!sk[107]) & (g194) & (g188)) + ((g125) & (sk[107]) & (!g194) & (g188)) + ((g125) & (sk[107]) & (g194) & (!g188)) + ((g125) & (sk[107]) & (g194) & (g188)));
	assign g206 = (((!sk[108]) & (!g131) & (g191) & (!g187)) + ((!sk[108]) & (!g131) & (g191) & (g187)) + ((!sk[108]) & (g131) & (!g191) & (g187)) + ((!sk[108]) & (g131) & (g191) & (!g187)) + ((!sk[108]) & (g131) & (g191) & (g187)) + ((sk[108]) & (!g131) & (!g191) & (g187)) + ((sk[108]) & (!g131) & (g191) & (!g187)) + ((sk[108]) & (!g131) & (g191) & (g187)));
	assign g207 = (((!g125) & (!sk[109]) & (g175) & (!g177)) + ((!g125) & (!sk[109]) & (g175) & (g177)) + ((g125) & (!sk[109]) & (!g175) & (g177)) + ((g125) & (!sk[109]) & (g175) & (!g177)) + ((g125) & (!sk[109]) & (g175) & (g177)) + ((g125) & (sk[109]) & (!g175) & (g177)) + ((g125) & (sk[109]) & (g175) & (!g177)) + ((g125) & (sk[109]) & (g175) & (g177)));
	assign g208 = (((!g131) & (!sk[110]) & (g179) & (!g177)) + ((!g131) & (!sk[110]) & (g179) & (g177)) + ((!g131) & (sk[110]) & (!g179) & (g177)) + ((!g131) & (sk[110]) & (g179) & (!g177)) + ((!g131) & (sk[110]) & (g179) & (g177)) + ((g131) & (!sk[110]) & (!g179) & (g177)) + ((g131) & (!sk[110]) & (g179) & (!g177)) + ((g131) & (!sk[110]) & (g179) & (g177)));
	assign g209 = (((!sk[111]) & (!g125) & (!g179) & (!g186) & (g187) & (!g182)) + ((!sk[111]) & (!g125) & (!g179) & (!g186) & (g187) & (g182)) + ((!sk[111]) & (!g125) & (!g179) & (g186) & (!g187) & (!g182)) + ((!sk[111]) & (!g125) & (!g179) & (g186) & (!g187) & (g182)) + ((!sk[111]) & (!g125) & (!g179) & (g186) & (g187) & (!g182)) + ((!sk[111]) & (!g125) & (!g179) & (g186) & (g187) & (g182)) + ((!sk[111]) & (!g125) & (g179) & (!g186) & (!g187) & (!g182)) + ((!sk[111]) & (!g125) & (g179) & (!g186) & (!g187) & (g182)) + ((!sk[111]) & (!g125) & (g179) & (!g186) & (g187) & (!g182)) + ((!sk[111]) & (!g125) & (g179) & (!g186) & (g187) & (g182)) + ((!sk[111]) & (!g125) & (g179) & (g186) & (!g187) & (!g182)) + ((!sk[111]) & (!g125) & (g179) & (g186) & (!g187) & (g182)) + ((!sk[111]) & (!g125) & (g179) & (g186) & (g187) & (!g182)) + ((!sk[111]) & (!g125) & (g179) & (g186) & (g187) & (g182)) + ((!sk[111]) & (g125) & (!g179) & (!g186) & (g187) & (!g182)) + ((!sk[111]) & (g125) & (!g179) & (!g186) & (g187) & (g182)) + ((!sk[111]) & (g125) & (!g179) & (g186) & (!g187) & (!g182)) + ((!sk[111]) & (g125) & (!g179) & (g186) & (!g187) & (g182)) + ((!sk[111]) & (g125) & (!g179) & (g186) & (g187) & (!g182)) + ((!sk[111]) & (g125) & (!g179) & (g186) & (g187) & (g182)) + ((!sk[111]) & (g125) & (g179) & (!g186) & (!g187) & (!g182)) + ((!sk[111]) & (g125) & (g179) & (!g186) & (!g187) & (g182)) + ((!sk[111]) & (g125) & (g179) & (!g186) & (g187) & (!g182)) + ((!sk[111]) & (g125) & (g179) & (!g186) & (g187) & (g182)) + ((!sk[111]) & (g125) & (g179) & (g186) & (!g187) & (!g182)) + ((!sk[111]) & (g125) & (g179) & (g186) & (!g187) & (g182)) + ((!sk[111]) & (g125) & (g179) & (g186) & (g187) & (!g182)) + ((!sk[111]) & (g125) & (g179) & (g186) & (g187) & (g182)) + ((sk[111]) & (g125) & (!g179) & (!g186) & (!g187) & (g182)) + ((sk[111]) & (g125) & (!g179) & (!g186) & (g187) & (!g182)) + ((sk[111]) & (g125) & (!g179) & (!g186) & (g187) & (g182)) + ((sk[111]) & (g125) & (!g179) & (g186) & (!g187) & (!g182)) + ((sk[111]) & (g125) & (!g179) & (g186) & (!g187) & (g182)) + ((sk[111]) & (g125) & (!g179) & (g186) & (g187) & (!g182)) + ((sk[111]) & (g125) & (!g179) & (g186) & (g187) & (g182)) + ((sk[111]) & (g125) & (g179) & (!g186) & (!g187) & (!g182)) + ((sk[111]) & (g125) & (g179) & (!g186) & (!g187) & (g182)) + ((sk[111]) & (g125) & (g179) & (!g186) & (g187) & (!g182)) + ((sk[111]) & (g125) & (g179) & (!g186) & (g187) & (g182)) + ((sk[111]) & (g125) & (g179) & (g186) & (!g187) & (!g182)) + ((sk[111]) & (g125) & (g179) & (g186) & (!g187) & (g182)) + ((sk[111]) & (g125) & (g179) & (g186) & (g187) & (!g182)) + ((sk[111]) & (g125) & (g179) & (g186) & (g187) & (g182)));
	assign g210 = (((!sk[112]) & (!g205) & (!g206) & (!g207) & (g208) & (!g209)) + ((!sk[112]) & (!g205) & (!g206) & (!g207) & (g208) & (g209)) + ((!sk[112]) & (!g205) & (!g206) & (g207) & (!g208) & (!g209)) + ((!sk[112]) & (!g205) & (!g206) & (g207) & (!g208) & (g209)) + ((!sk[112]) & (!g205) & (!g206) & (g207) & (g208) & (!g209)) + ((!sk[112]) & (!g205) & (!g206) & (g207) & (g208) & (g209)) + ((!sk[112]) & (!g205) & (g206) & (!g207) & (!g208) & (!g209)) + ((!sk[112]) & (!g205) & (g206) & (!g207) & (!g208) & (g209)) + ((!sk[112]) & (!g205) & (g206) & (!g207) & (g208) & (!g209)) + ((!sk[112]) & (!g205) & (g206) & (!g207) & (g208) & (g209)) + ((!sk[112]) & (!g205) & (g206) & (g207) & (!g208) & (!g209)) + ((!sk[112]) & (!g205) & (g206) & (g207) & (!g208) & (g209)) + ((!sk[112]) & (!g205) & (g206) & (g207) & (g208) & (!g209)) + ((!sk[112]) & (!g205) & (g206) & (g207) & (g208) & (g209)) + ((!sk[112]) & (g205) & (!g206) & (!g207) & (g208) & (!g209)) + ((!sk[112]) & (g205) & (!g206) & (!g207) & (g208) & (g209)) + ((!sk[112]) & (g205) & (!g206) & (g207) & (!g208) & (!g209)) + ((!sk[112]) & (g205) & (!g206) & (g207) & (!g208) & (g209)) + ((!sk[112]) & (g205) & (!g206) & (g207) & (g208) & (!g209)) + ((!sk[112]) & (g205) & (!g206) & (g207) & (g208) & (g209)) + ((!sk[112]) & (g205) & (g206) & (!g207) & (!g208) & (!g209)) + ((!sk[112]) & (g205) & (g206) & (!g207) & (!g208) & (g209)) + ((!sk[112]) & (g205) & (g206) & (!g207) & (g208) & (!g209)) + ((!sk[112]) & (g205) & (g206) & (!g207) & (g208) & (g209)) + ((!sk[112]) & (g205) & (g206) & (g207) & (!g208) & (!g209)) + ((!sk[112]) & (g205) & (g206) & (g207) & (!g208) & (g209)) + ((!sk[112]) & (g205) & (g206) & (g207) & (g208) & (!g209)) + ((!sk[112]) & (g205) & (g206) & (g207) & (g208) & (g209)) + ((sk[112]) & (!g205) & (!g206) & (!g207) & (!g208) & (!g209)));
	assign g211 = (((!g131) & (!sk[113]) & (!g182) & (!g183) & (g204) & (!g210)) + ((!g131) & (!sk[113]) & (!g182) & (!g183) & (g204) & (g210)) + ((!g131) & (!sk[113]) & (!g182) & (g183) & (!g204) & (!g210)) + ((!g131) & (!sk[113]) & (!g182) & (g183) & (!g204) & (g210)) + ((!g131) & (!sk[113]) & (!g182) & (g183) & (g204) & (!g210)) + ((!g131) & (!sk[113]) & (!g182) & (g183) & (g204) & (g210)) + ((!g131) & (!sk[113]) & (g182) & (!g183) & (!g204) & (!g210)) + ((!g131) & (!sk[113]) & (g182) & (!g183) & (!g204) & (g210)) + ((!g131) & (!sk[113]) & (g182) & (!g183) & (g204) & (!g210)) + ((!g131) & (!sk[113]) & (g182) & (!g183) & (g204) & (g210)) + ((!g131) & (!sk[113]) & (g182) & (g183) & (!g204) & (!g210)) + ((!g131) & (!sk[113]) & (g182) & (g183) & (!g204) & (g210)) + ((!g131) & (!sk[113]) & (g182) & (g183) & (g204) & (!g210)) + ((!g131) & (!sk[113]) & (g182) & (g183) & (g204) & (g210)) + ((!g131) & (sk[113]) & (!g182) & (!g183) & (g204) & (g210)) + ((g131) & (!sk[113]) & (!g182) & (!g183) & (g204) & (!g210)) + ((g131) & (!sk[113]) & (!g182) & (!g183) & (g204) & (g210)) + ((g131) & (!sk[113]) & (!g182) & (g183) & (!g204) & (!g210)) + ((g131) & (!sk[113]) & (!g182) & (g183) & (!g204) & (g210)) + ((g131) & (!sk[113]) & (!g182) & (g183) & (g204) & (!g210)) + ((g131) & (!sk[113]) & (!g182) & (g183) & (g204) & (g210)) + ((g131) & (!sk[113]) & (g182) & (!g183) & (!g204) & (!g210)) + ((g131) & (!sk[113]) & (g182) & (!g183) & (!g204) & (g210)) + ((g131) & (!sk[113]) & (g182) & (!g183) & (g204) & (!g210)) + ((g131) & (!sk[113]) & (g182) & (!g183) & (g204) & (g210)) + ((g131) & (!sk[113]) & (g182) & (g183) & (!g204) & (!g210)) + ((g131) & (!sk[113]) & (g182) & (g183) & (!g204) & (g210)) + ((g131) & (!sk[113]) & (g182) & (g183) & (g204) & (!g210)) + ((g131) & (!sk[113]) & (g182) & (g183) & (g204) & (g210)) + ((g131) & (sk[113]) & (!g182) & (!g183) & (g204) & (g210)) + ((g131) & (sk[113]) & (!g182) & (g183) & (g204) & (g210)) + ((g131) & (sk[113]) & (g182) & (!g183) & (g204) & (g210)) + ((g131) & (sk[113]) & (g182) & (g183) & (g204) & (g210)));
	assign g212 = (((!sk[114]) & (!g107) & (g174)) + ((!sk[114]) & (g107) & (g174)) + ((sk[114]) & (!g107) & (!g174)));
	assign g213 = (((!sk[115]) & (!g45) & (g118)) + ((!sk[115]) & (g45) & (g118)) + ((sk[115]) & (g45) & (g118)));
	assign g214 = (((!sk[116]) & (!g135) & (g159) & (!g183)) + ((!sk[116]) & (!g135) & (g159) & (g183)) + ((!sk[116]) & (g135) & (!g159) & (g183)) + ((!sk[116]) & (g135) & (g159) & (!g183)) + ((!sk[116]) & (g135) & (g159) & (g183)) + ((sk[116]) & (!g135) & (!g159) & (g183)) + ((sk[116]) & (!g135) & (g159) & (g183)) + ((sk[116]) & (g135) & (!g159) & (g183)));
	assign g215 = (((!g75) & (!g105) & (sk[117]) & (!g191) & (g180)) + ((!g75) & (!g105) & (sk[117]) & (g191) & (!g180)) + ((!g75) & (!g105) & (sk[117]) & (g191) & (g180)) + ((!g75) & (g105) & (!sk[117]) & (!g191) & (!g180)) + ((!g75) & (g105) & (!sk[117]) & (!g191) & (g180)) + ((!g75) & (g105) & (!sk[117]) & (g191) & (!g180)) + ((!g75) & (g105) & (!sk[117]) & (g191) & (g180)) + ((!g75) & (g105) & (sk[117]) & (g191) & (!g180)) + ((!g75) & (g105) & (sk[117]) & (g191) & (g180)) + ((g75) & (!g105) & (sk[117]) & (!g191) & (g180)) + ((g75) & (!g105) & (sk[117]) & (g191) & (g180)) + ((g75) & (g105) & (!sk[117]) & (!g191) & (!g180)) + ((g75) & (g105) & (!sk[117]) & (!g191) & (g180)) + ((g75) & (g105) & (!sk[117]) & (g191) & (!g180)) + ((g75) & (g105) & (!sk[117]) & (g191) & (g180)));
	assign g216 = (((!g131) & (!g194) & (!g212) & (!g213) & (!g214) & (!g215)) + ((!g131) & (!g194) & (!g212) & (g213) & (!g214) & (!g215)) + ((!g131) & (g194) & (!g212) & (!g213) & (!g214) & (!g215)) + ((g131) & (!g194) & (!g212) & (!g213) & (!g214) & (!g215)) + ((g131) & (!g194) & (!g212) & (g213) & (!g214) & (!g215)) + ((g131) & (!g194) & (g212) & (!g213) & (!g214) & (!g215)) + ((g131) & (!g194) & (g212) & (g213) & (!g214) & (!g215)) + ((g131) & (g194) & (!g212) & (!g213) & (!g214) & (!g215)) + ((g131) & (g194) & (g212) & (!g213) & (!g214) & (!g215)));
	assign g217 = (((!g10) & (!sk[119]) & (g120)) + ((g10) & (!sk[119]) & (g120)) + ((g10) & (sk[119]) & (g120)));
	assign g218 = (((!i_8_) & (!sk[120]) & (i_6_) & (!g120)) + ((!i_8_) & (!sk[120]) & (i_6_) & (g120)) + ((i_8_) & (!sk[120]) & (!i_6_) & (g120)) + ((i_8_) & (!sk[120]) & (i_6_) & (!g120)) + ((i_8_) & (!sk[120]) & (i_6_) & (g120)) + ((i_8_) & (sk[120]) & (!i_6_) & (g120)));
	assign g219 = (((!i_10_) & (i_11_) & (!i_15_) & (!sk[121]) & (!g174)) + ((!i_10_) & (i_11_) & (!i_15_) & (!sk[121]) & (g174)) + ((!i_10_) & (i_11_) & (i_15_) & (!sk[121]) & (!g174)) + ((!i_10_) & (i_11_) & (i_15_) & (!sk[121]) & (g174)) + ((i_10_) & (i_11_) & (!i_15_) & (!sk[121]) & (!g174)) + ((i_10_) & (i_11_) & (!i_15_) & (!sk[121]) & (g174)) + ((i_10_) & (i_11_) & (!i_15_) & (sk[121]) & (!g174)) + ((i_10_) & (i_11_) & (i_15_) & (!sk[121]) & (!g174)) + ((i_10_) & (i_11_) & (i_15_) & (!sk[121]) & (g174)));
	assign g220 = (((!g165) & (!g217) & (g200) & (!g212) & (g218) & (g219)) + ((!g165) & (!g217) & (g200) & (g212) & (g218) & (g219)) + ((!g165) & (g217) & (!g200) & (!g212) & (g218) & (g219)) + ((!g165) & (g217) & (!g200) & (g212) & (!g218) & (g219)) + ((!g165) & (g217) & (!g200) & (g212) & (g218) & (g219)) + ((!g165) & (g217) & (g200) & (!g212) & (g218) & (g219)) + ((!g165) & (g217) & (g200) & (g212) & (!g218) & (g219)) + ((!g165) & (g217) & (g200) & (g212) & (g218) & (g219)) + ((g165) & (!g217) & (!g200) & (!g212) & (g218) & (g219)) + ((g165) & (!g217) & (!g200) & (g212) & (!g218) & (g219)) + ((g165) & (!g217) & (!g200) & (g212) & (g218) & (g219)) + ((g165) & (!g217) & (g200) & (!g212) & (g218) & (g219)) + ((g165) & (!g217) & (g200) & (g212) & (!g218) & (g219)) + ((g165) & (!g217) & (g200) & (g212) & (g218) & (g219)) + ((g165) & (g217) & (!g200) & (!g212) & (g218) & (g219)) + ((g165) & (g217) & (!g200) & (g212) & (!g218) & (g219)) + ((g165) & (g217) & (!g200) & (g212) & (g218) & (g219)) + ((g165) & (g217) & (g200) & (!g212) & (g218) & (g219)) + ((g165) & (g217) & (g200) & (g212) & (!g218) & (g219)) + ((g165) & (g217) & (g200) & (g212) & (g218) & (g219)));
	assign g221 = (((!g165) & (!sk[123]) & (g179)) + ((g165) & (!sk[123]) & (g179)) + ((g165) & (sk[123]) & (g179)));
	assign g222 = (((!g122) & (g175) & (!sk[124]) & (!g177)) + ((!g122) & (g175) & (!sk[124]) & (g177)) + ((g122) & (!g175) & (!sk[124]) & (g177)) + ((g122) & (!g175) & (sk[124]) & (g177)) + ((g122) & (g175) & (!sk[124]) & (!g177)) + ((g122) & (g175) & (!sk[124]) & (g177)) + ((g122) & (g175) & (sk[124]) & (!g177)) + ((g122) & (g175) & (sk[124]) & (g177)));
	assign g223 = (((!g135) & (!sk[125]) & (g122) & (!g180) & (!g183)) + ((!g135) & (!sk[125]) & (g122) & (!g180) & (g183)) + ((!g135) & (!sk[125]) & (g122) & (g180) & (!g183)) + ((!g135) & (!sk[125]) & (g122) & (g180) & (g183)) + ((!g135) & (sk[125]) & (!g122) & (!g180) & (!g183)) + ((!g135) & (sk[125]) & (!g122) & (!g180) & (g183)) + ((!g135) & (sk[125]) & (g122) & (!g180) & (!g183)) + ((g135) & (!sk[125]) & (g122) & (!g180) & (!g183)) + ((g135) & (!sk[125]) & (g122) & (!g180) & (g183)) + ((g135) & (!sk[125]) & (g122) & (g180) & (!g183)) + ((g135) & (!sk[125]) & (g122) & (g180) & (g183)) + ((g135) & (sk[125]) & (!g122) & (!g180) & (!g183)) + ((g135) & (sk[125]) & (!g122) & (!g180) & (g183)) + ((g135) & (sk[125]) & (!g122) & (g180) & (!g183)) + ((g135) & (sk[125]) & (!g122) & (g180) & (g183)) + ((g135) & (sk[125]) & (g122) & (!g180) & (!g183)));
	assign g224 = (((!g135) & (!g122) & (!g185) & (!g191) & (!g186) & (!g187)) + ((!g135) & (!g122) & (g185) & (!g191) & (!g186) & (!g187)) + ((!g135) & (g122) & (!g185) & (!g191) & (!g186) & (!g187)) + ((g135) & (!g122) & (!g185) & (!g191) & (!g186) & (!g187)) + ((g135) & (!g122) & (!g185) & (!g191) & (!g186) & (g187)) + ((g135) & (!g122) & (!g185) & (!g191) & (g186) & (!g187)) + ((g135) & (!g122) & (!g185) & (!g191) & (g186) & (g187)) + ((g135) & (!g122) & (!g185) & (g191) & (!g186) & (!g187)) + ((g135) & (!g122) & (!g185) & (g191) & (!g186) & (g187)) + ((g135) & (!g122) & (!g185) & (g191) & (g186) & (!g187)) + ((g135) & (!g122) & (!g185) & (g191) & (g186) & (g187)) + ((g135) & (!g122) & (g185) & (!g191) & (!g186) & (!g187)) + ((g135) & (!g122) & (g185) & (!g191) & (!g186) & (g187)) + ((g135) & (!g122) & (g185) & (!g191) & (g186) & (!g187)) + ((g135) & (!g122) & (g185) & (!g191) & (g186) & (g187)) + ((g135) & (!g122) & (g185) & (g191) & (!g186) & (!g187)) + ((g135) & (!g122) & (g185) & (g191) & (!g186) & (g187)) + ((g135) & (!g122) & (g185) & (g191) & (g186) & (!g187)) + ((g135) & (!g122) & (g185) & (g191) & (g186) & (g187)) + ((g135) & (g122) & (!g185) & (!g191) & (!g186) & (!g187)) + ((g135) & (g122) & (!g185) & (!g191) & (!g186) & (g187)) + ((g135) & (g122) & (!g185) & (g191) & (!g186) & (!g187)) + ((g135) & (g122) & (!g185) & (g191) & (!g186) & (g187)));
	assign g225 = (((!sk[127]) & (g120) & (!g101)) + ((!sk[127]) & (g120) & (g101)) + ((sk[127]) & (g120) & (g101)));
	assign g226 = (((!sk[0]) & (!i_8_) & (!g45) & (g118)) + ((!sk[0]) & (!i_8_) & (g45) & (!g118)) + ((!sk[0]) & (!i_8_) & (g45) & (g118)) + ((!sk[0]) & (i_8_) & (!g45) & (g118)) + ((!sk[0]) & (i_8_) & (g45) & (!g118)) + ((!sk[0]) & (i_8_) & (g45) & (g118)) + ((sk[0]) & (!i_8_) & (!g45) & (!g118)) + ((sk[0]) & (!i_8_) & (!g45) & (g118)) + ((sk[0]) & (!i_8_) & (g45) & (!g118)) + ((sk[0]) & (!i_8_) & (g45) & (g118)) + ((sk[0]) & (i_8_) & (!g45) & (!g118)) + ((sk[0]) & (i_8_) & (!g45) & (g118)) + ((sk[0]) & (i_8_) & (g45) & (!g118)));
	assign g227 = (((!sk[1]) & (g101) & (!g118)) + ((!sk[1]) & (g101) & (g118)) + ((sk[1]) & (g101) & (g118)));
	assign g228 = (((!sk[2]) & (!g179) & (!g225) & (g226) & (!g227)) + ((!sk[2]) & (!g179) & (!g225) & (g226) & (g227)) + ((!sk[2]) & (!g179) & (g225) & (g226) & (!g227)) + ((!sk[2]) & (!g179) & (g225) & (g226) & (g227)) + ((!sk[2]) & (g179) & (!g225) & (g226) & (!g227)) + ((!sk[2]) & (g179) & (!g225) & (g226) & (g227)) + ((!sk[2]) & (g179) & (g225) & (g226) & (!g227)) + ((!sk[2]) & (g179) & (g225) & (g226) & (g227)) + ((sk[2]) & (g179) & (!g225) & (!g226) & (!g227)) + ((sk[2]) & (g179) & (!g225) & (!g226) & (g227)) + ((sk[2]) & (g179) & (!g225) & (g226) & (g227)) + ((sk[2]) & (g179) & (g225) & (!g226) & (!g227)) + ((sk[2]) & (g179) & (g225) & (!g226) & (g227)) + ((sk[2]) & (g179) & (g225) & (g226) & (!g227)) + ((sk[2]) & (g179) & (g225) & (g226) & (g227)));
	assign g229 = (((!sk[3]) & (!g221) & (!g222) & (g223) & (!g224) & (g228)) + ((!sk[3]) & (!g221) & (!g222) & (g223) & (g224) & (!g228)) + ((!sk[3]) & (!g221) & (!g222) & (g223) & (g224) & (g228)) + ((!sk[3]) & (!g221) & (g222) & (!g223) & (!g224) & (!g228)) + ((!sk[3]) & (!g221) & (g222) & (!g223) & (!g224) & (g228)) + ((!sk[3]) & (!g221) & (g222) & (!g223) & (g224) & (!g228)) + ((!sk[3]) & (!g221) & (g222) & (!g223) & (g224) & (g228)) + ((!sk[3]) & (!g221) & (g222) & (g223) & (!g224) & (!g228)) + ((!sk[3]) & (!g221) & (g222) & (g223) & (!g224) & (g228)) + ((!sk[3]) & (!g221) & (g222) & (g223) & (g224) & (!g228)) + ((!sk[3]) & (!g221) & (g222) & (g223) & (g224) & (g228)) + ((!sk[3]) & (g221) & (!g222) & (g223) & (!g224) & (g228)) + ((!sk[3]) & (g221) & (!g222) & (g223) & (g224) & (!g228)) + ((!sk[3]) & (g221) & (!g222) & (g223) & (g224) & (g228)) + ((!sk[3]) & (g221) & (g222) & (!g223) & (!g224) & (!g228)) + ((!sk[3]) & (g221) & (g222) & (!g223) & (!g224) & (g228)) + ((!sk[3]) & (g221) & (g222) & (!g223) & (g224) & (!g228)) + ((!sk[3]) & (g221) & (g222) & (!g223) & (g224) & (g228)) + ((!sk[3]) & (g221) & (g222) & (g223) & (!g224) & (!g228)) + ((!sk[3]) & (g221) & (g222) & (g223) & (!g224) & (g228)) + ((!sk[3]) & (g221) & (g222) & (g223) & (g224) & (!g228)) + ((!sk[3]) & (g221) & (g222) & (g223) & (g224) & (g228)) + ((sk[3]) & (!g221) & (!g222) & (g223) & (g224) & (!g228)));
	assign g230 = (((!g123) & (!g192) & (!g200) & (sk[4]) & (g212)) + ((!g123) & (!g192) & (g200) & (!sk[4]) & (!g212)) + ((!g123) & (!g192) & (g200) & (!sk[4]) & (g212)) + ((!g123) & (!g192) & (g200) & (sk[4]) & (!g212)) + ((!g123) & (!g192) & (g200) & (sk[4]) & (g212)) + ((!g123) & (g192) & (!g200) & (sk[4]) & (!g212)) + ((!g123) & (g192) & (!g200) & (sk[4]) & (g212)) + ((!g123) & (g192) & (g200) & (!sk[4]) & (!g212)) + ((!g123) & (g192) & (g200) & (!sk[4]) & (g212)) + ((!g123) & (g192) & (g200) & (sk[4]) & (!g212)) + ((!g123) & (g192) & (g200) & (sk[4]) & (g212)) + ((g123) & (!g192) & (g200) & (!sk[4]) & (!g212)) + ((g123) & (!g192) & (g200) & (!sk[4]) & (g212)) + ((g123) & (g192) & (g200) & (!sk[4]) & (!g212)) + ((g123) & (g192) & (g200) & (!sk[4]) & (g212)));
	assign g231 = (((!sk[5]) & (!g122) & (!g123) & (g191)) + ((!sk[5]) & (!g122) & (g123) & (!g191)) + ((!sk[5]) & (!g122) & (g123) & (g191)) + ((!sk[5]) & (g122) & (!g123) & (g191)) + ((!sk[5]) & (g122) & (g123) & (!g191)) + ((!sk[5]) & (g122) & (g123) & (g191)) + ((sk[5]) & (!g122) & (!g123) & (g191)) + ((sk[5]) & (g122) & (!g123) & (g191)) + ((sk[5]) & (g122) & (g123) & (g191)));
	assign g232 = (((!g161) & (!g122) & (!sk[6]) & (g187)) + ((!g161) & (g122) & (!sk[6]) & (!g187)) + ((!g161) & (g122) & (!sk[6]) & (g187)) + ((!g161) & (g122) & (sk[6]) & (g187)) + ((g161) & (!g122) & (!sk[6]) & (g187)) + ((g161) & (!g122) & (sk[6]) & (g187)) + ((g161) & (g122) & (!sk[6]) & (!g187)) + ((g161) & (g122) & (!sk[6]) & (g187)) + ((g161) & (g122) & (sk[6]) & (g187)));
	assign g233 = (((!g105) & (!g191) & (!sk[7]) & (g175) & (!g200)) + ((!g105) & (!g191) & (!sk[7]) & (g175) & (g200)) + ((!g105) & (!g191) & (sk[7]) & (!g175) & (g200)) + ((!g105) & (!g191) & (sk[7]) & (g175) & (!g200)) + ((!g105) & (!g191) & (sk[7]) & (g175) & (g200)) + ((!g105) & (g191) & (!sk[7]) & (g175) & (!g200)) + ((!g105) & (g191) & (!sk[7]) & (g175) & (g200)) + ((!g105) & (g191) & (sk[7]) & (!g175) & (!g200)) + ((!g105) & (g191) & (sk[7]) & (!g175) & (g200)) + ((!g105) & (g191) & (sk[7]) & (g175) & (!g200)) + ((!g105) & (g191) & (sk[7]) & (g175) & (g200)) + ((g105) & (!g191) & (!sk[7]) & (g175) & (!g200)) + ((g105) & (!g191) & (!sk[7]) & (g175) & (g200)) + ((g105) & (g191) & (!sk[7]) & (g175) & (!g200)) + ((g105) & (g191) & (!sk[7]) & (g175) & (g200)));
	assign g234 = (((!g142) & (!g130) & (!g180) & (!g182) & (sk[8]) & (!g183)) + ((!g142) & (!g130) & (g180) & (!g182) & (!sk[8]) & (g183)) + ((!g142) & (!g130) & (g180) & (g182) & (!sk[8]) & (!g183)) + ((!g142) & (!g130) & (g180) & (g182) & (!sk[8]) & (g183)) + ((!g142) & (g130) & (!g180) & (!g182) & (!sk[8]) & (!g183)) + ((!g142) & (g130) & (!g180) & (!g182) & (!sk[8]) & (g183)) + ((!g142) & (g130) & (!g180) & (!g182) & (sk[8]) & (!g183)) + ((!g142) & (g130) & (!g180) & (g182) & (!sk[8]) & (!g183)) + ((!g142) & (g130) & (!g180) & (g182) & (!sk[8]) & (g183)) + ((!g142) & (g130) & (!g180) & (g182) & (sk[8]) & (!g183)) + ((!g142) & (g130) & (g180) & (!g182) & (!sk[8]) & (!g183)) + ((!g142) & (g130) & (g180) & (!g182) & (!sk[8]) & (g183)) + ((!g142) & (g130) & (g180) & (g182) & (!sk[8]) & (!g183)) + ((!g142) & (g130) & (g180) & (g182) & (!sk[8]) & (g183)) + ((g142) & (!g130) & (!g180) & (!g182) & (sk[8]) & (!g183)) + ((g142) & (!g130) & (g180) & (!g182) & (!sk[8]) & (g183)) + ((g142) & (!g130) & (g180) & (!g182) & (sk[8]) & (!g183)) + ((g142) & (!g130) & (g180) & (g182) & (!sk[8]) & (!g183)) + ((g142) & (!g130) & (g180) & (g182) & (!sk[8]) & (g183)) + ((g142) & (g130) & (!g180) & (!g182) & (!sk[8]) & (!g183)) + ((g142) & (g130) & (!g180) & (!g182) & (!sk[8]) & (g183)) + ((g142) & (g130) & (!g180) & (!g182) & (sk[8]) & (!g183)) + ((g142) & (g130) & (!g180) & (!g182) & (sk[8]) & (g183)) + ((g142) & (g130) & (!g180) & (g182) & (!sk[8]) & (!g183)) + ((g142) & (g130) & (!g180) & (g182) & (!sk[8]) & (g183)) + ((g142) & (g130) & (!g180) & (g182) & (sk[8]) & (!g183)) + ((g142) & (g130) & (!g180) & (g182) & (sk[8]) & (g183)) + ((g142) & (g130) & (g180) & (!g182) & (!sk[8]) & (!g183)) + ((g142) & (g130) & (g180) & (!g182) & (!sk[8]) & (g183)) + ((g142) & (g130) & (g180) & (!g182) & (sk[8]) & (!g183)) + ((g142) & (g130) & (g180) & (!g182) & (sk[8]) & (g183)) + ((g142) & (g130) & (g180) & (g182) & (!sk[8]) & (!g183)) + ((g142) & (g130) & (g180) & (g182) & (!sk[8]) & (g183)) + ((g142) & (g130) & (g180) & (g182) & (sk[8]) & (!g183)) + ((g142) & (g130) & (g180) & (g182) & (sk[8]) & (g183)));
	assign g235 = (((!g230) & (!g231) & (!sk[9]) & (g232) & (!g233) & (g234)) + ((!g230) & (!g231) & (!sk[9]) & (g232) & (g233) & (!g234)) + ((!g230) & (!g231) & (!sk[9]) & (g232) & (g233) & (g234)) + ((!g230) & (!g231) & (sk[9]) & (!g232) & (!g233) & (g234)) + ((!g230) & (g231) & (!sk[9]) & (!g232) & (!g233) & (!g234)) + ((!g230) & (g231) & (!sk[9]) & (!g232) & (!g233) & (g234)) + ((!g230) & (g231) & (!sk[9]) & (!g232) & (g233) & (!g234)) + ((!g230) & (g231) & (!sk[9]) & (!g232) & (g233) & (g234)) + ((!g230) & (g231) & (!sk[9]) & (g232) & (!g233) & (!g234)) + ((!g230) & (g231) & (!sk[9]) & (g232) & (!g233) & (g234)) + ((!g230) & (g231) & (!sk[9]) & (g232) & (g233) & (!g234)) + ((!g230) & (g231) & (!sk[9]) & (g232) & (g233) & (g234)) + ((g230) & (!g231) & (!sk[9]) & (g232) & (!g233) & (g234)) + ((g230) & (!g231) & (!sk[9]) & (g232) & (g233) & (!g234)) + ((g230) & (!g231) & (!sk[9]) & (g232) & (g233) & (g234)) + ((g230) & (g231) & (!sk[9]) & (!g232) & (!g233) & (!g234)) + ((g230) & (g231) & (!sk[9]) & (!g232) & (!g233) & (g234)) + ((g230) & (g231) & (!sk[9]) & (!g232) & (g233) & (!g234)) + ((g230) & (g231) & (!sk[9]) & (!g232) & (g233) & (g234)) + ((g230) & (g231) & (!sk[9]) & (g232) & (!g233) & (!g234)) + ((g230) & (g231) & (!sk[9]) & (g232) & (!g233) & (g234)) + ((g230) & (g231) & (!sk[9]) & (g232) & (g233) & (!g234)) + ((g230) & (g231) & (!sk[9]) & (g232) & (g233) & (g234)));
	assign g236 = (((g102) & (!sk[10]) & (!g212)) + ((g102) & (!sk[10]) & (g212)) + ((g102) & (sk[10]) & (g212)));
	assign g237 = (((!g102) & (!g182) & (!sk[11]) & (g183)) + ((!g102) & (g182) & (!sk[11]) & (!g183)) + ((!g102) & (g182) & (!sk[11]) & (g183)) + ((g102) & (!g182) & (!sk[11]) & (g183)) + ((g102) & (!g182) & (sk[11]) & (g183)) + ((g102) & (g182) & (!sk[11]) & (!g183)) + ((g102) & (g182) & (!sk[11]) & (g183)) + ((g102) & (g182) & (sk[11]) & (!g183)) + ((g102) & (g182) & (sk[11]) & (g183)));
	assign g238 = (((!sk[12]) & (!g102) & (!g175) & (g177)) + ((!sk[12]) & (!g102) & (g175) & (!g177)) + ((!sk[12]) & (!g102) & (g175) & (g177)) + ((!sk[12]) & (g102) & (!g175) & (g177)) + ((!sk[12]) & (g102) & (g175) & (!g177)) + ((!sk[12]) & (g102) & (g175) & (g177)) + ((sk[12]) & (g102) & (!g175) & (g177)) + ((sk[12]) & (g102) & (g175) & (!g177)) + ((sk[12]) & (g102) & (g175) & (g177)));
	assign g239 = (((!sk[13]) & (!g130) & (!g185) & (g212)) + ((!sk[13]) & (!g130) & (g185) & (!g212)) + ((!sk[13]) & (!g130) & (g185) & (g212)) + ((!sk[13]) & (g130) & (!g185) & (g212)) + ((!sk[13]) & (g130) & (g185) & (!g212)) + ((!sk[13]) & (g130) & (g185) & (g212)) + ((sk[13]) & (!g130) & (!g185) & (g212)) + ((sk[13]) & (!g130) & (g185) & (!g212)) + ((sk[13]) & (!g130) & (g185) & (g212)));
	assign g240 = (((!sk[14]) & (!g102) & (!g105) & (g183) & (!g192)) + ((!sk[14]) & (!g102) & (!g105) & (g183) & (g192)) + ((!sk[14]) & (!g102) & (g105) & (g183) & (!g192)) + ((!sk[14]) & (!g102) & (g105) & (g183) & (g192)) + ((!sk[14]) & (g102) & (!g105) & (g183) & (!g192)) + ((!sk[14]) & (g102) & (!g105) & (g183) & (g192)) + ((!sk[14]) & (g102) & (g105) & (g183) & (!g192)) + ((!sk[14]) & (g102) & (g105) & (g183) & (g192)) + ((sk[14]) & (!g102) & (!g105) & (!g183) & (!g192)) + ((sk[14]) & (!g102) & (g105) & (!g183) & (!g192)) + ((sk[14]) & (!g102) & (g105) & (!g183) & (g192)) + ((sk[14]) & (!g102) & (g105) & (g183) & (!g192)) + ((sk[14]) & (!g102) & (g105) & (g183) & (g192)) + ((sk[14]) & (g102) & (!g105) & (!g183) & (!g192)) + ((sk[14]) & (g102) & (g105) & (!g183) & (!g192)) + ((sk[14]) & (g102) & (g105) & (g183) & (!g192)));
	assign g241 = (((!g102) & (!g191) & (g180) & (!sk[15]) & (!g200)) + ((!g102) & (!g191) & (g180) & (!sk[15]) & (g200)) + ((!g102) & (g191) & (g180) & (!sk[15]) & (!g200)) + ((!g102) & (g191) & (g180) & (!sk[15]) & (g200)) + ((g102) & (!g191) & (!g180) & (sk[15]) & (g200)) + ((g102) & (!g191) & (g180) & (!sk[15]) & (!g200)) + ((g102) & (!g191) & (g180) & (!sk[15]) & (g200)) + ((g102) & (!g191) & (g180) & (sk[15]) & (!g200)) + ((g102) & (!g191) & (g180) & (sk[15]) & (g200)) + ((g102) & (g191) & (!g180) & (sk[15]) & (!g200)) + ((g102) & (g191) & (!g180) & (sk[15]) & (g200)) + ((g102) & (g191) & (g180) & (!sk[15]) & (!g200)) + ((g102) & (g191) & (g180) & (!sk[15]) & (g200)) + ((g102) & (g191) & (g180) & (sk[15]) & (!g200)) + ((g102) & (g191) & (g180) & (sk[15]) & (g200)));
	assign g242 = (((!g236) & (!g237) & (!g238) & (!g239) & (g240) & (!g241)));
	assign g243 = (((!sk[17]) & (!g130) & (!g191) & (g187)) + ((!sk[17]) & (!g130) & (g191) & (!g187)) + ((!sk[17]) & (!g130) & (g191) & (g187)) + ((!sk[17]) & (g130) & (!g191) & (g187)) + ((!sk[17]) & (g130) & (g191) & (!g187)) + ((!sk[17]) & (g130) & (g191) & (g187)) + ((sk[17]) & (!g130) & (!g191) & (g187)) + ((sk[17]) & (!g130) & (g191) & (!g187)) + ((sk[17]) & (!g130) & (g191) & (g187)));
	assign g244 = (((!sk[18]) & (!g130) & (!g186) & (g192)) + ((!sk[18]) & (!g130) & (g186) & (!g192)) + ((!sk[18]) & (!g130) & (g186) & (g192)) + ((!sk[18]) & (g130) & (!g186) & (g192)) + ((!sk[18]) & (g130) & (g186) & (!g192)) + ((!sk[18]) & (g130) & (g186) & (g192)) + ((sk[18]) & (!g130) & (!g186) & (g192)) + ((sk[18]) & (!g130) & (g186) & (!g192)) + ((sk[18]) & (!g130) & (g186) & (g192)));
	assign g245 = (((!g123) & (!sk[19]) & (!g175) & (g177)) + ((!g123) & (!sk[19]) & (g175) & (!g177)) + ((!g123) & (!sk[19]) & (g175) & (g177)) + ((!g123) & (sk[19]) & (!g175) & (g177)) + ((!g123) & (sk[19]) & (g175) & (!g177)) + ((!g123) & (sk[19]) & (g175) & (g177)) + ((g123) & (!sk[19]) & (!g175) & (g177)) + ((g123) & (!sk[19]) & (g175) & (!g177)) + ((g123) & (!sk[19]) & (g175) & (g177)));
	assign g246 = (((!i_8_) & (!g73) & (g200) & (!sk[20]) & (!g212)) + ((!i_8_) & (!g73) & (g200) & (!sk[20]) & (g212)) + ((!i_8_) & (g73) & (!g200) & (sk[20]) & (g212)) + ((!i_8_) & (g73) & (g200) & (!sk[20]) & (!g212)) + ((!i_8_) & (g73) & (g200) & (!sk[20]) & (g212)) + ((!i_8_) & (g73) & (g200) & (sk[20]) & (!g212)) + ((!i_8_) & (g73) & (g200) & (sk[20]) & (g212)) + ((i_8_) & (!g73) & (g200) & (!sk[20]) & (!g212)) + ((i_8_) & (!g73) & (g200) & (!sk[20]) & (g212)) + ((i_8_) & (g73) & (g200) & (!sk[20]) & (!g212)) + ((i_8_) & (g73) & (g200) & (!sk[20]) & (g212)) + ((i_8_) & (g73) & (g200) & (sk[20]) & (!g212)) + ((i_8_) & (g73) & (g200) & (sk[20]) & (g212)));
	assign g247 = (((!i_8_) & (!g73) & (!g135) & (!g131) & (!g185) & (!g197)) + ((!i_8_) & (!g73) & (!g135) & (g131) & (!g185) & (!g197)) + ((!i_8_) & (!g73) & (!g135) & (g131) & (!g185) & (g197)) + ((!i_8_) & (!g73) & (g135) & (!g131) & (!g185) & (!g197)) + ((!i_8_) & (!g73) & (g135) & (g131) & (!g185) & (!g197)) + ((!i_8_) & (!g73) & (g135) & (g131) & (!g185) & (g197)) + ((!i_8_) & (!g73) & (g135) & (g131) & (g185) & (!g197)) + ((!i_8_) & (!g73) & (g135) & (g131) & (g185) & (g197)) + ((!i_8_) & (g73) & (!g135) & (!g131) & (!g185) & (!g197)) + ((!i_8_) & (g73) & (!g135) & (g131) & (!g185) & (!g197)) + ((!i_8_) & (g73) & (!g135) & (g131) & (!g185) & (g197)) + ((!i_8_) & (g73) & (g135) & (!g131) & (!g185) & (!g197)) + ((!i_8_) & (g73) & (g135) & (g131) & (!g185) & (!g197)) + ((!i_8_) & (g73) & (g135) & (g131) & (!g185) & (g197)) + ((i_8_) & (!g73) & (!g135) & (!g131) & (!g185) & (!g197)) + ((i_8_) & (!g73) & (!g135) & (g131) & (!g185) & (!g197)) + ((i_8_) & (!g73) & (!g135) & (g131) & (!g185) & (g197)) + ((i_8_) & (!g73) & (g135) & (!g131) & (!g185) & (!g197)) + ((i_8_) & (!g73) & (g135) & (g131) & (!g185) & (!g197)) + ((i_8_) & (!g73) & (g135) & (g131) & (!g185) & (g197)) + ((i_8_) & (!g73) & (g135) & (g131) & (g185) & (!g197)) + ((i_8_) & (!g73) & (g135) & (g131) & (g185) & (g197)) + ((i_8_) & (g73) & (!g135) & (!g131) & (!g185) & (!g197)) + ((i_8_) & (g73) & (!g135) & (g131) & (!g185) & (!g197)) + ((i_8_) & (g73) & (!g135) & (g131) & (!g185) & (g197)) + ((i_8_) & (g73) & (g135) & (!g131) & (!g185) & (!g197)) + ((i_8_) & (g73) & (g135) & (g131) & (!g185) & (!g197)) + ((i_8_) & (g73) & (g135) & (g131) & (!g185) & (g197)) + ((i_8_) & (g73) & (g135) & (g131) & (g185) & (!g197)) + ((i_8_) & (g73) & (g135) & (g131) & (g185) & (g197)));
	assign g248 = (((!g243) & (!g244) & (!g245) & (!g246) & (sk[22]) & (g247)) + ((!g243) & (!g244) & (g245) & (!g246) & (!sk[22]) & (g247)) + ((!g243) & (!g244) & (g245) & (g246) & (!sk[22]) & (!g247)) + ((!g243) & (!g244) & (g245) & (g246) & (!sk[22]) & (g247)) + ((!g243) & (g244) & (!g245) & (!g246) & (!sk[22]) & (!g247)) + ((!g243) & (g244) & (!g245) & (!g246) & (!sk[22]) & (g247)) + ((!g243) & (g244) & (!g245) & (g246) & (!sk[22]) & (!g247)) + ((!g243) & (g244) & (!g245) & (g246) & (!sk[22]) & (g247)) + ((!g243) & (g244) & (g245) & (!g246) & (!sk[22]) & (!g247)) + ((!g243) & (g244) & (g245) & (!g246) & (!sk[22]) & (g247)) + ((!g243) & (g244) & (g245) & (g246) & (!sk[22]) & (!g247)) + ((!g243) & (g244) & (g245) & (g246) & (!sk[22]) & (g247)) + ((g243) & (!g244) & (g245) & (!g246) & (!sk[22]) & (g247)) + ((g243) & (!g244) & (g245) & (g246) & (!sk[22]) & (!g247)) + ((g243) & (!g244) & (g245) & (g246) & (!sk[22]) & (g247)) + ((g243) & (g244) & (!g245) & (!g246) & (!sk[22]) & (!g247)) + ((g243) & (g244) & (!g245) & (!g246) & (!sk[22]) & (g247)) + ((g243) & (g244) & (!g245) & (g246) & (!sk[22]) & (!g247)) + ((g243) & (g244) & (!g245) & (g246) & (!sk[22]) & (g247)) + ((g243) & (g244) & (g245) & (!g246) & (!sk[22]) & (!g247)) + ((g243) & (g244) & (g245) & (!g246) & (!sk[22]) & (g247)) + ((g243) & (g244) & (g245) & (g246) & (!sk[22]) & (!g247)) + ((g243) & (g244) & (g245) & (g246) & (!sk[22]) & (g247)));
	assign g249 = (((!i_9_) & (!i_11_) & (!sk[23]) & (i_15_) & (!g174)) + ((!i_9_) & (!i_11_) & (!sk[23]) & (i_15_) & (g174)) + ((!i_9_) & (!i_11_) & (sk[23]) & (!i_15_) & (!g174)) + ((!i_9_) & (i_11_) & (!sk[23]) & (i_15_) & (!g174)) + ((!i_9_) & (i_11_) & (!sk[23]) & (i_15_) & (g174)) + ((i_9_) & (!i_11_) & (!sk[23]) & (i_15_) & (!g174)) + ((i_9_) & (!i_11_) & (!sk[23]) & (i_15_) & (g174)) + ((i_9_) & (i_11_) & (!sk[23]) & (i_15_) & (!g174)) + ((i_9_) & (i_11_) & (!sk[23]) & (i_15_) & (g174)));
	assign g250 = (((!g161) & (!g157) & (!g186) & (!g187) & (!g182) & (!g192)) + ((!g161) & (!g157) & (!g186) & (!g187) & (!g182) & (g192)) + ((!g161) & (!g157) & (!g186) & (!g187) & (g182) & (!g192)) + ((!g161) & (!g157) & (!g186) & (!g187) & (g182) & (g192)) + ((!g161) & (!g157) & (!g186) & (g187) & (!g182) & (!g192)) + ((!g161) & (!g157) & (!g186) & (g187) & (!g182) & (g192)) + ((!g161) & (!g157) & (!g186) & (g187) & (g182) & (!g192)) + ((!g161) & (!g157) & (!g186) & (g187) & (g182) & (g192)) + ((!g161) & (!g157) & (g186) & (!g187) & (!g182) & (!g192)) + ((!g161) & (!g157) & (g186) & (!g187) & (!g182) & (g192)) + ((!g161) & (!g157) & (g186) & (!g187) & (g182) & (!g192)) + ((!g161) & (!g157) & (g186) & (!g187) & (g182) & (g192)) + ((!g161) & (!g157) & (g186) & (g187) & (!g182) & (!g192)) + ((!g161) & (!g157) & (g186) & (g187) & (!g182) & (g192)) + ((!g161) & (!g157) & (g186) & (g187) & (g182) & (!g192)) + ((!g161) & (!g157) & (g186) & (g187) & (g182) & (g192)) + ((!g161) & (g157) & (!g186) & (!g187) & (!g182) & (!g192)) + ((!g161) & (g157) & (!g186) & (!g187) & (!g182) & (g192)) + ((!g161) & (g157) & (!g186) & (!g187) & (g182) & (!g192)) + ((!g161) & (g157) & (!g186) & (!g187) & (g182) & (g192)) + ((!g161) & (g157) & (g186) & (!g187) & (!g182) & (!g192)) + ((!g161) & (g157) & (g186) & (!g187) & (!g182) & (g192)) + ((!g161) & (g157) & (g186) & (!g187) & (g182) & (!g192)) + ((!g161) & (g157) & (g186) & (!g187) & (g182) & (g192)) + ((g161) & (!g157) & (!g186) & (!g187) & (!g182) & (!g192)) + ((g161) & (!g157) & (!g186) & (g187) & (!g182) & (!g192)) + ((g161) & (g157) & (!g186) & (!g187) & (!g182) & (!g192)));
	assign g251 = (((!g102) & (!g130) & (!g188) & (!g175) & (!g249) & (g250)) + ((!g102) & (!g130) & (!g188) & (!g175) & (g249) & (g250)) + ((!g102) & (!g130) & (!g188) & (g175) & (!g249) & (g250)) + ((!g102) & (!g130) & (g188) & (!g175) & (!g249) & (g250)) + ((!g102) & (!g130) & (g188) & (!g175) & (g249) & (g250)) + ((!g102) & (!g130) & (g188) & (g175) & (!g249) & (g250)) + ((!g102) & (g130) & (!g188) & (!g175) & (!g249) & (g250)) + ((!g102) & (g130) & (!g188) & (!g175) & (g249) & (g250)) + ((!g102) & (g130) & (!g188) & (g175) & (!g249) & (g250)) + ((!g102) & (g130) & (!g188) & (g175) & (g249) & (g250)) + ((!g102) & (g130) & (g188) & (!g175) & (!g249) & (g250)) + ((!g102) & (g130) & (g188) & (!g175) & (g249) & (g250)) + ((!g102) & (g130) & (g188) & (g175) & (!g249) & (g250)) + ((!g102) & (g130) & (g188) & (g175) & (g249) & (g250)) + ((g102) & (!g130) & (!g188) & (!g175) & (!g249) & (g250)) + ((g102) & (!g130) & (!g188) & (g175) & (!g249) & (g250)) + ((g102) & (!g130) & (g188) & (!g175) & (!g249) & (g250)) + ((g102) & (!g130) & (g188) & (g175) & (!g249) & (g250)) + ((g102) & (g130) & (!g188) & (!g175) & (!g249) & (g250)) + ((g102) & (g130) & (!g188) & (!g175) & (g249) & (g250)) + ((g102) & (g130) & (!g188) & (g175) & (!g249) & (g250)) + ((g102) & (g130) & (!g188) & (g175) & (g249) & (g250)) + ((g102) & (g130) & (g188) & (!g175) & (!g249) & (g250)) + ((g102) & (g130) & (g188) & (g175) & (!g249) & (g250)));
	assign g252 = (((!g220) & (g229) & (g235) & (g242) & (g248) & (g251)));
	assign g253 = (((!sk[27]) & (g2) & (!g120)) + ((!sk[27]) & (g2) & (g120)) + ((sk[27]) & (!g2) & (!g120)) + ((sk[27]) & (!g2) & (g120)) + ((sk[27]) & (g2) & (!g120)));
	assign g254 = (((!sk[28]) & (g30) & (!g166)) + ((!sk[28]) & (g30) & (g166)) + ((sk[28]) & (!g30) & (!g166)) + ((sk[28]) & (!g30) & (g166)) + ((sk[28]) & (g30) & (!g166)));
	assign g255 = (((!sk[29]) & (!g157) & (!g165) & (g182) & (!g253) & (g254)) + ((!sk[29]) & (!g157) & (!g165) & (g182) & (g253) & (!g254)) + ((!sk[29]) & (!g157) & (!g165) & (g182) & (g253) & (g254)) + ((!sk[29]) & (!g157) & (g165) & (!g182) & (!g253) & (!g254)) + ((!sk[29]) & (!g157) & (g165) & (!g182) & (!g253) & (g254)) + ((!sk[29]) & (!g157) & (g165) & (!g182) & (g253) & (!g254)) + ((!sk[29]) & (!g157) & (g165) & (!g182) & (g253) & (g254)) + ((!sk[29]) & (!g157) & (g165) & (g182) & (!g253) & (!g254)) + ((!sk[29]) & (!g157) & (g165) & (g182) & (!g253) & (g254)) + ((!sk[29]) & (!g157) & (g165) & (g182) & (g253) & (!g254)) + ((!sk[29]) & (!g157) & (g165) & (g182) & (g253) & (g254)) + ((!sk[29]) & (g157) & (!g165) & (g182) & (!g253) & (g254)) + ((!sk[29]) & (g157) & (!g165) & (g182) & (g253) & (!g254)) + ((!sk[29]) & (g157) & (!g165) & (g182) & (g253) & (g254)) + ((!sk[29]) & (g157) & (g165) & (!g182) & (!g253) & (!g254)) + ((!sk[29]) & (g157) & (g165) & (!g182) & (!g253) & (g254)) + ((!sk[29]) & (g157) & (g165) & (!g182) & (g253) & (!g254)) + ((!sk[29]) & (g157) & (g165) & (!g182) & (g253) & (g254)) + ((!sk[29]) & (g157) & (g165) & (g182) & (!g253) & (!g254)) + ((!sk[29]) & (g157) & (g165) & (g182) & (!g253) & (g254)) + ((!sk[29]) & (g157) & (g165) & (g182) & (g253) & (!g254)) + ((!sk[29]) & (g157) & (g165) & (g182) & (g253) & (g254)) + ((sk[29]) & (!g157) & (!g165) & (g182) & (!g253) & (!g254)) + ((sk[29]) & (!g157) & (!g165) & (g182) & (!g253) & (g254)) + ((sk[29]) & (!g157) & (!g165) & (g182) & (g253) & (!g254)) + ((sk[29]) & (!g157) & (g165) & (g182) & (!g253) & (!g254)) + ((sk[29]) & (!g157) & (g165) & (g182) & (!g253) & (g254)) + ((sk[29]) & (!g157) & (g165) & (g182) & (g253) & (!g254)) + ((sk[29]) & (!g157) & (g165) & (g182) & (g253) & (g254)) + ((sk[29]) & (g157) & (!g165) & (g182) & (!g253) & (!g254)) + ((sk[29]) & (g157) & (!g165) & (g182) & (!g253) & (g254)) + ((sk[29]) & (g157) & (!g165) & (g182) & (g253) & (!g254)) + ((sk[29]) & (g157) & (!g165) & (g182) & (g253) & (g254)) + ((sk[29]) & (g157) & (g165) & (g182) & (!g253) & (!g254)) + ((sk[29]) & (g157) & (g165) & (g182) & (!g253) & (g254)) + ((sk[29]) & (g157) & (g165) & (g182) & (g253) & (!g254)) + ((sk[29]) & (g157) & (g165) & (g182) & (g253) & (g254)));
	assign g256 = (((g80) & (!i_11_) & (!i_15_) & (!g157) & (g121) & (!g174)) + ((g80) & (!i_11_) & (!i_15_) & (g157) & (g121) & (!g174)) + ((g80) & (i_11_) & (!i_15_) & (g157) & (!g121) & (!g174)) + ((g80) & (i_11_) & (!i_15_) & (g157) & (g121) & (!g174)));
	assign g257 = (((!sk[31]) & (g2) & (!g166)) + ((!sk[31]) & (g2) & (g166)) + ((sk[31]) & (g2) & (g166)));
	assign g258 = (((!sk[32]) & (!i_8_) & (!g73) & (g135) & (!g257)) + ((!sk[32]) & (!i_8_) & (!g73) & (g135) & (g257)) + ((!sk[32]) & (!i_8_) & (g73) & (g135) & (!g257)) + ((!sk[32]) & (!i_8_) & (g73) & (g135) & (g257)) + ((!sk[32]) & (i_8_) & (!g73) & (g135) & (!g257)) + ((!sk[32]) & (i_8_) & (!g73) & (g135) & (g257)) + ((!sk[32]) & (i_8_) & (g73) & (g135) & (!g257)) + ((!sk[32]) & (i_8_) & (g73) & (g135) & (g257)) + ((sk[32]) & (!i_8_) & (!g73) & (g135) & (!g257)) + ((sk[32]) & (i_8_) & (!g73) & (g135) & (!g257)) + ((sk[32]) & (i_8_) & (g73) & (g135) & (!g257)));
	assign g259 = (((!g164) & (sk[33]) & (!g217)) + ((g164) & (!sk[33]) & (!g217)) + ((g164) & (!sk[33]) & (g217)));
	assign g260 = (((!i_9_) & (!sk[34]) & (!i_11_) & (i_15_) & (!g176)) + ((!i_9_) & (!sk[34]) & (!i_11_) & (i_15_) & (g176)) + ((!i_9_) & (!sk[34]) & (i_11_) & (i_15_) & (!g176)) + ((!i_9_) & (!sk[34]) & (i_11_) & (i_15_) & (g176)) + ((!i_9_) & (sk[34]) & (!i_11_) & (i_15_) & (!g176)) + ((i_9_) & (!sk[34]) & (!i_11_) & (i_15_) & (!g176)) + ((i_9_) & (!sk[34]) & (!i_11_) & (i_15_) & (g176)) + ((i_9_) & (!sk[34]) & (i_11_) & (i_15_) & (!g176)) + ((i_9_) & (!sk[34]) & (i_11_) & (i_15_) & (g176)));
	assign g261 = (((!g74) & (!g194) & (!g258) & (!g177) & (!g259) & (g260)) + ((!g74) & (!g194) & (!g258) & (g177) & (!g259) & (g260)) + ((!g74) & (!g194) & (!g258) & (g177) & (g259) & (g260)) + ((!g74) & (g194) & (!g258) & (!g177) & (!g259) & (g260)) + ((!g74) & (g194) & (!g258) & (g177) & (!g259) & (g260)) + ((!g74) & (g194) & (!g258) & (g177) & (g259) & (g260)) + ((!g74) & (g194) & (g258) & (!g177) & (!g259) & (g260)) + ((!g74) & (g194) & (g258) & (g177) & (!g259) & (g260)) + ((g74) & (!g194) & (!g258) & (!g177) & (!g259) & (g260)) + ((g74) & (!g194) & (!g258) & (!g177) & (g259) & (g260)) + ((g74) & (!g194) & (!g258) & (g177) & (!g259) & (g260)) + ((g74) & (!g194) & (!g258) & (g177) & (g259) & (g260)) + ((g74) & (g194) & (!g258) & (!g177) & (!g259) & (g260)) + ((g74) & (g194) & (!g258) & (!g177) & (g259) & (g260)) + ((g74) & (g194) & (!g258) & (g177) & (!g259) & (g260)) + ((g74) & (g194) & (!g258) & (g177) & (g259) & (g260)) + ((g74) & (g194) & (g258) & (!g177) & (!g259) & (g260)) + ((g74) & (g194) & (g258) & (g177) & (!g259) & (g260)));
	assign g262 = (((!i_8_) & (!sk[36]) & (!i_6_) & (i_7_) & (!g120)) + ((!i_8_) & (!sk[36]) & (!i_6_) & (i_7_) & (g120)) + ((!i_8_) & (!sk[36]) & (i_6_) & (i_7_) & (!g120)) + ((!i_8_) & (!sk[36]) & (i_6_) & (i_7_) & (g120)) + ((!i_8_) & (sk[36]) & (!i_6_) & (!i_7_) & (g120)) + ((i_8_) & (!sk[36]) & (!i_6_) & (i_7_) & (!g120)) + ((i_8_) & (!sk[36]) & (!i_6_) & (i_7_) & (g120)) + ((i_8_) & (!sk[36]) & (i_6_) & (i_7_) & (!g120)) + ((i_8_) & (!sk[36]) & (i_6_) & (i_7_) & (g120)) + ((i_8_) & (sk[36]) & (!i_6_) & (i_7_) & (g120)));
	assign g263 = (((!g159) & (!g185) & (!g262) & (sk[37]) & (g191)) + ((!g159) & (!g185) & (g262) & (!sk[37]) & (!g191)) + ((!g159) & (!g185) & (g262) & (!sk[37]) & (g191)) + ((!g159) & (!g185) & (g262) & (sk[37]) & (g191)) + ((!g159) & (g185) & (!g262) & (sk[37]) & (g191)) + ((!g159) & (g185) & (g262) & (!sk[37]) & (!g191)) + ((!g159) & (g185) & (g262) & (!sk[37]) & (g191)) + ((!g159) & (g185) & (g262) & (sk[37]) & (!g191)) + ((!g159) & (g185) & (g262) & (sk[37]) & (g191)) + ((g159) & (!g185) & (g262) & (!sk[37]) & (!g191)) + ((g159) & (!g185) & (g262) & (!sk[37]) & (g191)) + ((g159) & (g185) & (g262) & (!sk[37]) & (!g191)) + ((g159) & (g185) & (g262) & (!sk[37]) & (g191)) + ((g159) & (g185) & (g262) & (sk[37]) & (!g191)) + ((g159) & (g185) & (g262) & (sk[37]) & (g191)));
	assign g264 = (((!g165) & (!g154) & (!sk[38]) & (g192) & (!g263)) + ((!g165) & (!g154) & (!sk[38]) & (g192) & (g263)) + ((!g165) & (!g154) & (sk[38]) & (!g192) & (!g263)) + ((!g165) & (g154) & (!sk[38]) & (g192) & (!g263)) + ((!g165) & (g154) & (!sk[38]) & (g192) & (g263)) + ((!g165) & (g154) & (sk[38]) & (!g192) & (!g263)) + ((!g165) & (g154) & (sk[38]) & (g192) & (!g263)) + ((g165) & (!g154) & (!sk[38]) & (g192) & (!g263)) + ((g165) & (!g154) & (!sk[38]) & (g192) & (g263)) + ((g165) & (!g154) & (sk[38]) & (!g192) & (!g263)) + ((g165) & (g154) & (!sk[38]) & (g192) & (!g263)) + ((g165) & (g154) & (!sk[38]) & (g192) & (g263)) + ((g165) & (g154) & (sk[38]) & (!g192) & (!g263)));
	assign g265 = (((!sk[39]) & (!g144) & (!g130) & (g200)) + ((!sk[39]) & (!g144) & (g130) & (!g200)) + ((!sk[39]) & (!g144) & (g130) & (g200)) + ((!sk[39]) & (g144) & (!g130) & (g200)) + ((!sk[39]) & (g144) & (g130) & (!g200)) + ((!sk[39]) & (g144) & (g130) & (g200)) + ((sk[39]) & (!g144) & (!g130) & (!g200)) + ((sk[39]) & (!g144) & (g130) & (!g200)) + ((sk[39]) & (!g144) & (g130) & (g200)));
	assign g266 = (((!i_9_) & (i_10_) & (i_11_) & (!i_15_) & (!g130) & (!g174)) + ((i_9_) & (!i_10_) & (!i_11_) & (!i_15_) & (!g130) & (!g174)) + ((i_9_) & (!i_10_) & (!i_11_) & (!i_15_) & (g130) & (!g174)));
	assign g267 = (((!g159) & (!sk[41]) & (!g197) & (g258) & (!g265) & (g266)) + ((!g159) & (!sk[41]) & (!g197) & (g258) & (g265) & (!g266)) + ((!g159) & (!sk[41]) & (!g197) & (g258) & (g265) & (g266)) + ((!g159) & (!sk[41]) & (g197) & (!g258) & (!g265) & (!g266)) + ((!g159) & (!sk[41]) & (g197) & (!g258) & (!g265) & (g266)) + ((!g159) & (!sk[41]) & (g197) & (!g258) & (g265) & (!g266)) + ((!g159) & (!sk[41]) & (g197) & (!g258) & (g265) & (g266)) + ((!g159) & (!sk[41]) & (g197) & (g258) & (!g265) & (!g266)) + ((!g159) & (!sk[41]) & (g197) & (g258) & (!g265) & (g266)) + ((!g159) & (!sk[41]) & (g197) & (g258) & (g265) & (!g266)) + ((!g159) & (!sk[41]) & (g197) & (g258) & (g265) & (g266)) + ((!g159) & (sk[41]) & (!g197) & (!g258) & (!g265) & (!g266)) + ((!g159) & (sk[41]) & (!g197) & (!g258) & (g265) & (!g266)) + ((!g159) & (sk[41]) & (!g197) & (!g258) & (g265) & (g266)) + ((!g159) & (sk[41]) & (!g197) & (g258) & (!g265) & (!g266)) + ((!g159) & (sk[41]) & (!g197) & (g258) & (g265) & (!g266)) + ((!g159) & (sk[41]) & (!g197) & (g258) & (g265) & (g266)) + ((g159) & (!sk[41]) & (!g197) & (g258) & (!g265) & (g266)) + ((g159) & (!sk[41]) & (!g197) & (g258) & (g265) & (!g266)) + ((g159) & (!sk[41]) & (!g197) & (g258) & (g265) & (g266)) + ((g159) & (!sk[41]) & (g197) & (!g258) & (!g265) & (!g266)) + ((g159) & (!sk[41]) & (g197) & (!g258) & (!g265) & (g266)) + ((g159) & (!sk[41]) & (g197) & (!g258) & (g265) & (!g266)) + ((g159) & (!sk[41]) & (g197) & (!g258) & (g265) & (g266)) + ((g159) & (!sk[41]) & (g197) & (g258) & (!g265) & (!g266)) + ((g159) & (!sk[41]) & (g197) & (g258) & (!g265) & (g266)) + ((g159) & (!sk[41]) & (g197) & (g258) & (g265) & (!g266)) + ((g159) & (!sk[41]) & (g197) & (g258) & (g265) & (g266)) + ((g159) & (sk[41]) & (!g197) & (!g258) & (!g265) & (!g266)) + ((g159) & (sk[41]) & (!g197) & (!g258) & (g265) & (!g266)) + ((g159) & (sk[41]) & (!g197) & (!g258) & (g265) & (g266)) + ((g159) & (sk[41]) & (!g197) & (g258) & (!g265) & (!g266)) + ((g159) & (sk[41]) & (!g197) & (g258) & (g265) & (!g266)) + ((g159) & (sk[41]) & (!g197) & (g258) & (g265) & (g266)) + ((g159) & (sk[41]) & (g197) & (g258) & (!g265) & (!g266)) + ((g159) & (sk[41]) & (g197) & (g258) & (g265) & (!g266)) + ((g159) & (sk[41]) & (g197) & (g258) & (g265) & (g266)));
	assign g268 = (((!g255) & (!g256) & (!g261) & (g264) & (sk[42]) & (g267)) + ((!g255) & (!g256) & (g261) & (!g264) & (!sk[42]) & (g267)) + ((!g255) & (!g256) & (g261) & (g264) & (!sk[42]) & (!g267)) + ((!g255) & (!g256) & (g261) & (g264) & (!sk[42]) & (g267)) + ((!g255) & (g256) & (!g261) & (!g264) & (!sk[42]) & (!g267)) + ((!g255) & (g256) & (!g261) & (!g264) & (!sk[42]) & (g267)) + ((!g255) & (g256) & (!g261) & (g264) & (!sk[42]) & (!g267)) + ((!g255) & (g256) & (!g261) & (g264) & (!sk[42]) & (g267)) + ((!g255) & (g256) & (g261) & (!g264) & (!sk[42]) & (!g267)) + ((!g255) & (g256) & (g261) & (!g264) & (!sk[42]) & (g267)) + ((!g255) & (g256) & (g261) & (g264) & (!sk[42]) & (!g267)) + ((!g255) & (g256) & (g261) & (g264) & (!sk[42]) & (g267)) + ((g255) & (!g256) & (g261) & (!g264) & (!sk[42]) & (g267)) + ((g255) & (!g256) & (g261) & (g264) & (!sk[42]) & (!g267)) + ((g255) & (!g256) & (g261) & (g264) & (!sk[42]) & (g267)) + ((g255) & (g256) & (!g261) & (!g264) & (!sk[42]) & (!g267)) + ((g255) & (g256) & (!g261) & (!g264) & (!sk[42]) & (g267)) + ((g255) & (g256) & (!g261) & (g264) & (!sk[42]) & (!g267)) + ((g255) & (g256) & (!g261) & (g264) & (!sk[42]) & (g267)) + ((g255) & (g256) & (g261) & (!g264) & (!sk[42]) & (!g267)) + ((g255) & (g256) & (g261) & (!g264) & (!sk[42]) & (g267)) + ((g255) & (g256) & (g261) & (g264) & (!sk[42]) & (!g267)) + ((g255) & (g256) & (g261) & (g264) & (!sk[42]) & (g267)));
	assign g269 = (((g196) & (g203) & (g211) & (g216) & (g252) & (g268)));
	assign g270 = (((!sk[44]) & (g3) & (!g24)) + ((!sk[44]) & (g3) & (g24)) + ((sk[44]) & (g3) & (!g24)));
	assign g271 = (((!i_9_) & (!i_10_) & (!i_11_) & (!i_15_) & (!g68) & (g74)) + ((!i_9_) & (!i_10_) & (i_11_) & (!i_15_) & (!g68) & (g74)) + ((!i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (!g68) & (g74)) + ((i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (!g68) & (g74)) + ((i_9_) & (i_10_) & (i_11_) & (!i_15_) & (!g68) & (g74)));
	assign g272 = (((!sk[46]) & (g24) & (!g86)) + ((!sk[46]) & (g24) & (g86)) + ((sk[46]) & (!g24) & (g86)));
	assign g273 = (((!g68) & (sk[47]) & (g86)) + ((g68) & (!sk[47]) & (!g86)) + ((g68) & (!sk[47]) & (g86)));
	assign g274 = (((!i_8_) & (!sk[48]) & (!g73) & (g272) & (!g273)) + ((!i_8_) & (!sk[48]) & (!g73) & (g272) & (g273)) + ((!i_8_) & (!sk[48]) & (g73) & (g272) & (!g273)) + ((!i_8_) & (!sk[48]) & (g73) & (g272) & (g273)) + ((!i_8_) & (sk[48]) & (g73) & (!g272) & (g273)) + ((!i_8_) & (sk[48]) & (g73) & (g272) & (!g273)) + ((!i_8_) & (sk[48]) & (g73) & (g272) & (g273)) + ((i_8_) & (!sk[48]) & (!g73) & (g272) & (!g273)) + ((i_8_) & (!sk[48]) & (!g73) & (g272) & (g273)) + ((i_8_) & (!sk[48]) & (g73) & (g272) & (!g273)) + ((i_8_) & (!sk[48]) & (g73) & (g272) & (g273)));
	assign g275 = (((!sk[49]) & (g27) & (!g68)) + ((!sk[49]) & (g27) & (g68)) + ((sk[49]) & (g27) & (!g68)));
	assign g276 = (((!i_8_) & (!sk[50]) & (!g28) & (g73) & (!g275)) + ((!i_8_) & (!sk[50]) & (!g28) & (g73) & (g275)) + ((!i_8_) & (!sk[50]) & (g28) & (g73) & (!g275)) + ((!i_8_) & (!sk[50]) & (g28) & (g73) & (g275)) + ((i_8_) & (!sk[50]) & (!g28) & (g73) & (!g275)) + ((i_8_) & (!sk[50]) & (!g28) & (g73) & (g275)) + ((i_8_) & (!sk[50]) & (g28) & (g73) & (!g275)) + ((i_8_) & (!sk[50]) & (g28) & (g73) & (g275)) + ((i_8_) & (sk[50]) & (!g28) & (g73) & (g275)) + ((i_8_) & (sk[50]) & (g28) & (g73) & (!g275)) + ((i_8_) & (sk[50]) & (g28) & (g73) & (g275)));
	assign g277 = (((!i_8_) & (!sk[51]) & (!g28) & (g73) & (!g275)) + ((!i_8_) & (!sk[51]) & (!g28) & (g73) & (g275)) + ((!i_8_) & (!sk[51]) & (g28) & (g73) & (!g275)) + ((!i_8_) & (!sk[51]) & (g28) & (g73) & (g275)) + ((!i_8_) & (sk[51]) & (!g28) & (g73) & (g275)) + ((!i_8_) & (sk[51]) & (g28) & (g73) & (!g275)) + ((!i_8_) & (sk[51]) & (g28) & (g73) & (g275)) + ((i_8_) & (!sk[51]) & (!g28) & (g73) & (!g275)) + ((i_8_) & (!sk[51]) & (!g28) & (g73) & (g275)) + ((i_8_) & (!sk[51]) & (g28) & (g73) & (!g275)) + ((i_8_) & (!sk[51]) & (g28) & (g73) & (g275)));
	assign g278 = (((!sk[52]) & (g20) & (!g68)) + ((!sk[52]) & (g20) & (g68)) + ((sk[52]) & (g20) & (!g68)));
	assign g279 = (((!i_8_) & (!g25) & (g73) & (!sk[53]) & (!g278)) + ((!i_8_) & (!g25) & (g73) & (!sk[53]) & (g278)) + ((!i_8_) & (!g25) & (g73) & (sk[53]) & (!g278)) + ((!i_8_) & (!g25) & (g73) & (sk[53]) & (g278)) + ((!i_8_) & (g25) & (g73) & (!sk[53]) & (!g278)) + ((!i_8_) & (g25) & (g73) & (!sk[53]) & (g278)) + ((i_8_) & (!g25) & (g73) & (!sk[53]) & (!g278)) + ((i_8_) & (!g25) & (g73) & (!sk[53]) & (g278)) + ((i_8_) & (!g25) & (g73) & (sk[53]) & (!g278)) + ((i_8_) & (!g25) & (g73) & (sk[53]) & (g278)) + ((i_8_) & (g25) & (g73) & (!sk[53]) & (!g278)) + ((i_8_) & (g25) & (g73) & (!sk[53]) & (g278)) + ((i_8_) & (g25) & (g73) & (sk[53]) & (g278)));
	assign g280 = (((!i_8_) & (!g24) & (!sk[54]) & (g73) & (!g68) & (g83)) + ((!i_8_) & (!g24) & (!sk[54]) & (g73) & (g68) & (!g83)) + ((!i_8_) & (!g24) & (!sk[54]) & (g73) & (g68) & (g83)) + ((!i_8_) & (!g24) & (sk[54]) & (g73) & (!g68) & (g83)) + ((!i_8_) & (!g24) & (sk[54]) & (g73) & (g68) & (g83)) + ((!i_8_) & (g24) & (!sk[54]) & (!g73) & (!g68) & (!g83)) + ((!i_8_) & (g24) & (!sk[54]) & (!g73) & (!g68) & (g83)) + ((!i_8_) & (g24) & (!sk[54]) & (!g73) & (g68) & (!g83)) + ((!i_8_) & (g24) & (!sk[54]) & (!g73) & (g68) & (g83)) + ((!i_8_) & (g24) & (!sk[54]) & (g73) & (!g68) & (!g83)) + ((!i_8_) & (g24) & (!sk[54]) & (g73) & (!g68) & (g83)) + ((!i_8_) & (g24) & (!sk[54]) & (g73) & (g68) & (!g83)) + ((!i_8_) & (g24) & (!sk[54]) & (g73) & (g68) & (g83)) + ((i_8_) & (!g24) & (!sk[54]) & (g73) & (!g68) & (g83)) + ((i_8_) & (!g24) & (!sk[54]) & (g73) & (g68) & (!g83)) + ((i_8_) & (!g24) & (!sk[54]) & (g73) & (g68) & (g83)) + ((i_8_) & (!g24) & (sk[54]) & (g73) & (!g68) & (g83)) + ((i_8_) & (!g24) & (sk[54]) & (g73) & (g68) & (g83)) + ((i_8_) & (g24) & (!sk[54]) & (!g73) & (!g68) & (!g83)) + ((i_8_) & (g24) & (!sk[54]) & (!g73) & (!g68) & (g83)) + ((i_8_) & (g24) & (!sk[54]) & (!g73) & (g68) & (!g83)) + ((i_8_) & (g24) & (!sk[54]) & (!g73) & (g68) & (g83)) + ((i_8_) & (g24) & (!sk[54]) & (g73) & (!g68) & (!g83)) + ((i_8_) & (g24) & (!sk[54]) & (g73) & (!g68) & (g83)) + ((i_8_) & (g24) & (!sk[54]) & (g73) & (g68) & (!g83)) + ((i_8_) & (g24) & (!sk[54]) & (g73) & (g68) & (g83)) + ((i_8_) & (g24) & (sk[54]) & (g73) & (!g68) & (g83)));
	assign g281 = (((g35) & (!sk[55]) & (!g68)) + ((g35) & (!sk[55]) & (g68)) + ((g35) & (sk[55]) & (!g68)));
	assign g282 = (((!sk[56]) & (g3) & (!g68)) + ((!sk[56]) & (g3) & (g68)) + ((sk[56]) & (g3) & (!g68)));
	assign g283 = (((i_8_) & (g73) & (!g273) & (!g281) & (!g282) & (g270)) + ((i_8_) & (g73) & (!g273) & (!g281) & (g282) & (!g270)) + ((i_8_) & (g73) & (!g273) & (!g281) & (g282) & (g270)) + ((i_8_) & (g73) & (!g273) & (g281) & (!g282) & (!g270)) + ((i_8_) & (g73) & (!g273) & (g281) & (!g282) & (g270)) + ((i_8_) & (g73) & (!g273) & (g281) & (g282) & (!g270)) + ((i_8_) & (g73) & (!g273) & (g281) & (g282) & (g270)) + ((i_8_) & (g73) & (g273) & (!g281) & (!g282) & (!g270)) + ((i_8_) & (g73) & (g273) & (!g281) & (!g282) & (g270)) + ((i_8_) & (g73) & (g273) & (!g281) & (g282) & (!g270)) + ((i_8_) & (g73) & (g273) & (!g281) & (g282) & (g270)) + ((i_8_) & (g73) & (g273) & (g281) & (!g282) & (!g270)) + ((i_8_) & (g73) & (g273) & (g281) & (!g282) & (g270)) + ((i_8_) & (g73) & (g273) & (g281) & (g282) & (!g270)) + ((i_8_) & (g73) & (g273) & (g281) & (g282) & (g270)));
	assign g284 = (((!g274) & (!g276) & (!g277) & (!g279) & (!g280) & (!g283)));
	assign g285 = (((!g74) & (!sk[59]) & (!g270) & (g271) & (!g284)) + ((!g74) & (!sk[59]) & (!g270) & (g271) & (g284)) + ((!g74) & (!sk[59]) & (g270) & (g271) & (!g284)) + ((!g74) & (!sk[59]) & (g270) & (g271) & (g284)) + ((!g74) & (sk[59]) & (!g270) & (!g271) & (g284)) + ((!g74) & (sk[59]) & (g270) & (!g271) & (g284)) + ((g74) & (!sk[59]) & (!g270) & (g271) & (!g284)) + ((g74) & (!sk[59]) & (!g270) & (g271) & (g284)) + ((g74) & (!sk[59]) & (g270) & (g271) & (!g284)) + ((g74) & (!sk[59]) & (g270) & (g271) & (g284)) + ((g74) & (sk[59]) & (!g270) & (!g271) & (g284)));
	assign g286 = (((!g68) & (sk[60]) & (!g126)) + ((g68) & (!sk[60]) & (!g126)) + ((g68) & (!sk[60]) & (g126)));
	assign g287 = (((!g121) & (!g254) & (!sk[61]) & (g282)) + ((!g121) & (!g254) & (sk[61]) & (g282)) + ((!g121) & (g254) & (!sk[61]) & (!g282)) + ((!g121) & (g254) & (!sk[61]) & (g282)) + ((g121) & (!g254) & (!sk[61]) & (g282)) + ((g121) & (!g254) & (sk[61]) & (g282)) + ((g121) & (g254) & (!sk[61]) & (!g282)) + ((g121) & (g254) & (!sk[61]) & (g282)) + ((g121) & (g254) & (sk[61]) & (g282)));
	assign g288 = (((!g3) & (!g24) & (!sk[62]) & (g68) & (!g125) & (g126)) + ((!g3) & (!g24) & (!sk[62]) & (g68) & (g125) & (!g126)) + ((!g3) & (!g24) & (!sk[62]) & (g68) & (g125) & (g126)) + ((!g3) & (!g24) & (sk[62]) & (!g68) & (g125) & (!g126)) + ((!g3) & (!g24) & (sk[62]) & (g68) & (g125) & (!g126)) + ((!g3) & (g24) & (!sk[62]) & (!g68) & (!g125) & (!g126)) + ((!g3) & (g24) & (!sk[62]) & (!g68) & (!g125) & (g126)) + ((!g3) & (g24) & (!sk[62]) & (!g68) & (g125) & (!g126)) + ((!g3) & (g24) & (!sk[62]) & (!g68) & (g125) & (g126)) + ((!g3) & (g24) & (!sk[62]) & (g68) & (!g125) & (!g126)) + ((!g3) & (g24) & (!sk[62]) & (g68) & (!g125) & (g126)) + ((!g3) & (g24) & (!sk[62]) & (g68) & (g125) & (!g126)) + ((!g3) & (g24) & (!sk[62]) & (g68) & (g125) & (g126)) + ((!g3) & (g24) & (sk[62]) & (!g68) & (g125) & (!g126)) + ((g3) & (!g24) & (!sk[62]) & (g68) & (!g125) & (g126)) + ((g3) & (!g24) & (!sk[62]) & (g68) & (g125) & (!g126)) + ((g3) & (!g24) & (!sk[62]) & (g68) & (g125) & (g126)) + ((g3) & (!g24) & (sk[62]) & (!g68) & (g125) & (!g126)) + ((g3) & (!g24) & (sk[62]) & (!g68) & (g125) & (g126)) + ((g3) & (!g24) & (sk[62]) & (g68) & (g125) & (!g126)) + ((g3) & (g24) & (!sk[62]) & (!g68) & (!g125) & (!g126)) + ((g3) & (g24) & (!sk[62]) & (!g68) & (!g125) & (g126)) + ((g3) & (g24) & (!sk[62]) & (!g68) & (g125) & (!g126)) + ((g3) & (g24) & (!sk[62]) & (!g68) & (g125) & (g126)) + ((g3) & (g24) & (!sk[62]) & (g68) & (!g125) & (!g126)) + ((g3) & (g24) & (!sk[62]) & (g68) & (!g125) & (g126)) + ((g3) & (g24) & (!sk[62]) & (g68) & (g125) & (!g126)) + ((g3) & (g24) & (!sk[62]) & (g68) & (g125) & (g126)) + ((g3) & (g24) & (sk[62]) & (!g68) & (g125) & (!g126)) + ((g3) & (g24) & (sk[62]) & (!g68) & (g125) & (g126)));
	assign g289 = (((!g123) & (!g119) & (!g226) & (!g282) & (sk[63]) & (!g270)) + ((!g123) & (!g119) & (g226) & (!g282) & (!sk[63]) & (g270)) + ((!g123) & (!g119) & (g226) & (!g282) & (sk[63]) & (!g270)) + ((!g123) & (!g119) & (g226) & (g282) & (!sk[63]) & (!g270)) + ((!g123) & (!g119) & (g226) & (g282) & (!sk[63]) & (g270)) + ((!g123) & (!g119) & (g226) & (g282) & (sk[63]) & (!g270)) + ((!g123) & (g119) & (!g226) & (!g282) & (!sk[63]) & (!g270)) + ((!g123) & (g119) & (!g226) & (!g282) & (!sk[63]) & (g270)) + ((!g123) & (g119) & (!g226) & (!g282) & (sk[63]) & (!g270)) + ((!g123) & (g119) & (!g226) & (g282) & (!sk[63]) & (!g270)) + ((!g123) & (g119) & (!g226) & (g282) & (!sk[63]) & (g270)) + ((!g123) & (g119) & (g226) & (!g282) & (!sk[63]) & (!g270)) + ((!g123) & (g119) & (g226) & (!g282) & (!sk[63]) & (g270)) + ((!g123) & (g119) & (g226) & (!g282) & (sk[63]) & (!g270)) + ((!g123) & (g119) & (g226) & (g282) & (!sk[63]) & (!g270)) + ((!g123) & (g119) & (g226) & (g282) & (!sk[63]) & (g270)) + ((g123) & (!g119) & (!g226) & (!g282) & (sk[63]) & (!g270)) + ((g123) & (!g119) & (!g226) & (!g282) & (sk[63]) & (g270)) + ((g123) & (!g119) & (g226) & (!g282) & (!sk[63]) & (g270)) + ((g123) & (!g119) & (g226) & (!g282) & (sk[63]) & (!g270)) + ((g123) & (!g119) & (g226) & (!g282) & (sk[63]) & (g270)) + ((g123) & (!g119) & (g226) & (g282) & (!sk[63]) & (!g270)) + ((g123) & (!g119) & (g226) & (g282) & (!sk[63]) & (g270)) + ((g123) & (!g119) & (g226) & (g282) & (sk[63]) & (!g270)) + ((g123) & (!g119) & (g226) & (g282) & (sk[63]) & (g270)) + ((g123) & (g119) & (!g226) & (!g282) & (!sk[63]) & (!g270)) + ((g123) & (g119) & (!g226) & (!g282) & (!sk[63]) & (g270)) + ((g123) & (g119) & (!g226) & (!g282) & (sk[63]) & (!g270)) + ((g123) & (g119) & (!g226) & (g282) & (!sk[63]) & (!g270)) + ((g123) & (g119) & (!g226) & (g282) & (!sk[63]) & (g270)) + ((g123) & (g119) & (g226) & (!g282) & (!sk[63]) & (!g270)) + ((g123) & (g119) & (g226) & (!g282) & (!sk[63]) & (g270)) + ((g123) & (g119) & (g226) & (!g282) & (sk[63]) & (!g270)) + ((g123) & (g119) & (g226) & (g282) & (!sk[63]) & (!g270)) + ((g123) & (g119) & (g226) & (g282) & (!sk[63]) & (g270)));
	assign g290 = (((!g75) & (!g122) & (!g286) & (!g287) & (!g288) & (g289)) + ((!g75) & (g122) & (!g286) & (!g287) & (!g288) & (g289)) + ((g75) & (!g122) & (!g286) & (!g287) & (!g288) & (g289)) + ((g75) & (!g122) & (g286) & (!g287) & (!g288) & (g289)) + ((g75) & (g122) & (!g286) & (!g287) & (!g288) & (g289)));
	assign g291 = (((!i_8_) & (!sk[65]) & (!g73) & (g105) & (!g272)) + ((!i_8_) & (!sk[65]) & (!g73) & (g105) & (g272)) + ((!i_8_) & (!sk[65]) & (g73) & (g105) & (!g272)) + ((!i_8_) & (!sk[65]) & (g73) & (g105) & (g272)) + ((!i_8_) & (sk[65]) & (!g73) & (!g105) & (g272)) + ((!i_8_) & (sk[65]) & (g73) & (!g105) & (g272)) + ((i_8_) & (!sk[65]) & (!g73) & (g105) & (!g272)) + ((i_8_) & (!sk[65]) & (!g73) & (g105) & (g272)) + ((i_8_) & (!sk[65]) & (g73) & (g105) & (!g272)) + ((i_8_) & (!sk[65]) & (g73) & (g105) & (g272)) + ((i_8_) & (sk[65]) & (!g73) & (!g105) & (g272)) + ((i_8_) & (sk[65]) & (g73) & (!g105) & (g272)) + ((i_8_) & (sk[65]) & (g73) & (g105) & (g272)));
	assign g292 = (((!g142) & (!g227) & (!sk[66]) & (g275) & (!g282)) + ((!g142) & (!g227) & (!sk[66]) & (g275) & (g282)) + ((!g142) & (!g227) & (sk[66]) & (!g275) & (!g282)) + ((!g142) & (!g227) & (sk[66]) & (!g275) & (g282)) + ((!g142) & (g227) & (!sk[66]) & (g275) & (!g282)) + ((!g142) & (g227) & (!sk[66]) & (g275) & (g282)) + ((!g142) & (g227) & (sk[66]) & (!g275) & (!g282)) + ((g142) & (!g227) & (!sk[66]) & (g275) & (!g282)) + ((g142) & (!g227) & (!sk[66]) & (g275) & (g282)) + ((g142) & (!g227) & (sk[66]) & (!g275) & (!g282)) + ((g142) & (!g227) & (sk[66]) & (!g275) & (g282)) + ((g142) & (!g227) & (sk[66]) & (g275) & (!g282)) + ((g142) & (!g227) & (sk[66]) & (g275) & (g282)) + ((g142) & (g227) & (!sk[66]) & (g275) & (!g282)) + ((g142) & (g227) & (!sk[66]) & (g275) & (g282)) + ((g142) & (g227) & (sk[66]) & (!g275) & (!g282)));
	assign g293 = (((!i_8_) & (!sk[67]) & (!g24) & (g73) & (!g126) & (g105)) + ((!i_8_) & (!sk[67]) & (!g24) & (g73) & (g126) & (!g105)) + ((!i_8_) & (!sk[67]) & (!g24) & (g73) & (g126) & (g105)) + ((!i_8_) & (!sk[67]) & (g24) & (!g73) & (!g126) & (!g105)) + ((!i_8_) & (!sk[67]) & (g24) & (!g73) & (!g126) & (g105)) + ((!i_8_) & (!sk[67]) & (g24) & (!g73) & (g126) & (!g105)) + ((!i_8_) & (!sk[67]) & (g24) & (!g73) & (g126) & (g105)) + ((!i_8_) & (!sk[67]) & (g24) & (g73) & (!g126) & (!g105)) + ((!i_8_) & (!sk[67]) & (g24) & (g73) & (!g126) & (g105)) + ((!i_8_) & (!sk[67]) & (g24) & (g73) & (g126) & (!g105)) + ((!i_8_) & (!sk[67]) & (g24) & (g73) & (g126) & (g105)) + ((!i_8_) & (sk[67]) & (!g24) & (!g73) & (!g126) & (!g105)) + ((!i_8_) & (sk[67]) & (!g24) & (g73) & (!g126) & (!g105)) + ((i_8_) & (!sk[67]) & (!g24) & (g73) & (!g126) & (g105)) + ((i_8_) & (!sk[67]) & (!g24) & (g73) & (g126) & (!g105)) + ((i_8_) & (!sk[67]) & (!g24) & (g73) & (g126) & (g105)) + ((i_8_) & (!sk[67]) & (g24) & (!g73) & (!g126) & (!g105)) + ((i_8_) & (!sk[67]) & (g24) & (!g73) & (!g126) & (g105)) + ((i_8_) & (!sk[67]) & (g24) & (!g73) & (g126) & (!g105)) + ((i_8_) & (!sk[67]) & (g24) & (!g73) & (g126) & (g105)) + ((i_8_) & (!sk[67]) & (g24) & (g73) & (!g126) & (!g105)) + ((i_8_) & (!sk[67]) & (g24) & (g73) & (!g126) & (g105)) + ((i_8_) & (!sk[67]) & (g24) & (g73) & (g126) & (!g105)) + ((i_8_) & (!sk[67]) & (g24) & (g73) & (g126) & (g105)) + ((i_8_) & (sk[67]) & (!g24) & (!g73) & (!g126) & (!g105)) + ((i_8_) & (sk[67]) & (!g24) & (g73) & (!g126) & (!g105)) + ((i_8_) & (sk[67]) & (!g24) & (g73) & (!g126) & (g105)));
	assign g294 = (((!g25) & (!sk[68]) & (!g28) & (g105)) + ((!g25) & (!sk[68]) & (g28) & (!g105)) + ((!g25) & (!sk[68]) & (g28) & (g105)) + ((!g25) & (sk[68]) & (!g28) & (!g105)) + ((!g25) & (sk[68]) & (g28) & (!g105)) + ((g25) & (!sk[68]) & (!g28) & (g105)) + ((g25) & (!sk[68]) & (g28) & (!g105)) + ((g25) & (!sk[68]) & (g28) & (g105)) + ((g25) & (sk[68]) & (g28) & (!g105)));
	assign g295 = (((!sk[69]) & (g68) & (!g83)) + ((!sk[69]) & (g68) & (g83)) + ((sk[69]) & (!g68) & (g83)));
	assign g296 = (((!sk[70]) & (g107) & (!g68)) + ((!sk[70]) & (g107) & (g68)) + ((sk[70]) & (!g107) & (!g68)));
	assign g297 = (((!g125) & (!g142) & (!g295) & (!g296) & (sk[71]) & (!g278)) + ((!g125) & (!g142) & (!g295) & (g296) & (sk[71]) & (!g278)) + ((!g125) & (!g142) & (g295) & (!g296) & (!sk[71]) & (g278)) + ((!g125) & (!g142) & (g295) & (g296) & (!sk[71]) & (!g278)) + ((!g125) & (!g142) & (g295) & (g296) & (!sk[71]) & (g278)) + ((!g125) & (g142) & (!g295) & (!g296) & (!sk[71]) & (!g278)) + ((!g125) & (g142) & (!g295) & (!g296) & (!sk[71]) & (g278)) + ((!g125) & (g142) & (!g295) & (!g296) & (sk[71]) & (!g278)) + ((!g125) & (g142) & (!g295) & (!g296) & (sk[71]) & (g278)) + ((!g125) & (g142) & (!g295) & (g296) & (!sk[71]) & (!g278)) + ((!g125) & (g142) & (!g295) & (g296) & (!sk[71]) & (g278)) + ((!g125) & (g142) & (!g295) & (g296) & (sk[71]) & (!g278)) + ((!g125) & (g142) & (!g295) & (g296) & (sk[71]) & (g278)) + ((!g125) & (g142) & (g295) & (!g296) & (!sk[71]) & (!g278)) + ((!g125) & (g142) & (g295) & (!g296) & (!sk[71]) & (g278)) + ((!g125) & (g142) & (g295) & (!g296) & (sk[71]) & (!g278)) + ((!g125) & (g142) & (g295) & (!g296) & (sk[71]) & (g278)) + ((!g125) & (g142) & (g295) & (g296) & (!sk[71]) & (!g278)) + ((!g125) & (g142) & (g295) & (g296) & (!sk[71]) & (g278)) + ((!g125) & (g142) & (g295) & (g296) & (sk[71]) & (!g278)) + ((!g125) & (g142) & (g295) & (g296) & (sk[71]) & (g278)) + ((g125) & (!g142) & (!g295) & (!g296) & (sk[71]) & (!g278)) + ((g125) & (!g142) & (g295) & (!g296) & (!sk[71]) & (g278)) + ((g125) & (!g142) & (g295) & (g296) & (!sk[71]) & (!g278)) + ((g125) & (!g142) & (g295) & (g296) & (!sk[71]) & (g278)) + ((g125) & (g142) & (!g295) & (!g296) & (!sk[71]) & (!g278)) + ((g125) & (g142) & (!g295) & (!g296) & (!sk[71]) & (g278)) + ((g125) & (g142) & (!g295) & (!g296) & (sk[71]) & (!g278)) + ((g125) & (g142) & (!g295) & (!g296) & (sk[71]) & (g278)) + ((g125) & (g142) & (!g295) & (g296) & (!sk[71]) & (!g278)) + ((g125) & (g142) & (!g295) & (g296) & (!sk[71]) & (g278)) + ((g125) & (g142) & (g295) & (!g296) & (!sk[71]) & (!g278)) + ((g125) & (g142) & (g295) & (!g296) & (!sk[71]) & (g278)) + ((g125) & (g142) & (g295) & (g296) & (!sk[71]) & (!g278)) + ((g125) & (g142) & (g295) & (g296) & (!sk[71]) & (g278)));
	assign g298 = (((!g291) & (!g292) & (!sk[72]) & (g293) & (!g294) & (g297)) + ((!g291) & (!g292) & (!sk[72]) & (g293) & (g294) & (!g297)) + ((!g291) & (!g292) & (!sk[72]) & (g293) & (g294) & (g297)) + ((!g291) & (g292) & (!sk[72]) & (!g293) & (!g294) & (!g297)) + ((!g291) & (g292) & (!sk[72]) & (!g293) & (!g294) & (g297)) + ((!g291) & (g292) & (!sk[72]) & (!g293) & (g294) & (!g297)) + ((!g291) & (g292) & (!sk[72]) & (!g293) & (g294) & (g297)) + ((!g291) & (g292) & (!sk[72]) & (g293) & (!g294) & (!g297)) + ((!g291) & (g292) & (!sk[72]) & (g293) & (!g294) & (g297)) + ((!g291) & (g292) & (!sk[72]) & (g293) & (g294) & (!g297)) + ((!g291) & (g292) & (!sk[72]) & (g293) & (g294) & (g297)) + ((!g291) & (g292) & (sk[72]) & (!g293) & (!g294) & (g297)) + ((g291) & (!g292) & (!sk[72]) & (g293) & (!g294) & (g297)) + ((g291) & (!g292) & (!sk[72]) & (g293) & (g294) & (!g297)) + ((g291) & (!g292) & (!sk[72]) & (g293) & (g294) & (g297)) + ((g291) & (g292) & (!sk[72]) & (!g293) & (!g294) & (!g297)) + ((g291) & (g292) & (!sk[72]) & (!g293) & (!g294) & (g297)) + ((g291) & (g292) & (!sk[72]) & (!g293) & (g294) & (!g297)) + ((g291) & (g292) & (!sk[72]) & (!g293) & (g294) & (g297)) + ((g291) & (g292) & (!sk[72]) & (g293) & (!g294) & (!g297)) + ((g291) & (g292) & (!sk[72]) & (g293) & (!g294) & (g297)) + ((g291) & (g292) & (!sk[72]) & (g293) & (g294) & (!g297)) + ((g291) & (g292) & (!sk[72]) & (g293) & (g294) & (g297)));
	assign g299 = (((!sk[73]) & (!g24) & (!g68) & (g122) & (!g83)) + ((!sk[73]) & (!g24) & (!g68) & (g122) & (g83)) + ((!sk[73]) & (!g24) & (g68) & (g122) & (!g83)) + ((!sk[73]) & (!g24) & (g68) & (g122) & (g83)) + ((!sk[73]) & (g24) & (!g68) & (g122) & (!g83)) + ((!sk[73]) & (g24) & (!g68) & (g122) & (g83)) + ((!sk[73]) & (g24) & (g68) & (g122) & (!g83)) + ((!sk[73]) & (g24) & (g68) & (g122) & (g83)) + ((sk[73]) & (!g24) & (!g68) & (g122) & (g83)) + ((sk[73]) & (!g24) & (g68) & (g122) & (g83)) + ((sk[73]) & (g24) & (!g68) & (g122) & (g83)));
	assign g300 = (((!sk[74]) & (!i_8_) & (!g24) & (g73) & (!g68) & (g126)) + ((!sk[74]) & (!i_8_) & (!g24) & (g73) & (g68) & (!g126)) + ((!sk[74]) & (!i_8_) & (!g24) & (g73) & (g68) & (g126)) + ((!sk[74]) & (!i_8_) & (g24) & (!g73) & (!g68) & (!g126)) + ((!sk[74]) & (!i_8_) & (g24) & (!g73) & (!g68) & (g126)) + ((!sk[74]) & (!i_8_) & (g24) & (!g73) & (g68) & (!g126)) + ((!sk[74]) & (!i_8_) & (g24) & (!g73) & (g68) & (g126)) + ((!sk[74]) & (!i_8_) & (g24) & (g73) & (!g68) & (!g126)) + ((!sk[74]) & (!i_8_) & (g24) & (g73) & (!g68) & (g126)) + ((!sk[74]) & (!i_8_) & (g24) & (g73) & (g68) & (!g126)) + ((!sk[74]) & (!i_8_) & (g24) & (g73) & (g68) & (g126)) + ((!sk[74]) & (i_8_) & (!g24) & (g73) & (!g68) & (g126)) + ((!sk[74]) & (i_8_) & (!g24) & (g73) & (g68) & (!g126)) + ((!sk[74]) & (i_8_) & (!g24) & (g73) & (g68) & (g126)) + ((!sk[74]) & (i_8_) & (g24) & (!g73) & (!g68) & (!g126)) + ((!sk[74]) & (i_8_) & (g24) & (!g73) & (!g68) & (g126)) + ((!sk[74]) & (i_8_) & (g24) & (!g73) & (g68) & (!g126)) + ((!sk[74]) & (i_8_) & (g24) & (!g73) & (g68) & (g126)) + ((!sk[74]) & (i_8_) & (g24) & (g73) & (!g68) & (!g126)) + ((!sk[74]) & (i_8_) & (g24) & (g73) & (!g68) & (g126)) + ((!sk[74]) & (i_8_) & (g24) & (g73) & (g68) & (!g126)) + ((!sk[74]) & (i_8_) & (g24) & (g73) & (g68) & (g126)) + ((sk[74]) & (!i_8_) & (!g24) & (g73) & (!g68) & (!g126)) + ((sk[74]) & (!i_8_) & (!g24) & (g73) & (g68) & (!g126)) + ((sk[74]) & (!i_8_) & (g24) & (g73) & (!g68) & (!g126)));
	assign g301 = (((!g28) & (!sk[75]) & (!g135) & (g122) & (!g275)) + ((!g28) & (!sk[75]) & (!g135) & (g122) & (g275)) + ((!g28) & (!sk[75]) & (g135) & (g122) & (!g275)) + ((!g28) & (!sk[75]) & (g135) & (g122) & (g275)) + ((!g28) & (sk[75]) & (!g135) & (!g122) & (!g275)) + ((!g28) & (sk[75]) & (!g135) & (g122) & (!g275)) + ((!g28) & (sk[75]) & (g135) & (!g122) & (!g275)) + ((!g28) & (sk[75]) & (g135) & (!g122) & (g275)) + ((!g28) & (sk[75]) & (g135) & (g122) & (!g275)) + ((g28) & (!sk[75]) & (!g135) & (g122) & (!g275)) + ((g28) & (!sk[75]) & (!g135) & (g122) & (g275)) + ((g28) & (!sk[75]) & (g135) & (g122) & (!g275)) + ((g28) & (!sk[75]) & (g135) & (g122) & (g275)) + ((g28) & (sk[75]) & (g135) & (!g122) & (!g275)) + ((g28) & (sk[75]) & (g135) & (!g122) & (g275)));
	assign g302 = (((!g135) & (!g122) & (!g273) & (!g281) & (!g296) & (!g278)) + ((!g135) & (!g122) & (!g273) & (!g281) & (!g296) & (g278)) + ((!g135) & (g122) & (!g273) & (!g281) & (!g296) & (!g278)) + ((g135) & (!g122) & (!g273) & (!g281) & (!g296) & (!g278)) + ((g135) & (!g122) & (!g273) & (!g281) & (!g296) & (g278)) + ((g135) & (!g122) & (!g273) & (!g281) & (g296) & (!g278)) + ((g135) & (!g122) & (!g273) & (!g281) & (g296) & (g278)) + ((g135) & (!g122) & (!g273) & (g281) & (!g296) & (!g278)) + ((g135) & (!g122) & (!g273) & (g281) & (!g296) & (g278)) + ((g135) & (!g122) & (!g273) & (g281) & (g296) & (!g278)) + ((g135) & (!g122) & (!g273) & (g281) & (g296) & (g278)) + ((g135) & (!g122) & (g273) & (!g281) & (!g296) & (!g278)) + ((g135) & (!g122) & (g273) & (!g281) & (!g296) & (g278)) + ((g135) & (!g122) & (g273) & (!g281) & (g296) & (!g278)) + ((g135) & (!g122) & (g273) & (!g281) & (g296) & (g278)) + ((g135) & (!g122) & (g273) & (g281) & (!g296) & (!g278)) + ((g135) & (!g122) & (g273) & (g281) & (!g296) & (g278)) + ((g135) & (!g122) & (g273) & (g281) & (g296) & (!g278)) + ((g135) & (!g122) & (g273) & (g281) & (g296) & (g278)) + ((g135) & (g122) & (!g273) & (!g281) & (!g296) & (!g278)) + ((g135) & (g122) & (!g273) & (!g281) & (g296) & (!g278)) + ((g135) & (g122) & (!g273) & (g281) & (!g296) & (!g278)) + ((g135) & (g122) & (!g273) & (g281) & (g296) & (!g278)));
	assign g303 = (((!g24) & (!g35) & (!sk[77]) & (g107) & (!g123) & (g130)) + ((!g24) & (!g35) & (!sk[77]) & (g107) & (g123) & (!g130)) + ((!g24) & (!g35) & (!sk[77]) & (g107) & (g123) & (g130)) + ((!g24) & (!g35) & (sk[77]) & (!g107) & (!g123) & (!g130)) + ((!g24) & (!g35) & (sk[77]) & (!g107) & (!g123) & (g130)) + ((!g24) & (!g35) & (sk[77]) & (!g107) & (g123) & (!g130)) + ((!g24) & (g35) & (!sk[77]) & (!g107) & (!g123) & (!g130)) + ((!g24) & (g35) & (!sk[77]) & (!g107) & (!g123) & (g130)) + ((!g24) & (g35) & (!sk[77]) & (!g107) & (g123) & (!g130)) + ((!g24) & (g35) & (!sk[77]) & (!g107) & (g123) & (g130)) + ((!g24) & (g35) & (!sk[77]) & (g107) & (!g123) & (!g130)) + ((!g24) & (g35) & (!sk[77]) & (g107) & (!g123) & (g130)) + ((!g24) & (g35) & (!sk[77]) & (g107) & (g123) & (!g130)) + ((!g24) & (g35) & (!sk[77]) & (g107) & (g123) & (g130)) + ((!g24) & (g35) & (sk[77]) & (!g107) & (!g123) & (!g130)) + ((!g24) & (g35) & (sk[77]) & (!g107) & (!g123) & (g130)) + ((!g24) & (g35) & (sk[77]) & (!g107) & (g123) & (!g130)) + ((!g24) & (g35) & (sk[77]) & (g107) & (!g123) & (!g130)) + ((!g24) & (g35) & (sk[77]) & (g107) & (!g123) & (g130)) + ((!g24) & (g35) & (sk[77]) & (g107) & (g123) & (!g130)) + ((g24) & (!g35) & (!sk[77]) & (g107) & (!g123) & (g130)) + ((g24) & (!g35) & (!sk[77]) & (g107) & (g123) & (!g130)) + ((g24) & (!g35) & (!sk[77]) & (g107) & (g123) & (g130)) + ((g24) & (g35) & (!sk[77]) & (!g107) & (!g123) & (!g130)) + ((g24) & (g35) & (!sk[77]) & (!g107) & (!g123) & (g130)) + ((g24) & (g35) & (!sk[77]) & (!g107) & (g123) & (!g130)) + ((g24) & (g35) & (!sk[77]) & (!g107) & (g123) & (g130)) + ((g24) & (g35) & (!sk[77]) & (g107) & (!g123) & (!g130)) + ((g24) & (g35) & (!sk[77]) & (g107) & (!g123) & (g130)) + ((g24) & (g35) & (!sk[77]) & (g107) & (g123) & (!g130)) + ((g24) & (g35) & (!sk[77]) & (g107) & (g123) & (g130)));
	assign g304 = (((!g299) & (!g300) & (!sk[78]) & (g301) & (!g302) & (g303)) + ((!g299) & (!g300) & (!sk[78]) & (g301) & (g302) & (!g303)) + ((!g299) & (!g300) & (!sk[78]) & (g301) & (g302) & (g303)) + ((!g299) & (!g300) & (sk[78]) & (g301) & (g302) & (!g303)) + ((!g299) & (g300) & (!sk[78]) & (!g301) & (!g302) & (!g303)) + ((!g299) & (g300) & (!sk[78]) & (!g301) & (!g302) & (g303)) + ((!g299) & (g300) & (!sk[78]) & (!g301) & (g302) & (!g303)) + ((!g299) & (g300) & (!sk[78]) & (!g301) & (g302) & (g303)) + ((!g299) & (g300) & (!sk[78]) & (g301) & (!g302) & (!g303)) + ((!g299) & (g300) & (!sk[78]) & (g301) & (!g302) & (g303)) + ((!g299) & (g300) & (!sk[78]) & (g301) & (g302) & (!g303)) + ((!g299) & (g300) & (!sk[78]) & (g301) & (g302) & (g303)) + ((g299) & (!g300) & (!sk[78]) & (g301) & (!g302) & (g303)) + ((g299) & (!g300) & (!sk[78]) & (g301) & (g302) & (!g303)) + ((g299) & (!g300) & (!sk[78]) & (g301) & (g302) & (g303)) + ((g299) & (g300) & (!sk[78]) & (!g301) & (!g302) & (!g303)) + ((g299) & (g300) & (!sk[78]) & (!g301) & (!g302) & (g303)) + ((g299) & (g300) & (!sk[78]) & (!g301) & (g302) & (!g303)) + ((g299) & (g300) & (!sk[78]) & (!g301) & (g302) & (g303)) + ((g299) & (g300) & (!sk[78]) & (g301) & (!g302) & (!g303)) + ((g299) & (g300) & (!sk[78]) & (g301) & (!g302) & (g303)) + ((g299) & (g300) & (!sk[78]) & (g301) & (g302) & (!g303)) + ((g299) & (g300) & (!sk[78]) & (g301) & (g302) & (g303)));
	assign g305 = (((!sk[79]) & (!g25) & (!g102) & (g278)) + ((!sk[79]) & (!g25) & (g102) & (!g278)) + ((!sk[79]) & (!g25) & (g102) & (g278)) + ((!sk[79]) & (g25) & (!g102) & (g278)) + ((!sk[79]) & (g25) & (g102) & (!g278)) + ((!sk[79]) & (g25) & (g102) & (g278)) + ((sk[79]) & (!g25) & (g102) & (!g278)) + ((sk[79]) & (!g25) & (g102) & (g278)) + ((sk[79]) & (g25) & (g102) & (g278)));
	assign g306 = (((g225) & (!sk[80]) & (!g275)) + ((g225) & (!sk[80]) & (g275)) + ((g225) & (sk[80]) & (g275)));
	assign g307 = (((!g24) & (!g35) & (!g102) & (g83) & (sk[81]) & (!g105)) + ((!g24) & (!g35) & (g102) & (!g83) & (!sk[81]) & (g105)) + ((!g24) & (!g35) & (g102) & (g83) & (!sk[81]) & (!g105)) + ((!g24) & (!g35) & (g102) & (g83) & (!sk[81]) & (g105)) + ((!g24) & (!g35) & (g102) & (g83) & (sk[81]) & (!g105)) + ((!g24) & (g35) & (!g102) & (!g83) & (!sk[81]) & (!g105)) + ((!g24) & (g35) & (!g102) & (!g83) & (!sk[81]) & (g105)) + ((!g24) & (g35) & (!g102) & (!g83) & (sk[81]) & (!g105)) + ((!g24) & (g35) & (!g102) & (g83) & (!sk[81]) & (!g105)) + ((!g24) & (g35) & (!g102) & (g83) & (!sk[81]) & (g105)) + ((!g24) & (g35) & (!g102) & (g83) & (sk[81]) & (!g105)) + ((!g24) & (g35) & (g102) & (!g83) & (!sk[81]) & (!g105)) + ((!g24) & (g35) & (g102) & (!g83) & (!sk[81]) & (g105)) + ((!g24) & (g35) & (g102) & (!g83) & (sk[81]) & (!g105)) + ((!g24) & (g35) & (g102) & (!g83) & (sk[81]) & (g105)) + ((!g24) & (g35) & (g102) & (g83) & (!sk[81]) & (!g105)) + ((!g24) & (g35) & (g102) & (g83) & (!sk[81]) & (g105)) + ((!g24) & (g35) & (g102) & (g83) & (sk[81]) & (!g105)) + ((!g24) & (g35) & (g102) & (g83) & (sk[81]) & (g105)) + ((g24) & (!g35) & (g102) & (!g83) & (!sk[81]) & (g105)) + ((g24) & (!g35) & (g102) & (g83) & (!sk[81]) & (!g105)) + ((g24) & (!g35) & (g102) & (g83) & (!sk[81]) & (g105)) + ((g24) & (g35) & (!g102) & (!g83) & (!sk[81]) & (!g105)) + ((g24) & (g35) & (!g102) & (!g83) & (!sk[81]) & (g105)) + ((g24) & (g35) & (!g102) & (g83) & (!sk[81]) & (!g105)) + ((g24) & (g35) & (!g102) & (g83) & (!sk[81]) & (g105)) + ((g24) & (g35) & (g102) & (!g83) & (!sk[81]) & (!g105)) + ((g24) & (g35) & (g102) & (!g83) & (!sk[81]) & (g105)) + ((g24) & (g35) & (g102) & (g83) & (!sk[81]) & (!g105)) + ((g24) & (g35) & (g102) & (g83) & (!sk[81]) & (g105)));
	assign g308 = (((!sk[82]) & (!g24) & (!g27) & (g68) & (!g102) & (g83)) + ((!sk[82]) & (!g24) & (!g27) & (g68) & (g102) & (!g83)) + ((!sk[82]) & (!g24) & (!g27) & (g68) & (g102) & (g83)) + ((!sk[82]) & (!g24) & (g27) & (!g68) & (!g102) & (!g83)) + ((!sk[82]) & (!g24) & (g27) & (!g68) & (!g102) & (g83)) + ((!sk[82]) & (!g24) & (g27) & (!g68) & (g102) & (!g83)) + ((!sk[82]) & (!g24) & (g27) & (!g68) & (g102) & (g83)) + ((!sk[82]) & (!g24) & (g27) & (g68) & (!g102) & (!g83)) + ((!sk[82]) & (!g24) & (g27) & (g68) & (!g102) & (g83)) + ((!sk[82]) & (!g24) & (g27) & (g68) & (g102) & (!g83)) + ((!sk[82]) & (!g24) & (g27) & (g68) & (g102) & (g83)) + ((!sk[82]) & (g24) & (!g27) & (g68) & (!g102) & (g83)) + ((!sk[82]) & (g24) & (!g27) & (g68) & (g102) & (!g83)) + ((!sk[82]) & (g24) & (!g27) & (g68) & (g102) & (g83)) + ((!sk[82]) & (g24) & (g27) & (!g68) & (!g102) & (!g83)) + ((!sk[82]) & (g24) & (g27) & (!g68) & (!g102) & (g83)) + ((!sk[82]) & (g24) & (g27) & (!g68) & (g102) & (!g83)) + ((!sk[82]) & (g24) & (g27) & (!g68) & (g102) & (g83)) + ((!sk[82]) & (g24) & (g27) & (g68) & (!g102) & (!g83)) + ((!sk[82]) & (g24) & (g27) & (g68) & (!g102) & (g83)) + ((!sk[82]) & (g24) & (g27) & (g68) & (g102) & (!g83)) + ((!sk[82]) & (g24) & (g27) & (g68) & (g102) & (g83)) + ((sk[82]) & (!g24) & (!g27) & (!g68) & (g102) & (g83)) + ((sk[82]) & (!g24) & (!g27) & (g68) & (g102) & (g83)) + ((sk[82]) & (!g24) & (g27) & (!g68) & (g102) & (!g83)) + ((sk[82]) & (!g24) & (g27) & (!g68) & (g102) & (g83)) + ((sk[82]) & (!g24) & (g27) & (g68) & (g102) & (!g83)) + ((sk[82]) & (!g24) & (g27) & (g68) & (g102) & (g83)) + ((sk[82]) & (g24) & (!g27) & (!g68) & (g102) & (g83)) + ((sk[82]) & (g24) & (g27) & (!g68) & (g102) & (g83)));
	assign g309 = (((!g24) & (sk[83]) & (!g107)) + ((g24) & (!sk[83]) & (!g107)) + ((g24) & (!sk[83]) & (g107)));
	assign g310 = (((!g102) & (!g272) & (!sk[84]) & (g309)) + ((!g102) & (g272) & (!sk[84]) & (!g309)) + ((!g102) & (g272) & (!sk[84]) & (g309)) + ((g102) & (!g272) & (!sk[84]) & (g309)) + ((g102) & (!g272) & (sk[84]) & (g309)) + ((g102) & (g272) & (!sk[84]) & (!g309)) + ((g102) & (g272) & (!sk[84]) & (g309)) + ((g102) & (g272) & (sk[84]) & (!g309)) + ((g102) & (g272) & (sk[84]) & (g309)));
	assign g311 = (((!i_8_) & (!g73) & (!sk[85]) & (g309) & (!g296)) + ((!i_8_) & (!g73) & (!sk[85]) & (g309) & (g296)) + ((!i_8_) & (g73) & (!sk[85]) & (g309) & (!g296)) + ((!i_8_) & (g73) & (!sk[85]) & (g309) & (g296)) + ((!i_8_) & (g73) & (sk[85]) & (g309) & (!g296)) + ((!i_8_) & (g73) & (sk[85]) & (g309) & (g296)) + ((i_8_) & (!g73) & (!sk[85]) & (g309) & (!g296)) + ((i_8_) & (!g73) & (!sk[85]) & (g309) & (g296)) + ((i_8_) & (g73) & (!sk[85]) & (g309) & (!g296)) + ((i_8_) & (g73) & (!sk[85]) & (g309) & (g296)) + ((i_8_) & (g73) & (sk[85]) & (!g309) & (g296)) + ((i_8_) & (g73) & (sk[85]) & (g309) & (g296)));
	assign g312 = (((!g305) & (!g306) & (!g307) & (!g308) & (!g310) & (!g311)));
	assign g313 = (((g43) & (!sk[87]) & (!g166)) + ((g43) & (!sk[87]) & (g166)) + ((g43) & (sk[87]) & (g166)));
	assign g314 = (((!g24) & (!sk[88]) & (!g83) & (g130)) + ((!g24) & (!sk[88]) & (g83) & (!g130)) + ((!g24) & (!sk[88]) & (g83) & (g130)) + ((!g24) & (sk[88]) & (g83) & (!g130)) + ((g24) & (!sk[88]) & (!g83) & (g130)) + ((g24) & (!sk[88]) & (g83) & (!g130)) + ((g24) & (!sk[88]) & (g83) & (g130)));
	assign g315 = (((!sk[89]) & (i_15_) & (!g24)) + ((!sk[89]) & (i_15_) & (g24)) + ((sk[89]) & (!i_15_) & (!g24)));
	assign g316 = (((!g151) & (!g313) & (!g278) & (!g314) & (!g315) & (g1632)) + ((!g151) & (!g313) & (!g278) & (!g314) & (g315) & (g1632)) + ((!g151) & (!g313) & (g278) & (!g314) & (!g315) & (g1632)) + ((!g151) & (!g313) & (g278) & (!g314) & (g315) & (g1632)) + ((!g151) & (g313) & (!g278) & (!g314) & (!g315) & (g1632)) + ((!g151) & (g313) & (!g278) & (!g314) & (g315) & (g1632)) + ((g151) & (!g313) & (!g278) & (!g314) & (!g315) & (g1632)) + ((g151) & (!g313) & (g278) & (!g314) & (!g315) & (g1632)) + ((g151) & (g313) & (!g278) & (!g314) & (!g315) & (g1632)));
	assign g317 = (((!g131) & (!sk[91]) & (!g272) & (g273)) + ((!g131) & (!sk[91]) & (g272) & (!g273)) + ((!g131) & (!sk[91]) & (g272) & (g273)) + ((!g131) & (sk[91]) & (!g272) & (g273)) + ((!g131) & (sk[91]) & (g272) & (!g273)) + ((!g131) & (sk[91]) & (g272) & (g273)) + ((g131) & (!sk[91]) & (!g272) & (g273)) + ((g131) & (!sk[91]) & (g272) & (!g273)) + ((g131) & (!sk[91]) & (g272) & (g273)));
	assign g318 = (((!g25) & (!sk[92]) & (!g125) & (g278)) + ((!g25) & (!sk[92]) & (g125) & (!g278)) + ((!g25) & (!sk[92]) & (g125) & (g278)) + ((!g25) & (sk[92]) & (g125) & (!g278)) + ((!g25) & (sk[92]) & (g125) & (g278)) + ((g25) & (!sk[92]) & (!g125) & (g278)) + ((g25) & (!sk[92]) & (g125) & (!g278)) + ((g25) & (!sk[92]) & (g125) & (g278)) + ((g25) & (sk[92]) & (g125) & (g278)));
	assign g319 = (((!g131) & (!sk[93]) & (!g295) & (g281) & (!g296)) + ((!g131) & (!sk[93]) & (!g295) & (g281) & (g296)) + ((!g131) & (!sk[93]) & (g295) & (g281) & (!g296)) + ((!g131) & (!sk[93]) & (g295) & (g281) & (g296)) + ((!g131) & (sk[93]) & (!g295) & (!g281) & (g296)) + ((!g131) & (sk[93]) & (!g295) & (g281) & (!g296)) + ((!g131) & (sk[93]) & (!g295) & (g281) & (g296)) + ((!g131) & (sk[93]) & (g295) & (!g281) & (!g296)) + ((!g131) & (sk[93]) & (g295) & (!g281) & (g296)) + ((!g131) & (sk[93]) & (g295) & (g281) & (!g296)) + ((!g131) & (sk[93]) & (g295) & (g281) & (g296)) + ((g131) & (!sk[93]) & (!g295) & (g281) & (!g296)) + ((g131) & (!sk[93]) & (!g295) & (g281) & (g296)) + ((g131) & (!sk[93]) & (g295) & (g281) & (!g296)) + ((g131) & (!sk[93]) & (g295) & (g281) & (g296)));
	assign g320 = (((!g125) & (!g275) & (!sk[94]) & (g273) & (!g281)) + ((!g125) & (!g275) & (!sk[94]) & (g273) & (g281)) + ((!g125) & (g275) & (!sk[94]) & (g273) & (!g281)) + ((!g125) & (g275) & (!sk[94]) & (g273) & (g281)) + ((g125) & (!g275) & (!sk[94]) & (g273) & (!g281)) + ((g125) & (!g275) & (!sk[94]) & (g273) & (g281)) + ((g125) & (!g275) & (sk[94]) & (!g273) & (g281)) + ((g125) & (!g275) & (sk[94]) & (g273) & (!g281)) + ((g125) & (!g275) & (sk[94]) & (g273) & (g281)) + ((g125) & (g275) & (!sk[94]) & (g273) & (!g281)) + ((g125) & (g275) & (!sk[94]) & (g273) & (g281)) + ((g125) & (g275) & (sk[94]) & (!g273) & (!g281)) + ((g125) & (g275) & (sk[94]) & (!g273) & (g281)) + ((g125) & (g275) & (sk[94]) & (g273) & (!g281)) + ((g125) & (g275) & (sk[94]) & (g273) & (g281)));
	assign g321 = (((!g317) & (!g318) & (!sk[95]) & (g1625) & (!g319) & (g320)) + ((!g317) & (!g318) & (!sk[95]) & (g1625) & (g319) & (!g320)) + ((!g317) & (!g318) & (!sk[95]) & (g1625) & (g319) & (g320)) + ((!g317) & (!g318) & (sk[95]) & (g1625) & (!g319) & (!g320)) + ((!g317) & (g318) & (!sk[95]) & (!g1625) & (!g319) & (!g320)) + ((!g317) & (g318) & (!sk[95]) & (!g1625) & (!g319) & (g320)) + ((!g317) & (g318) & (!sk[95]) & (!g1625) & (g319) & (!g320)) + ((!g317) & (g318) & (!sk[95]) & (!g1625) & (g319) & (g320)) + ((!g317) & (g318) & (!sk[95]) & (g1625) & (!g319) & (!g320)) + ((!g317) & (g318) & (!sk[95]) & (g1625) & (!g319) & (g320)) + ((!g317) & (g318) & (!sk[95]) & (g1625) & (g319) & (!g320)) + ((!g317) & (g318) & (!sk[95]) & (g1625) & (g319) & (g320)) + ((g317) & (!g318) & (!sk[95]) & (g1625) & (!g319) & (g320)) + ((g317) & (!g318) & (!sk[95]) & (g1625) & (g319) & (!g320)) + ((g317) & (!g318) & (!sk[95]) & (g1625) & (g319) & (g320)) + ((g317) & (g318) & (!sk[95]) & (!g1625) & (!g319) & (!g320)) + ((g317) & (g318) & (!sk[95]) & (!g1625) & (!g319) & (g320)) + ((g317) & (g318) & (!sk[95]) & (!g1625) & (g319) & (!g320)) + ((g317) & (g318) & (!sk[95]) & (!g1625) & (g319) & (g320)) + ((g317) & (g318) & (!sk[95]) & (g1625) & (!g319) & (!g320)) + ((g317) & (g318) & (!sk[95]) & (g1625) & (!g319) & (g320)) + ((g317) & (g318) & (!sk[95]) & (g1625) & (g319) & (!g320)) + ((g317) & (g318) & (!sk[95]) & (g1625) & (g319) & (g320)));
	assign g322 = (((g290) & (g298) & (g304) & (g312) & (g316) & (g321)));
	assign g323 = (((!sk[97]) & (!i_10_) & (!i_11_) & (i_15_) & (!g24)) + ((!sk[97]) & (!i_10_) & (!i_11_) & (i_15_) & (g24)) + ((!sk[97]) & (!i_10_) & (i_11_) & (i_15_) & (!g24)) + ((!sk[97]) & (!i_10_) & (i_11_) & (i_15_) & (g24)) + ((!sk[97]) & (i_10_) & (!i_11_) & (i_15_) & (!g24)) + ((!sk[97]) & (i_10_) & (!i_11_) & (i_15_) & (g24)) + ((!sk[97]) & (i_10_) & (i_11_) & (i_15_) & (!g24)) + ((!sk[97]) & (i_10_) & (i_11_) & (i_15_) & (g24)) + ((sk[97]) & (!i_10_) & (!i_11_) & (!i_15_) & (!g24)) + ((sk[97]) & (!i_10_) & (!i_11_) & (!i_15_) & (g24)) + ((sk[97]) & (!i_10_) & (!i_11_) & (i_15_) & (!g24)) + ((sk[97]) & (!i_10_) & (!i_11_) & (i_15_) & (g24)) + ((sk[97]) & (!i_10_) & (i_11_) & (!i_15_) & (!g24)) + ((sk[97]) & (!i_10_) & (i_11_) & (!i_15_) & (g24)) + ((sk[97]) & (!i_10_) & (i_11_) & (i_15_) & (!g24)) + ((sk[97]) & (!i_10_) & (i_11_) & (i_15_) & (g24)) + ((sk[97]) & (i_10_) & (!i_11_) & (!i_15_) & (!g24)) + ((sk[97]) & (i_10_) & (!i_11_) & (!i_15_) & (g24)) + ((sk[97]) & (i_10_) & (!i_11_) & (i_15_) & (!g24)) + ((sk[97]) & (i_10_) & (!i_11_) & (i_15_) & (g24)) + ((sk[97]) & (i_10_) & (i_11_) & (!i_15_) & (g24)) + ((sk[97]) & (i_10_) & (i_11_) & (i_15_) & (!g24)) + ((sk[97]) & (i_10_) & (i_11_) & (i_15_) & (g24)));
	assign g324 = (((!i_8_) & (!i_9_) & (!sk[98]) & (i_10_) & (!i_11_) & (i_15_)) + ((!i_8_) & (!i_9_) & (!sk[98]) & (i_10_) & (i_11_) & (!i_15_)) + ((!i_8_) & (!i_9_) & (!sk[98]) & (i_10_) & (i_11_) & (i_15_)) + ((!i_8_) & (!i_9_) & (sk[98]) & (!i_10_) & (i_11_) & (!i_15_)) + ((!i_8_) & (i_9_) & (!sk[98]) & (!i_10_) & (!i_11_) & (!i_15_)) + ((!i_8_) & (i_9_) & (!sk[98]) & (!i_10_) & (!i_11_) & (i_15_)) + ((!i_8_) & (i_9_) & (!sk[98]) & (!i_10_) & (i_11_) & (!i_15_)) + ((!i_8_) & (i_9_) & (!sk[98]) & (!i_10_) & (i_11_) & (i_15_)) + ((!i_8_) & (i_9_) & (!sk[98]) & (i_10_) & (!i_11_) & (!i_15_)) + ((!i_8_) & (i_9_) & (!sk[98]) & (i_10_) & (!i_11_) & (i_15_)) + ((!i_8_) & (i_9_) & (!sk[98]) & (i_10_) & (i_11_) & (!i_15_)) + ((!i_8_) & (i_9_) & (!sk[98]) & (i_10_) & (i_11_) & (i_15_)) + ((i_8_) & (!i_9_) & (!sk[98]) & (i_10_) & (!i_11_) & (i_15_)) + ((i_8_) & (!i_9_) & (!sk[98]) & (i_10_) & (i_11_) & (!i_15_)) + ((i_8_) & (!i_9_) & (!sk[98]) & (i_10_) & (i_11_) & (i_15_)) + ((i_8_) & (i_9_) & (!sk[98]) & (!i_10_) & (!i_11_) & (!i_15_)) + ((i_8_) & (i_9_) & (!sk[98]) & (!i_10_) & (!i_11_) & (i_15_)) + ((i_8_) & (i_9_) & (!sk[98]) & (!i_10_) & (i_11_) & (!i_15_)) + ((i_8_) & (i_9_) & (!sk[98]) & (!i_10_) & (i_11_) & (i_15_)) + ((i_8_) & (i_9_) & (!sk[98]) & (i_10_) & (!i_11_) & (!i_15_)) + ((i_8_) & (i_9_) & (!sk[98]) & (i_10_) & (!i_11_) & (i_15_)) + ((i_8_) & (i_9_) & (!sk[98]) & (i_10_) & (i_11_) & (!i_15_)) + ((i_8_) & (i_9_) & (!sk[98]) & (i_10_) & (i_11_) & (i_15_)) + ((i_8_) & (i_9_) & (sk[98]) & (i_10_) & (!i_11_) & (!i_15_)));
	assign g325 = (((!sk[99]) & (!g68) & (!g165) & (g324)) + ((!sk[99]) & (!g68) & (g165) & (!g324)) + ((!sk[99]) & (!g68) & (g165) & (g324)) + ((!sk[99]) & (g68) & (!g165) & (g324)) + ((!sk[99]) & (g68) & (g165) & (!g324)) + ((!sk[99]) & (g68) & (g165) & (g324)) + ((sk[99]) & (!g68) & (g165) & (g324)));
	assign g326 = (((!i_9_) & (!i_10_) & (!sk[100]) & (i_11_) & (!i_15_) & (g68)) + ((!i_9_) & (!i_10_) & (!sk[100]) & (i_11_) & (i_15_) & (!g68)) + ((!i_9_) & (!i_10_) & (!sk[100]) & (i_11_) & (i_15_) & (g68)) + ((!i_9_) & (i_10_) & (!sk[100]) & (!i_11_) & (!i_15_) & (!g68)) + ((!i_9_) & (i_10_) & (!sk[100]) & (!i_11_) & (!i_15_) & (g68)) + ((!i_9_) & (i_10_) & (!sk[100]) & (!i_11_) & (i_15_) & (!g68)) + ((!i_9_) & (i_10_) & (!sk[100]) & (!i_11_) & (i_15_) & (g68)) + ((!i_9_) & (i_10_) & (!sk[100]) & (i_11_) & (!i_15_) & (!g68)) + ((!i_9_) & (i_10_) & (!sk[100]) & (i_11_) & (!i_15_) & (g68)) + ((!i_9_) & (i_10_) & (!sk[100]) & (i_11_) & (i_15_) & (!g68)) + ((!i_9_) & (i_10_) & (!sk[100]) & (i_11_) & (i_15_) & (g68)) + ((!i_9_) & (i_10_) & (sk[100]) & (!i_11_) & (!i_15_) & (!g68)) + ((!i_9_) & (i_10_) & (sk[100]) & (i_11_) & (!i_15_) & (!g68)) + ((i_9_) & (!i_10_) & (!sk[100]) & (i_11_) & (!i_15_) & (g68)) + ((i_9_) & (!i_10_) & (!sk[100]) & (i_11_) & (i_15_) & (!g68)) + ((i_9_) & (!i_10_) & (!sk[100]) & (i_11_) & (i_15_) & (g68)) + ((i_9_) & (!i_10_) & (sk[100]) & (i_11_) & (!i_15_) & (!g68)) + ((i_9_) & (i_10_) & (!sk[100]) & (!i_11_) & (!i_15_) & (!g68)) + ((i_9_) & (i_10_) & (!sk[100]) & (!i_11_) & (!i_15_) & (g68)) + ((i_9_) & (i_10_) & (!sk[100]) & (!i_11_) & (i_15_) & (!g68)) + ((i_9_) & (i_10_) & (!sk[100]) & (!i_11_) & (i_15_) & (g68)) + ((i_9_) & (i_10_) & (!sk[100]) & (i_11_) & (!i_15_) & (!g68)) + ((i_9_) & (i_10_) & (!sk[100]) & (i_11_) & (!i_15_) & (g68)) + ((i_9_) & (i_10_) & (!sk[100]) & (i_11_) & (i_15_) & (!g68)) + ((i_9_) & (i_10_) & (!sk[100]) & (i_11_) & (i_15_) & (g68)));
	assign g327 = (((!i_8_) & (!g24) & (g35) & (!g73) & (!sk[101]) & (g107)) + ((!i_8_) & (!g24) & (g35) & (g73) & (!sk[101]) & (!g107)) + ((!i_8_) & (!g24) & (g35) & (g73) & (!sk[101]) & (g107)) + ((!i_8_) & (g24) & (!g35) & (!g73) & (!sk[101]) & (!g107)) + ((!i_8_) & (g24) & (!g35) & (!g73) & (!sk[101]) & (g107)) + ((!i_8_) & (g24) & (!g35) & (g73) & (!sk[101]) & (!g107)) + ((!i_8_) & (g24) & (!g35) & (g73) & (!sk[101]) & (g107)) + ((!i_8_) & (g24) & (g35) & (!g73) & (!sk[101]) & (!g107)) + ((!i_8_) & (g24) & (g35) & (!g73) & (!sk[101]) & (g107)) + ((!i_8_) & (g24) & (g35) & (g73) & (!sk[101]) & (!g107)) + ((!i_8_) & (g24) & (g35) & (g73) & (!sk[101]) & (g107)) + ((i_8_) & (!g24) & (!g35) & (g73) & (sk[101]) & (!g107)) + ((i_8_) & (!g24) & (g35) & (!g73) & (!sk[101]) & (g107)) + ((i_8_) & (!g24) & (g35) & (g73) & (!sk[101]) & (!g107)) + ((i_8_) & (!g24) & (g35) & (g73) & (!sk[101]) & (g107)) + ((i_8_) & (!g24) & (g35) & (g73) & (sk[101]) & (!g107)) + ((i_8_) & (!g24) & (g35) & (g73) & (sk[101]) & (g107)) + ((i_8_) & (g24) & (!g35) & (!g73) & (!sk[101]) & (!g107)) + ((i_8_) & (g24) & (!g35) & (!g73) & (!sk[101]) & (g107)) + ((i_8_) & (g24) & (!g35) & (g73) & (!sk[101]) & (!g107)) + ((i_8_) & (g24) & (!g35) & (g73) & (!sk[101]) & (g107)) + ((i_8_) & (g24) & (g35) & (!g73) & (!sk[101]) & (!g107)) + ((i_8_) & (g24) & (g35) & (!g73) & (!sk[101]) & (g107)) + ((i_8_) & (g24) & (g35) & (g73) & (!sk[101]) & (!g107)) + ((i_8_) & (g24) & (g35) & (g73) & (!sk[101]) & (g107)));
	assign g328 = (((!g125) & (!g105) & (!g272) & (!g326) & (sk[102]) & (!g327)) + ((!g125) & (!g105) & (g272) & (!g326) & (!sk[102]) & (g327)) + ((!g125) & (!g105) & (g272) & (!g326) & (sk[102]) & (!g327)) + ((!g125) & (!g105) & (g272) & (g326) & (!sk[102]) & (!g327)) + ((!g125) & (!g105) & (g272) & (g326) & (!sk[102]) & (g327)) + ((!g125) & (g105) & (!g272) & (!g326) & (!sk[102]) & (!g327)) + ((!g125) & (g105) & (!g272) & (!g326) & (!sk[102]) & (g327)) + ((!g125) & (g105) & (!g272) & (!g326) & (sk[102]) & (!g327)) + ((!g125) & (g105) & (!g272) & (g326) & (!sk[102]) & (!g327)) + ((!g125) & (g105) & (!g272) & (g326) & (!sk[102]) & (g327)) + ((!g125) & (g105) & (!g272) & (g326) & (sk[102]) & (!g327)) + ((!g125) & (g105) & (g272) & (!g326) & (!sk[102]) & (!g327)) + ((!g125) & (g105) & (g272) & (!g326) & (!sk[102]) & (g327)) + ((!g125) & (g105) & (g272) & (!g326) & (sk[102]) & (!g327)) + ((!g125) & (g105) & (g272) & (g326) & (!sk[102]) & (!g327)) + ((!g125) & (g105) & (g272) & (g326) & (!sk[102]) & (g327)) + ((!g125) & (g105) & (g272) & (g326) & (sk[102]) & (!g327)) + ((g125) & (!g105) & (!g272) & (!g326) & (sk[102]) & (!g327)) + ((g125) & (!g105) & (g272) & (!g326) & (!sk[102]) & (g327)) + ((g125) & (!g105) & (g272) & (g326) & (!sk[102]) & (!g327)) + ((g125) & (!g105) & (g272) & (g326) & (!sk[102]) & (g327)) + ((g125) & (g105) & (!g272) & (!g326) & (!sk[102]) & (!g327)) + ((g125) & (g105) & (!g272) & (!g326) & (!sk[102]) & (g327)) + ((g125) & (g105) & (!g272) & (!g326) & (sk[102]) & (!g327)) + ((g125) & (g105) & (!g272) & (g326) & (!sk[102]) & (!g327)) + ((g125) & (g105) & (!g272) & (g326) & (!sk[102]) & (g327)) + ((g125) & (g105) & (!g272) & (g326) & (sk[102]) & (!g327)) + ((g125) & (g105) & (g272) & (!g326) & (!sk[102]) & (!g327)) + ((g125) & (g105) & (g272) & (!g326) & (!sk[102]) & (g327)) + ((g125) & (g105) & (g272) & (g326) & (!sk[102]) & (!g327)) + ((g125) & (g105) & (g272) & (g326) & (!sk[102]) & (g327)));
	assign g329 = (((!g25) & (!g102) & (g123) & (!g275) & (!g325) & (g328)) + ((!g25) & (!g102) & (g123) & (g275) & (!g325) & (g328)) + ((!g25) & (g102) & (g123) & (!g275) & (!g325) & (g328)) + ((g25) & (!g102) & (!g123) & (!g275) & (!g325) & (g328)) + ((g25) & (!g102) & (!g123) & (g275) & (!g325) & (g328)) + ((g25) & (!g102) & (g123) & (!g275) & (!g325) & (g328)) + ((g25) & (!g102) & (g123) & (g275) & (!g325) & (g328)) + ((g25) & (g102) & (!g123) & (!g275) & (!g325) & (g328)) + ((g25) & (g102) & (g123) & (!g275) & (!g325) & (g328)));
	assign g330 = (((!g24) & (!g35) & (!sk[104]) & (g157) & (!g74) & (g155)) + ((!g24) & (!g35) & (!sk[104]) & (g157) & (g74) & (!g155)) + ((!g24) & (!g35) & (!sk[104]) & (g157) & (g74) & (g155)) + ((!g24) & (g35) & (!sk[104]) & (!g157) & (!g74) & (!g155)) + ((!g24) & (g35) & (!sk[104]) & (!g157) & (!g74) & (g155)) + ((!g24) & (g35) & (!sk[104]) & (!g157) & (g74) & (!g155)) + ((!g24) & (g35) & (!sk[104]) & (!g157) & (g74) & (g155)) + ((!g24) & (g35) & (!sk[104]) & (g157) & (!g74) & (!g155)) + ((!g24) & (g35) & (!sk[104]) & (g157) & (!g74) & (g155)) + ((!g24) & (g35) & (!sk[104]) & (g157) & (g74) & (!g155)) + ((!g24) & (g35) & (!sk[104]) & (g157) & (g74) & (g155)) + ((!g24) & (g35) & (sk[104]) & (!g157) & (!g74) & (!g155)) + ((!g24) & (g35) & (sk[104]) & (!g157) & (g74) & (!g155)) + ((!g24) & (g35) & (sk[104]) & (!g157) & (g74) & (g155)) + ((!g24) & (g35) & (sk[104]) & (g157) & (!g74) & (!g155)) + ((!g24) & (g35) & (sk[104]) & (g157) & (!g74) & (g155)) + ((!g24) & (g35) & (sk[104]) & (g157) & (g74) & (!g155)) + ((!g24) & (g35) & (sk[104]) & (g157) & (g74) & (g155)) + ((g24) & (!g35) & (!sk[104]) & (g157) & (!g74) & (g155)) + ((g24) & (!g35) & (!sk[104]) & (g157) & (g74) & (!g155)) + ((g24) & (!g35) & (!sk[104]) & (g157) & (g74) & (g155)) + ((g24) & (g35) & (!sk[104]) & (!g157) & (!g74) & (!g155)) + ((g24) & (g35) & (!sk[104]) & (!g157) & (!g74) & (g155)) + ((g24) & (g35) & (!sk[104]) & (!g157) & (g74) & (!g155)) + ((g24) & (g35) & (!sk[104]) & (!g157) & (g74) & (g155)) + ((g24) & (g35) & (!sk[104]) & (g157) & (!g74) & (!g155)) + ((g24) & (g35) & (!sk[104]) & (g157) & (!g74) & (g155)) + ((g24) & (g35) & (!sk[104]) & (g157) & (g74) & (!g155)) + ((g24) & (g35) & (!sk[104]) & (g157) & (g74) & (g155)));
	assign g331 = (((!g125) & (!g168) & (!g121) & (!g270) & (!g330) & (g1606)) + ((!g125) & (!g168) & (!g121) & (g270) & (!g330) & (g1606)) + ((!g125) & (!g168) & (g121) & (!g270) & (!g330) & (g1606)) + ((!g125) & (g168) & (!g121) & (!g270) & (!g330) & (g1606)) + ((!g125) & (g168) & (g121) & (!g270) & (!g330) & (g1606)) + ((g125) & (!g168) & (!g121) & (!g270) & (!g330) & (g1606)) + ((g125) & (!g168) & (g121) & (!g270) & (!g330) & (g1606)) + ((g125) & (g168) & (!g121) & (!g270) & (!g330) & (g1606)) + ((g125) & (g168) & (g121) & (!g270) & (!g330) & (g1606)));
	assign g332 = (((!g285) & (!g322) & (g1613) & (!sk[106]) & (!g329) & (g331)) + ((!g285) & (!g322) & (g1613) & (!sk[106]) & (g329) & (!g331)) + ((!g285) & (!g322) & (g1613) & (!sk[106]) & (g329) & (g331)) + ((!g285) & (g322) & (!g1613) & (!sk[106]) & (!g329) & (!g331)) + ((!g285) & (g322) & (!g1613) & (!sk[106]) & (!g329) & (g331)) + ((!g285) & (g322) & (!g1613) & (!sk[106]) & (g329) & (!g331)) + ((!g285) & (g322) & (!g1613) & (!sk[106]) & (g329) & (g331)) + ((!g285) & (g322) & (g1613) & (!sk[106]) & (!g329) & (!g331)) + ((!g285) & (g322) & (g1613) & (!sk[106]) & (!g329) & (g331)) + ((!g285) & (g322) & (g1613) & (!sk[106]) & (g329) & (!g331)) + ((!g285) & (g322) & (g1613) & (!sk[106]) & (g329) & (g331)) + ((g285) & (!g322) & (g1613) & (!sk[106]) & (!g329) & (g331)) + ((g285) & (!g322) & (g1613) & (!sk[106]) & (g329) & (!g331)) + ((g285) & (!g322) & (g1613) & (!sk[106]) & (g329) & (g331)) + ((g285) & (g322) & (!g1613) & (!sk[106]) & (!g329) & (!g331)) + ((g285) & (g322) & (!g1613) & (!sk[106]) & (!g329) & (g331)) + ((g285) & (g322) & (!g1613) & (!sk[106]) & (g329) & (!g331)) + ((g285) & (g322) & (!g1613) & (!sk[106]) & (g329) & (g331)) + ((g285) & (g322) & (g1613) & (!sk[106]) & (!g329) & (!g331)) + ((g285) & (g322) & (g1613) & (!sk[106]) & (!g329) & (g331)) + ((g285) & (g322) & (g1613) & (!sk[106]) & (g329) & (!g331)) + ((g285) & (g322) & (g1613) & (!sk[106]) & (g329) & (g331)) + ((g285) & (g322) & (g1613) & (sk[106]) & (g329) & (g331)));
	assign g333 = (((!i_12_) & (!i_13_) & (i_14_) & (!sk[107]) & (!g20)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[107]) & (g20)) + ((!i_12_) & (!i_13_) & (i_14_) & (sk[107]) & (g20)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[107]) & (!g20)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[107]) & (g20)) + ((!i_12_) & (i_13_) & (i_14_) & (sk[107]) & (g20)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[107]) & (!g20)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[107]) & (g20)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[107]) & (!g20)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[107]) & (g20)) + ((i_12_) & (i_13_) & (i_14_) & (sk[107]) & (g20)));
	assign g334 = (((!g28) & (!sk[108]) & (!g98) & (g180)) + ((!g28) & (!sk[108]) & (g98) & (!g180)) + ((!g28) & (!sk[108]) & (g98) & (g180)) + ((!g28) & (sk[108]) & (!g98) & (!g180)) + ((g28) & (!sk[108]) & (!g98) & (g180)) + ((g28) & (!sk[108]) & (g98) & (!g180)) + ((g28) & (!sk[108]) & (g98) & (g180)));
	assign g335 = (((!sk[109]) & (!i_12_) & (!i_13_) & (i_14_) & (!g83)) + ((!sk[109]) & (!i_12_) & (!i_13_) & (i_14_) & (g83)) + ((!sk[109]) & (!i_12_) & (i_13_) & (i_14_) & (!g83)) + ((!sk[109]) & (!i_12_) & (i_13_) & (i_14_) & (g83)) + ((!sk[109]) & (i_12_) & (!i_13_) & (i_14_) & (!g83)) + ((!sk[109]) & (i_12_) & (!i_13_) & (i_14_) & (g83)) + ((!sk[109]) & (i_12_) & (i_13_) & (i_14_) & (!g83)) + ((!sk[109]) & (i_12_) & (i_13_) & (i_14_) & (g83)) + ((sk[109]) & (!i_12_) & (!i_13_) & (i_14_) & (g83)) + ((sk[109]) & (!i_12_) & (i_13_) & (i_14_) & (g83)) + ((sk[109]) & (i_12_) & (i_13_) & (i_14_) & (g83)));
	assign g336 = (((!sk[110]) & (!g87) & (!g191) & (g272)) + ((!sk[110]) & (!g87) & (g191) & (!g272)) + ((!sk[110]) & (!g87) & (g191) & (g272)) + ((!sk[110]) & (g87) & (!g191) & (g272)) + ((!sk[110]) & (g87) & (g191) & (!g272)) + ((!sk[110]) & (g87) & (g191) & (g272)) + ((sk[110]) & (g87) & (!g191) & (!g272)));
	assign g337 = (((g35) & (!sk[111]) & (!g176)) + ((g35) & (!sk[111]) & (g176)) + ((g35) & (sk[111]) & (!g176)));
	assign g338 = (((!i_12_) & (!i_13_) & (!sk[112]) & (i_14_) & (!g107)) + ((!i_12_) & (!i_13_) & (!sk[112]) & (i_14_) & (g107)) + ((!i_12_) & (!i_13_) & (sk[112]) & (i_14_) & (!g107)) + ((!i_12_) & (i_13_) & (!sk[112]) & (i_14_) & (!g107)) + ((!i_12_) & (i_13_) & (!sk[112]) & (i_14_) & (g107)) + ((!i_12_) & (i_13_) & (sk[112]) & (i_14_) & (!g107)) + ((i_12_) & (!i_13_) & (!sk[112]) & (i_14_) & (!g107)) + ((i_12_) & (!i_13_) & (!sk[112]) & (i_14_) & (g107)) + ((i_12_) & (i_13_) & (!sk[112]) & (i_14_) & (!g107)) + ((i_12_) & (i_13_) & (!sk[112]) & (i_14_) & (g107)) + ((i_12_) & (i_13_) & (sk[112]) & (i_14_) & (!g107)));
	assign g339 = (((!sk[113]) & (!i_12_) & (!i_13_) & (i_14_) & (!g35)) + ((!sk[113]) & (!i_12_) & (!i_13_) & (i_14_) & (g35)) + ((!sk[113]) & (!i_12_) & (i_13_) & (i_14_) & (!g35)) + ((!sk[113]) & (!i_12_) & (i_13_) & (i_14_) & (g35)) + ((!sk[113]) & (i_12_) & (!i_13_) & (i_14_) & (!g35)) + ((!sk[113]) & (i_12_) & (!i_13_) & (i_14_) & (g35)) + ((!sk[113]) & (i_12_) & (i_13_) & (i_14_) & (!g35)) + ((!sk[113]) & (i_12_) & (i_13_) & (i_14_) & (g35)) + ((sk[113]) & (!i_12_) & (!i_13_) & (i_14_) & (g35)) + ((sk[113]) & (!i_12_) & (i_13_) & (i_14_) & (g35)) + ((sk[113]) & (i_12_) & (i_13_) & (i_14_) & (g35)));
	assign g340 = (((!sk[114]) & (g83) & (!g176)) + ((!sk[114]) & (g83) & (g176)) + ((sk[114]) & (!g83) & (!g176)) + ((sk[114]) & (!g83) & (g176)) + ((sk[114]) & (g83) & (g176)));
	assign g341 = (((!sk[115]) & (!g77) & (!g188) & (g270)) + ((!sk[115]) & (!g77) & (g188) & (!g270)) + ((!sk[115]) & (!g77) & (g188) & (g270)) + ((!sk[115]) & (g77) & (!g188) & (g270)) + ((!sk[115]) & (g77) & (g188) & (!g270)) + ((!sk[115]) & (g77) & (g188) & (g270)) + ((sk[115]) & (!g77) & (!g188) & (!g270)));
	assign g342 = (((g86) & (!sk[116]) & (!g176)) + ((g86) & (!sk[116]) & (g176)) + ((g86) & (sk[116]) & (!g176)));
	assign g343 = (((!sk[117]) & (g20) & (!g176)) + ((!sk[117]) & (g20) & (g176)) + ((sk[117]) & (!g20) & (!g176)) + ((sk[117]) & (!g20) & (g176)) + ((sk[117]) & (g20) & (g176)));
	assign g344 = (((!sk[118]) & (!g164) & (!g340) & (g341) & (!g342) & (g343)) + ((!sk[118]) & (!g164) & (!g340) & (g341) & (g342) & (!g343)) + ((!sk[118]) & (!g164) & (!g340) & (g341) & (g342) & (g343)) + ((!sk[118]) & (!g164) & (g340) & (!g341) & (!g342) & (!g343)) + ((!sk[118]) & (!g164) & (g340) & (!g341) & (!g342) & (g343)) + ((!sk[118]) & (!g164) & (g340) & (!g341) & (g342) & (!g343)) + ((!sk[118]) & (!g164) & (g340) & (!g341) & (g342) & (g343)) + ((!sk[118]) & (!g164) & (g340) & (g341) & (!g342) & (!g343)) + ((!sk[118]) & (!g164) & (g340) & (g341) & (!g342) & (g343)) + ((!sk[118]) & (!g164) & (g340) & (g341) & (g342) & (!g343)) + ((!sk[118]) & (!g164) & (g340) & (g341) & (g342) & (g343)) + ((!sk[118]) & (g164) & (!g340) & (g341) & (!g342) & (g343)) + ((!sk[118]) & (g164) & (!g340) & (g341) & (g342) & (!g343)) + ((!sk[118]) & (g164) & (!g340) & (g341) & (g342) & (g343)) + ((!sk[118]) & (g164) & (g340) & (!g341) & (!g342) & (!g343)) + ((!sk[118]) & (g164) & (g340) & (!g341) & (!g342) & (g343)) + ((!sk[118]) & (g164) & (g340) & (!g341) & (g342) & (!g343)) + ((!sk[118]) & (g164) & (g340) & (!g341) & (g342) & (g343)) + ((!sk[118]) & (g164) & (g340) & (g341) & (!g342) & (!g343)) + ((!sk[118]) & (g164) & (g340) & (g341) & (!g342) & (g343)) + ((!sk[118]) & (g164) & (g340) & (g341) & (g342) & (!g343)) + ((!sk[118]) & (g164) & (g340) & (g341) & (g342) & (g343)) + ((sk[118]) & (g164) & (!g340) & (!g341) & (!g342) & (!g343)) + ((sk[118]) & (g164) & (!g340) & (!g341) & (!g342) & (g343)) + ((sk[118]) & (g164) & (!g340) & (!g341) & (g342) & (!g343)) + ((sk[118]) & (g164) & (!g340) & (!g341) & (g342) & (g343)) + ((sk[118]) & (g164) & (!g340) & (g341) & (!g342) & (!g343)) + ((sk[118]) & (g164) & (!g340) & (g341) & (!g342) & (g343)) + ((sk[118]) & (g164) & (!g340) & (g341) & (g342) & (!g343)) + ((sk[118]) & (g164) & (!g340) & (g341) & (g342) & (g343)) + ((sk[118]) & (g164) & (g340) & (!g341) & (!g342) & (!g343)) + ((sk[118]) & (g164) & (g340) & (!g341) & (!g342) & (g343)) + ((sk[118]) & (g164) & (g340) & (!g341) & (g342) & (!g343)) + ((sk[118]) & (g164) & (g340) & (!g341) & (g342) & (g343)) + ((sk[118]) & (g164) & (g340) & (g341) & (!g342) & (!g343)) + ((sk[118]) & (g164) & (g340) & (g341) & (g342) & (!g343)) + ((sk[118]) & (g164) & (g340) & (g341) & (g342) & (g343)));
	assign g345 = (((!g164) & (!g253) & (!g337) & (!g338) & (!g339) & (!g344)) + ((!g164) & (!g253) & (!g337) & (g338) & (!g339) & (!g344)) + ((!g164) & (g253) & (!g337) & (!g338) & (!g339) & (!g344)) + ((!g164) & (g253) & (!g337) & (!g338) & (g339) & (!g344)) + ((!g164) & (g253) & (!g337) & (g338) & (!g339) & (!g344)) + ((!g164) & (g253) & (!g337) & (g338) & (g339) & (!g344)) + ((!g164) & (g253) & (g337) & (!g338) & (!g339) & (!g344)) + ((!g164) & (g253) & (g337) & (!g338) & (g339) & (!g344)) + ((!g164) & (g253) & (g337) & (g338) & (!g339) & (!g344)) + ((!g164) & (g253) & (g337) & (g338) & (g339) & (!g344)) + ((g164) & (!g253) & (!g337) & (!g338) & (!g339) & (!g344)) + ((g164) & (g253) & (!g337) & (!g338) & (!g339) & (!g344)) + ((g164) & (g253) & (g337) & (!g338) & (!g339) & (!g344)));
	assign g346 = (((!g253) & (!g333) & (g334) & (!g335) & (g336) & (g345)) + ((g253) & (!g333) & (!g334) & (!g335) & (!g336) & (g345)) + ((g253) & (!g333) & (!g334) & (!g335) & (g336) & (g345)) + ((g253) & (!g333) & (!g334) & (g335) & (!g336) & (g345)) + ((g253) & (!g333) & (!g334) & (g335) & (g336) & (g345)) + ((g253) & (!g333) & (g334) & (!g335) & (!g336) & (g345)) + ((g253) & (!g333) & (g334) & (!g335) & (g336) & (g345)) + ((g253) & (!g333) & (g334) & (g335) & (!g336) & (g345)) + ((g253) & (!g333) & (g334) & (g335) & (g336) & (g345)) + ((g253) & (g333) & (!g334) & (!g335) & (!g336) & (g345)) + ((g253) & (g333) & (!g334) & (!g335) & (g336) & (g345)) + ((g253) & (g333) & (!g334) & (g335) & (!g336) & (g345)) + ((g253) & (g333) & (!g334) & (g335) & (g336) & (g345)) + ((g253) & (g333) & (g334) & (!g335) & (!g336) & (g345)) + ((g253) & (g333) & (g334) & (!g335) & (g336) & (g345)) + ((g253) & (g333) & (g334) & (g335) & (!g336) & (g345)) + ((g253) & (g333) & (g334) & (g335) & (g336) & (g345)));
	assign g347 = (((g154) & (!sk[121]) & (!g122)) + ((g154) & (!sk[121]) & (g122)) + ((g154) & (sk[121]) & (!g122)));
	assign g348 = (((!sk[122]) & (!i_8_) & (!g73) & (g130)) + ((!sk[122]) & (!i_8_) & (g73) & (!g130)) + ((!sk[122]) & (!i_8_) & (g73) & (g130)) + ((!sk[122]) & (i_8_) & (!g73) & (g130)) + ((!sk[122]) & (i_8_) & (g73) & (!g130)) + ((!sk[122]) & (i_8_) & (g73) & (g130)) + ((sk[122]) & (!i_8_) & (!g73) & (g130)) + ((sk[122]) & (i_8_) & (!g73) & (g130)) + ((sk[122]) & (i_8_) & (g73) & (g130)));
	assign g349 = (((!g144) & (!sk[123]) & (!g164) & (g347) & (!g105) & (g348)) + ((!g144) & (!sk[123]) & (!g164) & (g347) & (g105) & (!g348)) + ((!g144) & (!sk[123]) & (!g164) & (g347) & (g105) & (g348)) + ((!g144) & (!sk[123]) & (g164) & (!g347) & (!g105) & (!g348)) + ((!g144) & (!sk[123]) & (g164) & (!g347) & (!g105) & (g348)) + ((!g144) & (!sk[123]) & (g164) & (!g347) & (g105) & (!g348)) + ((!g144) & (!sk[123]) & (g164) & (!g347) & (g105) & (g348)) + ((!g144) & (!sk[123]) & (g164) & (g347) & (!g105) & (!g348)) + ((!g144) & (!sk[123]) & (g164) & (g347) & (!g105) & (g348)) + ((!g144) & (!sk[123]) & (g164) & (g347) & (g105) & (!g348)) + ((!g144) & (!sk[123]) & (g164) & (g347) & (g105) & (g348)) + ((!g144) & (sk[123]) & (!g164) & (g347) & (g105) & (g348)) + ((g144) & (!sk[123]) & (!g164) & (g347) & (!g105) & (g348)) + ((g144) & (!sk[123]) & (!g164) & (g347) & (g105) & (!g348)) + ((g144) & (!sk[123]) & (!g164) & (g347) & (g105) & (g348)) + ((g144) & (!sk[123]) & (g164) & (!g347) & (!g105) & (!g348)) + ((g144) & (!sk[123]) & (g164) & (!g347) & (!g105) & (g348)) + ((g144) & (!sk[123]) & (g164) & (!g347) & (g105) & (!g348)) + ((g144) & (!sk[123]) & (g164) & (!g347) & (g105) & (g348)) + ((g144) & (!sk[123]) & (g164) & (g347) & (!g105) & (!g348)) + ((g144) & (!sk[123]) & (g164) & (g347) & (!g105) & (g348)) + ((g144) & (!sk[123]) & (g164) & (g347) & (g105) & (!g348)) + ((g144) & (!sk[123]) & (g164) & (g347) & (g105) & (g348)));
	assign g350 = (((!i_8_) & (!i_6_) & (!i_7_) & (!g120) & (g166) & (!g118)) + ((!i_8_) & (!i_6_) & (!i_7_) & (!g120) & (g166) & (g118)) + ((!i_8_) & (!i_6_) & (!i_7_) & (g120) & (g166) & (!g118)) + ((!i_8_) & (!i_6_) & (!i_7_) & (g120) & (g166) & (g118)) + ((!i_8_) & (!i_6_) & (i_7_) & (g120) & (!g166) & (!g118)) + ((!i_8_) & (!i_6_) & (i_7_) & (g120) & (!g166) & (g118)) + ((!i_8_) & (!i_6_) & (i_7_) & (g120) & (g166) & (!g118)) + ((!i_8_) & (!i_6_) & (i_7_) & (g120) & (g166) & (g118)) + ((!i_8_) & (i_6_) & (!i_7_) & (!g120) & (g166) & (!g118)) + ((!i_8_) & (i_6_) & (!i_7_) & (!g120) & (g166) & (g118)) + ((!i_8_) & (i_6_) & (!i_7_) & (g120) & (g166) & (!g118)) + ((!i_8_) & (i_6_) & (!i_7_) & (g120) & (g166) & (g118)) + ((i_8_) & (!i_6_) & (!i_7_) & (!g120) & (g166) & (!g118)) + ((i_8_) & (!i_6_) & (!i_7_) & (!g120) & (g166) & (g118)) + ((i_8_) & (!i_6_) & (!i_7_) & (g120) & (g166) & (!g118)) + ((i_8_) & (!i_6_) & (!i_7_) & (g120) & (g166) & (g118)) + ((i_8_) & (!i_6_) & (i_7_) & (g120) & (!g166) & (!g118)) + ((i_8_) & (!i_6_) & (i_7_) & (g120) & (!g166) & (g118)) + ((i_8_) & (!i_6_) & (i_7_) & (g120) & (g166) & (!g118)) + ((i_8_) & (!i_6_) & (i_7_) & (g120) & (g166) & (g118)) + ((i_8_) & (i_6_) & (!i_7_) & (!g120) & (!g166) & (g118)) + ((i_8_) & (i_6_) & (!i_7_) & (!g120) & (g166) & (g118)) + ((i_8_) & (i_6_) & (!i_7_) & (g120) & (!g166) & (!g118)) + ((i_8_) & (i_6_) & (!i_7_) & (g120) & (!g166) & (g118)) + ((i_8_) & (i_6_) & (!i_7_) & (g120) & (g166) & (!g118)) + ((i_8_) & (i_6_) & (!i_7_) & (g120) & (g166) & (g118)));
	assign g351 = (((!i_7_) & (!g72) & (!sk[125]) & (g350)) + ((!i_7_) & (!g72) & (sk[125]) & (!g350)) + ((!i_7_) & (g72) & (!sk[125]) & (!g350)) + ((!i_7_) & (g72) & (!sk[125]) & (g350)) + ((!i_7_) & (g72) & (sk[125]) & (!g350)) + ((i_7_) & (!g72) & (!sk[125]) & (g350)) + ((i_7_) & (!g72) & (sk[125]) & (!g350)) + ((i_7_) & (g72) & (!sk[125]) & (!g350)) + ((i_7_) & (g72) & (!sk[125]) & (g350)));
	assign g352 = (((!g119) & (!g121) & (!g227) & (sk[126]) & (g351)) + ((!g119) & (!g121) & (g227) & (!sk[126]) & (!g351)) + ((!g119) & (!g121) & (g227) & (!sk[126]) & (g351)) + ((!g119) & (g121) & (g227) & (!sk[126]) & (!g351)) + ((!g119) & (g121) & (g227) & (!sk[126]) & (g351)) + ((g119) & (!g121) & (g227) & (!sk[126]) & (!g351)) + ((g119) & (!g121) & (g227) & (!sk[126]) & (g351)) + ((g119) & (g121) & (g227) & (!sk[126]) & (!g351)) + ((g119) & (g121) & (g227) & (!sk[126]) & (g351)));
	assign g353 = (((!i_11_) & (!i_15_) & (!sk[127]) & (g53)) + ((!i_11_) & (!i_15_) & (sk[127]) & (!g53)) + ((!i_11_) & (i_15_) & (!sk[127]) & (!g53)) + ((!i_11_) & (i_15_) & (!sk[127]) & (g53)) + ((i_11_) & (!i_15_) & (!sk[127]) & (g53)) + ((i_11_) & (i_15_) & (!sk[127]) & (!g53)) + ((i_11_) & (i_15_) & (!sk[127]) & (g53)));
	assign g354 = (((!g3) & (!g35) & (!g176) & (!g349) & (!g352) & (g353)) + ((!g3) & (g35) & (!g176) & (!g349) & (!g352) & (g353)) + ((!g3) & (g35) & (!g176) & (!g349) & (g352) & (g353)) + ((g3) & (!g35) & (!g176) & (!g349) & (!g352) & (g353)) + ((g3) & (!g35) & (!g176) & (g349) & (!g352) & (g353)) + ((g3) & (g35) & (!g176) & (!g349) & (!g352) & (g353)) + ((g3) & (g35) & (!g176) & (!g349) & (g352) & (g353)) + ((g3) & (g35) & (!g176) & (g349) & (!g352) & (g353)));
	assign g355 = (((!sk[1]) & (i_12_) & (!i_14_)) + ((!sk[1]) & (i_12_) & (i_14_)) + ((sk[1]) & (!i_12_) & (i_14_)));
	assign g356 = (((!g159) & (sk[2]) & (!g313)) + ((!g159) & (sk[2]) & (g313)) + ((g159) & (!sk[2]) & (!g313)) + ((g159) & (!sk[2]) & (g313)) + ((g159) & (sk[2]) & (g313)));
	assign g357 = (((!sk[3]) & (g27) & (!g176)) + ((!sk[3]) & (g27) & (g176)) + ((sk[3]) & (g27) & (!g176)));
	assign g358 = (((!g107) & (sk[4]) & (!g176)) + ((g107) & (!sk[4]) & (!g176)) + ((g107) & (!sk[4]) & (g176)));
	assign g359 = (((!g27) & (!g126) & (g102) & (!sk[5]) & (!g176)) + ((!g27) & (!g126) & (g102) & (!sk[5]) & (g176)) + ((!g27) & (!g126) & (g102) & (sk[5]) & (!g176)) + ((!g27) & (g126) & (g102) & (!sk[5]) & (!g176)) + ((!g27) & (g126) & (g102) & (!sk[5]) & (g176)) + ((g27) & (!g126) & (g102) & (!sk[5]) & (!g176)) + ((g27) & (!g126) & (g102) & (!sk[5]) & (g176)) + ((g27) & (!g126) & (g102) & (sk[5]) & (!g176)) + ((g27) & (g126) & (g102) & (!sk[5]) & (!g176)) + ((g27) & (g126) & (g102) & (!sk[5]) & (g176)) + ((g27) & (g126) & (g102) & (sk[5]) & (!g176)));
	assign g360 = (((!g105) & (!g342) & (!g358) & (sk[6]) & (!g359)) + ((!g105) & (!g342) & (g358) & (!sk[6]) & (!g359)) + ((!g105) & (!g342) & (g358) & (!sk[6]) & (g359)) + ((!g105) & (g342) & (g358) & (!sk[6]) & (!g359)) + ((!g105) & (g342) & (g358) & (!sk[6]) & (g359)) + ((g105) & (!g342) & (!g358) & (sk[6]) & (!g359)) + ((g105) & (!g342) & (g358) & (!sk[6]) & (!g359)) + ((g105) & (!g342) & (g358) & (!sk[6]) & (g359)) + ((g105) & (!g342) & (g358) & (sk[6]) & (!g359)) + ((g105) & (g342) & (!g358) & (sk[6]) & (!g359)) + ((g105) & (g342) & (g358) & (!sk[6]) & (!g359)) + ((g105) & (g342) & (g358) & (!sk[6]) & (g359)) + ((g105) & (g342) & (g358) & (sk[6]) & (!g359)));
	assign g361 = (((!g355) & (!g83) & (!g356) & (!g357) & (!g350) & (g360)) + ((!g355) & (!g83) & (!g356) & (!g357) & (g350) & (g360)) + ((!g355) & (!g83) & (!g356) & (g357) & (!g350) & (g360)) + ((!g355) & (!g83) & (g356) & (!g357) & (!g350) & (g360)) + ((!g355) & (!g83) & (g356) & (!g357) & (g350) & (g360)) + ((!g355) & (!g83) & (g356) & (g357) & (!g350) & (g360)) + ((!g355) & (g83) & (!g356) & (!g357) & (!g350) & (g360)) + ((!g355) & (g83) & (!g356) & (!g357) & (g350) & (g360)) + ((!g355) & (g83) & (!g356) & (g357) & (!g350) & (g360)) + ((!g355) & (g83) & (g356) & (!g357) & (!g350) & (g360)) + ((!g355) & (g83) & (g356) & (!g357) & (g350) & (g360)) + ((!g355) & (g83) & (g356) & (g357) & (!g350) & (g360)) + ((g355) & (!g83) & (!g356) & (!g357) & (!g350) & (g360)) + ((g355) & (!g83) & (!g356) & (!g357) & (g350) & (g360)) + ((g355) & (!g83) & (!g356) & (g357) & (!g350) & (g360)) + ((g355) & (!g83) & (g356) & (!g357) & (!g350) & (g360)) + ((g355) & (!g83) & (g356) & (!g357) & (g350) & (g360)) + ((g355) & (!g83) & (g356) & (g357) & (!g350) & (g360)) + ((g355) & (g83) & (!g356) & (!g357) & (!g350) & (g360)) + ((g355) & (g83) & (!g356) & (!g357) & (g350) & (g360)) + ((g355) & (g83) & (!g356) & (g357) & (!g350) & (g360)));
	assign g362 = (((!g154) & (!sk[8]) & (!g340) & (g335)) + ((!g154) & (!sk[8]) & (g340) & (!g335)) + ((!g154) & (!sk[8]) & (g340) & (g335)) + ((!g154) & (sk[8]) & (!g340) & (!g335)) + ((!g154) & (sk[8]) & (!g340) & (g335)) + ((!g154) & (sk[8]) & (g340) & (g335)) + ((g154) & (!sk[8]) & (!g340) & (g335)) + ((g154) & (!sk[8]) & (g340) & (!g335)) + ((g154) & (!sk[8]) & (g340) & (g335)));
	assign g363 = (((!g159) & (!sk[9]) & (!g154) & (g333) & (!g343)) + ((!g159) & (!sk[9]) & (!g154) & (g333) & (g343)) + ((!g159) & (!sk[9]) & (g154) & (g333) & (!g343)) + ((!g159) & (!sk[9]) & (g154) & (g333) & (g343)) + ((!g159) & (sk[9]) & (!g154) & (!g333) & (g343)) + ((!g159) & (sk[9]) & (g154) & (!g333) & (!g343)) + ((!g159) & (sk[9]) & (g154) & (!g333) & (g343)) + ((g159) & (!sk[9]) & (!g154) & (g333) & (!g343)) + ((g159) & (!sk[9]) & (!g154) & (g333) & (g343)) + ((g159) & (!sk[9]) & (g154) & (g333) & (!g343)) + ((g159) & (!sk[9]) & (g154) & (g333) & (g343)) + ((g159) & (sk[9]) & (!g154) & (!g333) & (g343)) + ((g159) & (sk[9]) & (g154) & (!g333) & (!g343)) + ((g159) & (sk[9]) & (g154) & (!g333) & (g343)) + ((g159) & (sk[9]) & (g154) & (g333) & (!g343)) + ((g159) & (sk[9]) & (g154) & (g333) & (g343)));
	assign g364 = (((!g159) & (!sk[10]) & (!g154) & (g337) & (!g334) & (g339)) + ((!g159) & (!sk[10]) & (!g154) & (g337) & (g334) & (!g339)) + ((!g159) & (!sk[10]) & (!g154) & (g337) & (g334) & (g339)) + ((!g159) & (!sk[10]) & (g154) & (!g337) & (!g334) & (!g339)) + ((!g159) & (!sk[10]) & (g154) & (!g337) & (!g334) & (g339)) + ((!g159) & (!sk[10]) & (g154) & (!g337) & (g334) & (!g339)) + ((!g159) & (!sk[10]) & (g154) & (!g337) & (g334) & (g339)) + ((!g159) & (!sk[10]) & (g154) & (g337) & (!g334) & (!g339)) + ((!g159) & (!sk[10]) & (g154) & (g337) & (!g334) & (g339)) + ((!g159) & (!sk[10]) & (g154) & (g337) & (g334) & (!g339)) + ((!g159) & (!sk[10]) & (g154) & (g337) & (g334) & (g339)) + ((!g159) & (sk[10]) & (!g154) & (!g337) & (g334) & (!g339)) + ((!g159) & (sk[10]) & (g154) & (!g337) & (g334) & (!g339)) + ((g159) & (!sk[10]) & (!g154) & (g337) & (!g334) & (g339)) + ((g159) & (!sk[10]) & (!g154) & (g337) & (g334) & (!g339)) + ((g159) & (!sk[10]) & (!g154) & (g337) & (g334) & (g339)) + ((g159) & (!sk[10]) & (g154) & (!g337) & (!g334) & (!g339)) + ((g159) & (!sk[10]) & (g154) & (!g337) & (!g334) & (g339)) + ((g159) & (!sk[10]) & (g154) & (!g337) & (g334) & (!g339)) + ((g159) & (!sk[10]) & (g154) & (!g337) & (g334) & (g339)) + ((g159) & (!sk[10]) & (g154) & (g337) & (!g334) & (!g339)) + ((g159) & (!sk[10]) & (g154) & (g337) & (!g334) & (g339)) + ((g159) & (!sk[10]) & (g154) & (g337) & (g334) & (!g339)) + ((g159) & (!sk[10]) & (g154) & (g337) & (g334) & (g339)) + ((g159) & (sk[10]) & (!g154) & (!g337) & (g334) & (!g339)) + ((g159) & (sk[10]) & (!g154) & (!g337) & (g334) & (g339)) + ((g159) & (sk[10]) & (!g154) & (g337) & (g334) & (!g339)) + ((g159) & (sk[10]) & (!g154) & (g337) & (g334) & (g339)) + ((g159) & (sk[10]) & (g154) & (!g337) & (!g334) & (!g339)) + ((g159) & (sk[10]) & (g154) & (!g337) & (!g334) & (g339)) + ((g159) & (sk[10]) & (g154) & (!g337) & (g334) & (!g339)) + ((g159) & (sk[10]) & (g154) & (!g337) & (g334) & (g339)) + ((g159) & (sk[10]) & (g154) & (g337) & (!g334) & (!g339)) + ((g159) & (sk[10]) & (g154) & (g337) & (!g334) & (g339)) + ((g159) & (sk[10]) & (g154) & (g337) & (g334) & (!g339)) + ((g159) & (sk[10]) & (g154) & (g337) & (g334) & (g339)));
	assign g365 = (((!g154) & (!g342) & (g336) & (!g362) & (g363) & (g364)) + ((g154) & (!g342) & (!g336) & (!g362) & (g363) & (g364)) + ((g154) & (!g342) & (g336) & (!g362) & (g363) & (g364)) + ((g154) & (g342) & (!g336) & (!g362) & (g363) & (g364)) + ((g154) & (g342) & (g336) & (!g362) & (g363) & (g364)));
	assign g366 = (((!g102) & (!g186) & (!sk[12]) & (g296) & (!g358)) + ((!g102) & (!g186) & (!sk[12]) & (g296) & (g358)) + ((!g102) & (g186) & (!sk[12]) & (g296) & (!g358)) + ((!g102) & (g186) & (!sk[12]) & (g296) & (g358)) + ((g102) & (!g186) & (!sk[12]) & (g296) & (!g358)) + ((g102) & (!g186) & (!sk[12]) & (g296) & (g358)) + ((g102) & (!g186) & (sk[12]) & (!g296) & (g358)) + ((g102) & (!g186) & (sk[12]) & (g296) & (!g358)) + ((g102) & (!g186) & (sk[12]) & (g296) & (g358)) + ((g102) & (g186) & (!sk[12]) & (g296) & (!g358)) + ((g102) & (g186) & (!sk[12]) & (g296) & (g358)) + ((g102) & (g186) & (sk[12]) & (!g296) & (!g358)) + ((g102) & (g186) & (sk[12]) & (!g296) & (g358)) + ((g102) & (g186) & (sk[12]) & (g296) & (!g358)) + ((g102) & (g186) & (sk[12]) & (g296) & (g358)));
	assign g367 = (((!g108) & (!g105) & (!g212) & (sk[13]) & (g309)) + ((!g108) & (!g105) & (g212) & (!sk[13]) & (!g309)) + ((!g108) & (!g105) & (g212) & (!sk[13]) & (g309)) + ((!g108) & (!g105) & (g212) & (sk[13]) & (!g309)) + ((!g108) & (!g105) & (g212) & (sk[13]) & (g309)) + ((!g108) & (g105) & (g212) & (!sk[13]) & (!g309)) + ((!g108) & (g105) & (g212) & (!sk[13]) & (g309)) + ((g108) & (!g105) & (!g212) & (sk[13]) & (!g309)) + ((g108) & (!g105) & (!g212) & (sk[13]) & (g309)) + ((g108) & (!g105) & (g212) & (!sk[13]) & (!g309)) + ((g108) & (!g105) & (g212) & (!sk[13]) & (g309)) + ((g108) & (!g105) & (g212) & (sk[13]) & (!g309)) + ((g108) & (!g105) & (g212) & (sk[13]) & (g309)) + ((g108) & (g105) & (g212) & (!sk[13]) & (!g309)) + ((g108) & (g105) & (g212) & (!sk[13]) & (g309)));
	assign g368 = (((!g123) & (!g185) & (!g187) & (sk[14]) & (g337)) + ((!g123) & (!g185) & (g187) & (!sk[14]) & (!g337)) + ((!g123) & (!g185) & (g187) & (!sk[14]) & (g337)) + ((!g123) & (!g185) & (g187) & (sk[14]) & (!g337)) + ((!g123) & (!g185) & (g187) & (sk[14]) & (g337)) + ((!g123) & (g185) & (!g187) & (sk[14]) & (!g337)) + ((!g123) & (g185) & (!g187) & (sk[14]) & (g337)) + ((!g123) & (g185) & (g187) & (!sk[14]) & (!g337)) + ((!g123) & (g185) & (g187) & (!sk[14]) & (g337)) + ((!g123) & (g185) & (g187) & (sk[14]) & (!g337)) + ((!g123) & (g185) & (g187) & (sk[14]) & (g337)) + ((g123) & (!g185) & (g187) & (!sk[14]) & (!g337)) + ((g123) & (!g185) & (g187) & (!sk[14]) & (g337)) + ((g123) & (g185) & (g187) & (!sk[14]) & (!g337)) + ((g123) & (g185) & (g187) & (!sk[14]) & (g337)));
	assign g369 = (((!i_12_) & (!i_13_) & (!sk[15]) & (i_14_) & (!g126)) + ((!i_12_) & (!i_13_) & (!sk[15]) & (i_14_) & (g126)) + ((!i_12_) & (!i_13_) & (sk[15]) & (i_14_) & (!g126)) + ((!i_12_) & (i_13_) & (!sk[15]) & (i_14_) & (!g126)) + ((!i_12_) & (i_13_) & (!sk[15]) & (i_14_) & (g126)) + ((!i_12_) & (i_13_) & (sk[15]) & (i_14_) & (!g126)) + ((i_12_) & (!i_13_) & (!sk[15]) & (i_14_) & (!g126)) + ((i_12_) & (!i_13_) & (!sk[15]) & (i_14_) & (g126)) + ((i_12_) & (i_13_) & (!sk[15]) & (i_14_) & (!g126)) + ((i_12_) & (i_13_) & (!sk[15]) & (i_14_) & (g126)) + ((i_12_) & (i_13_) & (sk[15]) & (i_14_) & (!g126)));
	assign g370 = (((!g253) & (!g369) & (!sk[16]) & (g338) & (!g358)) + ((!g253) & (!g369) & (!sk[16]) & (g338) & (g358)) + ((!g253) & (!g369) & (sk[16]) & (!g338) & (g358)) + ((!g253) & (!g369) & (sk[16]) & (g338) & (!g358)) + ((!g253) & (!g369) & (sk[16]) & (g338) & (g358)) + ((!g253) & (g369) & (!sk[16]) & (g338) & (!g358)) + ((!g253) & (g369) & (!sk[16]) & (g338) & (g358)) + ((!g253) & (g369) & (sk[16]) & (!g338) & (!g358)) + ((!g253) & (g369) & (sk[16]) & (!g338) & (g358)) + ((!g253) & (g369) & (sk[16]) & (g338) & (!g358)) + ((!g253) & (g369) & (sk[16]) & (g338) & (g358)) + ((g253) & (!g369) & (!sk[16]) & (g338) & (!g358)) + ((g253) & (!g369) & (!sk[16]) & (g338) & (g358)) + ((g253) & (g369) & (!sk[16]) & (g338) & (!g358)) + ((g253) & (g369) & (!sk[16]) & (g338) & (g358)));
	assign g371 = (((!g135) & (!g122) & (!g131) & (sk[17]) & (g342)) + ((!g135) & (!g122) & (g131) & (!sk[17]) & (!g342)) + ((!g135) & (!g122) & (g131) & (!sk[17]) & (g342)) + ((!g135) & (!g122) & (g131) & (sk[17]) & (g342)) + ((!g135) & (g122) & (!g131) & (sk[17]) & (g342)) + ((!g135) & (g122) & (g131) & (!sk[17]) & (!g342)) + ((!g135) & (g122) & (g131) & (!sk[17]) & (g342)) + ((!g135) & (g122) & (g131) & (sk[17]) & (g342)) + ((g135) & (!g122) & (!g131) & (sk[17]) & (g342)) + ((g135) & (!g122) & (g131) & (!sk[17]) & (!g342)) + ((g135) & (!g122) & (g131) & (!sk[17]) & (g342)) + ((g135) & (g122) & (!g131) & (sk[17]) & (g342)) + ((g135) & (g122) & (g131) & (!sk[17]) & (!g342)) + ((g135) & (g122) & (g131) & (!sk[17]) & (g342)) + ((g135) & (g122) & (g131) & (sk[17]) & (g342)));
	assign g372 = (((!sk[18]) & (!g123) & (!g130) & (g342) & (!g358)) + ((!sk[18]) & (!g123) & (!g130) & (g342) & (g358)) + ((!sk[18]) & (!g123) & (g130) & (g342) & (!g358)) + ((!sk[18]) & (!g123) & (g130) & (g342) & (g358)) + ((!sk[18]) & (g123) & (!g130) & (g342) & (!g358)) + ((!sk[18]) & (g123) & (!g130) & (g342) & (g358)) + ((!sk[18]) & (g123) & (g130) & (g342) & (!g358)) + ((!sk[18]) & (g123) & (g130) & (g342) & (g358)) + ((sk[18]) & (!g123) & (!g130) & (!g342) & (!g358)) + ((sk[18]) & (!g123) & (g130) & (!g342) & (!g358)) + ((sk[18]) & (!g123) & (g130) & (!g342) & (g358)) + ((sk[18]) & (g123) & (!g130) & (!g342) & (!g358)) + ((sk[18]) & (g123) & (g130) & (!g342) & (!g358)) + ((sk[18]) & (g123) & (g130) & (!g342) & (g358)) + ((sk[18]) & (g123) & (g130) & (g342) & (!g358)) + ((sk[18]) & (g123) & (g130) & (g342) & (g358)));
	assign g373 = (((!sk[19]) & (!g367) & (!g368) & (g370) & (!g371) & (g372)) + ((!sk[19]) & (!g367) & (!g368) & (g370) & (g371) & (!g372)) + ((!sk[19]) & (!g367) & (!g368) & (g370) & (g371) & (g372)) + ((!sk[19]) & (!g367) & (g368) & (!g370) & (!g371) & (!g372)) + ((!sk[19]) & (!g367) & (g368) & (!g370) & (!g371) & (g372)) + ((!sk[19]) & (!g367) & (g368) & (!g370) & (g371) & (!g372)) + ((!sk[19]) & (!g367) & (g368) & (!g370) & (g371) & (g372)) + ((!sk[19]) & (!g367) & (g368) & (g370) & (!g371) & (!g372)) + ((!sk[19]) & (!g367) & (g368) & (g370) & (!g371) & (g372)) + ((!sk[19]) & (!g367) & (g368) & (g370) & (g371) & (!g372)) + ((!sk[19]) & (!g367) & (g368) & (g370) & (g371) & (g372)) + ((!sk[19]) & (g367) & (!g368) & (g370) & (!g371) & (g372)) + ((!sk[19]) & (g367) & (!g368) & (g370) & (g371) & (!g372)) + ((!sk[19]) & (g367) & (!g368) & (g370) & (g371) & (g372)) + ((!sk[19]) & (g367) & (g368) & (!g370) & (!g371) & (!g372)) + ((!sk[19]) & (g367) & (g368) & (!g370) & (!g371) & (g372)) + ((!sk[19]) & (g367) & (g368) & (!g370) & (g371) & (!g372)) + ((!sk[19]) & (g367) & (g368) & (!g370) & (g371) & (g372)) + ((!sk[19]) & (g367) & (g368) & (g370) & (!g371) & (!g372)) + ((!sk[19]) & (g367) & (g368) & (g370) & (!g371) & (g372)) + ((!sk[19]) & (g367) & (g368) & (g370) & (g371) & (!g372)) + ((!sk[19]) & (g367) & (g368) & (g370) & (g371) & (g372)) + ((sk[19]) & (!g367) & (!g368) & (!g370) & (!g371) & (g372)));
	assign g374 = (((!g161) & (!g157) & (!sk[20]) & (g337) & (!g343)) + ((!g161) & (!g157) & (!sk[20]) & (g337) & (g343)) + ((!g161) & (!g157) & (sk[20]) & (!g337) & (!g343)) + ((!g161) & (!g157) & (sk[20]) & (!g337) & (g343)) + ((!g161) & (!g157) & (sk[20]) & (g337) & (!g343)) + ((!g161) & (!g157) & (sk[20]) & (g337) & (g343)) + ((!g161) & (g157) & (!sk[20]) & (g337) & (!g343)) + ((!g161) & (g157) & (!sk[20]) & (g337) & (g343)) + ((!g161) & (g157) & (sk[20]) & (!g337) & (!g343)) + ((!g161) & (g157) & (sk[20]) & (!g337) & (g343)) + ((g161) & (!g157) & (!sk[20]) & (g337) & (!g343)) + ((g161) & (!g157) & (!sk[20]) & (g337) & (g343)) + ((g161) & (!g157) & (sk[20]) & (!g337) & (g343)) + ((g161) & (g157) & (!sk[20]) & (g337) & (!g343)) + ((g161) & (g157) & (!sk[20]) & (g337) & (g343)) + ((g161) & (g157) & (sk[20]) & (!g337) & (g343)));
	assign g375 = (((!i_8_) & (!g73) & (!sk[21]) & (g192) & (!g212)) + ((!i_8_) & (!g73) & (!sk[21]) & (g192) & (g212)) + ((!i_8_) & (g73) & (!sk[21]) & (g192) & (!g212)) + ((!i_8_) & (g73) & (!sk[21]) & (g192) & (g212)) + ((i_8_) & (!g73) & (!sk[21]) & (g192) & (!g212)) + ((i_8_) & (!g73) & (!sk[21]) & (g192) & (g212)) + ((i_8_) & (g73) & (!sk[21]) & (g192) & (!g212)) + ((i_8_) & (g73) & (!sk[21]) & (g192) & (g212)) + ((i_8_) & (g73) & (sk[21]) & (!g192) & (g212)) + ((i_8_) & (g73) & (sk[21]) & (g192) & (!g212)) + ((i_8_) & (g73) & (sk[21]) & (g192) & (g212)));
	assign g376 = (((!g125) & (!g191) & (!sk[22]) & (g192) & (!g212)) + ((!g125) & (!g191) & (!sk[22]) & (g192) & (g212)) + ((!g125) & (g191) & (!sk[22]) & (g192) & (!g212)) + ((!g125) & (g191) & (!sk[22]) & (g192) & (g212)) + ((g125) & (!g191) & (!sk[22]) & (g192) & (!g212)) + ((g125) & (!g191) & (!sk[22]) & (g192) & (g212)) + ((g125) & (!g191) & (sk[22]) & (!g192) & (g212)) + ((g125) & (!g191) & (sk[22]) & (g192) & (!g212)) + ((g125) & (!g191) & (sk[22]) & (g192) & (g212)) + ((g125) & (g191) & (!sk[22]) & (g192) & (!g212)) + ((g125) & (g191) & (!sk[22]) & (g192) & (g212)) + ((g125) & (g191) & (sk[22]) & (!g192) & (!g212)) + ((g125) & (g191) & (sk[22]) & (!g192) & (g212)) + ((g125) & (g191) & (sk[22]) & (g192) & (!g212)) + ((g125) & (g191) & (sk[22]) & (g192) & (g212)));
	assign g377 = (((!sk[23]) & (!i_8_) & (!g73) & (g102) & (!g337)) + ((!sk[23]) & (!i_8_) & (!g73) & (g102) & (g337)) + ((!sk[23]) & (!i_8_) & (g73) & (g102) & (!g337)) + ((!sk[23]) & (!i_8_) & (g73) & (g102) & (g337)) + ((!sk[23]) & (i_8_) & (!g73) & (g102) & (!g337)) + ((!sk[23]) & (i_8_) & (!g73) & (g102) & (g337)) + ((!sk[23]) & (i_8_) & (g73) & (g102) & (!g337)) + ((!sk[23]) & (i_8_) & (g73) & (g102) & (g337)) + ((sk[23]) & (!i_8_) & (!g73) & (g102) & (g337)) + ((sk[23]) & (!i_8_) & (g73) & (g102) & (g337)) + ((sk[23]) & (i_8_) & (!g73) & (g102) & (g337)) + ((sk[23]) & (i_8_) & (g73) & (!g102) & (g337)) + ((sk[23]) & (i_8_) & (g73) & (g102) & (g337)));
	assign g378 = (((!g102) & (!g105) & (!g186) & (!g182) & (!g295) & (!g281)) + ((!g102) & (g105) & (!g186) & (!g182) & (!g295) & (!g281)) + ((!g102) & (g105) & (!g186) & (!g182) & (!g295) & (g281)) + ((!g102) & (g105) & (!g186) & (!g182) & (g295) & (!g281)) + ((!g102) & (g105) & (!g186) & (!g182) & (g295) & (g281)) + ((!g102) & (g105) & (!g186) & (g182) & (!g295) & (!g281)) + ((!g102) & (g105) & (!g186) & (g182) & (!g295) & (g281)) + ((!g102) & (g105) & (!g186) & (g182) & (g295) & (!g281)) + ((!g102) & (g105) & (!g186) & (g182) & (g295) & (g281)) + ((!g102) & (g105) & (g186) & (!g182) & (!g295) & (!g281)) + ((!g102) & (g105) & (g186) & (!g182) & (!g295) & (g281)) + ((!g102) & (g105) & (g186) & (!g182) & (g295) & (!g281)) + ((!g102) & (g105) & (g186) & (!g182) & (g295) & (g281)) + ((!g102) & (g105) & (g186) & (g182) & (!g295) & (!g281)) + ((!g102) & (g105) & (g186) & (g182) & (!g295) & (g281)) + ((!g102) & (g105) & (g186) & (g182) & (g295) & (!g281)) + ((!g102) & (g105) & (g186) & (g182) & (g295) & (g281)) + ((g102) & (!g105) & (!g186) & (!g182) & (!g295) & (!g281)) + ((g102) & (g105) & (!g186) & (!g182) & (!g295) & (!g281)) + ((g102) & (g105) & (!g186) & (!g182) & (g295) & (!g281)) + ((g102) & (g105) & (!g186) & (g182) & (!g295) & (!g281)) + ((g102) & (g105) & (!g186) & (g182) & (g295) & (!g281)) + ((g102) & (g105) & (g186) & (!g182) & (!g295) & (!g281)) + ((g102) & (g105) & (g186) & (!g182) & (g295) & (!g281)) + ((g102) & (g105) & (g186) & (g182) & (!g295) & (!g281)) + ((g102) & (g105) & (g186) & (g182) & (g295) & (!g281)));
	assign g379 = (((!sk[25]) & (!g374) & (!g375) & (g376) & (!g377) & (g378)) + ((!sk[25]) & (!g374) & (!g375) & (g376) & (g377) & (!g378)) + ((!sk[25]) & (!g374) & (!g375) & (g376) & (g377) & (g378)) + ((!sk[25]) & (!g374) & (g375) & (!g376) & (!g377) & (!g378)) + ((!sk[25]) & (!g374) & (g375) & (!g376) & (!g377) & (g378)) + ((!sk[25]) & (!g374) & (g375) & (!g376) & (g377) & (!g378)) + ((!sk[25]) & (!g374) & (g375) & (!g376) & (g377) & (g378)) + ((!sk[25]) & (!g374) & (g375) & (g376) & (!g377) & (!g378)) + ((!sk[25]) & (!g374) & (g375) & (g376) & (!g377) & (g378)) + ((!sk[25]) & (!g374) & (g375) & (g376) & (g377) & (!g378)) + ((!sk[25]) & (!g374) & (g375) & (g376) & (g377) & (g378)) + ((!sk[25]) & (g374) & (!g375) & (g376) & (!g377) & (g378)) + ((!sk[25]) & (g374) & (!g375) & (g376) & (g377) & (!g378)) + ((!sk[25]) & (g374) & (!g375) & (g376) & (g377) & (g378)) + ((!sk[25]) & (g374) & (g375) & (!g376) & (!g377) & (!g378)) + ((!sk[25]) & (g374) & (g375) & (!g376) & (!g377) & (g378)) + ((!sk[25]) & (g374) & (g375) & (!g376) & (g377) & (!g378)) + ((!sk[25]) & (g374) & (g375) & (!g376) & (g377) & (g378)) + ((!sk[25]) & (g374) & (g375) & (g376) & (!g377) & (!g378)) + ((!sk[25]) & (g374) & (g375) & (g376) & (!g377) & (g378)) + ((!sk[25]) & (g374) & (g375) & (g376) & (g377) & (!g378)) + ((!sk[25]) & (g374) & (g375) & (g376) & (g377) & (g378)) + ((sk[25]) & (g374) & (!g375) & (!g376) & (!g377) & (g378)));
	assign g380 = (((!g164) & (!sk[26]) & (!g123) & (g333) & (!g335)) + ((!g164) & (!sk[26]) & (!g123) & (g333) & (g335)) + ((!g164) & (!sk[26]) & (g123) & (g333) & (!g335)) + ((!g164) & (!sk[26]) & (g123) & (g333) & (g335)) + ((!g164) & (sk[26]) & (!g123) & (!g333) & (!g335)) + ((!g164) & (sk[26]) & (!g123) & (g333) & (!g335)) + ((!g164) & (sk[26]) & (g123) & (!g333) & (!g335)) + ((!g164) & (sk[26]) & (g123) & (!g333) & (g335)) + ((!g164) & (sk[26]) & (g123) & (g333) & (!g335)) + ((!g164) & (sk[26]) & (g123) & (g333) & (g335)) + ((g164) & (!sk[26]) & (!g123) & (g333) & (!g335)) + ((g164) & (!sk[26]) & (!g123) & (g333) & (g335)) + ((g164) & (!sk[26]) & (g123) & (g333) & (!g335)) + ((g164) & (!sk[26]) & (g123) & (g333) & (g335)) + ((g164) & (sk[26]) & (!g123) & (!g333) & (!g335)) + ((g164) & (sk[26]) & (g123) & (!g333) & (!g335)));
	assign g381 = (((!sk[27]) & (!g226) & (!g227) & (g275) & (!g357) & (g334)) + ((!sk[27]) & (!g226) & (!g227) & (g275) & (g357) & (!g334)) + ((!sk[27]) & (!g226) & (!g227) & (g275) & (g357) & (g334)) + ((!sk[27]) & (!g226) & (g227) & (!g275) & (!g357) & (!g334)) + ((!sk[27]) & (!g226) & (g227) & (!g275) & (!g357) & (g334)) + ((!sk[27]) & (!g226) & (g227) & (!g275) & (g357) & (!g334)) + ((!sk[27]) & (!g226) & (g227) & (!g275) & (g357) & (g334)) + ((!sk[27]) & (!g226) & (g227) & (g275) & (!g357) & (!g334)) + ((!sk[27]) & (!g226) & (g227) & (g275) & (!g357) & (g334)) + ((!sk[27]) & (!g226) & (g227) & (g275) & (g357) & (!g334)) + ((!sk[27]) & (!g226) & (g227) & (g275) & (g357) & (g334)) + ((!sk[27]) & (g226) & (!g227) & (g275) & (!g357) & (g334)) + ((!sk[27]) & (g226) & (!g227) & (g275) & (g357) & (!g334)) + ((!sk[27]) & (g226) & (!g227) & (g275) & (g357) & (g334)) + ((!sk[27]) & (g226) & (g227) & (!g275) & (!g357) & (!g334)) + ((!sk[27]) & (g226) & (g227) & (!g275) & (!g357) & (g334)) + ((!sk[27]) & (g226) & (g227) & (!g275) & (g357) & (!g334)) + ((!sk[27]) & (g226) & (g227) & (!g275) & (g357) & (g334)) + ((!sk[27]) & (g226) & (g227) & (g275) & (!g357) & (!g334)) + ((!sk[27]) & (g226) & (g227) & (g275) & (!g357) & (g334)) + ((!sk[27]) & (g226) & (g227) & (g275) & (g357) & (!g334)) + ((!sk[27]) & (g226) & (g227) & (g275) & (g357) & (g334)) + ((sk[27]) & (!g226) & (!g227) & (!g275) & (!g357) & (g334)) + ((sk[27]) & (!g226) & (!g227) & (!g275) & (g357) & (g334)) + ((sk[27]) & (!g226) & (g227) & (!g275) & (!g357) & (g334)) + ((sk[27]) & (g226) & (!g227) & (!g275) & (!g357) & (!g334)) + ((sk[27]) & (g226) & (!g227) & (!g275) & (!g357) & (g334)) + ((sk[27]) & (g226) & (!g227) & (!g275) & (g357) & (!g334)) + ((sk[27]) & (g226) & (!g227) & (!g275) & (g357) & (g334)) + ((sk[27]) & (g226) & (!g227) & (g275) & (!g357) & (!g334)) + ((sk[27]) & (g226) & (!g227) & (g275) & (!g357) & (g334)) + ((sk[27]) & (g226) & (!g227) & (g275) & (g357) & (!g334)) + ((sk[27]) & (g226) & (!g227) & (g275) & (g357) & (g334)) + ((sk[27]) & (g226) & (g227) & (!g275) & (!g357) & (g334)) + ((sk[27]) & (g226) & (g227) & (g275) & (!g357) & (g334)));
	assign g382 = (((!g164) & (!g225) & (!g334) & (!g336) & (g380) & (g381)) + ((!g164) & (!g225) & (!g334) & (g336) & (g380) & (g381)) + ((!g164) & (!g225) & (g334) & (!g336) & (g380) & (g381)) + ((!g164) & (!g225) & (g334) & (g336) & (g380) & (g381)) + ((!g164) & (g225) & (g334) & (!g336) & (g380) & (g381)) + ((!g164) & (g225) & (g334) & (g336) & (g380) & (g381)) + ((g164) & (!g225) & (g334) & (g336) & (g380) & (g381)) + ((g164) & (g225) & (g334) & (g336) & (g380) & (g381)));
	assign g383 = (((!sk[29]) & (g125) & (!g254)) + ((!sk[29]) & (g125) & (g254)) + ((sk[29]) & (!g125) & (g254)));
	assign g384 = (((!g142) & (!g257) & (g179) & (!g254) & (!sk[30]) & (g217)) + ((!g142) & (!g257) & (g179) & (!g254) & (sk[30]) & (!g217)) + ((!g142) & (!g257) & (g179) & (!g254) & (sk[30]) & (g217)) + ((!g142) & (!g257) & (g179) & (g254) & (!sk[30]) & (!g217)) + ((!g142) & (!g257) & (g179) & (g254) & (!sk[30]) & (g217)) + ((!g142) & (!g257) & (g179) & (g254) & (sk[30]) & (!g217)) + ((!g142) & (!g257) & (g179) & (g254) & (sk[30]) & (g217)) + ((!g142) & (g257) & (!g179) & (!g254) & (!sk[30]) & (!g217)) + ((!g142) & (g257) & (!g179) & (!g254) & (!sk[30]) & (g217)) + ((!g142) & (g257) & (!g179) & (g254) & (!sk[30]) & (!g217)) + ((!g142) & (g257) & (!g179) & (g254) & (!sk[30]) & (g217)) + ((!g142) & (g257) & (g179) & (!g254) & (!sk[30]) & (!g217)) + ((!g142) & (g257) & (g179) & (!g254) & (!sk[30]) & (g217)) + ((!g142) & (g257) & (g179) & (!g254) & (sk[30]) & (!g217)) + ((!g142) & (g257) & (g179) & (!g254) & (sk[30]) & (g217)) + ((!g142) & (g257) & (g179) & (g254) & (!sk[30]) & (!g217)) + ((!g142) & (g257) & (g179) & (g254) & (!sk[30]) & (g217)) + ((!g142) & (g257) & (g179) & (g254) & (sk[30]) & (!g217)) + ((!g142) & (g257) & (g179) & (g254) & (sk[30]) & (g217)) + ((g142) & (!g257) & (g179) & (!g254) & (!sk[30]) & (g217)) + ((g142) & (!g257) & (g179) & (!g254) & (sk[30]) & (!g217)) + ((g142) & (!g257) & (g179) & (!g254) & (sk[30]) & (g217)) + ((g142) & (!g257) & (g179) & (g254) & (!sk[30]) & (!g217)) + ((g142) & (!g257) & (g179) & (g254) & (!sk[30]) & (g217)) + ((g142) & (!g257) & (g179) & (g254) & (sk[30]) & (g217)) + ((g142) & (g257) & (!g179) & (!g254) & (!sk[30]) & (!g217)) + ((g142) & (g257) & (!g179) & (!g254) & (!sk[30]) & (g217)) + ((g142) & (g257) & (!g179) & (g254) & (!sk[30]) & (!g217)) + ((g142) & (g257) & (!g179) & (g254) & (!sk[30]) & (g217)) + ((g142) & (g257) & (g179) & (!g254) & (!sk[30]) & (!g217)) + ((g142) & (g257) & (g179) & (!g254) & (!sk[30]) & (g217)) + ((g142) & (g257) & (g179) & (!g254) & (sk[30]) & (!g217)) + ((g142) & (g257) & (g179) & (!g254) & (sk[30]) & (g217)) + ((g142) & (g257) & (g179) & (g254) & (!sk[30]) & (!g217)) + ((g142) & (g257) & (g179) & (g254) & (!sk[30]) & (g217)) + ((g142) & (g257) & (g179) & (g254) & (sk[30]) & (!g217)) + ((g142) & (g257) & (g179) & (g254) & (sk[30]) & (g217)));
	assign g385 = (((!sk[31]) & (!i_8_) & (!g73) & (g357) & (!g358)) + ((!sk[31]) & (!i_8_) & (!g73) & (g357) & (g358)) + ((!sk[31]) & (!i_8_) & (g73) & (g357) & (!g358)) + ((!sk[31]) & (!i_8_) & (g73) & (g357) & (g358)) + ((!sk[31]) & (i_8_) & (!g73) & (g357) & (!g358)) + ((!sk[31]) & (i_8_) & (!g73) & (g357) & (g358)) + ((!sk[31]) & (i_8_) & (g73) & (g357) & (!g358)) + ((!sk[31]) & (i_8_) & (g73) & (g357) & (g358)) + ((sk[31]) & (!i_8_) & (g73) & (!g357) & (g358)) + ((sk[31]) & (!i_8_) & (g73) & (g357) & (g358)) + ((sk[31]) & (i_8_) & (g73) & (!g357) & (g358)) + ((sk[31]) & (i_8_) & (g73) & (g357) & (!g358)) + ((sk[31]) & (i_8_) & (g73) & (g357) & (g358)));
	assign g386 = (((!g347) & (!g356) & (!g383) & (!g384) & (!g358) & (!g385)) + ((!g347) & (!g356) & (g383) & (!g384) & (!g358) & (!g385)) + ((!g347) & (g356) & (!g383) & (!g384) & (!g358) & (!g385)) + ((!g347) & (g356) & (g383) & (!g384) & (!g358) & (!g385)) + ((g347) & (!g356) & (!g383) & (!g384) & (!g358) & (!g385)) + ((g347) & (!g356) & (g383) & (!g384) & (!g358) & (!g385)) + ((g347) & (!g356) & (g383) & (!g384) & (g358) & (!g385)) + ((g347) & (g356) & (!g383) & (!g384) & (!g358) & (!g385)) + ((g347) & (g356) & (g383) & (!g384) & (!g358) & (!g385)));
	assign g387 = (((g365) & (!g366) & (g373) & (g379) & (g382) & (g386)));
	assign g388 = (((!i_12_) & (i_13_) & (i_14_) & (g20) & (!g157) & (!g130)) + ((!i_12_) & (i_13_) & (i_14_) & (g20) & (g157) & (!g130)) + ((i_12_) & (!i_13_) & (i_14_) & (g20) & (g157) & (!g130)) + ((i_12_) & (!i_13_) & (i_14_) & (g20) & (g157) & (g130)));
	assign g389 = (((!g3) & (!g176) & (!sk[35]) & (g226) & (!g341)) + ((!g3) & (!g176) & (!sk[35]) & (g226) & (g341)) + ((!g3) & (!g176) & (sk[35]) & (!g226) & (!g341)) + ((!g3) & (g176) & (!sk[35]) & (g226) & (!g341)) + ((!g3) & (g176) & (!sk[35]) & (g226) & (g341)) + ((!g3) & (g176) & (sk[35]) & (!g226) & (!g341)) + ((g3) & (!g176) & (!sk[35]) & (g226) & (!g341)) + ((g3) & (!g176) & (!sk[35]) & (g226) & (g341)) + ((g3) & (!g176) & (sk[35]) & (!g226) & (!g341)) + ((g3) & (!g176) & (sk[35]) & (!g226) & (g341)) + ((g3) & (g176) & (!sk[35]) & (g226) & (!g341)) + ((g3) & (g176) & (!sk[35]) & (g226) & (g341)) + ((g3) & (g176) & (sk[35]) & (!g226) & (!g341)));
	assign g390 = (((!g20) & (!g126) & (!g122) & (!g123) & (!g105) & (!g176)) + ((!g20) & (!g126) & (!g122) & (!g123) & (g105) & (!g176)) + ((!g20) & (!g126) & (!g122) & (g123) & (!g105) & (!g176)) + ((!g20) & (!g126) & (g122) & (!g123) & (!g105) & (!g176)) + ((!g20) & (!g126) & (g122) & (!g123) & (g105) & (!g176)) + ((!g20) & (!g126) & (g122) & (g123) & (!g105) & (!g176)) + ((g20) & (!g126) & (!g122) & (!g123) & (!g105) & (!g176)) + ((g20) & (!g126) & (!g122) & (!g123) & (g105) & (!g176)) + ((g20) & (!g126) & (!g122) & (g123) & (!g105) & (!g176)) + ((g20) & (!g126) & (g122) & (!g123) & (!g105) & (!g176)) + ((g20) & (!g126) & (g122) & (!g123) & (g105) & (!g176)) + ((g20) & (!g126) & (g122) & (g123) & (!g105) & (!g176)) + ((g20) & (!g126) & (g122) & (g123) & (g105) & (!g176)) + ((g20) & (g126) & (!g122) & (!g123) & (!g105) & (!g176)) + ((g20) & (g126) & (!g122) & (g123) & (!g105) & (!g176)) + ((g20) & (g126) & (g122) & (!g123) & (!g105) & (!g176)) + ((g20) & (g126) & (g122) & (!g123) & (g105) & (!g176)) + ((g20) & (g126) & (g122) & (g123) & (!g105) & (!g176)) + ((g20) & (g126) & (g122) & (g123) & (g105) & (!g176)));
	assign g391 = (((!g125) & (!g126) & (!g176) & (sk[37]) & (!g389) & (!g390)) + ((!g125) & (!g126) & (g176) & (!sk[37]) & (!g389) & (g390)) + ((!g125) & (!g126) & (g176) & (!sk[37]) & (g389) & (!g390)) + ((!g125) & (!g126) & (g176) & (!sk[37]) & (g389) & (g390)) + ((!g125) & (!g126) & (g176) & (sk[37]) & (!g389) & (!g390)) + ((!g125) & (g126) & (!g176) & (!sk[37]) & (!g389) & (!g390)) + ((!g125) & (g126) & (!g176) & (!sk[37]) & (!g389) & (g390)) + ((!g125) & (g126) & (!g176) & (!sk[37]) & (g389) & (!g390)) + ((!g125) & (g126) & (!g176) & (!sk[37]) & (g389) & (g390)) + ((!g125) & (g126) & (!g176) & (sk[37]) & (!g389) & (!g390)) + ((!g125) & (g126) & (g176) & (!sk[37]) & (!g389) & (!g390)) + ((!g125) & (g126) & (g176) & (!sk[37]) & (!g389) & (g390)) + ((!g125) & (g126) & (g176) & (!sk[37]) & (g389) & (!g390)) + ((!g125) & (g126) & (g176) & (!sk[37]) & (g389) & (g390)) + ((!g125) & (g126) & (g176) & (sk[37]) & (!g389) & (!g390)) + ((g125) & (!g126) & (g176) & (!sk[37]) & (!g389) & (g390)) + ((g125) & (!g126) & (g176) & (!sk[37]) & (g389) & (!g390)) + ((g125) & (!g126) & (g176) & (!sk[37]) & (g389) & (g390)) + ((g125) & (!g126) & (g176) & (sk[37]) & (!g389) & (!g390)) + ((g125) & (g126) & (!g176) & (!sk[37]) & (!g389) & (!g390)) + ((g125) & (g126) & (!g176) & (!sk[37]) & (!g389) & (g390)) + ((g125) & (g126) & (!g176) & (!sk[37]) & (g389) & (!g390)) + ((g125) & (g126) & (!g176) & (!sk[37]) & (g389) & (g390)) + ((g125) & (g126) & (!g176) & (sk[37]) & (!g389) & (!g390)) + ((g125) & (g126) & (g176) & (!sk[37]) & (!g389) & (!g390)) + ((g125) & (g126) & (g176) & (!sk[37]) & (!g389) & (g390)) + ((g125) & (g126) & (g176) & (!sk[37]) & (g389) & (!g390)) + ((g125) & (g126) & (g176) & (!sk[37]) & (g389) & (g390)) + ((g125) & (g126) & (g176) & (sk[37]) & (!g389) & (!g390)));
	assign g392 = (((g42) & (!sk[38]) & (!g72)) + ((g42) & (!sk[38]) & (g72)) + ((g42) & (sk[38]) & (g72)));
	assign g393 = (((!g102) & (!sk[39]) & (!g191) & (g273) & (!g392)) + ((!g102) & (!sk[39]) & (!g191) & (g273) & (g392)) + ((!g102) & (!sk[39]) & (g191) & (g273) & (!g392)) + ((!g102) & (!sk[39]) & (g191) & (g273) & (g392)) + ((!g102) & (sk[39]) & (g191) & (!g273) & (g392)) + ((!g102) & (sk[39]) & (g191) & (g273) & (g392)) + ((g102) & (!sk[39]) & (!g191) & (g273) & (!g392)) + ((g102) & (!sk[39]) & (!g191) & (g273) & (g392)) + ((g102) & (!sk[39]) & (g191) & (g273) & (!g392)) + ((g102) & (!sk[39]) & (g191) & (g273) & (g392)) + ((g102) & (sk[39]) & (!g191) & (g273) & (!g392)) + ((g102) & (sk[39]) & (!g191) & (g273) & (g392)) + ((g102) & (sk[39]) & (g191) & (!g273) & (g392)) + ((g102) & (sk[39]) & (g191) & (g273) & (!g392)) + ((g102) & (sk[39]) & (g191) & (g273) & (g392)));
	assign g394 = (((!sk[40]) & (g15) & (!g71)) + ((!sk[40]) & (g15) & (g71)) + ((sk[40]) & (g15) & (g71)));
	assign g395 = (((!i_6_) & (!i_7_) & (i_10_) & (!sk[41]) & (!i_11_) & (g394)) + ((!i_6_) & (!i_7_) & (i_10_) & (!sk[41]) & (i_11_) & (!g394)) + ((!i_6_) & (!i_7_) & (i_10_) & (!sk[41]) & (i_11_) & (g394)) + ((!i_6_) & (i_7_) & (!i_10_) & (!sk[41]) & (!i_11_) & (!g394)) + ((!i_6_) & (i_7_) & (!i_10_) & (!sk[41]) & (!i_11_) & (g394)) + ((!i_6_) & (i_7_) & (!i_10_) & (!sk[41]) & (i_11_) & (!g394)) + ((!i_6_) & (i_7_) & (!i_10_) & (!sk[41]) & (i_11_) & (g394)) + ((!i_6_) & (i_7_) & (i_10_) & (!sk[41]) & (!i_11_) & (!g394)) + ((!i_6_) & (i_7_) & (i_10_) & (!sk[41]) & (!i_11_) & (g394)) + ((!i_6_) & (i_7_) & (i_10_) & (!sk[41]) & (i_11_) & (!g394)) + ((!i_6_) & (i_7_) & (i_10_) & (!sk[41]) & (i_11_) & (g394)) + ((!i_6_) & (i_7_) & (i_10_) & (sk[41]) & (!i_11_) & (g394)) + ((i_6_) & (!i_7_) & (i_10_) & (!sk[41]) & (!i_11_) & (g394)) + ((i_6_) & (!i_7_) & (i_10_) & (!sk[41]) & (i_11_) & (!g394)) + ((i_6_) & (!i_7_) & (i_10_) & (!sk[41]) & (i_11_) & (g394)) + ((i_6_) & (!i_7_) & (i_10_) & (sk[41]) & (!i_11_) & (g394)) + ((i_6_) & (i_7_) & (!i_10_) & (!sk[41]) & (!i_11_) & (!g394)) + ((i_6_) & (i_7_) & (!i_10_) & (!sk[41]) & (!i_11_) & (g394)) + ((i_6_) & (i_7_) & (!i_10_) & (!sk[41]) & (i_11_) & (!g394)) + ((i_6_) & (i_7_) & (!i_10_) & (!sk[41]) & (i_11_) & (g394)) + ((i_6_) & (i_7_) & (i_10_) & (!sk[41]) & (!i_11_) & (!g394)) + ((i_6_) & (i_7_) & (i_10_) & (!sk[41]) & (!i_11_) & (g394)) + ((i_6_) & (i_7_) & (i_10_) & (!sk[41]) & (i_11_) & (!g394)) + ((i_6_) & (i_7_) & (i_10_) & (!sk[41]) & (i_11_) & (g394)));
	assign g396 = (((!sk[42]) & (!g142) & (!g333) & (g395)) + ((!sk[42]) & (!g142) & (g333) & (!g395)) + ((!sk[42]) & (!g142) & (g333) & (g395)) + ((!sk[42]) & (g142) & (!g333) & (g395)) + ((!sk[42]) & (g142) & (g333) & (!g395)) + ((!sk[42]) & (g142) & (g333) & (g395)) + ((sk[42]) & (!g142) & (!g333) & (!g395)) + ((sk[42]) & (g142) & (!g333) & (!g395)) + ((sk[42]) & (g142) & (g333) & (!g395)));
	assign g397 = (((g355) & (!sk[43]) & (!g126)) + ((g355) & (!sk[43]) & (g126)) + ((g355) & (sk[43]) & (!g126)));
	assign g398 = (((!i_14_) & (!g125) & (!g154) & (!g122) & (!g83) & (g397)) + ((!i_14_) & (!g125) & (!g154) & (!g122) & (g83) & (g397)) + ((!i_14_) & (!g125) & (!g154) & (g122) & (!g83) & (g397)) + ((!i_14_) & (!g125) & (!g154) & (g122) & (g83) & (g397)) + ((!i_14_) & (!g125) & (g154) & (g122) & (!g83) & (g397)) + ((!i_14_) & (!g125) & (g154) & (g122) & (g83) & (g397)) + ((!i_14_) & (g125) & (!g154) & (!g122) & (!g83) & (g397)) + ((!i_14_) & (g125) & (!g154) & (!g122) & (g83) & (g397)) + ((!i_14_) & (g125) & (!g154) & (g122) & (!g83) & (g397)) + ((!i_14_) & (g125) & (!g154) & (g122) & (g83) & (g397)) + ((!i_14_) & (g125) & (g154) & (g122) & (!g83) & (g397)) + ((!i_14_) & (g125) & (g154) & (g122) & (g83) & (g397)) + ((i_14_) & (!g125) & (!g154) & (!g122) & (!g83) & (g397)) + ((i_14_) & (!g125) & (!g154) & (!g122) & (g83) & (g397)) + ((i_14_) & (!g125) & (!g154) & (g122) & (!g83) & (g397)) + ((i_14_) & (!g125) & (!g154) & (g122) & (g83) & (g397)) + ((i_14_) & (!g125) & (g154) & (g122) & (!g83) & (g397)) + ((i_14_) & (!g125) & (g154) & (g122) & (g83) & (g397)) + ((i_14_) & (g125) & (!g154) & (!g122) & (!g83) & (g397)) + ((i_14_) & (g125) & (!g154) & (!g122) & (g83) & (!g397)) + ((i_14_) & (g125) & (!g154) & (!g122) & (g83) & (g397)) + ((i_14_) & (g125) & (!g154) & (g122) & (!g83) & (g397)) + ((i_14_) & (g125) & (!g154) & (g122) & (g83) & (!g397)) + ((i_14_) & (g125) & (!g154) & (g122) & (g83) & (g397)) + ((i_14_) & (g125) & (g154) & (!g122) & (g83) & (!g397)) + ((i_14_) & (g125) & (g154) & (!g122) & (g83) & (g397)) + ((i_14_) & (g125) & (g154) & (g122) & (!g83) & (g397)) + ((i_14_) & (g125) & (g154) & (g122) & (g83) & (!g397)) + ((i_14_) & (g125) & (g154) & (g122) & (g83) & (g397)));
	assign g399 = (((!g135) & (!g123) & (!g186) & (!g227) & (!g341) & (!g337)) + ((!g135) & (!g123) & (!g186) & (!g227) & (g341) & (!g337)) + ((!g135) & (!g123) & (!g186) & (g227) & (g341) & (!g337)) + ((!g135) & (g123) & (!g186) & (!g227) & (!g341) & (!g337)) + ((!g135) & (g123) & (!g186) & (!g227) & (g341) & (!g337)) + ((!g135) & (g123) & (!g186) & (g227) & (g341) & (!g337)) + ((!g135) & (g123) & (g186) & (!g227) & (!g341) & (!g337)) + ((!g135) & (g123) & (g186) & (!g227) & (g341) & (!g337)) + ((!g135) & (g123) & (g186) & (g227) & (g341) & (!g337)) + ((g135) & (!g123) & (!g186) & (!g227) & (!g341) & (!g337)) + ((g135) & (!g123) & (!g186) & (!g227) & (!g341) & (g337)) + ((g135) & (!g123) & (!g186) & (!g227) & (g341) & (!g337)) + ((g135) & (!g123) & (!g186) & (!g227) & (g341) & (g337)) + ((g135) & (!g123) & (!g186) & (g227) & (g341) & (!g337)) + ((g135) & (!g123) & (!g186) & (g227) & (g341) & (g337)) + ((g135) & (g123) & (!g186) & (!g227) & (!g341) & (!g337)) + ((g135) & (g123) & (!g186) & (!g227) & (!g341) & (g337)) + ((g135) & (g123) & (!g186) & (!g227) & (g341) & (!g337)) + ((g135) & (g123) & (!g186) & (!g227) & (g341) & (g337)) + ((g135) & (g123) & (!g186) & (g227) & (g341) & (!g337)) + ((g135) & (g123) & (!g186) & (g227) & (g341) & (g337)) + ((g135) & (g123) & (g186) & (!g227) & (!g341) & (!g337)) + ((g135) & (g123) & (g186) & (!g227) & (!g341) & (g337)) + ((g135) & (g123) & (g186) & (!g227) & (g341) & (!g337)) + ((g135) & (g123) & (g186) & (!g227) & (g341) & (g337)) + ((g135) & (g123) & (g186) & (g227) & (g341) & (!g337)) + ((g135) & (g123) & (g186) & (g227) & (g341) & (g337)));
	assign g400 = (((!g356) & (!g369) & (!g393) & (g396) & (!g398) & (g399)) + ((!g356) & (g369) & (!g393) & (g396) & (!g398) & (g399)) + ((g356) & (!g369) & (!g393) & (g396) & (!g398) & (g399)));
	assign g401 = (((!g105) & (!g257) & (!sk[47]) & (g254) & (!g217)) + ((!g105) & (!g257) & (!sk[47]) & (g254) & (g217)) + ((!g105) & (g257) & (!sk[47]) & (g254) & (!g217)) + ((!g105) & (g257) & (!sk[47]) & (g254) & (g217)) + ((g105) & (!g257) & (!sk[47]) & (g254) & (!g217)) + ((g105) & (!g257) & (!sk[47]) & (g254) & (g217)) + ((g105) & (!g257) & (sk[47]) & (g254) & (!g217)) + ((g105) & (g257) & (!sk[47]) & (g254) & (!g217)) + ((g105) & (g257) & (!sk[47]) & (g254) & (g217)));
	assign g402 = (((!g159) & (!g154) & (g122) & (!sk[48]) & (!g257) & (g313)) + ((!g159) & (!g154) & (g122) & (!sk[48]) & (g257) & (!g313)) + ((!g159) & (!g154) & (g122) & (!sk[48]) & (g257) & (g313)) + ((!g159) & (g154) & (!g122) & (!sk[48]) & (!g257) & (!g313)) + ((!g159) & (g154) & (!g122) & (!sk[48]) & (!g257) & (g313)) + ((!g159) & (g154) & (!g122) & (!sk[48]) & (g257) & (!g313)) + ((!g159) & (g154) & (!g122) & (!sk[48]) & (g257) & (g313)) + ((!g159) & (g154) & (g122) & (!sk[48]) & (!g257) & (!g313)) + ((!g159) & (g154) & (g122) & (!sk[48]) & (!g257) & (g313)) + ((!g159) & (g154) & (g122) & (!sk[48]) & (g257) & (!g313)) + ((!g159) & (g154) & (g122) & (!sk[48]) & (g257) & (g313)) + ((g159) & (!g154) & (g122) & (!sk[48]) & (!g257) & (g313)) + ((g159) & (!g154) & (g122) & (!sk[48]) & (g257) & (!g313)) + ((g159) & (!g154) & (g122) & (!sk[48]) & (g257) & (g313)) + ((g159) & (g154) & (!g122) & (!sk[48]) & (!g257) & (!g313)) + ((g159) & (g154) & (!g122) & (!sk[48]) & (!g257) & (g313)) + ((g159) & (g154) & (!g122) & (!sk[48]) & (g257) & (!g313)) + ((g159) & (g154) & (!g122) & (!sk[48]) & (g257) & (g313)) + ((g159) & (g154) & (!g122) & (sk[48]) & (!g257) & (!g313)) + ((g159) & (g154) & (g122) & (!sk[48]) & (!g257) & (!g313)) + ((g159) & (g154) & (g122) & (!sk[48]) & (!g257) & (g313)) + ((g159) & (g154) & (g122) & (!sk[48]) & (g257) & (!g313)) + ((g159) & (g154) & (g122) & (!sk[48]) & (g257) & (g313)));
	assign g403 = (((!i_9_) & (!i_10_) & (!sk[49]) & (i_11_)) + ((!i_9_) & (!i_10_) & (sk[49]) & (i_11_)) + ((!i_9_) & (i_10_) & (!sk[49]) & (!i_11_)) + ((!i_9_) & (i_10_) & (!sk[49]) & (i_11_)) + ((i_9_) & (!i_10_) & (!sk[49]) & (i_11_)) + ((i_9_) & (i_10_) & (!sk[49]) & (!i_11_)) + ((i_9_) & (i_10_) & (!sk[49]) & (i_11_)) + ((i_9_) & (i_10_) & (sk[49]) & (!i_11_)));
	assign g404 = (((!i_15_) & (!g68) & (!g257) & (!g254) & (!g217) & (g403)) + ((!i_15_) & (!g68) & (!g257) & (!g254) & (g217) & (g403)) + ((!i_15_) & (!g68) & (!g257) & (g254) & (g217) & (g403)) + ((!i_15_) & (!g68) & (g257) & (!g254) & (!g217) & (g403)) + ((!i_15_) & (!g68) & (g257) & (!g254) & (g217) & (g403)) + ((!i_15_) & (!g68) & (g257) & (g254) & (!g217) & (g403)) + ((!i_15_) & (!g68) & (g257) & (g254) & (g217) & (g403)));
	assign g405 = (((!g296) & (!g282) & (!sk[51]) & (g401) & (!g402) & (g404)) + ((!g296) & (!g282) & (!sk[51]) & (g401) & (g402) & (!g404)) + ((!g296) & (!g282) & (!sk[51]) & (g401) & (g402) & (g404)) + ((!g296) & (!g282) & (sk[51]) & (!g401) & (!g402) & (!g404)) + ((!g296) & (!g282) & (sk[51]) & (!g401) & (g402) & (!g404)) + ((!g296) & (!g282) & (sk[51]) & (g401) & (!g402) & (!g404)) + ((!g296) & (!g282) & (sk[51]) & (g401) & (g402) & (!g404)) + ((!g296) & (g282) & (!sk[51]) & (!g401) & (!g402) & (!g404)) + ((!g296) & (g282) & (!sk[51]) & (!g401) & (!g402) & (g404)) + ((!g296) & (g282) & (!sk[51]) & (!g401) & (g402) & (!g404)) + ((!g296) & (g282) & (!sk[51]) & (!g401) & (g402) & (g404)) + ((!g296) & (g282) & (!sk[51]) & (g401) & (!g402) & (!g404)) + ((!g296) & (g282) & (!sk[51]) & (g401) & (!g402) & (g404)) + ((!g296) & (g282) & (!sk[51]) & (g401) & (g402) & (!g404)) + ((!g296) & (g282) & (!sk[51]) & (g401) & (g402) & (g404)) + ((!g296) & (g282) & (sk[51]) & (!g401) & (g402) & (!g404)) + ((!g296) & (g282) & (sk[51]) & (g401) & (g402) & (!g404)) + ((g296) & (!g282) & (!sk[51]) & (g401) & (!g402) & (g404)) + ((g296) & (!g282) & (!sk[51]) & (g401) & (g402) & (!g404)) + ((g296) & (!g282) & (!sk[51]) & (g401) & (g402) & (g404)) + ((g296) & (!g282) & (sk[51]) & (g401) & (!g402) & (!g404)) + ((g296) & (!g282) & (sk[51]) & (g401) & (g402) & (!g404)) + ((g296) & (g282) & (!sk[51]) & (!g401) & (!g402) & (!g404)) + ((g296) & (g282) & (!sk[51]) & (!g401) & (!g402) & (g404)) + ((g296) & (g282) & (!sk[51]) & (!g401) & (g402) & (!g404)) + ((g296) & (g282) & (!sk[51]) & (!g401) & (g402) & (g404)) + ((g296) & (g282) & (!sk[51]) & (g401) & (!g402) & (!g404)) + ((g296) & (g282) & (!sk[51]) & (g401) & (!g402) & (g404)) + ((g296) & (g282) & (!sk[51]) & (g401) & (g402) & (!g404)) + ((g296) & (g282) & (!sk[51]) & (g401) & (g402) & (g404)) + ((g296) & (g282) & (sk[51]) & (g401) & (g402) & (!g404)));
	assign g406 = (((!g185) & (!sk[52]) & (!g197) & (g179) & (!g187) & (g282)) + ((!g185) & (!sk[52]) & (!g197) & (g179) & (g187) & (!g282)) + ((!g185) & (!sk[52]) & (!g197) & (g179) & (g187) & (g282)) + ((!g185) & (!sk[52]) & (g197) & (!g179) & (!g187) & (!g282)) + ((!g185) & (!sk[52]) & (g197) & (!g179) & (!g187) & (g282)) + ((!g185) & (!sk[52]) & (g197) & (!g179) & (g187) & (!g282)) + ((!g185) & (!sk[52]) & (g197) & (!g179) & (g187) & (g282)) + ((!g185) & (!sk[52]) & (g197) & (g179) & (!g187) & (!g282)) + ((!g185) & (!sk[52]) & (g197) & (g179) & (!g187) & (g282)) + ((!g185) & (!sk[52]) & (g197) & (g179) & (g187) & (!g282)) + ((!g185) & (!sk[52]) & (g197) & (g179) & (g187) & (g282)) + ((!g185) & (sk[52]) & (!g197) & (!g179) & (!g187) & (!g282)) + ((g185) & (!sk[52]) & (!g197) & (g179) & (!g187) & (g282)) + ((g185) & (!sk[52]) & (!g197) & (g179) & (g187) & (!g282)) + ((g185) & (!sk[52]) & (!g197) & (g179) & (g187) & (g282)) + ((g185) & (!sk[52]) & (g197) & (!g179) & (!g187) & (!g282)) + ((g185) & (!sk[52]) & (g197) & (!g179) & (!g187) & (g282)) + ((g185) & (!sk[52]) & (g197) & (!g179) & (g187) & (!g282)) + ((g185) & (!sk[52]) & (g197) & (!g179) & (g187) & (g282)) + ((g185) & (!sk[52]) & (g197) & (g179) & (!g187) & (!g282)) + ((g185) & (!sk[52]) & (g197) & (g179) & (!g187) & (g282)) + ((g185) & (!sk[52]) & (g197) & (g179) & (g187) & (!g282)) + ((g185) & (!sk[52]) & (g197) & (g179) & (g187) & (g282)));
	assign g407 = (((!i_8_) & (!i_6_) & (!sk[53]) & (i_7_) & (!g72) & (g120)) + ((!i_8_) & (!i_6_) & (!sk[53]) & (i_7_) & (g72) & (!g120)) + ((!i_8_) & (!i_6_) & (!sk[53]) & (i_7_) & (g72) & (g120)) + ((!i_8_) & (!i_6_) & (sk[53]) & (!i_7_) & (!g72) & (g120)) + ((!i_8_) & (!i_6_) & (sk[53]) & (!i_7_) & (g72) & (g120)) + ((!i_8_) & (!i_6_) & (sk[53]) & (i_7_) & (!g72) & (g120)) + ((!i_8_) & (!i_6_) & (sk[53]) & (i_7_) & (g72) & (!g120)) + ((!i_8_) & (!i_6_) & (sk[53]) & (i_7_) & (g72) & (g120)) + ((!i_8_) & (i_6_) & (!sk[53]) & (!i_7_) & (!g72) & (!g120)) + ((!i_8_) & (i_6_) & (!sk[53]) & (!i_7_) & (!g72) & (g120)) + ((!i_8_) & (i_6_) & (!sk[53]) & (!i_7_) & (g72) & (!g120)) + ((!i_8_) & (i_6_) & (!sk[53]) & (!i_7_) & (g72) & (g120)) + ((!i_8_) & (i_6_) & (!sk[53]) & (i_7_) & (!g72) & (!g120)) + ((!i_8_) & (i_6_) & (!sk[53]) & (i_7_) & (!g72) & (g120)) + ((!i_8_) & (i_6_) & (!sk[53]) & (i_7_) & (g72) & (!g120)) + ((!i_8_) & (i_6_) & (!sk[53]) & (i_7_) & (g72) & (g120)) + ((!i_8_) & (i_6_) & (sk[53]) & (i_7_) & (g72) & (!g120)) + ((!i_8_) & (i_6_) & (sk[53]) & (i_7_) & (g72) & (g120)) + ((i_8_) & (!i_6_) & (!sk[53]) & (i_7_) & (!g72) & (g120)) + ((i_8_) & (!i_6_) & (!sk[53]) & (i_7_) & (g72) & (!g120)) + ((i_8_) & (!i_6_) & (!sk[53]) & (i_7_) & (g72) & (g120)) + ((i_8_) & (!i_6_) & (sk[53]) & (i_7_) & (g72) & (!g120)) + ((i_8_) & (!i_6_) & (sk[53]) & (i_7_) & (g72) & (g120)) + ((i_8_) & (i_6_) & (!sk[53]) & (!i_7_) & (!g72) & (!g120)) + ((i_8_) & (i_6_) & (!sk[53]) & (!i_7_) & (!g72) & (g120)) + ((i_8_) & (i_6_) & (!sk[53]) & (!i_7_) & (g72) & (!g120)) + ((i_8_) & (i_6_) & (!sk[53]) & (!i_7_) & (g72) & (g120)) + ((i_8_) & (i_6_) & (!sk[53]) & (i_7_) & (!g72) & (!g120)) + ((i_8_) & (i_6_) & (!sk[53]) & (i_7_) & (!g72) & (g120)) + ((i_8_) & (i_6_) & (!sk[53]) & (i_7_) & (g72) & (!g120)) + ((i_8_) & (i_6_) & (!sk[53]) & (i_7_) & (g72) & (g120)) + ((i_8_) & (i_6_) & (sk[53]) & (!i_7_) & (!g72) & (g120)) + ((i_8_) & (i_6_) & (sk[53]) & (!i_7_) & (g72) & (g120)));
	assign g408 = (((!sk[54]) & (g1) & (!g118)) + ((!sk[54]) & (g1) & (g118)) + ((sk[54]) & (!g1) & (!g118)) + ((sk[54]) & (!g1) & (g118)) + ((sk[54]) & (g1) & (!g118)));
	assign g409 = (((!g272) & (!sk[55]) & (!g334) & (g408)) + ((!g272) & (!sk[55]) & (g334) & (!g408)) + ((!g272) & (!sk[55]) & (g334) & (g408)) + ((!g272) & (sk[55]) & (!g334) & (!g408)) + ((g272) & (!sk[55]) & (!g334) & (g408)) + ((g272) & (!sk[55]) & (g334) & (!g408)) + ((g272) & (!sk[55]) & (g334) & (g408)) + ((g272) & (sk[55]) & (!g334) & (!g408)) + ((g272) & (sk[55]) & (g334) & (!g408)));
	assign g410 = (((!g168) & (!g342) & (!sk[56]) & (g406) & (!g407) & (g409)) + ((!g168) & (!g342) & (!sk[56]) & (g406) & (g407) & (!g409)) + ((!g168) & (!g342) & (!sk[56]) & (g406) & (g407) & (g409)) + ((!g168) & (!g342) & (sk[56]) & (!g406) & (!g407) & (!g409)) + ((!g168) & (!g342) & (sk[56]) & (!g406) & (g407) & (!g409)) + ((!g168) & (!g342) & (sk[56]) & (g406) & (!g407) & (!g409)) + ((!g168) & (!g342) & (sk[56]) & (g406) & (g407) & (!g409)) + ((!g168) & (g342) & (!sk[56]) & (!g406) & (!g407) & (!g409)) + ((!g168) & (g342) & (!sk[56]) & (!g406) & (!g407) & (g409)) + ((!g168) & (g342) & (!sk[56]) & (!g406) & (g407) & (!g409)) + ((!g168) & (g342) & (!sk[56]) & (!g406) & (g407) & (g409)) + ((!g168) & (g342) & (!sk[56]) & (g406) & (!g407) & (!g409)) + ((!g168) & (g342) & (!sk[56]) & (g406) & (!g407) & (g409)) + ((!g168) & (g342) & (!sk[56]) & (g406) & (g407) & (!g409)) + ((!g168) & (g342) & (!sk[56]) & (g406) & (g407) & (g409)) + ((!g168) & (g342) & (sk[56]) & (!g406) & (!g407) & (!g409)) + ((!g168) & (g342) & (sk[56]) & (g406) & (!g407) & (!g409)) + ((g168) & (!g342) & (!sk[56]) & (g406) & (!g407) & (g409)) + ((g168) & (!g342) & (!sk[56]) & (g406) & (g407) & (!g409)) + ((g168) & (!g342) & (!sk[56]) & (g406) & (g407) & (g409)) + ((g168) & (!g342) & (sk[56]) & (g406) & (!g407) & (!g409)) + ((g168) & (!g342) & (sk[56]) & (g406) & (g407) & (!g409)) + ((g168) & (g342) & (!sk[56]) & (!g406) & (!g407) & (!g409)) + ((g168) & (g342) & (!sk[56]) & (!g406) & (!g407) & (g409)) + ((g168) & (g342) & (!sk[56]) & (!g406) & (g407) & (!g409)) + ((g168) & (g342) & (!sk[56]) & (!g406) & (g407) & (g409)) + ((g168) & (g342) & (!sk[56]) & (g406) & (!g407) & (!g409)) + ((g168) & (g342) & (!sk[56]) & (g406) & (!g407) & (g409)) + ((g168) & (g342) & (!sk[56]) & (g406) & (g407) & (!g409)) + ((g168) & (g342) & (!sk[56]) & (g406) & (g407) & (g409)) + ((g168) & (g342) & (sk[56]) & (g406) & (!g407) & (!g409)));
	assign g411 = (((!g388) & (!g391) & (!sk[57]) & (g400) & (!g405) & (g410)) + ((!g388) & (!g391) & (!sk[57]) & (g400) & (g405) & (!g410)) + ((!g388) & (!g391) & (!sk[57]) & (g400) & (g405) & (g410)) + ((!g388) & (g391) & (!sk[57]) & (!g400) & (!g405) & (!g410)) + ((!g388) & (g391) & (!sk[57]) & (!g400) & (!g405) & (g410)) + ((!g388) & (g391) & (!sk[57]) & (!g400) & (g405) & (!g410)) + ((!g388) & (g391) & (!sk[57]) & (!g400) & (g405) & (g410)) + ((!g388) & (g391) & (!sk[57]) & (g400) & (!g405) & (!g410)) + ((!g388) & (g391) & (!sk[57]) & (g400) & (!g405) & (g410)) + ((!g388) & (g391) & (!sk[57]) & (g400) & (g405) & (!g410)) + ((!g388) & (g391) & (!sk[57]) & (g400) & (g405) & (g410)) + ((!g388) & (g391) & (sk[57]) & (g400) & (g405) & (g410)) + ((g388) & (!g391) & (!sk[57]) & (g400) & (!g405) & (g410)) + ((g388) & (!g391) & (!sk[57]) & (g400) & (g405) & (!g410)) + ((g388) & (!g391) & (!sk[57]) & (g400) & (g405) & (g410)) + ((g388) & (g391) & (!sk[57]) & (!g400) & (!g405) & (!g410)) + ((g388) & (g391) & (!sk[57]) & (!g400) & (!g405) & (g410)) + ((g388) & (g391) & (!sk[57]) & (!g400) & (g405) & (!g410)) + ((g388) & (g391) & (!sk[57]) & (!g400) & (g405) & (g410)) + ((g388) & (g391) & (!sk[57]) & (g400) & (!g405) & (!g410)) + ((g388) & (g391) & (!sk[57]) & (g400) & (!g405) & (g410)) + ((g388) & (g391) & (!sk[57]) & (g400) & (g405) & (!g410)) + ((g388) & (g391) & (!sk[57]) & (g400) & (g405) & (g410)));
	assign g412 = (((!g346) & (!sk[58]) & (!g354) & (g361) & (!g387) & (g411)) + ((!g346) & (!sk[58]) & (!g354) & (g361) & (g387) & (!g411)) + ((!g346) & (!sk[58]) & (!g354) & (g361) & (g387) & (g411)) + ((!g346) & (!sk[58]) & (g354) & (!g361) & (!g387) & (!g411)) + ((!g346) & (!sk[58]) & (g354) & (!g361) & (!g387) & (g411)) + ((!g346) & (!sk[58]) & (g354) & (!g361) & (g387) & (!g411)) + ((!g346) & (!sk[58]) & (g354) & (!g361) & (g387) & (g411)) + ((!g346) & (!sk[58]) & (g354) & (g361) & (!g387) & (!g411)) + ((!g346) & (!sk[58]) & (g354) & (g361) & (!g387) & (g411)) + ((!g346) & (!sk[58]) & (g354) & (g361) & (g387) & (!g411)) + ((!g346) & (!sk[58]) & (g354) & (g361) & (g387) & (g411)) + ((g346) & (!sk[58]) & (!g354) & (g361) & (!g387) & (g411)) + ((g346) & (!sk[58]) & (!g354) & (g361) & (g387) & (!g411)) + ((g346) & (!sk[58]) & (!g354) & (g361) & (g387) & (g411)) + ((g346) & (!sk[58]) & (g354) & (!g361) & (!g387) & (!g411)) + ((g346) & (!sk[58]) & (g354) & (!g361) & (!g387) & (g411)) + ((g346) & (!sk[58]) & (g354) & (!g361) & (g387) & (!g411)) + ((g346) & (!sk[58]) & (g354) & (!g361) & (g387) & (g411)) + ((g346) & (!sk[58]) & (g354) & (g361) & (!g387) & (!g411)) + ((g346) & (!sk[58]) & (g354) & (g361) & (!g387) & (g411)) + ((g346) & (!sk[58]) & (g354) & (g361) & (g387) & (!g411)) + ((g346) & (!sk[58]) & (g354) & (g361) & (g387) & (g411)) + ((g346) & (sk[58]) & (!g354) & (g361) & (g387) & (g411)));
	assign g413 = (((!g102) & (!g257) & (!sk[59]) & (g313)) + ((!g102) & (!g257) & (sk[59]) & (!g313)) + ((!g102) & (g257) & (!sk[59]) & (!g313)) + ((!g102) & (g257) & (!sk[59]) & (g313)) + ((g102) & (!g257) & (!sk[59]) & (g313)) + ((g102) & (g257) & (!sk[59]) & (!g313)) + ((g102) & (g257) & (!sk[59]) & (g313)));
	assign g414 = (((!g105) & (!sk[60]) & (!g119) & (g413)) + ((!g105) & (!sk[60]) & (g119) & (!g413)) + ((!g105) & (!sk[60]) & (g119) & (g413)) + ((g105) & (!sk[60]) & (!g119) & (g413)) + ((g105) & (!sk[60]) & (g119) & (!g413)) + ((g105) & (!sk[60]) & (g119) & (g413)) + ((g105) & (sk[60]) & (!g119) & (g413)));
	assign g415 = (((!sk[61]) & (!g78) & (!g131) & (g333)) + ((!sk[61]) & (!g78) & (g131) & (!g333)) + ((!sk[61]) & (!g78) & (g131) & (g333)) + ((!sk[61]) & (g78) & (!g131) & (g333)) + ((!sk[61]) & (g78) & (g131) & (!g333)) + ((!sk[61]) & (g78) & (g131) & (g333)) + ((sk[61]) & (!g78) & (!g131) & (!g333)) + ((sk[61]) & (!g78) & (!g131) & (g333)) + ((sk[61]) & (g78) & (!g131) & (g333)));
	assign g416 = (((!i_9_) & (!i_10_) & (i_11_) & (!i_15_) & (!sk[62]) & (g176)) + ((!i_9_) & (!i_10_) & (i_11_) & (i_15_) & (!sk[62]) & (!g176)) + ((!i_9_) & (!i_10_) & (i_11_) & (i_15_) & (!sk[62]) & (g176)) + ((!i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (!sk[62]) & (!g176)) + ((!i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (!sk[62]) & (g176)) + ((!i_9_) & (i_10_) & (!i_11_) & (i_15_) & (!sk[62]) & (!g176)) + ((!i_9_) & (i_10_) & (!i_11_) & (i_15_) & (!sk[62]) & (g176)) + ((!i_9_) & (i_10_) & (i_11_) & (!i_15_) & (!sk[62]) & (!g176)) + ((!i_9_) & (i_10_) & (i_11_) & (!i_15_) & (!sk[62]) & (g176)) + ((!i_9_) & (i_10_) & (i_11_) & (i_15_) & (!sk[62]) & (!g176)) + ((!i_9_) & (i_10_) & (i_11_) & (i_15_) & (!sk[62]) & (g176)) + ((i_9_) & (!i_10_) & (i_11_) & (!i_15_) & (!sk[62]) & (g176)) + ((i_9_) & (!i_10_) & (i_11_) & (i_15_) & (!sk[62]) & (!g176)) + ((i_9_) & (!i_10_) & (i_11_) & (i_15_) & (!sk[62]) & (g176)) + ((i_9_) & (!i_10_) & (i_11_) & (i_15_) & (sk[62]) & (!g176)) + ((i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (!sk[62]) & (!g176)) + ((i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (!sk[62]) & (g176)) + ((i_9_) & (i_10_) & (!i_11_) & (i_15_) & (!sk[62]) & (!g176)) + ((i_9_) & (i_10_) & (!i_11_) & (i_15_) & (!sk[62]) & (g176)) + ((i_9_) & (i_10_) & (!i_11_) & (i_15_) & (sk[62]) & (!g176)) + ((i_9_) & (i_10_) & (i_11_) & (!i_15_) & (!sk[62]) & (!g176)) + ((i_9_) & (i_10_) & (i_11_) & (!i_15_) & (!sk[62]) & (g176)) + ((i_9_) & (i_10_) & (i_11_) & (i_15_) & (!sk[62]) & (!g176)) + ((i_9_) & (i_10_) & (i_11_) & (i_15_) & (!sk[62]) & (g176)));
	assign g417 = (((!sk[63]) & (!i_6_) & (!g120) & (g154) & (!g197) & (g416)) + ((!sk[63]) & (!i_6_) & (!g120) & (g154) & (g197) & (!g416)) + ((!sk[63]) & (!i_6_) & (!g120) & (g154) & (g197) & (g416)) + ((!sk[63]) & (!i_6_) & (g120) & (!g154) & (!g197) & (!g416)) + ((!sk[63]) & (!i_6_) & (g120) & (!g154) & (!g197) & (g416)) + ((!sk[63]) & (!i_6_) & (g120) & (!g154) & (g197) & (!g416)) + ((!sk[63]) & (!i_6_) & (g120) & (!g154) & (g197) & (g416)) + ((!sk[63]) & (!i_6_) & (g120) & (g154) & (!g197) & (!g416)) + ((!sk[63]) & (!i_6_) & (g120) & (g154) & (!g197) & (g416)) + ((!sk[63]) & (!i_6_) & (g120) & (g154) & (g197) & (!g416)) + ((!sk[63]) & (!i_6_) & (g120) & (g154) & (g197) & (g416)) + ((!sk[63]) & (i_6_) & (!g120) & (g154) & (!g197) & (g416)) + ((!sk[63]) & (i_6_) & (!g120) & (g154) & (g197) & (!g416)) + ((!sk[63]) & (i_6_) & (!g120) & (g154) & (g197) & (g416)) + ((!sk[63]) & (i_6_) & (g120) & (!g154) & (!g197) & (!g416)) + ((!sk[63]) & (i_6_) & (g120) & (!g154) & (!g197) & (g416)) + ((!sk[63]) & (i_6_) & (g120) & (!g154) & (g197) & (!g416)) + ((!sk[63]) & (i_6_) & (g120) & (!g154) & (g197) & (g416)) + ((!sk[63]) & (i_6_) & (g120) & (g154) & (!g197) & (!g416)) + ((!sk[63]) & (i_6_) & (g120) & (g154) & (!g197) & (g416)) + ((!sk[63]) & (i_6_) & (g120) & (g154) & (g197) & (!g416)) + ((!sk[63]) & (i_6_) & (g120) & (g154) & (g197) & (g416)) + ((sk[63]) & (!i_6_) & (!g120) & (!g154) & (g197) & (!g416)) + ((sk[63]) & (!i_6_) & (!g120) & (!g154) & (g197) & (g416)) + ((sk[63]) & (!i_6_) & (g120) & (!g154) & (!g197) & (g416)) + ((sk[63]) & (!i_6_) & (g120) & (!g154) & (g197) & (!g416)) + ((sk[63]) & (!i_6_) & (g120) & (!g154) & (g197) & (g416)) + ((sk[63]) & (!i_6_) & (g120) & (g154) & (!g197) & (g416)) + ((sk[63]) & (!i_6_) & (g120) & (g154) & (g197) & (g416)) + ((sk[63]) & (i_6_) & (!g120) & (!g154) & (g197) & (!g416)) + ((sk[63]) & (i_6_) & (!g120) & (!g154) & (g197) & (g416)) + ((sk[63]) & (i_6_) & (g120) & (!g154) & (g197) & (!g416)) + ((sk[63]) & (i_6_) & (g120) & (!g154) & (g197) & (g416)));
	assign g418 = (((!g355) & (!g35) & (!sk[64]) & (g107) & (!g159) & (g313)) + ((!g355) & (!g35) & (!sk[64]) & (g107) & (g159) & (!g313)) + ((!g355) & (!g35) & (!sk[64]) & (g107) & (g159) & (g313)) + ((!g355) & (g35) & (!sk[64]) & (!g107) & (!g159) & (!g313)) + ((!g355) & (g35) & (!sk[64]) & (!g107) & (!g159) & (g313)) + ((!g355) & (g35) & (!sk[64]) & (!g107) & (g159) & (!g313)) + ((!g355) & (g35) & (!sk[64]) & (!g107) & (g159) & (g313)) + ((!g355) & (g35) & (!sk[64]) & (g107) & (!g159) & (!g313)) + ((!g355) & (g35) & (!sk[64]) & (g107) & (!g159) & (g313)) + ((!g355) & (g35) & (!sk[64]) & (g107) & (g159) & (!g313)) + ((!g355) & (g35) & (!sk[64]) & (g107) & (g159) & (g313)) + ((g355) & (!g35) & (!sk[64]) & (g107) & (!g159) & (g313)) + ((g355) & (!g35) & (!sk[64]) & (g107) & (g159) & (!g313)) + ((g355) & (!g35) & (!sk[64]) & (g107) & (g159) & (g313)) + ((g355) & (!g35) & (sk[64]) & (!g107) & (!g159) & (!g313)) + ((g355) & (!g35) & (sk[64]) & (!g107) & (!g159) & (g313)) + ((g355) & (!g35) & (sk[64]) & (!g107) & (g159) & (g313)) + ((g355) & (g35) & (!sk[64]) & (!g107) & (!g159) & (!g313)) + ((g355) & (g35) & (!sk[64]) & (!g107) & (!g159) & (g313)) + ((g355) & (g35) & (!sk[64]) & (!g107) & (g159) & (!g313)) + ((g355) & (g35) & (!sk[64]) & (!g107) & (g159) & (g313)) + ((g355) & (g35) & (!sk[64]) & (g107) & (!g159) & (!g313)) + ((g355) & (g35) & (!sk[64]) & (g107) & (!g159) & (g313)) + ((g355) & (g35) & (!sk[64]) & (g107) & (g159) & (!g313)) + ((g355) & (g35) & (!sk[64]) & (g107) & (g159) & (g313)) + ((g355) & (g35) & (sk[64]) & (!g107) & (!g159) & (!g313)) + ((g355) & (g35) & (sk[64]) & (!g107) & (!g159) & (g313)) + ((g355) & (g35) & (sk[64]) & (!g107) & (g159) & (g313)) + ((g355) & (g35) & (sk[64]) & (g107) & (!g159) & (g313)) + ((g355) & (g35) & (sk[64]) & (g107) & (g159) & (g313)));
	assign g419 = (((!g20) & (!sk[65]) & (!g355) & (g135) & (!g165) & (g174)) + ((!g20) & (!sk[65]) & (!g355) & (g135) & (g165) & (!g174)) + ((!g20) & (!sk[65]) & (!g355) & (g135) & (g165) & (g174)) + ((!g20) & (!sk[65]) & (g355) & (!g135) & (!g165) & (!g174)) + ((!g20) & (!sk[65]) & (g355) & (!g135) & (!g165) & (g174)) + ((!g20) & (!sk[65]) & (g355) & (!g135) & (g165) & (!g174)) + ((!g20) & (!sk[65]) & (g355) & (!g135) & (g165) & (g174)) + ((!g20) & (!sk[65]) & (g355) & (g135) & (!g165) & (!g174)) + ((!g20) & (!sk[65]) & (g355) & (g135) & (!g165) & (g174)) + ((!g20) & (!sk[65]) & (g355) & (g135) & (g165) & (!g174)) + ((!g20) & (!sk[65]) & (g355) & (g135) & (g165) & (g174)) + ((g20) & (!sk[65]) & (!g355) & (g135) & (!g165) & (g174)) + ((g20) & (!sk[65]) & (!g355) & (g135) & (g165) & (!g174)) + ((g20) & (!sk[65]) & (!g355) & (g135) & (g165) & (g174)) + ((g20) & (!sk[65]) & (g355) & (!g135) & (!g165) & (!g174)) + ((g20) & (!sk[65]) & (g355) & (!g135) & (!g165) & (g174)) + ((g20) & (!sk[65]) & (g355) & (!g135) & (g165) & (!g174)) + ((g20) & (!sk[65]) & (g355) & (!g135) & (g165) & (g174)) + ((g20) & (!sk[65]) & (g355) & (g135) & (!g165) & (!g174)) + ((g20) & (!sk[65]) & (g355) & (g135) & (!g165) & (g174)) + ((g20) & (!sk[65]) & (g355) & (g135) & (g165) & (!g174)) + ((g20) & (!sk[65]) & (g355) & (g135) & (g165) & (g174)) + ((g20) & (sk[65]) & (!g355) & (!g135) & (!g165) & (!g174)) + ((g20) & (sk[65]) & (!g355) & (!g135) & (g165) & (!g174)) + ((g20) & (sk[65]) & (g355) & (!g135) & (!g165) & (!g174)) + ((g20) & (sk[65]) & (g355) & (!g135) & (g165) & (!g174)) + ((g20) & (sk[65]) & (g355) & (!g135) & (g165) & (g174)) + ((g20) & (sk[65]) & (g355) & (g135) & (g165) & (!g174)) + ((g20) & (sk[65]) & (g355) & (g135) & (g165) & (g174)));
	assign g420 = (((!g194) & (!g414) & (!g415) & (!g417) & (!g418) & (!g419)) + ((!g194) & (g414) & (!g415) & (!g417) & (!g418) & (!g419)) + ((g194) & (g414) & (!g415) & (!g417) & (!g418) & (!g419)));
	assign g421 = (((!sk[67]) & (g1) & (!g120)) + ((!sk[67]) & (g1) & (g120)) + ((sk[67]) & (g1) & (g120)));
	assign g422 = (((!g159) & (!g313) & (!sk[68]) & (g421)) + ((!g159) & (!g313) & (sk[68]) & (!g421)) + ((!g159) & (!g313) & (sk[68]) & (g421)) + ((!g159) & (g313) & (!sk[68]) & (!g421)) + ((!g159) & (g313) & (!sk[68]) & (g421)) + ((!g159) & (g313) & (sk[68]) & (!g421)) + ((!g159) & (g313) & (sk[68]) & (g421)) + ((g159) & (!g313) & (!sk[68]) & (g421)) + ((g159) & (!g313) & (sk[68]) & (g421)) + ((g159) & (g313) & (!sk[68]) & (!g421)) + ((g159) & (g313) & (!sk[68]) & (g421)) + ((g159) & (g313) & (sk[68]) & (!g421)) + ((g159) & (g313) & (sk[68]) & (g421)));
	assign g423 = (((!sk[69]) & (!i_15_) & (!g34) & (g68) & (!g422)) + ((!sk[69]) & (!i_15_) & (!g34) & (g68) & (g422)) + ((!sk[69]) & (!i_15_) & (g34) & (g68) & (!g422)) + ((!sk[69]) & (!i_15_) & (g34) & (g68) & (g422)) + ((!sk[69]) & (i_15_) & (!g34) & (g68) & (!g422)) + ((!sk[69]) & (i_15_) & (!g34) & (g68) & (g422)) + ((!sk[69]) & (i_15_) & (g34) & (g68) & (!g422)) + ((!sk[69]) & (i_15_) & (g34) & (g68) & (g422)) + ((sk[69]) & (i_15_) & (g34) & (!g68) & (g422)));
	assign g424 = (((!g25) & (!sk[70]) & (!g130) & (g397)) + ((!g25) & (!sk[70]) & (g130) & (!g397)) + ((!g25) & (!sk[70]) & (g130) & (g397)) + ((!g25) & (sk[70]) & (!g130) & (!g397)) + ((!g25) & (sk[70]) & (!g130) & (g397)) + ((g25) & (!sk[70]) & (!g130) & (g397)) + ((g25) & (!sk[70]) & (g130) & (!g397)) + ((g25) & (!sk[70]) & (g130) & (g397)) + ((g25) & (sk[70]) & (!g130) & (g397)));
	assign g425 = (((!g257) & (!g254) & (!sk[71]) & (g217)) + ((!g257) & (g254) & (!sk[71]) & (!g217)) + ((!g257) & (g254) & (!sk[71]) & (g217)) + ((!g257) & (g254) & (sk[71]) & (!g217)) + ((g257) & (!g254) & (!sk[71]) & (g217)) + ((g257) & (g254) & (!sk[71]) & (!g217)) + ((g257) & (g254) & (!sk[71]) & (g217)));
	assign g426 = (((!g92) & (!g105) & (!sk[72]) & (g275) & (!g425)) + ((!g92) & (!g105) & (!sk[72]) & (g275) & (g425)) + ((!g92) & (!g105) & (sk[72]) & (!g275) & (!g425)) + ((!g92) & (!g105) & (sk[72]) & (!g275) & (g425)) + ((!g92) & (g105) & (!sk[72]) & (g275) & (!g425)) + ((!g92) & (g105) & (!sk[72]) & (g275) & (g425)) + ((!g92) & (g105) & (sk[72]) & (!g275) & (!g425)) + ((!g92) & (g105) & (sk[72]) & (!g275) & (g425)) + ((!g92) & (g105) & (sk[72]) & (g275) & (g425)) + ((g92) & (!g105) & (!sk[72]) & (g275) & (!g425)) + ((g92) & (!g105) & (!sk[72]) & (g275) & (g425)) + ((g92) & (g105) & (!sk[72]) & (g275) & (!g425)) + ((g92) & (g105) & (!sk[72]) & (g275) & (g425)) + ((g92) & (g105) & (sk[72]) & (!g275) & (!g425)) + ((g92) & (g105) & (sk[72]) & (!g275) & (g425)) + ((g92) & (g105) & (sk[72]) & (g275) & (g425)));
	assign g427 = (((!sk[73]) & (!g161) & (!g183) & (g423) & (!g424) & (g426)) + ((!sk[73]) & (!g161) & (!g183) & (g423) & (g424) & (!g426)) + ((!sk[73]) & (!g161) & (!g183) & (g423) & (g424) & (g426)) + ((!sk[73]) & (!g161) & (g183) & (!g423) & (!g424) & (!g426)) + ((!sk[73]) & (!g161) & (g183) & (!g423) & (!g424) & (g426)) + ((!sk[73]) & (!g161) & (g183) & (!g423) & (g424) & (!g426)) + ((!sk[73]) & (!g161) & (g183) & (!g423) & (g424) & (g426)) + ((!sk[73]) & (!g161) & (g183) & (g423) & (!g424) & (!g426)) + ((!sk[73]) & (!g161) & (g183) & (g423) & (!g424) & (g426)) + ((!sk[73]) & (!g161) & (g183) & (g423) & (g424) & (!g426)) + ((!sk[73]) & (!g161) & (g183) & (g423) & (g424) & (g426)) + ((!sk[73]) & (g161) & (!g183) & (g423) & (!g424) & (g426)) + ((!sk[73]) & (g161) & (!g183) & (g423) & (g424) & (!g426)) + ((!sk[73]) & (g161) & (!g183) & (g423) & (g424) & (g426)) + ((!sk[73]) & (g161) & (g183) & (!g423) & (!g424) & (!g426)) + ((!sk[73]) & (g161) & (g183) & (!g423) & (!g424) & (g426)) + ((!sk[73]) & (g161) & (g183) & (!g423) & (g424) & (!g426)) + ((!sk[73]) & (g161) & (g183) & (!g423) & (g424) & (g426)) + ((!sk[73]) & (g161) & (g183) & (g423) & (!g424) & (!g426)) + ((!sk[73]) & (g161) & (g183) & (g423) & (!g424) & (g426)) + ((!sk[73]) & (g161) & (g183) & (g423) & (g424) & (!g426)) + ((!sk[73]) & (g161) & (g183) & (g423) & (g424) & (g426)) + ((sk[73]) & (!g161) & (!g183) & (!g423) & (!g424) & (g426)) + ((sk[73]) & (!g161) & (g183) & (!g423) & (!g424) & (g426)) + ((sk[73]) & (g161) & (!g183) & (!g423) & (!g424) & (g426)));
	assign g428 = (((!i_9_) & (!sk[74]) & (!i_10_) & (i_11_)) + ((!i_9_) & (!sk[74]) & (i_10_) & (!i_11_)) + ((!i_9_) & (!sk[74]) & (i_10_) & (i_11_)) + ((!i_9_) & (sk[74]) & (!i_10_) & (!i_11_)) + ((!i_9_) & (sk[74]) & (!i_10_) & (i_11_)) + ((!i_9_) & (sk[74]) & (i_10_) & (i_11_)) + ((i_9_) & (!sk[74]) & (!i_10_) & (i_11_)) + ((i_9_) & (!sk[74]) & (i_10_) & (!i_11_)) + ((i_9_) & (!sk[74]) & (i_10_) & (i_11_)) + ((i_9_) & (sk[74]) & (!i_10_) & (!i_11_)) + ((i_9_) & (sk[74]) & (!i_10_) & (i_11_)) + ((i_9_) & (sk[74]) & (i_10_) & (!i_11_)) + ((i_9_) & (sk[74]) & (i_10_) & (i_11_)));
	assign g429 = (((!i_9_) & (!i_10_) & (!sk[75]) & (i_11_)) + ((!i_9_) & (i_10_) & (!sk[75]) & (!i_11_)) + ((!i_9_) & (i_10_) & (!sk[75]) & (i_11_)) + ((i_9_) & (!i_10_) & (!sk[75]) & (i_11_)) + ((i_9_) & (!i_10_) & (sk[75]) & (i_11_)) + ((i_9_) & (i_10_) & (!sk[75]) & (!i_11_)) + ((i_9_) & (i_10_) & (!sk[75]) & (i_11_)));
	assign g430 = (((!i_15_) & (!g428) & (!sk[76]) & (g68) & (!g429)) + ((!i_15_) & (!g428) & (!sk[76]) & (g68) & (g429)) + ((!i_15_) & (!g428) & (sk[76]) & (!g68) & (!g429)) + ((!i_15_) & (!g428) & (sk[76]) & (!g68) & (g429)) + ((!i_15_) & (g428) & (!sk[76]) & (g68) & (!g429)) + ((!i_15_) & (g428) & (!sk[76]) & (g68) & (g429)) + ((!i_15_) & (g428) & (sk[76]) & (!g68) & (g429)) + ((i_15_) & (!g428) & (!sk[76]) & (g68) & (!g429)) + ((i_15_) & (!g428) & (!sk[76]) & (g68) & (g429)) + ((i_15_) & (!g428) & (sk[76]) & (!g68) & (g429)) + ((i_15_) & (g428) & (!sk[76]) & (g68) & (!g429)) + ((i_15_) & (g428) & (!sk[76]) & (g68) & (g429)) + ((i_15_) & (g428) & (sk[76]) & (!g68) & (g429)));
	assign g431 = (((!i_8_) & (!sk[77]) & (!i_6_) & (i_7_) & (!g120)) + ((!i_8_) & (!sk[77]) & (!i_6_) & (i_7_) & (g120)) + ((!i_8_) & (!sk[77]) & (i_6_) & (i_7_) & (!g120)) + ((!i_8_) & (!sk[77]) & (i_6_) & (i_7_) & (g120)) + ((!i_8_) & (sk[77]) & (!i_6_) & (i_7_) & (g120)) + ((i_8_) & (!sk[77]) & (!i_6_) & (i_7_) & (!g120)) + ((i_8_) & (!sk[77]) & (!i_6_) & (i_7_) & (g120)) + ((i_8_) & (!sk[77]) & (i_6_) & (i_7_) & (!g120)) + ((i_8_) & (!sk[77]) & (i_6_) & (i_7_) & (g120)) + ((i_8_) & (sk[77]) & (!i_6_) & (!i_7_) & (g120)));
	assign g432 = (((!g159) & (!sk[78]) & (!g185) & (g272) & (!g431)) + ((!g159) & (!sk[78]) & (!g185) & (g272) & (g431)) + ((!g159) & (!sk[78]) & (g185) & (g272) & (!g431)) + ((!g159) & (!sk[78]) & (g185) & (g272) & (g431)) + ((!g159) & (sk[78]) & (!g185) & (g272) & (!g431)) + ((!g159) & (sk[78]) & (!g185) & (g272) & (g431)) + ((!g159) & (sk[78]) & (g185) & (!g272) & (g431)) + ((!g159) & (sk[78]) & (g185) & (g272) & (!g431)) + ((!g159) & (sk[78]) & (g185) & (g272) & (g431)) + ((g159) & (!sk[78]) & (!g185) & (g272) & (!g431)) + ((g159) & (!sk[78]) & (!g185) & (g272) & (g431)) + ((g159) & (!sk[78]) & (g185) & (g272) & (!g431)) + ((g159) & (!sk[78]) & (g185) & (g272) & (g431)) + ((g159) & (sk[78]) & (g185) & (!g272) & (g431)) + ((g159) & (sk[78]) & (g185) & (g272) & (g431)));
	assign g433 = (((!g425) & (!g402) & (!sk[79]) & (g341) & (!g430) & (g432)) + ((!g425) & (!g402) & (!sk[79]) & (g341) & (g430) & (!g432)) + ((!g425) & (!g402) & (!sk[79]) & (g341) & (g430) & (g432)) + ((!g425) & (!g402) & (sk[79]) & (g341) & (!g430) & (!g432)) + ((!g425) & (g402) & (!sk[79]) & (!g341) & (!g430) & (!g432)) + ((!g425) & (g402) & (!sk[79]) & (!g341) & (!g430) & (g432)) + ((!g425) & (g402) & (!sk[79]) & (!g341) & (g430) & (!g432)) + ((!g425) & (g402) & (!sk[79]) & (!g341) & (g430) & (g432)) + ((!g425) & (g402) & (!sk[79]) & (g341) & (!g430) & (!g432)) + ((!g425) & (g402) & (!sk[79]) & (g341) & (!g430) & (g432)) + ((!g425) & (g402) & (!sk[79]) & (g341) & (g430) & (!g432)) + ((!g425) & (g402) & (!sk[79]) & (g341) & (g430) & (g432)) + ((!g425) & (g402) & (sk[79]) & (!g341) & (!g430) & (!g432)) + ((!g425) & (g402) & (sk[79]) & (g341) & (!g430) & (!g432)) + ((g425) & (!g402) & (!sk[79]) & (g341) & (!g430) & (g432)) + ((g425) & (!g402) & (!sk[79]) & (g341) & (g430) & (!g432)) + ((g425) & (!g402) & (!sk[79]) & (g341) & (g430) & (g432)) + ((g425) & (!g402) & (sk[79]) & (g341) & (!g430) & (!g432)) + ((g425) & (!g402) & (sk[79]) & (g341) & (g430) & (!g432)) + ((g425) & (g402) & (!sk[79]) & (!g341) & (!g430) & (!g432)) + ((g425) & (g402) & (!sk[79]) & (!g341) & (!g430) & (g432)) + ((g425) & (g402) & (!sk[79]) & (!g341) & (g430) & (!g432)) + ((g425) & (g402) & (!sk[79]) & (!g341) & (g430) & (g432)) + ((g425) & (g402) & (!sk[79]) & (g341) & (!g430) & (!g432)) + ((g425) & (g402) & (!sk[79]) & (g341) & (!g430) & (g432)) + ((g425) & (g402) & (!sk[79]) & (g341) & (g430) & (!g432)) + ((g425) & (g402) & (!sk[79]) & (g341) & (g430) & (g432)) + ((g425) & (g402) & (sk[79]) & (!g341) & (!g430) & (!g432)) + ((g425) & (g402) & (sk[79]) & (!g341) & (g430) & (!g432)) + ((g425) & (g402) & (sk[79]) & (g341) & (!g430) & (!g432)) + ((g425) & (g402) & (sk[79]) & (g341) & (g430) & (!g432)));
	assign g434 = (((!i_8_) & (!i_6_) & (i_7_) & (!g72) & (!g120) & (g118)) + ((!i_8_) & (!i_6_) & (i_7_) & (!g72) & (g120) & (g118)) + ((!i_8_) & (!i_6_) & (i_7_) & (g72) & (!g120) & (!g118)) + ((!i_8_) & (!i_6_) & (i_7_) & (g72) & (!g120) & (g118)) + ((!i_8_) & (!i_6_) & (i_7_) & (g72) & (g120) & (!g118)) + ((!i_8_) & (!i_6_) & (i_7_) & (g72) & (g120) & (g118)) + ((!i_8_) & (i_6_) & (i_7_) & (!g72) & (g120) & (!g118)) + ((!i_8_) & (i_6_) & (i_7_) & (!g72) & (g120) & (g118)) + ((!i_8_) & (i_6_) & (i_7_) & (g72) & (g120) & (!g118)) + ((!i_8_) & (i_6_) & (i_7_) & (g72) & (g120) & (g118)) + ((i_8_) & (i_6_) & (i_7_) & (!g72) & (!g120) & (g118)) + ((i_8_) & (i_6_) & (i_7_) & (!g72) & (g120) & (g118)) + ((i_8_) & (i_6_) & (i_7_) & (g72) & (!g120) & (!g118)) + ((i_8_) & (i_6_) & (i_7_) & (g72) & (!g120) & (g118)) + ((i_8_) & (i_6_) & (i_7_) & (g72) & (g120) & (!g118)) + ((i_8_) & (i_6_) & (i_7_) & (g72) & (g120) & (g118)));
	assign g435 = (((!sk[81]) & (!g154) & (!g253) & (g356) & (!g383)) + ((!sk[81]) & (!g154) & (!g253) & (g356) & (g383)) + ((!sk[81]) & (!g154) & (g253) & (g356) & (!g383)) + ((!sk[81]) & (!g154) & (g253) & (g356) & (g383)) + ((!sk[81]) & (g154) & (!g253) & (g356) & (!g383)) + ((!sk[81]) & (g154) & (!g253) & (g356) & (g383)) + ((!sk[81]) & (g154) & (g253) & (g356) & (!g383)) + ((!sk[81]) & (g154) & (g253) & (g356) & (g383)) + ((sk[81]) & (g154) & (g253) & (!g356) & (g383)));
	assign g436 = (((!g164) & (!g213) & (!sk[82]) & (g402)) + ((!g164) & (!g213) & (sk[82]) & (!g402)) + ((!g164) & (g213) & (!sk[82]) & (!g402)) + ((!g164) & (g213) & (!sk[82]) & (g402)) + ((!g164) & (g213) & (sk[82]) & (!g402)) + ((!g164) & (g213) & (sk[82]) & (g402)) + ((g164) & (!g213) & (!sk[82]) & (g402)) + ((g164) & (!g213) & (sk[82]) & (!g402)) + ((g164) & (!g213) & (sk[82]) & (g402)) + ((g164) & (g213) & (!sk[82]) & (!g402)) + ((g164) & (g213) & (!sk[82]) & (g402)) + ((g164) & (g213) & (sk[82]) & (!g402)) + ((g164) & (g213) & (sk[82]) & (g402)));
	assign g437 = (((!g70) & (!g82) & (!g357) & (!g434) & (!g435) & (!g436)) + ((!g70) & (!g82) & (!g357) & (!g434) & (!g435) & (g436)) + ((!g70) & (!g82) & (!g357) & (!g434) & (g435) & (!g436)) + ((!g70) & (!g82) & (!g357) & (!g434) & (g435) & (g436)) + ((!g70) & (!g82) & (!g357) & (g434) & (!g435) & (!g436)) + ((!g70) & (!g82) & (!g357) & (g434) & (!g435) & (g436)) + ((!g70) & (!g82) & (!g357) & (g434) & (g435) & (!g436)) + ((!g70) & (!g82) & (!g357) & (g434) & (g435) & (g436)) + ((!g70) & (!g82) & (g357) & (!g434) & (!g435) & (!g436)) + ((!g70) & (!g82) & (g357) & (!g434) & (!g435) & (g436)) + ((!g70) & (!g82) & (g357) & (!g434) & (g435) & (!g436)) + ((!g70) & (!g82) & (g357) & (!g434) & (g435) & (g436)) + ((!g70) & (g82) & (!g357) & (!g434) & (g435) & (!g436)) + ((!g70) & (g82) & (!g357) & (!g434) & (g435) & (g436)) + ((!g70) & (g82) & (!g357) & (g434) & (g435) & (!g436)) + ((!g70) & (g82) & (!g357) & (g434) & (g435) & (g436)) + ((!g70) & (g82) & (g357) & (!g434) & (g435) & (!g436)) + ((!g70) & (g82) & (g357) & (!g434) & (g435) & (g436)) + ((g70) & (!g82) & (!g357) & (!g434) & (!g435) & (!g436)) + ((g70) & (!g82) & (!g357) & (!g434) & (g435) & (!g436)) + ((g70) & (!g82) & (!g357) & (g434) & (!g435) & (!g436)) + ((g70) & (!g82) & (!g357) & (g434) & (g435) & (!g436)) + ((g70) & (!g82) & (g357) & (!g434) & (!g435) & (!g436)) + ((g70) & (!g82) & (g357) & (!g434) & (g435) & (!g436)) + ((g70) & (g82) & (!g357) & (!g434) & (g435) & (!g436)) + ((g70) & (g82) & (!g357) & (g434) & (g435) & (!g436)) + ((g70) & (g82) & (g357) & (!g434) & (g435) & (!g436)));
	assign g438 = (((!g102) & (!g122) & (!g257) & (sk[84]) & (!g313)) + ((!g102) & (!g122) & (g257) & (!sk[84]) & (!g313)) + ((!g102) & (!g122) & (g257) & (!sk[84]) & (g313)) + ((!g102) & (g122) & (g257) & (!sk[84]) & (!g313)) + ((!g102) & (g122) & (g257) & (!sk[84]) & (g313)) + ((g102) & (!g122) & (g257) & (!sk[84]) & (!g313)) + ((g102) & (!g122) & (g257) & (!sk[84]) & (g313)) + ((g102) & (g122) & (g257) & (!sk[84]) & (!g313)) + ((g102) & (g122) & (g257) & (!sk[84]) & (g313)));
	assign g439 = (((!g73) & (!sk[85]) & (!g159) & (g123) & (!g142)) + ((!g73) & (!sk[85]) & (!g159) & (g123) & (g142)) + ((!g73) & (!sk[85]) & (g159) & (g123) & (!g142)) + ((!g73) & (!sk[85]) & (g159) & (g123) & (g142)) + ((!g73) & (sk[85]) & (g159) & (g123) & (g142)) + ((g73) & (!sk[85]) & (!g159) & (g123) & (!g142)) + ((g73) & (!sk[85]) & (!g159) & (g123) & (g142)) + ((g73) & (!sk[85]) & (g159) & (g123) & (!g142)) + ((g73) & (!sk[85]) & (g159) & (g123) & (g142)));
	assign g440 = (((!g105) & (!sk[86]) & (!g438) & (g439)) + ((!g105) & (!sk[86]) & (g438) & (!g439)) + ((!g105) & (!sk[86]) & (g438) & (g439)) + ((g105) & (!sk[86]) & (!g438) & (g439)) + ((g105) & (!sk[86]) & (g438) & (!g439)) + ((g105) & (!sk[86]) & (g438) & (g439)) + ((g105) & (sk[86]) & (g438) & (g439)));
	assign g441 = (((!sk[87]) & (!g413) & (!g217) & (g286) & (!g340) & (g440)) + ((!sk[87]) & (!g413) & (!g217) & (g286) & (g340) & (!g440)) + ((!sk[87]) & (!g413) & (!g217) & (g286) & (g340) & (g440)) + ((!sk[87]) & (!g413) & (g217) & (!g286) & (!g340) & (!g440)) + ((!sk[87]) & (!g413) & (g217) & (!g286) & (!g340) & (g440)) + ((!sk[87]) & (!g413) & (g217) & (!g286) & (g340) & (!g440)) + ((!sk[87]) & (!g413) & (g217) & (!g286) & (g340) & (g440)) + ((!sk[87]) & (!g413) & (g217) & (g286) & (!g340) & (!g440)) + ((!sk[87]) & (!g413) & (g217) & (g286) & (!g340) & (g440)) + ((!sk[87]) & (!g413) & (g217) & (g286) & (g340) & (!g440)) + ((!sk[87]) & (!g413) & (g217) & (g286) & (g340) & (g440)) + ((!sk[87]) & (g413) & (!g217) & (g286) & (!g340) & (g440)) + ((!sk[87]) & (g413) & (!g217) & (g286) & (g340) & (!g440)) + ((!sk[87]) & (g413) & (!g217) & (g286) & (g340) & (g440)) + ((!sk[87]) & (g413) & (g217) & (!g286) & (!g340) & (!g440)) + ((!sk[87]) & (g413) & (g217) & (!g286) & (!g340) & (g440)) + ((!sk[87]) & (g413) & (g217) & (!g286) & (g340) & (!g440)) + ((!sk[87]) & (g413) & (g217) & (!g286) & (g340) & (g440)) + ((!sk[87]) & (g413) & (g217) & (g286) & (!g340) & (!g440)) + ((!sk[87]) & (g413) & (g217) & (g286) & (!g340) & (g440)) + ((!sk[87]) & (g413) & (g217) & (g286) & (g340) & (!g440)) + ((!sk[87]) & (g413) & (g217) & (g286) & (g340) & (g440)) + ((sk[87]) & (!g413) & (!g217) & (!g286) & (!g340) & (g440)) + ((sk[87]) & (!g413) & (!g217) & (!g286) & (g340) & (!g440)) + ((sk[87]) & (!g413) & (!g217) & (!g286) & (g340) & (g440)) + ((sk[87]) & (!g413) & (g217) & (!g286) & (!g340) & (g440)) + ((sk[87]) & (!g413) & (g217) & (!g286) & (g340) & (!g440)) + ((sk[87]) & (!g413) & (g217) & (!g286) & (g340) & (g440)) + ((sk[87]) & (g413) & (!g217) & (!g286) & (!g340) & (g440)) + ((sk[87]) & (g413) & (!g217) & (!g286) & (g340) & (!g440)) + ((sk[87]) & (g413) & (!g217) & (!g286) & (g340) & (g440)) + ((sk[87]) & (g413) & (!g217) & (g286) & (!g340) & (g440)) + ((sk[87]) & (g413) & (!g217) & (g286) & (g340) & (!g440)) + ((sk[87]) & (g413) & (!g217) & (g286) & (g340) & (g440)) + ((sk[87]) & (g413) & (g217) & (!g286) & (!g340) & (g440)) + ((sk[87]) & (g413) & (g217) & (!g286) & (g340) & (!g440)) + ((sk[87]) & (g413) & (g217) & (!g286) & (g340) & (g440)));
	assign g442 = (((g420) & (g427) & (g433) & (g437) & (g441) & (g1593)));
	assign g443 = (((!sk[89]) & (!g73) & (!g164) & (g402)) + ((!sk[89]) & (!g73) & (g164) & (!g402)) + ((!sk[89]) & (!g73) & (g164) & (g402)) + ((!sk[89]) & (g73) & (!g164) & (g402)) + ((!sk[89]) & (g73) & (g164) & (!g402)) + ((!sk[89]) & (g73) & (g164) & (g402)) + ((sk[89]) & (!g73) & (!g164) & (g402)));
	assign g444 = (((!sk[90]) & (!g142) & (!g105) & (g259)) + ((!sk[90]) & (!g142) & (g105) & (!g259)) + ((!sk[90]) & (!g142) & (g105) & (g259)) + ((!sk[90]) & (g142) & (!g105) & (g259)) + ((!sk[90]) & (g142) & (g105) & (!g259)) + ((!sk[90]) & (g142) & (g105) & (g259)) + ((sk[90]) & (g142) & (g105) & (g259)));
	assign g445 = (((!sk[91]) & (g80) & (!i_11_)) + ((!sk[91]) & (g80) & (i_11_)) + ((sk[91]) & (g80) & (i_11_)));
	assign g446 = (((!g125) & (!sk[92]) & (!g413) & (g439)) + ((!g125) & (!sk[92]) & (g413) & (!g439)) + ((!g125) & (!sk[92]) & (g413) & (g439)) + ((!g125) & (sk[92]) & (g413) & (g439)) + ((g125) & (!sk[92]) & (!g413) & (g439)) + ((g125) & (!sk[92]) & (g413) & (!g439)) + ((g125) & (!sk[92]) & (g413) & (g439)));
	assign g447 = (((g142) & (!sk[93]) & (!g217)) + ((g142) & (!sk[93]) & (g217)) + ((g142) & (sk[93]) & (!g217)));
	assign g448 = (((!i_15_) & (!g428) & (!g445) & (!g176) & (!g446) & (!g447)) + ((!i_15_) & (!g428) & (!g445) & (!g176) & (!g446) & (g447)) + ((!i_15_) & (!g428) & (g445) & (!g176) & (!g446) & (!g447)) + ((!i_15_) & (!g428) & (g445) & (!g176) & (!g446) & (g447)) + ((i_15_) & (!g428) & (g445) & (!g176) & (!g446) & (!g447)) + ((i_15_) & (!g428) & (g445) & (!g176) & (g446) & (!g447)) + ((i_15_) & (g428) & (g445) & (!g176) & (!g446) & (!g447)) + ((i_15_) & (g428) & (g445) & (!g176) & (g446) & (!g447)));
	assign g449 = (((!g78) & (!g177) & (g278) & (!sk[95]) & (!g333)) + ((!g78) & (!g177) & (g278) & (!sk[95]) & (g333)) + ((!g78) & (g177) & (g278) & (!sk[95]) & (!g333)) + ((!g78) & (g177) & (g278) & (!sk[95]) & (g333)) + ((g78) & (!g177) & (!g278) & (sk[95]) & (!g333)) + ((g78) & (!g177) & (g278) & (!sk[95]) & (!g333)) + ((g78) & (!g177) & (g278) & (!sk[95]) & (g333)) + ((g78) & (g177) & (g278) & (!sk[95]) & (!g333)) + ((g78) & (g177) & (g278) & (!sk[95]) & (g333)));
	assign g450 = (((!g24) & (!g35) & (!sk[96]) & (g36) & (!g161) & (g68)) + ((!g24) & (!g35) & (!sk[96]) & (g36) & (g161) & (!g68)) + ((!g24) & (!g35) & (!sk[96]) & (g36) & (g161) & (g68)) + ((!g24) & (!g35) & (sk[96]) & (g36) & (!g161) & (!g68)) + ((!g24) & (!g35) & (sk[96]) & (g36) & (g161) & (!g68)) + ((!g24) & (g35) & (!sk[96]) & (!g36) & (!g161) & (!g68)) + ((!g24) & (g35) & (!sk[96]) & (!g36) & (!g161) & (g68)) + ((!g24) & (g35) & (!sk[96]) & (!g36) & (g161) & (!g68)) + ((!g24) & (g35) & (!sk[96]) & (!g36) & (g161) & (g68)) + ((!g24) & (g35) & (!sk[96]) & (g36) & (!g161) & (!g68)) + ((!g24) & (g35) & (!sk[96]) & (g36) & (!g161) & (g68)) + ((!g24) & (g35) & (!sk[96]) & (g36) & (g161) & (!g68)) + ((!g24) & (g35) & (!sk[96]) & (g36) & (g161) & (g68)) + ((!g24) & (g35) & (sk[96]) & (!g36) & (!g161) & (!g68)) + ((!g24) & (g35) & (sk[96]) & (!g36) & (!g161) & (g68)) + ((!g24) & (g35) & (sk[96]) & (!g36) & (g161) & (!g68)) + ((!g24) & (g35) & (sk[96]) & (!g36) & (g161) & (g68)) + ((!g24) & (g35) & (sk[96]) & (g36) & (!g161) & (!g68)) + ((!g24) & (g35) & (sk[96]) & (g36) & (!g161) & (g68)) + ((!g24) & (g35) & (sk[96]) & (g36) & (g161) & (!g68)) + ((!g24) & (g35) & (sk[96]) & (g36) & (g161) & (g68)) + ((g24) & (!g35) & (!sk[96]) & (g36) & (!g161) & (g68)) + ((g24) & (!g35) & (!sk[96]) & (g36) & (g161) & (!g68)) + ((g24) & (!g35) & (!sk[96]) & (g36) & (g161) & (g68)) + ((g24) & (!g35) & (sk[96]) & (g36) & (!g161) & (!g68)) + ((g24) & (!g35) & (sk[96]) & (g36) & (g161) & (!g68)) + ((g24) & (g35) & (!sk[96]) & (!g36) & (!g161) & (!g68)) + ((g24) & (g35) & (!sk[96]) & (!g36) & (!g161) & (g68)) + ((g24) & (g35) & (!sk[96]) & (!g36) & (g161) & (!g68)) + ((g24) & (g35) & (!sk[96]) & (!g36) & (g161) & (g68)) + ((g24) & (g35) & (!sk[96]) & (g36) & (!g161) & (!g68)) + ((g24) & (g35) & (!sk[96]) & (g36) & (!g161) & (g68)) + ((g24) & (g35) & (!sk[96]) & (g36) & (g161) & (!g68)) + ((g24) & (g35) & (!sk[96]) & (g36) & (g161) & (g68)) + ((g24) & (g35) & (sk[96]) & (!g36) & (g161) & (!g68)) + ((g24) & (g35) & (sk[96]) & (g36) & (!g161) & (!g68)) + ((g24) & (g35) & (sk[96]) & (g36) & (g161) & (!g68)));
	assign g451 = (((!g20) & (!g355) & (!sk[97]) & (g78)) + ((!g20) & (!g355) & (sk[97]) & (g78)) + ((!g20) & (g355) & (!sk[97]) & (!g78)) + ((!g20) & (g355) & (!sk[97]) & (g78)) + ((!g20) & (g355) & (sk[97]) & (g78)) + ((g20) & (!g355) & (!sk[97]) & (g78)) + ((g20) & (!g355) & (sk[97]) & (g78)) + ((g20) & (g355) & (!sk[97]) & (!g78)) + ((g20) & (g355) & (!sk[97]) & (g78)));
	assign g452 = (((!g161) & (!g175) & (g177) & (!g278) & (!sk[98]) & (g451)) + ((!g161) & (!g175) & (g177) & (g278) & (!sk[98]) & (!g451)) + ((!g161) & (!g175) & (g177) & (g278) & (!sk[98]) & (g451)) + ((!g161) & (g175) & (!g177) & (!g278) & (!sk[98]) & (!g451)) + ((!g161) & (g175) & (!g177) & (!g278) & (!sk[98]) & (g451)) + ((!g161) & (g175) & (!g177) & (g278) & (!sk[98]) & (!g451)) + ((!g161) & (g175) & (!g177) & (g278) & (!sk[98]) & (g451)) + ((!g161) & (g175) & (g177) & (!g278) & (!sk[98]) & (!g451)) + ((!g161) & (g175) & (g177) & (!g278) & (!sk[98]) & (g451)) + ((!g161) & (g175) & (g177) & (g278) & (!sk[98]) & (!g451)) + ((!g161) & (g175) & (g177) & (g278) & (!sk[98]) & (g451)) + ((g161) & (!g175) & (!g177) & (!g278) & (sk[98]) & (!g451)) + ((g161) & (!g175) & (!g177) & (g278) & (sk[98]) & (!g451)) + ((g161) & (!g175) & (!g177) & (g278) & (sk[98]) & (g451)) + ((g161) & (!g175) & (g177) & (!g278) & (!sk[98]) & (g451)) + ((g161) & (!g175) & (g177) & (!g278) & (sk[98]) & (!g451)) + ((g161) & (!g175) & (g177) & (!g278) & (sk[98]) & (g451)) + ((g161) & (!g175) & (g177) & (g278) & (!sk[98]) & (!g451)) + ((g161) & (!g175) & (g177) & (g278) & (!sk[98]) & (g451)) + ((g161) & (!g175) & (g177) & (g278) & (sk[98]) & (!g451)) + ((g161) & (!g175) & (g177) & (g278) & (sk[98]) & (g451)) + ((g161) & (g175) & (!g177) & (!g278) & (!sk[98]) & (!g451)) + ((g161) & (g175) & (!g177) & (!g278) & (!sk[98]) & (g451)) + ((g161) & (g175) & (!g177) & (!g278) & (sk[98]) & (!g451)) + ((g161) & (g175) & (!g177) & (!g278) & (sk[98]) & (g451)) + ((g161) & (g175) & (!g177) & (g278) & (!sk[98]) & (!g451)) + ((g161) & (g175) & (!g177) & (g278) & (!sk[98]) & (g451)) + ((g161) & (g175) & (!g177) & (g278) & (sk[98]) & (!g451)) + ((g161) & (g175) & (!g177) & (g278) & (sk[98]) & (g451)) + ((g161) & (g175) & (g177) & (!g278) & (!sk[98]) & (!g451)) + ((g161) & (g175) & (g177) & (!g278) & (!sk[98]) & (g451)) + ((g161) & (g175) & (g177) & (!g278) & (sk[98]) & (!g451)) + ((g161) & (g175) & (g177) & (!g278) & (sk[98]) & (g451)) + ((g161) & (g175) & (g177) & (g278) & (!sk[98]) & (!g451)) + ((g161) & (g175) & (g177) & (g278) & (!sk[98]) & (g451)) + ((g161) & (g175) & (g177) & (g278) & (sk[98]) & (!g451)) + ((g161) & (g175) & (g177) & (g278) & (sk[98]) & (g451)));
	assign g453 = (((!g109) & (!g157) & (!sk[99]) & (g186) & (!g192) & (g452)) + ((!g109) & (!g157) & (!sk[99]) & (g186) & (g192) & (!g452)) + ((!g109) & (!g157) & (!sk[99]) & (g186) & (g192) & (g452)) + ((!g109) & (!g157) & (sk[99]) & (!g186) & (!g192) & (!g452)) + ((!g109) & (!g157) & (sk[99]) & (!g186) & (g192) & (!g452)) + ((!g109) & (!g157) & (sk[99]) & (g186) & (!g192) & (!g452)) + ((!g109) & (!g157) & (sk[99]) & (g186) & (g192) & (!g452)) + ((!g109) & (g157) & (!sk[99]) & (!g186) & (!g192) & (!g452)) + ((!g109) & (g157) & (!sk[99]) & (!g186) & (!g192) & (g452)) + ((!g109) & (g157) & (!sk[99]) & (!g186) & (g192) & (!g452)) + ((!g109) & (g157) & (!sk[99]) & (!g186) & (g192) & (g452)) + ((!g109) & (g157) & (!sk[99]) & (g186) & (!g192) & (!g452)) + ((!g109) & (g157) & (!sk[99]) & (g186) & (!g192) & (g452)) + ((!g109) & (g157) & (!sk[99]) & (g186) & (g192) & (!g452)) + ((!g109) & (g157) & (!sk[99]) & (g186) & (g192) & (g452)) + ((!g109) & (g157) & (sk[99]) & (!g186) & (!g192) & (!g452)) + ((g109) & (!g157) & (!sk[99]) & (g186) & (!g192) & (g452)) + ((g109) & (!g157) & (!sk[99]) & (g186) & (g192) & (!g452)) + ((g109) & (!g157) & (!sk[99]) & (g186) & (g192) & (g452)) + ((g109) & (!g157) & (sk[99]) & (!g186) & (!g192) & (!g452)) + ((g109) & (!g157) & (sk[99]) & (!g186) & (g192) & (!g452)) + ((g109) & (!g157) & (sk[99]) & (g186) & (!g192) & (!g452)) + ((g109) & (!g157) & (sk[99]) & (g186) & (g192) & (!g452)) + ((g109) & (g157) & (!sk[99]) & (!g186) & (!g192) & (!g452)) + ((g109) & (g157) & (!sk[99]) & (!g186) & (!g192) & (g452)) + ((g109) & (g157) & (!sk[99]) & (!g186) & (g192) & (!g452)) + ((g109) & (g157) & (!sk[99]) & (!g186) & (g192) & (g452)) + ((g109) & (g157) & (!sk[99]) & (g186) & (!g192) & (!g452)) + ((g109) & (g157) & (!sk[99]) & (g186) & (!g192) & (g452)) + ((g109) & (g157) & (!sk[99]) & (g186) & (g192) & (!g452)) + ((g109) & (g157) & (!sk[99]) & (g186) & (g192) & (g452)));
	assign g454 = (((!i_8_) & (!sk[100]) & (!g392) & (g449) & (!g450) & (g453)) + ((!i_8_) & (!sk[100]) & (!g392) & (g449) & (g450) & (!g453)) + ((!i_8_) & (!sk[100]) & (!g392) & (g449) & (g450) & (g453)) + ((!i_8_) & (!sk[100]) & (g392) & (!g449) & (!g450) & (!g453)) + ((!i_8_) & (!sk[100]) & (g392) & (!g449) & (!g450) & (g453)) + ((!i_8_) & (!sk[100]) & (g392) & (!g449) & (g450) & (!g453)) + ((!i_8_) & (!sk[100]) & (g392) & (!g449) & (g450) & (g453)) + ((!i_8_) & (!sk[100]) & (g392) & (g449) & (!g450) & (!g453)) + ((!i_8_) & (!sk[100]) & (g392) & (g449) & (!g450) & (g453)) + ((!i_8_) & (!sk[100]) & (g392) & (g449) & (g450) & (!g453)) + ((!i_8_) & (!sk[100]) & (g392) & (g449) & (g450) & (g453)) + ((!i_8_) & (sk[100]) & (!g392) & (!g449) & (!g450) & (g453)) + ((!i_8_) & (sk[100]) & (!g392) & (!g449) & (g450) & (g453)) + ((!i_8_) & (sk[100]) & (!g392) & (g449) & (!g450) & (g453)) + ((!i_8_) & (sk[100]) & (!g392) & (g449) & (g450) & (g453)) + ((!i_8_) & (sk[100]) & (g392) & (g449) & (!g450) & (g453)) + ((!i_8_) & (sk[100]) & (g392) & (g449) & (g450) & (g453)) + ((i_8_) & (!sk[100]) & (!g392) & (g449) & (!g450) & (g453)) + ((i_8_) & (!sk[100]) & (!g392) & (g449) & (g450) & (!g453)) + ((i_8_) & (!sk[100]) & (!g392) & (g449) & (g450) & (g453)) + ((i_8_) & (!sk[100]) & (g392) & (!g449) & (!g450) & (!g453)) + ((i_8_) & (!sk[100]) & (g392) & (!g449) & (!g450) & (g453)) + ((i_8_) & (!sk[100]) & (g392) & (!g449) & (g450) & (!g453)) + ((i_8_) & (!sk[100]) & (g392) & (!g449) & (g450) & (g453)) + ((i_8_) & (!sk[100]) & (g392) & (g449) & (!g450) & (!g453)) + ((i_8_) & (!sk[100]) & (g392) & (g449) & (!g450) & (g453)) + ((i_8_) & (!sk[100]) & (g392) & (g449) & (g450) & (!g453)) + ((i_8_) & (!sk[100]) & (g392) & (g449) & (g450) & (g453)) + ((i_8_) & (sk[100]) & (!g392) & (!g449) & (!g450) & (g453)) + ((i_8_) & (sk[100]) & (!g392) & (!g449) & (g450) & (g453)) + ((i_8_) & (sk[100]) & (!g392) & (g449) & (!g450) & (g453)) + ((i_8_) & (sk[100]) & (!g392) & (g449) & (g450) & (g453)) + ((i_8_) & (sk[100]) & (g392) & (!g449) & (!g450) & (g453)) + ((i_8_) & (sk[100]) & (g392) & (g449) & (!g450) & (g453)));
	assign g455 = (((!g66) & (!g1584) & (g448) & (!sk[101]) & (!g454)) + ((!g66) & (!g1584) & (g448) & (!sk[101]) & (g454)) + ((!g66) & (g1584) & (g448) & (!sk[101]) & (!g454)) + ((!g66) & (g1584) & (g448) & (!sk[101]) & (g454)) + ((g66) & (!g1584) & (g448) & (!sk[101]) & (!g454)) + ((g66) & (!g1584) & (g448) & (!sk[101]) & (g454)) + ((g66) & (g1584) & (!g448) & (sk[101]) & (g454)) + ((g66) & (g1584) & (g448) & (!sk[101]) & (!g454)) + ((g66) & (g1584) & (g448) & (!sk[101]) & (g454)));
	assign g456 = (((g173) & (g269) & (g332) & (g412) & (g442) & (g455)));
	assign g457 = (((!i_0_) & (!i_1_) & (!sk[103]) & (g6)) + ((!i_0_) & (i_1_) & (!sk[103]) & (!g6)) + ((!i_0_) & (i_1_) & (!sk[103]) & (g6)) + ((i_0_) & (!i_1_) & (!sk[103]) & (g6)) + ((i_0_) & (!i_1_) & (sk[103]) & (g6)) + ((i_0_) & (i_1_) & (!sk[103]) & (!g6)) + ((i_0_) & (i_1_) & (!sk[103]) & (g6)));
	assign g458 = (((!g457) & (sk[104]) & (g51)) + ((g457) & (!sk[104]) & (!g51)) + ((g457) & (!sk[104]) & (g51)));
	assign g459 = (((!g24) & (!g74) & (!g91) & (sk[105]) & (g257)) + ((!g24) & (!g74) & (g91) & (!sk[105]) & (!g257)) + ((!g24) & (!g74) & (g91) & (!sk[105]) & (g257)) + ((!g24) & (g74) & (!g91) & (sk[105]) & (!g257)) + ((!g24) & (g74) & (!g91) & (sk[105]) & (g257)) + ((!g24) & (g74) & (g91) & (!sk[105]) & (!g257)) + ((!g24) & (g74) & (g91) & (!sk[105]) & (g257)) + ((g24) & (!g74) & (g91) & (!sk[105]) & (!g257)) + ((g24) & (!g74) & (g91) & (!sk[105]) & (g257)) + ((g24) & (g74) & (g91) & (!sk[105]) & (!g257)) + ((g24) & (g74) & (g91) & (!sk[105]) & (g257)));
	assign g460 = (((!i_12_) & (!sk[106]) & (!i_13_) & (i_14_)) + ((!i_12_) & (!sk[106]) & (i_13_) & (!i_14_)) + ((!i_12_) & (!sk[106]) & (i_13_) & (i_14_)) + ((!i_12_) & (sk[106]) & (!i_13_) & (!i_14_)) + ((!i_12_) & (sk[106]) & (!i_13_) & (i_14_)) + ((!i_12_) & (sk[106]) & (i_13_) & (!i_14_)) + ((!i_12_) & (sk[106]) & (i_13_) & (i_14_)) + ((i_12_) & (!sk[106]) & (!i_13_) & (i_14_)) + ((i_12_) & (!sk[106]) & (i_13_) & (!i_14_)) + ((i_12_) & (!sk[106]) & (i_13_) & (i_14_)) + ((i_12_) & (sk[106]) & (!i_13_) & (!i_14_)) + ((i_12_) & (sk[106]) & (!i_13_) & (i_14_)) + ((i_12_) & (sk[106]) & (i_13_) & (i_14_)));
	assign g461 = (((!sk[107]) & (g27) & (!g460)) + ((!sk[107]) & (g27) & (g460)) + ((sk[107]) & (g27) & (!g460)));
	assign g462 = (((!g75) & (!sk[108]) & (!g107) & (g460)) + ((!g75) & (!sk[108]) & (g107) & (!g460)) + ((!g75) & (!sk[108]) & (g107) & (g460)) + ((!g75) & (sk[108]) & (!g107) & (!g460)) + ((g75) & (!sk[108]) & (!g107) & (g460)) + ((g75) & (!sk[108]) & (g107) & (!g460)) + ((g75) & (!sk[108]) & (g107) & (g460)));
	assign g463 = (((!i_8_) & (!g27) & (g73) & (!g86) & (!sk[109]) & (g460)) + ((!i_8_) & (!g27) & (g73) & (g86) & (!sk[109]) & (!g460)) + ((!i_8_) & (!g27) & (g73) & (g86) & (!sk[109]) & (g460)) + ((!i_8_) & (!g27) & (g73) & (g86) & (sk[109]) & (!g460)) + ((!i_8_) & (g27) & (!g73) & (!g86) & (!sk[109]) & (!g460)) + ((!i_8_) & (g27) & (!g73) & (!g86) & (!sk[109]) & (g460)) + ((!i_8_) & (g27) & (!g73) & (g86) & (!sk[109]) & (!g460)) + ((!i_8_) & (g27) & (!g73) & (g86) & (!sk[109]) & (g460)) + ((!i_8_) & (g27) & (g73) & (!g86) & (!sk[109]) & (!g460)) + ((!i_8_) & (g27) & (g73) & (!g86) & (!sk[109]) & (g460)) + ((!i_8_) & (g27) & (g73) & (!g86) & (sk[109]) & (!g460)) + ((!i_8_) & (g27) & (g73) & (g86) & (!sk[109]) & (!g460)) + ((!i_8_) & (g27) & (g73) & (g86) & (!sk[109]) & (g460)) + ((!i_8_) & (g27) & (g73) & (g86) & (sk[109]) & (!g460)) + ((i_8_) & (!g27) & (g73) & (!g86) & (!sk[109]) & (g460)) + ((i_8_) & (!g27) & (g73) & (g86) & (!sk[109]) & (!g460)) + ((i_8_) & (!g27) & (g73) & (g86) & (!sk[109]) & (g460)) + ((i_8_) & (g27) & (!g73) & (!g86) & (!sk[109]) & (!g460)) + ((i_8_) & (g27) & (!g73) & (!g86) & (!sk[109]) & (g460)) + ((i_8_) & (g27) & (!g73) & (g86) & (!sk[109]) & (!g460)) + ((i_8_) & (g27) & (!g73) & (g86) & (!sk[109]) & (g460)) + ((i_8_) & (g27) & (g73) & (!g86) & (!sk[109]) & (!g460)) + ((i_8_) & (g27) & (g73) & (!g86) & (!sk[109]) & (g460)) + ((i_8_) & (g27) & (g73) & (!g86) & (sk[109]) & (!g460)) + ((i_8_) & (g27) & (g73) & (g86) & (!sk[109]) & (!g460)) + ((i_8_) & (g27) & (g73) & (g86) & (!sk[109]) & (g460)) + ((i_8_) & (g27) & (g73) & (g86) & (sk[109]) & (!g460)));
	assign g464 = (((!i_8_) & (!g3) & (g73) & (!sk[110]) & (!g83) & (g460)) + ((!i_8_) & (!g3) & (g73) & (!sk[110]) & (g83) & (!g460)) + ((!i_8_) & (!g3) & (g73) & (!sk[110]) & (g83) & (g460)) + ((!i_8_) & (!g3) & (g73) & (sk[110]) & (g83) & (!g460)) + ((!i_8_) & (g3) & (!g73) & (!sk[110]) & (!g83) & (!g460)) + ((!i_8_) & (g3) & (!g73) & (!sk[110]) & (!g83) & (g460)) + ((!i_8_) & (g3) & (!g73) & (!sk[110]) & (g83) & (!g460)) + ((!i_8_) & (g3) & (!g73) & (!sk[110]) & (g83) & (g460)) + ((!i_8_) & (g3) & (g73) & (!sk[110]) & (!g83) & (!g460)) + ((!i_8_) & (g3) & (g73) & (!sk[110]) & (!g83) & (g460)) + ((!i_8_) & (g3) & (g73) & (!sk[110]) & (g83) & (!g460)) + ((!i_8_) & (g3) & (g73) & (!sk[110]) & (g83) & (g460)) + ((!i_8_) & (g3) & (g73) & (sk[110]) & (g83) & (!g460)) + ((i_8_) & (!g3) & (g73) & (!sk[110]) & (!g83) & (g460)) + ((i_8_) & (!g3) & (g73) & (!sk[110]) & (g83) & (!g460)) + ((i_8_) & (!g3) & (g73) & (!sk[110]) & (g83) & (g460)) + ((i_8_) & (!g3) & (g73) & (sk[110]) & (g83) & (!g460)) + ((i_8_) & (g3) & (!g73) & (!sk[110]) & (!g83) & (!g460)) + ((i_8_) & (g3) & (!g73) & (!sk[110]) & (!g83) & (g460)) + ((i_8_) & (g3) & (!g73) & (!sk[110]) & (g83) & (!g460)) + ((i_8_) & (g3) & (!g73) & (!sk[110]) & (g83) & (g460)) + ((i_8_) & (g3) & (g73) & (!sk[110]) & (!g83) & (!g460)) + ((i_8_) & (g3) & (g73) & (!sk[110]) & (!g83) & (g460)) + ((i_8_) & (g3) & (g73) & (!sk[110]) & (g83) & (!g460)) + ((i_8_) & (g3) & (g73) & (!sk[110]) & (g83) & (g460)) + ((i_8_) & (g3) & (g73) & (sk[110]) & (!g83) & (!g460)) + ((i_8_) & (g3) & (g73) & (sk[110]) & (g83) & (!g460)));
	assign g465 = (((!i_8_) & (!sk[111]) & (!g20) & (g35) & (!g73) & (g460)) + ((!i_8_) & (!sk[111]) & (!g20) & (g35) & (g73) & (!g460)) + ((!i_8_) & (!sk[111]) & (!g20) & (g35) & (g73) & (g460)) + ((!i_8_) & (!sk[111]) & (g20) & (!g35) & (!g73) & (!g460)) + ((!i_8_) & (!sk[111]) & (g20) & (!g35) & (!g73) & (g460)) + ((!i_8_) & (!sk[111]) & (g20) & (!g35) & (g73) & (!g460)) + ((!i_8_) & (!sk[111]) & (g20) & (!g35) & (g73) & (g460)) + ((!i_8_) & (!sk[111]) & (g20) & (g35) & (!g73) & (!g460)) + ((!i_8_) & (!sk[111]) & (g20) & (g35) & (!g73) & (g460)) + ((!i_8_) & (!sk[111]) & (g20) & (g35) & (g73) & (!g460)) + ((!i_8_) & (!sk[111]) & (g20) & (g35) & (g73) & (g460)) + ((!i_8_) & (sk[111]) & (g20) & (!g35) & (g73) & (!g460)) + ((!i_8_) & (sk[111]) & (g20) & (g35) & (g73) & (!g460)) + ((i_8_) & (!sk[111]) & (!g20) & (g35) & (!g73) & (g460)) + ((i_8_) & (!sk[111]) & (!g20) & (g35) & (g73) & (!g460)) + ((i_8_) & (!sk[111]) & (!g20) & (g35) & (g73) & (g460)) + ((i_8_) & (!sk[111]) & (g20) & (!g35) & (!g73) & (!g460)) + ((i_8_) & (!sk[111]) & (g20) & (!g35) & (!g73) & (g460)) + ((i_8_) & (!sk[111]) & (g20) & (!g35) & (g73) & (!g460)) + ((i_8_) & (!sk[111]) & (g20) & (!g35) & (g73) & (g460)) + ((i_8_) & (!sk[111]) & (g20) & (g35) & (!g73) & (!g460)) + ((i_8_) & (!sk[111]) & (g20) & (g35) & (!g73) & (g460)) + ((i_8_) & (!sk[111]) & (g20) & (g35) & (g73) & (!g460)) + ((i_8_) & (!sk[111]) & (g20) & (g35) & (g73) & (g460)) + ((i_8_) & (sk[111]) & (!g20) & (g35) & (g73) & (!g460)) + ((i_8_) & (sk[111]) & (g20) & (!g35) & (g73) & (!g460)) + ((i_8_) & (sk[111]) & (g20) & (g35) & (g73) & (!g460)));
	assign g466 = (((!i_8_) & (!sk[112]) & (!g73) & (g107) & (!g353) & (g460)) + ((!i_8_) & (!sk[112]) & (!g73) & (g107) & (g353) & (!g460)) + ((!i_8_) & (!sk[112]) & (!g73) & (g107) & (g353) & (g460)) + ((!i_8_) & (!sk[112]) & (g73) & (!g107) & (!g353) & (!g460)) + ((!i_8_) & (!sk[112]) & (g73) & (!g107) & (!g353) & (g460)) + ((!i_8_) & (!sk[112]) & (g73) & (!g107) & (g353) & (!g460)) + ((!i_8_) & (!sk[112]) & (g73) & (!g107) & (g353) & (g460)) + ((!i_8_) & (!sk[112]) & (g73) & (g107) & (!g353) & (!g460)) + ((!i_8_) & (!sk[112]) & (g73) & (g107) & (!g353) & (g460)) + ((!i_8_) & (!sk[112]) & (g73) & (g107) & (g353) & (!g460)) + ((!i_8_) & (!sk[112]) & (g73) & (g107) & (g353) & (g460)) + ((!i_8_) & (sk[112]) & (g73) & (!g107) & (!g353) & (!g460)) + ((!i_8_) & (sk[112]) & (g73) & (!g107) & (g353) & (!g460)) + ((!i_8_) & (sk[112]) & (g73) & (g107) & (g353) & (!g460)) + ((i_8_) & (!sk[112]) & (!g73) & (g107) & (!g353) & (g460)) + ((i_8_) & (!sk[112]) & (!g73) & (g107) & (g353) & (!g460)) + ((i_8_) & (!sk[112]) & (!g73) & (g107) & (g353) & (g460)) + ((i_8_) & (!sk[112]) & (g73) & (!g107) & (!g353) & (!g460)) + ((i_8_) & (!sk[112]) & (g73) & (!g107) & (!g353) & (g460)) + ((i_8_) & (!sk[112]) & (g73) & (!g107) & (g353) & (!g460)) + ((i_8_) & (!sk[112]) & (g73) & (!g107) & (g353) & (g460)) + ((i_8_) & (!sk[112]) & (g73) & (g107) & (!g353) & (!g460)) + ((i_8_) & (!sk[112]) & (g73) & (g107) & (!g353) & (g460)) + ((i_8_) & (!sk[112]) & (g73) & (g107) & (g353) & (!g460)) + ((i_8_) & (!sk[112]) & (g73) & (g107) & (g353) & (g460)));
	assign g467 = (((!g463) & (!g464) & (!sk[113]) & (g465) & (!g466)) + ((!g463) & (!g464) & (!sk[113]) & (g465) & (g466)) + ((!g463) & (!g464) & (sk[113]) & (!g465) & (!g466)) + ((!g463) & (g464) & (!sk[113]) & (g465) & (!g466)) + ((!g463) & (g464) & (!sk[113]) & (g465) & (g466)) + ((g463) & (!g464) & (!sk[113]) & (g465) & (!g466)) + ((g463) & (!g464) & (!sk[113]) & (g465) & (g466)) + ((g463) & (g464) & (!sk[113]) & (g465) & (!g466)) + ((g463) & (g464) & (!sk[113]) & (g465) & (g466)));
	assign g468 = (((!g24) & (sk[114]) & (g69)) + ((g24) & (!sk[114]) & (!g69)) + ((g24) & (!sk[114]) & (g69)));
	assign g469 = (((!g3) & (!g460) & (!sk[115]) & (g468)) + ((!g3) & (!g460) & (sk[115]) & (!g468)) + ((!g3) & (g460) & (!sk[115]) & (!g468)) + ((!g3) & (g460) & (!sk[115]) & (g468)) + ((!g3) & (g460) & (sk[115]) & (!g468)) + ((g3) & (!g460) & (!sk[115]) & (g468)) + ((g3) & (g460) & (!sk[115]) & (!g468)) + ((g3) & (g460) & (!sk[115]) & (g468)) + ((g3) & (g460) & (sk[115]) & (!g468)));
	assign g470 = (((!g121) & (!g213) & (!sk[116]) & (g469)) + ((!g121) & (g213) & (!sk[116]) & (!g469)) + ((!g121) & (g213) & (!sk[116]) & (g469)) + ((!g121) & (g213) & (sk[116]) & (!g469)) + ((g121) & (!g213) & (!sk[116]) & (g469)) + ((g121) & (!g213) & (sk[116]) & (!g469)) + ((g121) & (g213) & (!sk[116]) & (!g469)) + ((g121) & (g213) & (!sk[116]) & (g469)) + ((g121) & (g213) & (sk[116]) & (!g469)));
	assign g471 = (((!sk[117]) & (!g161) & (!g86) & (g460)) + ((!sk[117]) & (!g161) & (g86) & (!g460)) + ((!sk[117]) & (!g161) & (g86) & (g460)) + ((!sk[117]) & (g161) & (!g86) & (g460)) + ((!sk[117]) & (g161) & (g86) & (!g460)) + ((!sk[117]) & (g161) & (g86) & (g460)) + ((sk[117]) & (g161) & (g86) & (!g460)));
	assign g472 = (((!g20) & (!g27) & (g83) & (!sk[118]) & (!g460)) + ((!g20) & (!g27) & (g83) & (!sk[118]) & (g460)) + ((!g20) & (!g27) & (g83) & (sk[118]) & (!g460)) + ((!g20) & (g27) & (!g83) & (sk[118]) & (!g460)) + ((!g20) & (g27) & (g83) & (!sk[118]) & (!g460)) + ((!g20) & (g27) & (g83) & (!sk[118]) & (g460)) + ((!g20) & (g27) & (g83) & (sk[118]) & (!g460)) + ((g20) & (!g27) & (!g83) & (sk[118]) & (!g460)) + ((g20) & (!g27) & (g83) & (!sk[118]) & (!g460)) + ((g20) & (!g27) & (g83) & (!sk[118]) & (g460)) + ((g20) & (!g27) & (g83) & (sk[118]) & (!g460)) + ((g20) & (g27) & (!g83) & (sk[118]) & (!g460)) + ((g20) & (g27) & (g83) & (!sk[118]) & (!g460)) + ((g20) & (g27) & (g83) & (!sk[118]) & (g460)) + ((g20) & (g27) & (g83) & (sk[118]) & (!g460)));
	assign g473 = (((!sk[119]) & (g24) & (!g81)) + ((!sk[119]) & (g24) & (g81)) + ((sk[119]) & (!g24) & (g81)));
	assign g474 = (((!sk[120]) & (!g157) & (!g86) & (g460) & (!g473)) + ((!sk[120]) & (!g157) & (!g86) & (g460) & (g473)) + ((!sk[120]) & (!g157) & (g86) & (g460) & (!g473)) + ((!sk[120]) & (!g157) & (g86) & (g460) & (g473)) + ((!sk[120]) & (g157) & (!g86) & (g460) & (!g473)) + ((!sk[120]) & (g157) & (!g86) & (g460) & (g473)) + ((!sk[120]) & (g157) & (g86) & (g460) & (!g473)) + ((!sk[120]) & (g157) & (g86) & (g460) & (g473)) + ((sk[120]) & (g157) & (!g86) & (!g460) & (g473)) + ((sk[120]) & (g157) & (!g86) & (g460) & (g473)) + ((sk[120]) & (g157) & (g86) & (!g460) & (!g473)) + ((sk[120]) & (g157) & (g86) & (!g460) & (g473)) + ((sk[120]) & (g157) & (g86) & (g460) & (g473)));
	assign g475 = (((!i_8_) & (!g73) & (g86) & (!sk[121]) & (!g126) & (g460)) + ((!i_8_) & (!g73) & (g86) & (!sk[121]) & (g126) & (!g460)) + ((!i_8_) & (!g73) & (g86) & (!sk[121]) & (g126) & (g460)) + ((!i_8_) & (g73) & (!g86) & (!sk[121]) & (!g126) & (!g460)) + ((!i_8_) & (g73) & (!g86) & (!sk[121]) & (!g126) & (g460)) + ((!i_8_) & (g73) & (!g86) & (!sk[121]) & (g126) & (!g460)) + ((!i_8_) & (g73) & (!g86) & (!sk[121]) & (g126) & (g460)) + ((!i_8_) & (g73) & (!g86) & (sk[121]) & (!g126) & (!g460)) + ((!i_8_) & (g73) & (g86) & (!sk[121]) & (!g126) & (!g460)) + ((!i_8_) & (g73) & (g86) & (!sk[121]) & (!g126) & (g460)) + ((!i_8_) & (g73) & (g86) & (!sk[121]) & (g126) & (!g460)) + ((!i_8_) & (g73) & (g86) & (!sk[121]) & (g126) & (g460)) + ((!i_8_) & (g73) & (g86) & (sk[121]) & (!g126) & (!g460)) + ((i_8_) & (!g73) & (g86) & (!sk[121]) & (!g126) & (g460)) + ((i_8_) & (!g73) & (g86) & (!sk[121]) & (g126) & (!g460)) + ((i_8_) & (!g73) & (g86) & (!sk[121]) & (g126) & (g460)) + ((i_8_) & (g73) & (!g86) & (!sk[121]) & (!g126) & (!g460)) + ((i_8_) & (g73) & (!g86) & (!sk[121]) & (!g126) & (g460)) + ((i_8_) & (g73) & (!g86) & (!sk[121]) & (g126) & (!g460)) + ((i_8_) & (g73) & (!g86) & (!sk[121]) & (g126) & (g460)) + ((i_8_) & (g73) & (!g86) & (sk[121]) & (!g126) & (!g460)) + ((i_8_) & (g73) & (g86) & (!sk[121]) & (!g126) & (!g460)) + ((i_8_) & (g73) & (g86) & (!sk[121]) & (!g126) & (g460)) + ((i_8_) & (g73) & (g86) & (!sk[121]) & (g126) & (!g460)) + ((i_8_) & (g73) & (g86) & (!sk[121]) & (g126) & (g460)) + ((i_8_) & (g73) & (g86) & (sk[121]) & (!g126) & (!g460)) + ((i_8_) & (g73) & (g86) & (sk[121]) & (g126) & (!g460)));
	assign g476 = (((!g142) & (!g470) & (!g471) & (!g472) & (!g474) & (!g475)) + ((g142) & (!g470) & (!g471) & (!g472) & (!g474) & (!g475)) + ((g142) & (!g470) & (!g471) & (g472) & (!g474) & (!g475)));
	assign g477 = (((g17) & (!sk[123]) & (!g24)) + ((g17) & (!sk[123]) & (g24)) + ((g17) & (sk[123]) & (!g24)));
	assign g478 = (((g80) & (!i_11_) & (!i_15_) & (g119) & (!g392) & (!g460)) + ((g80) & (!i_11_) & (!i_15_) & (g119) & (g392) & (!g460)) + ((g80) & (i_11_) & (!i_15_) & (!g119) & (g392) & (!g460)) + ((g80) & (i_11_) & (!i_15_) & (g119) & (g392) & (!g460)));
	assign g479 = (((!g225) & (!sk[125]) & (!g213) & (g477) & (!g478)) + ((!g225) & (!sk[125]) & (!g213) & (g477) & (g478)) + ((!g225) & (!sk[125]) & (g213) & (g477) & (!g478)) + ((!g225) & (!sk[125]) & (g213) & (g477) & (g478)) + ((!g225) & (sk[125]) & (!g213) & (!g477) & (!g478)) + ((!g225) & (sk[125]) & (!g213) & (g477) & (!g478)) + ((!g225) & (sk[125]) & (g213) & (!g477) & (!g478)) + ((g225) & (!sk[125]) & (!g213) & (g477) & (!g478)) + ((g225) & (!sk[125]) & (!g213) & (g477) & (g478)) + ((g225) & (!sk[125]) & (g213) & (g477) & (!g478)) + ((g225) & (!sk[125]) & (g213) & (g477) & (g478)) + ((g225) & (sk[125]) & (!g213) & (!g477) & (!g478)) + ((g225) & (sk[125]) & (g213) & (!g477) & (!g478)));
	assign g480 = (((!g167) & (!g461) & (!g462) & (g467) & (g476) & (g479)) + ((!g167) & (g461) & (!g462) & (g467) & (g476) & (g479)) + ((g167) & (!g461) & (!g462) & (g467) & (g476) & (g479)));
	assign g481 = (((!sk[127]) & (!g24) & (!g154) & (g91) & (!g175)) + ((!sk[127]) & (!g24) & (!g154) & (g91) & (g175)) + ((!sk[127]) & (!g24) & (g154) & (g91) & (!g175)) + ((!sk[127]) & (!g24) & (g154) & (g91) & (g175)) + ((!sk[127]) & (g24) & (!g154) & (g91) & (!g175)) + ((!sk[127]) & (g24) & (!g154) & (g91) & (g175)) + ((!sk[127]) & (g24) & (g154) & (g91) & (!g175)) + ((!sk[127]) & (g24) & (g154) & (g91) & (g175)) + ((sk[127]) & (!g24) & (!g154) & (!g91) & (!g175)) + ((sk[127]) & (!g24) & (!g154) & (!g91) & (g175)) + ((sk[127]) & (!g24) & (!g154) & (g91) & (g175)) + ((sk[127]) & (g24) & (!g154) & (!g91) & (g175)) + ((sk[127]) & (g24) & (!g154) & (g91) & (g175)));
	assign g482 = (((!i_12_) & (!sk[0]) & (!i_13_) & (i_14_)) + ((!i_12_) & (!sk[0]) & (i_13_) & (!i_14_)) + ((!i_12_) & (!sk[0]) & (i_13_) & (i_14_)) + ((!i_12_) & (sk[0]) & (!i_13_) & (i_14_)) + ((!i_12_) & (sk[0]) & (i_13_) & (i_14_)) + ((i_12_) & (!sk[0]) & (!i_13_) & (i_14_)) + ((i_12_) & (!sk[0]) & (i_13_) & (!i_14_)) + ((i_12_) & (!sk[0]) & (i_13_) & (i_14_)) + ((i_12_) & (sk[0]) & (!i_13_) & (i_14_)));
	assign g483 = (((!sk[1]) & (g36) & (!g482)) + ((!sk[1]) & (g36) & (g482)) + ((sk[1]) & (g36) & (g482)));
	assign g484 = (((!sk[2]) & (g91) & (!g482)) + ((!sk[2]) & (g91) & (g482)) + ((sk[2]) & (!g91) & (g482)));
	assign g485 = (((!sk[3]) & (!g159) & (!g154) & (g483) & (!g484)) + ((!sk[3]) & (!g159) & (!g154) & (g483) & (g484)) + ((!sk[3]) & (!g159) & (g154) & (g483) & (!g484)) + ((!sk[3]) & (!g159) & (g154) & (g483) & (g484)) + ((!sk[3]) & (g159) & (!g154) & (g483) & (!g484)) + ((!sk[3]) & (g159) & (!g154) & (g483) & (g484)) + ((!sk[3]) & (g159) & (g154) & (g483) & (!g484)) + ((!sk[3]) & (g159) & (g154) & (g483) & (g484)) + ((sk[3]) & (!g159) & (!g154) & (!g483) & (g484)) + ((sk[3]) & (!g159) & (!g154) & (g483) & (!g484)) + ((sk[3]) & (!g159) & (!g154) & (g483) & (g484)) + ((sk[3]) & (!g159) & (g154) & (!g483) & (g484)) + ((sk[3]) & (!g159) & (g154) & (g483) & (g484)) + ((sk[3]) & (g159) & (!g154) & (g483) & (!g484)) + ((sk[3]) & (g159) & (!g154) & (g483) & (g484)));
	assign g486 = (((!g91) & (sk[4]) & (!g460)) + ((g91) & (!sk[4]) & (!g460)) + ((g91) & (!sk[4]) & (g460)));
	assign g487 = (((!g91) & (sk[5]) & (!g174)) + ((g91) & (!sk[5]) & (!g174)) + ((g91) & (!sk[5]) & (g174)));
	assign g488 = (((!g102) & (!sk[6]) & (!g105) & (g486) & (!g487)) + ((!g102) & (!sk[6]) & (!g105) & (g486) & (g487)) + ((!g102) & (!sk[6]) & (g105) & (g486) & (!g487)) + ((!g102) & (!sk[6]) & (g105) & (g486) & (g487)) + ((!g102) & (sk[6]) & (!g105) & (g486) & (!g487)) + ((!g102) & (sk[6]) & (!g105) & (g486) & (g487)) + ((g102) & (!sk[6]) & (!g105) & (g486) & (!g487)) + ((g102) & (!sk[6]) & (!g105) & (g486) & (g487)) + ((g102) & (!sk[6]) & (g105) & (g486) & (!g487)) + ((g102) & (!sk[6]) & (g105) & (g486) & (g487)) + ((g102) & (sk[6]) & (!g105) & (!g486) & (g487)) + ((g102) & (sk[6]) & (!g105) & (g486) & (!g487)) + ((g102) & (sk[6]) & (!g105) & (g486) & (g487)) + ((g102) & (sk[6]) & (g105) & (!g486) & (g487)) + ((g102) & (sk[6]) & (g105) & (g486) & (g487)));
	assign g489 = (((g17) & (!sk[7]) & (!g482)) + ((g17) & (!sk[7]) & (g482)) + ((g17) & (sk[7]) & (g482)));
	assign g490 = (((!g105) & (!g253) & (!g200) & (!g212) & (!g356) & (!g489)) + ((!g105) & (!g253) & (!g200) & (!g212) & (g356) & (!g489)) + ((!g105) & (g253) & (!g200) & (!g212) & (!g356) & (!g489)) + ((!g105) & (g253) & (!g200) & (!g212) & (g356) & (!g489)) + ((!g105) & (g253) & (g200) & (!g212) & (!g356) & (!g489)) + ((g105) & (!g253) & (!g200) & (!g212) & (!g356) & (!g489)) + ((g105) & (!g253) & (!g200) & (!g212) & (!g356) & (g489)) + ((g105) & (!g253) & (!g200) & (!g212) & (g356) & (!g489)) + ((g105) & (!g253) & (!g200) & (!g212) & (g356) & (g489)) + ((g105) & (!g253) & (!g200) & (g212) & (!g356) & (!g489)) + ((g105) & (!g253) & (!g200) & (g212) & (!g356) & (g489)) + ((g105) & (!g253) & (!g200) & (g212) & (g356) & (!g489)) + ((g105) & (!g253) & (!g200) & (g212) & (g356) & (g489)) + ((g105) & (g253) & (!g200) & (!g212) & (!g356) & (!g489)) + ((g105) & (g253) & (!g200) & (!g212) & (!g356) & (g489)) + ((g105) & (g253) & (!g200) & (!g212) & (g356) & (!g489)) + ((g105) & (g253) & (!g200) & (!g212) & (g356) & (g489)) + ((g105) & (g253) & (!g200) & (g212) & (!g356) & (!g489)) + ((g105) & (g253) & (!g200) & (g212) & (!g356) & (g489)) + ((g105) & (g253) & (!g200) & (g212) & (g356) & (!g489)) + ((g105) & (g253) & (!g200) & (g212) & (g356) & (g489)) + ((g105) & (g253) & (g200) & (!g212) & (!g356) & (!g489)) + ((g105) & (g253) & (g200) & (!g212) & (!g356) & (g489)) + ((g105) & (g253) & (g200) & (g212) & (!g356) & (!g489)) + ((g105) & (g253) & (g200) & (g212) & (!g356) & (g489)));
	assign g491 = (((!sk[9]) & (!g481) & (!g485) & (g488) & (!g490)) + ((!sk[9]) & (!g481) & (!g485) & (g488) & (g490)) + ((!sk[9]) & (!g481) & (g485) & (g488) & (!g490)) + ((!sk[9]) & (!g481) & (g485) & (g488) & (g490)) + ((!sk[9]) & (g481) & (!g485) & (g488) & (!g490)) + ((!sk[9]) & (g481) & (!g485) & (g488) & (g490)) + ((!sk[9]) & (g481) & (g485) & (g488) & (!g490)) + ((!sk[9]) & (g481) & (g485) & (g488) & (g490)) + ((sk[9]) & (!g481) & (!g485) & (!g488) & (g490)));
	assign g492 = (((!sk[10]) & (!g24) & (!g36) & (g91) & (!g88)) + ((!sk[10]) & (!g24) & (!g36) & (g91) & (g88)) + ((!sk[10]) & (!g24) & (g36) & (g91) & (!g88)) + ((!sk[10]) & (!g24) & (g36) & (g91) & (g88)) + ((!sk[10]) & (g24) & (!g36) & (g91) & (!g88)) + ((!sk[10]) & (g24) & (!g36) & (g91) & (g88)) + ((!sk[10]) & (g24) & (g36) & (g91) & (!g88)) + ((!sk[10]) & (g24) & (g36) & (g91) & (g88)) + ((sk[10]) & (!g24) & (!g36) & (!g91) & (!g88)) + ((sk[10]) & (!g24) & (!g36) & (!g91) & (g88)) + ((sk[10]) & (!g24) & (!g36) & (g91) & (g88)) + ((sk[10]) & (!g24) & (g36) & (!g91) & (!g88)) + ((sk[10]) & (!g24) & (g36) & (!g91) & (g88)) + ((sk[10]) & (!g24) & (g36) & (g91) & (!g88)) + ((sk[10]) & (!g24) & (g36) & (g91) & (g88)));
	assign g493 = (((!g165) & (!g131) & (!g257) & (!g383) & (!g477) & (!g492)) + ((!g165) & (!g131) & (!g257) & (g383) & (!g477) & (!g492)) + ((!g165) & (!g131) & (g257) & (!g383) & (!g477) & (!g492)) + ((!g165) & (!g131) & (g257) & (g383) & (!g477) & (!g492)) + ((!g165) & (g131) & (!g257) & (!g383) & (!g477) & (!g492)) + ((!g165) & (g131) & (!g257) & (!g383) & (!g477) & (g492)) + ((!g165) & (g131) & (!g257) & (g383) & (!g477) & (!g492)) + ((!g165) & (g131) & (!g257) & (g383) & (!g477) & (g492)) + ((!g165) & (g131) & (!g257) & (g383) & (g477) & (!g492)) + ((!g165) & (g131) & (!g257) & (g383) & (g477) & (g492)) + ((!g165) & (g131) & (g257) & (!g383) & (!g477) & (!g492)) + ((!g165) & (g131) & (g257) & (!g383) & (!g477) & (g492)) + ((!g165) & (g131) & (g257) & (g383) & (!g477) & (!g492)) + ((!g165) & (g131) & (g257) & (g383) & (!g477) & (g492)) + ((g165) & (!g131) & (!g257) & (!g383) & (!g477) & (!g492)) + ((g165) & (!g131) & (!g257) & (g383) & (!g477) & (!g492)) + ((g165) & (!g131) & (g257) & (!g383) & (!g477) & (!g492)) + ((g165) & (!g131) & (g257) & (g383) & (!g477) & (!g492)) + ((g165) & (g131) & (!g257) & (!g383) & (!g477) & (!g492)) + ((g165) & (g131) & (!g257) & (g383) & (!g477) & (!g492)) + ((g165) & (g131) & (g257) & (!g383) & (!g477) & (!g492)) + ((g165) & (g131) & (g257) & (g383) & (!g477) & (!g492)));
	assign g494 = (((!i_9_) & (!i_10_) & (!i_11_) & (!i_15_) & (!g174) & (!g460)) + ((!i_9_) & (!i_10_) & (!i_11_) & (!i_15_) & (g174) & (!g460)) + ((!i_9_) & (!i_10_) & (i_11_) & (!i_15_) & (!g174) & (!g460)) + ((!i_9_) & (!i_10_) & (i_11_) & (!i_15_) & (g174) & (!g460)) + ((!i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (!g174) & (!g460)) + ((!i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (g174) & (!g460)) + ((!i_9_) & (i_10_) & (!i_11_) & (i_15_) & (!g174) & (!g460)) + ((!i_9_) & (i_10_) & (!i_11_) & (i_15_) & (g174) & (!g460)) + ((!i_9_) & (i_10_) & (i_11_) & (!i_15_) & (!g174) & (!g460)) + ((!i_9_) & (i_10_) & (i_11_) & (!i_15_) & (g174) & (!g460)) + ((!i_9_) & (i_10_) & (i_11_) & (i_15_) & (!g174) & (!g460)) + ((!i_9_) & (i_10_) & (i_11_) & (i_15_) & (!g174) & (g460)) + ((!i_9_) & (i_10_) & (i_11_) & (i_15_) & (g174) & (!g460)) + ((i_9_) & (!i_10_) & (!i_11_) & (!i_15_) & (!g174) & (!g460)) + ((i_9_) & (!i_10_) & (!i_11_) & (!i_15_) & (g174) & (!g460)) + ((i_9_) & (!i_10_) & (i_11_) & (!i_15_) & (!g174) & (!g460)) + ((i_9_) & (!i_10_) & (i_11_) & (!i_15_) & (g174) & (!g460)) + ((i_9_) & (!i_10_) & (i_11_) & (i_15_) & (!g174) & (!g460)) + ((i_9_) & (!i_10_) & (i_11_) & (i_15_) & (g174) & (!g460)) + ((i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (!g174) & (!g460)) + ((i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (g174) & (!g460)) + ((i_9_) & (i_10_) & (!i_11_) & (i_15_) & (!g174) & (!g460)) + ((i_9_) & (i_10_) & (!i_11_) & (i_15_) & (!g174) & (g460)) + ((i_9_) & (i_10_) & (i_11_) & (!i_15_) & (!g174) & (!g460)) + ((i_9_) & (i_10_) & (i_11_) & (!i_15_) & (g174) & (!g460)));
	assign g495 = (((!g22) & (sk[13]) & (!g460)) + ((g22) & (!sk[13]) & (!g460)) + ((g22) & (!sk[13]) & (g460)));
	assign g496 = (((!g24) & (sk[14]) & (g88)) + ((g24) & (!sk[14]) & (!g88)) + ((g24) & (!sk[14]) & (g88)));
	assign g497 = (((!i_8_) & (!i_6_) & (!i_7_) & (g118) & (!g495) & (g496)) + ((!i_8_) & (!i_6_) & (!i_7_) & (g118) & (g495) & (g496)) + ((!i_8_) & (!i_6_) & (i_7_) & (g118) & (g495) & (!g496)));
	assign g498 = (((!g102) & (!g350) & (!g468) & (sk[16]) & (!g494) & (!g497)) + ((!g102) & (!g350) & (!g468) & (sk[16]) & (g494) & (!g497)) + ((!g102) & (!g350) & (g468) & (!sk[16]) & (!g494) & (g497)) + ((!g102) & (!g350) & (g468) & (!sk[16]) & (g494) & (!g497)) + ((!g102) & (!g350) & (g468) & (!sk[16]) & (g494) & (g497)) + ((!g102) & (!g350) & (g468) & (sk[16]) & (!g494) & (!g497)) + ((!g102) & (!g350) & (g468) & (sk[16]) & (g494) & (!g497)) + ((!g102) & (g350) & (!g468) & (!sk[16]) & (!g494) & (!g497)) + ((!g102) & (g350) & (!g468) & (!sk[16]) & (!g494) & (g497)) + ((!g102) & (g350) & (!g468) & (!sk[16]) & (g494) & (!g497)) + ((!g102) & (g350) & (!g468) & (!sk[16]) & (g494) & (g497)) + ((!g102) & (g350) & (!g468) & (sk[16]) & (!g494) & (!g497)) + ((!g102) & (g350) & (g468) & (!sk[16]) & (!g494) & (!g497)) + ((!g102) & (g350) & (g468) & (!sk[16]) & (!g494) & (g497)) + ((!g102) & (g350) & (g468) & (!sk[16]) & (g494) & (!g497)) + ((!g102) & (g350) & (g468) & (!sk[16]) & (g494) & (g497)) + ((g102) & (!g350) & (!g468) & (sk[16]) & (!g494) & (!g497)) + ((g102) & (!g350) & (!g468) & (sk[16]) & (g494) & (!g497)) + ((g102) & (!g350) & (g468) & (!sk[16]) & (!g494) & (g497)) + ((g102) & (!g350) & (g468) & (!sk[16]) & (g494) & (!g497)) + ((g102) & (!g350) & (g468) & (!sk[16]) & (g494) & (g497)) + ((g102) & (g350) & (!g468) & (!sk[16]) & (!g494) & (!g497)) + ((g102) & (g350) & (!g468) & (!sk[16]) & (!g494) & (g497)) + ((g102) & (g350) & (!g468) & (!sk[16]) & (g494) & (!g497)) + ((g102) & (g350) & (!g468) & (!sk[16]) & (g494) & (g497)) + ((g102) & (g350) & (!g468) & (sk[16]) & (!g494) & (!g497)) + ((g102) & (g350) & (g468) & (!sk[16]) & (!g494) & (!g497)) + ((g102) & (g350) & (g468) & (!sk[16]) & (!g494) & (g497)) + ((g102) & (g350) & (g468) & (!sk[16]) & (g494) & (!g497)) + ((g102) & (g350) & (g468) & (!sk[16]) & (g494) & (g497)));
	assign g499 = (((!g459) & (!g480) & (g491) & (!sk[17]) & (!g493) & (g498)) + ((!g459) & (!g480) & (g491) & (!sk[17]) & (g493) & (!g498)) + ((!g459) & (!g480) & (g491) & (!sk[17]) & (g493) & (g498)) + ((!g459) & (g480) & (!g491) & (!sk[17]) & (!g493) & (!g498)) + ((!g459) & (g480) & (!g491) & (!sk[17]) & (!g493) & (g498)) + ((!g459) & (g480) & (!g491) & (!sk[17]) & (g493) & (!g498)) + ((!g459) & (g480) & (!g491) & (!sk[17]) & (g493) & (g498)) + ((!g459) & (g480) & (g491) & (!sk[17]) & (!g493) & (!g498)) + ((!g459) & (g480) & (g491) & (!sk[17]) & (!g493) & (g498)) + ((!g459) & (g480) & (g491) & (!sk[17]) & (g493) & (!g498)) + ((!g459) & (g480) & (g491) & (!sk[17]) & (g493) & (g498)) + ((!g459) & (g480) & (g491) & (sk[17]) & (g493) & (g498)) + ((g459) & (!g480) & (g491) & (!sk[17]) & (!g493) & (g498)) + ((g459) & (!g480) & (g491) & (!sk[17]) & (g493) & (!g498)) + ((g459) & (!g480) & (g491) & (!sk[17]) & (g493) & (g498)) + ((g459) & (g480) & (!g491) & (!sk[17]) & (!g493) & (!g498)) + ((g459) & (g480) & (!g491) & (!sk[17]) & (!g493) & (g498)) + ((g459) & (g480) & (!g491) & (!sk[17]) & (g493) & (!g498)) + ((g459) & (g480) & (!g491) & (!sk[17]) & (g493) & (g498)) + ((g459) & (g480) & (g491) & (!sk[17]) & (!g493) & (!g498)) + ((g459) & (g480) & (g491) & (!sk[17]) & (!g493) & (g498)) + ((g459) & (g480) & (g491) & (!sk[17]) & (g493) & (!g498)) + ((g459) & (g480) & (g491) & (!sk[17]) & (g493) & (g498)));
	assign g500 = (((!i_12_) & (!i_13_) & (!sk[18]) & (i_14_) & (!g88)) + ((!i_12_) & (!i_13_) & (!sk[18]) & (i_14_) & (g88)) + ((!i_12_) & (!i_13_) & (sk[18]) & (i_14_) & (g88)) + ((!i_12_) & (i_13_) & (!sk[18]) & (i_14_) & (!g88)) + ((!i_12_) & (i_13_) & (!sk[18]) & (i_14_) & (g88)) + ((!i_12_) & (i_13_) & (sk[18]) & (i_14_) & (g88)) + ((i_12_) & (!i_13_) & (!sk[18]) & (i_14_) & (!g88)) + ((i_12_) & (!i_13_) & (!sk[18]) & (i_14_) & (g88)) + ((i_12_) & (!i_13_) & (sk[18]) & (i_14_) & (g88)) + ((i_12_) & (i_13_) & (!sk[18]) & (i_14_) & (!g88)) + ((i_12_) & (i_13_) & (!sk[18]) & (i_14_) & (g88)));
	assign g501 = (((g81) & (!sk[19]) & (!g460)) + ((g81) & (!sk[19]) & (g460)) + ((g81) & (sk[19]) & (!g460)));
	assign g502 = (((!g161) & (!sk[20]) & (!g183) & (g501) & (!g473)) + ((!g161) & (!sk[20]) & (!g183) & (g501) & (g473)) + ((!g161) & (!sk[20]) & (g183) & (g501) & (!g473)) + ((!g161) & (!sk[20]) & (g183) & (g501) & (g473)) + ((g161) & (!sk[20]) & (!g183) & (g501) & (!g473)) + ((g161) & (!sk[20]) & (!g183) & (g501) & (g473)) + ((g161) & (!sk[20]) & (g183) & (g501) & (!g473)) + ((g161) & (!sk[20]) & (g183) & (g501) & (g473)) + ((g161) & (sk[20]) & (!g183) & (!g501) & (g473)) + ((g161) & (sk[20]) & (!g183) & (g501) & (!g473)) + ((g161) & (sk[20]) & (!g183) & (g501) & (g473)) + ((g161) & (sk[20]) & (g183) & (!g501) & (!g473)) + ((g161) & (sk[20]) & (g183) & (!g501) & (g473)) + ((g161) & (sk[20]) & (g183) & (g501) & (!g473)) + ((g161) & (sk[20]) & (g183) & (g501) & (g473)));
	assign g503 = (((!g125) & (!g164) & (!g105) & (!g487) & (!g500) & (!g502)) + ((!g125) & (!g164) & (!g105) & (g487) & (!g500) & (!g502)) + ((!g125) & (!g164) & (g105) & (!g487) & (!g500) & (!g502)) + ((!g125) & (!g164) & (g105) & (!g487) & (g500) & (!g502)) + ((!g125) & (!g164) & (g105) & (g487) & (!g500) & (!g502)) + ((!g125) & (!g164) & (g105) & (g487) & (g500) & (!g502)) + ((!g125) & (g164) & (!g105) & (!g487) & (!g500) & (!g502)) + ((!g125) & (g164) & (!g105) & (g487) & (!g500) & (!g502)) + ((!g125) & (g164) & (g105) & (!g487) & (!g500) & (!g502)) + ((!g125) & (g164) & (g105) & (g487) & (!g500) & (!g502)) + ((g125) & (!g164) & (!g105) & (!g487) & (!g500) & (!g502)) + ((g125) & (!g164) & (g105) & (!g487) & (!g500) & (!g502)) + ((g125) & (!g164) & (g105) & (!g487) & (g500) & (!g502)) + ((g125) & (g164) & (!g105) & (!g487) & (!g500) & (!g502)) + ((g125) & (g164) & (g105) & (!g487) & (!g500) & (!g502)));
	assign g504 = (((!sk[22]) & (!g355) & (!g91) & (g212)) + ((!sk[22]) & (!g355) & (g91) & (!g212)) + ((!sk[22]) & (!g355) & (g91) & (g212)) + ((!sk[22]) & (g355) & (!g91) & (g212)) + ((!sk[22]) & (g355) & (g91) & (!g212)) + ((!sk[22]) & (g355) & (g91) & (g212)) + ((sk[22]) & (!g355) & (!g91) & (!g212)) + ((sk[22]) & (!g355) & (g91) & (!g212)) + ((sk[22]) & (g355) & (g91) & (!g212)));
	assign g505 = (((!g157) & (!sk[23]) & (!g186) & (g192)) + ((!g157) & (!sk[23]) & (g186) & (!g192)) + ((!g157) & (!sk[23]) & (g186) & (g192)) + ((g157) & (!sk[23]) & (!g186) & (g192)) + ((g157) & (!sk[23]) & (g186) & (!g192)) + ((g157) & (!sk[23]) & (g186) & (g192)) + ((g157) & (sk[23]) & (!g186) & (g192)) + ((g157) & (sk[23]) & (g186) & (!g192)) + ((g157) & (sk[23]) & (g186) & (g192)));
	assign g506 = (((!g125) & (!g253) & (!g483) & (sk[24]) & (!g504) & (!g505)) + ((!g125) & (!g253) & (!g483) & (sk[24]) & (g504) & (!g505)) + ((!g125) & (!g253) & (g483) & (!sk[24]) & (!g504) & (g505)) + ((!g125) & (!g253) & (g483) & (!sk[24]) & (g504) & (!g505)) + ((!g125) & (!g253) & (g483) & (!sk[24]) & (g504) & (g505)) + ((!g125) & (g253) & (!g483) & (!sk[24]) & (!g504) & (!g505)) + ((!g125) & (g253) & (!g483) & (!sk[24]) & (!g504) & (g505)) + ((!g125) & (g253) & (!g483) & (!sk[24]) & (g504) & (!g505)) + ((!g125) & (g253) & (!g483) & (!sk[24]) & (g504) & (g505)) + ((!g125) & (g253) & (!g483) & (sk[24]) & (!g504) & (!g505)) + ((!g125) & (g253) & (!g483) & (sk[24]) & (g504) & (!g505)) + ((!g125) & (g253) & (g483) & (!sk[24]) & (!g504) & (!g505)) + ((!g125) & (g253) & (g483) & (!sk[24]) & (!g504) & (g505)) + ((!g125) & (g253) & (g483) & (!sk[24]) & (g504) & (!g505)) + ((!g125) & (g253) & (g483) & (!sk[24]) & (g504) & (g505)) + ((!g125) & (g253) & (g483) & (sk[24]) & (!g504) & (!g505)) + ((!g125) & (g253) & (g483) & (sk[24]) & (g504) & (!g505)) + ((g125) & (!g253) & (!g483) & (sk[24]) & (g504) & (!g505)) + ((g125) & (!g253) & (g483) & (!sk[24]) & (!g504) & (g505)) + ((g125) & (!g253) & (g483) & (!sk[24]) & (g504) & (!g505)) + ((g125) & (!g253) & (g483) & (!sk[24]) & (g504) & (g505)) + ((g125) & (g253) & (!g483) & (!sk[24]) & (!g504) & (!g505)) + ((g125) & (g253) & (!g483) & (!sk[24]) & (!g504) & (g505)) + ((g125) & (g253) & (!g483) & (!sk[24]) & (g504) & (!g505)) + ((g125) & (g253) & (!g483) & (!sk[24]) & (g504) & (g505)) + ((g125) & (g253) & (!g483) & (sk[24]) & (g504) & (!g505)) + ((g125) & (g253) & (g483) & (!sk[24]) & (!g504) & (!g505)) + ((g125) & (g253) & (g483) & (!sk[24]) & (!g504) & (g505)) + ((g125) & (g253) & (g483) & (!sk[24]) & (g504) & (!g505)) + ((g125) & (g253) & (g483) & (!sk[24]) & (g504) & (g505)) + ((g125) & (g253) & (g483) & (sk[24]) & (g504) & (!g505)));
	assign g507 = (((!i_12_) & (!i_13_) & (!sk[25]) & (i_14_)) + ((!i_12_) & (i_13_) & (!sk[25]) & (!i_14_)) + ((!i_12_) & (i_13_) & (!sk[25]) & (i_14_)) + ((!i_12_) & (i_13_) & (sk[25]) & (i_14_)) + ((i_12_) & (!i_13_) & (!sk[25]) & (i_14_)) + ((i_12_) & (!i_13_) & (sk[25]) & (i_14_)) + ((i_12_) & (i_13_) & (!sk[25]) & (!i_14_)) + ((i_12_) & (i_13_) & (!sk[25]) & (i_14_)));
	assign g508 = (((g69) & (!sk[26]) & (!g507)) + ((g69) & (!sk[26]) & (g507)) + ((g69) & (sk[26]) & (g507)));
	assign g509 = (((!g355) & (!g125) & (!sk[27]) & (g88) & (!g191)) + ((!g355) & (!g125) & (!sk[27]) & (g88) & (g191)) + ((!g355) & (g125) & (!sk[27]) & (g88) & (!g191)) + ((!g355) & (g125) & (!sk[27]) & (g88) & (g191)) + ((!g355) & (g125) & (sk[27]) & (!g88) & (g191)) + ((!g355) & (g125) & (sk[27]) & (g88) & (g191)) + ((g355) & (!g125) & (!sk[27]) & (g88) & (!g191)) + ((g355) & (!g125) & (!sk[27]) & (g88) & (g191)) + ((g355) & (g125) & (!sk[27]) & (g88) & (!g191)) + ((g355) & (g125) & (!sk[27]) & (g88) & (g191)) + ((g355) & (g125) & (sk[27]) & (!g88) & (g191)) + ((g355) & (g125) & (sk[27]) & (g88) & (!g191)) + ((g355) & (g125) & (sk[27]) & (g88) & (g191)));
	assign g510 = (((!g122) & (!g413) & (!g473) & (sk[28]) & (!g508) & (!g509)) + ((!g122) & (!g413) & (g473) & (!sk[28]) & (!g508) & (g509)) + ((!g122) & (!g413) & (g473) & (!sk[28]) & (g508) & (!g509)) + ((!g122) & (!g413) & (g473) & (!sk[28]) & (g508) & (g509)) + ((!g122) & (g413) & (!g473) & (!sk[28]) & (!g508) & (!g509)) + ((!g122) & (g413) & (!g473) & (!sk[28]) & (!g508) & (g509)) + ((!g122) & (g413) & (!g473) & (!sk[28]) & (g508) & (!g509)) + ((!g122) & (g413) & (!g473) & (!sk[28]) & (g508) & (g509)) + ((!g122) & (g413) & (!g473) & (sk[28]) & (!g508) & (!g509)) + ((!g122) & (g413) & (!g473) & (sk[28]) & (g508) & (!g509)) + ((!g122) & (g413) & (g473) & (!sk[28]) & (!g508) & (!g509)) + ((!g122) & (g413) & (g473) & (!sk[28]) & (!g508) & (g509)) + ((!g122) & (g413) & (g473) & (!sk[28]) & (g508) & (!g509)) + ((!g122) & (g413) & (g473) & (!sk[28]) & (g508) & (g509)) + ((!g122) & (g413) & (g473) & (sk[28]) & (!g508) & (!g509)) + ((!g122) & (g413) & (g473) & (sk[28]) & (g508) & (!g509)) + ((g122) & (!g413) & (!g473) & (sk[28]) & (!g508) & (!g509)) + ((g122) & (!g413) & (g473) & (!sk[28]) & (!g508) & (g509)) + ((g122) & (!g413) & (g473) & (!sk[28]) & (g508) & (!g509)) + ((g122) & (!g413) & (g473) & (!sk[28]) & (g508) & (g509)) + ((g122) & (g413) & (!g473) & (!sk[28]) & (!g508) & (!g509)) + ((g122) & (g413) & (!g473) & (!sk[28]) & (!g508) & (g509)) + ((g122) & (g413) & (!g473) & (!sk[28]) & (g508) & (!g509)) + ((g122) & (g413) & (!g473) & (!sk[28]) & (g508) & (g509)) + ((g122) & (g413) & (!g473) & (sk[28]) & (!g508) & (!g509)) + ((g122) & (g413) & (!g473) & (sk[28]) & (g508) & (!g509)) + ((g122) & (g413) & (g473) & (!sk[28]) & (!g508) & (!g509)) + ((g122) & (g413) & (g473) & (!sk[28]) & (!g508) & (g509)) + ((g122) & (g413) & (g473) & (!sk[28]) & (g508) & (!g509)) + ((g122) & (g413) & (g473) & (!sk[28]) & (g508) & (g509)));
	assign g511 = (((g69) & (!sk[29]) & (!g460)) + ((g69) & (!sk[29]) & (g460)) + ((g69) & (sk[29]) & (!g460)));
	assign g512 = (((!g180) & (!g225) & (!sk[30]) & (g213) & (!g425)) + ((!g180) & (!g225) & (!sk[30]) & (g213) & (g425)) + ((!g180) & (g225) & (!sk[30]) & (g213) & (!g425)) + ((!g180) & (g225) & (!sk[30]) & (g213) & (g425)) + ((g180) & (!g225) & (!sk[30]) & (g213) & (!g425)) + ((g180) & (!g225) & (!sk[30]) & (g213) & (g425)) + ((g180) & (!g225) & (sk[30]) & (!g213) & (!g425)) + ((g180) & (!g225) & (sk[30]) & (g213) & (!g425)) + ((g180) & (!g225) & (sk[30]) & (g213) & (g425)) + ((g180) & (g225) & (!sk[30]) & (g213) & (!g425)) + ((g180) & (g225) & (!sk[30]) & (g213) & (g425)) + ((g180) & (g225) & (sk[30]) & (!g213) & (!g425)) + ((g180) & (g225) & (sk[30]) & (!g213) & (g425)) + ((g180) & (g225) & (sk[30]) & (g213) & (!g425)) + ((g180) & (g225) & (sk[30]) & (g213) & (g425)));
	assign g513 = (((!g36) & (sk[31]) & (!g76)) + ((!g36) & (sk[31]) & (g76)) + ((g36) & (!sk[31]) & (!g76)) + ((g36) & (!sk[31]) & (g76)) + ((g36) & (sk[31]) & (g76)));
	assign g514 = (((!g24) & (sk[32]) & (g36)) + ((g24) & (!sk[32]) & (!g36)) + ((g24) & (!sk[32]) & (g36)));
	assign g515 = (((!g125) & (!g192) & (g513) & (!sk[33]) & (!g514)) + ((!g125) & (!g192) & (g513) & (!sk[33]) & (g514)) + ((!g125) & (g192) & (g513) & (!sk[33]) & (!g514)) + ((!g125) & (g192) & (g513) & (!sk[33]) & (g514)) + ((g125) & (!g192) & (!g513) & (sk[33]) & (!g514)) + ((g125) & (!g192) & (!g513) & (sk[33]) & (g514)) + ((g125) & (!g192) & (g513) & (!sk[33]) & (!g514)) + ((g125) & (!g192) & (g513) & (!sk[33]) & (g514)) + ((g125) & (!g192) & (g513) & (sk[33]) & (g514)) + ((g125) & (g192) & (!g513) & (sk[33]) & (!g514)) + ((g125) & (g192) & (!g513) & (sk[33]) & (g514)) + ((g125) & (g192) & (g513) & (!sk[33]) & (!g514)) + ((g125) & (g192) & (g513) & (!sk[33]) & (g514)) + ((g125) & (g192) & (g513) & (sk[33]) & (!g514)) + ((g125) & (g192) & (g513) & (sk[33]) & (g514)));
	assign g516 = (((!g188) & (!g436) & (!g511) & (sk[34]) & (!g512) & (!g515)) + ((!g188) & (!g436) & (g511) & (!sk[34]) & (!g512) & (g515)) + ((!g188) & (!g436) & (g511) & (!sk[34]) & (g512) & (!g515)) + ((!g188) & (!g436) & (g511) & (!sk[34]) & (g512) & (g515)) + ((!g188) & (!g436) & (g511) & (sk[34]) & (!g512) & (!g515)) + ((!g188) & (g436) & (!g511) & (!sk[34]) & (!g512) & (!g515)) + ((!g188) & (g436) & (!g511) & (!sk[34]) & (!g512) & (g515)) + ((!g188) & (g436) & (!g511) & (!sk[34]) & (g512) & (!g515)) + ((!g188) & (g436) & (!g511) & (!sk[34]) & (g512) & (g515)) + ((!g188) & (g436) & (!g511) & (sk[34]) & (!g512) & (!g515)) + ((!g188) & (g436) & (g511) & (!sk[34]) & (!g512) & (!g515)) + ((!g188) & (g436) & (g511) & (!sk[34]) & (!g512) & (g515)) + ((!g188) & (g436) & (g511) & (!sk[34]) & (g512) & (!g515)) + ((!g188) & (g436) & (g511) & (!sk[34]) & (g512) & (g515)) + ((g188) & (!g436) & (!g511) & (sk[34]) & (!g512) & (!g515)) + ((g188) & (!g436) & (g511) & (!sk[34]) & (!g512) & (g515)) + ((g188) & (!g436) & (g511) & (!sk[34]) & (g512) & (!g515)) + ((g188) & (!g436) & (g511) & (!sk[34]) & (g512) & (g515)) + ((g188) & (!g436) & (g511) & (sk[34]) & (!g512) & (!g515)) + ((g188) & (g436) & (!g511) & (!sk[34]) & (!g512) & (!g515)) + ((g188) & (g436) & (!g511) & (!sk[34]) & (!g512) & (g515)) + ((g188) & (g436) & (!g511) & (!sk[34]) & (g512) & (!g515)) + ((g188) & (g436) & (!g511) & (!sk[34]) & (g512) & (g515)) + ((g188) & (g436) & (g511) & (!sk[34]) & (!g512) & (!g515)) + ((g188) & (g436) & (g511) & (!sk[34]) & (!g512) & (g515)) + ((g188) & (g436) & (g511) & (!sk[34]) & (g512) & (!g515)) + ((g188) & (g436) & (g511) & (!sk[34]) & (g512) & (g515)));
	assign g517 = (((!g24) & (!g113) & (!g257) & (sk[35]) & (g356)) + ((!g24) & (!g113) & (g257) & (!sk[35]) & (!g356)) + ((!g24) & (!g113) & (g257) & (!sk[35]) & (g356)) + ((!g24) & (!g113) & (g257) & (sk[35]) & (!g356)) + ((!g24) & (!g113) & (g257) & (sk[35]) & (g356)) + ((!g24) & (g113) & (g257) & (!sk[35]) & (!g356)) + ((!g24) & (g113) & (g257) & (!sk[35]) & (g356)) + ((g24) & (!g113) & (g257) & (!sk[35]) & (!g356)) + ((g24) & (!g113) & (g257) & (!sk[35]) & (g356)) + ((g24) & (g113) & (g257) & (!sk[35]) & (!g356)) + ((g24) & (g113) & (g257) & (!sk[35]) & (g356)));
	assign g518 = (((!i_8_) & (!sk[36]) & (!i_6_) & (i_7_) & (!g120)) + ((!i_8_) & (!sk[36]) & (!i_6_) & (i_7_) & (g120)) + ((!i_8_) & (!sk[36]) & (i_6_) & (i_7_) & (!g120)) + ((!i_8_) & (!sk[36]) & (i_6_) & (i_7_) & (g120)) + ((!i_8_) & (sk[36]) & (!i_6_) & (!i_7_) & (g120)) + ((i_8_) & (!sk[36]) & (!i_6_) & (i_7_) & (!g120)) + ((i_8_) & (!sk[36]) & (!i_6_) & (i_7_) & (g120)) + ((i_8_) & (!sk[36]) & (i_6_) & (i_7_) & (!g120)) + ((i_8_) & (!sk[36]) & (i_6_) & (i_7_) & (g120)) + ((i_8_) & (sk[36]) & (!i_6_) & (!i_7_) & (g120)) + ((i_8_) & (sk[36]) & (!i_6_) & (i_7_) & (g120)));
	assign g519 = (((!g348) & (!sk[37]) & (!g514) & (g517) & (!g1577)) + ((!g348) & (!sk[37]) & (!g514) & (g517) & (g1577)) + ((!g348) & (!sk[37]) & (g514) & (g517) & (!g1577)) + ((!g348) & (!sk[37]) & (g514) & (g517) & (g1577)) + ((!g348) & (sk[37]) & (!g514) & (!g517) & (g1577)) + ((g348) & (!sk[37]) & (!g514) & (g517) & (!g1577)) + ((g348) & (!sk[37]) & (!g514) & (g517) & (g1577)) + ((g348) & (!sk[37]) & (g514) & (g517) & (!g1577)) + ((g348) & (!sk[37]) & (g514) & (g517) & (g1577)) + ((g348) & (sk[37]) & (!g514) & (!g517) & (g1577)) + ((g348) & (sk[37]) & (g514) & (!g517) & (g1577)));
	assign g520 = (((!i_9_) & (!i_10_) & (!i_11_) & (sk[38]) & (!g225) & (!g213)) + ((!i_9_) & (!i_10_) & (!i_11_) & (sk[38]) & (!g225) & (g213)) + ((!i_9_) & (!i_10_) & (!i_11_) & (sk[38]) & (g225) & (!g213)) + ((!i_9_) & (!i_10_) & (!i_11_) & (sk[38]) & (g225) & (g213)) + ((!i_9_) & (!i_10_) & (i_11_) & (!sk[38]) & (!g225) & (g213)) + ((!i_9_) & (!i_10_) & (i_11_) & (!sk[38]) & (g225) & (!g213)) + ((!i_9_) & (!i_10_) & (i_11_) & (!sk[38]) & (g225) & (g213)) + ((!i_9_) & (!i_10_) & (i_11_) & (sk[38]) & (!g225) & (!g213)) + ((!i_9_) & (!i_10_) & (i_11_) & (sk[38]) & (!g225) & (g213)) + ((!i_9_) & (!i_10_) & (i_11_) & (sk[38]) & (g225) & (!g213)) + ((!i_9_) & (!i_10_) & (i_11_) & (sk[38]) & (g225) & (g213)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[38]) & (!g225) & (!g213)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[38]) & (!g225) & (g213)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[38]) & (g225) & (!g213)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[38]) & (g225) & (g213)) + ((!i_9_) & (i_10_) & (!i_11_) & (sk[38]) & (!g225) & (!g213)) + ((!i_9_) & (i_10_) & (!i_11_) & (sk[38]) & (!g225) & (g213)) + ((!i_9_) & (i_10_) & (!i_11_) & (sk[38]) & (g225) & (!g213)) + ((!i_9_) & (i_10_) & (!i_11_) & (sk[38]) & (g225) & (g213)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[38]) & (!g225) & (!g213)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[38]) & (!g225) & (g213)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[38]) & (g225) & (!g213)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[38]) & (g225) & (g213)) + ((!i_9_) & (i_10_) & (i_11_) & (sk[38]) & (!g225) & (!g213)) + ((!i_9_) & (i_10_) & (i_11_) & (sk[38]) & (!g225) & (g213)) + ((!i_9_) & (i_10_) & (i_11_) & (sk[38]) & (g225) & (!g213)) + ((!i_9_) & (i_10_) & (i_11_) & (sk[38]) & (g225) & (g213)) + ((i_9_) & (!i_10_) & (!i_11_) & (sk[38]) & (!g225) & (!g213)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[38]) & (!g225) & (g213)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[38]) & (g225) & (!g213)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[38]) & (g225) & (g213)) + ((i_9_) & (!i_10_) & (i_11_) & (sk[38]) & (!g225) & (!g213)) + ((i_9_) & (!i_10_) & (i_11_) & (sk[38]) & (!g225) & (g213)) + ((i_9_) & (!i_10_) & (i_11_) & (sk[38]) & (g225) & (!g213)) + ((i_9_) & (!i_10_) & (i_11_) & (sk[38]) & (g225) & (g213)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[38]) & (!g225) & (!g213)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[38]) & (!g225) & (g213)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[38]) & (g225) & (!g213)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[38]) & (g225) & (g213)) + ((i_9_) & (i_10_) & (!i_11_) & (sk[38]) & (!g225) & (!g213)) + ((i_9_) & (i_10_) & (!i_11_) & (sk[38]) & (!g225) & (g213)) + ((i_9_) & (i_10_) & (!i_11_) & (sk[38]) & (g225) & (!g213)) + ((i_9_) & (i_10_) & (!i_11_) & (sk[38]) & (g225) & (g213)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[38]) & (!g225) & (!g213)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[38]) & (!g225) & (g213)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[38]) & (g225) & (!g213)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[38]) & (g225) & (g213)) + ((i_9_) & (i_10_) & (i_11_) & (sk[38]) & (!g225) & (!g213)) + ((i_9_) & (i_10_) & (i_11_) & (sk[38]) & (!g225) & (g213)) + ((i_9_) & (i_10_) & (i_11_) & (sk[38]) & (g225) & (!g213)) + ((i_9_) & (i_10_) & (i_11_) & (sk[38]) & (g225) & (g213)));
	assign g521 = (((!sk[39]) & (g22) & (!g482)) + ((!sk[39]) & (g22) & (g482)) + ((sk[39]) & (!g22) & (g482)));
	assign g522 = (((g88) & (!sk[40]) & (!g174)) + ((g88) & (!sk[40]) & (g174)) + ((g88) & (sk[40]) & (!g174)));
	assign g523 = (((!g164) & (!sk[41]) & (!g253) & (g483) & (!g484) & (g500)) + ((!g164) & (!sk[41]) & (!g253) & (g483) & (g484) & (!g500)) + ((!g164) & (!sk[41]) & (!g253) & (g483) & (g484) & (g500)) + ((!g164) & (!sk[41]) & (g253) & (!g483) & (!g484) & (!g500)) + ((!g164) & (!sk[41]) & (g253) & (!g483) & (!g484) & (g500)) + ((!g164) & (!sk[41]) & (g253) & (!g483) & (g484) & (!g500)) + ((!g164) & (!sk[41]) & (g253) & (!g483) & (g484) & (g500)) + ((!g164) & (!sk[41]) & (g253) & (g483) & (!g484) & (!g500)) + ((!g164) & (!sk[41]) & (g253) & (g483) & (!g484) & (g500)) + ((!g164) & (!sk[41]) & (g253) & (g483) & (g484) & (!g500)) + ((!g164) & (!sk[41]) & (g253) & (g483) & (g484) & (g500)) + ((!g164) & (sk[41]) & (!g253) & (!g483) & (!g484) & (!g500)) + ((!g164) & (sk[41]) & (!g253) & (!g483) & (g484) & (!g500)) + ((!g164) & (sk[41]) & (!g253) & (g483) & (!g484) & (!g500)) + ((!g164) & (sk[41]) & (!g253) & (g483) & (g484) & (!g500)) + ((!g164) & (sk[41]) & (g253) & (!g483) & (!g484) & (!g500)) + ((!g164) & (sk[41]) & (g253) & (!g483) & (!g484) & (g500)) + ((!g164) & (sk[41]) & (g253) & (!g483) & (g484) & (!g500)) + ((!g164) & (sk[41]) & (g253) & (!g483) & (g484) & (g500)) + ((!g164) & (sk[41]) & (g253) & (g483) & (!g484) & (!g500)) + ((!g164) & (sk[41]) & (g253) & (g483) & (!g484) & (g500)) + ((!g164) & (sk[41]) & (g253) & (g483) & (g484) & (!g500)) + ((!g164) & (sk[41]) & (g253) & (g483) & (g484) & (g500)) + ((g164) & (!sk[41]) & (!g253) & (g483) & (!g484) & (g500)) + ((g164) & (!sk[41]) & (!g253) & (g483) & (g484) & (!g500)) + ((g164) & (!sk[41]) & (!g253) & (g483) & (g484) & (g500)) + ((g164) & (!sk[41]) & (g253) & (!g483) & (!g484) & (!g500)) + ((g164) & (!sk[41]) & (g253) & (!g483) & (!g484) & (g500)) + ((g164) & (!sk[41]) & (g253) & (!g483) & (g484) & (!g500)) + ((g164) & (!sk[41]) & (g253) & (!g483) & (g484) & (g500)) + ((g164) & (!sk[41]) & (g253) & (g483) & (!g484) & (!g500)) + ((g164) & (!sk[41]) & (g253) & (g483) & (!g484) & (g500)) + ((g164) & (!sk[41]) & (g253) & (g483) & (g484) & (!g500)) + ((g164) & (!sk[41]) & (g253) & (g483) & (g484) & (g500)) + ((g164) & (sk[41]) & (!g253) & (!g483) & (!g484) & (!g500)) + ((g164) & (sk[41]) & (g253) & (!g483) & (!g484) & (!g500)) + ((g164) & (sk[41]) & (g253) & (!g483) & (!g484) & (g500)));
	assign g524 = (((!sk[42]) & (!g164) & (!g521) & (g522) & (!g523)) + ((!sk[42]) & (!g164) & (!g521) & (g522) & (g523)) + ((!sk[42]) & (!g164) & (g521) & (g522) & (!g523)) + ((!sk[42]) & (!g164) & (g521) & (g522) & (g523)) + ((!sk[42]) & (g164) & (!g521) & (g522) & (!g523)) + ((!sk[42]) & (g164) & (!g521) & (g522) & (g523)) + ((!sk[42]) & (g164) & (g521) & (g522) & (!g523)) + ((!sk[42]) & (g164) & (g521) & (g522) & (g523)) + ((sk[42]) & (!g164) & (!g521) & (!g522) & (g523)) + ((sk[42]) & (!g164) & (!g521) & (g522) & (g523)) + ((sk[42]) & (!g164) & (g521) & (!g522) & (g523)) + ((sk[42]) & (!g164) & (g521) & (g522) & (g523)) + ((sk[42]) & (g164) & (!g521) & (!g522) & (g523)));
	assign g525 = (((g503) & (g506) & (g510) & (g516) & (g519) & (g1564)));
	assign g526 = (((!g22) & (!g24) & (!g125) & (!g123) & (sk[44]) & (!g438)) + ((!g22) & (!g24) & (!g125) & (!g123) & (sk[44]) & (g438)) + ((!g22) & (!g24) & (!g125) & (g123) & (sk[44]) & (!g438)) + ((!g22) & (!g24) & (g125) & (!g123) & (!sk[44]) & (g438)) + ((!g22) & (!g24) & (g125) & (!g123) & (sk[44]) & (!g438)) + ((!g22) & (!g24) & (g125) & (!g123) & (sk[44]) & (g438)) + ((!g22) & (!g24) & (g125) & (g123) & (!sk[44]) & (!g438)) + ((!g22) & (!g24) & (g125) & (g123) & (!sk[44]) & (g438)) + ((!g22) & (!g24) & (g125) & (g123) & (sk[44]) & (!g438)) + ((!g22) & (!g24) & (g125) & (g123) & (sk[44]) & (g438)) + ((!g22) & (g24) & (!g125) & (!g123) & (!sk[44]) & (!g438)) + ((!g22) & (g24) & (!g125) & (!g123) & (!sk[44]) & (g438)) + ((!g22) & (g24) & (!g125) & (g123) & (!sk[44]) & (!g438)) + ((!g22) & (g24) & (!g125) & (g123) & (!sk[44]) & (g438)) + ((!g22) & (g24) & (g125) & (!g123) & (!sk[44]) & (!g438)) + ((!g22) & (g24) & (g125) & (!g123) & (!sk[44]) & (g438)) + ((!g22) & (g24) & (g125) & (g123) & (!sk[44]) & (!g438)) + ((!g22) & (g24) & (g125) & (g123) & (!sk[44]) & (g438)) + ((g22) & (!g24) & (g125) & (!g123) & (!sk[44]) & (g438)) + ((g22) & (!g24) & (g125) & (g123) & (!sk[44]) & (!g438)) + ((g22) & (!g24) & (g125) & (g123) & (!sk[44]) & (g438)) + ((g22) & (g24) & (!g125) & (!g123) & (!sk[44]) & (!g438)) + ((g22) & (g24) & (!g125) & (!g123) & (!sk[44]) & (g438)) + ((g22) & (g24) & (!g125) & (g123) & (!sk[44]) & (!g438)) + ((g22) & (g24) & (!g125) & (g123) & (!sk[44]) & (g438)) + ((g22) & (g24) & (g125) & (!g123) & (!sk[44]) & (!g438)) + ((g22) & (g24) & (g125) & (!g123) & (!sk[44]) & (g438)) + ((g22) & (g24) & (g125) & (g123) & (!sk[44]) & (!g438)) + ((g22) & (g24) & (g125) & (g123) & (!sk[44]) & (g438)));
	assign g527 = (((!sk[45]) & (!g355) & (!g75) & (g91) & (!g212)) + ((!sk[45]) & (!g355) & (!g75) & (g91) & (g212)) + ((!sk[45]) & (!g355) & (g75) & (g91) & (!g212)) + ((!sk[45]) & (!g355) & (g75) & (g91) & (g212)) + ((!sk[45]) & (g355) & (!g75) & (g91) & (!g212)) + ((!sk[45]) & (g355) & (!g75) & (g91) & (g212)) + ((!sk[45]) & (g355) & (g75) & (g91) & (!g212)) + ((!sk[45]) & (g355) & (g75) & (g91) & (g212)) + ((sk[45]) & (!g355) & (!g75) & (!g91) & (g212)) + ((sk[45]) & (!g355) & (!g75) & (g91) & (g212)) + ((sk[45]) & (g355) & (!g75) & (!g91) & (!g212)) + ((sk[45]) & (g355) & (!g75) & (!g91) & (g212)) + ((sk[45]) & (g355) & (!g75) & (g91) & (g212)));
	assign g528 = (((!g17) & (!sk[46]) & (!g22) & (g24) & (!g81)) + ((!g17) & (!sk[46]) & (!g22) & (g24) & (g81)) + ((!g17) & (!sk[46]) & (g22) & (g24) & (!g81)) + ((!g17) & (!sk[46]) & (g22) & (g24) & (g81)) + ((!g17) & (sk[46]) & (!g22) & (!g24) & (!g81)) + ((!g17) & (sk[46]) & (!g22) & (!g24) & (g81)) + ((!g17) & (sk[46]) & (g22) & (!g24) & (g81)) + ((g17) & (!sk[46]) & (!g22) & (g24) & (!g81)) + ((g17) & (!sk[46]) & (!g22) & (g24) & (g81)) + ((g17) & (!sk[46]) & (g22) & (g24) & (!g81)) + ((g17) & (!sk[46]) & (g22) & (g24) & (g81)) + ((g17) & (sk[46]) & (!g22) & (!g24) & (!g81)) + ((g17) & (sk[46]) & (!g22) & (!g24) & (g81)) + ((g17) & (sk[46]) & (g22) & (!g24) & (!g81)) + ((g17) & (sk[46]) & (g22) & (!g24) & (g81)));
	assign g529 = (((!g73) & (!g468) & (!sk[47]) & (g487) & (!g528)) + ((!g73) & (!g468) & (!sk[47]) & (g487) & (g528)) + ((!g73) & (g468) & (!sk[47]) & (g487) & (!g528)) + ((!g73) & (g468) & (!sk[47]) & (g487) & (g528)) + ((g73) & (!g468) & (!sk[47]) & (g487) & (!g528)) + ((g73) & (!g468) & (!sk[47]) & (g487) & (g528)) + ((g73) & (!g468) & (sk[47]) & (!g487) & (g528)) + ((g73) & (!g468) & (sk[47]) & (g487) & (!g528)) + ((g73) & (!g468) & (sk[47]) & (g487) & (g528)) + ((g73) & (g468) & (!sk[47]) & (g487) & (!g528)) + ((g73) & (g468) & (!sk[47]) & (g487) & (g528)) + ((g73) & (g468) & (sk[47]) & (!g487) & (!g528)) + ((g73) & (g468) & (sk[47]) & (!g487) & (g528)) + ((g73) & (g468) & (sk[47]) & (g487) & (!g528)) + ((g73) & (g468) & (sk[47]) & (g487) & (g528)));
	assign g530 = (((!g75) & (!g192) & (g513) & (!g514) & (!g527) & (!g529)) + ((g75) & (!g192) & (!g513) & (!g514) & (!g527) & (!g529)) + ((g75) & (!g192) & (!g513) & (g514) & (!g527) & (!g529)) + ((g75) & (!g192) & (g513) & (!g514) & (!g527) & (!g529)) + ((g75) & (!g192) & (g513) & (g514) & (!g527) & (!g529)) + ((g75) & (g192) & (!g513) & (!g514) & (!g527) & (!g529)) + ((g75) & (g192) & (!g513) & (g514) & (!g527) & (!g529)) + ((g75) & (g192) & (g513) & (!g514) & (!g527) & (!g529)) + ((g75) & (g192) & (g513) & (g514) & (!g527) & (!g529)));
	assign g531 = (((!g69) & (!sk[49]) & (!g154) & (g113) & (!g119) & (g482)) + ((!g69) & (!sk[49]) & (!g154) & (g113) & (g119) & (!g482)) + ((!g69) & (!sk[49]) & (!g154) & (g113) & (g119) & (g482)) + ((!g69) & (!sk[49]) & (g154) & (!g113) & (!g119) & (!g482)) + ((!g69) & (!sk[49]) & (g154) & (!g113) & (!g119) & (g482)) + ((!g69) & (!sk[49]) & (g154) & (!g113) & (g119) & (!g482)) + ((!g69) & (!sk[49]) & (g154) & (!g113) & (g119) & (g482)) + ((!g69) & (!sk[49]) & (g154) & (g113) & (!g119) & (!g482)) + ((!g69) & (!sk[49]) & (g154) & (g113) & (!g119) & (g482)) + ((!g69) & (!sk[49]) & (g154) & (g113) & (g119) & (!g482)) + ((!g69) & (!sk[49]) & (g154) & (g113) & (g119) & (g482)) + ((!g69) & (sk[49]) & (!g154) & (!g113) & (!g119) & (g482)) + ((!g69) & (sk[49]) & (!g154) & (!g113) & (g119) & (g482)) + ((g69) & (!sk[49]) & (!g154) & (g113) & (!g119) & (g482)) + ((g69) & (!sk[49]) & (!g154) & (g113) & (g119) & (!g482)) + ((g69) & (!sk[49]) & (!g154) & (g113) & (g119) & (g482)) + ((g69) & (!sk[49]) & (g154) & (!g113) & (!g119) & (!g482)) + ((g69) & (!sk[49]) & (g154) & (!g113) & (!g119) & (g482)) + ((g69) & (!sk[49]) & (g154) & (!g113) & (g119) & (!g482)) + ((g69) & (!sk[49]) & (g154) & (!g113) & (g119) & (g482)) + ((g69) & (!sk[49]) & (g154) & (g113) & (!g119) & (!g482)) + ((g69) & (!sk[49]) & (g154) & (g113) & (!g119) & (g482)) + ((g69) & (!sk[49]) & (g154) & (g113) & (g119) & (!g482)) + ((g69) & (!sk[49]) & (g154) & (g113) & (g119) & (g482)) + ((g69) & (sk[49]) & (!g154) & (!g113) & (!g119) & (g482)) + ((g69) & (sk[49]) & (!g154) & (!g113) & (g119) & (g482)) + ((g69) & (sk[49]) & (!g154) & (g113) & (g119) & (g482)) + ((g69) & (sk[49]) & (g154) & (!g113) & (g119) & (g482)) + ((g69) & (sk[49]) & (g154) & (g113) & (g119) & (g482)));
	assign g532 = (((!g24) & (!g122) & (!g113) & (!g105) & (g174) & (!g531)) + ((!g24) & (!g122) & (!g113) & (g105) & (!g174) & (!g531)) + ((!g24) & (!g122) & (!g113) & (g105) & (g174) & (!g531)) + ((!g24) & (!g122) & (g113) & (!g105) & (!g174) & (!g531)) + ((!g24) & (!g122) & (g113) & (!g105) & (g174) & (!g531)) + ((!g24) & (!g122) & (g113) & (g105) & (!g174) & (!g531)) + ((!g24) & (!g122) & (g113) & (g105) & (g174) & (!g531)) + ((!g24) & (g122) & (g113) & (!g105) & (!g174) & (!g531)) + ((!g24) & (g122) & (g113) & (!g105) & (g174) & (!g531)) + ((!g24) & (g122) & (g113) & (g105) & (!g174) & (!g531)) + ((!g24) & (g122) & (g113) & (g105) & (g174) & (!g531)) + ((g24) & (!g122) & (!g113) & (!g105) & (g174) & (!g531)) + ((g24) & (!g122) & (!g113) & (g105) & (!g174) & (!g531)) + ((g24) & (!g122) & (!g113) & (g105) & (g174) & (!g531)) + ((g24) & (!g122) & (g113) & (!g105) & (!g174) & (!g531)) + ((g24) & (!g122) & (g113) & (!g105) & (g174) & (!g531)) + ((g24) & (!g122) & (g113) & (g105) & (!g174) & (!g531)) + ((g24) & (!g122) & (g113) & (g105) & (g174) & (!g531)) + ((g24) & (g122) & (!g113) & (!g105) & (g174) & (!g531)) + ((g24) & (g122) & (!g113) & (g105) & (!g174) & (!g531)) + ((g24) & (g122) & (!g113) & (g105) & (g174) & (!g531)) + ((g24) & (g122) & (g113) & (!g105) & (!g174) & (!g531)) + ((g24) & (g122) & (g113) & (!g105) & (g174) & (!g531)) + ((g24) & (g122) & (g113) & (g105) & (!g174) & (!g531)) + ((g24) & (g122) & (g113) & (g105) & (g174) & (!g531)));
	assign g533 = (((!i_9_) & (!i_10_) & (!i_11_) & (!i_15_) & (!g174) & (!g460)) + ((!i_9_) & (!i_10_) & (!i_11_) & (!i_15_) & (g174) & (!g460)) + ((!i_9_) & (!i_10_) & (i_11_) & (!i_15_) & (!g174) & (!g460)) + ((!i_9_) & (!i_10_) & (i_11_) & (!i_15_) & (g174) & (!g460)) + ((!i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (!g174) & (!g460)) + ((!i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (g174) & (!g460)) + ((!i_9_) & (i_10_) & (i_11_) & (!i_15_) & (!g174) & (!g460)) + ((!i_9_) & (i_10_) & (i_11_) & (!i_15_) & (g174) & (!g460)) + ((i_9_) & (!i_10_) & (!i_11_) & (!i_15_) & (!g174) & (!g460)) + ((i_9_) & (!i_10_) & (!i_11_) & (!i_15_) & (g174) & (!g460)) + ((i_9_) & (!i_10_) & (i_11_) & (!i_15_) & (!g174) & (!g460)) + ((i_9_) & (!i_10_) & (i_11_) & (!i_15_) & (g174) & (!g460)) + ((i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (!g174) & (!g460)) + ((i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (g174) & (!g460)) + ((i_9_) & (i_10_) & (!i_11_) & (i_15_) & (!g174) & (!g460)) + ((i_9_) & (i_10_) & (!i_11_) & (i_15_) & (!g174) & (g460)) + ((i_9_) & (i_10_) & (i_11_) & (!i_15_) & (!g174) & (!g460)) + ((i_9_) & (i_10_) & (i_11_) & (!i_15_) & (g174) & (!g460)));
	assign g534 = (((g88) & (!sk[52]) & (!g460)) + ((g88) & (!sk[52]) & (g460)) + ((g88) & (sk[52]) & (!g460)));
	assign g535 = (((!g157) & (!g191) & (g534) & (!g496) & (!sk[53]) & (g522)) + ((!g157) & (!g191) & (g534) & (g496) & (!sk[53]) & (!g522)) + ((!g157) & (!g191) & (g534) & (g496) & (!sk[53]) & (g522)) + ((!g157) & (g191) & (!g534) & (!g496) & (!sk[53]) & (!g522)) + ((!g157) & (g191) & (!g534) & (!g496) & (!sk[53]) & (g522)) + ((!g157) & (g191) & (!g534) & (g496) & (!sk[53]) & (!g522)) + ((!g157) & (g191) & (!g534) & (g496) & (!sk[53]) & (g522)) + ((!g157) & (g191) & (g534) & (!g496) & (!sk[53]) & (!g522)) + ((!g157) & (g191) & (g534) & (!g496) & (!sk[53]) & (g522)) + ((!g157) & (g191) & (g534) & (g496) & (!sk[53]) & (!g522)) + ((!g157) & (g191) & (g534) & (g496) & (!sk[53]) & (g522)) + ((g157) & (!g191) & (!g534) & (!g496) & (sk[53]) & (g522)) + ((g157) & (!g191) & (!g534) & (g496) & (sk[53]) & (!g522)) + ((g157) & (!g191) & (!g534) & (g496) & (sk[53]) & (g522)) + ((g157) & (!g191) & (g534) & (!g496) & (!sk[53]) & (g522)) + ((g157) & (!g191) & (g534) & (!g496) & (sk[53]) & (!g522)) + ((g157) & (!g191) & (g534) & (!g496) & (sk[53]) & (g522)) + ((g157) & (!g191) & (g534) & (g496) & (!sk[53]) & (!g522)) + ((g157) & (!g191) & (g534) & (g496) & (!sk[53]) & (g522)) + ((g157) & (!g191) & (g534) & (g496) & (sk[53]) & (!g522)) + ((g157) & (!g191) & (g534) & (g496) & (sk[53]) & (g522)) + ((g157) & (g191) & (!g534) & (!g496) & (!sk[53]) & (!g522)) + ((g157) & (g191) & (!g534) & (!g496) & (!sk[53]) & (g522)) + ((g157) & (g191) & (!g534) & (!g496) & (sk[53]) & (!g522)) + ((g157) & (g191) & (!g534) & (!g496) & (sk[53]) & (g522)) + ((g157) & (g191) & (!g534) & (g496) & (!sk[53]) & (!g522)) + ((g157) & (g191) & (!g534) & (g496) & (!sk[53]) & (g522)) + ((g157) & (g191) & (!g534) & (g496) & (sk[53]) & (!g522)) + ((g157) & (g191) & (!g534) & (g496) & (sk[53]) & (g522)) + ((g157) & (g191) & (g534) & (!g496) & (!sk[53]) & (!g522)) + ((g157) & (g191) & (g534) & (!g496) & (!sk[53]) & (g522)) + ((g157) & (g191) & (g534) & (!g496) & (sk[53]) & (!g522)) + ((g157) & (g191) & (g534) & (!g496) & (sk[53]) & (g522)) + ((g157) & (g191) & (g534) & (g496) & (!sk[53]) & (!g522)) + ((g157) & (g191) & (g534) & (g496) & (!sk[53]) & (g522)) + ((g157) & (g191) & (g534) & (g496) & (sk[53]) & (!g522)) + ((g157) & (g191) & (g534) & (g496) & (sk[53]) & (g522)));
	assign g536 = (((!sk[54]) & (!g168) & (!g435) & (g501) & (!g533) & (g535)) + ((!sk[54]) & (!g168) & (!g435) & (g501) & (g533) & (!g535)) + ((!sk[54]) & (!g168) & (!g435) & (g501) & (g533) & (g535)) + ((!sk[54]) & (!g168) & (g435) & (!g501) & (!g533) & (!g535)) + ((!sk[54]) & (!g168) & (g435) & (!g501) & (!g533) & (g535)) + ((!sk[54]) & (!g168) & (g435) & (!g501) & (g533) & (!g535)) + ((!sk[54]) & (!g168) & (g435) & (!g501) & (g533) & (g535)) + ((!sk[54]) & (!g168) & (g435) & (g501) & (!g533) & (!g535)) + ((!sk[54]) & (!g168) & (g435) & (g501) & (!g533) & (g535)) + ((!sk[54]) & (!g168) & (g435) & (g501) & (g533) & (!g535)) + ((!sk[54]) & (!g168) & (g435) & (g501) & (g533) & (g535)) + ((!sk[54]) & (g168) & (!g435) & (g501) & (!g533) & (g535)) + ((!sk[54]) & (g168) & (!g435) & (g501) & (g533) & (!g535)) + ((!sk[54]) & (g168) & (!g435) & (g501) & (g533) & (g535)) + ((!sk[54]) & (g168) & (g435) & (!g501) & (!g533) & (!g535)) + ((!sk[54]) & (g168) & (g435) & (!g501) & (!g533) & (g535)) + ((!sk[54]) & (g168) & (g435) & (!g501) & (g533) & (!g535)) + ((!sk[54]) & (g168) & (g435) & (!g501) & (g533) & (g535)) + ((!sk[54]) & (g168) & (g435) & (g501) & (!g533) & (!g535)) + ((!sk[54]) & (g168) & (g435) & (g501) & (!g533) & (g535)) + ((!sk[54]) & (g168) & (g435) & (g501) & (g533) & (!g535)) + ((!sk[54]) & (g168) & (g435) & (g501) & (g533) & (g535)) + ((sk[54]) & (!g168) & (!g435) & (!g501) & (!g533) & (!g535)) + ((sk[54]) & (!g168) & (!g435) & (!g501) & (g533) & (!g535)) + ((sk[54]) & (!g168) & (g435) & (!g501) & (!g533) & (!g535)) + ((sk[54]) & (!g168) & (g435) & (!g501) & (g533) & (!g535)) + ((sk[54]) & (!g168) & (g435) & (g501) & (!g533) & (!g535)) + ((sk[54]) & (!g168) & (g435) & (g501) & (g533) & (!g535)) + ((sk[54]) & (g168) & (!g435) & (!g501) & (!g533) & (!g535)) + ((sk[54]) & (g168) & (g435) & (!g501) & (!g533) & (!g535)) + ((sk[54]) & (g168) & (g435) & (g501) & (!g533) & (!g535)));
	assign g537 = (((!sk[55]) & (!g526) & (!g1459) & (g530) & (!g532) & (g536)) + ((!sk[55]) & (!g526) & (!g1459) & (g530) & (g532) & (!g536)) + ((!sk[55]) & (!g526) & (!g1459) & (g530) & (g532) & (g536)) + ((!sk[55]) & (!g526) & (g1459) & (!g530) & (!g532) & (!g536)) + ((!sk[55]) & (!g526) & (g1459) & (!g530) & (!g532) & (g536)) + ((!sk[55]) & (!g526) & (g1459) & (!g530) & (g532) & (!g536)) + ((!sk[55]) & (!g526) & (g1459) & (!g530) & (g532) & (g536)) + ((!sk[55]) & (!g526) & (g1459) & (g530) & (!g532) & (!g536)) + ((!sk[55]) & (!g526) & (g1459) & (g530) & (!g532) & (g536)) + ((!sk[55]) & (!g526) & (g1459) & (g530) & (g532) & (!g536)) + ((!sk[55]) & (!g526) & (g1459) & (g530) & (g532) & (g536)) + ((!sk[55]) & (g526) & (!g1459) & (g530) & (!g532) & (g536)) + ((!sk[55]) & (g526) & (!g1459) & (g530) & (g532) & (!g536)) + ((!sk[55]) & (g526) & (!g1459) & (g530) & (g532) & (g536)) + ((!sk[55]) & (g526) & (g1459) & (!g530) & (!g532) & (!g536)) + ((!sk[55]) & (g526) & (g1459) & (!g530) & (!g532) & (g536)) + ((!sk[55]) & (g526) & (g1459) & (!g530) & (g532) & (!g536)) + ((!sk[55]) & (g526) & (g1459) & (!g530) & (g532) & (g536)) + ((!sk[55]) & (g526) & (g1459) & (g530) & (!g532) & (!g536)) + ((!sk[55]) & (g526) & (g1459) & (g530) & (!g532) & (g536)) + ((!sk[55]) & (g526) & (g1459) & (g530) & (g532) & (!g536)) + ((!sk[55]) & (g526) & (g1459) & (g530) & (g532) & (g536)) + ((sk[55]) & (!g526) & (!g1459) & (g530) & (g532) & (g536)));
	assign g538 = (((!i_14_) & (!sk[56]) & (!g102) & (g113)) + ((!i_14_) & (!sk[56]) & (g102) & (!g113)) + ((!i_14_) & (!sk[56]) & (g102) & (g113)) + ((i_14_) & (!sk[56]) & (!g102) & (g113)) + ((i_14_) & (!sk[56]) & (g102) & (!g113)) + ((i_14_) & (!sk[56]) & (g102) & (g113)) + ((i_14_) & (sk[56]) & (g102) & (!g113)));
	assign g539 = (((!g119) & (!sk[57]) & (!g121) & (g213) & (!g351)) + ((!g119) & (!sk[57]) & (!g121) & (g213) & (g351)) + ((!g119) & (!sk[57]) & (g121) & (g213) & (!g351)) + ((!g119) & (!sk[57]) & (g121) & (g213) & (g351)) + ((!g119) & (sk[57]) & (!g121) & (!g213) & (g351)) + ((g119) & (!sk[57]) & (!g121) & (g213) & (!g351)) + ((g119) & (!sk[57]) & (!g121) & (g213) & (g351)) + ((g119) & (!sk[57]) & (g121) & (g213) & (!g351)) + ((g119) & (!sk[57]) & (g121) & (g213) & (g351)));
	assign g540 = (((!i_9_) & (!i_10_) & (!sk[58]) & (i_11_) & (!i_15_) & (g174)) + ((!i_9_) & (!i_10_) & (!sk[58]) & (i_11_) & (i_15_) & (!g174)) + ((!i_9_) & (!i_10_) & (!sk[58]) & (i_11_) & (i_15_) & (g174)) + ((!i_9_) & (!i_10_) & (sk[58]) & (!i_11_) & (i_15_) & (!g174)) + ((!i_9_) & (i_10_) & (!sk[58]) & (!i_11_) & (!i_15_) & (!g174)) + ((!i_9_) & (i_10_) & (!sk[58]) & (!i_11_) & (!i_15_) & (g174)) + ((!i_9_) & (i_10_) & (!sk[58]) & (!i_11_) & (i_15_) & (!g174)) + ((!i_9_) & (i_10_) & (!sk[58]) & (!i_11_) & (i_15_) & (g174)) + ((!i_9_) & (i_10_) & (!sk[58]) & (i_11_) & (!i_15_) & (!g174)) + ((!i_9_) & (i_10_) & (!sk[58]) & (i_11_) & (!i_15_) & (g174)) + ((!i_9_) & (i_10_) & (!sk[58]) & (i_11_) & (i_15_) & (!g174)) + ((!i_9_) & (i_10_) & (!sk[58]) & (i_11_) & (i_15_) & (g174)) + ((i_9_) & (!i_10_) & (!sk[58]) & (i_11_) & (!i_15_) & (g174)) + ((i_9_) & (!i_10_) & (!sk[58]) & (i_11_) & (i_15_) & (!g174)) + ((i_9_) & (!i_10_) & (!sk[58]) & (i_11_) & (i_15_) & (g174)) + ((i_9_) & (i_10_) & (!sk[58]) & (!i_11_) & (!i_15_) & (!g174)) + ((i_9_) & (i_10_) & (!sk[58]) & (!i_11_) & (!i_15_) & (g174)) + ((i_9_) & (i_10_) & (!sk[58]) & (!i_11_) & (i_15_) & (!g174)) + ((i_9_) & (i_10_) & (!sk[58]) & (!i_11_) & (i_15_) & (g174)) + ((i_9_) & (i_10_) & (!sk[58]) & (i_11_) & (!i_15_) & (!g174)) + ((i_9_) & (i_10_) & (!sk[58]) & (i_11_) & (!i_15_) & (g174)) + ((i_9_) & (i_10_) & (!sk[58]) & (i_11_) & (i_15_) & (!g174)) + ((i_9_) & (i_10_) & (!sk[58]) & (i_11_) & (i_15_) & (g174)) + ((i_9_) & (i_10_) & (sk[58]) & (i_11_) & (i_15_) & (!g174)));
	assign g541 = (((!g69) & (!g254) & (!g402) & (!g487) & (!g539) & (g540)) + ((!g69) & (!g254) & (!g402) & (g487) & (!g539) & (g540)) + ((!g69) & (!g254) & (!g402) & (g487) & (g539) & (g540)) + ((!g69) & (!g254) & (g402) & (!g487) & (!g539) & (g540)) + ((!g69) & (!g254) & (g402) & (g487) & (!g539) & (g540)) + ((!g69) & (!g254) & (g402) & (g487) & (g539) & (g540)) + ((!g69) & (g254) & (!g402) & (!g487) & (!g539) & (g540)) + ((!g69) & (g254) & (!g402) & (g487) & (!g539) & (g540)) + ((!g69) & (g254) & (!g402) & (g487) & (g539) & (g540)) + ((g69) & (!g254) & (!g402) & (!g487) & (!g539) & (g540)) + ((g69) & (!g254) & (!g402) & (g487) & (!g539) & (g540)) + ((g69) & (!g254) & (!g402) & (g487) & (g539) & (g540)) + ((g69) & (!g254) & (g402) & (!g487) & (!g539) & (g540)) + ((g69) & (!g254) & (g402) & (g487) & (!g539) & (g540)) + ((g69) & (!g254) & (g402) & (g487) & (g539) & (g540)) + ((g69) & (g254) & (!g402) & (!g487) & (!g539) & (g540)) + ((g69) & (g254) & (!g402) & (g487) & (!g539) & (g540)) + ((g69) & (g254) & (!g402) & (g487) & (g539) & (g540)) + ((g69) & (g254) & (g402) & (!g487) & (!g539) & (g540)) + ((g69) & (g254) & (g402) & (g487) & (!g539) & (g540)));
	assign g542 = (((!g105) & (!g186) & (!g513) & (sk[60]) & (!g514)) + ((!g105) & (!g186) & (!g513) & (sk[60]) & (g514)) + ((!g105) & (!g186) & (g513) & (!sk[60]) & (!g514)) + ((!g105) & (!g186) & (g513) & (!sk[60]) & (g514)) + ((!g105) & (!g186) & (g513) & (sk[60]) & (g514)) + ((!g105) & (g186) & (!g513) & (sk[60]) & (!g514)) + ((!g105) & (g186) & (!g513) & (sk[60]) & (g514)) + ((!g105) & (g186) & (g513) & (!sk[60]) & (!g514)) + ((!g105) & (g186) & (g513) & (!sk[60]) & (g514)) + ((!g105) & (g186) & (g513) & (sk[60]) & (!g514)) + ((!g105) & (g186) & (g513) & (sk[60]) & (g514)) + ((g105) & (!g186) & (g513) & (!sk[60]) & (!g514)) + ((g105) & (!g186) & (g513) & (!sk[60]) & (g514)) + ((g105) & (g186) & (g513) & (!sk[60]) & (!g514)) + ((g105) & (g186) & (g513) & (!sk[60]) & (g514)));
	assign g543 = (((!sk[61]) & (g76) & (!g81)) + ((!sk[61]) & (g76) & (g81)) + ((sk[61]) & (!g76) & (g81)));
	assign g544 = (((!g105) & (!sk[62]) & (!g182) & (g543) & (!g473)) + ((!g105) & (!sk[62]) & (!g182) & (g543) & (g473)) + ((!g105) & (!sk[62]) & (g182) & (g543) & (!g473)) + ((!g105) & (!sk[62]) & (g182) & (g543) & (g473)) + ((!g105) & (sk[62]) & (!g182) & (!g543) & (g473)) + ((!g105) & (sk[62]) & (!g182) & (g543) & (!g473)) + ((!g105) & (sk[62]) & (!g182) & (g543) & (g473)) + ((!g105) & (sk[62]) & (g182) & (!g543) & (!g473)) + ((!g105) & (sk[62]) & (g182) & (!g543) & (g473)) + ((!g105) & (sk[62]) & (g182) & (g543) & (!g473)) + ((!g105) & (sk[62]) & (g182) & (g543) & (g473)) + ((g105) & (!sk[62]) & (!g182) & (g543) & (!g473)) + ((g105) & (!sk[62]) & (!g182) & (g543) & (g473)) + ((g105) & (!sk[62]) & (g182) & (g543) & (!g473)) + ((g105) & (!sk[62]) & (g182) & (g543) & (g473)));
	assign g545 = (((!g22) & (!g69) & (!g113) & (sk[63]) & (!g105) & (g482)) + ((!g22) & (!g69) & (g113) & (!sk[63]) & (!g105) & (g482)) + ((!g22) & (!g69) & (g113) & (!sk[63]) & (g105) & (!g482)) + ((!g22) & (!g69) & (g113) & (!sk[63]) & (g105) & (g482)) + ((!g22) & (!g69) & (g113) & (sk[63]) & (!g105) & (g482)) + ((!g22) & (g69) & (!g113) & (!sk[63]) & (!g105) & (!g482)) + ((!g22) & (g69) & (!g113) & (!sk[63]) & (!g105) & (g482)) + ((!g22) & (g69) & (!g113) & (!sk[63]) & (g105) & (!g482)) + ((!g22) & (g69) & (!g113) & (!sk[63]) & (g105) & (g482)) + ((!g22) & (g69) & (!g113) & (sk[63]) & (!g105) & (g482)) + ((!g22) & (g69) & (g113) & (!sk[63]) & (!g105) & (!g482)) + ((!g22) & (g69) & (g113) & (!sk[63]) & (!g105) & (g482)) + ((!g22) & (g69) & (g113) & (!sk[63]) & (g105) & (!g482)) + ((!g22) & (g69) & (g113) & (!sk[63]) & (g105) & (g482)) + ((!g22) & (g69) & (g113) & (sk[63]) & (!g105) & (g482)) + ((g22) & (!g69) & (!g113) & (sk[63]) & (!g105) & (g482)) + ((g22) & (!g69) & (g113) & (!sk[63]) & (!g105) & (g482)) + ((g22) & (!g69) & (g113) & (!sk[63]) & (g105) & (!g482)) + ((g22) & (!g69) & (g113) & (!sk[63]) & (g105) & (g482)) + ((g22) & (g69) & (!g113) & (!sk[63]) & (!g105) & (!g482)) + ((g22) & (g69) & (!g113) & (!sk[63]) & (!g105) & (g482)) + ((g22) & (g69) & (!g113) & (!sk[63]) & (g105) & (!g482)) + ((g22) & (g69) & (!g113) & (!sk[63]) & (g105) & (g482)) + ((g22) & (g69) & (!g113) & (sk[63]) & (!g105) & (g482)) + ((g22) & (g69) & (g113) & (!sk[63]) & (!g105) & (!g482)) + ((g22) & (g69) & (g113) & (!sk[63]) & (!g105) & (g482)) + ((g22) & (g69) & (g113) & (!sk[63]) & (g105) & (!g482)) + ((g22) & (g69) & (g113) & (!sk[63]) & (g105) & (g482)) + ((g22) & (g69) & (g113) & (sk[63]) & (!g105) & (g482)));
	assign g546 = (((!g105) & (!sk[64]) & (!g487) & (g484) & (!g522)) + ((!g105) & (!sk[64]) & (!g487) & (g484) & (g522)) + ((!g105) & (!sk[64]) & (g487) & (g484) & (!g522)) + ((!g105) & (!sk[64]) & (g487) & (g484) & (g522)) + ((!g105) & (sk[64]) & (!g487) & (!g484) & (g522)) + ((!g105) & (sk[64]) & (!g487) & (g484) & (!g522)) + ((!g105) & (sk[64]) & (!g487) & (g484) & (g522)) + ((!g105) & (sk[64]) & (g487) & (!g484) & (!g522)) + ((!g105) & (sk[64]) & (g487) & (!g484) & (g522)) + ((!g105) & (sk[64]) & (g487) & (g484) & (!g522)) + ((!g105) & (sk[64]) & (g487) & (g484) & (g522)) + ((g105) & (!sk[64]) & (!g487) & (g484) & (!g522)) + ((g105) & (!sk[64]) & (!g487) & (g484) & (g522)) + ((g105) & (!sk[64]) & (g487) & (g484) & (!g522)) + ((g105) & (!sk[64]) & (g487) & (g484) & (g522)));
	assign g547 = (((!g102) & (!g483) & (!sk[65]) & (g489) & (!g484) & (g500)) + ((!g102) & (!g483) & (!sk[65]) & (g489) & (g484) & (!g500)) + ((!g102) & (!g483) & (!sk[65]) & (g489) & (g484) & (g500)) + ((!g102) & (g483) & (!sk[65]) & (!g489) & (!g484) & (!g500)) + ((!g102) & (g483) & (!sk[65]) & (!g489) & (!g484) & (g500)) + ((!g102) & (g483) & (!sk[65]) & (!g489) & (g484) & (!g500)) + ((!g102) & (g483) & (!sk[65]) & (!g489) & (g484) & (g500)) + ((!g102) & (g483) & (!sk[65]) & (g489) & (!g484) & (!g500)) + ((!g102) & (g483) & (!sk[65]) & (g489) & (!g484) & (g500)) + ((!g102) & (g483) & (!sk[65]) & (g489) & (g484) & (!g500)) + ((!g102) & (g483) & (!sk[65]) & (g489) & (g484) & (g500)) + ((g102) & (!g483) & (!sk[65]) & (g489) & (!g484) & (g500)) + ((g102) & (!g483) & (!sk[65]) & (g489) & (g484) & (!g500)) + ((g102) & (!g483) & (!sk[65]) & (g489) & (g484) & (g500)) + ((g102) & (!g483) & (sk[65]) & (!g489) & (!g484) & (g500)) + ((g102) & (!g483) & (sk[65]) & (!g489) & (g484) & (!g500)) + ((g102) & (!g483) & (sk[65]) & (!g489) & (g484) & (g500)) + ((g102) & (!g483) & (sk[65]) & (g489) & (!g484) & (!g500)) + ((g102) & (!g483) & (sk[65]) & (g489) & (!g484) & (g500)) + ((g102) & (!g483) & (sk[65]) & (g489) & (g484) & (!g500)) + ((g102) & (!g483) & (sk[65]) & (g489) & (g484) & (g500)) + ((g102) & (g483) & (!sk[65]) & (!g489) & (!g484) & (!g500)) + ((g102) & (g483) & (!sk[65]) & (!g489) & (!g484) & (g500)) + ((g102) & (g483) & (!sk[65]) & (!g489) & (g484) & (!g500)) + ((g102) & (g483) & (!sk[65]) & (!g489) & (g484) & (g500)) + ((g102) & (g483) & (!sk[65]) & (g489) & (!g484) & (!g500)) + ((g102) & (g483) & (!sk[65]) & (g489) & (!g484) & (g500)) + ((g102) & (g483) & (!sk[65]) & (g489) & (g484) & (!g500)) + ((g102) & (g483) & (!sk[65]) & (g489) & (g484) & (g500)) + ((g102) & (g483) & (sk[65]) & (!g489) & (!g484) & (!g500)) + ((g102) & (g483) & (sk[65]) & (!g489) & (!g484) & (g500)) + ((g102) & (g483) & (sk[65]) & (!g489) & (g484) & (!g500)) + ((g102) & (g483) & (sk[65]) & (!g489) & (g484) & (g500)) + ((g102) & (g483) & (sk[65]) & (g489) & (!g484) & (!g500)) + ((g102) & (g483) & (sk[65]) & (g489) & (!g484) & (g500)) + ((g102) & (g483) & (sk[65]) & (g489) & (g484) & (!g500)) + ((g102) & (g483) & (sk[65]) & (g489) & (g484) & (g500)));
	assign g548 = (((!g542) & (!g544) & (!sk[66]) & (g545) & (!g546) & (g547)) + ((!g542) & (!g544) & (!sk[66]) & (g545) & (g546) & (!g547)) + ((!g542) & (!g544) & (!sk[66]) & (g545) & (g546) & (g547)) + ((!g542) & (!g544) & (sk[66]) & (!g545) & (!g546) & (!g547)) + ((!g542) & (g544) & (!sk[66]) & (!g545) & (!g546) & (!g547)) + ((!g542) & (g544) & (!sk[66]) & (!g545) & (!g546) & (g547)) + ((!g542) & (g544) & (!sk[66]) & (!g545) & (g546) & (!g547)) + ((!g542) & (g544) & (!sk[66]) & (!g545) & (g546) & (g547)) + ((!g542) & (g544) & (!sk[66]) & (g545) & (!g546) & (!g547)) + ((!g542) & (g544) & (!sk[66]) & (g545) & (!g546) & (g547)) + ((!g542) & (g544) & (!sk[66]) & (g545) & (g546) & (!g547)) + ((!g542) & (g544) & (!sk[66]) & (g545) & (g546) & (g547)) + ((g542) & (!g544) & (!sk[66]) & (g545) & (!g546) & (g547)) + ((g542) & (!g544) & (!sk[66]) & (g545) & (g546) & (!g547)) + ((g542) & (!g544) & (!sk[66]) & (g545) & (g546) & (g547)) + ((g542) & (g544) & (!sk[66]) & (!g545) & (!g546) & (!g547)) + ((g542) & (g544) & (!sk[66]) & (!g545) & (!g546) & (g547)) + ((g542) & (g544) & (!sk[66]) & (!g545) & (g546) & (!g547)) + ((g542) & (g544) & (!sk[66]) & (!g545) & (g546) & (g547)) + ((g542) & (g544) & (!sk[66]) & (g545) & (!g546) & (!g547)) + ((g542) & (g544) & (!sk[66]) & (g545) & (!g546) & (g547)) + ((g542) & (g544) & (!sk[66]) & (g545) & (g546) & (!g547)) + ((g542) & (g544) & (!sk[66]) & (g545) & (g546) & (g547)));
	assign g549 = (((!g538) & (!sk[67]) & (!g541) & (g548)) + ((!g538) & (!sk[67]) & (g541) & (!g548)) + ((!g538) & (!sk[67]) & (g541) & (g548)) + ((!g538) & (sk[67]) & (!g541) & (g548)) + ((g538) & (!sk[67]) & (!g541) & (g548)) + ((g538) & (!sk[67]) & (g541) & (!g548)) + ((g538) & (!sk[67]) & (g541) & (g548)));
	assign g550 = (((!g17) & (!g22) & (!g81) & (!g142) & (!g174) & (!g351)) + ((!g17) & (!g22) & (!g81) & (!g142) & (!g174) & (g351)) + ((!g17) & (!g22) & (!g81) & (g142) & (!g174) & (!g351)) + ((!g17) & (!g22) & (g81) & (!g142) & (!g174) & (!g351)) + ((!g17) & (!g22) & (g81) & (!g142) & (!g174) & (g351)) + ((!g17) & (!g22) & (g81) & (g142) & (!g174) & (!g351)) + ((!g17) & (g22) & (g81) & (!g142) & (!g174) & (!g351)) + ((!g17) & (g22) & (g81) & (!g142) & (!g174) & (g351)) + ((!g17) & (g22) & (g81) & (g142) & (!g174) & (!g351)) + ((g17) & (!g22) & (!g81) & (!g142) & (!g174) & (!g351)) + ((g17) & (!g22) & (!g81) & (!g142) & (!g174) & (g351)) + ((g17) & (!g22) & (!g81) & (g142) & (!g174) & (!g351)) + ((g17) & (!g22) & (g81) & (!g142) & (!g174) & (!g351)) + ((g17) & (!g22) & (g81) & (!g142) & (!g174) & (g351)) + ((g17) & (!g22) & (g81) & (g142) & (!g174) & (!g351)) + ((g17) & (g22) & (!g81) & (!g142) & (!g174) & (!g351)) + ((g17) & (g22) & (!g81) & (!g142) & (!g174) & (g351)) + ((g17) & (g22) & (!g81) & (g142) & (!g174) & (!g351)) + ((g17) & (g22) & (g81) & (!g142) & (!g174) & (!g351)) + ((g17) & (g22) & (g81) & (!g142) & (!g174) & (g351)) + ((g17) & (g22) & (g81) & (g142) & (!g174) & (!g351)));
	assign g551 = (((!sk[69]) & (g22) & (!g76)) + ((!sk[69]) & (g22) & (g76)) + ((sk[69]) & (!g22) & (g76)) + ((sk[69]) & (g22) & (!g76)) + ((sk[69]) & (g22) & (g76)));
	assign g552 = (((!g76) & (sk[70]) & (!g69)) + ((g76) & (!sk[70]) & (!g69)) + ((g76) & (!sk[70]) & (g69)) + ((g76) & (sk[70]) & (!g69)) + ((g76) & (sk[70]) & (g69)));
	assign g553 = (((!g17) & (!sk[71]) & (!g76) & (g135) & (!g88) & (g460)) + ((!g17) & (!sk[71]) & (!g76) & (g135) & (g88) & (!g460)) + ((!g17) & (!sk[71]) & (!g76) & (g135) & (g88) & (g460)) + ((!g17) & (!sk[71]) & (g76) & (!g135) & (!g88) & (!g460)) + ((!g17) & (!sk[71]) & (g76) & (!g135) & (!g88) & (g460)) + ((!g17) & (!sk[71]) & (g76) & (!g135) & (g88) & (!g460)) + ((!g17) & (!sk[71]) & (g76) & (!g135) & (g88) & (g460)) + ((!g17) & (!sk[71]) & (g76) & (g135) & (!g88) & (!g460)) + ((!g17) & (!sk[71]) & (g76) & (g135) & (!g88) & (g460)) + ((!g17) & (!sk[71]) & (g76) & (g135) & (g88) & (!g460)) + ((!g17) & (!sk[71]) & (g76) & (g135) & (g88) & (g460)) + ((!g17) & (sk[71]) & (!g76) & (!g135) & (!g88) & (!g460)) + ((!g17) & (sk[71]) & (!g76) & (!g135) & (!g88) & (g460)) + ((!g17) & (sk[71]) & (!g76) & (g135) & (!g88) & (!g460)) + ((!g17) & (sk[71]) & (!g76) & (g135) & (!g88) & (g460)) + ((!g17) & (sk[71]) & (!g76) & (g135) & (g88) & (!g460)) + ((!g17) & (sk[71]) & (!g76) & (g135) & (g88) & (g460)) + ((!g17) & (sk[71]) & (g76) & (!g135) & (!g88) & (!g460)) + ((!g17) & (sk[71]) & (g76) & (!g135) & (!g88) & (g460)) + ((!g17) & (sk[71]) & (g76) & (!g135) & (g88) & (!g460)) + ((!g17) & (sk[71]) & (g76) & (!g135) & (g88) & (g460)) + ((!g17) & (sk[71]) & (g76) & (g135) & (!g88) & (!g460)) + ((!g17) & (sk[71]) & (g76) & (g135) & (!g88) & (g460)) + ((!g17) & (sk[71]) & (g76) & (g135) & (g88) & (!g460)) + ((!g17) & (sk[71]) & (g76) & (g135) & (g88) & (g460)) + ((g17) & (!sk[71]) & (!g76) & (g135) & (!g88) & (g460)) + ((g17) & (!sk[71]) & (!g76) & (g135) & (g88) & (!g460)) + ((g17) & (!sk[71]) & (!g76) & (g135) & (g88) & (g460)) + ((g17) & (!sk[71]) & (g76) & (!g135) & (!g88) & (!g460)) + ((g17) & (!sk[71]) & (g76) & (!g135) & (!g88) & (g460)) + ((g17) & (!sk[71]) & (g76) & (!g135) & (g88) & (!g460)) + ((g17) & (!sk[71]) & (g76) & (!g135) & (g88) & (g460)) + ((g17) & (!sk[71]) & (g76) & (g135) & (!g88) & (!g460)) + ((g17) & (!sk[71]) & (g76) & (g135) & (!g88) & (g460)) + ((g17) & (!sk[71]) & (g76) & (g135) & (g88) & (!g460)) + ((g17) & (!sk[71]) & (g76) & (g135) & (g88) & (g460)) + ((g17) & (sk[71]) & (!g76) & (g135) & (!g88) & (!g460)) + ((g17) & (sk[71]) & (!g76) & (g135) & (!g88) & (g460)) + ((g17) & (sk[71]) & (!g76) & (g135) & (g88) & (!g460)) + ((g17) & (sk[71]) & (!g76) & (g135) & (g88) & (g460)) + ((g17) & (sk[71]) & (g76) & (!g135) & (!g88) & (g460)) + ((g17) & (sk[71]) & (g76) & (!g135) & (g88) & (g460)) + ((g17) & (sk[71]) & (g76) & (g135) & (!g88) & (!g460)) + ((g17) & (sk[71]) & (g76) & (g135) & (!g88) & (g460)) + ((g17) & (sk[71]) & (g76) & (g135) & (g88) & (!g460)) + ((g17) & (sk[71]) & (g76) & (g135) & (g88) & (g460)));
	assign g554 = (((!g17) & (!g76) & (!g122) & (!g81) & (sk[72]) & (!g460)) + ((!g17) & (!g76) & (!g122) & (!g81) & (sk[72]) & (g460)) + ((!g17) & (!g76) & (!g122) & (g81) & (sk[72]) & (!g460)) + ((!g17) & (!g76) & (!g122) & (g81) & (sk[72]) & (g460)) + ((!g17) & (!g76) & (g122) & (!g81) & (!sk[72]) & (g460)) + ((!g17) & (!g76) & (g122) & (!g81) & (sk[72]) & (!g460)) + ((!g17) & (!g76) & (g122) & (!g81) & (sk[72]) & (g460)) + ((!g17) & (!g76) & (g122) & (g81) & (!sk[72]) & (!g460)) + ((!g17) & (!g76) & (g122) & (g81) & (!sk[72]) & (g460)) + ((!g17) & (g76) & (!g122) & (!g81) & (!sk[72]) & (!g460)) + ((!g17) & (g76) & (!g122) & (!g81) & (!sk[72]) & (g460)) + ((!g17) & (g76) & (!g122) & (!g81) & (sk[72]) & (!g460)) + ((!g17) & (g76) & (!g122) & (!g81) & (sk[72]) & (g460)) + ((!g17) & (g76) & (!g122) & (g81) & (!sk[72]) & (!g460)) + ((!g17) & (g76) & (!g122) & (g81) & (!sk[72]) & (g460)) + ((!g17) & (g76) & (!g122) & (g81) & (sk[72]) & (!g460)) + ((!g17) & (g76) & (!g122) & (g81) & (sk[72]) & (g460)) + ((!g17) & (g76) & (g122) & (!g81) & (!sk[72]) & (!g460)) + ((!g17) & (g76) & (g122) & (!g81) & (!sk[72]) & (g460)) + ((!g17) & (g76) & (g122) & (!g81) & (sk[72]) & (!g460)) + ((!g17) & (g76) & (g122) & (!g81) & (sk[72]) & (g460)) + ((!g17) & (g76) & (g122) & (g81) & (!sk[72]) & (!g460)) + ((!g17) & (g76) & (g122) & (g81) & (!sk[72]) & (g460)) + ((!g17) & (g76) & (g122) & (g81) & (sk[72]) & (g460)) + ((g17) & (!g76) & (!g122) & (!g81) & (sk[72]) & (!g460)) + ((g17) & (!g76) & (!g122) & (!g81) & (sk[72]) & (g460)) + ((g17) & (!g76) & (!g122) & (g81) & (sk[72]) & (!g460)) + ((g17) & (!g76) & (!g122) & (g81) & (sk[72]) & (g460)) + ((g17) & (!g76) & (g122) & (!g81) & (!sk[72]) & (g460)) + ((g17) & (!g76) & (g122) & (g81) & (!sk[72]) & (!g460)) + ((g17) & (!g76) & (g122) & (g81) & (!sk[72]) & (g460)) + ((g17) & (g76) & (!g122) & (!g81) & (!sk[72]) & (!g460)) + ((g17) & (g76) & (!g122) & (!g81) & (!sk[72]) & (g460)) + ((g17) & (g76) & (!g122) & (!g81) & (sk[72]) & (!g460)) + ((g17) & (g76) & (!g122) & (!g81) & (sk[72]) & (g460)) + ((g17) & (g76) & (!g122) & (g81) & (!sk[72]) & (!g460)) + ((g17) & (g76) & (!g122) & (g81) & (!sk[72]) & (g460)) + ((g17) & (g76) & (!g122) & (g81) & (sk[72]) & (!g460)) + ((g17) & (g76) & (!g122) & (g81) & (sk[72]) & (g460)) + ((g17) & (g76) & (g122) & (!g81) & (!sk[72]) & (!g460)) + ((g17) & (g76) & (g122) & (!g81) & (!sk[72]) & (g460)) + ((g17) & (g76) & (g122) & (!g81) & (sk[72]) & (g460)) + ((g17) & (g76) & (g122) & (g81) & (!sk[72]) & (!g460)) + ((g17) & (g76) & (g122) & (g81) & (!sk[72]) & (g460)) + ((g17) & (g76) & (g122) & (g81) & (sk[72]) & (g460)));
	assign g555 = (((g36) & (!sk[73]) & (!g460)) + ((g36) & (!sk[73]) & (g460)) + ((g36) & (sk[73]) & (!g460)));
	assign g556 = (((!g102) & (!g105) & (!g555) & (!g501) & (!g543) & (!g534)) + ((!g102) & (!g105) & (!g555) & (!g501) & (!g543) & (g534)) + ((!g102) & (!g105) & (!g555) & (!g501) & (g543) & (!g534)) + ((!g102) & (!g105) & (!g555) & (!g501) & (g543) & (g534)) + ((!g102) & (g105) & (!g555) & (!g501) & (!g543) & (!g534)) + ((!g102) & (g105) & (!g555) & (!g501) & (!g543) & (g534)) + ((!g102) & (g105) & (!g555) & (!g501) & (g543) & (!g534)) + ((!g102) & (g105) & (!g555) & (!g501) & (g543) & (g534)) + ((!g102) & (g105) & (!g555) & (g501) & (!g543) & (!g534)) + ((!g102) & (g105) & (!g555) & (g501) & (!g543) & (g534)) + ((!g102) & (g105) & (!g555) & (g501) & (g543) & (!g534)) + ((!g102) & (g105) & (!g555) & (g501) & (g543) & (g534)) + ((!g102) & (g105) & (g555) & (!g501) & (!g543) & (!g534)) + ((!g102) & (g105) & (g555) & (!g501) & (!g543) & (g534)) + ((!g102) & (g105) & (g555) & (!g501) & (g543) & (!g534)) + ((!g102) & (g105) & (g555) & (!g501) & (g543) & (g534)) + ((!g102) & (g105) & (g555) & (g501) & (!g543) & (!g534)) + ((!g102) & (g105) & (g555) & (g501) & (!g543) & (g534)) + ((!g102) & (g105) & (g555) & (g501) & (g543) & (!g534)) + ((!g102) & (g105) & (g555) & (g501) & (g543) & (g534)) + ((g102) & (!g105) & (!g555) & (!g501) & (!g543) & (!g534)) + ((g102) & (g105) & (!g555) & (!g501) & (!g543) & (!g534)));
	assign g557 = (((!sk[75]) & (g76) & (!g113)) + ((!sk[75]) & (g76) & (g113)) + ((sk[75]) & (!g76) & (!g113)));
	assign g558 = (((!g125) & (!g122) & (!g123) & (g552) & (!g511) & (!g557)) + ((!g125) & (!g122) & (g123) & (!g552) & (!g511) & (!g557)) + ((!g125) & (!g122) & (g123) & (!g552) & (!g511) & (g557)) + ((!g125) & (!g122) & (g123) & (!g552) & (g511) & (!g557)) + ((!g125) & (!g122) & (g123) & (!g552) & (g511) & (g557)) + ((!g125) & (!g122) & (g123) & (g552) & (!g511) & (!g557)) + ((!g125) & (!g122) & (g123) & (g552) & (!g511) & (g557)) + ((!g125) & (!g122) & (g123) & (g552) & (g511) & (!g557)) + ((!g125) & (!g122) & (g123) & (g552) & (g511) & (g557)) + ((!g125) & (g122) & (!g123) & (g552) & (!g511) & (!g557)) + ((!g125) & (g122) & (g123) & (!g552) & (!g511) & (!g557)) + ((!g125) & (g122) & (g123) & (!g552) & (g511) & (!g557)) + ((!g125) & (g122) & (g123) & (g552) & (!g511) & (!g557)) + ((!g125) & (g122) & (g123) & (g552) & (g511) & (!g557)) + ((g125) & (!g122) & (!g123) & (g552) & (!g511) & (!g557)) + ((g125) & (!g122) & (g123) & (g552) & (!g511) & (!g557)) + ((g125) & (!g122) & (g123) & (g552) & (g511) & (!g557)) + ((g125) & (g122) & (!g123) & (g552) & (!g511) & (!g557)) + ((g125) & (g122) & (g123) & (g552) & (!g511) & (!g557)) + ((g125) & (g122) & (g123) & (g552) & (g511) & (!g557)));
	assign g559 = (((!sk[77]) & (!g119) & (!g121) & (g552) & (!g511) & (g558)) + ((!sk[77]) & (!g119) & (!g121) & (g552) & (g511) & (!g558)) + ((!sk[77]) & (!g119) & (!g121) & (g552) & (g511) & (g558)) + ((!sk[77]) & (!g119) & (g121) & (!g552) & (!g511) & (!g558)) + ((!sk[77]) & (!g119) & (g121) & (!g552) & (!g511) & (g558)) + ((!sk[77]) & (!g119) & (g121) & (!g552) & (g511) & (!g558)) + ((!sk[77]) & (!g119) & (g121) & (!g552) & (g511) & (g558)) + ((!sk[77]) & (!g119) & (g121) & (g552) & (!g511) & (!g558)) + ((!sk[77]) & (!g119) & (g121) & (g552) & (!g511) & (g558)) + ((!sk[77]) & (!g119) & (g121) & (g552) & (g511) & (!g558)) + ((!sk[77]) & (!g119) & (g121) & (g552) & (g511) & (g558)) + ((!sk[77]) & (g119) & (!g121) & (g552) & (!g511) & (g558)) + ((!sk[77]) & (g119) & (!g121) & (g552) & (g511) & (!g558)) + ((!sk[77]) & (g119) & (!g121) & (g552) & (g511) & (g558)) + ((!sk[77]) & (g119) & (g121) & (!g552) & (!g511) & (!g558)) + ((!sk[77]) & (g119) & (g121) & (!g552) & (!g511) & (g558)) + ((!sk[77]) & (g119) & (g121) & (!g552) & (g511) & (!g558)) + ((!sk[77]) & (g119) & (g121) & (!g552) & (g511) & (g558)) + ((!sk[77]) & (g119) & (g121) & (g552) & (!g511) & (!g558)) + ((!sk[77]) & (g119) & (g121) & (g552) & (!g511) & (g558)) + ((!sk[77]) & (g119) & (g121) & (g552) & (g511) & (!g558)) + ((!sk[77]) & (g119) & (g121) & (g552) & (g511) & (g558)) + ((sk[77]) & (!g119) & (!g121) & (!g552) & (!g511) & (g558)) + ((sk[77]) & (!g119) & (!g121) & (!g552) & (g511) & (g558)) + ((sk[77]) & (!g119) & (!g121) & (g552) & (!g511) & (g558)) + ((sk[77]) & (!g119) & (!g121) & (g552) & (g511) & (g558)) + ((sk[77]) & (!g119) & (g121) & (g552) & (!g511) & (g558)) + ((sk[77]) & (g119) & (!g121) & (!g552) & (!g511) & (g558)) + ((sk[77]) & (g119) & (!g121) & (g552) & (!g511) & (g558)) + ((sk[77]) & (g119) & (g121) & (g552) & (!g511) & (g558)));
	assign g560 = (((!g76) & (!sk[78]) & (!g161) & (g122) & (!g91) & (g88)) + ((!g76) & (!sk[78]) & (!g161) & (g122) & (g91) & (!g88)) + ((!g76) & (!sk[78]) & (!g161) & (g122) & (g91) & (g88)) + ((!g76) & (!sk[78]) & (g161) & (!g122) & (!g91) & (!g88)) + ((!g76) & (!sk[78]) & (g161) & (!g122) & (!g91) & (g88)) + ((!g76) & (!sk[78]) & (g161) & (!g122) & (g91) & (!g88)) + ((!g76) & (!sk[78]) & (g161) & (!g122) & (g91) & (g88)) + ((!g76) & (!sk[78]) & (g161) & (g122) & (!g91) & (!g88)) + ((!g76) & (!sk[78]) & (g161) & (g122) & (!g91) & (g88)) + ((!g76) & (!sk[78]) & (g161) & (g122) & (g91) & (!g88)) + ((!g76) & (!sk[78]) & (g161) & (g122) & (g91) & (g88)) + ((!g76) & (sk[78]) & (!g161) & (g122) & (!g91) & (!g88)) + ((!g76) & (sk[78]) & (!g161) & (g122) & (!g91) & (g88)) + ((!g76) & (sk[78]) & (!g161) & (g122) & (g91) & (g88)) + ((!g76) & (sk[78]) & (g161) & (!g122) & (!g91) & (g88)) + ((!g76) & (sk[78]) & (g161) & (!g122) & (g91) & (g88)) + ((!g76) & (sk[78]) & (g161) & (g122) & (!g91) & (!g88)) + ((!g76) & (sk[78]) & (g161) & (g122) & (!g91) & (g88)) + ((!g76) & (sk[78]) & (g161) & (g122) & (g91) & (g88)) + ((g76) & (!sk[78]) & (!g161) & (g122) & (!g91) & (g88)) + ((g76) & (!sk[78]) & (!g161) & (g122) & (g91) & (!g88)) + ((g76) & (!sk[78]) & (!g161) & (g122) & (g91) & (g88)) + ((g76) & (!sk[78]) & (g161) & (!g122) & (!g91) & (!g88)) + ((g76) & (!sk[78]) & (g161) & (!g122) & (!g91) & (g88)) + ((g76) & (!sk[78]) & (g161) & (!g122) & (g91) & (!g88)) + ((g76) & (!sk[78]) & (g161) & (!g122) & (g91) & (g88)) + ((g76) & (!sk[78]) & (g161) & (g122) & (!g91) & (!g88)) + ((g76) & (!sk[78]) & (g161) & (g122) & (!g91) & (g88)) + ((g76) & (!sk[78]) & (g161) & (g122) & (g91) & (!g88)) + ((g76) & (!sk[78]) & (g161) & (g122) & (g91) & (g88)));
	assign g561 = (((!g17) & (!g88) & (!sk[79]) & (g113) & (!g105) & (g460)) + ((!g17) & (!g88) & (!sk[79]) & (g113) & (g105) & (!g460)) + ((!g17) & (!g88) & (!sk[79]) & (g113) & (g105) & (g460)) + ((!g17) & (!g88) & (sk[79]) & (!g113) & (!g105) & (!g460)) + ((!g17) & (g88) & (!sk[79]) & (!g113) & (!g105) & (!g460)) + ((!g17) & (g88) & (!sk[79]) & (!g113) & (!g105) & (g460)) + ((!g17) & (g88) & (!sk[79]) & (!g113) & (g105) & (!g460)) + ((!g17) & (g88) & (!sk[79]) & (!g113) & (g105) & (g460)) + ((!g17) & (g88) & (!sk[79]) & (g113) & (!g105) & (!g460)) + ((!g17) & (g88) & (!sk[79]) & (g113) & (!g105) & (g460)) + ((!g17) & (g88) & (!sk[79]) & (g113) & (g105) & (!g460)) + ((!g17) & (g88) & (!sk[79]) & (g113) & (g105) & (g460)) + ((!g17) & (g88) & (sk[79]) & (!g113) & (!g105) & (!g460)) + ((!g17) & (g88) & (sk[79]) & (g113) & (!g105) & (!g460)) + ((g17) & (!g88) & (!sk[79]) & (g113) & (!g105) & (g460)) + ((g17) & (!g88) & (!sk[79]) & (g113) & (g105) & (!g460)) + ((g17) & (!g88) & (!sk[79]) & (g113) & (g105) & (g460)) + ((g17) & (!g88) & (sk[79]) & (!g113) & (!g105) & (!g460)) + ((g17) & (!g88) & (sk[79]) & (g113) & (!g105) & (!g460)) + ((g17) & (g88) & (!sk[79]) & (!g113) & (!g105) & (!g460)) + ((g17) & (g88) & (!sk[79]) & (!g113) & (!g105) & (g460)) + ((g17) & (g88) & (!sk[79]) & (!g113) & (g105) & (!g460)) + ((g17) & (g88) & (!sk[79]) & (!g113) & (g105) & (g460)) + ((g17) & (g88) & (!sk[79]) & (g113) & (!g105) & (!g460)) + ((g17) & (g88) & (!sk[79]) & (g113) & (!g105) & (g460)) + ((g17) & (g88) & (!sk[79]) & (g113) & (g105) & (!g460)) + ((g17) & (g88) & (!sk[79]) & (g113) & (g105) & (g460)) + ((g17) & (g88) & (sk[79]) & (!g113) & (!g105) & (!g460)) + ((g17) & (g88) & (sk[79]) & (g113) & (!g105) & (!g460)));
	assign g562 = (((!sk[80]) & (g76) & (!g91)) + ((!sk[80]) & (g76) & (g91)) + ((sk[80]) & (!g76) & (!g91)));
	assign g563 = (((!i_8_) & (!sk[81]) & (!g73) & (g486) & (!g562)) + ((!i_8_) & (!sk[81]) & (!g73) & (g486) & (g562)) + ((!i_8_) & (!sk[81]) & (g73) & (g486) & (!g562)) + ((!i_8_) & (!sk[81]) & (g73) & (g486) & (g562)) + ((!i_8_) & (sk[81]) & (g73) & (!g486) & (g562)) + ((!i_8_) & (sk[81]) & (g73) & (g486) & (!g562)) + ((!i_8_) & (sk[81]) & (g73) & (g486) & (g562)) + ((i_8_) & (!sk[81]) & (!g73) & (g486) & (!g562)) + ((i_8_) & (!sk[81]) & (!g73) & (g486) & (g562)) + ((i_8_) & (!sk[81]) & (g73) & (g486) & (!g562)) + ((i_8_) & (!sk[81]) & (g73) & (g486) & (g562)));
	assign g564 = (((!g123) & (!g555) & (!sk[82]) & (g486)) + ((!g123) & (!g555) & (sk[82]) & (g486)) + ((!g123) & (g555) & (!sk[82]) & (!g486)) + ((!g123) & (g555) & (!sk[82]) & (g486)) + ((!g123) & (g555) & (sk[82]) & (!g486)) + ((!g123) & (g555) & (sk[82]) & (g486)) + ((g123) & (!g555) & (!sk[82]) & (g486)) + ((g123) & (g555) & (!sk[82]) & (!g486)) + ((g123) & (g555) & (!sk[82]) & (g486)));
	assign g565 = (((!g36) & (!g76) & (!sk[83]) & (g88) & (!g130) & (g460)) + ((!g36) & (!g76) & (!sk[83]) & (g88) & (g130) & (!g460)) + ((!g36) & (!g76) & (!sk[83]) & (g88) & (g130) & (g460)) + ((!g36) & (!g76) & (sk[83]) & (g88) & (!g130) & (!g460)) + ((!g36) & (!g76) & (sk[83]) & (g88) & (!g130) & (g460)) + ((!g36) & (g76) & (!sk[83]) & (!g88) & (!g130) & (!g460)) + ((!g36) & (g76) & (!sk[83]) & (!g88) & (!g130) & (g460)) + ((!g36) & (g76) & (!sk[83]) & (!g88) & (g130) & (!g460)) + ((!g36) & (g76) & (!sk[83]) & (!g88) & (g130) & (g460)) + ((!g36) & (g76) & (!sk[83]) & (g88) & (!g130) & (!g460)) + ((!g36) & (g76) & (!sk[83]) & (g88) & (!g130) & (g460)) + ((!g36) & (g76) & (!sk[83]) & (g88) & (g130) & (!g460)) + ((!g36) & (g76) & (!sk[83]) & (g88) & (g130) & (g460)) + ((g36) & (!g76) & (!sk[83]) & (g88) & (!g130) & (g460)) + ((g36) & (!g76) & (!sk[83]) & (g88) & (g130) & (!g460)) + ((g36) & (!g76) & (!sk[83]) & (g88) & (g130) & (g460)) + ((g36) & (!g76) & (sk[83]) & (!g88) & (!g130) & (!g460)) + ((g36) & (!g76) & (sk[83]) & (!g88) & (!g130) & (g460)) + ((g36) & (!g76) & (sk[83]) & (g88) & (!g130) & (!g460)) + ((g36) & (!g76) & (sk[83]) & (g88) & (!g130) & (g460)) + ((g36) & (g76) & (!sk[83]) & (!g88) & (!g130) & (!g460)) + ((g36) & (g76) & (!sk[83]) & (!g88) & (!g130) & (g460)) + ((g36) & (g76) & (!sk[83]) & (!g88) & (g130) & (!g460)) + ((g36) & (g76) & (!sk[83]) & (!g88) & (g130) & (g460)) + ((g36) & (g76) & (!sk[83]) & (g88) & (!g130) & (!g460)) + ((g36) & (g76) & (!sk[83]) & (g88) & (!g130) & (g460)) + ((g36) & (g76) & (!sk[83]) & (g88) & (g130) & (!g460)) + ((g36) & (g76) & (!sk[83]) & (g88) & (g130) & (g460)) + ((g36) & (g76) & (sk[83]) & (!g88) & (!g130) & (!g460)) + ((g36) & (g76) & (sk[83]) & (g88) & (!g130) & (!g460)));
	assign g566 = (((!g76) & (!sk[84]) & (!g81) & (g91) & (!g130) & (g460)) + ((!g76) & (!sk[84]) & (!g81) & (g91) & (g130) & (!g460)) + ((!g76) & (!sk[84]) & (!g81) & (g91) & (g130) & (g460)) + ((!g76) & (!sk[84]) & (g81) & (!g91) & (!g130) & (!g460)) + ((!g76) & (!sk[84]) & (g81) & (!g91) & (!g130) & (g460)) + ((!g76) & (!sk[84]) & (g81) & (!g91) & (g130) & (!g460)) + ((!g76) & (!sk[84]) & (g81) & (!g91) & (g130) & (g460)) + ((!g76) & (!sk[84]) & (g81) & (g91) & (!g130) & (!g460)) + ((!g76) & (!sk[84]) & (g81) & (g91) & (!g130) & (g460)) + ((!g76) & (!sk[84]) & (g81) & (g91) & (g130) & (!g460)) + ((!g76) & (!sk[84]) & (g81) & (g91) & (g130) & (g460)) + ((!g76) & (sk[84]) & (!g81) & (!g91) & (!g130) & (!g460)) + ((!g76) & (sk[84]) & (!g81) & (!g91) & (!g130) & (g460)) + ((!g76) & (sk[84]) & (g81) & (!g91) & (!g130) & (!g460)) + ((!g76) & (sk[84]) & (g81) & (!g91) & (!g130) & (g460)) + ((!g76) & (sk[84]) & (g81) & (g91) & (!g130) & (!g460)) + ((!g76) & (sk[84]) & (g81) & (g91) & (!g130) & (g460)) + ((g76) & (!sk[84]) & (!g81) & (g91) & (!g130) & (g460)) + ((g76) & (!sk[84]) & (!g81) & (g91) & (g130) & (!g460)) + ((g76) & (!sk[84]) & (!g81) & (g91) & (g130) & (g460)) + ((g76) & (!sk[84]) & (g81) & (!g91) & (!g130) & (!g460)) + ((g76) & (!sk[84]) & (g81) & (!g91) & (!g130) & (g460)) + ((g76) & (!sk[84]) & (g81) & (!g91) & (g130) & (!g460)) + ((g76) & (!sk[84]) & (g81) & (!g91) & (g130) & (g460)) + ((g76) & (!sk[84]) & (g81) & (g91) & (!g130) & (!g460)) + ((g76) & (!sk[84]) & (g81) & (g91) & (!g130) & (g460)) + ((g76) & (!sk[84]) & (g81) & (g91) & (g130) & (!g460)) + ((g76) & (!sk[84]) & (g81) & (g91) & (g130) & (g460)) + ((g76) & (sk[84]) & (!g81) & (!g91) & (!g130) & (!g460)) + ((g76) & (sk[84]) & (g81) & (!g91) & (!g130) & (!g460)) + ((g76) & (sk[84]) & (g81) & (g91) & (!g130) & (!g460)));
	assign g567 = (((!g560) & (!g561) & (!g563) & (!g564) & (!g565) & (!g566)));
	assign g568 = (((!i_8_) & (!sk[86]) & (!g73) & (g76) & (!g88) & (g460)) + ((!i_8_) & (!sk[86]) & (!g73) & (g76) & (g88) & (!g460)) + ((!i_8_) & (!sk[86]) & (!g73) & (g76) & (g88) & (g460)) + ((!i_8_) & (!sk[86]) & (g73) & (!g76) & (!g88) & (!g460)) + ((!i_8_) & (!sk[86]) & (g73) & (!g76) & (!g88) & (g460)) + ((!i_8_) & (!sk[86]) & (g73) & (!g76) & (g88) & (!g460)) + ((!i_8_) & (!sk[86]) & (g73) & (!g76) & (g88) & (g460)) + ((!i_8_) & (!sk[86]) & (g73) & (g76) & (!g88) & (!g460)) + ((!i_8_) & (!sk[86]) & (g73) & (g76) & (!g88) & (g460)) + ((!i_8_) & (!sk[86]) & (g73) & (g76) & (g88) & (!g460)) + ((!i_8_) & (!sk[86]) & (g73) & (g76) & (g88) & (g460)) + ((i_8_) & (!sk[86]) & (!g73) & (g76) & (!g88) & (g460)) + ((i_8_) & (!sk[86]) & (!g73) & (g76) & (g88) & (!g460)) + ((i_8_) & (!sk[86]) & (!g73) & (g76) & (g88) & (g460)) + ((i_8_) & (!sk[86]) & (g73) & (!g76) & (!g88) & (!g460)) + ((i_8_) & (!sk[86]) & (g73) & (!g76) & (!g88) & (g460)) + ((i_8_) & (!sk[86]) & (g73) & (!g76) & (g88) & (!g460)) + ((i_8_) & (!sk[86]) & (g73) & (!g76) & (g88) & (g460)) + ((i_8_) & (!sk[86]) & (g73) & (g76) & (!g88) & (!g460)) + ((i_8_) & (!sk[86]) & (g73) & (g76) & (!g88) & (g460)) + ((i_8_) & (!sk[86]) & (g73) & (g76) & (g88) & (!g460)) + ((i_8_) & (!sk[86]) & (g73) & (g76) & (g88) & (g460)) + ((i_8_) & (sk[86]) & (g73) & (!g76) & (g88) & (!g460)) + ((i_8_) & (sk[86]) & (g73) & (!g76) & (g88) & (g460)) + ((i_8_) & (sk[86]) & (g73) & (g76) & (g88) & (!g460)));
	assign g569 = (((!g76) & (!sk[87]) & (!g161) & (g157) & (!g81) & (g88)) + ((!g76) & (!sk[87]) & (!g161) & (g157) & (g81) & (!g88)) + ((!g76) & (!sk[87]) & (!g161) & (g157) & (g81) & (g88)) + ((!g76) & (!sk[87]) & (g161) & (!g157) & (!g81) & (!g88)) + ((!g76) & (!sk[87]) & (g161) & (!g157) & (!g81) & (g88)) + ((!g76) & (!sk[87]) & (g161) & (!g157) & (g81) & (!g88)) + ((!g76) & (!sk[87]) & (g161) & (!g157) & (g81) & (g88)) + ((!g76) & (!sk[87]) & (g161) & (g157) & (!g81) & (!g88)) + ((!g76) & (!sk[87]) & (g161) & (g157) & (!g81) & (g88)) + ((!g76) & (!sk[87]) & (g161) & (g157) & (g81) & (!g88)) + ((!g76) & (!sk[87]) & (g161) & (g157) & (g81) & (g88)) + ((!g76) & (sk[87]) & (!g161) & (g157) & (!g81) & (g88)) + ((!g76) & (sk[87]) & (!g161) & (g157) & (g81) & (g88)) + ((!g76) & (sk[87]) & (g161) & (!g157) & (g81) & (!g88)) + ((!g76) & (sk[87]) & (g161) & (!g157) & (g81) & (g88)) + ((!g76) & (sk[87]) & (g161) & (g157) & (!g81) & (g88)) + ((!g76) & (sk[87]) & (g161) & (g157) & (g81) & (!g88)) + ((!g76) & (sk[87]) & (g161) & (g157) & (g81) & (g88)) + ((g76) & (!sk[87]) & (!g161) & (g157) & (!g81) & (g88)) + ((g76) & (!sk[87]) & (!g161) & (g157) & (g81) & (!g88)) + ((g76) & (!sk[87]) & (!g161) & (g157) & (g81) & (g88)) + ((g76) & (!sk[87]) & (g161) & (!g157) & (!g81) & (!g88)) + ((g76) & (!sk[87]) & (g161) & (!g157) & (!g81) & (g88)) + ((g76) & (!sk[87]) & (g161) & (!g157) & (g81) & (!g88)) + ((g76) & (!sk[87]) & (g161) & (!g157) & (g81) & (g88)) + ((g76) & (!sk[87]) & (g161) & (g157) & (!g81) & (!g88)) + ((g76) & (!sk[87]) & (g161) & (g157) & (!g81) & (g88)) + ((g76) & (!sk[87]) & (g161) & (g157) & (g81) & (!g88)) + ((g76) & (!sk[87]) & (g161) & (g157) & (g81) & (g88)));
	assign g570 = (((!i_10_) & (!sk[88]) & (!i_11_) & (i_15_) & (!g76)) + ((!i_10_) & (!sk[88]) & (!i_11_) & (i_15_) & (g76)) + ((!i_10_) & (!sk[88]) & (i_11_) & (i_15_) & (!g76)) + ((!i_10_) & (!sk[88]) & (i_11_) & (i_15_) & (g76)) + ((!i_10_) & (sk[88]) & (!i_11_) & (i_15_) & (!g76)) + ((i_10_) & (!sk[88]) & (!i_11_) & (i_15_) & (!g76)) + ((i_10_) & (!sk[88]) & (!i_11_) & (i_15_) & (g76)) + ((i_10_) & (!sk[88]) & (i_11_) & (i_15_) & (!g76)) + ((i_10_) & (!sk[88]) & (i_11_) & (i_15_) & (g76)));
	assign g571 = (((!sk[89]) & (!g123) & (!g213) & (g551) & (!g570)) + ((!sk[89]) & (!g123) & (!g213) & (g551) & (g570)) + ((!sk[89]) & (!g123) & (g213) & (g551) & (!g570)) + ((!sk[89]) & (!g123) & (g213) & (g551) & (g570)) + ((!sk[89]) & (g123) & (!g213) & (g551) & (!g570)) + ((!sk[89]) & (g123) & (!g213) & (g551) & (g570)) + ((!sk[89]) & (g123) & (g213) & (g551) & (!g570)) + ((!sk[89]) & (g123) & (g213) & (g551) & (g570)) + ((sk[89]) & (!g123) & (!g213) & (!g551) & (!g570)) + ((sk[89]) & (!g123) & (!g213) & (!g551) & (g570)) + ((sk[89]) & (!g123) & (g213) & (!g551) & (!g570)) + ((sk[89]) & (!g123) & (g213) & (!g551) & (g570)) + ((sk[89]) & (!g123) & (g213) & (g551) & (g570)) + ((sk[89]) & (g123) & (g213) & (!g551) & (g570)) + ((sk[89]) & (g123) & (g213) & (g551) & (g570)));
	assign g572 = (((!g17) & (!g76) & (g125) & (!sk[90]) & (!g81) & (g225)) + ((!g17) & (!g76) & (g125) & (!sk[90]) & (g81) & (!g225)) + ((!g17) & (!g76) & (g125) & (!sk[90]) & (g81) & (g225)) + ((!g17) & (!g76) & (g125) & (sk[90]) & (g81) & (!g225)) + ((!g17) & (!g76) & (g125) & (sk[90]) & (g81) & (g225)) + ((!g17) & (g76) & (!g125) & (!sk[90]) & (!g81) & (!g225)) + ((!g17) & (g76) & (!g125) & (!sk[90]) & (!g81) & (g225)) + ((!g17) & (g76) & (!g125) & (!sk[90]) & (g81) & (!g225)) + ((!g17) & (g76) & (!g125) & (!sk[90]) & (g81) & (g225)) + ((!g17) & (g76) & (g125) & (!sk[90]) & (!g81) & (!g225)) + ((!g17) & (g76) & (g125) & (!sk[90]) & (!g81) & (g225)) + ((!g17) & (g76) & (g125) & (!sk[90]) & (g81) & (!g225)) + ((!g17) & (g76) & (g125) & (!sk[90]) & (g81) & (g225)) + ((g17) & (!g76) & (!g125) & (sk[90]) & (!g81) & (g225)) + ((g17) & (!g76) & (!g125) & (sk[90]) & (g81) & (g225)) + ((g17) & (!g76) & (g125) & (!sk[90]) & (!g81) & (g225)) + ((g17) & (!g76) & (g125) & (!sk[90]) & (g81) & (!g225)) + ((g17) & (!g76) & (g125) & (!sk[90]) & (g81) & (g225)) + ((g17) & (!g76) & (g125) & (sk[90]) & (!g81) & (!g225)) + ((g17) & (!g76) & (g125) & (sk[90]) & (!g81) & (g225)) + ((g17) & (!g76) & (g125) & (sk[90]) & (g81) & (!g225)) + ((g17) & (!g76) & (g125) & (sk[90]) & (g81) & (g225)) + ((g17) & (g76) & (!g125) & (!sk[90]) & (!g81) & (!g225)) + ((g17) & (g76) & (!g125) & (!sk[90]) & (!g81) & (g225)) + ((g17) & (g76) & (!g125) & (!sk[90]) & (g81) & (!g225)) + ((g17) & (g76) & (!g125) & (!sk[90]) & (g81) & (g225)) + ((g17) & (g76) & (g125) & (!sk[90]) & (!g81) & (!g225)) + ((g17) & (g76) & (g125) & (!sk[90]) & (!g81) & (g225)) + ((g17) & (g76) & (g125) & (!sk[90]) & (g81) & (!g225)) + ((g17) & (g76) & (g125) & (!sk[90]) & (g81) & (g225)));
	assign g573 = (((!g135) & (!g131) & (!g562) & (sk[91]) & (!g557)) + ((!g135) & (!g131) & (g562) & (!sk[91]) & (!g557)) + ((!g135) & (!g131) & (g562) & (!sk[91]) & (g557)) + ((!g135) & (g131) & (!g562) & (sk[91]) & (!g557)) + ((!g135) & (g131) & (!g562) & (sk[91]) & (g557)) + ((!g135) & (g131) & (g562) & (!sk[91]) & (!g557)) + ((!g135) & (g131) & (g562) & (!sk[91]) & (g557)) + ((g135) & (!g131) & (!g562) & (sk[91]) & (!g557)) + ((g135) & (!g131) & (g562) & (!sk[91]) & (!g557)) + ((g135) & (!g131) & (g562) & (!sk[91]) & (g557)) + ((g135) & (g131) & (!g562) & (sk[91]) & (!g557)) + ((g135) & (g131) & (!g562) & (sk[91]) & (g557)) + ((g135) & (g131) & (g562) & (!sk[91]) & (!g557)) + ((g135) & (g131) & (g562) & (!sk[91]) & (g557)) + ((g135) & (g131) & (g562) & (sk[91]) & (!g557)) + ((g135) & (g131) & (g562) & (sk[91]) & (g557)));
	assign g574 = (((!i_8_) & (!g73) & (g76) & (!sk[92]) & (!g113) & (g460)) + ((!i_8_) & (!g73) & (g76) & (!sk[92]) & (g113) & (!g460)) + ((!i_8_) & (!g73) & (g76) & (!sk[92]) & (g113) & (g460)) + ((!i_8_) & (g73) & (!g76) & (!sk[92]) & (!g113) & (!g460)) + ((!i_8_) & (g73) & (!g76) & (!sk[92]) & (!g113) & (g460)) + ((!i_8_) & (g73) & (!g76) & (!sk[92]) & (g113) & (!g460)) + ((!i_8_) & (g73) & (!g76) & (!sk[92]) & (g113) & (g460)) + ((!i_8_) & (g73) & (!g76) & (sk[92]) & (!g113) & (!g460)) + ((!i_8_) & (g73) & (g76) & (!sk[92]) & (!g113) & (!g460)) + ((!i_8_) & (g73) & (g76) & (!sk[92]) & (!g113) & (g460)) + ((!i_8_) & (g73) & (g76) & (!sk[92]) & (g113) & (!g460)) + ((!i_8_) & (g73) & (g76) & (!sk[92]) & (g113) & (g460)) + ((!i_8_) & (g73) & (g76) & (sk[92]) & (!g113) & (!g460)) + ((i_8_) & (!g73) & (g76) & (!sk[92]) & (!g113) & (g460)) + ((i_8_) & (!g73) & (g76) & (!sk[92]) & (g113) & (!g460)) + ((i_8_) & (!g73) & (g76) & (!sk[92]) & (g113) & (g460)) + ((i_8_) & (g73) & (!g76) & (!sk[92]) & (!g113) & (!g460)) + ((i_8_) & (g73) & (!g76) & (!sk[92]) & (!g113) & (g460)) + ((i_8_) & (g73) & (!g76) & (!sk[92]) & (g113) & (!g460)) + ((i_8_) & (g73) & (!g76) & (!sk[92]) & (g113) & (g460)) + ((i_8_) & (g73) & (!g76) & (sk[92]) & (!g113) & (!g460)) + ((i_8_) & (g73) & (!g76) & (sk[92]) & (!g113) & (g460)) + ((i_8_) & (g73) & (g76) & (!sk[92]) & (!g113) & (!g460)) + ((i_8_) & (g73) & (g76) & (!sk[92]) & (!g113) & (g460)) + ((i_8_) & (g73) & (g76) & (!sk[92]) & (g113) & (!g460)) + ((i_8_) & (g73) & (g76) & (!sk[92]) & (g113) & (g460)) + ((i_8_) & (g73) & (g76) & (sk[92]) & (!g113) & (!g460)));
	assign g575 = (((!g568) & (!g569) & (!g571) & (!g572) & (g573) & (!g574)));
	assign g576 = (((!g17) & (!g36) & (!g76) & (sk[94]) & (g88) & (!g131)) + ((!g17) & (!g36) & (g76) & (!sk[94]) & (!g88) & (g131)) + ((!g17) & (!g36) & (g76) & (!sk[94]) & (g88) & (!g131)) + ((!g17) & (!g36) & (g76) & (!sk[94]) & (g88) & (g131)) + ((!g17) & (g36) & (!g76) & (!sk[94]) & (!g88) & (!g131)) + ((!g17) & (g36) & (!g76) & (!sk[94]) & (!g88) & (g131)) + ((!g17) & (g36) & (!g76) & (!sk[94]) & (g88) & (!g131)) + ((!g17) & (g36) & (!g76) & (!sk[94]) & (g88) & (g131)) + ((!g17) & (g36) & (!g76) & (sk[94]) & (!g88) & (!g131)) + ((!g17) & (g36) & (!g76) & (sk[94]) & (g88) & (!g131)) + ((!g17) & (g36) & (g76) & (!sk[94]) & (!g88) & (!g131)) + ((!g17) & (g36) & (g76) & (!sk[94]) & (!g88) & (g131)) + ((!g17) & (g36) & (g76) & (!sk[94]) & (g88) & (!g131)) + ((!g17) & (g36) & (g76) & (!sk[94]) & (g88) & (g131)) + ((g17) & (!g36) & (!g76) & (sk[94]) & (!g88) & (!g131)) + ((g17) & (!g36) & (!g76) & (sk[94]) & (g88) & (!g131)) + ((g17) & (!g36) & (g76) & (!sk[94]) & (!g88) & (g131)) + ((g17) & (!g36) & (g76) & (!sk[94]) & (g88) & (!g131)) + ((g17) & (!g36) & (g76) & (!sk[94]) & (g88) & (g131)) + ((g17) & (g36) & (!g76) & (!sk[94]) & (!g88) & (!g131)) + ((g17) & (g36) & (!g76) & (!sk[94]) & (!g88) & (g131)) + ((g17) & (g36) & (!g76) & (!sk[94]) & (g88) & (!g131)) + ((g17) & (g36) & (!g76) & (!sk[94]) & (g88) & (g131)) + ((g17) & (g36) & (!g76) & (sk[94]) & (!g88) & (!g131)) + ((g17) & (g36) & (!g76) & (sk[94]) & (g88) & (!g131)) + ((g17) & (g36) & (g76) & (!sk[94]) & (!g88) & (!g131)) + ((g17) & (g36) & (g76) & (!sk[94]) & (!g88) & (g131)) + ((g17) & (g36) & (g76) & (!sk[94]) & (g88) & (!g131)) + ((g17) & (g36) & (g76) & (!sk[94]) & (g88) & (g131)));
	assign g577 = (((!g125) & (!g131) & (!sk[95]) & (g551) & (!g543)) + ((!g125) & (!g131) & (!sk[95]) & (g551) & (g543)) + ((!g125) & (!g131) & (sk[95]) & (g551) & (!g543)) + ((!g125) & (g131) & (!sk[95]) & (g551) & (!g543)) + ((!g125) & (g131) & (!sk[95]) & (g551) & (g543)) + ((!g125) & (g131) & (sk[95]) & (!g551) & (!g543)) + ((!g125) & (g131) & (sk[95]) & (!g551) & (g543)) + ((!g125) & (g131) & (sk[95]) & (g551) & (!g543)) + ((!g125) & (g131) & (sk[95]) & (g551) & (g543)) + ((g125) & (!g131) & (!sk[95]) & (g551) & (!g543)) + ((g125) & (!g131) & (!sk[95]) & (g551) & (g543)) + ((g125) & (!g131) & (sk[95]) & (g551) & (!g543)) + ((g125) & (g131) & (!sk[95]) & (g551) & (!g543)) + ((g125) & (g131) & (!sk[95]) & (g551) & (g543)) + ((g125) & (g131) & (sk[95]) & (g551) & (!g543)) + ((g125) & (g131) & (sk[95]) & (g551) & (g543)));
	assign g578 = (((g17) & (!sk[96]) & (!g460)) + ((g17) & (!sk[96]) & (g460)) + ((g17) & (sk[96]) & (!g460)));
	assign g579 = (((!g102) & (!sk[97]) & (!g105) & (g578) & (!g495)) + ((!g102) & (!sk[97]) & (!g105) & (g578) & (g495)) + ((!g102) & (!sk[97]) & (g105) & (g578) & (!g495)) + ((!g102) & (!sk[97]) & (g105) & (g578) & (g495)) + ((!g102) & (sk[97]) & (!g105) & (!g578) & (g495)) + ((!g102) & (sk[97]) & (!g105) & (g578) & (g495)) + ((g102) & (!sk[97]) & (!g105) & (g578) & (!g495)) + ((g102) & (!sk[97]) & (!g105) & (g578) & (g495)) + ((g102) & (!sk[97]) & (g105) & (g578) & (!g495)) + ((g102) & (!sk[97]) & (g105) & (g578) & (g495)) + ((g102) & (sk[97]) & (!g105) & (!g578) & (g495)) + ((g102) & (sk[97]) & (!g105) & (g578) & (!g495)) + ((g102) & (sk[97]) & (!g105) & (g578) & (g495)) + ((g102) & (sk[97]) & (g105) & (g578) & (!g495)) + ((g102) & (sk[97]) & (g105) & (g578) & (g495)));
	assign g580 = (((!i_15_) & (!g151) & (!g460) & (!g576) & (g577) & (!g579)) + ((!i_15_) & (!g151) & (g460) & (!g576) & (g577) & (!g579)) + ((!i_15_) & (g151) & (!g460) & (!g576) & (g577) & (!g579)) + ((!i_15_) & (g151) & (g460) & (!g576) & (g577) & (!g579)) + ((i_15_) & (!g151) & (!g460) & (!g576) & (g577) & (!g579)) + ((i_15_) & (!g151) & (g460) & (!g576) & (g577) & (!g579)) + ((i_15_) & (g151) & (g460) & (!g576) & (g577) & (!g579)));
	assign g581 = (((g1554) & (g1543) & (g559) & (g567) & (g575) & (g580)));
	assign g582 = (((!i_12_) & (!sk[100]) & (!i_13_) & (i_14_) & (!g75) & (g81)) + ((!i_12_) & (!sk[100]) & (!i_13_) & (i_14_) & (g75) & (!g81)) + ((!i_12_) & (!sk[100]) & (!i_13_) & (i_14_) & (g75) & (g81)) + ((!i_12_) & (!sk[100]) & (i_13_) & (!i_14_) & (!g75) & (!g81)) + ((!i_12_) & (!sk[100]) & (i_13_) & (!i_14_) & (!g75) & (g81)) + ((!i_12_) & (!sk[100]) & (i_13_) & (!i_14_) & (g75) & (!g81)) + ((!i_12_) & (!sk[100]) & (i_13_) & (!i_14_) & (g75) & (g81)) + ((!i_12_) & (!sk[100]) & (i_13_) & (i_14_) & (!g75) & (!g81)) + ((!i_12_) & (!sk[100]) & (i_13_) & (i_14_) & (!g75) & (g81)) + ((!i_12_) & (!sk[100]) & (i_13_) & (i_14_) & (g75) & (!g81)) + ((!i_12_) & (!sk[100]) & (i_13_) & (i_14_) & (g75) & (g81)) + ((!i_12_) & (sk[100]) & (i_13_) & (i_14_) & (!g75) & (g81)) + ((i_12_) & (!sk[100]) & (!i_13_) & (i_14_) & (!g75) & (g81)) + ((i_12_) & (!sk[100]) & (!i_13_) & (i_14_) & (g75) & (!g81)) + ((i_12_) & (!sk[100]) & (!i_13_) & (i_14_) & (g75) & (g81)) + ((i_12_) & (!sk[100]) & (i_13_) & (!i_14_) & (!g75) & (!g81)) + ((i_12_) & (!sk[100]) & (i_13_) & (!i_14_) & (!g75) & (g81)) + ((i_12_) & (!sk[100]) & (i_13_) & (!i_14_) & (g75) & (!g81)) + ((i_12_) & (!sk[100]) & (i_13_) & (!i_14_) & (g75) & (g81)) + ((i_12_) & (!sk[100]) & (i_13_) & (i_14_) & (!g75) & (!g81)) + ((i_12_) & (!sk[100]) & (i_13_) & (i_14_) & (!g75) & (g81)) + ((i_12_) & (!sk[100]) & (i_13_) & (i_14_) & (g75) & (!g81)) + ((i_12_) & (!sk[100]) & (i_13_) & (i_14_) & (g75) & (g81)) + ((i_12_) & (sk[100]) & (i_13_) & (!i_14_) & (!g75) & (g81)));
	assign g583 = (((!sk[101]) & (!i_8_) & (!g73) & (g501) & (!g543)) + ((!sk[101]) & (!i_8_) & (!g73) & (g501) & (g543)) + ((!sk[101]) & (!i_8_) & (g73) & (g501) & (!g543)) + ((!sk[101]) & (!i_8_) & (g73) & (g501) & (g543)) + ((!sk[101]) & (i_8_) & (!g73) & (g501) & (!g543)) + ((!sk[101]) & (i_8_) & (!g73) & (g501) & (g543)) + ((!sk[101]) & (i_8_) & (g73) & (g501) & (!g543)) + ((!sk[101]) & (i_8_) & (g73) & (g501) & (g543)) + ((sk[101]) & (!i_8_) & (g73) & (!g501) & (g543)) + ((sk[101]) & (!i_8_) & (g73) & (g501) & (!g543)) + ((sk[101]) & (!i_8_) & (g73) & (g501) & (g543)));
	assign g584 = (((!i_8_) & (!sk[102]) & (!g73) & (g76) & (!g88) & (g460)) + ((!i_8_) & (!sk[102]) & (!g73) & (g76) & (g88) & (!g460)) + ((!i_8_) & (!sk[102]) & (!g73) & (g76) & (g88) & (g460)) + ((!i_8_) & (!sk[102]) & (g73) & (!g76) & (!g88) & (!g460)) + ((!i_8_) & (!sk[102]) & (g73) & (!g76) & (!g88) & (g460)) + ((!i_8_) & (!sk[102]) & (g73) & (!g76) & (g88) & (!g460)) + ((!i_8_) & (!sk[102]) & (g73) & (!g76) & (g88) & (g460)) + ((!i_8_) & (!sk[102]) & (g73) & (g76) & (!g88) & (!g460)) + ((!i_8_) & (!sk[102]) & (g73) & (g76) & (!g88) & (g460)) + ((!i_8_) & (!sk[102]) & (g73) & (g76) & (g88) & (!g460)) + ((!i_8_) & (!sk[102]) & (g73) & (g76) & (g88) & (g460)) + ((!i_8_) & (sk[102]) & (g73) & (!g76) & (g88) & (!g460)) + ((!i_8_) & (sk[102]) & (g73) & (!g76) & (g88) & (g460)) + ((!i_8_) & (sk[102]) & (g73) & (g76) & (g88) & (!g460)) + ((i_8_) & (!sk[102]) & (!g73) & (g76) & (!g88) & (g460)) + ((i_8_) & (!sk[102]) & (!g73) & (g76) & (g88) & (!g460)) + ((i_8_) & (!sk[102]) & (!g73) & (g76) & (g88) & (g460)) + ((i_8_) & (!sk[102]) & (g73) & (!g76) & (!g88) & (!g460)) + ((i_8_) & (!sk[102]) & (g73) & (!g76) & (!g88) & (g460)) + ((i_8_) & (!sk[102]) & (g73) & (!g76) & (g88) & (!g460)) + ((i_8_) & (!sk[102]) & (g73) & (!g76) & (g88) & (g460)) + ((i_8_) & (!sk[102]) & (g73) & (g76) & (!g88) & (!g460)) + ((i_8_) & (!sk[102]) & (g73) & (g76) & (!g88) & (g460)) + ((i_8_) & (!sk[102]) & (g73) & (g76) & (g88) & (!g460)) + ((i_8_) & (!sk[102]) & (g73) & (g76) & (g88) & (g460)));
	assign g585 = (((!i_8_) & (!g73) & (g552) & (!sk[103]) & (!g511)) + ((!i_8_) & (!g73) & (g552) & (!sk[103]) & (g511)) + ((!i_8_) & (g73) & (g552) & (!sk[103]) & (!g511)) + ((!i_8_) & (g73) & (g552) & (!sk[103]) & (g511)) + ((i_8_) & (!g73) & (g552) & (!sk[103]) & (!g511)) + ((i_8_) & (!g73) & (g552) & (!sk[103]) & (g511)) + ((i_8_) & (g73) & (!g552) & (sk[103]) & (!g511)) + ((i_8_) & (g73) & (!g552) & (sk[103]) & (g511)) + ((i_8_) & (g73) & (g552) & (!sk[103]) & (!g511)) + ((i_8_) & (g73) & (g552) & (!sk[103]) & (g511)) + ((i_8_) & (g73) & (g552) & (sk[103]) & (g511)));
	assign g586 = (((!i_8_) & (!g73) & (g551) & (!sk[104]) & (!g578) & (g495)) + ((!i_8_) & (!g73) & (g551) & (!sk[104]) & (g578) & (!g495)) + ((!i_8_) & (!g73) & (g551) & (!sk[104]) & (g578) & (g495)) + ((!i_8_) & (g73) & (!g551) & (!sk[104]) & (!g578) & (!g495)) + ((!i_8_) & (g73) & (!g551) & (!sk[104]) & (!g578) & (g495)) + ((!i_8_) & (g73) & (!g551) & (!sk[104]) & (g578) & (!g495)) + ((!i_8_) & (g73) & (!g551) & (!sk[104]) & (g578) & (g495)) + ((!i_8_) & (g73) & (!g551) & (sk[104]) & (!g578) & (g495)) + ((!i_8_) & (g73) & (!g551) & (sk[104]) & (g578) & (!g495)) + ((!i_8_) & (g73) & (!g551) & (sk[104]) & (g578) & (g495)) + ((!i_8_) & (g73) & (g551) & (!sk[104]) & (!g578) & (!g495)) + ((!i_8_) & (g73) & (g551) & (!sk[104]) & (!g578) & (g495)) + ((!i_8_) & (g73) & (g551) & (!sk[104]) & (g578) & (!g495)) + ((!i_8_) & (g73) & (g551) & (!sk[104]) & (g578) & (g495)) + ((!i_8_) & (g73) & (g551) & (sk[104]) & (!g578) & (g495)) + ((!i_8_) & (g73) & (g551) & (sk[104]) & (g578) & (!g495)) + ((!i_8_) & (g73) & (g551) & (sk[104]) & (g578) & (g495)) + ((i_8_) & (!g73) & (g551) & (!sk[104]) & (!g578) & (g495)) + ((i_8_) & (!g73) & (g551) & (!sk[104]) & (g578) & (!g495)) + ((i_8_) & (!g73) & (g551) & (!sk[104]) & (g578) & (g495)) + ((i_8_) & (g73) & (!g551) & (!sk[104]) & (!g578) & (!g495)) + ((i_8_) & (g73) & (!g551) & (!sk[104]) & (!g578) & (g495)) + ((i_8_) & (g73) & (!g551) & (!sk[104]) & (g578) & (!g495)) + ((i_8_) & (g73) & (!g551) & (!sk[104]) & (g578) & (g495)) + ((i_8_) & (g73) & (!g551) & (sk[104]) & (!g578) & (!g495)) + ((i_8_) & (g73) & (!g551) & (sk[104]) & (!g578) & (g495)) + ((i_8_) & (g73) & (!g551) & (sk[104]) & (g578) & (!g495)) + ((i_8_) & (g73) & (!g551) & (sk[104]) & (g578) & (g495)) + ((i_8_) & (g73) & (g551) & (!sk[104]) & (!g578) & (!g495)) + ((i_8_) & (g73) & (g551) & (!sk[104]) & (!g578) & (g495)) + ((i_8_) & (g73) & (g551) & (!sk[104]) & (g578) & (!g495)) + ((i_8_) & (g73) & (g551) & (!sk[104]) & (g578) & (g495)) + ((i_8_) & (g73) & (g551) & (sk[104]) & (!g578) & (g495)) + ((i_8_) & (g73) & (g551) & (sk[104]) & (g578) & (!g495)) + ((i_8_) & (g73) & (g551) & (sk[104]) & (g578) & (g495)));
	assign g587 = (((!g74) & (!g513) & (!g583) & (!g584) & (!g585) & (!g586)) + ((!g74) & (g513) & (!g583) & (!g584) & (!g585) & (!g586)) + ((g74) & (g513) & (!g583) & (!g584) & (!g585) & (!g586)));
	assign g588 = (((!i_8_) & (!sk[106]) & (!g17) & (g73) & (!g76) & (g511)) + ((!i_8_) & (!sk[106]) & (!g17) & (g73) & (g76) & (!g511)) + ((!i_8_) & (!sk[106]) & (!g17) & (g73) & (g76) & (g511)) + ((!i_8_) & (!sk[106]) & (g17) & (!g73) & (!g76) & (!g511)) + ((!i_8_) & (!sk[106]) & (g17) & (!g73) & (!g76) & (g511)) + ((!i_8_) & (!sk[106]) & (g17) & (!g73) & (g76) & (!g511)) + ((!i_8_) & (!sk[106]) & (g17) & (!g73) & (g76) & (g511)) + ((!i_8_) & (!sk[106]) & (g17) & (g73) & (!g76) & (!g511)) + ((!i_8_) & (!sk[106]) & (g17) & (g73) & (!g76) & (g511)) + ((!i_8_) & (!sk[106]) & (g17) & (g73) & (g76) & (!g511)) + ((!i_8_) & (!sk[106]) & (g17) & (g73) & (g76) & (g511)) + ((!i_8_) & (sk[106]) & (!g17) & (g73) & (!g76) & (g511)) + ((!i_8_) & (sk[106]) & (!g17) & (g73) & (g76) & (g511)) + ((!i_8_) & (sk[106]) & (g17) & (g73) & (!g76) & (!g511)) + ((!i_8_) & (sk[106]) & (g17) & (g73) & (!g76) & (g511)) + ((!i_8_) & (sk[106]) & (g17) & (g73) & (g76) & (g511)) + ((i_8_) & (!sk[106]) & (!g17) & (g73) & (!g76) & (g511)) + ((i_8_) & (!sk[106]) & (!g17) & (g73) & (g76) & (!g511)) + ((i_8_) & (!sk[106]) & (!g17) & (g73) & (g76) & (g511)) + ((i_8_) & (!sk[106]) & (g17) & (!g73) & (!g76) & (!g511)) + ((i_8_) & (!sk[106]) & (g17) & (!g73) & (!g76) & (g511)) + ((i_8_) & (!sk[106]) & (g17) & (!g73) & (g76) & (!g511)) + ((i_8_) & (!sk[106]) & (g17) & (!g73) & (g76) & (g511)) + ((i_8_) & (!sk[106]) & (g17) & (g73) & (!g76) & (!g511)) + ((i_8_) & (!sk[106]) & (g17) & (g73) & (!g76) & (g511)) + ((i_8_) & (!sk[106]) & (g17) & (g73) & (g76) & (!g511)) + ((i_8_) & (!sk[106]) & (g17) & (g73) & (g76) & (g511)) + ((i_8_) & (sk[106]) & (g17) & (g73) & (!g76) & (!g511)) + ((i_8_) & (sk[106]) & (g17) & (g73) & (!g76) & (g511)));
	assign g589 = (((!g582) & (!g587) & (!sk[107]) & (g588)) + ((!g582) & (g587) & (!sk[107]) & (!g588)) + ((!g582) & (g587) & (!sk[107]) & (g588)) + ((!g582) & (g587) & (sk[107]) & (!g588)) + ((g582) & (!g587) & (!sk[107]) & (g588)) + ((g582) & (g587) & (!sk[107]) & (!g588)) + ((g582) & (g587) & (!sk[107]) & (g588)));
	assign g590 = (((!g74) & (!sk[108]) & (!g259) & (g552)) + ((!g74) & (!sk[108]) & (g259) & (!g552)) + ((!g74) & (!sk[108]) & (g259) & (g552)) + ((!g74) & (sk[108]) & (!g259) & (!g552)) + ((g74) & (!sk[108]) & (!g259) & (g552)) + ((g74) & (!sk[108]) & (g259) & (!g552)) + ((g74) & (!sk[108]) & (g259) & (g552)) + ((g74) & (sk[108]) & (!g259) & (!g552)) + ((g74) & (sk[108]) & (g259) & (!g552)));
	assign g591 = (((!g125) & (!g168) & (!sk[109]) & (g511)) + ((!g125) & (g168) & (!sk[109]) & (!g511)) + ((!g125) & (g168) & (!sk[109]) & (g511)) + ((!g125) & (g168) & (sk[109]) & (g511)) + ((g125) & (!g168) & (!sk[109]) & (g511)) + ((g125) & (!g168) & (sk[109]) & (g511)) + ((g125) & (g168) & (!sk[109]) & (!g511)) + ((g125) & (g168) & (!sk[109]) & (g511)) + ((g125) & (g168) & (sk[109]) & (g511)));
	assign g592 = (((!i_8_) & (!g73) & (!g155) & (!g555) & (!g486) & (!g591)) + ((!i_8_) & (!g73) & (g155) & (!g555) & (!g486) & (!g591)) + ((!i_8_) & (!g73) & (g155) & (!g555) & (g486) & (!g591)) + ((!i_8_) & (!g73) & (g155) & (g555) & (!g486) & (!g591)) + ((!i_8_) & (!g73) & (g155) & (g555) & (g486) & (!g591)) + ((!i_8_) & (g73) & (!g155) & (!g555) & (!g486) & (!g591)) + ((!i_8_) & (g73) & (g155) & (!g555) & (!g486) & (!g591)) + ((!i_8_) & (g73) & (g155) & (!g555) & (g486) & (!g591)) + ((i_8_) & (!g73) & (!g155) & (!g555) & (!g486) & (!g591)) + ((i_8_) & (!g73) & (g155) & (!g555) & (!g486) & (!g591)) + ((i_8_) & (!g73) & (g155) & (!g555) & (g486) & (!g591)) + ((i_8_) & (!g73) & (g155) & (g555) & (!g486) & (!g591)) + ((i_8_) & (!g73) & (g155) & (g555) & (g486) & (!g591)) + ((i_8_) & (g73) & (!g155) & (!g555) & (!g486) & (!g591)) + ((i_8_) & (g73) & (g155) & (!g555) & (!g486) & (!g591)));
	assign g593 = (((!g157) & (!g262) & (!g258) & (g551) & (!g562) & (!g501)) + ((!g157) & (!g262) & (!g258) & (g551) & (!g562) & (g501)) + ((!g157) & (!g262) & (!g258) & (g551) & (g562) & (!g501)) + ((!g157) & (!g262) & (!g258) & (g551) & (g562) & (g501)) + ((!g157) & (!g262) & (g258) & (!g551) & (!g562) & (!g501)) + ((!g157) & (!g262) & (g258) & (!g551) & (!g562) & (g501)) + ((!g157) & (!g262) & (g258) & (!g551) & (g562) & (!g501)) + ((!g157) & (!g262) & (g258) & (!g551) & (g562) & (g501)) + ((!g157) & (!g262) & (g258) & (g551) & (!g562) & (!g501)) + ((!g157) & (!g262) & (g258) & (g551) & (!g562) & (g501)) + ((!g157) & (!g262) & (g258) & (g551) & (g562) & (!g501)) + ((!g157) & (!g262) & (g258) & (g551) & (g562) & (g501)) + ((!g157) & (g262) & (!g258) & (g551) & (!g562) & (!g501)) + ((!g157) & (g262) & (!g258) & (g551) & (!g562) & (g501)) + ((!g157) & (g262) & (g258) & (!g551) & (!g562) & (!g501)) + ((!g157) & (g262) & (g258) & (!g551) & (!g562) & (g501)) + ((!g157) & (g262) & (g258) & (g551) & (!g562) & (!g501)) + ((!g157) & (g262) & (g258) & (g551) & (!g562) & (g501)) + ((g157) & (!g262) & (!g258) & (g551) & (!g562) & (!g501)) + ((g157) & (!g262) & (!g258) & (g551) & (g562) & (!g501)) + ((g157) & (!g262) & (g258) & (!g551) & (!g562) & (!g501)) + ((g157) & (!g262) & (g258) & (!g551) & (g562) & (!g501)) + ((g157) & (!g262) & (g258) & (g551) & (!g562) & (!g501)) + ((g157) & (!g262) & (g258) & (g551) & (g562) & (!g501)) + ((g157) & (g262) & (!g258) & (g551) & (!g562) & (!g501)) + ((g157) & (g262) & (g258) & (!g551) & (!g562) & (!g501)) + ((g157) & (g262) & (g258) & (g551) & (!g562) & (!g501)));
	assign g594 = (((!g157) & (!g135) & (!sk[112]) & (g253) & (!g254)) + ((!g157) & (!g135) & (!sk[112]) & (g253) & (g254)) + ((!g157) & (g135) & (!sk[112]) & (g253) & (!g254)) + ((!g157) & (g135) & (!sk[112]) & (g253) & (g254)) + ((!g157) & (g135) & (sk[112]) & (g253) & (g254)) + ((g157) & (!g135) & (!sk[112]) & (g253) & (!g254)) + ((g157) & (!g135) & (!sk[112]) & (g253) & (g254)) + ((g157) & (g135) & (!sk[112]) & (g253) & (!g254)) + ((g157) & (g135) & (!sk[112]) & (g253) & (g254)));
	assign g595 = (((!sk[113]) & (!g258) & (!g431) & (g543) & (!g557) & (g594)) + ((!sk[113]) & (!g258) & (!g431) & (g543) & (g557) & (!g594)) + ((!sk[113]) & (!g258) & (!g431) & (g543) & (g557) & (g594)) + ((!sk[113]) & (!g258) & (g431) & (!g543) & (!g557) & (!g594)) + ((!sk[113]) & (!g258) & (g431) & (!g543) & (!g557) & (g594)) + ((!sk[113]) & (!g258) & (g431) & (!g543) & (g557) & (!g594)) + ((!sk[113]) & (!g258) & (g431) & (!g543) & (g557) & (g594)) + ((!sk[113]) & (!g258) & (g431) & (g543) & (!g557) & (!g594)) + ((!sk[113]) & (!g258) & (g431) & (g543) & (!g557) & (g594)) + ((!sk[113]) & (!g258) & (g431) & (g543) & (g557) & (!g594)) + ((!sk[113]) & (!g258) & (g431) & (g543) & (g557) & (g594)) + ((!sk[113]) & (g258) & (!g431) & (g543) & (!g557) & (g594)) + ((!sk[113]) & (g258) & (!g431) & (g543) & (g557) & (!g594)) + ((!sk[113]) & (g258) & (!g431) & (g543) & (g557) & (g594)) + ((!sk[113]) & (g258) & (g431) & (!g543) & (!g557) & (!g594)) + ((!sk[113]) & (g258) & (g431) & (!g543) & (!g557) & (g594)) + ((!sk[113]) & (g258) & (g431) & (!g543) & (g557) & (!g594)) + ((!sk[113]) & (g258) & (g431) & (!g543) & (g557) & (g594)) + ((!sk[113]) & (g258) & (g431) & (g543) & (!g557) & (!g594)) + ((!sk[113]) & (g258) & (g431) & (g543) & (!g557) & (g594)) + ((!sk[113]) & (g258) & (g431) & (g543) & (g557) & (!g594)) + ((!sk[113]) & (g258) & (g431) & (g543) & (g557) & (g594)) + ((sk[113]) & (!g258) & (!g431) & (!g543) & (!g557) & (!g594)) + ((sk[113]) & (!g258) & (!g431) & (!g543) & (!g557) & (g594)) + ((sk[113]) & (!g258) & (!g431) & (g543) & (!g557) & (g594)) + ((sk[113]) & (!g258) & (g431) & (!g543) & (!g557) & (!g594)) + ((sk[113]) & (!g258) & (g431) & (!g543) & (!g557) & (g594)) + ((sk[113]) & (!g258) & (g431) & (g543) & (!g557) & (g594)) + ((sk[113]) & (g258) & (!g431) & (!g543) & (!g557) & (!g594)) + ((sk[113]) & (g258) & (!g431) & (!g543) & (!g557) & (g594)) + ((sk[113]) & (g258) & (!g431) & (!g543) & (g557) & (!g594)) + ((sk[113]) & (g258) & (!g431) & (!g543) & (g557) & (g594)) + ((sk[113]) & (g258) & (!g431) & (g543) & (!g557) & (g594)) + ((sk[113]) & (g258) & (!g431) & (g543) & (g557) & (g594)) + ((sk[113]) & (g258) & (g431) & (!g543) & (!g557) & (!g594)) + ((sk[113]) & (g258) & (g431) & (!g543) & (!g557) & (g594)) + ((sk[113]) & (g258) & (g431) & (g543) & (!g557) & (g594)));
	assign g596 = (((!g167) & (!g578) & (!g590) & (g592) & (g593) & (g595)) + ((!g167) & (g578) & (!g590) & (g592) & (g593) & (g595)) + ((g167) & (!g578) & (!g590) & (g592) & (g593) & (g595)));
	assign g597 = (((g81) & (!sk[115]) & (!g482)) + ((g81) & (!sk[115]) & (g482)) + ((g81) & (sk[115]) & (g482)));
	assign g598 = (((!g159) & (!g521) & (!sk[116]) & (g597) & (!g483) & (g489)) + ((!g159) & (!g521) & (!sk[116]) & (g597) & (g483) & (!g489)) + ((!g159) & (!g521) & (!sk[116]) & (g597) & (g483) & (g489)) + ((!g159) & (!g521) & (sk[116]) & (!g597) & (!g483) & (g489)) + ((!g159) & (!g521) & (sk[116]) & (!g597) & (g483) & (!g489)) + ((!g159) & (!g521) & (sk[116]) & (!g597) & (g483) & (g489)) + ((!g159) & (!g521) & (sk[116]) & (g597) & (!g483) & (!g489)) + ((!g159) & (!g521) & (sk[116]) & (g597) & (!g483) & (g489)) + ((!g159) & (!g521) & (sk[116]) & (g597) & (g483) & (!g489)) + ((!g159) & (!g521) & (sk[116]) & (g597) & (g483) & (g489)) + ((!g159) & (g521) & (!sk[116]) & (!g597) & (!g483) & (!g489)) + ((!g159) & (g521) & (!sk[116]) & (!g597) & (!g483) & (g489)) + ((!g159) & (g521) & (!sk[116]) & (!g597) & (g483) & (!g489)) + ((!g159) & (g521) & (!sk[116]) & (!g597) & (g483) & (g489)) + ((!g159) & (g521) & (!sk[116]) & (g597) & (!g483) & (!g489)) + ((!g159) & (g521) & (!sk[116]) & (g597) & (!g483) & (g489)) + ((!g159) & (g521) & (!sk[116]) & (g597) & (g483) & (!g489)) + ((!g159) & (g521) & (!sk[116]) & (g597) & (g483) & (g489)) + ((!g159) & (g521) & (sk[116]) & (!g597) & (!g483) & (!g489)) + ((!g159) & (g521) & (sk[116]) & (!g597) & (!g483) & (g489)) + ((!g159) & (g521) & (sk[116]) & (!g597) & (g483) & (!g489)) + ((!g159) & (g521) & (sk[116]) & (!g597) & (g483) & (g489)) + ((!g159) & (g521) & (sk[116]) & (g597) & (!g483) & (!g489)) + ((!g159) & (g521) & (sk[116]) & (g597) & (!g483) & (g489)) + ((!g159) & (g521) & (sk[116]) & (g597) & (g483) & (!g489)) + ((!g159) & (g521) & (sk[116]) & (g597) & (g483) & (g489)) + ((g159) & (!g521) & (!sk[116]) & (g597) & (!g483) & (g489)) + ((g159) & (!g521) & (!sk[116]) & (g597) & (g483) & (!g489)) + ((g159) & (!g521) & (!sk[116]) & (g597) & (g483) & (g489)) + ((g159) & (g521) & (!sk[116]) & (!g597) & (!g483) & (!g489)) + ((g159) & (g521) & (!sk[116]) & (!g597) & (!g483) & (g489)) + ((g159) & (g521) & (!sk[116]) & (!g597) & (g483) & (!g489)) + ((g159) & (g521) & (!sk[116]) & (!g597) & (g483) & (g489)) + ((g159) & (g521) & (!sk[116]) & (g597) & (!g483) & (!g489)) + ((g159) & (g521) & (!sk[116]) & (g597) & (!g483) & (g489)) + ((g159) & (g521) & (!sk[116]) & (g597) & (g483) & (!g489)) + ((g159) & (g521) & (!sk[116]) & (g597) & (g483) & (g489)));
	assign g599 = (((!g159) & (!g154) & (!g500) & (sk[117]) & (!g522) & (!g598)) + ((!g159) & (!g154) & (g500) & (!sk[117]) & (!g522) & (g598)) + ((!g159) & (!g154) & (g500) & (!sk[117]) & (g522) & (!g598)) + ((!g159) & (!g154) & (g500) & (!sk[117]) & (g522) & (g598)) + ((!g159) & (g154) & (!g500) & (!sk[117]) & (!g522) & (!g598)) + ((!g159) & (g154) & (!g500) & (!sk[117]) & (!g522) & (g598)) + ((!g159) & (g154) & (!g500) & (!sk[117]) & (g522) & (!g598)) + ((!g159) & (g154) & (!g500) & (!sk[117]) & (g522) & (g598)) + ((!g159) & (g154) & (!g500) & (sk[117]) & (!g522) & (!g598)) + ((!g159) & (g154) & (!g500) & (sk[117]) & (g522) & (!g598)) + ((!g159) & (g154) & (g500) & (!sk[117]) & (!g522) & (!g598)) + ((!g159) & (g154) & (g500) & (!sk[117]) & (!g522) & (g598)) + ((!g159) & (g154) & (g500) & (!sk[117]) & (g522) & (!g598)) + ((!g159) & (g154) & (g500) & (!sk[117]) & (g522) & (g598)) + ((g159) & (!g154) & (!g500) & (sk[117]) & (!g522) & (!g598)) + ((g159) & (!g154) & (g500) & (!sk[117]) & (!g522) & (g598)) + ((g159) & (!g154) & (g500) & (!sk[117]) & (g522) & (!g598)) + ((g159) & (!g154) & (g500) & (!sk[117]) & (g522) & (g598)) + ((g159) & (g154) & (!g500) & (!sk[117]) & (!g522) & (!g598)) + ((g159) & (g154) & (!g500) & (!sk[117]) & (!g522) & (g598)) + ((g159) & (g154) & (!g500) & (!sk[117]) & (g522) & (!g598)) + ((g159) & (g154) & (!g500) & (!sk[117]) & (g522) & (g598)) + ((g159) & (g154) & (!g500) & (sk[117]) & (!g522) & (!g598)) + ((g159) & (g154) & (!g500) & (sk[117]) & (g522) & (!g598)) + ((g159) & (g154) & (g500) & (!sk[117]) & (!g522) & (!g598)) + ((g159) & (g154) & (g500) & (!sk[117]) & (!g522) & (g598)) + ((g159) & (g154) & (g500) & (!sk[117]) & (g522) & (!g598)) + ((g159) & (g154) & (g500) & (!sk[117]) & (g522) & (g598)) + ((g159) & (g154) & (g500) & (sk[117]) & (!g522) & (!g598)) + ((g159) & (g154) & (g500) & (sk[117]) & (g522) & (!g598)));
	assign g600 = (((!g154) & (!g521) & (!g597) & (!g489) & (sk[118]) & (g599)) + ((!g154) & (!g521) & (g597) & (!g489) & (!sk[118]) & (g599)) + ((!g154) & (!g521) & (g597) & (g489) & (!sk[118]) & (!g599)) + ((!g154) & (!g521) & (g597) & (g489) & (!sk[118]) & (g599)) + ((!g154) & (g521) & (!g597) & (!g489) & (!sk[118]) & (!g599)) + ((!g154) & (g521) & (!g597) & (!g489) & (!sk[118]) & (g599)) + ((!g154) & (g521) & (!g597) & (g489) & (!sk[118]) & (!g599)) + ((!g154) & (g521) & (!g597) & (g489) & (!sk[118]) & (g599)) + ((!g154) & (g521) & (g597) & (!g489) & (!sk[118]) & (!g599)) + ((!g154) & (g521) & (g597) & (!g489) & (!sk[118]) & (g599)) + ((!g154) & (g521) & (g597) & (g489) & (!sk[118]) & (!g599)) + ((!g154) & (g521) & (g597) & (g489) & (!sk[118]) & (g599)) + ((g154) & (!g521) & (!g597) & (!g489) & (sk[118]) & (g599)) + ((g154) & (!g521) & (!g597) & (g489) & (sk[118]) & (g599)) + ((g154) & (!g521) & (g597) & (!g489) & (!sk[118]) & (g599)) + ((g154) & (!g521) & (g597) & (!g489) & (sk[118]) & (g599)) + ((g154) & (!g521) & (g597) & (g489) & (!sk[118]) & (!g599)) + ((g154) & (!g521) & (g597) & (g489) & (!sk[118]) & (g599)) + ((g154) & (!g521) & (g597) & (g489) & (sk[118]) & (g599)) + ((g154) & (g521) & (!g597) & (!g489) & (!sk[118]) & (!g599)) + ((g154) & (g521) & (!g597) & (!g489) & (!sk[118]) & (g599)) + ((g154) & (g521) & (!g597) & (!g489) & (sk[118]) & (g599)) + ((g154) & (g521) & (!g597) & (g489) & (!sk[118]) & (!g599)) + ((g154) & (g521) & (!g597) & (g489) & (!sk[118]) & (g599)) + ((g154) & (g521) & (!g597) & (g489) & (sk[118]) & (g599)) + ((g154) & (g521) & (g597) & (!g489) & (!sk[118]) & (!g599)) + ((g154) & (g521) & (g597) & (!g489) & (!sk[118]) & (g599)) + ((g154) & (g521) & (g597) & (!g489) & (sk[118]) & (g599)) + ((g154) & (g521) & (g597) & (g489) & (!sk[118]) & (!g599)) + ((g154) & (g521) & (g597) & (g489) & (!sk[118]) & (g599)) + ((g154) & (g521) & (g597) & (g489) & (sk[118]) & (g599)));
	assign g601 = (((!i_14_) & (!sk[119]) & (!g88) & (g123)) + ((!i_14_) & (!sk[119]) & (g88) & (!g123)) + ((!i_14_) & (!sk[119]) & (g88) & (g123)) + ((i_14_) & (!sk[119]) & (!g88) & (g123)) + ((i_14_) & (!sk[119]) & (g88) & (!g123)) + ((i_14_) & (!sk[119]) & (g88) & (g123)) + ((i_14_) & (sk[119]) & (g88) & (!g123)));
	assign g602 = (((!g123) & (!g186) & (!sk[120]) & (g513) & (!g514)) + ((!g123) & (!g186) & (!sk[120]) & (g513) & (g514)) + ((!g123) & (!g186) & (sk[120]) & (!g513) & (!g514)) + ((!g123) & (!g186) & (sk[120]) & (!g513) & (g514)) + ((!g123) & (!g186) & (sk[120]) & (g513) & (g514)) + ((!g123) & (g186) & (!sk[120]) & (g513) & (!g514)) + ((!g123) & (g186) & (!sk[120]) & (g513) & (g514)) + ((!g123) & (g186) & (sk[120]) & (!g513) & (!g514)) + ((!g123) & (g186) & (sk[120]) & (!g513) & (g514)) + ((!g123) & (g186) & (sk[120]) & (g513) & (!g514)) + ((!g123) & (g186) & (sk[120]) & (g513) & (g514)) + ((g123) & (!g186) & (!sk[120]) & (g513) & (!g514)) + ((g123) & (!g186) & (!sk[120]) & (g513) & (g514)) + ((g123) & (g186) & (!sk[120]) & (g513) & (!g514)) + ((g123) & (g186) & (!sk[120]) & (g513) & (g514)));
	assign g603 = (((!i_12_) & (!i_13_) & (i_14_) & (!sk[121]) & (!g91) & (g123)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[121]) & (g91) & (!g123)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[121]) & (g91) & (g123)) + ((!i_12_) & (!i_13_) & (i_14_) & (sk[121]) & (!g91) & (!g123)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[121]) & (!g91) & (!g123)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[121]) & (!g91) & (g123)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[121]) & (g91) & (!g123)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[121]) & (g91) & (g123)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[121]) & (!g91) & (!g123)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[121]) & (!g91) & (g123)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[121]) & (g91) & (!g123)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[121]) & (g91) & (g123)) + ((!i_12_) & (i_13_) & (i_14_) & (sk[121]) & (!g91) & (!g123)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[121]) & (!g91) & (g123)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[121]) & (g91) & (!g123)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[121]) & (g91) & (g123)) + ((i_12_) & (!i_13_) & (i_14_) & (sk[121]) & (!g91) & (!g123)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[121]) & (!g91) & (!g123)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[121]) & (!g91) & (g123)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[121]) & (g91) & (!g123)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[121]) & (g91) & (g123)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[121]) & (!g91) & (!g123)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[121]) & (!g91) & (g123)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[121]) & (g91) & (!g123)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[121]) & (g91) & (g123)));
	assign g604 = (((!sk[122]) & (!g142) & (!g521) & (g597) & (!g489)) + ((!sk[122]) & (!g142) & (!g521) & (g597) & (g489)) + ((!sk[122]) & (!g142) & (g521) & (g597) & (!g489)) + ((!sk[122]) & (!g142) & (g521) & (g597) & (g489)) + ((!sk[122]) & (g142) & (!g521) & (g597) & (!g489)) + ((!sk[122]) & (g142) & (!g521) & (g597) & (g489)) + ((!sk[122]) & (g142) & (g521) & (g597) & (!g489)) + ((!sk[122]) & (g142) & (g521) & (g597) & (g489)) + ((sk[122]) & (!g142) & (!g521) & (!g597) & (g489)) + ((sk[122]) & (!g142) & (!g521) & (g597) & (!g489)) + ((sk[122]) & (!g142) & (!g521) & (g597) & (g489)) + ((sk[122]) & (!g142) & (g521) & (!g597) & (!g489)) + ((sk[122]) & (!g142) & (g521) & (!g597) & (g489)) + ((sk[122]) & (!g142) & (g521) & (g597) & (!g489)) + ((sk[122]) & (!g142) & (g521) & (g597) & (g489)));
	assign g605 = (((!sk[123]) & (g36) & (!g174)) + ((!sk[123]) & (g36) & (g174)) + ((sk[123]) & (g36) & (!g174)));
	assign g606 = (((!g17) & (!sk[124]) & (!g421) & (g408) & (!g507)) + ((!g17) & (!sk[124]) & (!g421) & (g408) & (g507)) + ((!g17) & (!sk[124]) & (g421) & (g408) & (!g507)) + ((!g17) & (!sk[124]) & (g421) & (g408) & (g507)) + ((g17) & (!sk[124]) & (!g421) & (g408) & (!g507)) + ((g17) & (!sk[124]) & (!g421) & (g408) & (g507)) + ((g17) & (!sk[124]) & (g421) & (g408) & (!g507)) + ((g17) & (!sk[124]) & (g421) & (g408) & (g507)) + ((g17) & (sk[124]) & (!g421) & (!g408) & (g507)) + ((g17) & (sk[124]) & (g421) & (!g408) & (g507)) + ((g17) & (sk[124]) & (g421) & (g408) & (g507)));
	assign g607 = (((!sk[125]) & (g226) & (!g461)) + ((!sk[125]) & (g226) & (g461)) + ((sk[125]) & (!g226) & (g461)));
	assign g608 = (((!sk[126]) & (g81) & (!g174)) + ((!sk[126]) & (g81) & (g174)) + ((sk[126]) & (!g81) & (!g174)) + ((sk[126]) & (!g81) & (g174)) + ((sk[126]) & (g81) & (g174)));
	assign g609 = (((!sk[127]) & (!g177) & (!g392) & (g608)) + ((!sk[127]) & (!g177) & (g392) & (!g608)) + ((!sk[127]) & (!g177) & (g392) & (g608)) + ((!sk[127]) & (g177) & (!g392) & (g608)) + ((!sk[127]) & (g177) & (g392) & (!g608)) + ((!sk[127]) & (g177) & (g392) & (g608)) + ((sk[127]) & (!g177) & (g392) & (!g608)) + ((sk[127]) & (g177) & (g392) & (!g608)) + ((sk[127]) & (g177) & (g392) & (g608)));
	assign g610 = (((!sk[0]) & (!i_9_) & (!i_11_) & (i_15_) & (!g24)) + ((!sk[0]) & (!i_9_) & (!i_11_) & (i_15_) & (g24)) + ((!sk[0]) & (!i_9_) & (i_11_) & (i_15_) & (!g24)) + ((!sk[0]) & (!i_9_) & (i_11_) & (i_15_) & (g24)) + ((!sk[0]) & (i_9_) & (!i_11_) & (i_15_) & (!g24)) + ((!sk[0]) & (i_9_) & (!i_11_) & (i_15_) & (g24)) + ((!sk[0]) & (i_9_) & (i_11_) & (i_15_) & (!g24)) + ((!sk[0]) & (i_9_) & (i_11_) & (i_15_) & (g24)) + ((sk[0]) & (!i_9_) & (i_11_) & (i_15_) & (!g24)));
	assign g611 = (((!g24) & (!sk[1]) & (!g88) & (g113) & (!g174)) + ((!g24) & (!sk[1]) & (!g88) & (g113) & (g174)) + ((!g24) & (!sk[1]) & (g88) & (g113) & (!g174)) + ((!g24) & (!sk[1]) & (g88) & (g113) & (g174)) + ((!g24) & (sk[1]) & (!g88) & (g113) & (!g174)) + ((!g24) & (sk[1]) & (!g88) & (g113) & (g174)) + ((g24) & (!sk[1]) & (!g88) & (g113) & (!g174)) + ((g24) & (!sk[1]) & (!g88) & (g113) & (g174)) + ((g24) & (!sk[1]) & (g88) & (g113) & (!g174)) + ((g24) & (!sk[1]) & (g88) & (g113) & (g174)) + ((g24) & (sk[1]) & (!g88) & (!g113) & (g174)) + ((g24) & (sk[1]) & (!g88) & (g113) & (!g174)) + ((g24) & (sk[1]) & (!g88) & (g113) & (g174)) + ((g24) & (sk[1]) & (g88) & (!g113) & (g174)) + ((g24) & (sk[1]) & (g88) & (g113) & (g174)));
	assign g612 = (((!g1) & (!sk[2]) & (!i_15_) & (g34) & (!g120) & (g174)) + ((!g1) & (!sk[2]) & (!i_15_) & (g34) & (g120) & (!g174)) + ((!g1) & (!sk[2]) & (!i_15_) & (g34) & (g120) & (g174)) + ((!g1) & (!sk[2]) & (i_15_) & (!g34) & (!g120) & (!g174)) + ((!g1) & (!sk[2]) & (i_15_) & (!g34) & (!g120) & (g174)) + ((!g1) & (!sk[2]) & (i_15_) & (!g34) & (g120) & (!g174)) + ((!g1) & (!sk[2]) & (i_15_) & (!g34) & (g120) & (g174)) + ((!g1) & (!sk[2]) & (i_15_) & (g34) & (!g120) & (!g174)) + ((!g1) & (!sk[2]) & (i_15_) & (g34) & (!g120) & (g174)) + ((!g1) & (!sk[2]) & (i_15_) & (g34) & (g120) & (!g174)) + ((!g1) & (!sk[2]) & (i_15_) & (g34) & (g120) & (g174)) + ((g1) & (!sk[2]) & (!i_15_) & (g34) & (!g120) & (g174)) + ((g1) & (!sk[2]) & (!i_15_) & (g34) & (g120) & (!g174)) + ((g1) & (!sk[2]) & (!i_15_) & (g34) & (g120) & (g174)) + ((g1) & (!sk[2]) & (i_15_) & (!g34) & (!g120) & (!g174)) + ((g1) & (!sk[2]) & (i_15_) & (!g34) & (!g120) & (g174)) + ((g1) & (!sk[2]) & (i_15_) & (!g34) & (g120) & (!g174)) + ((g1) & (!sk[2]) & (i_15_) & (!g34) & (g120) & (g174)) + ((g1) & (!sk[2]) & (i_15_) & (g34) & (!g120) & (!g174)) + ((g1) & (!sk[2]) & (i_15_) & (g34) & (!g120) & (g174)) + ((g1) & (!sk[2]) & (i_15_) & (g34) & (g120) & (!g174)) + ((g1) & (!sk[2]) & (i_15_) & (g34) & (g120) & (g174)) + ((g1) & (sk[2]) & (!i_15_) & (g34) & (g120) & (!g174)));
	assign g613 = (((!g73) & (!g159) & (!g192) & (!g611) & (sk[3]) & (!g612)) + ((!g73) & (!g159) & (!g192) & (g611) & (sk[3]) & (!g612)) + ((!g73) & (!g159) & (g192) & (!g611) & (!sk[3]) & (g612)) + ((!g73) & (!g159) & (g192) & (g611) & (!sk[3]) & (!g612)) + ((!g73) & (!g159) & (g192) & (g611) & (!sk[3]) & (g612)) + ((!g73) & (g159) & (!g192) & (!g611) & (!sk[3]) & (!g612)) + ((!g73) & (g159) & (!g192) & (!g611) & (!sk[3]) & (g612)) + ((!g73) & (g159) & (!g192) & (!g611) & (sk[3]) & (!g612)) + ((!g73) & (g159) & (!g192) & (g611) & (!sk[3]) & (!g612)) + ((!g73) & (g159) & (!g192) & (g611) & (!sk[3]) & (g612)) + ((!g73) & (g159) & (!g192) & (g611) & (sk[3]) & (!g612)) + ((!g73) & (g159) & (g192) & (!g611) & (!sk[3]) & (!g612)) + ((!g73) & (g159) & (g192) & (!g611) & (!sk[3]) & (g612)) + ((!g73) & (g159) & (g192) & (!g611) & (sk[3]) & (!g612)) + ((!g73) & (g159) & (g192) & (g611) & (!sk[3]) & (!g612)) + ((!g73) & (g159) & (g192) & (g611) & (!sk[3]) & (g612)) + ((!g73) & (g159) & (g192) & (g611) & (sk[3]) & (!g612)) + ((g73) & (!g159) & (!g192) & (g611) & (sk[3]) & (!g612)) + ((g73) & (!g159) & (g192) & (!g611) & (!sk[3]) & (g612)) + ((g73) & (!g159) & (g192) & (g611) & (!sk[3]) & (!g612)) + ((g73) & (!g159) & (g192) & (g611) & (!sk[3]) & (g612)) + ((g73) & (g159) & (!g192) & (!g611) & (!sk[3]) & (!g612)) + ((g73) & (g159) & (!g192) & (!g611) & (!sk[3]) & (g612)) + ((g73) & (g159) & (!g192) & (g611) & (!sk[3]) & (!g612)) + ((g73) & (g159) & (!g192) & (g611) & (!sk[3]) & (g612)) + ((g73) & (g159) & (!g192) & (g611) & (sk[3]) & (!g612)) + ((g73) & (g159) & (g192) & (!g611) & (!sk[3]) & (!g612)) + ((g73) & (g159) & (g192) & (!g611) & (!sk[3]) & (g612)) + ((g73) & (g159) & (g192) & (g611) & (!sk[3]) & (!g612)) + ((g73) & (g159) & (g192) & (g611) & (!sk[3]) & (g612)) + ((g73) & (g159) & (g192) & (g611) & (sk[3]) & (!g612)));
	assign g614 = (((!g183) & (!g383) & (!g607) & (!g609) & (!g610) & (g613)) + ((!g183) & (g383) & (!g607) & (!g609) & (!g610) & (g613)) + ((!g183) & (g383) & (!g607) & (!g609) & (g610) & (g613)) + ((g183) & (g383) & (!g607) & (!g609) & (!g610) & (g613)) + ((g183) & (g383) & (!g607) & (!g609) & (g610) & (g613)));
	assign g615 = (((!g144) & (!g257) & (!sk[5]) & (g254) & (!g217) & (g226)) + ((!g144) & (!g257) & (!sk[5]) & (g254) & (g217) & (!g226)) + ((!g144) & (!g257) & (!sk[5]) & (g254) & (g217) & (g226)) + ((!g144) & (!g257) & (sk[5]) & (g254) & (!g217) & (g226)) + ((!g144) & (g257) & (!sk[5]) & (!g254) & (!g217) & (!g226)) + ((!g144) & (g257) & (!sk[5]) & (!g254) & (!g217) & (g226)) + ((!g144) & (g257) & (!sk[5]) & (!g254) & (g217) & (!g226)) + ((!g144) & (g257) & (!sk[5]) & (!g254) & (g217) & (g226)) + ((!g144) & (g257) & (!sk[5]) & (g254) & (!g217) & (!g226)) + ((!g144) & (g257) & (!sk[5]) & (g254) & (!g217) & (g226)) + ((!g144) & (g257) & (!sk[5]) & (g254) & (g217) & (!g226)) + ((!g144) & (g257) & (!sk[5]) & (g254) & (g217) & (g226)) + ((g144) & (!g257) & (!sk[5]) & (g254) & (!g217) & (g226)) + ((g144) & (!g257) & (!sk[5]) & (g254) & (g217) & (!g226)) + ((g144) & (!g257) & (!sk[5]) & (g254) & (g217) & (g226)) + ((g144) & (g257) & (!sk[5]) & (!g254) & (!g217) & (!g226)) + ((g144) & (g257) & (!sk[5]) & (!g254) & (!g217) & (g226)) + ((g144) & (g257) & (!sk[5]) & (!g254) & (g217) & (!g226)) + ((g144) & (g257) & (!sk[5]) & (!g254) & (g217) & (g226)) + ((g144) & (g257) & (!sk[5]) & (g254) & (!g217) & (!g226)) + ((g144) & (g257) & (!sk[5]) & (g254) & (!g217) & (g226)) + ((g144) & (g257) & (!sk[5]) & (g254) & (g217) & (!g226)) + ((g144) & (g257) & (!sk[5]) & (g254) & (g217) & (g226)));
	assign g616 = (((!g175) & (!g422) & (!g615) & (!g555) & (!g486) & (!g578)) + ((!g175) & (!g422) & (!g615) & (!g555) & (g486) & (!g578)) + ((!g175) & (!g422) & (!g615) & (g555) & (!g486) & (!g578)) + ((!g175) & (!g422) & (!g615) & (g555) & (g486) & (!g578)) + ((!g175) & (!g422) & (g615) & (!g555) & (!g486) & (!g578)) + ((!g175) & (!g422) & (g615) & (!g555) & (!g486) & (g578)) + ((!g175) & (!g422) & (g615) & (!g555) & (g486) & (!g578)) + ((!g175) & (!g422) & (g615) & (!g555) & (g486) & (g578)) + ((!g175) & (!g422) & (g615) & (g555) & (!g486) & (!g578)) + ((!g175) & (!g422) & (g615) & (g555) & (!g486) & (g578)) + ((!g175) & (!g422) & (g615) & (g555) & (g486) & (!g578)) + ((!g175) & (!g422) & (g615) & (g555) & (g486) & (g578)) + ((!g175) & (g422) & (!g615) & (!g555) & (!g486) & (!g578)) + ((!g175) & (g422) & (g615) & (!g555) & (!g486) & (!g578)) + ((!g175) & (g422) & (g615) & (!g555) & (!g486) & (g578)) + ((g175) & (!g422) & (!g615) & (!g555) & (!g486) & (!g578)) + ((g175) & (!g422) & (!g615) & (!g555) & (g486) & (!g578)) + ((g175) & (!g422) & (!g615) & (g555) & (!g486) & (!g578)) + ((g175) & (!g422) & (!g615) & (g555) & (g486) & (!g578)) + ((g175) & (!g422) & (g615) & (!g555) & (!g486) & (!g578)) + ((g175) & (!g422) & (g615) & (!g555) & (!g486) & (g578)) + ((g175) & (!g422) & (g615) & (!g555) & (g486) & (!g578)) + ((g175) & (!g422) & (g615) & (!g555) & (g486) & (g578)) + ((g175) & (!g422) & (g615) & (g555) & (!g486) & (!g578)) + ((g175) & (!g422) & (g615) & (g555) & (!g486) & (g578)) + ((g175) & (!g422) & (g615) & (g555) & (g486) & (!g578)) + ((g175) & (!g422) & (g615) & (g555) & (g486) & (g578)));
	assign g617 = (((!g161) & (!g191) & (g534) & (!sk[7]) & (!g496) & (g522)) + ((!g161) & (!g191) & (g534) & (!sk[7]) & (g496) & (!g522)) + ((!g161) & (!g191) & (g534) & (!sk[7]) & (g496) & (g522)) + ((!g161) & (g191) & (!g534) & (!sk[7]) & (!g496) & (!g522)) + ((!g161) & (g191) & (!g534) & (!sk[7]) & (!g496) & (g522)) + ((!g161) & (g191) & (!g534) & (!sk[7]) & (g496) & (!g522)) + ((!g161) & (g191) & (!g534) & (!sk[7]) & (g496) & (g522)) + ((!g161) & (g191) & (g534) & (!sk[7]) & (!g496) & (!g522)) + ((!g161) & (g191) & (g534) & (!sk[7]) & (!g496) & (g522)) + ((!g161) & (g191) & (g534) & (!sk[7]) & (g496) & (!g522)) + ((!g161) & (g191) & (g534) & (!sk[7]) & (g496) & (g522)) + ((g161) & (!g191) & (!g534) & (sk[7]) & (!g496) & (g522)) + ((g161) & (!g191) & (!g534) & (sk[7]) & (g496) & (!g522)) + ((g161) & (!g191) & (!g534) & (sk[7]) & (g496) & (g522)) + ((g161) & (!g191) & (g534) & (!sk[7]) & (!g496) & (g522)) + ((g161) & (!g191) & (g534) & (!sk[7]) & (g496) & (!g522)) + ((g161) & (!g191) & (g534) & (!sk[7]) & (g496) & (g522)) + ((g161) & (!g191) & (g534) & (sk[7]) & (!g496) & (!g522)) + ((g161) & (!g191) & (g534) & (sk[7]) & (!g496) & (g522)) + ((g161) & (!g191) & (g534) & (sk[7]) & (g496) & (!g522)) + ((g161) & (!g191) & (g534) & (sk[7]) & (g496) & (g522)) + ((g161) & (g191) & (!g534) & (!sk[7]) & (!g496) & (!g522)) + ((g161) & (g191) & (!g534) & (!sk[7]) & (!g496) & (g522)) + ((g161) & (g191) & (!g534) & (!sk[7]) & (g496) & (!g522)) + ((g161) & (g191) & (!g534) & (!sk[7]) & (g496) & (g522)) + ((g161) & (g191) & (!g534) & (sk[7]) & (!g496) & (!g522)) + ((g161) & (g191) & (!g534) & (sk[7]) & (!g496) & (g522)) + ((g161) & (g191) & (!g534) & (sk[7]) & (g496) & (!g522)) + ((g161) & (g191) & (!g534) & (sk[7]) & (g496) & (g522)) + ((g161) & (g191) & (g534) & (!sk[7]) & (!g496) & (!g522)) + ((g161) & (g191) & (g534) & (!sk[7]) & (!g496) & (g522)) + ((g161) & (g191) & (g534) & (!sk[7]) & (g496) & (!g522)) + ((g161) & (g191) & (g534) & (!sk[7]) & (g496) & (g522)) + ((g161) & (g191) & (g534) & (sk[7]) & (!g496) & (!g522)) + ((g161) & (g191) & (g534) & (sk[7]) & (!g496) & (g522)) + ((g161) & (g191) & (g534) & (sk[7]) & (g496) & (!g522)) + ((g161) & (g191) & (g534) & (sk[7]) & (g496) & (g522)));
	assign g618 = (((!g125) & (!g159) & (!g438) & (sk[8]) & (!g522) & (!g617)) + ((!g125) & (!g159) & (g438) & (!sk[8]) & (!g522) & (g617)) + ((!g125) & (!g159) & (g438) & (!sk[8]) & (g522) & (!g617)) + ((!g125) & (!g159) & (g438) & (!sk[8]) & (g522) & (g617)) + ((!g125) & (!g159) & (g438) & (sk[8]) & (!g522) & (!g617)) + ((!g125) & (g159) & (!g438) & (!sk[8]) & (!g522) & (!g617)) + ((!g125) & (g159) & (!g438) & (!sk[8]) & (!g522) & (g617)) + ((!g125) & (g159) & (!g438) & (!sk[8]) & (g522) & (!g617)) + ((!g125) & (g159) & (!g438) & (!sk[8]) & (g522) & (g617)) + ((!g125) & (g159) & (!g438) & (sk[8]) & (!g522) & (!g617)) + ((!g125) & (g159) & (g438) & (!sk[8]) & (!g522) & (!g617)) + ((!g125) & (g159) & (g438) & (!sk[8]) & (!g522) & (g617)) + ((!g125) & (g159) & (g438) & (!sk[8]) & (g522) & (!g617)) + ((!g125) & (g159) & (g438) & (!sk[8]) & (g522) & (g617)) + ((!g125) & (g159) & (g438) & (sk[8]) & (!g522) & (!g617)) + ((!g125) & (g159) & (g438) & (sk[8]) & (g522) & (!g617)) + ((g125) & (!g159) & (!g438) & (sk[8]) & (!g522) & (!g617)) + ((g125) & (!g159) & (g438) & (!sk[8]) & (!g522) & (g617)) + ((g125) & (!g159) & (g438) & (!sk[8]) & (g522) & (!g617)) + ((g125) & (!g159) & (g438) & (!sk[8]) & (g522) & (g617)) + ((g125) & (!g159) & (g438) & (sk[8]) & (!g522) & (!g617)) + ((g125) & (g159) & (!g438) & (!sk[8]) & (!g522) & (!g617)) + ((g125) & (g159) & (!g438) & (!sk[8]) & (!g522) & (g617)) + ((g125) & (g159) & (!g438) & (!sk[8]) & (g522) & (!g617)) + ((g125) & (g159) & (!g438) & (!sk[8]) & (g522) & (g617)) + ((g125) & (g159) & (!g438) & (sk[8]) & (!g522) & (!g617)) + ((g125) & (g159) & (g438) & (!sk[8]) & (!g522) & (!g617)) + ((g125) & (g159) & (g438) & (!sk[8]) & (!g522) & (g617)) + ((g125) & (g159) & (g438) & (!sk[8]) & (g522) & (!g617)) + ((g125) & (g159) & (g438) & (!sk[8]) & (g522) & (g617)) + ((g125) & (g159) & (g438) & (sk[8]) & (!g522) & (!g617)));
	assign g619 = (((!g601) & (!sk[9]) & (!g1458) & (g614) & (!g616) & (g618)) + ((!g601) & (!sk[9]) & (!g1458) & (g614) & (g616) & (!g618)) + ((!g601) & (!sk[9]) & (!g1458) & (g614) & (g616) & (g618)) + ((!g601) & (!sk[9]) & (g1458) & (!g614) & (!g616) & (!g618)) + ((!g601) & (!sk[9]) & (g1458) & (!g614) & (!g616) & (g618)) + ((!g601) & (!sk[9]) & (g1458) & (!g614) & (g616) & (!g618)) + ((!g601) & (!sk[9]) & (g1458) & (!g614) & (g616) & (g618)) + ((!g601) & (!sk[9]) & (g1458) & (g614) & (!g616) & (!g618)) + ((!g601) & (!sk[9]) & (g1458) & (g614) & (!g616) & (g618)) + ((!g601) & (!sk[9]) & (g1458) & (g614) & (g616) & (!g618)) + ((!g601) & (!sk[9]) & (g1458) & (g614) & (g616) & (g618)) + ((!g601) & (sk[9]) & (g1458) & (g614) & (g616) & (g618)) + ((g601) & (!sk[9]) & (!g1458) & (g614) & (!g616) & (g618)) + ((g601) & (!sk[9]) & (!g1458) & (g614) & (g616) & (!g618)) + ((g601) & (!sk[9]) & (!g1458) & (g614) & (g616) & (g618)) + ((g601) & (!sk[9]) & (g1458) & (!g614) & (!g616) & (!g618)) + ((g601) & (!sk[9]) & (g1458) & (!g614) & (!g616) & (g618)) + ((g601) & (!sk[9]) & (g1458) & (!g614) & (g616) & (!g618)) + ((g601) & (!sk[9]) & (g1458) & (!g614) & (g616) & (g618)) + ((g601) & (!sk[9]) & (g1458) & (g614) & (!g616) & (!g618)) + ((g601) & (!sk[9]) & (g1458) & (g614) & (!g616) & (g618)) + ((g601) & (!sk[9]) & (g1458) & (g614) & (g616) & (!g618)) + ((g601) & (!sk[9]) & (g1458) & (g614) & (g616) & (g618)));
	assign g620 = (((!g550) & (g581) & (g589) & (g596) & (g600) & (g619)));
	assign g621 = (((g269) & (g499) & (g525) & (g537) & (g549) & (g620)));
	assign o_8_ = (((!i_0_) & (!sk[12]) & (!i_1_) & (i_3_)) + ((!i_0_) & (!sk[12]) & (i_1_) & (!i_3_)) + ((!i_0_) & (!sk[12]) & (i_1_) & (i_3_)) + ((!i_0_) & (sk[12]) & (!i_1_) & (i_3_)) + ((i_0_) & (!sk[12]) & (!i_1_) & (i_3_)) + ((i_0_) & (!sk[12]) & (i_1_) & (!i_3_)) + ((i_0_) & (!sk[12]) & (i_1_) & (i_3_)));
	assign g623 = (((!g117) & (!g129) & (!sk[13]) & (g132) & (!g153)) + ((!g117) & (!g129) & (!sk[13]) & (g132) & (g153)) + ((!g117) & (g129) & (!sk[13]) & (g132) & (!g153)) + ((!g117) & (g129) & (!sk[13]) & (g132) & (g153)) + ((g117) & (!g129) & (!sk[13]) & (g132) & (!g153)) + ((g117) & (!g129) & (!sk[13]) & (g132) & (g153)) + ((g117) & (g129) & (!sk[13]) & (g132) & (!g153)) + ((g117) & (g129) & (!sk[13]) & (g132) & (g153)) + ((g117) & (g129) & (sk[13]) & (g132) & (g153)));
	assign g624 = (((!g18) & (!sk[14]) & (!g97) & (g578)) + ((!g18) & (!sk[14]) & (g97) & (!g578)) + ((!g18) & (!sk[14]) & (g97) & (g578)) + ((!g18) & (sk[14]) & (g97) & (!g578)) + ((g18) & (!sk[14]) & (!g97) & (g578)) + ((g18) & (!sk[14]) & (g97) & (!g578)) + ((g18) & (!sk[14]) & (g97) & (g578)));
	assign g625 = (((!i_12_) & (!sk[15]) & (!i_13_) & (i_14_) & (!g22)) + ((!i_12_) & (!sk[15]) & (!i_13_) & (i_14_) & (g22)) + ((!i_12_) & (!sk[15]) & (i_13_) & (i_14_) & (!g22)) + ((!i_12_) & (!sk[15]) & (i_13_) & (i_14_) & (g22)) + ((!i_12_) & (sk[15]) & (!i_13_) & (!i_14_) & (!g22)) + ((i_12_) & (!sk[15]) & (!i_13_) & (i_14_) & (!g22)) + ((i_12_) & (!sk[15]) & (!i_13_) & (i_14_) & (g22)) + ((i_12_) & (!sk[15]) & (i_13_) & (i_14_) & (!g22)) + ((i_12_) & (!sk[15]) & (i_13_) & (i_14_) & (g22)) + ((i_12_) & (sk[15]) & (!i_13_) & (!i_14_) & (!g22)) + ((i_12_) & (sk[15]) & (i_13_) & (!i_14_) & (!g22)));
	assign g626 = (((g19) & (!sk[16]) & (!g22)) + ((g19) & (!sk[16]) & (g22)) + ((g19) & (sk[16]) & (!g22)));
	assign g627 = (((!i_12_) & (!sk[17]) & (!i_13_) & (i_14_) & (!g88)) + ((!i_12_) & (!sk[17]) & (!i_13_) & (i_14_) & (g88)) + ((!i_12_) & (!sk[17]) & (i_13_) & (i_14_) & (!g88)) + ((!i_12_) & (!sk[17]) & (i_13_) & (i_14_) & (g88)) + ((!i_12_) & (sk[17]) & (!i_13_) & (!i_14_) & (g88)) + ((i_12_) & (!sk[17]) & (!i_13_) & (i_14_) & (!g88)) + ((i_12_) & (!sk[17]) & (!i_13_) & (i_14_) & (g88)) + ((i_12_) & (!sk[17]) & (i_13_) & (i_14_) & (!g88)) + ((i_12_) & (!sk[17]) & (i_13_) & (i_14_) & (g88)) + ((i_12_) & (sk[17]) & (!i_13_) & (!i_14_) & (g88)) + ((i_12_) & (sk[17]) & (i_13_) & (!i_14_) & (g88)));
	assign g628 = (((!g19) & (sk[18]) & (!g81)) + ((!g19) & (sk[18]) & (g81)) + ((g19) & (!sk[18]) & (!g81)) + ((g19) & (!sk[18]) & (g81)) + ((g19) & (sk[18]) & (!g81)));
	assign g629 = (((!i_12_) & (!i_13_) & (!i_14_) & (sk[19]) & (g81)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[19]) & (!g81)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[19]) & (g81)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[19]) & (!g81)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[19]) & (g81)) + ((i_12_) & (!i_13_) & (!i_14_) & (sk[19]) & (g81)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[19]) & (!g81)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[19]) & (g81)) + ((i_12_) & (i_13_) & (!i_14_) & (sk[19]) & (g81)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[19]) & (!g81)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[19]) & (g81)));
	assign g630 = (((g19) & (!sk[20]) & (!g88)) + ((g19) & (!sk[20]) & (g88)) + ((g19) & (sk[20]) & (g88)));
	assign g631 = (((!g154) & (!g624) & (!g627) & (!g628) & (!g629) & (!g630)) + ((!g154) & (!g624) & (!g627) & (!g628) & (!g629) & (g630)) + ((!g154) & (!g624) & (!g627) & (!g628) & (g629) & (!g630)) + ((!g154) & (!g624) & (!g627) & (!g628) & (g629) & (g630)) + ((!g154) & (!g624) & (!g627) & (g628) & (!g629) & (!g630)) + ((!g154) & (!g624) & (!g627) & (g628) & (!g629) & (g630)) + ((!g154) & (!g624) & (!g627) & (g628) & (g629) & (!g630)) + ((!g154) & (!g624) & (!g627) & (g628) & (g629) & (g630)) + ((!g154) & (!g624) & (g627) & (!g628) & (!g629) & (!g630)) + ((!g154) & (!g624) & (g627) & (!g628) & (!g629) & (g630)) + ((!g154) & (!g624) & (g627) & (!g628) & (g629) & (!g630)) + ((!g154) & (!g624) & (g627) & (!g628) & (g629) & (g630)) + ((!g154) & (!g624) & (g627) & (g628) & (!g629) & (!g630)) + ((!g154) & (!g624) & (g627) & (g628) & (!g629) & (g630)) + ((!g154) & (!g624) & (g627) & (g628) & (g629) & (!g630)) + ((!g154) & (!g624) & (g627) & (g628) & (g629) & (g630)) + ((!g154) & (g624) & (!g627) & (!g628) & (!g629) & (!g630)) + ((!g154) & (g624) & (!g627) & (!g628) & (!g629) & (g630)) + ((!g154) & (g624) & (!g627) & (!g628) & (g629) & (!g630)) + ((!g154) & (g624) & (!g627) & (!g628) & (g629) & (g630)) + ((!g154) & (g624) & (!g627) & (g628) & (!g629) & (g630)) + ((!g154) & (g624) & (!g627) & (g628) & (g629) & (!g630)) + ((!g154) & (g624) & (!g627) & (g628) & (g629) & (g630)) + ((!g154) & (g624) & (g627) & (!g628) & (!g629) & (!g630)) + ((!g154) & (g624) & (g627) & (!g628) & (!g629) & (g630)) + ((!g154) & (g624) & (g627) & (!g628) & (g629) & (!g630)) + ((!g154) & (g624) & (g627) & (!g628) & (g629) & (g630)) + ((!g154) & (g624) & (g627) & (g628) & (!g629) & (!g630)) + ((!g154) & (g624) & (g627) & (g628) & (!g629) & (g630)) + ((!g154) & (g624) & (g627) & (g628) & (g629) & (!g630)) + ((!g154) & (g624) & (g627) & (g628) & (g629) & (g630)));
	assign g632 = (((!g159) & (!g154) & (g624) & (!g625) & (!g626) & (!g631)) + ((!g159) & (g154) & (g624) & (!g625) & (!g626) & (!g631)) + ((!g159) & (g154) & (g624) & (!g625) & (g626) & (!g631)) + ((g159) & (!g154) & (!g624) & (!g625) & (!g626) & (!g631)) + ((g159) & (!g154) & (g624) & (!g625) & (!g626) & (!g631)) + ((g159) & (g154) & (!g624) & (!g625) & (!g626) & (!g631)) + ((g159) & (g154) & (!g624) & (!g625) & (g626) & (!g631)) + ((g159) & (g154) & (!g624) & (g625) & (!g626) & (!g631)) + ((g159) & (g154) & (!g624) & (g625) & (g626) & (!g631)) + ((g159) & (g154) & (g624) & (!g625) & (!g626) & (!g631)) + ((g159) & (g154) & (g624) & (!g625) & (g626) & (!g631)) + ((g159) & (g154) & (g624) & (g625) & (!g626) & (!g631)) + ((g159) & (g154) & (g624) & (g625) & (g626) & (!g631)));
	assign g633 = (((!g75) & (!sk[23]) & (!g102) & (g513) & (!g632)) + ((!g75) & (!sk[23]) & (!g102) & (g513) & (g632)) + ((!g75) & (!sk[23]) & (g102) & (g513) & (!g632)) + ((!g75) & (!sk[23]) & (g102) & (g513) & (g632)) + ((!g75) & (sk[23]) & (!g102) & (g513) & (g632)) + ((!g75) & (sk[23]) & (g102) & (g513) & (g632)) + ((g75) & (!sk[23]) & (!g102) & (g513) & (!g632)) + ((g75) & (!sk[23]) & (!g102) & (g513) & (g632)) + ((g75) & (!sk[23]) & (g102) & (g513) & (!g632)) + ((g75) & (!sk[23]) & (g102) & (g513) & (g632)) + ((g75) & (sk[23]) & (!g102) & (!g513) & (g632)) + ((g75) & (sk[23]) & (!g102) & (g513) & (g632)) + ((g75) & (sk[23]) & (g102) & (g513) & (g632)));
	assign g634 = (((!sk[24]) & (g19) & (!g35)) + ((!sk[24]) & (g19) & (g35)) + ((sk[24]) & (!g19) & (!g35)) + ((sk[24]) & (!g19) & (g35)) + ((sk[24]) & (g19) & (!g35)));
	assign g635 = (((g19) & (!sk[25]) & (!g36)) + ((g19) & (!sk[25]) & (g36)) + ((g19) & (sk[25]) & (g36)));
	assign g636 = (((!sk[26]) & (!i_8_) & (!g45) & (g394)) + ((!sk[26]) & (!i_8_) & (g45) & (!g394)) + ((!sk[26]) & (!i_8_) & (g45) & (g394)) + ((!sk[26]) & (i_8_) & (!g45) & (g394)) + ((!sk[26]) & (i_8_) & (g45) & (!g394)) + ((!sk[26]) & (i_8_) & (g45) & (g394)) + ((sk[26]) & (i_8_) & (g45) & (g394)));
	assign g637 = (((!i_9_) & (!i_10_) & (!i_11_) & (!g135) & (g630) & (!g636)) + ((!i_9_) & (!i_10_) & (!i_11_) & (!g135) & (g630) & (g636)) + ((!i_9_) & (!i_10_) & (i_11_) & (!g135) & (!g630) & (g636)) + ((!i_9_) & (!i_10_) & (i_11_) & (!g135) & (g630) & (!g636)) + ((!i_9_) & (!i_10_) & (i_11_) & (!g135) & (g630) & (g636)) + ((!i_9_) & (!i_10_) & (i_11_) & (g135) & (!g630) & (g636)) + ((!i_9_) & (!i_10_) & (i_11_) & (g135) & (g630) & (g636)) + ((!i_9_) & (i_10_) & (!i_11_) & (!g135) & (!g630) & (g636)) + ((!i_9_) & (i_10_) & (!i_11_) & (!g135) & (g630) & (!g636)) + ((!i_9_) & (i_10_) & (!i_11_) & (!g135) & (g630) & (g636)) + ((!i_9_) & (i_10_) & (!i_11_) & (g135) & (!g630) & (g636)) + ((!i_9_) & (i_10_) & (!i_11_) & (g135) & (g630) & (g636)) + ((!i_9_) & (i_10_) & (i_11_) & (!g135) & (!g630) & (g636)) + ((!i_9_) & (i_10_) & (i_11_) & (!g135) & (g630) & (!g636)) + ((!i_9_) & (i_10_) & (i_11_) & (!g135) & (g630) & (g636)) + ((!i_9_) & (i_10_) & (i_11_) & (g135) & (!g630) & (g636)) + ((!i_9_) & (i_10_) & (i_11_) & (g135) & (g630) & (g636)) + ((i_9_) & (!i_10_) & (!i_11_) & (!g135) & (g630) & (!g636)) + ((i_9_) & (!i_10_) & (!i_11_) & (!g135) & (g630) & (g636)) + ((i_9_) & (!i_10_) & (i_11_) & (!g135) & (g630) & (!g636)) + ((i_9_) & (!i_10_) & (i_11_) & (!g135) & (g630) & (g636)) + ((i_9_) & (i_10_) & (!i_11_) & (!g135) & (g630) & (!g636)) + ((i_9_) & (i_10_) & (!i_11_) & (!g135) & (g630) & (g636)) + ((i_9_) & (i_10_) & (i_11_) & (!g135) & (g630) & (!g636)) + ((i_9_) & (i_10_) & (i_11_) & (!g135) & (g630) & (g636)));
	assign g638 = (((!g17) & (g19) & (!g102) & (!g91) & (!g88) & (!g105)) + ((!g17) & (g19) & (!g102) & (!g91) & (g88) & (!g105)) + ((!g17) & (g19) & (!g102) & (g91) & (g88) & (!g105)) + ((!g17) & (g19) & (g102) & (!g91) & (!g88) & (!g105)) + ((!g17) & (g19) & (g102) & (!g91) & (g88) & (!g105)) + ((!g17) & (g19) & (g102) & (g91) & (g88) & (!g105)) + ((g17) & (g19) & (!g102) & (!g91) & (!g88) & (!g105)) + ((g17) & (g19) & (!g102) & (!g91) & (g88) & (!g105)) + ((g17) & (g19) & (!g102) & (g91) & (g88) & (!g105)) + ((g17) & (g19) & (g102) & (!g91) & (!g88) & (!g105)) + ((g17) & (g19) & (g102) & (!g91) & (!g88) & (g105)) + ((g17) & (g19) & (g102) & (!g91) & (g88) & (!g105)) + ((g17) & (g19) & (g102) & (!g91) & (g88) & (g105)) + ((g17) & (g19) & (g102) & (g91) & (!g88) & (!g105)) + ((g17) & (g19) & (g102) & (g91) & (!g88) & (g105)) + ((g17) & (g19) & (g102) & (g91) & (g88) & (!g105)) + ((g17) & (g19) & (g102) & (g91) & (g88) & (g105)));
	assign g639 = (((!g634) & (g105) & (!g383) & (!g635) & (!g637) & (!g638)) + ((!g634) & (g105) & (g383) & (!g635) & (!g637) & (!g638)) + ((!g634) & (g105) & (g383) & (g635) & (!g637) & (!g638)) + ((g634) & (!g105) & (!g383) & (!g635) & (!g637) & (!g638)) + ((g634) & (!g105) & (g383) & (!g635) & (!g637) & (!g638)) + ((g634) & (!g105) & (g383) & (g635) & (!g637) & (!g638)) + ((g634) & (g105) & (!g383) & (!g635) & (!g637) & (!g638)) + ((g634) & (g105) & (g383) & (!g635) & (!g637) & (!g638)) + ((g634) & (g105) & (g383) & (g635) & (!g637) & (!g638)));
	assign g640 = (((!i_13_) & (!sk[30]) & (!i_14_) & (g91)) + ((!i_13_) & (!sk[30]) & (i_14_) & (!g91)) + ((!i_13_) & (!sk[30]) & (i_14_) & (g91)) + ((!i_13_) & (sk[30]) & (!i_14_) & (!g91)) + ((i_13_) & (!sk[30]) & (!i_14_) & (g91)) + ((i_13_) & (!sk[30]) & (i_14_) & (!g91)) + ((i_13_) & (!sk[30]) & (i_14_) & (g91)));
	assign g641 = (((!sk[31]) & (!i_12_) & (!i_13_) & (i_14_) & (!g36)) + ((!sk[31]) & (!i_12_) & (!i_13_) & (i_14_) & (g36)) + ((!sk[31]) & (!i_12_) & (i_13_) & (i_14_) & (!g36)) + ((!sk[31]) & (!i_12_) & (i_13_) & (i_14_) & (g36)) + ((!sk[31]) & (i_12_) & (!i_13_) & (i_14_) & (!g36)) + ((!sk[31]) & (i_12_) & (!i_13_) & (i_14_) & (g36)) + ((!sk[31]) & (i_12_) & (i_13_) & (i_14_) & (!g36)) + ((!sk[31]) & (i_12_) & (i_13_) & (i_14_) & (g36)) + ((sk[31]) & (!i_12_) & (!i_13_) & (!i_14_) & (g36)) + ((sk[31]) & (i_12_) & (!i_13_) & (!i_14_) & (g36)) + ((sk[31]) & (i_12_) & (i_13_) & (!i_14_) & (g36)));
	assign g642 = (((!sk[32]) & (g19) & (!g113)) + ((!sk[32]) & (g19) & (g113)) + ((sk[32]) & (g19) & (!g113)));
	assign g643 = (((!g125) & (!g642) & (!sk[33]) & (g628) & (!g629)) + ((!g125) & (!g642) & (!sk[33]) & (g628) & (g629)) + ((!g125) & (g642) & (!sk[33]) & (g628) & (!g629)) + ((!g125) & (g642) & (!sk[33]) & (g628) & (g629)) + ((g125) & (!g642) & (!sk[33]) & (g628) & (!g629)) + ((g125) & (!g642) & (!sk[33]) & (g628) & (g629)) + ((g125) & (!g642) & (sk[33]) & (!g628) & (!g629)) + ((g125) & (!g642) & (sk[33]) & (!g628) & (g629)) + ((g125) & (!g642) & (sk[33]) & (g628) & (g629)) + ((g125) & (g642) & (!sk[33]) & (g628) & (!g629)) + ((g125) & (g642) & (!sk[33]) & (g628) & (g629)) + ((g125) & (g642) & (sk[33]) & (!g628) & (!g629)) + ((g125) & (g642) & (sk[33]) & (!g628) & (g629)) + ((g125) & (g642) & (sk[33]) & (g628) & (!g629)) + ((g125) & (g642) & (sk[33]) & (g628) & (g629)));
	assign g644 = (((!g356) & (!g640) & (!sk[34]) & (g641) & (!g629) & (g643)) + ((!g356) & (!g640) & (!sk[34]) & (g641) & (g629) & (!g643)) + ((!g356) & (!g640) & (!sk[34]) & (g641) & (g629) & (g643)) + ((!g356) & (!g640) & (sk[34]) & (!g641) & (!g629) & (!g643)) + ((!g356) & (!g640) & (sk[34]) & (!g641) & (g629) & (!g643)) + ((!g356) & (!g640) & (sk[34]) & (g641) & (!g629) & (!g643)) + ((!g356) & (!g640) & (sk[34]) & (g641) & (g629) & (!g643)) + ((!g356) & (g640) & (!sk[34]) & (!g641) & (!g629) & (!g643)) + ((!g356) & (g640) & (!sk[34]) & (!g641) & (!g629) & (g643)) + ((!g356) & (g640) & (!sk[34]) & (!g641) & (g629) & (!g643)) + ((!g356) & (g640) & (!sk[34]) & (!g641) & (g629) & (g643)) + ((!g356) & (g640) & (!sk[34]) & (g641) & (!g629) & (!g643)) + ((!g356) & (g640) & (!sk[34]) & (g641) & (!g629) & (g643)) + ((!g356) & (g640) & (!sk[34]) & (g641) & (g629) & (!g643)) + ((!g356) & (g640) & (!sk[34]) & (g641) & (g629) & (g643)) + ((!g356) & (g640) & (sk[34]) & (!g641) & (!g629) & (!g643)) + ((!g356) & (g640) & (sk[34]) & (!g641) & (g629) & (!g643)) + ((!g356) & (g640) & (sk[34]) & (g641) & (!g629) & (!g643)) + ((!g356) & (g640) & (sk[34]) & (g641) & (g629) & (!g643)) + ((g356) & (!g640) & (!sk[34]) & (g641) & (!g629) & (g643)) + ((g356) & (!g640) & (!sk[34]) & (g641) & (g629) & (!g643)) + ((g356) & (!g640) & (!sk[34]) & (g641) & (g629) & (g643)) + ((g356) & (!g640) & (sk[34]) & (!g641) & (!g629) & (!g643)) + ((g356) & (g640) & (!sk[34]) & (!g641) & (!g629) & (!g643)) + ((g356) & (g640) & (!sk[34]) & (!g641) & (!g629) & (g643)) + ((g356) & (g640) & (!sk[34]) & (!g641) & (g629) & (!g643)) + ((g356) & (g640) & (!sk[34]) & (!g641) & (g629) & (g643)) + ((g356) & (g640) & (!sk[34]) & (g641) & (!g629) & (!g643)) + ((g356) & (g640) & (!sk[34]) & (g641) & (!g629) & (g643)) + ((g356) & (g640) & (!sk[34]) & (g641) & (g629) & (!g643)) + ((g356) & (g640) & (!sk[34]) & (g641) & (g629) & (g643)));
	assign g645 = (((!sk[35]) & (!g164) & (!g625) & (g627)) + ((!sk[35]) & (!g164) & (g625) & (!g627)) + ((!sk[35]) & (!g164) & (g625) & (g627)) + ((!sk[35]) & (g164) & (!g625) & (g627)) + ((!sk[35]) & (g164) & (g625) & (!g627)) + ((!sk[35]) & (g164) & (g625) & (g627)) + ((sk[35]) & (g164) & (!g625) & (g627)) + ((sk[35]) & (g164) & (g625) & (!g627)) + ((sk[35]) & (g164) & (g625) & (g627)));
	assign g646 = (((!sk[36]) & (!g122) & (!g217) & (g635)) + ((!sk[36]) & (!g122) & (g217) & (!g635)) + ((!sk[36]) & (!g122) & (g217) & (g635)) + ((!sk[36]) & (g122) & (!g217) & (g635)) + ((!sk[36]) & (g122) & (g217) & (!g635)) + ((!sk[36]) & (g122) & (g217) & (g635)) + ((sk[36]) & (!g122) & (g217) & (g635)) + ((sk[36]) & (g122) & (!g217) & (g635)) + ((sk[36]) & (g122) & (g217) & (g635)));
	assign g647 = (((!i_12_) & (!i_13_) & (!sk[37]) & (i_14_) & (!g91) & (g105)) + ((!i_12_) & (!i_13_) & (!sk[37]) & (i_14_) & (g91) & (!g105)) + ((!i_12_) & (!i_13_) & (!sk[37]) & (i_14_) & (g91) & (g105)) + ((!i_12_) & (!i_13_) & (sk[37]) & (!i_14_) & (!g91) & (!g105)) + ((!i_12_) & (i_13_) & (!sk[37]) & (!i_14_) & (!g91) & (!g105)) + ((!i_12_) & (i_13_) & (!sk[37]) & (!i_14_) & (!g91) & (g105)) + ((!i_12_) & (i_13_) & (!sk[37]) & (!i_14_) & (g91) & (!g105)) + ((!i_12_) & (i_13_) & (!sk[37]) & (!i_14_) & (g91) & (g105)) + ((!i_12_) & (i_13_) & (!sk[37]) & (i_14_) & (!g91) & (!g105)) + ((!i_12_) & (i_13_) & (!sk[37]) & (i_14_) & (!g91) & (g105)) + ((!i_12_) & (i_13_) & (!sk[37]) & (i_14_) & (g91) & (!g105)) + ((!i_12_) & (i_13_) & (!sk[37]) & (i_14_) & (g91) & (g105)) + ((i_12_) & (!i_13_) & (!sk[37]) & (i_14_) & (!g91) & (g105)) + ((i_12_) & (!i_13_) & (!sk[37]) & (i_14_) & (g91) & (!g105)) + ((i_12_) & (!i_13_) & (!sk[37]) & (i_14_) & (g91) & (g105)) + ((i_12_) & (!i_13_) & (sk[37]) & (!i_14_) & (!g91) & (!g105)) + ((i_12_) & (i_13_) & (!sk[37]) & (!i_14_) & (!g91) & (!g105)) + ((i_12_) & (i_13_) & (!sk[37]) & (!i_14_) & (!g91) & (g105)) + ((i_12_) & (i_13_) & (!sk[37]) & (!i_14_) & (g91) & (!g105)) + ((i_12_) & (i_13_) & (!sk[37]) & (!i_14_) & (g91) & (g105)) + ((i_12_) & (i_13_) & (!sk[37]) & (i_14_) & (!g91) & (!g105)) + ((i_12_) & (i_13_) & (!sk[37]) & (i_14_) & (!g91) & (g105)) + ((i_12_) & (i_13_) & (!sk[37]) & (i_14_) & (g91) & (!g105)) + ((i_12_) & (i_13_) & (!sk[37]) & (i_14_) & (g91) & (g105)) + ((i_12_) & (i_13_) & (sk[37]) & (!i_14_) & (!g91) & (!g105)));
	assign g648 = (((g19) & (!sk[38]) & (!g86)) + ((g19) & (!sk[38]) & (g86)) + ((g19) & (sk[38]) & (g86)));
	assign g649 = (((!g102) & (!g642) & (g635) & (!sk[39]) & (!g648)) + ((!g102) & (!g642) & (g635) & (!sk[39]) & (g648)) + ((!g102) & (g642) & (g635) & (!sk[39]) & (!g648)) + ((!g102) & (g642) & (g635) & (!sk[39]) & (g648)) + ((g102) & (!g642) & (!g635) & (sk[39]) & (g648)) + ((g102) & (!g642) & (g635) & (!sk[39]) & (!g648)) + ((g102) & (!g642) & (g635) & (!sk[39]) & (g648)) + ((g102) & (!g642) & (g635) & (sk[39]) & (!g648)) + ((g102) & (!g642) & (g635) & (sk[39]) & (g648)) + ((g102) & (g642) & (!g635) & (sk[39]) & (!g648)) + ((g102) & (g642) & (!g635) & (sk[39]) & (g648)) + ((g102) & (g642) & (g635) & (!sk[39]) & (!g648)) + ((g102) & (g642) & (g635) & (!sk[39]) & (g648)) + ((g102) & (g642) & (g635) & (sk[39]) & (!g648)) + ((g102) & (g642) & (g635) & (sk[39]) & (g648)));
	assign g650 = (((!g36) & (!sk[40]) & (!g76) & (g91) & (!g88) & (g123)) + ((!g36) & (!sk[40]) & (!g76) & (g91) & (g88) & (!g123)) + ((!g36) & (!sk[40]) & (!g76) & (g91) & (g88) & (g123)) + ((!g36) & (!sk[40]) & (g76) & (!g91) & (!g88) & (!g123)) + ((!g36) & (!sk[40]) & (g76) & (!g91) & (!g88) & (g123)) + ((!g36) & (!sk[40]) & (g76) & (!g91) & (g88) & (!g123)) + ((!g36) & (!sk[40]) & (g76) & (!g91) & (g88) & (g123)) + ((!g36) & (!sk[40]) & (g76) & (g91) & (!g88) & (!g123)) + ((!g36) & (!sk[40]) & (g76) & (g91) & (!g88) & (g123)) + ((!g36) & (!sk[40]) & (g76) & (g91) & (g88) & (!g123)) + ((!g36) & (!sk[40]) & (g76) & (g91) & (g88) & (g123)) + ((!g36) & (sk[40]) & (!g76) & (!g91) & (!g88) & (!g123)) + ((!g36) & (sk[40]) & (!g76) & (!g91) & (g88) & (!g123)) + ((!g36) & (sk[40]) & (!g76) & (g91) & (g88) & (!g123)) + ((g36) & (!sk[40]) & (!g76) & (g91) & (!g88) & (g123)) + ((g36) & (!sk[40]) & (!g76) & (g91) & (g88) & (!g123)) + ((g36) & (!sk[40]) & (!g76) & (g91) & (g88) & (g123)) + ((g36) & (!sk[40]) & (g76) & (!g91) & (!g88) & (!g123)) + ((g36) & (!sk[40]) & (g76) & (!g91) & (!g88) & (g123)) + ((g36) & (!sk[40]) & (g76) & (!g91) & (g88) & (!g123)) + ((g36) & (!sk[40]) & (g76) & (!g91) & (g88) & (g123)) + ((g36) & (!sk[40]) & (g76) & (g91) & (!g88) & (!g123)) + ((g36) & (!sk[40]) & (g76) & (g91) & (!g88) & (g123)) + ((g36) & (!sk[40]) & (g76) & (g91) & (g88) & (!g123)) + ((g36) & (!sk[40]) & (g76) & (g91) & (g88) & (g123)) + ((g36) & (sk[40]) & (!g76) & (!g91) & (!g88) & (!g123)) + ((g36) & (sk[40]) & (!g76) & (!g91) & (g88) & (!g123)) + ((g36) & (sk[40]) & (!g76) & (g91) & (!g88) & (!g123)) + ((g36) & (sk[40]) & (!g76) & (g91) & (g88) & (!g123)));
	assign g651 = (((g19) & (!sk[41]) & (!g107)) + ((g19) & (!sk[41]) & (g107)) + ((g19) & (sk[41]) & (!g107)));
	assign g652 = (((!sk[42]) & (g19) & (!g91)) + ((!sk[42]) & (g19) & (g91)) + ((sk[42]) & (g19) & (!g91)));
	assign g653 = (((!g634) & (!g102) & (g651) & (!sk[43]) & (!g652)) + ((!g634) & (!g102) & (g651) & (!sk[43]) & (g652)) + ((!g634) & (g102) & (!g651) & (sk[43]) & (!g652)) + ((!g634) & (g102) & (!g651) & (sk[43]) & (g652)) + ((!g634) & (g102) & (g651) & (!sk[43]) & (!g652)) + ((!g634) & (g102) & (g651) & (!sk[43]) & (g652)) + ((!g634) & (g102) & (g651) & (sk[43]) & (!g652)) + ((!g634) & (g102) & (g651) & (sk[43]) & (g652)) + ((g634) & (!g102) & (g651) & (!sk[43]) & (!g652)) + ((g634) & (!g102) & (g651) & (!sk[43]) & (g652)) + ((g634) & (g102) & (!g651) & (sk[43]) & (g652)) + ((g634) & (g102) & (g651) & (!sk[43]) & (!g652)) + ((g634) & (g102) & (g651) & (!sk[43]) & (g652)) + ((g634) & (g102) & (g651) & (sk[43]) & (!g652)) + ((g634) & (g102) & (g651) & (sk[43]) & (g652)));
	assign g654 = (((!sk[44]) & (g4) & (!g69)) + ((!sk[44]) & (g4) & (g69)) + ((sk[44]) & (g4) & (g69)));
	assign g655 = (((!sk[45]) & (!g70) & (!g511) & (g654)) + ((!sk[45]) & (!g70) & (g511) & (!g654)) + ((!sk[45]) & (!g70) & (g511) & (g654)) + ((!sk[45]) & (g70) & (!g511) & (g654)) + ((!sk[45]) & (g70) & (g511) & (!g654)) + ((!sk[45]) & (g70) & (g511) & (g654)) + ((sk[45]) & (!g70) & (!g511) & (!g654)));
	assign g656 = (((!i_8_) & (!i_6_) & (!i_7_) & (g118) & (!g655) & (g630)) + ((!i_8_) & (!i_6_) & (!i_7_) & (g118) & (g655) & (g630)) + ((!i_8_) & (i_6_) & (i_7_) & (g118) & (!g655) & (!g630)) + ((!i_8_) & (i_6_) & (i_7_) & (g118) & (!g655) & (g630)) + ((i_8_) & (!i_6_) & (!i_7_) & (g118) & (!g655) & (g630)) + ((i_8_) & (!i_6_) & (!i_7_) & (g118) & (g655) & (g630)) + ((i_8_) & (i_6_) & (!i_7_) & (g118) & (!g655) & (g630)) + ((i_8_) & (i_6_) & (!i_7_) & (g118) & (g655) & (g630)));
	assign g657 = (((!g647) & (!g649) & (!g650) & (!g653) & (sk[47]) & (!g656)) + ((!g647) & (!g649) & (g650) & (!g653) & (!sk[47]) & (g656)) + ((!g647) & (!g649) & (g650) & (g653) & (!sk[47]) & (!g656)) + ((!g647) & (!g649) & (g650) & (g653) & (!sk[47]) & (g656)) + ((!g647) & (g649) & (!g650) & (!g653) & (!sk[47]) & (!g656)) + ((!g647) & (g649) & (!g650) & (!g653) & (!sk[47]) & (g656)) + ((!g647) & (g649) & (!g650) & (g653) & (!sk[47]) & (!g656)) + ((!g647) & (g649) & (!g650) & (g653) & (!sk[47]) & (g656)) + ((!g647) & (g649) & (g650) & (!g653) & (!sk[47]) & (!g656)) + ((!g647) & (g649) & (g650) & (!g653) & (!sk[47]) & (g656)) + ((!g647) & (g649) & (g650) & (g653) & (!sk[47]) & (!g656)) + ((!g647) & (g649) & (g650) & (g653) & (!sk[47]) & (g656)) + ((g647) & (!g649) & (g650) & (!g653) & (!sk[47]) & (g656)) + ((g647) & (!g649) & (g650) & (g653) & (!sk[47]) & (!g656)) + ((g647) & (!g649) & (g650) & (g653) & (!sk[47]) & (g656)) + ((g647) & (g649) & (!g650) & (!g653) & (!sk[47]) & (!g656)) + ((g647) & (g649) & (!g650) & (!g653) & (!sk[47]) & (g656)) + ((g647) & (g649) & (!g650) & (g653) & (!sk[47]) & (!g656)) + ((g647) & (g649) & (!g650) & (g653) & (!sk[47]) & (g656)) + ((g647) & (g649) & (g650) & (!g653) & (!sk[47]) & (!g656)) + ((g647) & (g649) & (g650) & (!g653) & (!sk[47]) & (g656)) + ((g647) & (g649) & (g650) & (g653) & (!sk[47]) & (!g656)) + ((g647) & (g649) & (g650) & (g653) & (!sk[47]) & (g656)));
	assign g658 = (((!g17) & (!g19) & (g27) & (!g226) & (!sk[48]) & (g227)) + ((!g17) & (!g19) & (g27) & (g226) & (!sk[48]) & (!g227)) + ((!g17) & (!g19) & (g27) & (g226) & (!sk[48]) & (g227)) + ((!g17) & (g19) & (!g27) & (!g226) & (!sk[48]) & (!g227)) + ((!g17) & (g19) & (!g27) & (!g226) & (!sk[48]) & (g227)) + ((!g17) & (g19) & (!g27) & (g226) & (!sk[48]) & (!g227)) + ((!g17) & (g19) & (!g27) & (g226) & (!sk[48]) & (g227)) + ((!g17) & (g19) & (g27) & (!g226) & (!sk[48]) & (!g227)) + ((!g17) & (g19) & (g27) & (!g226) & (!sk[48]) & (g227)) + ((!g17) & (g19) & (g27) & (!g226) & (sk[48]) & (!g227)) + ((!g17) & (g19) & (g27) & (!g226) & (sk[48]) & (g227)) + ((!g17) & (g19) & (g27) & (g226) & (!sk[48]) & (!g227)) + ((!g17) & (g19) & (g27) & (g226) & (!sk[48]) & (g227)) + ((g17) & (!g19) & (g27) & (!g226) & (!sk[48]) & (g227)) + ((g17) & (!g19) & (g27) & (g226) & (!sk[48]) & (!g227)) + ((g17) & (!g19) & (g27) & (g226) & (!sk[48]) & (g227)) + ((g17) & (g19) & (!g27) & (!g226) & (!sk[48]) & (!g227)) + ((g17) & (g19) & (!g27) & (!g226) & (!sk[48]) & (g227)) + ((g17) & (g19) & (!g27) & (!g226) & (sk[48]) & (g227)) + ((g17) & (g19) & (!g27) & (g226) & (!sk[48]) & (!g227)) + ((g17) & (g19) & (!g27) & (g226) & (!sk[48]) & (g227)) + ((g17) & (g19) & (!g27) & (g226) & (sk[48]) & (g227)) + ((g17) & (g19) & (g27) & (!g226) & (!sk[48]) & (!g227)) + ((g17) & (g19) & (g27) & (!g226) & (!sk[48]) & (g227)) + ((g17) & (g19) & (g27) & (!g226) & (sk[48]) & (!g227)) + ((g17) & (g19) & (g27) & (!g226) & (sk[48]) & (g227)) + ((g17) & (g19) & (g27) & (g226) & (!sk[48]) & (!g227)) + ((g17) & (g19) & (g27) & (g226) & (!sk[48]) & (g227)) + ((g17) & (g19) & (g27) & (g226) & (sk[48]) & (g227)));
	assign g659 = (((!i_8_) & (!sk[49]) & (!g17) & (g19) & (!g36) & (g73)) + ((!i_8_) & (!sk[49]) & (!g17) & (g19) & (g36) & (!g73)) + ((!i_8_) & (!sk[49]) & (!g17) & (g19) & (g36) & (g73)) + ((!i_8_) & (!sk[49]) & (g17) & (!g19) & (!g36) & (!g73)) + ((!i_8_) & (!sk[49]) & (g17) & (!g19) & (!g36) & (g73)) + ((!i_8_) & (!sk[49]) & (g17) & (!g19) & (g36) & (!g73)) + ((!i_8_) & (!sk[49]) & (g17) & (!g19) & (g36) & (g73)) + ((!i_8_) & (!sk[49]) & (g17) & (g19) & (!g36) & (!g73)) + ((!i_8_) & (!sk[49]) & (g17) & (g19) & (!g36) & (g73)) + ((!i_8_) & (!sk[49]) & (g17) & (g19) & (g36) & (!g73)) + ((!i_8_) & (!sk[49]) & (g17) & (g19) & (g36) & (g73)) + ((i_8_) & (!sk[49]) & (!g17) & (g19) & (!g36) & (g73)) + ((i_8_) & (!sk[49]) & (!g17) & (g19) & (g36) & (!g73)) + ((i_8_) & (!sk[49]) & (!g17) & (g19) & (g36) & (g73)) + ((i_8_) & (!sk[49]) & (g17) & (!g19) & (!g36) & (!g73)) + ((i_8_) & (!sk[49]) & (g17) & (!g19) & (!g36) & (g73)) + ((i_8_) & (!sk[49]) & (g17) & (!g19) & (g36) & (!g73)) + ((i_8_) & (!sk[49]) & (g17) & (!g19) & (g36) & (g73)) + ((i_8_) & (!sk[49]) & (g17) & (g19) & (!g36) & (!g73)) + ((i_8_) & (!sk[49]) & (g17) & (g19) & (!g36) & (g73)) + ((i_8_) & (!sk[49]) & (g17) & (g19) & (g36) & (!g73)) + ((i_8_) & (!sk[49]) & (g17) & (g19) & (g36) & (g73)) + ((i_8_) & (sk[49]) & (!g17) & (g19) & (g36) & (g73)) + ((i_8_) & (sk[49]) & (g17) & (g19) & (!g36) & (g73)) + ((i_8_) & (sk[49]) & (g17) & (g19) & (g36) & (g73)));
	assign g660 = (((!g135) & (!g130) & (!g131) & (sk[50]) & (g635)) + ((!g135) & (!g130) & (g131) & (!sk[50]) & (!g635)) + ((!g135) & (!g130) & (g131) & (!sk[50]) & (g635)) + ((!g135) & (!g130) & (g131) & (sk[50]) & (g635)) + ((!g135) & (g130) & (!g131) & (sk[50]) & (g635)) + ((!g135) & (g130) & (g131) & (!sk[50]) & (!g635)) + ((!g135) & (g130) & (g131) & (!sk[50]) & (g635)) + ((!g135) & (g130) & (g131) & (sk[50]) & (g635)) + ((g135) & (!g130) & (!g131) & (sk[50]) & (g635)) + ((g135) & (!g130) & (g131) & (!sk[50]) & (!g635)) + ((g135) & (!g130) & (g131) & (!sk[50]) & (g635)) + ((g135) & (!g130) & (g131) & (sk[50]) & (g635)) + ((g135) & (g130) & (!g131) & (sk[50]) & (g635)) + ((g135) & (g130) & (g131) & (!sk[50]) & (!g635)) + ((g135) & (g130) & (g131) & (!sk[50]) & (g635)));
	assign g661 = (((!g105) & (!g543) & (!g513) & (sk[51]) & (!g635)) + ((!g105) & (!g543) & (!g513) & (sk[51]) & (g635)) + ((!g105) & (!g543) & (g513) & (!sk[51]) & (!g635)) + ((!g105) & (!g543) & (g513) & (!sk[51]) & (g635)) + ((!g105) & (!g543) & (g513) & (sk[51]) & (g635)) + ((!g105) & (g543) & (!g513) & (sk[51]) & (!g635)) + ((!g105) & (g543) & (!g513) & (sk[51]) & (g635)) + ((!g105) & (g543) & (g513) & (!sk[51]) & (!g635)) + ((!g105) & (g543) & (g513) & (!sk[51]) & (g635)) + ((!g105) & (g543) & (g513) & (sk[51]) & (!g635)) + ((!g105) & (g543) & (g513) & (sk[51]) & (g635)) + ((g105) & (!g543) & (g513) & (!sk[51]) & (!g635)) + ((g105) & (!g543) & (g513) & (!sk[51]) & (g635)) + ((g105) & (g543) & (g513) & (!sk[51]) & (!g635)) + ((g105) & (g543) & (g513) & (!sk[51]) & (g635)));
	assign g662 = (((!g36) & (!sk[52]) & (!g76) & (g125) & (!g91) & (g88)) + ((!g36) & (!sk[52]) & (!g76) & (g125) & (g91) & (!g88)) + ((!g36) & (!sk[52]) & (!g76) & (g125) & (g91) & (g88)) + ((!g36) & (!sk[52]) & (g76) & (!g125) & (!g91) & (!g88)) + ((!g36) & (!sk[52]) & (g76) & (!g125) & (!g91) & (g88)) + ((!g36) & (!sk[52]) & (g76) & (!g125) & (g91) & (!g88)) + ((!g36) & (!sk[52]) & (g76) & (!g125) & (g91) & (g88)) + ((!g36) & (!sk[52]) & (g76) & (g125) & (!g91) & (!g88)) + ((!g36) & (!sk[52]) & (g76) & (g125) & (!g91) & (g88)) + ((!g36) & (!sk[52]) & (g76) & (g125) & (g91) & (!g88)) + ((!g36) & (!sk[52]) & (g76) & (g125) & (g91) & (g88)) + ((!g36) & (sk[52]) & (!g76) & (g125) & (!g91) & (!g88)) + ((!g36) & (sk[52]) & (!g76) & (g125) & (!g91) & (g88)) + ((!g36) & (sk[52]) & (!g76) & (g125) & (g91) & (g88)) + ((g36) & (!sk[52]) & (!g76) & (g125) & (!g91) & (g88)) + ((g36) & (!sk[52]) & (!g76) & (g125) & (g91) & (!g88)) + ((g36) & (!sk[52]) & (!g76) & (g125) & (g91) & (g88)) + ((g36) & (!sk[52]) & (g76) & (!g125) & (!g91) & (!g88)) + ((g36) & (!sk[52]) & (g76) & (!g125) & (!g91) & (g88)) + ((g36) & (!sk[52]) & (g76) & (!g125) & (g91) & (!g88)) + ((g36) & (!sk[52]) & (g76) & (!g125) & (g91) & (g88)) + ((g36) & (!sk[52]) & (g76) & (g125) & (!g91) & (!g88)) + ((g36) & (!sk[52]) & (g76) & (g125) & (!g91) & (g88)) + ((g36) & (!sk[52]) & (g76) & (g125) & (g91) & (!g88)) + ((g36) & (!sk[52]) & (g76) & (g125) & (g91) & (g88)) + ((g36) & (sk[52]) & (!g76) & (g125) & (!g91) & (!g88)) + ((g36) & (sk[52]) & (!g76) & (g125) & (!g91) & (g88)) + ((g36) & (sk[52]) & (!g76) & (g125) & (g91) & (!g88)) + ((g36) & (sk[52]) & (!g76) & (g125) & (g91) & (g88)));
	assign g663 = (((!g658) & (!g659) & (!g660) & (!g661) & (sk[53]) & (!g662)) + ((!g658) & (!g659) & (g660) & (!g661) & (!sk[53]) & (g662)) + ((!g658) & (!g659) & (g660) & (g661) & (!sk[53]) & (!g662)) + ((!g658) & (!g659) & (g660) & (g661) & (!sk[53]) & (g662)) + ((!g658) & (g659) & (!g660) & (!g661) & (!sk[53]) & (!g662)) + ((!g658) & (g659) & (!g660) & (!g661) & (!sk[53]) & (g662)) + ((!g658) & (g659) & (!g660) & (g661) & (!sk[53]) & (!g662)) + ((!g658) & (g659) & (!g660) & (g661) & (!sk[53]) & (g662)) + ((!g658) & (g659) & (g660) & (!g661) & (!sk[53]) & (!g662)) + ((!g658) & (g659) & (g660) & (!g661) & (!sk[53]) & (g662)) + ((!g658) & (g659) & (g660) & (g661) & (!sk[53]) & (!g662)) + ((!g658) & (g659) & (g660) & (g661) & (!sk[53]) & (g662)) + ((g658) & (!g659) & (g660) & (!g661) & (!sk[53]) & (g662)) + ((g658) & (!g659) & (g660) & (g661) & (!sk[53]) & (!g662)) + ((g658) & (!g659) & (g660) & (g661) & (!sk[53]) & (g662)) + ((g658) & (g659) & (!g660) & (!g661) & (!sk[53]) & (!g662)) + ((g658) & (g659) & (!g660) & (!g661) & (!sk[53]) & (g662)) + ((g658) & (g659) & (!g660) & (g661) & (!sk[53]) & (!g662)) + ((g658) & (g659) & (!g660) & (g661) & (!sk[53]) & (g662)) + ((g658) & (g659) & (g660) & (!g661) & (!sk[53]) & (!g662)) + ((g658) & (g659) & (g660) & (!g661) & (!sk[53]) & (g662)) + ((g658) & (g659) & (g660) & (g661) & (!sk[53]) & (!g662)) + ((g658) & (g659) & (g660) & (g661) & (!sk[53]) & (g662)));
	assign g664 = (((!i_12_) & (!sk[54]) & (!i_13_) & (i_14_) & (!g113)) + ((!i_12_) & (!sk[54]) & (!i_13_) & (i_14_) & (g113)) + ((!i_12_) & (!sk[54]) & (i_13_) & (i_14_) & (!g113)) + ((!i_12_) & (!sk[54]) & (i_13_) & (i_14_) & (g113)) + ((!i_12_) & (sk[54]) & (!i_13_) & (!i_14_) & (!g113)) + ((i_12_) & (!sk[54]) & (!i_13_) & (i_14_) & (!g113)) + ((i_12_) & (!sk[54]) & (!i_13_) & (i_14_) & (g113)) + ((i_12_) & (!sk[54]) & (i_13_) & (i_14_) & (!g113)) + ((i_12_) & (!sk[54]) & (i_13_) & (i_14_) & (g113)) + ((i_12_) & (sk[54]) & (!i_13_) & (!i_14_) & (!g113)) + ((i_12_) & (sk[54]) & (i_13_) & (!i_14_) & (!g113)));
	assign g665 = (((!i_12_) & (!i_13_) & (!sk[55]) & (i_14_) & (!g91)) + ((!i_12_) & (!i_13_) & (!sk[55]) & (i_14_) & (g91)) + ((!i_12_) & (!i_13_) & (sk[55]) & (!i_14_) & (!g91)) + ((!i_12_) & (i_13_) & (!sk[55]) & (i_14_) & (!g91)) + ((!i_12_) & (i_13_) & (!sk[55]) & (i_14_) & (g91)) + ((i_12_) & (!i_13_) & (!sk[55]) & (i_14_) & (!g91)) + ((i_12_) & (!i_13_) & (!sk[55]) & (i_14_) & (g91)) + ((i_12_) & (!i_13_) & (sk[55]) & (!i_14_) & (!g91)) + ((i_12_) & (i_13_) & (!sk[55]) & (i_14_) & (!g91)) + ((i_12_) & (i_13_) & (!sk[55]) & (i_14_) & (g91)) + ((i_12_) & (i_13_) & (sk[55]) & (!i_14_) & (!g91)));
	assign g666 = (((!g164) & (!g253) & (g624) & (!sk[56]) & (!g664) & (g665)) + ((!g164) & (!g253) & (g624) & (!sk[56]) & (g664) & (!g665)) + ((!g164) & (!g253) & (g624) & (!sk[56]) & (g664) & (g665)) + ((!g164) & (!g253) & (g624) & (sk[56]) & (!g664) & (!g665)) + ((!g164) & (g253) & (!g624) & (!sk[56]) & (!g664) & (!g665)) + ((!g164) & (g253) & (!g624) & (!sk[56]) & (!g664) & (g665)) + ((!g164) & (g253) & (!g624) & (!sk[56]) & (g664) & (!g665)) + ((!g164) & (g253) & (!g624) & (!sk[56]) & (g664) & (g665)) + ((!g164) & (g253) & (!g624) & (sk[56]) & (!g664) & (!g665)) + ((!g164) & (g253) & (!g624) & (sk[56]) & (!g664) & (g665)) + ((!g164) & (g253) & (!g624) & (sk[56]) & (g664) & (!g665)) + ((!g164) & (g253) & (!g624) & (sk[56]) & (g664) & (g665)) + ((!g164) & (g253) & (g624) & (!sk[56]) & (!g664) & (!g665)) + ((!g164) & (g253) & (g624) & (!sk[56]) & (!g664) & (g665)) + ((!g164) & (g253) & (g624) & (!sk[56]) & (g664) & (!g665)) + ((!g164) & (g253) & (g624) & (!sk[56]) & (g664) & (g665)) + ((!g164) & (g253) & (g624) & (sk[56]) & (!g664) & (!g665)) + ((!g164) & (g253) & (g624) & (sk[56]) & (!g664) & (g665)) + ((!g164) & (g253) & (g624) & (sk[56]) & (g664) & (!g665)) + ((!g164) & (g253) & (g624) & (sk[56]) & (g664) & (g665)) + ((g164) & (!g253) & (g624) & (!sk[56]) & (!g664) & (g665)) + ((g164) & (!g253) & (g624) & (!sk[56]) & (g664) & (!g665)) + ((g164) & (!g253) & (g624) & (!sk[56]) & (g664) & (g665)) + ((g164) & (!g253) & (g624) & (sk[56]) & (!g664) & (!g665)) + ((g164) & (g253) & (!g624) & (!sk[56]) & (!g664) & (!g665)) + ((g164) & (g253) & (!g624) & (!sk[56]) & (!g664) & (g665)) + ((g164) & (g253) & (!g624) & (!sk[56]) & (g664) & (!g665)) + ((g164) & (g253) & (!g624) & (!sk[56]) & (g664) & (g665)) + ((g164) & (g253) & (g624) & (!sk[56]) & (!g664) & (!g665)) + ((g164) & (g253) & (g624) & (!sk[56]) & (!g664) & (g665)) + ((g164) & (g253) & (g624) & (!sk[56]) & (g664) & (!g665)) + ((g164) & (g253) & (g624) & (!sk[56]) & (g664) & (g665)) + ((g164) & (g253) & (g624) & (sk[56]) & (!g664) & (!g665)) + ((g164) & (g253) & (g624) & (sk[56]) & (!g664) & (g665)) + ((g164) & (g253) & (g624) & (sk[56]) & (g664) & (!g665)) + ((g164) & (g253) & (g624) & (sk[56]) & (g664) & (g665)));
	assign g667 = (((!g125) & (!sk[57]) & (!g226) & (g408) & (!g624) & (g666)) + ((!g125) & (!sk[57]) & (!g226) & (g408) & (g624) & (!g666)) + ((!g125) & (!sk[57]) & (!g226) & (g408) & (g624) & (g666)) + ((!g125) & (!sk[57]) & (g226) & (!g408) & (!g624) & (!g666)) + ((!g125) & (!sk[57]) & (g226) & (!g408) & (!g624) & (g666)) + ((!g125) & (!sk[57]) & (g226) & (!g408) & (g624) & (!g666)) + ((!g125) & (!sk[57]) & (g226) & (!g408) & (g624) & (g666)) + ((!g125) & (!sk[57]) & (g226) & (g408) & (!g624) & (!g666)) + ((!g125) & (!sk[57]) & (g226) & (g408) & (!g624) & (g666)) + ((!g125) & (!sk[57]) & (g226) & (g408) & (g624) & (!g666)) + ((!g125) & (!sk[57]) & (g226) & (g408) & (g624) & (g666)) + ((!g125) & (sk[57]) & (!g226) & (!g408) & (g624) & (g666)) + ((!g125) & (sk[57]) & (!g226) & (g408) & (g624) & (g666)) + ((!g125) & (sk[57]) & (g226) & (!g408) & (g624) & (g666)) + ((!g125) & (sk[57]) & (g226) & (g408) & (!g624) & (g666)) + ((!g125) & (sk[57]) & (g226) & (g408) & (g624) & (g666)) + ((g125) & (!sk[57]) & (!g226) & (g408) & (!g624) & (g666)) + ((g125) & (!sk[57]) & (!g226) & (g408) & (g624) & (!g666)) + ((g125) & (!sk[57]) & (!g226) & (g408) & (g624) & (g666)) + ((g125) & (!sk[57]) & (g226) & (!g408) & (!g624) & (!g666)) + ((g125) & (!sk[57]) & (g226) & (!g408) & (!g624) & (g666)) + ((g125) & (!sk[57]) & (g226) & (!g408) & (g624) & (!g666)) + ((g125) & (!sk[57]) & (g226) & (!g408) & (g624) & (g666)) + ((g125) & (!sk[57]) & (g226) & (g408) & (!g624) & (!g666)) + ((g125) & (!sk[57]) & (g226) & (g408) & (!g624) & (g666)) + ((g125) & (!sk[57]) & (g226) & (g408) & (g624) & (!g666)) + ((g125) & (!sk[57]) & (g226) & (g408) & (g624) & (g666)) + ((g125) & (sk[57]) & (!g226) & (!g408) & (g624) & (g666)) + ((g125) & (sk[57]) & (!g226) & (g408) & (g624) & (g666)) + ((g125) & (sk[57]) & (g226) & (!g408) & (g624) & (g666)) + ((g125) & (sk[57]) & (g226) & (g408) & (g624) & (g666)));
	assign g668 = (((g3) & (!sk[58]) & (!g19)) + ((g3) & (!sk[58]) & (g19)) + ((g3) & (sk[58]) & (g19)));
	assign g669 = (((!i_11_) & (!sk[59]) & (!i_15_) & (g53) & (!g76) & (g668)) + ((!i_11_) & (!sk[59]) & (!i_15_) & (g53) & (g76) & (!g668)) + ((!i_11_) & (!sk[59]) & (!i_15_) & (g53) & (g76) & (g668)) + ((!i_11_) & (!sk[59]) & (i_15_) & (!g53) & (!g76) & (!g668)) + ((!i_11_) & (!sk[59]) & (i_15_) & (!g53) & (!g76) & (g668)) + ((!i_11_) & (!sk[59]) & (i_15_) & (!g53) & (g76) & (!g668)) + ((!i_11_) & (!sk[59]) & (i_15_) & (!g53) & (g76) & (g668)) + ((!i_11_) & (!sk[59]) & (i_15_) & (g53) & (!g76) & (!g668)) + ((!i_11_) & (!sk[59]) & (i_15_) & (g53) & (!g76) & (g668)) + ((!i_11_) & (!sk[59]) & (i_15_) & (g53) & (g76) & (!g668)) + ((!i_11_) & (!sk[59]) & (i_15_) & (g53) & (g76) & (g668)) + ((!i_11_) & (sk[59]) & (!i_15_) & (!g53) & (!g76) & (!g668)) + ((!i_11_) & (sk[59]) & (!i_15_) & (!g53) & (g76) & (!g668)) + ((!i_11_) & (sk[59]) & (!i_15_) & (g53) & (!g76) & (!g668)) + ((!i_11_) & (sk[59]) & (!i_15_) & (g53) & (g76) & (!g668)) + ((!i_11_) & (sk[59]) & (i_15_) & (!g53) & (!g76) & (!g668)) + ((!i_11_) & (sk[59]) & (i_15_) & (!g53) & (g76) & (!g668)) + ((!i_11_) & (sk[59]) & (i_15_) & (g53) & (!g76) & (!g668)) + ((!i_11_) & (sk[59]) & (i_15_) & (g53) & (g76) & (!g668)) + ((i_11_) & (!sk[59]) & (!i_15_) & (g53) & (!g76) & (g668)) + ((i_11_) & (!sk[59]) & (!i_15_) & (g53) & (g76) & (!g668)) + ((i_11_) & (!sk[59]) & (!i_15_) & (g53) & (g76) & (g668)) + ((i_11_) & (!sk[59]) & (i_15_) & (!g53) & (!g76) & (!g668)) + ((i_11_) & (!sk[59]) & (i_15_) & (!g53) & (!g76) & (g668)) + ((i_11_) & (!sk[59]) & (i_15_) & (!g53) & (g76) & (!g668)) + ((i_11_) & (!sk[59]) & (i_15_) & (!g53) & (g76) & (g668)) + ((i_11_) & (!sk[59]) & (i_15_) & (g53) & (!g76) & (!g668)) + ((i_11_) & (!sk[59]) & (i_15_) & (g53) & (!g76) & (g668)) + ((i_11_) & (!sk[59]) & (i_15_) & (g53) & (g76) & (!g668)) + ((i_11_) & (!sk[59]) & (i_15_) & (g53) & (g76) & (g668)) + ((i_11_) & (sk[59]) & (!i_15_) & (!g53) & (!g76) & (!g668)) + ((i_11_) & (sk[59]) & (!i_15_) & (!g53) & (g76) & (!g668)) + ((i_11_) & (sk[59]) & (!i_15_) & (g53) & (!g76) & (!g668)) + ((i_11_) & (sk[59]) & (!i_15_) & (g53) & (g76) & (!g668)) + ((i_11_) & (sk[59]) & (i_15_) & (!g53) & (!g76) & (!g668)) + ((i_11_) & (sk[59]) & (i_15_) & (!g53) & (g76) & (!g668)) + ((i_11_) & (sk[59]) & (i_15_) & (g53) & (g76) & (!g668)));
	assign g670 = (((!i_8_) & (!g73) & (g635) & (!sk[60]) & (!g652)) + ((!i_8_) & (!g73) & (g635) & (!sk[60]) & (g652)) + ((!i_8_) & (g73) & (!g635) & (sk[60]) & (g652)) + ((!i_8_) & (g73) & (g635) & (!sk[60]) & (!g652)) + ((!i_8_) & (g73) & (g635) & (!sk[60]) & (g652)) + ((!i_8_) & (g73) & (g635) & (sk[60]) & (!g652)) + ((!i_8_) & (g73) & (g635) & (sk[60]) & (g652)) + ((i_8_) & (!g73) & (g635) & (!sk[60]) & (!g652)) + ((i_8_) & (!g73) & (g635) & (!sk[60]) & (g652)) + ((i_8_) & (g73) & (g635) & (!sk[60]) & (!g652)) + ((i_8_) & (g73) & (g635) & (!sk[60]) & (g652)));
	assign g671 = (((!g75) & (!g168) & (!g350) & (!g652) & (!g669) & (!g670)) + ((!g75) & (!g168) & (!g350) & (!g652) & (g669) & (!g670)) + ((!g75) & (!g168) & (g350) & (!g652) & (!g669) & (!g670)) + ((!g75) & (!g168) & (g350) & (!g652) & (g669) & (!g670)) + ((!g75) & (g168) & (!g350) & (!g652) & (g669) & (!g670)) + ((!g75) & (g168) & (g350) & (!g652) & (g669) & (!g670)) + ((g75) & (!g168) & (!g350) & (!g652) & (!g669) & (!g670)) + ((g75) & (!g168) & (!g350) & (!g652) & (g669) & (!g670)) + ((g75) & (!g168) & (!g350) & (g652) & (!g669) & (!g670)) + ((g75) & (!g168) & (!g350) & (g652) & (g669) & (!g670)) + ((g75) & (!g168) & (g350) & (!g652) & (!g669) & (!g670)) + ((g75) & (!g168) & (g350) & (!g652) & (g669) & (!g670)) + ((g75) & (g168) & (!g350) & (!g652) & (g669) & (!g670)) + ((g75) & (g168) & (!g350) & (g652) & (g669) & (!g670)) + ((g75) & (g168) & (g350) & (!g652) & (g669) & (!g670)));
	assign g672 = (((!g645) & (!g646) & (g657) & (g663) & (g667) & (g671)));
	assign g673 = (((!sk[63]) & (!g253) & (!g641) & (g635)) + ((!sk[63]) & (!g253) & (g641) & (!g635)) + ((!sk[63]) & (!g253) & (g641) & (g635)) + ((!sk[63]) & (g253) & (!g641) & (g635)) + ((!sk[63]) & (g253) & (g641) & (!g635)) + ((!sk[63]) & (g253) & (g641) & (g635)) + ((sk[63]) & (!g253) & (!g641) & (g635)) + ((sk[63]) & (!g253) & (g641) & (!g635)) + ((sk[63]) & (!g253) & (g641) & (g635)));
	assign g674 = (((!g30) & (!g120) & (!sk[64]) & (g626) & (!g630)) + ((!g30) & (!g120) & (!sk[64]) & (g626) & (g630)) + ((!g30) & (g120) & (!sk[64]) & (g626) & (!g630)) + ((!g30) & (g120) & (!sk[64]) & (g626) & (g630)) + ((g30) & (!g120) & (!sk[64]) & (g626) & (!g630)) + ((g30) & (!g120) & (!sk[64]) & (g626) & (g630)) + ((g30) & (g120) & (!sk[64]) & (g626) & (!g630)) + ((g30) & (g120) & (!sk[64]) & (g626) & (g630)) + ((g30) & (g120) & (sk[64]) & (!g626) & (g630)) + ((g30) & (g120) & (sk[64]) & (g626) & (!g630)) + ((g30) & (g120) & (sk[64]) & (g626) & (g630)));
	assign g675 = (((!g164) & (!g641) & (!g628) & (!g655) & (!g665) & (!g674)) + ((!g164) & (!g641) & (!g628) & (!g655) & (g665) & (!g674)) + ((!g164) & (!g641) & (!g628) & (g655) & (!g665) & (!g674)) + ((!g164) & (!g641) & (!g628) & (g655) & (g665) & (!g674)) + ((!g164) & (!g641) & (g628) & (!g655) & (!g665) & (!g674)) + ((!g164) & (!g641) & (g628) & (!g655) & (g665) & (!g674)) + ((!g164) & (!g641) & (g628) & (g655) & (!g665) & (!g674)) + ((!g164) & (!g641) & (g628) & (g655) & (g665) & (!g674)) + ((!g164) & (g641) & (!g628) & (!g655) & (!g665) & (!g674)) + ((!g164) & (g641) & (!g628) & (!g655) & (g665) & (!g674)) + ((!g164) & (g641) & (!g628) & (g655) & (!g665) & (!g674)) + ((!g164) & (g641) & (!g628) & (g655) & (g665) & (!g674)) + ((!g164) & (g641) & (g628) & (!g655) & (!g665) & (!g674)) + ((!g164) & (g641) & (g628) & (!g655) & (g665) & (!g674)) + ((!g164) & (g641) & (g628) & (g655) & (!g665) & (!g674)) + ((!g164) & (g641) & (g628) & (g655) & (g665) & (!g674)) + ((g164) & (!g641) & (g628) & (g655) & (!g665) & (!g674)));
	assign g676 = (((!g253) & (!g625) & (!g627) & (!g629) & (!g673) & (g675)) + ((g253) & (!g625) & (!g627) & (!g629) & (!g673) & (g675)) + ((g253) & (!g625) & (!g627) & (g629) & (!g673) & (g675)) + ((g253) & (!g625) & (g627) & (!g629) & (!g673) & (g675)) + ((g253) & (!g625) & (g627) & (g629) & (!g673) & (g675)) + ((g253) & (g625) & (!g627) & (!g629) & (!g673) & (g675)) + ((g253) & (g625) & (!g627) & (g629) & (!g673) & (g675)) + ((g253) & (g625) & (g627) & (!g629) & (!g673) & (g675)) + ((g253) & (g625) & (g627) & (g629) & (!g673) & (g675)));
	assign g677 = (((!i_12_) & (!i_13_) & (!sk[67]) & (g17)) + ((!i_12_) & (i_13_) & (!sk[67]) & (!g17)) + ((!i_12_) & (i_13_) & (!sk[67]) & (g17)) + ((!i_12_) & (i_13_) & (sk[67]) & (g17)) + ((i_12_) & (!i_13_) & (!sk[67]) & (g17)) + ((i_12_) & (i_13_) & (!sk[67]) & (!g17)) + ((i_12_) & (i_13_) & (!sk[67]) & (g17)));
	assign g678 = (((!i_14_) & (!g142) & (!g254) & (!g425) & (!g402) & (g677)) + ((!i_14_) & (!g142) & (!g254) & (!g425) & (g402) & (g677)) + ((!i_14_) & (!g142) & (!g254) & (g425) & (!g402) & (g677)) + ((!i_14_) & (!g142) & (!g254) & (g425) & (g402) & (g677)) + ((!i_14_) & (!g142) & (g254) & (!g425) & (!g402) & (g677)) + ((!i_14_) & (!g142) & (g254) & (g425) & (!g402) & (g677)) + ((!i_14_) & (g142) & (!g254) & (!g425) & (!g402) & (g677)) + ((!i_14_) & (g142) & (!g254) & (!g425) & (g402) & (g677)) + ((!i_14_) & (g142) & (!g254) & (g425) & (!g402) & (g677)) + ((!i_14_) & (g142) & (!g254) & (g425) & (g402) & (g677)) + ((!i_14_) & (g142) & (g254) & (!g425) & (!g402) & (g677)) + ((!i_14_) & (g142) & (g254) & (g425) & (!g402) & (g677)) + ((i_14_) & (!g142) & (!g254) & (!g425) & (!g402) & (g677)) + ((i_14_) & (!g142) & (!g254) & (!g425) & (g402) & (g677)) + ((i_14_) & (!g142) & (!g254) & (g425) & (!g402) & (g677)) + ((i_14_) & (!g142) & (!g254) & (g425) & (g402) & (g677)) + ((i_14_) & (!g142) & (g254) & (!g425) & (!g402) & (g677)) + ((i_14_) & (!g142) & (g254) & (!g425) & (g402) & (g677)) + ((i_14_) & (!g142) & (g254) & (g425) & (!g402) & (g677)) + ((i_14_) & (!g142) & (g254) & (g425) & (g402) & (g677)) + ((i_14_) & (g142) & (!g254) & (!g425) & (!g402) & (g677)) + ((i_14_) & (g142) & (!g254) & (!g425) & (g402) & (g677)) + ((i_14_) & (g142) & (g254) & (!g425) & (!g402) & (g677)) + ((i_14_) & (g142) & (g254) & (!g425) & (g402) & (g677)));
	assign g679 = (((!sk[69]) & (!i_11_) & (!i_15_) & (g19) & (!g53) & (g401)) + ((!sk[69]) & (!i_11_) & (!i_15_) & (g19) & (g53) & (!g401)) + ((!sk[69]) & (!i_11_) & (!i_15_) & (g19) & (g53) & (g401)) + ((!sk[69]) & (!i_11_) & (i_15_) & (!g19) & (!g53) & (!g401)) + ((!sk[69]) & (!i_11_) & (i_15_) & (!g19) & (!g53) & (g401)) + ((!sk[69]) & (!i_11_) & (i_15_) & (!g19) & (g53) & (!g401)) + ((!sk[69]) & (!i_11_) & (i_15_) & (!g19) & (g53) & (g401)) + ((!sk[69]) & (!i_11_) & (i_15_) & (g19) & (!g53) & (!g401)) + ((!sk[69]) & (!i_11_) & (i_15_) & (g19) & (!g53) & (g401)) + ((!sk[69]) & (!i_11_) & (i_15_) & (g19) & (g53) & (!g401)) + ((!sk[69]) & (!i_11_) & (i_15_) & (g19) & (g53) & (g401)) + ((!sk[69]) & (i_11_) & (!i_15_) & (g19) & (!g53) & (g401)) + ((!sk[69]) & (i_11_) & (!i_15_) & (g19) & (g53) & (!g401)) + ((!sk[69]) & (i_11_) & (!i_15_) & (g19) & (g53) & (g401)) + ((!sk[69]) & (i_11_) & (i_15_) & (!g19) & (!g53) & (!g401)) + ((!sk[69]) & (i_11_) & (i_15_) & (!g19) & (!g53) & (g401)) + ((!sk[69]) & (i_11_) & (i_15_) & (!g19) & (g53) & (!g401)) + ((!sk[69]) & (i_11_) & (i_15_) & (!g19) & (g53) & (g401)) + ((!sk[69]) & (i_11_) & (i_15_) & (g19) & (!g53) & (!g401)) + ((!sk[69]) & (i_11_) & (i_15_) & (g19) & (!g53) & (g401)) + ((!sk[69]) & (i_11_) & (i_15_) & (g19) & (g53) & (!g401)) + ((!sk[69]) & (i_11_) & (i_15_) & (g19) & (g53) & (g401)) + ((sk[69]) & (i_11_) & (!i_15_) & (g19) & (!g53) & (!g401)));
	assign g680 = (((!g3) & (g19) & (!g35) & (!g425) & (!g402) & (g353)) + ((!g3) & (g19) & (g35) & (!g425) & (!g402) & (g353)) + ((!g3) & (g19) & (g35) & (!g425) & (g402) & (g353)) + ((g3) & (g19) & (!g35) & (!g425) & (!g402) & (g353)) + ((g3) & (g19) & (!g35) & (g425) & (!g402) & (g353)) + ((g3) & (g19) & (g35) & (!g425) & (!g402) & (g353)) + ((g3) & (g19) & (g35) & (!g425) & (g402) & (g353)) + ((g3) & (g19) & (g35) & (g425) & (!g402) & (g353)));
	assign g681 = (((!g80) & (!sk[71]) & (!i_11_) & (g636)) + ((!g80) & (!sk[71]) & (i_11_) & (!g636)) + ((!g80) & (!sk[71]) & (i_11_) & (g636)) + ((g80) & (!sk[71]) & (!i_11_) & (g636)) + ((g80) & (!sk[71]) & (i_11_) & (!g636)) + ((g80) & (!sk[71]) & (i_11_) & (g636)) + ((g80) & (sk[71]) & (!i_11_) & (g636)));
	assign g682 = (((!g122) & (!sk[72]) & (!g123) & (g105) & (!g642) & (g626)) + ((!g122) & (!sk[72]) & (!g123) & (g105) & (g642) & (!g626)) + ((!g122) & (!sk[72]) & (!g123) & (g105) & (g642) & (g626)) + ((!g122) & (!sk[72]) & (g123) & (!g105) & (!g642) & (!g626)) + ((!g122) & (!sk[72]) & (g123) & (!g105) & (!g642) & (g626)) + ((!g122) & (!sk[72]) & (g123) & (!g105) & (g642) & (!g626)) + ((!g122) & (!sk[72]) & (g123) & (!g105) & (g642) & (g626)) + ((!g122) & (!sk[72]) & (g123) & (g105) & (!g642) & (!g626)) + ((!g122) & (!sk[72]) & (g123) & (g105) & (!g642) & (g626)) + ((!g122) & (!sk[72]) & (g123) & (g105) & (g642) & (!g626)) + ((!g122) & (!sk[72]) & (g123) & (g105) & (g642) & (g626)) + ((!g122) & (sk[72]) & (!g123) & (!g105) & (!g642) & (!g626)) + ((!g122) & (sk[72]) & (!g123) & (g105) & (!g642) & (!g626)) + ((!g122) & (sk[72]) & (!g123) & (g105) & (!g642) & (g626)) + ((!g122) & (sk[72]) & (g123) & (!g105) & (!g642) & (!g626)) + ((!g122) & (sk[72]) & (g123) & (g105) & (!g642) & (!g626)) + ((!g122) & (sk[72]) & (g123) & (g105) & (!g642) & (g626)) + ((!g122) & (sk[72]) & (g123) & (g105) & (g642) & (!g626)) + ((!g122) & (sk[72]) & (g123) & (g105) & (g642) & (g626)) + ((g122) & (!sk[72]) & (!g123) & (g105) & (!g642) & (g626)) + ((g122) & (!sk[72]) & (!g123) & (g105) & (g642) & (!g626)) + ((g122) & (!sk[72]) & (!g123) & (g105) & (g642) & (g626)) + ((g122) & (!sk[72]) & (g123) & (!g105) & (!g642) & (!g626)) + ((g122) & (!sk[72]) & (g123) & (!g105) & (!g642) & (g626)) + ((g122) & (!sk[72]) & (g123) & (!g105) & (g642) & (!g626)) + ((g122) & (!sk[72]) & (g123) & (!g105) & (g642) & (g626)) + ((g122) & (!sk[72]) & (g123) & (g105) & (!g642) & (!g626)) + ((g122) & (!sk[72]) & (g123) & (g105) & (!g642) & (g626)) + ((g122) & (!sk[72]) & (g123) & (g105) & (g642) & (!g626)) + ((g122) & (!sk[72]) & (g123) & (g105) & (g642) & (g626)) + ((g122) & (sk[72]) & (!g123) & (!g105) & (!g642) & (!g626)) + ((g122) & (sk[72]) & (!g123) & (g105) & (!g642) & (!g626)) + ((g122) & (sk[72]) & (g123) & (!g105) & (!g642) & (!g626)) + ((g122) & (sk[72]) & (g123) & (g105) & (!g642) & (!g626)) + ((g122) & (sk[72]) & (g123) & (g105) & (g642) & (!g626)));
	assign g683 = (((!i_12_) & (!i_14_) & (g88) & (!sk[73]) & (!g408)) + ((!i_12_) & (!i_14_) & (g88) & (!sk[73]) & (g408)) + ((!i_12_) & (i_14_) & (g88) & (!sk[73]) & (!g408)) + ((!i_12_) & (i_14_) & (g88) & (!sk[73]) & (g408)) + ((i_12_) & (!i_14_) & (g88) & (!sk[73]) & (!g408)) + ((i_12_) & (!i_14_) & (g88) & (!sk[73]) & (g408)) + ((i_12_) & (!i_14_) & (g88) & (sk[73]) & (!g408)) + ((i_12_) & (i_14_) & (g88) & (!sk[73]) & (!g408)) + ((i_12_) & (i_14_) & (g88) & (!sk[73]) & (g408)));
	assign g684 = (((!sk[74]) & (g4) & (!g113)) + ((!sk[74]) & (g4) & (g113)) + ((sk[74]) & (!g4) & (!g113)) + ((sk[74]) & (!g4) & (g113)) + ((sk[74]) & (g4) & (g113)));
	assign g685 = (((!sk[75]) & (!g135) & (!g131) & (g664) & (!g684)) + ((!sk[75]) & (!g135) & (!g131) & (g664) & (g684)) + ((!sk[75]) & (!g135) & (g131) & (g664) & (!g684)) + ((!sk[75]) & (!g135) & (g131) & (g664) & (g684)) + ((!sk[75]) & (g135) & (!g131) & (g664) & (!g684)) + ((!sk[75]) & (g135) & (!g131) & (g664) & (g684)) + ((!sk[75]) & (g135) & (g131) & (g664) & (!g684)) + ((!sk[75]) & (g135) & (g131) & (g664) & (g684)) + ((sk[75]) & (!g135) & (!g131) & (!g664) & (!g684)) + ((sk[75]) & (!g135) & (!g131) & (g664) & (!g684)) + ((sk[75]) & (!g135) & (!g131) & (g664) & (g684)) + ((sk[75]) & (!g135) & (g131) & (!g664) & (!g684)) + ((sk[75]) & (!g135) & (g131) & (g664) & (!g684)) + ((sk[75]) & (g135) & (!g131) & (g664) & (!g684)) + ((sk[75]) & (g135) & (!g131) & (g664) & (g684)));
	assign g686 = (((!i_12_) & (!i_13_) & (!i_14_) & (!g22) & (!g142) & (!g408)) + ((!i_12_) & (!i_13_) & (!i_14_) & (!g22) & (!g142) & (g408)) + ((i_12_) & (!i_13_) & (!i_14_) & (!g22) & (!g142) & (!g408)) + ((i_12_) & (!i_13_) & (!i_14_) & (!g22) & (!g142) & (g408)) + ((i_12_) & (!i_13_) & (!i_14_) & (!g22) & (g142) & (!g408)) + ((i_12_) & (i_13_) & (!i_14_) & (!g22) & (!g142) & (!g408)) + ((i_12_) & (i_13_) & (!i_14_) & (!g22) & (!g142) & (g408)) + ((i_12_) & (i_13_) & (!i_14_) & (!g22) & (g142) & (!g408)));
	assign g687 = (((!i_8_) & (!g73) & (!sk[77]) & (g102) & (!g562)) + ((!i_8_) & (!g73) & (!sk[77]) & (g102) & (g562)) + ((!i_8_) & (!g73) & (sk[77]) & (g102) & (g562)) + ((!i_8_) & (g73) & (!sk[77]) & (g102) & (!g562)) + ((!i_8_) & (g73) & (!sk[77]) & (g102) & (g562)) + ((!i_8_) & (g73) & (sk[77]) & (g102) & (g562)) + ((i_8_) & (!g73) & (!sk[77]) & (g102) & (!g562)) + ((i_8_) & (!g73) & (!sk[77]) & (g102) & (g562)) + ((i_8_) & (!g73) & (sk[77]) & (g102) & (g562)) + ((i_8_) & (g73) & (!sk[77]) & (g102) & (!g562)) + ((i_8_) & (g73) & (!sk[77]) & (g102) & (g562)) + ((i_8_) & (g73) & (sk[77]) & (!g102) & (g562)) + ((i_8_) & (g73) & (sk[77]) & (g102) & (g562)));
	assign g688 = (((!i_12_) & (!sk[78]) & (!i_14_) & (g113)) + ((!i_12_) & (!sk[78]) & (i_14_) & (!g113)) + ((!i_12_) & (!sk[78]) & (i_14_) & (g113)) + ((i_12_) & (!sk[78]) & (!i_14_) & (g113)) + ((i_12_) & (!sk[78]) & (i_14_) & (!g113)) + ((i_12_) & (!sk[78]) & (i_14_) & (g113)) + ((i_12_) & (sk[78]) & (!i_14_) & (!g113)));
	assign g689 = (((!g125) & (!g164) & (!g254) & (!g217) & (!g629) & (!g688)) + ((!g125) & (!g164) & (!g254) & (!g217) & (g629) & (!g688)) + ((!g125) & (!g164) & (!g254) & (g217) & (!g629) & (!g688)) + ((!g125) & (!g164) & (!g254) & (g217) & (g629) & (!g688)) + ((!g125) & (!g164) & (g254) & (!g217) & (!g629) & (!g688)) + ((!g125) & (!g164) & (g254) & (!g217) & (!g629) & (g688)) + ((!g125) & (!g164) & (g254) & (!g217) & (g629) & (!g688)) + ((!g125) & (!g164) & (g254) & (!g217) & (g629) & (g688)) + ((!g125) & (!g164) & (g254) & (g217) & (!g629) & (!g688)) + ((!g125) & (!g164) & (g254) & (g217) & (g629) & (!g688)) + ((!g125) & (g164) & (!g254) & (!g217) & (!g629) & (!g688)) + ((!g125) & (g164) & (!g254) & (g217) & (!g629) & (!g688)) + ((!g125) & (g164) & (g254) & (!g217) & (!g629) & (!g688)) + ((!g125) & (g164) & (g254) & (!g217) & (!g629) & (g688)) + ((!g125) & (g164) & (g254) & (g217) & (!g629) & (!g688)) + ((g125) & (!g164) & (!g254) & (!g217) & (!g629) & (!g688)) + ((g125) & (!g164) & (!g254) & (!g217) & (g629) & (!g688)) + ((g125) & (!g164) & (!g254) & (g217) & (!g629) & (!g688)) + ((g125) & (!g164) & (!g254) & (g217) & (g629) & (!g688)) + ((g125) & (!g164) & (g254) & (!g217) & (!g629) & (!g688)) + ((g125) & (!g164) & (g254) & (!g217) & (g629) & (!g688)) + ((g125) & (!g164) & (g254) & (g217) & (!g629) & (!g688)) + ((g125) & (!g164) & (g254) & (g217) & (g629) & (!g688)) + ((g125) & (g164) & (!g254) & (!g217) & (!g629) & (!g688)) + ((g125) & (g164) & (!g254) & (g217) & (!g629) & (!g688)) + ((g125) & (g164) & (g254) & (!g217) & (!g629) & (!g688)) + ((g125) & (g164) & (g254) & (g217) & (!g629) & (!g688)));
	assign g690 = (((!g683) & (!g685) & (!g686) & (sk[80]) & (!g687) & (g689)) + ((!g683) & (!g685) & (g686) & (!sk[80]) & (!g687) & (g689)) + ((!g683) & (!g685) & (g686) & (!sk[80]) & (g687) & (!g689)) + ((!g683) & (!g685) & (g686) & (!sk[80]) & (g687) & (g689)) + ((!g683) & (g685) & (!g686) & (!sk[80]) & (!g687) & (!g689)) + ((!g683) & (g685) & (!g686) & (!sk[80]) & (!g687) & (g689)) + ((!g683) & (g685) & (!g686) & (!sk[80]) & (g687) & (!g689)) + ((!g683) & (g685) & (!g686) & (!sk[80]) & (g687) & (g689)) + ((!g683) & (g685) & (g686) & (!sk[80]) & (!g687) & (!g689)) + ((!g683) & (g685) & (g686) & (!sk[80]) & (!g687) & (g689)) + ((!g683) & (g685) & (g686) & (!sk[80]) & (g687) & (!g689)) + ((!g683) & (g685) & (g686) & (!sk[80]) & (g687) & (g689)) + ((g683) & (!g685) & (g686) & (!sk[80]) & (!g687) & (g689)) + ((g683) & (!g685) & (g686) & (!sk[80]) & (g687) & (!g689)) + ((g683) & (!g685) & (g686) & (!sk[80]) & (g687) & (g689)) + ((g683) & (g685) & (!g686) & (!sk[80]) & (!g687) & (!g689)) + ((g683) & (g685) & (!g686) & (!sk[80]) & (!g687) & (g689)) + ((g683) & (g685) & (!g686) & (!sk[80]) & (g687) & (!g689)) + ((g683) & (g685) & (!g686) & (!sk[80]) & (g687) & (g689)) + ((g683) & (g685) & (g686) & (!sk[80]) & (!g687) & (!g689)) + ((g683) & (g685) & (g686) & (!sk[80]) & (!g687) & (g689)) + ((g683) & (g685) & (g686) & (!sk[80]) & (g687) & (!g689)) + ((g683) & (g685) & (g686) & (!sk[80]) & (g687) & (g689)));
	assign g691 = (((g676) & (!g678) & (!g679) & (!g680) & (g1457) & (g690)));
	assign g692 = (((!g30) & (g42) & (g118) & (!g113) & (!g460) & (!g629)) + ((!g30) & (g42) & (g118) & (!g113) & (!g460) & (g629)) + ((g30) & (!g42) & (g118) & (!g113) & (!g460) & (g629)) + ((g30) & (!g42) & (g118) & (!g113) & (g460) & (g629)) + ((g30) & (!g42) & (g118) & (g113) & (!g460) & (g629)) + ((g30) & (!g42) & (g118) & (g113) & (g460) & (g629)) + ((g30) & (g42) & (g118) & (!g113) & (!g460) & (!g629)) + ((g30) & (g42) & (g118) & (!g113) & (!g460) & (g629)) + ((g30) & (g42) & (g118) & (!g113) & (g460) & (g629)) + ((g30) & (g42) & (g118) & (g113) & (!g460) & (g629)) + ((g30) & (g42) & (g118) & (g113) & (g460) & (g629)));
	assign g693 = (((!i_12_) & (i_13_) & (!i_14_) & (g88) & (!g392) & (g407)) + ((!i_12_) & (i_13_) & (!i_14_) & (g88) & (g392) & (g407)) + ((i_12_) & (i_13_) & (!i_14_) & (g88) & (g392) & (!g407)) + ((i_12_) & (i_13_) & (!i_14_) & (g88) & (g392) & (g407)));
	assign g694 = (((!g131) & (!g624) & (!g625) & (sk[84]) & (!g630)) + ((!g131) & (!g624) & (!g625) & (sk[84]) & (g630)) + ((!g131) & (!g624) & (g625) & (!sk[84]) & (!g630)) + ((!g131) & (!g624) & (g625) & (!sk[84]) & (g630)) + ((!g131) & (!g624) & (g625) & (sk[84]) & (!g630)) + ((!g131) & (!g624) & (g625) & (sk[84]) & (g630)) + ((!g131) & (g624) & (!g625) & (sk[84]) & (g630)) + ((!g131) & (g624) & (g625) & (!sk[84]) & (!g630)) + ((!g131) & (g624) & (g625) & (!sk[84]) & (g630)) + ((!g131) & (g624) & (g625) & (sk[84]) & (!g630)) + ((!g131) & (g624) & (g625) & (sk[84]) & (g630)) + ((g131) & (!g624) & (g625) & (!sk[84]) & (!g630)) + ((g131) & (!g624) & (g625) & (!sk[84]) & (g630)) + ((g131) & (g624) & (g625) & (!sk[84]) & (!g630)) + ((g131) & (g624) & (g625) & (!sk[84]) & (g630)));
	assign g695 = (((!g17) & (!g19) & (!sk[85]) & (g125) & (!g694)) + ((!g17) & (!g19) & (!sk[85]) & (g125) & (g694)) + ((!g17) & (!g19) & (sk[85]) & (!g125) & (!g694)) + ((!g17) & (!g19) & (sk[85]) & (g125) & (!g694)) + ((!g17) & (g19) & (!sk[85]) & (g125) & (!g694)) + ((!g17) & (g19) & (!sk[85]) & (g125) & (g694)) + ((!g17) & (g19) & (sk[85]) & (!g125) & (!g694)) + ((!g17) & (g19) & (sk[85]) & (g125) & (!g694)) + ((g17) & (!g19) & (!sk[85]) & (g125) & (!g694)) + ((g17) & (!g19) & (!sk[85]) & (g125) & (g694)) + ((g17) & (!g19) & (sk[85]) & (!g125) & (!g694)) + ((g17) & (!g19) & (sk[85]) & (g125) & (!g694)) + ((g17) & (g19) & (!sk[85]) & (g125) & (!g694)) + ((g17) & (g19) & (!sk[85]) & (g125) & (g694)) + ((g17) & (g19) & (sk[85]) & (!g125) & (!g694)));
	assign g696 = (((!g19) & (!g69) & (!g352) & (!g692) & (!g693) & (g695)) + ((!g19) & (!g69) & (g352) & (!g692) & (!g693) & (g695)) + ((!g19) & (g69) & (!g352) & (!g692) & (!g693) & (g695)) + ((!g19) & (g69) & (g352) & (!g692) & (!g693) & (g695)) + ((g19) & (!g69) & (!g352) & (!g692) & (!g693) & (g695)) + ((g19) & (!g69) & (g352) & (!g692) & (!g693) & (g695)) + ((g19) & (g69) & (g352) & (!g692) & (!g693) & (g695)));
	assign g697 = (((g633) & (g639) & (g644) & (g672) & (g691) & (g696)));
	assign g698 = (((!sk[88]) & (!g355) & (!g35) & (g555)) + ((!sk[88]) & (!g355) & (g35) & (!g555)) + ((!sk[88]) & (!g355) & (g35) & (g555)) + ((!sk[88]) & (g355) & (!g35) & (g555)) + ((!sk[88]) & (g355) & (g35) & (!g555)) + ((!sk[88]) & (g355) & (g35) & (g555)) + ((sk[88]) & (!g355) & (!g35) & (!g555)) + ((sk[88]) & (!g355) & (g35) & (!g555)) + ((sk[88]) & (g355) & (!g35) & (!g555)));
	assign g699 = (((!g4) & (sk[89]) & (!g81)) + ((!g4) & (sk[89]) & (g81)) + ((g4) & (!sk[89]) & (!g81)) + ((g4) & (!sk[89]) & (g81)) + ((g4) & (sk[89]) & (!g81)));
	assign g700 = (((!g19) & (sk[90]) & (!g83)) + ((!g19) & (sk[90]) & (g83)) + ((g19) & (!sk[90]) & (!g83)) + ((g19) & (!sk[90]) & (g83)) + ((g19) & (sk[90]) & (!g83)));
	assign g701 = (((!g4) & (!sk[91]) & (!g69) & (g91) & (!g668)) + ((!g4) & (!sk[91]) & (!g69) & (g91) & (g668)) + ((!g4) & (!sk[91]) & (g69) & (g91) & (!g668)) + ((!g4) & (!sk[91]) & (g69) & (g91) & (g668)) + ((!g4) & (sk[91]) & (!g69) & (!g91) & (!g668)) + ((!g4) & (sk[91]) & (!g69) & (g91) & (!g668)) + ((!g4) & (sk[91]) & (g69) & (!g91) & (!g668)) + ((!g4) & (sk[91]) & (g69) & (g91) & (!g668)) + ((g4) & (!sk[91]) & (!g69) & (g91) & (!g668)) + ((g4) & (!sk[91]) & (!g69) & (g91) & (g668)) + ((g4) & (!sk[91]) & (g69) & (g91) & (!g668)) + ((g4) & (!sk[91]) & (g69) & (g91) & (g668)) + ((g4) & (sk[91]) & (!g69) & (g91) & (!g668)));
	assign g702 = (((!g634) & (!g37) & (!sk[92]) & (g75) & (!g654) & (g668)) + ((!g634) & (!g37) & (!sk[92]) & (g75) & (g654) & (!g668)) + ((!g634) & (!g37) & (!sk[92]) & (g75) & (g654) & (g668)) + ((!g634) & (!g37) & (sk[92]) & (!g75) & (!g654) & (!g668)) + ((!g634) & (!g37) & (sk[92]) & (!g75) & (!g654) & (g668)) + ((!g634) & (!g37) & (sk[92]) & (!g75) & (g654) & (!g668)) + ((!g634) & (!g37) & (sk[92]) & (!g75) & (g654) & (g668)) + ((!g634) & (g37) & (!sk[92]) & (!g75) & (!g654) & (!g668)) + ((!g634) & (g37) & (!sk[92]) & (!g75) & (!g654) & (g668)) + ((!g634) & (g37) & (!sk[92]) & (!g75) & (g654) & (!g668)) + ((!g634) & (g37) & (!sk[92]) & (!g75) & (g654) & (g668)) + ((!g634) & (g37) & (!sk[92]) & (g75) & (!g654) & (!g668)) + ((!g634) & (g37) & (!sk[92]) & (g75) & (!g654) & (g668)) + ((!g634) & (g37) & (!sk[92]) & (g75) & (g654) & (!g668)) + ((!g634) & (g37) & (!sk[92]) & (g75) & (g654) & (g668)) + ((!g634) & (g37) & (sk[92]) & (!g75) & (!g654) & (!g668)) + ((!g634) & (g37) & (sk[92]) & (!g75) & (!g654) & (g668)) + ((!g634) & (g37) & (sk[92]) & (!g75) & (g654) & (!g668)) + ((!g634) & (g37) & (sk[92]) & (!g75) & (g654) & (g668)) + ((g634) & (!g37) & (!sk[92]) & (g75) & (!g654) & (g668)) + ((g634) & (!g37) & (!sk[92]) & (g75) & (g654) & (!g668)) + ((g634) & (!g37) & (!sk[92]) & (g75) & (g654) & (g668)) + ((g634) & (!g37) & (sk[92]) & (!g75) & (!g654) & (!g668)) + ((g634) & (!g37) & (sk[92]) & (!g75) & (!g654) & (g668)) + ((g634) & (!g37) & (sk[92]) & (!g75) & (g654) & (!g668)) + ((g634) & (!g37) & (sk[92]) & (!g75) & (g654) & (g668)) + ((g634) & (g37) & (!sk[92]) & (!g75) & (!g654) & (!g668)) + ((g634) & (g37) & (!sk[92]) & (!g75) & (!g654) & (g668)) + ((g634) & (g37) & (!sk[92]) & (!g75) & (g654) & (!g668)) + ((g634) & (g37) & (!sk[92]) & (!g75) & (g654) & (g668)) + ((g634) & (g37) & (!sk[92]) & (g75) & (!g654) & (!g668)) + ((g634) & (g37) & (!sk[92]) & (g75) & (!g654) & (g668)) + ((g634) & (g37) & (!sk[92]) & (g75) & (g654) & (!g668)) + ((g634) & (g37) & (!sk[92]) & (g75) & (g654) & (g668)) + ((g634) & (g37) & (sk[92]) & (!g75) & (!g654) & (g668)) + ((g634) & (g37) & (sk[92]) & (!g75) & (g654) & (!g668)) + ((g634) & (g37) & (sk[92]) & (!g75) & (g654) & (g668)));
	assign g703 = (((!g4) & (sk[93]) & (!g88)) + ((!g4) & (sk[93]) & (g88)) + ((g4) & (!sk[93]) & (!g88)) + ((g4) & (!sk[93]) & (g88)) + ((g4) & (sk[93]) & (!g88)));
	assign g704 = (((!i_8_) & (g73) & (!g651) & (!g699) & (!g648) & (!g703)) + ((!i_8_) & (g73) & (!g651) & (!g699) & (!g648) & (g703)) + ((!i_8_) & (g73) & (!g651) & (!g699) & (g648) & (!g703)) + ((!i_8_) & (g73) & (!g651) & (!g699) & (g648) & (g703)) + ((!i_8_) & (g73) & (!g651) & (g699) & (!g648) & (!g703)) + ((!i_8_) & (g73) & (!g651) & (g699) & (g648) & (!g703)) + ((!i_8_) & (g73) & (!g651) & (g699) & (g648) & (g703)) + ((!i_8_) & (g73) & (g651) & (!g699) & (!g648) & (!g703)) + ((!i_8_) & (g73) & (g651) & (!g699) & (!g648) & (g703)) + ((!i_8_) & (g73) & (g651) & (!g699) & (g648) & (!g703)) + ((!i_8_) & (g73) & (g651) & (!g699) & (g648) & (g703)) + ((!i_8_) & (g73) & (g651) & (g699) & (!g648) & (!g703)) + ((!i_8_) & (g73) & (g651) & (g699) & (!g648) & (g703)) + ((!i_8_) & (g73) & (g651) & (g699) & (g648) & (!g703)) + ((!i_8_) & (g73) & (g651) & (g699) & (g648) & (g703)) + ((i_8_) & (g73) & (!g651) & (!g699) & (g648) & (!g703)) + ((i_8_) & (g73) & (!g651) & (!g699) & (g648) & (g703)) + ((i_8_) & (g73) & (!g651) & (g699) & (g648) & (!g703)) + ((i_8_) & (g73) & (!g651) & (g699) & (g648) & (g703)) + ((i_8_) & (g73) & (g651) & (!g699) & (g648) & (!g703)) + ((i_8_) & (g73) & (g651) & (!g699) & (g648) & (g703)) + ((i_8_) & (g73) & (g651) & (g699) & (g648) & (!g703)) + ((i_8_) & (g73) & (g651) & (g699) & (g648) & (g703)));
	assign g705 = (((!g18) & (!g33) & (!sk[95]) & (g73)) + ((!g18) & (g33) & (!sk[95]) & (!g73)) + ((!g18) & (g33) & (!sk[95]) & (g73)) + ((!g18) & (g33) & (sk[95]) & (g73)) + ((g18) & (!g33) & (!sk[95]) & (g73)) + ((g18) & (!g33) & (sk[95]) & (g73)) + ((g18) & (g33) & (!sk[95]) & (!g73)) + ((g18) & (g33) & (!sk[95]) & (g73)) + ((g18) & (g33) & (sk[95]) & (g73)));
	assign g706 = (((!g21) & (!g23) & (!sk[96]) & (g74) & (!g704) & (g705)) + ((!g21) & (!g23) & (!sk[96]) & (g74) & (g704) & (!g705)) + ((!g21) & (!g23) & (!sk[96]) & (g74) & (g704) & (g705)) + ((!g21) & (!g23) & (sk[96]) & (!g74) & (!g704) & (!g705)) + ((!g21) & (g23) & (!sk[96]) & (!g74) & (!g704) & (!g705)) + ((!g21) & (g23) & (!sk[96]) & (!g74) & (!g704) & (g705)) + ((!g21) & (g23) & (!sk[96]) & (!g74) & (g704) & (!g705)) + ((!g21) & (g23) & (!sk[96]) & (!g74) & (g704) & (g705)) + ((!g21) & (g23) & (!sk[96]) & (g74) & (!g704) & (!g705)) + ((!g21) & (g23) & (!sk[96]) & (g74) & (!g704) & (g705)) + ((!g21) & (g23) & (!sk[96]) & (g74) & (g704) & (!g705)) + ((!g21) & (g23) & (!sk[96]) & (g74) & (g704) & (g705)) + ((!g21) & (g23) & (sk[96]) & (!g74) & (!g704) & (!g705)) + ((!g21) & (g23) & (sk[96]) & (g74) & (!g704) & (!g705)) + ((g21) & (!g23) & (!sk[96]) & (g74) & (!g704) & (g705)) + ((g21) & (!g23) & (!sk[96]) & (g74) & (g704) & (!g705)) + ((g21) & (!g23) & (!sk[96]) & (g74) & (g704) & (g705)) + ((g21) & (!g23) & (sk[96]) & (!g74) & (!g704) & (!g705)) + ((g21) & (g23) & (!sk[96]) & (!g74) & (!g704) & (!g705)) + ((g21) & (g23) & (!sk[96]) & (!g74) & (!g704) & (g705)) + ((g21) & (g23) & (!sk[96]) & (!g74) & (g704) & (!g705)) + ((g21) & (g23) & (!sk[96]) & (!g74) & (g704) & (g705)) + ((g21) & (g23) & (!sk[96]) & (g74) & (!g704) & (!g705)) + ((g21) & (g23) & (!sk[96]) & (g74) & (!g704) & (g705)) + ((g21) & (g23) & (!sk[96]) & (g74) & (g704) & (!g705)) + ((g21) & (g23) & (!sk[96]) & (g74) & (g704) & (g705)) + ((g21) & (g23) & (sk[96]) & (!g74) & (!g704) & (!g705)));
	assign g707 = (((!g21) & (!g23) & (g75) & (g1531) & (!g702) & (g706)) + ((!g21) & (g23) & (!g75) & (g1531) & (!g702) & (g706)) + ((!g21) & (g23) & (g75) & (g1531) & (!g702) & (g706)) + ((g21) & (!g23) & (g75) & (g1531) & (!g702) & (g706)) + ((g21) & (g23) & (g75) & (g1531) & (!g702) & (g706)));
	assign g708 = (((!sk[98]) & (!i_8_) & (!g73) & (g108) & (!g309)) + ((!sk[98]) & (!i_8_) & (!g73) & (g108) & (g309)) + ((!sk[98]) & (!i_8_) & (g73) & (g108) & (!g309)) + ((!sk[98]) & (!i_8_) & (g73) & (g108) & (g309)) + ((!sk[98]) & (i_8_) & (!g73) & (g108) & (!g309)) + ((!sk[98]) & (i_8_) & (!g73) & (g108) & (g309)) + ((!sk[98]) & (i_8_) & (g73) & (g108) & (!g309)) + ((!sk[98]) & (i_8_) & (g73) & (g108) & (g309)) + ((sk[98]) & (i_8_) & (g73) & (!g108) & (g309)) + ((sk[98]) & (i_8_) & (g73) & (g108) & (!g309)) + ((sk[98]) & (i_8_) & (g73) & (g108) & (g309)));
	assign g709 = (((!g75) & (!g486) & (!sk[99]) & (g708)) + ((!g75) & (!g486) & (sk[99]) & (!g708)) + ((!g75) & (g486) & (!sk[99]) & (!g708)) + ((!g75) & (g486) & (!sk[99]) & (g708)) + ((g75) & (!g486) & (!sk[99]) & (g708)) + ((g75) & (!g486) & (sk[99]) & (!g708)) + ((g75) & (g486) & (!sk[99]) & (!g708)) + ((g75) & (g486) & (!sk[99]) & (g708)) + ((g75) & (g486) & (sk[99]) & (!g708)));
	assign g710 = (((!sk[100]) & (!g355) & (!g35) & (g75) & (!g555)) + ((!sk[100]) & (!g355) & (!g35) & (g75) & (g555)) + ((!sk[100]) & (!g355) & (g35) & (g75) & (!g555)) + ((!sk[100]) & (!g355) & (g35) & (g75) & (g555)) + ((!sk[100]) & (g355) & (!g35) & (g75) & (!g555)) + ((!sk[100]) & (g355) & (!g35) & (g75) & (g555)) + ((!sk[100]) & (g355) & (g35) & (g75) & (!g555)) + ((!sk[100]) & (g355) & (g35) & (g75) & (g555)) + ((sk[100]) & (!g355) & (!g35) & (!g75) & (g555)) + ((sk[100]) & (!g355) & (g35) & (!g75) & (g555)) + ((sk[100]) & (g355) & (!g35) & (!g75) & (g555)) + ((sk[100]) & (g355) & (g35) & (!g75) & (!g555)) + ((sk[100]) & (g355) & (g35) & (!g75) & (g555)));
	assign g711 = (((!g74) & (!g698) & (g196) & (g707) & (g709) & (!g710)) + ((!g74) & (g698) & (g196) & (g707) & (g709) & (!g710)) + ((g74) & (g698) & (g196) & (g707) & (g709) & (!g710)));
	assign g712 = (((!sk[102]) & (!g119) & (!g254) & (g668)) + ((!sk[102]) & (!g119) & (g254) & (!g668)) + ((!sk[102]) & (!g119) & (g254) & (g668)) + ((!sk[102]) & (g119) & (!g254) & (g668)) + ((!sk[102]) & (g119) & (g254) & (!g668)) + ((!sk[102]) & (g119) & (g254) & (g668)) + ((sk[102]) & (!g119) & (!g254) & (g668)) + ((sk[102]) & (g119) & (!g254) & (g668)) + ((sk[102]) & (g119) & (g254) & (g668)));
	assign g713 = (((!sk[103]) & (!g123) & (!g119) & (g654)) + ((!sk[103]) & (!g123) & (g119) & (!g654)) + ((!sk[103]) & (!g123) & (g119) & (g654)) + ((!sk[103]) & (g123) & (!g119) & (g654)) + ((!sk[103]) & (g123) & (g119) & (!g654)) + ((!sk[103]) & (g123) & (g119) & (g654)) + ((sk[103]) & (!g123) & (!g119) & (g654)) + ((sk[103]) & (!g123) & (g119) & (g654)) + ((sk[103]) & (g123) & (g119) & (g654)));
	assign g714 = (((!sk[104]) & (!g105) & (!g121) & (g654)) + ((!sk[104]) & (!g105) & (g121) & (!g654)) + ((!sk[104]) & (!g105) & (g121) & (g654)) + ((!sk[104]) & (g105) & (!g121) & (g654)) + ((!sk[104]) & (g105) & (g121) & (!g654)) + ((!sk[104]) & (g105) & (g121) & (g654)) + ((sk[104]) & (!g105) & (!g121) & (g654)) + ((sk[104]) & (!g105) & (g121) & (g654)) + ((sk[104]) & (g105) & (g121) & (g654)));
	assign g715 = (((!sk[105]) & (!g19) & (!g126) & (g122) & (!g684)) + ((!sk[105]) & (!g19) & (!g126) & (g122) & (g684)) + ((!sk[105]) & (!g19) & (g126) & (g122) & (!g684)) + ((!sk[105]) & (!g19) & (g126) & (g122) & (g684)) + ((!sk[105]) & (g19) & (!g126) & (g122) & (!g684)) + ((!sk[105]) & (g19) & (!g126) & (g122) & (g684)) + ((!sk[105]) & (g19) & (g126) & (g122) & (!g684)) + ((!sk[105]) & (g19) & (g126) & (g122) & (g684)) + ((sk[105]) & (!g19) & (!g126) & (g122) & (!g684)) + ((sk[105]) & (!g19) & (g126) & (g122) & (!g684)) + ((sk[105]) & (g19) & (!g126) & (g122) & (!g684)) + ((sk[105]) & (g19) & (!g126) & (g122) & (g684)) + ((sk[105]) & (g19) & (g126) & (g122) & (!g684)));
	assign g716 = (((!g3) & (!g19) & (g125) & (!g126) & (!sk[106]) & (g121)) + ((!g3) & (!g19) & (g125) & (g126) & (!sk[106]) & (!g121)) + ((!g3) & (!g19) & (g125) & (g126) & (!sk[106]) & (g121)) + ((!g3) & (g19) & (!g125) & (!g126) & (!sk[106]) & (!g121)) + ((!g3) & (g19) & (!g125) & (!g126) & (!sk[106]) & (g121)) + ((!g3) & (g19) & (!g125) & (g126) & (!sk[106]) & (!g121)) + ((!g3) & (g19) & (!g125) & (g126) & (!sk[106]) & (g121)) + ((!g3) & (g19) & (g125) & (!g126) & (!sk[106]) & (!g121)) + ((!g3) & (g19) & (g125) & (!g126) & (!sk[106]) & (g121)) + ((!g3) & (g19) & (g125) & (!g126) & (sk[106]) & (!g121)) + ((!g3) & (g19) & (g125) & (!g126) & (sk[106]) & (g121)) + ((!g3) & (g19) & (g125) & (g126) & (!sk[106]) & (!g121)) + ((!g3) & (g19) & (g125) & (g126) & (!sk[106]) & (g121)) + ((g3) & (!g19) & (g125) & (!g126) & (!sk[106]) & (g121)) + ((g3) & (!g19) & (g125) & (g126) & (!sk[106]) & (!g121)) + ((g3) & (!g19) & (g125) & (g126) & (!sk[106]) & (g121)) + ((g3) & (g19) & (!g125) & (!g126) & (!sk[106]) & (!g121)) + ((g3) & (g19) & (!g125) & (!g126) & (!sk[106]) & (g121)) + ((g3) & (g19) & (!g125) & (!g126) & (sk[106]) & (g121)) + ((g3) & (g19) & (!g125) & (g126) & (!sk[106]) & (!g121)) + ((g3) & (g19) & (!g125) & (g126) & (!sk[106]) & (g121)) + ((g3) & (g19) & (!g125) & (g126) & (sk[106]) & (g121)) + ((g3) & (g19) & (g125) & (!g126) & (!sk[106]) & (!g121)) + ((g3) & (g19) & (g125) & (!g126) & (!sk[106]) & (g121)) + ((g3) & (g19) & (g125) & (!g126) & (sk[106]) & (!g121)) + ((g3) & (g19) & (g125) & (!g126) & (sk[106]) & (g121)) + ((g3) & (g19) & (g125) & (g126) & (!sk[106]) & (!g121)) + ((g3) & (g19) & (g125) & (g126) & (!sk[106]) & (g121)) + ((g3) & (g19) & (g125) & (g126) & (sk[106]) & (!g121)) + ((g3) & (g19) & (g125) & (g126) & (sk[106]) & (g121)));
	assign g717 = (((!g19) & (!g75) & (!g126) & (!g715) & (sk[107]) & (!g716)) + ((!g19) & (!g75) & (g126) & (!g715) & (!sk[107]) & (g716)) + ((!g19) & (!g75) & (g126) & (!g715) & (sk[107]) & (!g716)) + ((!g19) & (!g75) & (g126) & (g715) & (!sk[107]) & (!g716)) + ((!g19) & (!g75) & (g126) & (g715) & (!sk[107]) & (g716)) + ((!g19) & (g75) & (!g126) & (!g715) & (!sk[107]) & (!g716)) + ((!g19) & (g75) & (!g126) & (!g715) & (!sk[107]) & (g716)) + ((!g19) & (g75) & (!g126) & (!g715) & (sk[107]) & (!g716)) + ((!g19) & (g75) & (!g126) & (g715) & (!sk[107]) & (!g716)) + ((!g19) & (g75) & (!g126) & (g715) & (!sk[107]) & (g716)) + ((!g19) & (g75) & (g126) & (!g715) & (!sk[107]) & (!g716)) + ((!g19) & (g75) & (g126) & (!g715) & (!sk[107]) & (g716)) + ((!g19) & (g75) & (g126) & (!g715) & (sk[107]) & (!g716)) + ((!g19) & (g75) & (g126) & (g715) & (!sk[107]) & (!g716)) + ((!g19) & (g75) & (g126) & (g715) & (!sk[107]) & (g716)) + ((g19) & (!g75) & (g126) & (!g715) & (!sk[107]) & (g716)) + ((g19) & (!g75) & (g126) & (!g715) & (sk[107]) & (!g716)) + ((g19) & (!g75) & (g126) & (g715) & (!sk[107]) & (!g716)) + ((g19) & (!g75) & (g126) & (g715) & (!sk[107]) & (g716)) + ((g19) & (g75) & (!g126) & (!g715) & (!sk[107]) & (!g716)) + ((g19) & (g75) & (!g126) & (!g715) & (!sk[107]) & (g716)) + ((g19) & (g75) & (!g126) & (!g715) & (sk[107]) & (!g716)) + ((g19) & (g75) & (!g126) & (g715) & (!sk[107]) & (!g716)) + ((g19) & (g75) & (!g126) & (g715) & (!sk[107]) & (g716)) + ((g19) & (g75) & (g126) & (!g715) & (!sk[107]) & (!g716)) + ((g19) & (g75) & (g126) & (!g715) & (!sk[107]) & (g716)) + ((g19) & (g75) & (g126) & (!g715) & (sk[107]) & (!g716)) + ((g19) & (g75) & (g126) & (g715) & (!sk[107]) & (!g716)) + ((g19) & (g75) & (g126) & (g715) & (!sk[107]) & (g716)));
	assign g718 = (((!sk[108]) & (!g125) & (!g226) & (g684) & (!g668)) + ((!sk[108]) & (!g125) & (!g226) & (g684) & (g668)) + ((!sk[108]) & (!g125) & (g226) & (g684) & (!g668)) + ((!sk[108]) & (!g125) & (g226) & (g684) & (g668)) + ((!sk[108]) & (g125) & (!g226) & (g684) & (!g668)) + ((!sk[108]) & (g125) & (!g226) & (g684) & (g668)) + ((!sk[108]) & (g125) & (g226) & (g684) & (!g668)) + ((!sk[108]) & (g125) & (g226) & (g684) & (g668)) + ((sk[108]) & (!g125) & (!g226) & (!g684) & (g668)) + ((sk[108]) & (!g125) & (!g226) & (g684) & (g668)) + ((sk[108]) & (g125) & (!g226) & (!g684) & (!g668)) + ((sk[108]) & (g125) & (!g226) & (!g684) & (g668)) + ((sk[108]) & (g125) & (!g226) & (g684) & (g668)) + ((sk[108]) & (g125) & (g226) & (!g684) & (!g668)) + ((sk[108]) & (g125) & (g226) & (!g684) & (g668)));
	assign g719 = (((!sk[109]) & (!g70) & (!g270) & (g511)) + ((!sk[109]) & (!g70) & (g270) & (!g511)) + ((!sk[109]) & (!g70) & (g270) & (g511)) + ((!sk[109]) & (g70) & (!g270) & (g511)) + ((!sk[109]) & (g70) & (g270) & (!g511)) + ((!sk[109]) & (g70) & (g270) & (g511)) + ((sk[109]) & (!g70) & (!g270) & (!g511)));
	assign g720 = (((!g77) & (!g719) & (!sk[110]) & (g654)) + ((!g77) & (g719) & (!sk[110]) & (!g654)) + ((!g77) & (g719) & (!sk[110]) & (g654)) + ((!g77) & (g719) & (sk[110]) & (!g654)) + ((g77) & (!g719) & (!sk[110]) & (g654)) + ((g77) & (g719) & (!sk[110]) & (!g654)) + ((g77) & (g719) & (!sk[110]) & (g654)));
	assign g721 = (((i_8_) & (!i_6_) & (!i_7_) & (g120) & (g508) & (!g720)) + ((i_8_) & (!i_6_) & (!i_7_) & (g120) & (g508) & (g720)) + ((i_8_) & (i_6_) & (!i_7_) & (g120) & (!g508) & (!g720)));
	assign g722 = (((!g712) & (!g713) & (!g714) & (g717) & (!g718) & (!g721)));
	assign g723 = (((g81) & (!sk[113]) & (!g507)) + ((g81) & (!sk[113]) & (g507)) + ((g81) & (sk[113]) & (g507)));
	assign g724 = (((!i_9_) & (!i_10_) & (!g123) & (!g315) & (!g408) & (g723)) + ((!i_9_) & (!i_10_) & (!g123) & (!g315) & (g408) & (g723)) + ((!i_9_) & (!i_10_) & (!g123) & (g315) & (!g408) & (g723)) + ((!i_9_) & (!i_10_) & (!g123) & (g315) & (g408) & (g723)) + ((!i_9_) & (i_10_) & (!g123) & (!g315) & (!g408) & (g723)) + ((!i_9_) & (i_10_) & (!g123) & (!g315) & (g408) & (g723)) + ((!i_9_) & (i_10_) & (!g123) & (g315) & (!g408) & (!g723)) + ((!i_9_) & (i_10_) & (!g123) & (g315) & (!g408) & (g723)) + ((!i_9_) & (i_10_) & (!g123) & (g315) & (g408) & (g723)) + ((!i_9_) & (i_10_) & (g123) & (g315) & (!g408) & (!g723)) + ((!i_9_) & (i_10_) & (g123) & (g315) & (!g408) & (g723)) + ((i_9_) & (!i_10_) & (!g123) & (!g315) & (!g408) & (g723)) + ((i_9_) & (!i_10_) & (!g123) & (!g315) & (g408) & (g723)) + ((i_9_) & (!i_10_) & (!g123) & (g315) & (!g408) & (g723)) + ((i_9_) & (!i_10_) & (!g123) & (g315) & (g408) & (g723)) + ((i_9_) & (i_10_) & (!g123) & (!g315) & (!g408) & (g723)) + ((i_9_) & (i_10_) & (!g123) & (!g315) & (g408) & (g723)) + ((i_9_) & (i_10_) & (!g123) & (g315) & (!g408) & (g723)) + ((i_9_) & (i_10_) & (!g123) & (g315) & (g408) & (g723)));
	assign g725 = (((!g17) & (!g19) & (!sk[115]) & (g357)) + ((!g17) & (!g19) & (sk[115]) & (!g357)) + ((!g17) & (g19) & (!sk[115]) & (!g357)) + ((!g17) & (g19) & (!sk[115]) & (g357)) + ((!g17) & (g19) & (sk[115]) & (!g357)) + ((g17) & (!g19) & (!sk[115]) & (g357)) + ((g17) & (!g19) & (sk[115]) & (!g357)) + ((g17) & (g19) & (!sk[115]) & (!g357)) + ((g17) & (g19) & (!sk[115]) & (g357)));
	assign g726 = (((!g121) & (!g434) & (g341) & (!sk[116]) & (!g725)) + ((!g121) & (!g434) & (g341) & (!sk[116]) & (g725)) + ((!g121) & (g434) & (!g341) & (sk[116]) & (!g725)) + ((!g121) & (g434) & (g341) & (!sk[116]) & (!g725)) + ((!g121) & (g434) & (g341) & (!sk[116]) & (g725)) + ((!g121) & (g434) & (g341) & (sk[116]) & (!g725)) + ((g121) & (!g434) & (!g341) & (sk[116]) & (!g725)) + ((g121) & (!g434) & (!g341) & (sk[116]) & (g725)) + ((g121) & (!g434) & (g341) & (!sk[116]) & (!g725)) + ((g121) & (!g434) & (g341) & (!sk[116]) & (g725)) + ((g121) & (g434) & (!g341) & (sk[116]) & (!g725)) + ((g121) & (g434) & (!g341) & (sk[116]) & (g725)) + ((g121) & (g434) & (g341) & (!sk[116]) & (!g725)) + ((g121) & (g434) & (g341) & (!sk[116]) & (g725)) + ((g121) & (g434) & (g341) & (sk[116]) & (!g725)));
	assign g727 = (((!g167) & (!g144) & (!g334) & (!g624) & (!g724) & (!g726)) + ((!g167) & (!g144) & (!g334) & (g624) & (!g724) & (!g726)) + ((!g167) & (!g144) & (g334) & (!g624) & (!g724) & (!g726)) + ((!g167) & (!g144) & (g334) & (g624) & (!g724) & (!g726)) + ((!g167) & (g144) & (g334) & (!g624) & (!g724) & (!g726)) + ((!g167) & (g144) & (g334) & (g624) & (!g724) & (!g726)) + ((g167) & (!g144) & (!g334) & (g624) & (!g724) & (!g726)) + ((g167) & (!g144) & (g334) & (g624) & (!g724) & (!g726)) + ((g167) & (g144) & (g334) & (g624) & (!g724) & (!g726)));
	assign g728 = (((!sk[118]) & (g355) & (!g35)) + ((!sk[118]) & (g355) & (g35)) + ((sk[118]) & (g355) & (g35)));
	assign g729 = (((!g355) & (!sk[119]) & (!g107) & (g486)) + ((!g355) & (!sk[119]) & (g107) & (!g486)) + ((!g355) & (!sk[119]) & (g107) & (g486)) + ((!g355) & (sk[119]) & (!g107) & (!g486)) + ((!g355) & (sk[119]) & (g107) & (!g486)) + ((g355) & (!sk[119]) & (!g107) & (g486)) + ((g355) & (!sk[119]) & (g107) & (!g486)) + ((g355) & (!sk[119]) & (g107) & (g486)) + ((g355) & (sk[119]) & (g107) & (!g486)));
	assign g730 = (((!sk[120]) & (!i_13_) & (!i_14_) & (g36) & (!g625)) + ((!sk[120]) & (!i_13_) & (!i_14_) & (g36) & (g625)) + ((!sk[120]) & (!i_13_) & (i_14_) & (g36) & (!g625)) + ((!sk[120]) & (!i_13_) & (i_14_) & (g36) & (g625)) + ((!sk[120]) & (i_13_) & (!i_14_) & (g36) & (!g625)) + ((!sk[120]) & (i_13_) & (!i_14_) & (g36) & (g625)) + ((!sk[120]) & (i_13_) & (i_14_) & (g36) & (!g625)) + ((!sk[120]) & (i_13_) & (i_14_) & (g36) & (g625)) + ((sk[120]) & (!i_13_) & (!i_14_) & (!g36) & (!g625)) + ((sk[120]) & (!i_13_) & (i_14_) & (!g36) & (!g625)) + ((sk[120]) & (!i_13_) & (i_14_) & (g36) & (!g625)) + ((sk[120]) & (i_13_) & (!i_14_) & (!g36) & (!g625)) + ((sk[120]) & (i_13_) & (!i_14_) & (g36) & (!g625)) + ((sk[120]) & (i_13_) & (i_14_) & (!g36) & (!g625)) + ((sk[120]) & (i_13_) & (i_14_) & (g36) & (!g625)));
	assign g731 = (((!g125) & (!g131) & (!g728) & (!g534) & (g729) & (!g730)) + ((!g125) & (!g131) & (!g728) & (!g534) & (g729) & (g730)) + ((!g125) & (g131) & (!g728) & (!g534) & (!g729) & (!g730)) + ((!g125) & (g131) & (!g728) & (!g534) & (!g729) & (g730)) + ((!g125) & (g131) & (!g728) & (!g534) & (g729) & (!g730)) + ((!g125) & (g131) & (!g728) & (!g534) & (g729) & (g730)) + ((!g125) & (g131) & (!g728) & (g534) & (!g729) & (!g730)) + ((!g125) & (g131) & (!g728) & (g534) & (!g729) & (g730)) + ((!g125) & (g131) & (!g728) & (g534) & (g729) & (!g730)) + ((!g125) & (g131) & (!g728) & (g534) & (g729) & (g730)) + ((!g125) & (g131) & (g728) & (!g534) & (!g729) & (!g730)) + ((!g125) & (g131) & (g728) & (!g534) & (!g729) & (g730)) + ((!g125) & (g131) & (g728) & (!g534) & (g729) & (!g730)) + ((!g125) & (g131) & (g728) & (!g534) & (g729) & (g730)) + ((!g125) & (g131) & (g728) & (g534) & (!g729) & (!g730)) + ((!g125) & (g131) & (g728) & (g534) & (!g729) & (g730)) + ((!g125) & (g131) & (g728) & (g534) & (g729) & (!g730)) + ((!g125) & (g131) & (g728) & (g534) & (g729) & (g730)) + ((g125) & (!g131) & (!g728) & (!g534) & (g729) & (g730)) + ((g125) & (g131) & (!g728) & (!g534) & (!g729) & (g730)) + ((g125) & (g131) & (!g728) & (!g534) & (g729) & (g730)) + ((g125) & (g131) & (!g728) & (g534) & (!g729) & (g730)) + ((g125) & (g131) & (!g728) & (g534) & (g729) & (g730)) + ((g125) & (g131) & (g728) & (!g534) & (!g729) & (g730)) + ((g125) & (g131) & (g728) & (!g534) & (g729) & (g730)) + ((g125) & (g131) & (g728) & (g534) & (!g729) & (g730)) + ((g125) & (g131) & (g728) & (g534) & (g729) & (g730)));
	assign g732 = (((!sk[122]) & (!g21) & (!g313) & (g254) & (!g333)) + ((!sk[122]) & (!g21) & (!g313) & (g254) & (g333)) + ((!sk[122]) & (!g21) & (g313) & (g254) & (!g333)) + ((!sk[122]) & (!g21) & (g313) & (g254) & (g333)) + ((!sk[122]) & (g21) & (!g313) & (g254) & (!g333)) + ((!sk[122]) & (g21) & (!g313) & (g254) & (g333)) + ((!sk[122]) & (g21) & (g313) & (g254) & (!g333)) + ((!sk[122]) & (g21) & (g313) & (g254) & (g333)) + ((sk[122]) & (!g21) & (g313) & (!g254) & (g333)) + ((sk[122]) & (!g21) & (g313) & (g254) & (g333)) + ((sk[122]) & (g21) & (!g313) & (!g254) & (!g333)) + ((sk[122]) & (g21) & (!g313) & (!g254) & (g333)) + ((sk[122]) & (g21) & (g313) & (!g254) & (!g333)) + ((sk[122]) & (g21) & (g313) & (!g254) & (g333)) + ((sk[122]) & (g21) & (g313) & (g254) & (g333)));
	assign g733 = (((!g87) & (!g125) & (!g122) & (sk[123]) & (!g272) & (!g534)) + ((!g87) & (!g125) & (!g122) & (sk[123]) & (!g272) & (g534)) + ((!g87) & (!g125) & (!g122) & (sk[123]) & (g272) & (!g534)) + ((!g87) & (!g125) & (!g122) & (sk[123]) & (g272) & (g534)) + ((!g87) & (!g125) & (g122) & (!sk[123]) & (!g272) & (g534)) + ((!g87) & (!g125) & (g122) & (!sk[123]) & (g272) & (!g534)) + ((!g87) & (!g125) & (g122) & (!sk[123]) & (g272) & (g534)) + ((!g87) & (g125) & (!g122) & (!sk[123]) & (!g272) & (!g534)) + ((!g87) & (g125) & (!g122) & (!sk[123]) & (!g272) & (g534)) + ((!g87) & (g125) & (!g122) & (!sk[123]) & (g272) & (!g534)) + ((!g87) & (g125) & (!g122) & (!sk[123]) & (g272) & (g534)) + ((!g87) & (g125) & (g122) & (!sk[123]) & (!g272) & (!g534)) + ((!g87) & (g125) & (g122) & (!sk[123]) & (!g272) & (g534)) + ((!g87) & (g125) & (g122) & (!sk[123]) & (g272) & (!g534)) + ((!g87) & (g125) & (g122) & (!sk[123]) & (g272) & (g534)) + ((g87) & (!g125) & (!g122) & (sk[123]) & (!g272) & (!g534)) + ((g87) & (!g125) & (!g122) & (sk[123]) & (!g272) & (g534)) + ((g87) & (!g125) & (!g122) & (sk[123]) & (g272) & (!g534)) + ((g87) & (!g125) & (!g122) & (sk[123]) & (g272) & (g534)) + ((g87) & (!g125) & (g122) & (!sk[123]) & (!g272) & (g534)) + ((g87) & (!g125) & (g122) & (!sk[123]) & (g272) & (!g534)) + ((g87) & (!g125) & (g122) & (!sk[123]) & (g272) & (g534)) + ((g87) & (!g125) & (g122) & (sk[123]) & (!g272) & (!g534)) + ((g87) & (g125) & (!g122) & (!sk[123]) & (!g272) & (!g534)) + ((g87) & (g125) & (!g122) & (!sk[123]) & (!g272) & (g534)) + ((g87) & (g125) & (!g122) & (!sk[123]) & (g272) & (!g534)) + ((g87) & (g125) & (!g122) & (!sk[123]) & (g272) & (g534)) + ((g87) & (g125) & (!g122) & (sk[123]) & (!g272) & (!g534)) + ((g87) & (g125) & (g122) & (!sk[123]) & (!g272) & (!g534)) + ((g87) & (g125) & (g122) & (!sk[123]) & (!g272) & (g534)) + ((g87) & (g125) & (g122) & (!sk[123]) & (g272) & (!g534)) + ((g87) & (g125) & (g122) & (!sk[123]) & (g272) & (g534)) + ((g87) & (g125) & (g122) & (sk[123]) & (!g272) & (!g534)));
	assign g734 = (((!g161) & (!g451) & (!g732) & (sk[124]) & (g733)) + ((!g161) & (!g451) & (g732) & (!sk[124]) & (!g733)) + ((!g161) & (!g451) & (g732) & (!sk[124]) & (g733)) + ((!g161) & (g451) & (!g732) & (sk[124]) & (g733)) + ((!g161) & (g451) & (g732) & (!sk[124]) & (!g733)) + ((!g161) & (g451) & (g732) & (!sk[124]) & (g733)) + ((g161) & (!g451) & (g732) & (!sk[124]) & (!g733)) + ((g161) & (!g451) & (g732) & (!sk[124]) & (g733)) + ((g161) & (g451) & (!g732) & (sk[124]) & (g733)) + ((g161) & (g451) & (g732) & (!sk[124]) & (!g733)) + ((g161) & (g451) & (g732) & (!sk[124]) & (g733)));
	assign g735 = (((!i_12_) & (!sk[125]) & (!i_13_) & (i_14_)) + ((!i_12_) & (!sk[125]) & (i_13_) & (!i_14_)) + ((!i_12_) & (!sk[125]) & (i_13_) & (i_14_)) + ((!i_12_) & (sk[125]) & (i_13_) & (!i_14_)) + ((i_12_) & (!sk[125]) & (!i_13_) & (i_14_)) + ((i_12_) & (!sk[125]) & (i_13_) & (!i_14_)) + ((i_12_) & (!sk[125]) & (i_13_) & (i_14_)) + ((i_12_) & (sk[125]) & (!i_13_) & (!i_14_)));
	assign g736 = (((!i_9_) & (!sk[126]) & (!i_10_) & (i_15_) & (!g19)) + ((!i_9_) & (!sk[126]) & (!i_10_) & (i_15_) & (g19)) + ((!i_9_) & (!sk[126]) & (i_10_) & (i_15_) & (!g19)) + ((!i_9_) & (!sk[126]) & (i_10_) & (i_15_) & (g19)) + ((!i_9_) & (sk[126]) & (i_10_) & (!i_15_) & (g19)) + ((i_9_) & (!sk[126]) & (!i_10_) & (i_15_) & (!g19)) + ((i_9_) & (!sk[126]) & (!i_10_) & (i_15_) & (g19)) + ((i_9_) & (!sk[126]) & (i_10_) & (i_15_) & (!g19)) + ((i_9_) & (!sk[126]) & (i_10_) & (i_15_) & (g19)));
	assign g737 = (((!sk[127]) & (!g68) & (!g126) & (g508) & (!g736)) + ((!sk[127]) & (!g68) & (!g126) & (g508) & (g736)) + ((!sk[127]) & (!g68) & (g126) & (g508) & (!g736)) + ((!sk[127]) & (!g68) & (g126) & (g508) & (g736)) + ((!sk[127]) & (g68) & (!g126) & (g508) & (!g736)) + ((!sk[127]) & (g68) & (!g126) & (g508) & (g736)) + ((!sk[127]) & (g68) & (g126) & (g508) & (!g736)) + ((!sk[127]) & (g68) & (g126) & (g508) & (g736)) + ((sk[127]) & (!g68) & (g126) & (!g508) & (!g736)) + ((sk[127]) & (g68) & (!g126) & (!g508) & (!g736)) + ((sk[127]) & (g68) & (g126) & (!g508) & (!g736)));
	assign g738 = (((!g22) & (sk[0]) & (g507)) + ((g22) & (!sk[0]) & (!g507)) + ((g22) & (!sk[0]) & (g507)));
	assign g739 = (((!sk[1]) & (!g562) & (!g737) & (g738)) + ((!sk[1]) & (!g562) & (g737) & (!g738)) + ((!sk[1]) & (!g562) & (g737) & (g738)) + ((!sk[1]) & (g562) & (!g737) & (g738)) + ((!sk[1]) & (g562) & (g737) & (!g738)) + ((!sk[1]) & (g562) & (g737) & (g738)) + ((sk[1]) & (!g562) & (g737) & (!g738)));
	assign g740 = (((!sk[2]) & (!i_15_) & (!g19) & (g428) & (!g68) & (g429)) + ((!sk[2]) & (!i_15_) & (!g19) & (g428) & (g68) & (!g429)) + ((!sk[2]) & (!i_15_) & (!g19) & (g428) & (g68) & (g429)) + ((!sk[2]) & (!i_15_) & (g19) & (!g428) & (!g68) & (!g429)) + ((!sk[2]) & (!i_15_) & (g19) & (!g428) & (!g68) & (g429)) + ((!sk[2]) & (!i_15_) & (g19) & (!g428) & (g68) & (!g429)) + ((!sk[2]) & (!i_15_) & (g19) & (!g428) & (g68) & (g429)) + ((!sk[2]) & (!i_15_) & (g19) & (g428) & (!g68) & (!g429)) + ((!sk[2]) & (!i_15_) & (g19) & (g428) & (!g68) & (g429)) + ((!sk[2]) & (!i_15_) & (g19) & (g428) & (g68) & (!g429)) + ((!sk[2]) & (!i_15_) & (g19) & (g428) & (g68) & (g429)) + ((!sk[2]) & (i_15_) & (!g19) & (g428) & (!g68) & (g429)) + ((!sk[2]) & (i_15_) & (!g19) & (g428) & (g68) & (!g429)) + ((!sk[2]) & (i_15_) & (!g19) & (g428) & (g68) & (g429)) + ((!sk[2]) & (i_15_) & (g19) & (!g428) & (!g68) & (!g429)) + ((!sk[2]) & (i_15_) & (g19) & (!g428) & (!g68) & (g429)) + ((!sk[2]) & (i_15_) & (g19) & (!g428) & (g68) & (!g429)) + ((!sk[2]) & (i_15_) & (g19) & (!g428) & (g68) & (g429)) + ((!sk[2]) & (i_15_) & (g19) & (g428) & (!g68) & (!g429)) + ((!sk[2]) & (i_15_) & (g19) & (g428) & (!g68) & (g429)) + ((!sk[2]) & (i_15_) & (g19) & (g428) & (g68) & (!g429)) + ((!sk[2]) & (i_15_) & (g19) & (g428) & (g68) & (g429)) + ((sk[2]) & (!i_15_) & (!g19) & (!g428) & (!g68) & (!g429)) + ((sk[2]) & (!i_15_) & (!g19) & (!g428) & (!g68) & (g429)) + ((sk[2]) & (!i_15_) & (!g19) & (g428) & (!g68) & (g429)) + ((sk[2]) & (!i_15_) & (g19) & (!g428) & (!g68) & (!g429)) + ((sk[2]) & (!i_15_) & (g19) & (!g428) & (!g68) & (g429)) + ((sk[2]) & (!i_15_) & (g19) & (!g428) & (g68) & (g429)) + ((sk[2]) & (!i_15_) & (g19) & (g428) & (!g68) & (g429)) + ((sk[2]) & (!i_15_) & (g19) & (g428) & (g68) & (g429)));
	assign g741 = (((!g27) & (!g105) & (!g425) & (!g735) & (g739) & (!g740)) + ((!g27) & (!g105) & (!g425) & (g735) & (g739) & (!g740)) + ((!g27) & (!g105) & (g425) & (!g735) & (g739) & (!g740)) + ((!g27) & (!g105) & (g425) & (g735) & (g739) & (!g740)) + ((!g27) & (g105) & (!g425) & (!g735) & (!g739) & (!g740)) + ((!g27) & (g105) & (!g425) & (!g735) & (g739) & (!g740)) + ((!g27) & (g105) & (!g425) & (g735) & (!g739) & (!g740)) + ((!g27) & (g105) & (!g425) & (g735) & (g739) & (!g740)) + ((!g27) & (g105) & (g425) & (!g735) & (!g739) & (!g740)) + ((!g27) & (g105) & (g425) & (!g735) & (!g739) & (g740)) + ((!g27) & (g105) & (g425) & (!g735) & (g739) & (!g740)) + ((!g27) & (g105) & (g425) & (!g735) & (g739) & (g740)) + ((!g27) & (g105) & (g425) & (g735) & (!g739) & (!g740)) + ((!g27) & (g105) & (g425) & (g735) & (!g739) & (g740)) + ((!g27) & (g105) & (g425) & (g735) & (g739) & (!g740)) + ((!g27) & (g105) & (g425) & (g735) & (g739) & (g740)) + ((g27) & (!g105) & (!g425) & (!g735) & (g739) & (!g740)) + ((g27) & (!g105) & (g425) & (!g735) & (g739) & (!g740)) + ((g27) & (!g105) & (g425) & (g735) & (g739) & (!g740)) + ((g27) & (g105) & (!g425) & (!g735) & (!g739) & (!g740)) + ((g27) & (g105) & (!g425) & (!g735) & (g739) & (!g740)) + ((g27) & (g105) & (g425) & (!g735) & (!g739) & (!g740)) + ((g27) & (g105) & (g425) & (!g735) & (!g739) & (g740)) + ((g27) & (g105) & (g425) & (!g735) & (g739) & (!g740)) + ((g27) & (g105) & (g425) & (!g735) & (g739) & (g740)) + ((g27) & (g105) & (g425) & (g735) & (!g739) & (!g740)) + ((g27) & (g105) & (g425) & (g735) & (!g739) & (g740)) + ((g27) & (g105) & (g425) & (g735) & (g739) & (!g740)) + ((g27) & (g105) & (g425) & (g735) & (g739) & (g740)));
	assign g742 = (((!g126) & (!g176) & (!sk[4]) & (g642)) + ((!g126) & (g176) & (!sk[4]) & (!g642)) + ((!g126) & (g176) & (!sk[4]) & (g642)) + ((!g126) & (g176) & (sk[4]) & (!g642)) + ((g126) & (!g176) & (!sk[4]) & (g642)) + ((g126) & (!g176) & (sk[4]) & (!g642)) + ((g126) & (g176) & (!sk[4]) & (!g642)) + ((g126) & (g176) & (!sk[4]) & (g642)) + ((g126) & (g176) & (sk[4]) & (!g642)));
	assign g743 = (((!g3) & (!i_12_) & (!i_13_) & (!i_14_) & (sk[5]) & (g69)) + ((!g3) & (!i_12_) & (i_13_) & (!i_14_) & (!sk[5]) & (g69)) + ((!g3) & (!i_12_) & (i_13_) & (i_14_) & (!sk[5]) & (!g69)) + ((!g3) & (!i_12_) & (i_13_) & (i_14_) & (!sk[5]) & (g69)) + ((!g3) & (i_12_) & (!i_13_) & (!i_14_) & (!sk[5]) & (!g69)) + ((!g3) & (i_12_) & (!i_13_) & (!i_14_) & (!sk[5]) & (g69)) + ((!g3) & (i_12_) & (!i_13_) & (!i_14_) & (sk[5]) & (g69)) + ((!g3) & (i_12_) & (!i_13_) & (i_14_) & (!sk[5]) & (!g69)) + ((!g3) & (i_12_) & (!i_13_) & (i_14_) & (!sk[5]) & (g69)) + ((!g3) & (i_12_) & (i_13_) & (!i_14_) & (!sk[5]) & (!g69)) + ((!g3) & (i_12_) & (i_13_) & (!i_14_) & (!sk[5]) & (g69)) + ((!g3) & (i_12_) & (i_13_) & (!i_14_) & (sk[5]) & (g69)) + ((!g3) & (i_12_) & (i_13_) & (i_14_) & (!sk[5]) & (!g69)) + ((!g3) & (i_12_) & (i_13_) & (i_14_) & (!sk[5]) & (g69)) + ((g3) & (!i_12_) & (!i_13_) & (!i_14_) & (sk[5]) & (g69)) + ((g3) & (!i_12_) & (!i_13_) & (i_14_) & (sk[5]) & (!g69)) + ((g3) & (!i_12_) & (!i_13_) & (i_14_) & (sk[5]) & (g69)) + ((g3) & (!i_12_) & (i_13_) & (!i_14_) & (!sk[5]) & (g69)) + ((g3) & (!i_12_) & (i_13_) & (i_14_) & (!sk[5]) & (!g69)) + ((g3) & (!i_12_) & (i_13_) & (i_14_) & (!sk[5]) & (g69)) + ((g3) & (!i_12_) & (i_13_) & (i_14_) & (sk[5]) & (!g69)) + ((g3) & (!i_12_) & (i_13_) & (i_14_) & (sk[5]) & (g69)) + ((g3) & (i_12_) & (!i_13_) & (!i_14_) & (!sk[5]) & (!g69)) + ((g3) & (i_12_) & (!i_13_) & (!i_14_) & (!sk[5]) & (g69)) + ((g3) & (i_12_) & (!i_13_) & (!i_14_) & (sk[5]) & (g69)) + ((g3) & (i_12_) & (!i_13_) & (i_14_) & (!sk[5]) & (!g69)) + ((g3) & (i_12_) & (!i_13_) & (i_14_) & (!sk[5]) & (g69)) + ((g3) & (i_12_) & (i_13_) & (!i_14_) & (!sk[5]) & (!g69)) + ((g3) & (i_12_) & (i_13_) & (!i_14_) & (!sk[5]) & (g69)) + ((g3) & (i_12_) & (i_13_) & (!i_14_) & (sk[5]) & (g69)) + ((g3) & (i_12_) & (i_13_) & (i_14_) & (!sk[5]) & (!g69)) + ((g3) & (i_12_) & (i_13_) & (i_14_) & (!sk[5]) & (g69)) + ((g3) & (i_12_) & (i_13_) & (i_14_) & (sk[5]) & (!g69)) + ((g3) & (i_12_) & (i_13_) & (i_14_) & (sk[5]) & (g69)));
	assign g744 = (((!g73) & (!g164) & (!g402) & (sk[6]) & (g742) & (!g743)) + ((!g73) & (!g164) & (g402) & (!sk[6]) & (!g742) & (g743)) + ((!g73) & (!g164) & (g402) & (!sk[6]) & (g742) & (!g743)) + ((!g73) & (!g164) & (g402) & (!sk[6]) & (g742) & (g743)) + ((!g73) & (!g164) & (g402) & (sk[6]) & (!g742) & (!g743)) + ((!g73) & (!g164) & (g402) & (sk[6]) & (!g742) & (g743)) + ((!g73) & (!g164) & (g402) & (sk[6]) & (g742) & (!g743)) + ((!g73) & (!g164) & (g402) & (sk[6]) & (g742) & (g743)) + ((!g73) & (g164) & (!g402) & (!sk[6]) & (!g742) & (!g743)) + ((!g73) & (g164) & (!g402) & (!sk[6]) & (!g742) & (g743)) + ((!g73) & (g164) & (!g402) & (!sk[6]) & (g742) & (!g743)) + ((!g73) & (g164) & (!g402) & (!sk[6]) & (g742) & (g743)) + ((!g73) & (g164) & (!g402) & (sk[6]) & (g742) & (!g743)) + ((!g73) & (g164) & (g402) & (!sk[6]) & (!g742) & (!g743)) + ((!g73) & (g164) & (g402) & (!sk[6]) & (!g742) & (g743)) + ((!g73) & (g164) & (g402) & (!sk[6]) & (g742) & (!g743)) + ((!g73) & (g164) & (g402) & (!sk[6]) & (g742) & (g743)) + ((!g73) & (g164) & (g402) & (sk[6]) & (g742) & (!g743)) + ((!g73) & (g164) & (g402) & (sk[6]) & (g742) & (g743)) + ((g73) & (!g164) & (!g402) & (sk[6]) & (g742) & (!g743)) + ((g73) & (!g164) & (g402) & (!sk[6]) & (!g742) & (g743)) + ((g73) & (!g164) & (g402) & (!sk[6]) & (g742) & (!g743)) + ((g73) & (!g164) & (g402) & (!sk[6]) & (g742) & (g743)) + ((g73) & (!g164) & (g402) & (sk[6]) & (g742) & (!g743)) + ((g73) & (!g164) & (g402) & (sk[6]) & (g742) & (g743)) + ((g73) & (g164) & (!g402) & (!sk[6]) & (!g742) & (!g743)) + ((g73) & (g164) & (!g402) & (!sk[6]) & (!g742) & (g743)) + ((g73) & (g164) & (!g402) & (!sk[6]) & (g742) & (!g743)) + ((g73) & (g164) & (!g402) & (!sk[6]) & (g742) & (g743)) + ((g73) & (g164) & (!g402) & (sk[6]) & (g742) & (!g743)) + ((g73) & (g164) & (g402) & (!sk[6]) & (!g742) & (!g743)) + ((g73) & (g164) & (g402) & (!sk[6]) & (!g742) & (g743)) + ((g73) & (g164) & (g402) & (!sk[6]) & (g742) & (!g743)) + ((g73) & (g164) & (g402) & (!sk[6]) & (g742) & (g743)) + ((g73) & (g164) & (g402) & (sk[6]) & (g742) & (!g743)) + ((g73) & (g164) & (g402) & (sk[6]) & (g742) & (g743)));
	assign g745 = (((!g157) & (!sk[7]) & (!g78) & (g333) & (!g723)) + ((!g157) & (!sk[7]) & (!g78) & (g333) & (g723)) + ((!g157) & (!sk[7]) & (g78) & (g333) & (!g723)) + ((!g157) & (!sk[7]) & (g78) & (g333) & (g723)) + ((g157) & (!sk[7]) & (!g78) & (g333) & (!g723)) + ((g157) & (!sk[7]) & (!g78) & (g333) & (g723)) + ((g157) & (!sk[7]) & (g78) & (g333) & (!g723)) + ((g157) & (!sk[7]) & (g78) & (g333) & (g723)) + ((g157) & (sk[7]) & (!g78) & (!g333) & (!g723)) + ((g157) & (sk[7]) & (!g78) & (!g333) & (g723)) + ((g157) & (sk[7]) & (!g78) & (g333) & (!g723)) + ((g157) & (sk[7]) & (!g78) & (g333) & (g723)) + ((g157) & (sk[7]) & (g78) & (!g333) & (g723)) + ((g157) & (sk[7]) & (g78) & (g333) & (!g723)) + ((g157) & (sk[7]) & (g78) & (g333) & (g723)));
	assign g746 = (((!g157) & (!g90) & (!g125) & (sk[8]) & (!g728) & (!g729)) + ((!g157) & (!g90) & (!g125) & (sk[8]) & (!g728) & (g729)) + ((!g157) & (!g90) & (!g125) & (sk[8]) & (g728) & (!g729)) + ((!g157) & (!g90) & (!g125) & (sk[8]) & (g728) & (g729)) + ((!g157) & (!g90) & (g125) & (!sk[8]) & (!g728) & (g729)) + ((!g157) & (!g90) & (g125) & (!sk[8]) & (g728) & (!g729)) + ((!g157) & (!g90) & (g125) & (!sk[8]) & (g728) & (g729)) + ((!g157) & (!g90) & (g125) & (sk[8]) & (!g728) & (g729)) + ((!g157) & (!g90) & (g125) & (sk[8]) & (g728) & (g729)) + ((!g157) & (g90) & (!g125) & (!sk[8]) & (!g728) & (!g729)) + ((!g157) & (g90) & (!g125) & (!sk[8]) & (!g728) & (g729)) + ((!g157) & (g90) & (!g125) & (!sk[8]) & (g728) & (!g729)) + ((!g157) & (g90) & (!g125) & (!sk[8]) & (g728) & (g729)) + ((!g157) & (g90) & (!g125) & (sk[8]) & (!g728) & (!g729)) + ((!g157) & (g90) & (!g125) & (sk[8]) & (!g728) & (g729)) + ((!g157) & (g90) & (!g125) & (sk[8]) & (g728) & (!g729)) + ((!g157) & (g90) & (!g125) & (sk[8]) & (g728) & (g729)) + ((!g157) & (g90) & (g125) & (!sk[8]) & (!g728) & (!g729)) + ((!g157) & (g90) & (g125) & (!sk[8]) & (!g728) & (g729)) + ((!g157) & (g90) & (g125) & (!sk[8]) & (g728) & (!g729)) + ((!g157) & (g90) & (g125) & (!sk[8]) & (g728) & (g729)) + ((!g157) & (g90) & (g125) & (sk[8]) & (!g728) & (g729)) + ((!g157) & (g90) & (g125) & (sk[8]) & (g728) & (g729)) + ((g157) & (!g90) & (!g125) & (sk[8]) & (!g728) & (!g729)) + ((g157) & (!g90) & (!g125) & (sk[8]) & (!g728) & (g729)) + ((g157) & (!g90) & (g125) & (!sk[8]) & (!g728) & (g729)) + ((g157) & (!g90) & (g125) & (!sk[8]) & (g728) & (!g729)) + ((g157) & (!g90) & (g125) & (!sk[8]) & (g728) & (g729)) + ((g157) & (!g90) & (g125) & (sk[8]) & (!g728) & (g729)) + ((g157) & (g90) & (!g125) & (!sk[8]) & (!g728) & (!g729)) + ((g157) & (g90) & (!g125) & (!sk[8]) & (!g728) & (g729)) + ((g157) & (g90) & (!g125) & (!sk[8]) & (g728) & (!g729)) + ((g157) & (g90) & (!g125) & (!sk[8]) & (g728) & (g729)) + ((g157) & (g90) & (g125) & (!sk[8]) & (!g728) & (!g729)) + ((g157) & (g90) & (g125) & (!sk[8]) & (!g728) & (g729)) + ((g157) & (g90) & (g125) & (!sk[8]) & (g728) & (!g729)) + ((g157) & (g90) & (g125) & (!sk[8]) & (g728) & (g729)));
	assign g747 = (((!sk[9]) & (!g165) & (!g217) & (g729) & (!g745) & (g746)) + ((!sk[9]) & (!g165) & (!g217) & (g729) & (g745) & (!g746)) + ((!sk[9]) & (!g165) & (!g217) & (g729) & (g745) & (g746)) + ((!sk[9]) & (!g165) & (g217) & (!g729) & (!g745) & (!g746)) + ((!sk[9]) & (!g165) & (g217) & (!g729) & (!g745) & (g746)) + ((!sk[9]) & (!g165) & (g217) & (!g729) & (g745) & (!g746)) + ((!sk[9]) & (!g165) & (g217) & (!g729) & (g745) & (g746)) + ((!sk[9]) & (!g165) & (g217) & (g729) & (!g745) & (!g746)) + ((!sk[9]) & (!g165) & (g217) & (g729) & (!g745) & (g746)) + ((!sk[9]) & (!g165) & (g217) & (g729) & (g745) & (!g746)) + ((!sk[9]) & (!g165) & (g217) & (g729) & (g745) & (g746)) + ((!sk[9]) & (g165) & (!g217) & (g729) & (!g745) & (g746)) + ((!sk[9]) & (g165) & (!g217) & (g729) & (g745) & (!g746)) + ((!sk[9]) & (g165) & (!g217) & (g729) & (g745) & (g746)) + ((!sk[9]) & (g165) & (g217) & (!g729) & (!g745) & (!g746)) + ((!sk[9]) & (g165) & (g217) & (!g729) & (!g745) & (g746)) + ((!sk[9]) & (g165) & (g217) & (!g729) & (g745) & (!g746)) + ((!sk[9]) & (g165) & (g217) & (!g729) & (g745) & (g746)) + ((!sk[9]) & (g165) & (g217) & (g729) & (!g745) & (!g746)) + ((!sk[9]) & (g165) & (g217) & (g729) & (!g745) & (g746)) + ((!sk[9]) & (g165) & (g217) & (g729) & (g745) & (!g746)) + ((!sk[9]) & (g165) & (g217) & (g729) & (g745) & (g746)) + ((sk[9]) & (!g165) & (!g217) & (!g729) & (!g745) & (g746)) + ((sk[9]) & (!g165) & (!g217) & (g729) & (!g745) & (g746)) + ((sk[9]) & (!g165) & (g217) & (g729) & (!g745) & (g746)) + ((sk[9]) & (g165) & (!g217) & (g729) & (!g745) & (g746)) + ((sk[9]) & (g165) & (g217) & (g729) & (!g745) & (g746)));
	assign g748 = (((g727) & (g1518) & (g734) & (g741) & (g744) & (g747)));
	assign g749 = (((!i_9_) & (!i_10_) & (i_11_) & (!sk[11]) & (!i_15_) & (g507)) + ((!i_9_) & (!i_10_) & (i_11_) & (!sk[11]) & (i_15_) & (!g507)) + ((!i_9_) & (!i_10_) & (i_11_) & (!sk[11]) & (i_15_) & (g507)) + ((!i_9_) & (!i_10_) & (i_11_) & (sk[11]) & (i_15_) & (g507)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[11]) & (!i_15_) & (!g507)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[11]) & (!i_15_) & (g507)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[11]) & (i_15_) & (!g507)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[11]) & (i_15_) & (g507)) + ((!i_9_) & (i_10_) & (!i_11_) & (sk[11]) & (i_15_) & (g507)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[11]) & (!i_15_) & (!g507)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[11]) & (!i_15_) & (g507)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[11]) & (i_15_) & (!g507)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[11]) & (i_15_) & (g507)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[11]) & (!i_15_) & (g507)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[11]) & (i_15_) & (!g507)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[11]) & (i_15_) & (g507)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[11]) & (!i_15_) & (!g507)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[11]) & (!i_15_) & (g507)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[11]) & (i_15_) & (!g507)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[11]) & (i_15_) & (g507)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[11]) & (!i_15_) & (!g507)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[11]) & (!i_15_) & (g507)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[11]) & (i_15_) & (!g507)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[11]) & (i_15_) & (g507)));
	assign g750 = (((!i_6_) & (!sk[12]) & (!g120) & (g135) & (!g113) & (g507)) + ((!i_6_) & (!sk[12]) & (!g120) & (g135) & (g113) & (!g507)) + ((!i_6_) & (!sk[12]) & (!g120) & (g135) & (g113) & (g507)) + ((!i_6_) & (!sk[12]) & (g120) & (!g135) & (!g113) & (!g507)) + ((!i_6_) & (!sk[12]) & (g120) & (!g135) & (!g113) & (g507)) + ((!i_6_) & (!sk[12]) & (g120) & (!g135) & (g113) & (!g507)) + ((!i_6_) & (!sk[12]) & (g120) & (!g135) & (g113) & (g507)) + ((!i_6_) & (!sk[12]) & (g120) & (g135) & (!g113) & (!g507)) + ((!i_6_) & (!sk[12]) & (g120) & (g135) & (!g113) & (g507)) + ((!i_6_) & (!sk[12]) & (g120) & (g135) & (g113) & (!g507)) + ((!i_6_) & (!sk[12]) & (g120) & (g135) & (g113) & (g507)) + ((!i_6_) & (sk[12]) & (!g120) & (!g135) & (!g113) & (g507)) + ((!i_6_) & (sk[12]) & (g120) & (!g135) & (!g113) & (!g507)) + ((!i_6_) & (sk[12]) & (g120) & (!g135) & (!g113) & (g507)) + ((!i_6_) & (sk[12]) & (g120) & (!g135) & (g113) & (!g507)) + ((!i_6_) & (sk[12]) & (g120) & (!g135) & (g113) & (g507)) + ((!i_6_) & (sk[12]) & (g120) & (g135) & (!g113) & (!g507)) + ((!i_6_) & (sk[12]) & (g120) & (g135) & (!g113) & (g507)) + ((!i_6_) & (sk[12]) & (g120) & (g135) & (g113) & (!g507)) + ((!i_6_) & (sk[12]) & (g120) & (g135) & (g113) & (g507)) + ((i_6_) & (!sk[12]) & (!g120) & (g135) & (!g113) & (g507)) + ((i_6_) & (!sk[12]) & (!g120) & (g135) & (g113) & (!g507)) + ((i_6_) & (!sk[12]) & (!g120) & (g135) & (g113) & (g507)) + ((i_6_) & (!sk[12]) & (g120) & (!g135) & (!g113) & (!g507)) + ((i_6_) & (!sk[12]) & (g120) & (!g135) & (!g113) & (g507)) + ((i_6_) & (!sk[12]) & (g120) & (!g135) & (g113) & (!g507)) + ((i_6_) & (!sk[12]) & (g120) & (!g135) & (g113) & (g507)) + ((i_6_) & (!sk[12]) & (g120) & (g135) & (!g113) & (!g507)) + ((i_6_) & (!sk[12]) & (g120) & (g135) & (!g113) & (g507)) + ((i_6_) & (!sk[12]) & (g120) & (g135) & (g113) & (!g507)) + ((i_6_) & (!sk[12]) & (g120) & (g135) & (g113) & (g507)) + ((i_6_) & (sk[12]) & (!g120) & (!g135) & (!g113) & (g507)) + ((i_6_) & (sk[12]) & (g120) & (!g135) & (!g113) & (g507)));
	assign g751 = (((!i_9_) & (!i_10_) & (i_11_) & (!i_15_) & (!sk[13]) & (g76)) + ((!i_9_) & (!i_10_) & (i_11_) & (i_15_) & (!sk[13]) & (!g76)) + ((!i_9_) & (!i_10_) & (i_11_) & (i_15_) & (!sk[13]) & (g76)) + ((!i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (!sk[13]) & (!g76)) + ((!i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (!sk[13]) & (g76)) + ((!i_9_) & (i_10_) & (!i_11_) & (i_15_) & (!sk[13]) & (!g76)) + ((!i_9_) & (i_10_) & (!i_11_) & (i_15_) & (!sk[13]) & (g76)) + ((!i_9_) & (i_10_) & (i_11_) & (!i_15_) & (!sk[13]) & (!g76)) + ((!i_9_) & (i_10_) & (i_11_) & (!i_15_) & (!sk[13]) & (g76)) + ((!i_9_) & (i_10_) & (i_11_) & (i_15_) & (!sk[13]) & (!g76)) + ((!i_9_) & (i_10_) & (i_11_) & (i_15_) & (!sk[13]) & (g76)) + ((i_9_) & (!i_10_) & (i_11_) & (!i_15_) & (!sk[13]) & (g76)) + ((i_9_) & (!i_10_) & (i_11_) & (i_15_) & (!sk[13]) & (!g76)) + ((i_9_) & (!i_10_) & (i_11_) & (i_15_) & (!sk[13]) & (g76)) + ((i_9_) & (!i_10_) & (i_11_) & (i_15_) & (sk[13]) & (!g76)) + ((i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (!sk[13]) & (!g76)) + ((i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (!sk[13]) & (g76)) + ((i_9_) & (i_10_) & (!i_11_) & (i_15_) & (!sk[13]) & (!g76)) + ((i_9_) & (i_10_) & (!i_11_) & (i_15_) & (!sk[13]) & (g76)) + ((i_9_) & (i_10_) & (!i_11_) & (i_15_) & (sk[13]) & (!g76)) + ((i_9_) & (i_10_) & (i_11_) & (!i_15_) & (!sk[13]) & (!g76)) + ((i_9_) & (i_10_) & (i_11_) & (!i_15_) & (!sk[13]) & (g76)) + ((i_9_) & (i_10_) & (i_11_) & (i_15_) & (!sk[13]) & (!g76)) + ((i_9_) & (i_10_) & (i_11_) & (i_15_) & (!sk[13]) & (g76)));
	assign g752 = (((!g185) & (!g416) & (!g562) & (sk[14]) & (!g751)) + ((!g185) & (!g416) & (g562) & (!sk[14]) & (!g751)) + ((!g185) & (!g416) & (g562) & (!sk[14]) & (g751)) + ((!g185) & (g416) & (g562) & (!sk[14]) & (!g751)) + ((!g185) & (g416) & (g562) & (!sk[14]) & (g751)) + ((g185) & (!g416) & (g562) & (!sk[14]) & (!g751)) + ((g185) & (!g416) & (g562) & (!sk[14]) & (g751)) + ((g185) & (g416) & (g562) & (!sk[14]) & (!g751)) + ((g185) & (g416) & (g562) & (!sk[14]) & (g751)));
	assign g753 = (((!g113) & (!sk[15]) & (!g507) & (g749) & (!g750) & (g752)) + ((!g113) & (!sk[15]) & (!g507) & (g749) & (g750) & (!g752)) + ((!g113) & (!sk[15]) & (!g507) & (g749) & (g750) & (g752)) + ((!g113) & (!sk[15]) & (g507) & (!g749) & (!g750) & (!g752)) + ((!g113) & (!sk[15]) & (g507) & (!g749) & (!g750) & (g752)) + ((!g113) & (!sk[15]) & (g507) & (!g749) & (g750) & (!g752)) + ((!g113) & (!sk[15]) & (g507) & (!g749) & (g750) & (g752)) + ((!g113) & (!sk[15]) & (g507) & (g749) & (!g750) & (!g752)) + ((!g113) & (!sk[15]) & (g507) & (g749) & (!g750) & (g752)) + ((!g113) & (!sk[15]) & (g507) & (g749) & (g750) & (!g752)) + ((!g113) & (!sk[15]) & (g507) & (g749) & (g750) & (g752)) + ((!g113) & (sk[15]) & (!g507) & (!g749) & (g750) & (!g752)) + ((!g113) & (sk[15]) & (!g507) & (g749) & (g750) & (!g752)) + ((!g113) & (sk[15]) & (!g507) & (g749) & (g750) & (g752)) + ((!g113) & (sk[15]) & (g507) & (!g749) & (g750) & (!g752)) + ((!g113) & (sk[15]) & (g507) & (!g749) & (g750) & (g752)) + ((!g113) & (sk[15]) & (g507) & (g749) & (g750) & (!g752)) + ((!g113) & (sk[15]) & (g507) & (g749) & (g750) & (g752)) + ((g113) & (!sk[15]) & (!g507) & (g749) & (!g750) & (g752)) + ((g113) & (!sk[15]) & (!g507) & (g749) & (g750) & (!g752)) + ((g113) & (!sk[15]) & (!g507) & (g749) & (g750) & (g752)) + ((g113) & (!sk[15]) & (g507) & (!g749) & (!g750) & (!g752)) + ((g113) & (!sk[15]) & (g507) & (!g749) & (!g750) & (g752)) + ((g113) & (!sk[15]) & (g507) & (!g749) & (g750) & (!g752)) + ((g113) & (!sk[15]) & (g507) & (!g749) & (g750) & (g752)) + ((g113) & (!sk[15]) & (g507) & (g749) & (!g750) & (!g752)) + ((g113) & (!sk[15]) & (g507) & (g749) & (!g750) & (g752)) + ((g113) & (!sk[15]) & (g507) & (g749) & (g750) & (!g752)) + ((g113) & (!sk[15]) & (g507) & (g749) & (g750) & (g752)) + ((g113) & (sk[15]) & (!g507) & (!g749) & (g750) & (!g752)) + ((g113) & (sk[15]) & (!g507) & (g749) & (g750) & (!g752)) + ((g113) & (sk[15]) & (!g507) & (g749) & (g750) & (g752)) + ((g113) & (sk[15]) & (g507) & (!g749) & (g750) & (!g752)) + ((g113) & (sk[15]) & (g507) & (g749) & (g750) & (!g752)) + ((g113) & (sk[15]) & (g507) & (g749) & (g750) & (g752)));
	assign g754 = (((!sk[16]) & (!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[16]) & (!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[16]) & (!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g112)) + ((!sk[16]) & (!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g112)) + ((!sk[16]) & (!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((!sk[16]) & (!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g112)) + ((!sk[16]) & (!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g112)) + ((!sk[16]) & (!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g112)) + ((!sk[16]) & (!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[16]) & (!i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[16]) & (!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g112)) + ((!sk[16]) & (i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[16]) & (i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[16]) & (i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g112)) + ((!sk[16]) & (i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g112)) + ((!sk[16]) & (i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((!sk[16]) & (i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g112)) + ((!sk[16]) & (i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g112)) + ((!sk[16]) & (i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g112)) + ((!sk[16]) & (i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[16]) & (i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[16]) & (i_15_) & (i_12_) & (i_13_) & (i_14_) & (g112)) + ((sk[16]) & (!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g112)) + ((sk[16]) & (!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g112)) + ((sk[16]) & (i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((sk[16]) & (i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((sk[16]) & (i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112)));
	assign g755 = (((!i_9_) & (!i_10_) & (i_15_) & (!sk[17]) & (!g507)) + ((!i_9_) & (!i_10_) & (i_15_) & (!sk[17]) & (g507)) + ((!i_9_) & (i_10_) & (i_15_) & (!sk[17]) & (!g507)) + ((!i_9_) & (i_10_) & (i_15_) & (!sk[17]) & (g507)) + ((!i_9_) & (i_10_) & (i_15_) & (sk[17]) & (g507)) + ((i_9_) & (!i_10_) & (i_15_) & (!sk[17]) & (!g507)) + ((i_9_) & (!i_10_) & (i_15_) & (!sk[17]) & (g507)) + ((i_9_) & (i_10_) & (i_15_) & (!sk[17]) & (!g507)) + ((i_9_) & (i_10_) & (i_15_) & (!sk[17]) & (g507)));
	assign g756 = (((!i_8_) & (!g73) & (!g130) & (!g754) & (sk[18]) & (g755)) + ((!i_8_) & (!g73) & (!g130) & (g754) & (sk[18]) & (!g755)) + ((!i_8_) & (!g73) & (!g130) & (g754) & (sk[18]) & (g755)) + ((!i_8_) & (!g73) & (g130) & (!g754) & (!sk[18]) & (g755)) + ((!i_8_) & (!g73) & (g130) & (g754) & (!sk[18]) & (!g755)) + ((!i_8_) & (!g73) & (g130) & (g754) & (!sk[18]) & (g755)) + ((!i_8_) & (g73) & (!g130) & (!g754) & (!sk[18]) & (!g755)) + ((!i_8_) & (g73) & (!g130) & (!g754) & (!sk[18]) & (g755)) + ((!i_8_) & (g73) & (!g130) & (!g754) & (sk[18]) & (g755)) + ((!i_8_) & (g73) & (!g130) & (g754) & (!sk[18]) & (!g755)) + ((!i_8_) & (g73) & (!g130) & (g754) & (!sk[18]) & (g755)) + ((!i_8_) & (g73) & (!g130) & (g754) & (sk[18]) & (!g755)) + ((!i_8_) & (g73) & (!g130) & (g754) & (sk[18]) & (g755)) + ((!i_8_) & (g73) & (g130) & (!g754) & (!sk[18]) & (!g755)) + ((!i_8_) & (g73) & (g130) & (!g754) & (!sk[18]) & (g755)) + ((!i_8_) & (g73) & (g130) & (!g754) & (sk[18]) & (g755)) + ((!i_8_) & (g73) & (g130) & (g754) & (!sk[18]) & (!g755)) + ((!i_8_) & (g73) & (g130) & (g754) & (!sk[18]) & (g755)) + ((!i_8_) & (g73) & (g130) & (g754) & (sk[18]) & (g755)) + ((i_8_) & (!g73) & (!g130) & (!g754) & (sk[18]) & (g755)) + ((i_8_) & (!g73) & (!g130) & (g754) & (sk[18]) & (!g755)) + ((i_8_) & (!g73) & (!g130) & (g754) & (sk[18]) & (g755)) + ((i_8_) & (!g73) & (g130) & (!g754) & (!sk[18]) & (g755)) + ((i_8_) & (!g73) & (g130) & (g754) & (!sk[18]) & (!g755)) + ((i_8_) & (!g73) & (g130) & (g754) & (!sk[18]) & (g755)) + ((i_8_) & (g73) & (!g130) & (!g754) & (!sk[18]) & (!g755)) + ((i_8_) & (g73) & (!g130) & (!g754) & (!sk[18]) & (g755)) + ((i_8_) & (g73) & (!g130) & (!g754) & (sk[18]) & (g755)) + ((i_8_) & (g73) & (!g130) & (g754) & (!sk[18]) & (!g755)) + ((i_8_) & (g73) & (!g130) & (g754) & (!sk[18]) & (g755)) + ((i_8_) & (g73) & (!g130) & (g754) & (sk[18]) & (!g755)) + ((i_8_) & (g73) & (!g130) & (g754) & (sk[18]) & (g755)) + ((i_8_) & (g73) & (g130) & (!g754) & (!sk[18]) & (!g755)) + ((i_8_) & (g73) & (g130) & (!g754) & (!sk[18]) & (g755)) + ((i_8_) & (g73) & (g130) & (g754) & (!sk[18]) & (!g755)) + ((i_8_) & (g73) & (g130) & (g754) & (!sk[18]) & (g755)));
	assign g757 = (((!g161) & (!g119) & (!g175) & (!g508) & (!g505) & (!g756)) + ((!g161) & (!g119) & (!g175) & (g508) & (!g505) & (!g756)) + ((!g161) & (!g119) & (g175) & (!g508) & (!g505) & (!g756)) + ((!g161) & (!g119) & (g175) & (g508) & (!g505) & (!g756)) + ((!g161) & (g119) & (!g175) & (!g508) & (!g505) & (!g756)) + ((!g161) & (g119) & (g175) & (!g508) & (!g505) & (!g756)) + ((g161) & (!g119) & (!g175) & (!g508) & (!g505) & (!g756)) + ((g161) & (!g119) & (!g175) & (g508) & (!g505) & (!g756)) + ((g161) & (g119) & (!g175) & (!g508) & (!g505) & (!g756)));
	assign g758 = (((!sk[20]) & (!g177) & (!g183) & (g278) & (!g392) & (g501)) + ((!sk[20]) & (!g177) & (!g183) & (g278) & (g392) & (!g501)) + ((!sk[20]) & (!g177) & (!g183) & (g278) & (g392) & (g501)) + ((!sk[20]) & (!g177) & (g183) & (!g278) & (!g392) & (!g501)) + ((!sk[20]) & (!g177) & (g183) & (!g278) & (!g392) & (g501)) + ((!sk[20]) & (!g177) & (g183) & (!g278) & (g392) & (!g501)) + ((!sk[20]) & (!g177) & (g183) & (!g278) & (g392) & (g501)) + ((!sk[20]) & (!g177) & (g183) & (g278) & (!g392) & (!g501)) + ((!sk[20]) & (!g177) & (g183) & (g278) & (!g392) & (g501)) + ((!sk[20]) & (!g177) & (g183) & (g278) & (g392) & (!g501)) + ((!sk[20]) & (!g177) & (g183) & (g278) & (g392) & (g501)) + ((!sk[20]) & (g177) & (!g183) & (g278) & (!g392) & (g501)) + ((!sk[20]) & (g177) & (!g183) & (g278) & (g392) & (!g501)) + ((!sk[20]) & (g177) & (!g183) & (g278) & (g392) & (g501)) + ((!sk[20]) & (g177) & (g183) & (!g278) & (!g392) & (!g501)) + ((!sk[20]) & (g177) & (g183) & (!g278) & (!g392) & (g501)) + ((!sk[20]) & (g177) & (g183) & (!g278) & (g392) & (!g501)) + ((!sk[20]) & (g177) & (g183) & (!g278) & (g392) & (g501)) + ((!sk[20]) & (g177) & (g183) & (g278) & (!g392) & (!g501)) + ((!sk[20]) & (g177) & (g183) & (g278) & (!g392) & (g501)) + ((!sk[20]) & (g177) & (g183) & (g278) & (g392) & (!g501)) + ((!sk[20]) & (g177) & (g183) & (g278) & (g392) & (g501)) + ((sk[20]) & (!g177) & (!g183) & (!g278) & (g392) & (g501)) + ((sk[20]) & (!g177) & (!g183) & (g278) & (g392) & (!g501)) + ((sk[20]) & (!g177) & (!g183) & (g278) & (g392) & (g501)) + ((sk[20]) & (!g177) & (g183) & (!g278) & (g392) & (!g501)) + ((sk[20]) & (!g177) & (g183) & (!g278) & (g392) & (g501)) + ((sk[20]) & (!g177) & (g183) & (g278) & (g392) & (!g501)) + ((sk[20]) & (!g177) & (g183) & (g278) & (g392) & (g501)) + ((sk[20]) & (g177) & (!g183) & (!g278) & (g392) & (!g501)) + ((sk[20]) & (g177) & (!g183) & (!g278) & (g392) & (g501)) + ((sk[20]) & (g177) & (!g183) & (g278) & (g392) & (!g501)) + ((sk[20]) & (g177) & (!g183) & (g278) & (g392) & (g501)) + ((sk[20]) & (g177) & (g183) & (!g278) & (g392) & (!g501)) + ((sk[20]) & (g177) & (g183) & (!g278) & (g392) & (g501)) + ((sk[20]) & (g177) & (g183) & (g278) & (g392) & (!g501)) + ((sk[20]) & (g177) & (g183) & (g278) & (g392) & (g501)));
	assign g759 = (((!g161) & (!g90) & (!g125) & (!g281) & (!g728) & (!g555)) + ((!g161) & (!g90) & (!g125) & (!g281) & (!g728) & (g555)) + ((!g161) & (!g90) & (!g125) & (!g281) & (g728) & (!g555)) + ((!g161) & (!g90) & (!g125) & (!g281) & (g728) & (g555)) + ((!g161) & (!g90) & (!g125) & (g281) & (!g728) & (!g555)) + ((!g161) & (!g90) & (!g125) & (g281) & (!g728) & (g555)) + ((!g161) & (!g90) & (!g125) & (g281) & (g728) & (!g555)) + ((!g161) & (!g90) & (!g125) & (g281) & (g728) & (g555)) + ((!g161) & (!g90) & (g125) & (!g281) & (!g728) & (!g555)) + ((!g161) & (!g90) & (g125) & (g281) & (!g728) & (!g555)) + ((!g161) & (g90) & (!g125) & (!g281) & (!g728) & (!g555)) + ((!g161) & (g90) & (!g125) & (!g281) & (!g728) & (g555)) + ((!g161) & (g90) & (!g125) & (!g281) & (g728) & (!g555)) + ((!g161) & (g90) & (!g125) & (!g281) & (g728) & (g555)) + ((!g161) & (g90) & (!g125) & (g281) & (!g728) & (!g555)) + ((!g161) & (g90) & (!g125) & (g281) & (!g728) & (g555)) + ((!g161) & (g90) & (!g125) & (g281) & (g728) & (!g555)) + ((!g161) & (g90) & (!g125) & (g281) & (g728) & (g555)) + ((!g161) & (g90) & (g125) & (!g281) & (!g728) & (!g555)) + ((!g161) & (g90) & (g125) & (g281) & (!g728) & (!g555)) + ((g161) & (!g90) & (!g125) & (!g281) & (!g728) & (!g555)) + ((g161) & (!g90) & (!g125) & (!g281) & (!g728) & (g555)) + ((g161) & (!g90) & (g125) & (!g281) & (!g728) & (!g555)));
	assign g760 = (((!g159) & (!g336) & (g627) & (!sk[22]) & (!g758) & (g759)) + ((!g159) & (!g336) & (g627) & (!sk[22]) & (g758) & (!g759)) + ((!g159) & (!g336) & (g627) & (!sk[22]) & (g758) & (g759)) + ((!g159) & (g336) & (!g627) & (!sk[22]) & (!g758) & (!g759)) + ((!g159) & (g336) & (!g627) & (!sk[22]) & (!g758) & (g759)) + ((!g159) & (g336) & (!g627) & (!sk[22]) & (g758) & (!g759)) + ((!g159) & (g336) & (!g627) & (!sk[22]) & (g758) & (g759)) + ((!g159) & (g336) & (!g627) & (sk[22]) & (!g758) & (g759)) + ((!g159) & (g336) & (g627) & (!sk[22]) & (!g758) & (!g759)) + ((!g159) & (g336) & (g627) & (!sk[22]) & (!g758) & (g759)) + ((!g159) & (g336) & (g627) & (!sk[22]) & (g758) & (!g759)) + ((!g159) & (g336) & (g627) & (!sk[22]) & (g758) & (g759)) + ((g159) & (!g336) & (!g627) & (sk[22]) & (!g758) & (g759)) + ((g159) & (!g336) & (g627) & (!sk[22]) & (!g758) & (g759)) + ((g159) & (!g336) & (g627) & (!sk[22]) & (g758) & (!g759)) + ((g159) & (!g336) & (g627) & (!sk[22]) & (g758) & (g759)) + ((g159) & (!g336) & (g627) & (sk[22]) & (!g758) & (g759)) + ((g159) & (g336) & (!g627) & (!sk[22]) & (!g758) & (!g759)) + ((g159) & (g336) & (!g627) & (!sk[22]) & (!g758) & (g759)) + ((g159) & (g336) & (!g627) & (!sk[22]) & (g758) & (!g759)) + ((g159) & (g336) & (!g627) & (!sk[22]) & (g758) & (g759)) + ((g159) & (g336) & (!g627) & (sk[22]) & (!g758) & (g759)) + ((g159) & (g336) & (g627) & (!sk[22]) & (!g758) & (!g759)) + ((g159) & (g336) & (g627) & (!sk[22]) & (!g758) & (g759)) + ((g159) & (g336) & (g627) & (!sk[22]) & (g758) & (!g759)) + ((g159) & (g336) & (g627) & (!sk[22]) & (g758) & (g759)) + ((g159) & (g336) & (g627) & (sk[22]) & (!g758) & (g759)));
	assign g761 = (((!sk[23]) & (g343) & (!g626)) + ((!sk[23]) & (g343) & (g626)) + ((sk[23]) & (g343) & (!g626)));
	assign g762 = (((!g27) & (!g168) & (!sk[24]) & (g735) & (!g719)) + ((!g27) & (!g168) & (!sk[24]) & (g735) & (g719)) + ((!g27) & (g168) & (!sk[24]) & (g735) & (!g719)) + ((!g27) & (g168) & (!sk[24]) & (g735) & (g719)) + ((!g27) & (g168) & (sk[24]) & (!g735) & (!g719)) + ((!g27) & (g168) & (sk[24]) & (g735) & (!g719)) + ((g27) & (!g168) & (!sk[24]) & (g735) & (!g719)) + ((g27) & (!g168) & (!sk[24]) & (g735) & (g719)) + ((g27) & (g168) & (!sk[24]) & (g735) & (!g719)) + ((g27) & (g168) & (!sk[24]) & (g735) & (g719)) + ((g27) & (g168) & (sk[24]) & (!g735) & (!g719)) + ((g27) & (g168) & (sk[24]) & (g735) & (!g719)) + ((g27) & (g168) & (sk[24]) & (g735) & (g719)));
	assign g763 = (((!g125) & (!g413) & (!g439) & (g761) & (sk[25]) & (!g762)) + ((!g125) & (!g413) & (g439) & (!g761) & (!sk[25]) & (g762)) + ((!g125) & (!g413) & (g439) & (g761) & (!sk[25]) & (!g762)) + ((!g125) & (!g413) & (g439) & (g761) & (!sk[25]) & (g762)) + ((!g125) & (!g413) & (g439) & (g761) & (sk[25]) & (!g762)) + ((!g125) & (g413) & (!g439) & (!g761) & (!sk[25]) & (!g762)) + ((!g125) & (g413) & (!g439) & (!g761) & (!sk[25]) & (g762)) + ((!g125) & (g413) & (!g439) & (g761) & (!sk[25]) & (!g762)) + ((!g125) & (g413) & (!g439) & (g761) & (!sk[25]) & (g762)) + ((!g125) & (g413) & (!g439) & (g761) & (sk[25]) & (!g762)) + ((!g125) & (g413) & (g439) & (!g761) & (!sk[25]) & (!g762)) + ((!g125) & (g413) & (g439) & (!g761) & (!sk[25]) & (g762)) + ((!g125) & (g413) & (g439) & (!g761) & (sk[25]) & (!g762)) + ((!g125) & (g413) & (g439) & (g761) & (!sk[25]) & (!g762)) + ((!g125) & (g413) & (g439) & (g761) & (!sk[25]) & (g762)) + ((!g125) & (g413) & (g439) & (g761) & (sk[25]) & (!g762)) + ((g125) & (!g413) & (!g439) & (g761) & (sk[25]) & (!g762)) + ((g125) & (!g413) & (g439) & (!g761) & (!sk[25]) & (g762)) + ((g125) & (!g413) & (g439) & (g761) & (!sk[25]) & (!g762)) + ((g125) & (!g413) & (g439) & (g761) & (!sk[25]) & (g762)) + ((g125) & (!g413) & (g439) & (g761) & (sk[25]) & (!g762)) + ((g125) & (g413) & (!g439) & (!g761) & (!sk[25]) & (!g762)) + ((g125) & (g413) & (!g439) & (!g761) & (!sk[25]) & (g762)) + ((g125) & (g413) & (!g439) & (g761) & (!sk[25]) & (!g762)) + ((g125) & (g413) & (!g439) & (g761) & (!sk[25]) & (g762)) + ((g125) & (g413) & (!g439) & (g761) & (sk[25]) & (!g762)) + ((g125) & (g413) & (g439) & (!g761) & (!sk[25]) & (!g762)) + ((g125) & (g413) & (g439) & (!g761) & (!sk[25]) & (g762)) + ((g125) & (g413) & (g439) & (g761) & (!sk[25]) & (!g762)) + ((g125) & (g413) & (g439) & (g761) & (!sk[25]) & (g762)) + ((g125) & (g413) & (g439) & (g761) & (sk[25]) & (!g762)));
	assign g764 = (((!g753) & (!g582) & (g587) & (g757) & (g760) & (g763)));
	assign g765 = (((!g75) & (sk[27]) & (g197)) + ((g75) & (!sk[27]) & (!g197)) + ((g75) & (!sk[27]) & (g197)));
	assign g766 = (((!g164) & (!sk[28]) & (!g102) & (g397)) + ((!g164) & (!sk[28]) & (g102) & (!g397)) + ((!g164) & (!sk[28]) & (g102) & (g397)) + ((!g164) & (sk[28]) & (g102) & (g397)) + ((g164) & (!sk[28]) & (!g102) & (g397)) + ((g164) & (!sk[28]) & (g102) & (!g397)) + ((g164) & (!sk[28]) & (g102) & (g397)) + ((g164) & (sk[28]) & (!g102) & (g397)) + ((g164) & (sk[28]) & (g102) & (g397)));
	assign g767 = (((!i_7_) & (!g17) & (g72) & (!sk[29]) & (!g76)) + ((!i_7_) & (!g17) & (g72) & (!sk[29]) & (g76)) + ((!i_7_) & (g17) & (g72) & (!sk[29]) & (!g76)) + ((!i_7_) & (g17) & (g72) & (!sk[29]) & (g76)) + ((i_7_) & (!g17) & (g72) & (!sk[29]) & (!g76)) + ((i_7_) & (!g17) & (g72) & (!sk[29]) & (g76)) + ((i_7_) & (g17) & (g72) & (!sk[29]) & (!g76)) + ((i_7_) & (g17) & (g72) & (!sk[29]) & (g76)) + ((i_7_) & (g17) & (g72) & (sk[29]) & (!g76)));
	assign g768 = (((!g102) & (!g257) & (!g313) & (!g217) & (!g737) & (!g684)) + ((!g102) & (!g257) & (!g313) & (!g217) & (!g737) & (g684)) + ((!g102) & (!g257) & (!g313) & (!g217) & (g737) & (!g684)) + ((!g102) & (!g257) & (!g313) & (!g217) & (g737) & (g684)) + ((!g102) & (!g257) & (!g313) & (g217) & (g737) & (g684)) + ((!g102) & (!g257) & (g313) & (!g217) & (g737) & (!g684)) + ((!g102) & (!g257) & (g313) & (!g217) & (g737) & (g684)) + ((!g102) & (!g257) & (g313) & (g217) & (g737) & (g684)) + ((!g102) & (g257) & (!g313) & (!g217) & (g737) & (!g684)) + ((!g102) & (g257) & (!g313) & (!g217) & (g737) & (g684)) + ((!g102) & (g257) & (!g313) & (g217) & (g737) & (g684)) + ((!g102) & (g257) & (g313) & (!g217) & (g737) & (!g684)) + ((!g102) & (g257) & (g313) & (!g217) & (g737) & (g684)) + ((!g102) & (g257) & (g313) & (g217) & (g737) & (g684)) + ((g102) & (!g257) & (!g313) & (!g217) & (g737) & (!g684)) + ((g102) & (!g257) & (!g313) & (!g217) & (g737) & (g684)) + ((g102) & (!g257) & (!g313) & (g217) & (g737) & (g684)) + ((g102) & (!g257) & (g313) & (!g217) & (g737) & (!g684)) + ((g102) & (!g257) & (g313) & (!g217) & (g737) & (g684)) + ((g102) & (!g257) & (g313) & (g217) & (g737) & (g684)) + ((g102) & (g257) & (!g313) & (!g217) & (g737) & (!g684)) + ((g102) & (g257) & (!g313) & (!g217) & (g737) & (g684)) + ((g102) & (g257) & (!g313) & (g217) & (g737) & (g684)) + ((g102) & (g257) & (g313) & (!g217) & (g737) & (!g684)) + ((g102) & (g257) & (g313) & (!g217) & (g737) & (g684)) + ((g102) & (g257) & (g313) & (g217) & (g737) & (g684)));
	assign g769 = (((!g142) & (!g749) & (!g766) & (sk[31]) & (!g767) & (g768)) + ((!g142) & (!g749) & (g766) & (!sk[31]) & (!g767) & (g768)) + ((!g142) & (!g749) & (g766) & (!sk[31]) & (g767) & (!g768)) + ((!g142) & (!g749) & (g766) & (!sk[31]) & (g767) & (g768)) + ((!g142) & (g749) & (!g766) & (!sk[31]) & (!g767) & (!g768)) + ((!g142) & (g749) & (!g766) & (!sk[31]) & (!g767) & (g768)) + ((!g142) & (g749) & (!g766) & (!sk[31]) & (g767) & (!g768)) + ((!g142) & (g749) & (!g766) & (!sk[31]) & (g767) & (g768)) + ((!g142) & (g749) & (g766) & (!sk[31]) & (!g767) & (!g768)) + ((!g142) & (g749) & (g766) & (!sk[31]) & (!g767) & (g768)) + ((!g142) & (g749) & (g766) & (!sk[31]) & (g767) & (!g768)) + ((!g142) & (g749) & (g766) & (!sk[31]) & (g767) & (g768)) + ((g142) & (!g749) & (!g766) & (sk[31]) & (!g767) & (g768)) + ((g142) & (!g749) & (g766) & (!sk[31]) & (!g767) & (g768)) + ((g142) & (!g749) & (g766) & (!sk[31]) & (g767) & (!g768)) + ((g142) & (!g749) & (g766) & (!sk[31]) & (g767) & (g768)) + ((g142) & (g749) & (!g766) & (!sk[31]) & (!g767) & (!g768)) + ((g142) & (g749) & (!g766) & (!sk[31]) & (!g767) & (g768)) + ((g142) & (g749) & (!g766) & (!sk[31]) & (g767) & (!g768)) + ((g142) & (g749) & (!g766) & (!sk[31]) & (g767) & (g768)) + ((g142) & (g749) & (!g766) & (sk[31]) & (!g767) & (g768)) + ((g142) & (g749) & (g766) & (!sk[31]) & (!g767) & (!g768)) + ((g142) & (g749) & (g766) & (!sk[31]) & (!g767) & (g768)) + ((g142) & (g749) & (g766) & (!sk[31]) & (g767) & (!g768)) + ((g142) & (g749) & (g766) & (!sk[31]) & (g767) & (g768)));
	assign g770 = (((!sk[32]) & (!i_15_) & (!g19) & (g445) & (!g176)) + ((!sk[32]) & (!i_15_) & (!g19) & (g445) & (g176)) + ((!sk[32]) & (!i_15_) & (g19) & (g445) & (!g176)) + ((!sk[32]) & (!i_15_) & (g19) & (g445) & (g176)) + ((!sk[32]) & (i_15_) & (!g19) & (g445) & (!g176)) + ((!sk[32]) & (i_15_) & (!g19) & (g445) & (g176)) + ((!sk[32]) & (i_15_) & (g19) & (g445) & (!g176)) + ((!sk[32]) & (i_15_) & (g19) & (g445) & (g176)) + ((sk[32]) & (!i_15_) & (!g19) & (g445) & (!g176)) + ((sk[32]) & (!i_15_) & (g19) & (g445) & (!g176)) + ((sk[32]) & (i_15_) & (g19) & (g445) & (!g176)) + ((sk[32]) & (i_15_) & (g19) & (g445) & (g176)));
	assign g771 = (((!i_8_) & (!sk[33]) & (!g73) & (g508) & (!g719)) + ((!i_8_) & (!sk[33]) & (!g73) & (g508) & (g719)) + ((!i_8_) & (!sk[33]) & (g73) & (g508) & (!g719)) + ((!i_8_) & (!sk[33]) & (g73) & (g508) & (g719)) + ((!i_8_) & (sk[33]) & (g73) & (!g508) & (!g719)) + ((!i_8_) & (sk[33]) & (g73) & (g508) & (!g719)) + ((!i_8_) & (sk[33]) & (g73) & (g508) & (g719)) + ((i_8_) & (!sk[33]) & (!g73) & (g508) & (!g719)) + ((i_8_) & (!sk[33]) & (!g73) & (g508) & (g719)) + ((i_8_) & (!sk[33]) & (g73) & (g508) & (!g719)) + ((i_8_) & (!sk[33]) & (g73) & (g508) & (g719)));
	assign g772 = (((!g105) & (!g438) & (!sk[34]) & (g439) & (!g770) & (g771)) + ((!g105) & (!g438) & (!sk[34]) & (g439) & (g770) & (!g771)) + ((!g105) & (!g438) & (!sk[34]) & (g439) & (g770) & (g771)) + ((!g105) & (!g438) & (sk[34]) & (!g439) & (!g770) & (!g771)) + ((!g105) & (!g438) & (sk[34]) & (g439) & (!g770) & (!g771)) + ((!g105) & (g438) & (!sk[34]) & (!g439) & (!g770) & (!g771)) + ((!g105) & (g438) & (!sk[34]) & (!g439) & (!g770) & (g771)) + ((!g105) & (g438) & (!sk[34]) & (!g439) & (g770) & (!g771)) + ((!g105) & (g438) & (!sk[34]) & (!g439) & (g770) & (g771)) + ((!g105) & (g438) & (!sk[34]) & (g439) & (!g770) & (!g771)) + ((!g105) & (g438) & (!sk[34]) & (g439) & (!g770) & (g771)) + ((!g105) & (g438) & (!sk[34]) & (g439) & (g770) & (!g771)) + ((!g105) & (g438) & (!sk[34]) & (g439) & (g770) & (g771)) + ((!g105) & (g438) & (sk[34]) & (!g439) & (!g770) & (!g771)) + ((!g105) & (g438) & (sk[34]) & (g439) & (!g770) & (!g771)) + ((g105) & (!g438) & (!sk[34]) & (g439) & (!g770) & (g771)) + ((g105) & (!g438) & (!sk[34]) & (g439) & (g770) & (!g771)) + ((g105) & (!g438) & (!sk[34]) & (g439) & (g770) & (g771)) + ((g105) & (!g438) & (sk[34]) & (!g439) & (!g770) & (!g771)) + ((g105) & (!g438) & (sk[34]) & (g439) & (!g770) & (!g771)) + ((g105) & (g438) & (!sk[34]) & (!g439) & (!g770) & (!g771)) + ((g105) & (g438) & (!sk[34]) & (!g439) & (!g770) & (g771)) + ((g105) & (g438) & (!sk[34]) & (!g439) & (g770) & (!g771)) + ((g105) & (g438) & (!sk[34]) & (!g439) & (g770) & (g771)) + ((g105) & (g438) & (!sk[34]) & (g439) & (!g770) & (!g771)) + ((g105) & (g438) & (!sk[34]) & (g439) & (!g770) & (g771)) + ((g105) & (g438) & (!sk[34]) & (g439) & (g770) & (!g771)) + ((g105) & (g438) & (!sk[34]) & (g439) & (g770) & (g771)) + ((g105) & (g438) & (sk[34]) & (!g439) & (!g770) & (!g771)) + ((g105) & (g438) & (sk[34]) & (g439) & (!g770) & (!g771)) + ((g105) & (g438) & (sk[34]) & (g439) & (g770) & (!g771)));
	assign g773 = (((!g765) & (!g271) & (g284) & (g202) & (g769) & (g772)));
	assign g774 = (((!i_8_) & (g165) & (!g83) & (!g182) & (!g735) & (g723)) + ((!i_8_) & (g165) & (!g83) & (!g182) & (g735) & (g723)) + ((!i_8_) & (g165) & (!g83) & (g182) & (!g735) & (g723)) + ((!i_8_) & (g165) & (!g83) & (g182) & (g735) & (g723)) + ((!i_8_) & (g165) & (g83) & (!g182) & (!g735) & (g723)) + ((!i_8_) & (g165) & (g83) & (!g182) & (g735) & (!g723)) + ((!i_8_) & (g165) & (g83) & (!g182) & (g735) & (g723)) + ((!i_8_) & (g165) & (g83) & (g182) & (!g735) & (g723)) + ((!i_8_) & (g165) & (g83) & (g182) & (g735) & (!g723)) + ((!i_8_) & (g165) & (g83) & (g182) & (g735) & (g723)) + ((i_8_) & (g165) & (!g83) & (g182) & (!g735) & (!g723)) + ((i_8_) & (g165) & (!g83) & (g182) & (!g735) & (g723)) + ((i_8_) & (g165) & (!g83) & (g182) & (g735) & (!g723)) + ((i_8_) & (g165) & (!g83) & (g182) & (g735) & (g723)) + ((i_8_) & (g165) & (g83) & (g182) & (!g735) & (!g723)) + ((i_8_) & (g165) & (g83) & (g182) & (!g735) & (g723)) + ((i_8_) & (g165) & (g83) & (g182) & (g735) & (!g723)) + ((i_8_) & (g165) & (g83) & (g182) & (g735) & (g723)));
	assign g775 = (((!sk[37]) & (!g87) & (!g135) & (g272) & (!g534)) + ((!sk[37]) & (!g87) & (!g135) & (g272) & (g534)) + ((!sk[37]) & (!g87) & (g135) & (g272) & (!g534)) + ((!sk[37]) & (!g87) & (g135) & (g272) & (g534)) + ((!sk[37]) & (g87) & (!g135) & (g272) & (!g534)) + ((!sk[37]) & (g87) & (!g135) & (g272) & (g534)) + ((!sk[37]) & (g87) & (g135) & (g272) & (!g534)) + ((!sk[37]) & (g87) & (g135) & (g272) & (g534)) + ((sk[37]) & (!g87) & (!g135) & (!g272) & (!g534)) + ((sk[37]) & (!g87) & (!g135) & (!g272) & (g534)) + ((sk[37]) & (!g87) & (!g135) & (g272) & (!g534)) + ((sk[37]) & (!g87) & (!g135) & (g272) & (g534)) + ((sk[37]) & (g87) & (!g135) & (!g272) & (g534)) + ((sk[37]) & (g87) & (!g135) & (g272) & (!g534)) + ((sk[37]) & (g87) & (!g135) & (g272) & (g534)));
	assign g776 = (((!g20) & (!g355) & (!sk[38]) & (g122) & (!g495)) + ((!g20) & (!g355) & (!sk[38]) & (g122) & (g495)) + ((!g20) & (!g355) & (sk[38]) & (g122) & (g495)) + ((!g20) & (g355) & (!sk[38]) & (g122) & (!g495)) + ((!g20) & (g355) & (!sk[38]) & (g122) & (g495)) + ((!g20) & (g355) & (sk[38]) & (g122) & (g495)) + ((g20) & (!g355) & (!sk[38]) & (g122) & (!g495)) + ((g20) & (!g355) & (!sk[38]) & (g122) & (g495)) + ((g20) & (!g355) & (sk[38]) & (g122) & (g495)) + ((g20) & (g355) & (!sk[38]) & (g122) & (!g495)) + ((g20) & (g355) & (!sk[38]) & (g122) & (g495)) + ((g20) & (g355) & (sk[38]) & (g122) & (!g495)) + ((g20) & (g355) & (sk[38]) & (g122) & (g495)));
	assign g777 = (((!i_8_) & (!i_12_) & (!i_13_) & (!i_14_) & (!g22) & (!g35)) + ((!i_8_) & (!i_12_) & (!i_13_) & (!i_14_) & (!g22) & (g35)) + ((!i_8_) & (!i_12_) & (i_13_) & (i_14_) & (!g22) & (!g35)) + ((!i_8_) & (!i_12_) & (i_13_) & (i_14_) & (!g22) & (g35)) + ((!i_8_) & (i_12_) & (!i_13_) & (!i_14_) & (!g22) & (!g35)) + ((!i_8_) & (i_12_) & (!i_13_) & (!i_14_) & (!g22) & (g35)) + ((!i_8_) & (i_12_) & (!i_13_) & (i_14_) & (!g22) & (!g35)) + ((!i_8_) & (i_12_) & (!i_13_) & (i_14_) & (!g22) & (g35)) + ((!i_8_) & (i_12_) & (i_13_) & (!i_14_) & (!g22) & (!g35)) + ((!i_8_) & (i_12_) & (i_13_) & (!i_14_) & (!g22) & (g35)) + ((i_8_) & (!i_12_) & (i_13_) & (!i_14_) & (!g22) & (g35)) + ((i_8_) & (!i_12_) & (i_13_) & (!i_14_) & (g22) & (g35)) + ((i_8_) & (i_12_) & (!i_13_) & (!i_14_) & (!g22) & (g35)) + ((i_8_) & (i_12_) & (!i_13_) & (!i_14_) & (g22) & (g35)));
	assign g778 = (((!g165) & (!sk[40]) & (!g339) & (g777)) + ((!g165) & (!sk[40]) & (g339) & (!g777)) + ((!g165) & (!sk[40]) & (g339) & (g777)) + ((g165) & (!sk[40]) & (!g339) & (g777)) + ((g165) & (!sk[40]) & (g339) & (!g777)) + ((g165) & (!sk[40]) & (g339) & (g777)) + ((g165) & (sk[40]) & (!g339) & (g777)) + ((g165) & (sk[40]) & (g339) & (!g777)) + ((g165) & (sk[40]) & (g339) & (g777)));
	assign g779 = (((!g122) & (!g194) & (!sk[41]) & (g775) & (!g776) & (g778)) + ((!g122) & (!g194) & (!sk[41]) & (g775) & (g776) & (!g778)) + ((!g122) & (!g194) & (!sk[41]) & (g775) & (g776) & (g778)) + ((!g122) & (!g194) & (sk[41]) & (!g775) & (!g776) & (!g778)) + ((!g122) & (g194) & (!sk[41]) & (!g775) & (!g776) & (!g778)) + ((!g122) & (g194) & (!sk[41]) & (!g775) & (!g776) & (g778)) + ((!g122) & (g194) & (!sk[41]) & (!g775) & (g776) & (!g778)) + ((!g122) & (g194) & (!sk[41]) & (!g775) & (g776) & (g778)) + ((!g122) & (g194) & (!sk[41]) & (g775) & (!g776) & (!g778)) + ((!g122) & (g194) & (!sk[41]) & (g775) & (!g776) & (g778)) + ((!g122) & (g194) & (!sk[41]) & (g775) & (g776) & (!g778)) + ((!g122) & (g194) & (!sk[41]) & (g775) & (g776) & (g778)) + ((!g122) & (g194) & (sk[41]) & (!g775) & (!g776) & (!g778)) + ((g122) & (!g194) & (!sk[41]) & (g775) & (!g776) & (g778)) + ((g122) & (!g194) & (!sk[41]) & (g775) & (g776) & (!g778)) + ((g122) & (!g194) & (!sk[41]) & (g775) & (g776) & (g778)) + ((g122) & (!g194) & (sk[41]) & (!g775) & (!g776) & (!g778)) + ((g122) & (g194) & (!sk[41]) & (!g775) & (!g776) & (!g778)) + ((g122) & (g194) & (!sk[41]) & (!g775) & (!g776) & (g778)) + ((g122) & (g194) & (!sk[41]) & (!g775) & (g776) & (!g778)) + ((g122) & (g194) & (!sk[41]) & (!g775) & (g776) & (g778)) + ((g122) & (g194) & (!sk[41]) & (g775) & (!g776) & (!g778)) + ((g122) & (g194) & (!sk[41]) & (g775) & (!g776) & (g778)) + ((g122) & (g194) & (!sk[41]) & (g775) & (g776) & (!g778)) + ((g122) & (g194) & (!sk[41]) & (g775) & (g776) & (g778)));
	assign g780 = (((!sk[42]) & (!g85) & (!g96) & (g99) & (!g774) & (g779)) + ((!sk[42]) & (!g85) & (!g96) & (g99) & (g774) & (!g779)) + ((!sk[42]) & (!g85) & (!g96) & (g99) & (g774) & (g779)) + ((!sk[42]) & (!g85) & (g96) & (!g99) & (!g774) & (!g779)) + ((!sk[42]) & (!g85) & (g96) & (!g99) & (!g774) & (g779)) + ((!sk[42]) & (!g85) & (g96) & (!g99) & (g774) & (!g779)) + ((!sk[42]) & (!g85) & (g96) & (!g99) & (g774) & (g779)) + ((!sk[42]) & (!g85) & (g96) & (g99) & (!g774) & (!g779)) + ((!sk[42]) & (!g85) & (g96) & (g99) & (!g774) & (g779)) + ((!sk[42]) & (!g85) & (g96) & (g99) & (g774) & (!g779)) + ((!sk[42]) & (!g85) & (g96) & (g99) & (g774) & (g779)) + ((!sk[42]) & (g85) & (!g96) & (g99) & (!g774) & (g779)) + ((!sk[42]) & (g85) & (!g96) & (g99) & (g774) & (!g779)) + ((!sk[42]) & (g85) & (!g96) & (g99) & (g774) & (g779)) + ((!sk[42]) & (g85) & (g96) & (!g99) & (!g774) & (!g779)) + ((!sk[42]) & (g85) & (g96) & (!g99) & (!g774) & (g779)) + ((!sk[42]) & (g85) & (g96) & (!g99) & (g774) & (!g779)) + ((!sk[42]) & (g85) & (g96) & (!g99) & (g774) & (g779)) + ((!sk[42]) & (g85) & (g96) & (g99) & (!g774) & (!g779)) + ((!sk[42]) & (g85) & (g96) & (g99) & (!g774) & (g779)) + ((!sk[42]) & (g85) & (g96) & (g99) & (g774) & (!g779)) + ((!sk[42]) & (g85) & (g96) & (g99) & (g774) & (g779)) + ((sk[42]) & (g85) & (g96) & (!g99) & (!g774) & (g779)));
	assign g781 = (((g722) & (g322) & (g748) & (g764) & (g773) & (g780)));
	assign g782 = (((g346) & (!g354) & (g361) & (g387) & (g411) & (g581)));
	assign g783 = (((!g21) & (!sk[45]) & (!g23) & (g122)) + ((!g21) & (!sk[45]) & (g23) & (!g122)) + ((!g21) & (!sk[45]) & (g23) & (g122)) + ((!g21) & (sk[45]) & (!g23) & (g122)) + ((g21) & (!sk[45]) & (!g23) & (g122)) + ((g21) & (!sk[45]) & (g23) & (!g122)) + ((g21) & (!sk[45]) & (g23) & (g122)) + ((g21) & (sk[45]) & (!g23) & (g122)) + ((g21) & (sk[45]) & (g23) & (g122)));
	assign g784 = (((!g122) & (!g699) & (!sk[46]) & (g700)) + ((!g122) & (g699) & (!sk[46]) & (!g700)) + ((!g122) & (g699) & (!sk[46]) & (g700)) + ((g122) & (!g699) & (!sk[46]) & (g700)) + ((g122) & (!g699) & (sk[46]) & (!g700)) + ((g122) & (!g699) & (sk[46]) & (g700)) + ((g122) & (g699) & (!sk[46]) & (!g700)) + ((g122) & (g699) & (!sk[46]) & (g700)) + ((g122) & (g699) & (sk[46]) & (!g700)));
	assign g785 = (((!g634) & (!g135) & (!g651) & (!g648) & (sk[47]) & (!g703)) + ((!g634) & (!g135) & (!g651) & (!g648) & (sk[47]) & (g703)) + ((!g634) & (!g135) & (!g651) & (g648) & (sk[47]) & (!g703)) + ((!g634) & (!g135) & (!g651) & (g648) & (sk[47]) & (g703)) + ((!g634) & (!g135) & (g651) & (!g648) & (!sk[47]) & (g703)) + ((!g634) & (!g135) & (g651) & (!g648) & (sk[47]) & (!g703)) + ((!g634) & (!g135) & (g651) & (!g648) & (sk[47]) & (g703)) + ((!g634) & (!g135) & (g651) & (g648) & (!sk[47]) & (!g703)) + ((!g634) & (!g135) & (g651) & (g648) & (!sk[47]) & (g703)) + ((!g634) & (!g135) & (g651) & (g648) & (sk[47]) & (!g703)) + ((!g634) & (!g135) & (g651) & (g648) & (sk[47]) & (g703)) + ((!g634) & (g135) & (!g651) & (!g648) & (!sk[47]) & (!g703)) + ((!g634) & (g135) & (!g651) & (!g648) & (!sk[47]) & (g703)) + ((!g634) & (g135) & (!g651) & (g648) & (!sk[47]) & (!g703)) + ((!g634) & (g135) & (!g651) & (g648) & (!sk[47]) & (g703)) + ((!g634) & (g135) & (g651) & (!g648) & (!sk[47]) & (!g703)) + ((!g634) & (g135) & (g651) & (!g648) & (!sk[47]) & (g703)) + ((!g634) & (g135) & (g651) & (g648) & (!sk[47]) & (!g703)) + ((!g634) & (g135) & (g651) & (g648) & (!sk[47]) & (g703)) + ((g634) & (!g135) & (!g651) & (!g648) & (sk[47]) & (!g703)) + ((g634) & (!g135) & (!g651) & (g648) & (sk[47]) & (!g703)) + ((g634) & (!g135) & (!g651) & (g648) & (sk[47]) & (g703)) + ((g634) & (!g135) & (g651) & (!g648) & (!sk[47]) & (g703)) + ((g634) & (!g135) & (g651) & (!g648) & (sk[47]) & (!g703)) + ((g634) & (!g135) & (g651) & (!g648) & (sk[47]) & (g703)) + ((g634) & (!g135) & (g651) & (g648) & (!sk[47]) & (!g703)) + ((g634) & (!g135) & (g651) & (g648) & (!sk[47]) & (g703)) + ((g634) & (!g135) & (g651) & (g648) & (sk[47]) & (!g703)) + ((g634) & (!g135) & (g651) & (g648) & (sk[47]) & (g703)) + ((g634) & (g135) & (!g651) & (!g648) & (!sk[47]) & (!g703)) + ((g634) & (g135) & (!g651) & (!g648) & (!sk[47]) & (g703)) + ((g634) & (g135) & (!g651) & (g648) & (!sk[47]) & (!g703)) + ((g634) & (g135) & (!g651) & (g648) & (!sk[47]) & (g703)) + ((g634) & (g135) & (g651) & (!g648) & (!sk[47]) & (!g703)) + ((g634) & (g135) & (g651) & (!g648) & (!sk[47]) & (g703)) + ((g634) & (g135) & (g651) & (g648) & (!sk[47]) & (!g703)) + ((g634) & (g135) & (g651) & (g648) & (!sk[47]) & (g703)));
	assign g786 = (((!g18) & (!g33) & (!sk[48]) & (g135) & (!g122) & (g785)) + ((!g18) & (!g33) & (!sk[48]) & (g135) & (g122) & (!g785)) + ((!g18) & (!g33) & (!sk[48]) & (g135) & (g122) & (g785)) + ((!g18) & (!g33) & (sk[48]) & (!g135) & (!g122) & (!g785)) + ((!g18) & (!g33) & (sk[48]) & (!g135) & (g122) & (!g785)) + ((!g18) & (!g33) & (sk[48]) & (g135) & (!g122) & (!g785)) + ((!g18) & (!g33) & (sk[48]) & (g135) & (g122) & (!g785)) + ((!g18) & (g33) & (!sk[48]) & (!g135) & (!g122) & (!g785)) + ((!g18) & (g33) & (!sk[48]) & (!g135) & (!g122) & (g785)) + ((!g18) & (g33) & (!sk[48]) & (!g135) & (g122) & (!g785)) + ((!g18) & (g33) & (!sk[48]) & (!g135) & (g122) & (g785)) + ((!g18) & (g33) & (!sk[48]) & (g135) & (!g122) & (!g785)) + ((!g18) & (g33) & (!sk[48]) & (g135) & (!g122) & (g785)) + ((!g18) & (g33) & (!sk[48]) & (g135) & (g122) & (!g785)) + ((!g18) & (g33) & (!sk[48]) & (g135) & (g122) & (g785)) + ((!g18) & (g33) & (sk[48]) & (g135) & (!g122) & (!g785)) + ((g18) & (!g33) & (!sk[48]) & (g135) & (!g122) & (g785)) + ((g18) & (!g33) & (!sk[48]) & (g135) & (g122) & (!g785)) + ((g18) & (!g33) & (!sk[48]) & (g135) & (g122) & (g785)) + ((g18) & (!g33) & (sk[48]) & (g135) & (!g122) & (!g785)) + ((g18) & (g33) & (!sk[48]) & (!g135) & (!g122) & (!g785)) + ((g18) & (g33) & (!sk[48]) & (!g135) & (!g122) & (g785)) + ((g18) & (g33) & (!sk[48]) & (!g135) & (g122) & (!g785)) + ((g18) & (g33) & (!sk[48]) & (!g135) & (g122) & (g785)) + ((g18) & (g33) & (!sk[48]) & (g135) & (!g122) & (!g785)) + ((g18) & (g33) & (!sk[48]) & (g135) & (!g122) & (g785)) + ((g18) & (g33) & (!sk[48]) & (g135) & (g122) & (!g785)) + ((g18) & (g33) & (!sk[48]) & (g135) & (g122) & (g785)) + ((g18) & (g33) & (sk[48]) & (g135) & (!g122) & (!g785)));
	assign g787 = (((!g122) & (!g648) & (!g783) & (!g784) & (sk[49]) & (g786)) + ((!g122) & (!g648) & (g783) & (!g784) & (!sk[49]) & (g786)) + ((!g122) & (!g648) & (g783) & (g784) & (!sk[49]) & (!g786)) + ((!g122) & (!g648) & (g783) & (g784) & (!sk[49]) & (g786)) + ((!g122) & (g648) & (!g783) & (!g784) & (!sk[49]) & (!g786)) + ((!g122) & (g648) & (!g783) & (!g784) & (!sk[49]) & (g786)) + ((!g122) & (g648) & (!g783) & (!g784) & (sk[49]) & (g786)) + ((!g122) & (g648) & (!g783) & (g784) & (!sk[49]) & (!g786)) + ((!g122) & (g648) & (!g783) & (g784) & (!sk[49]) & (g786)) + ((!g122) & (g648) & (g783) & (!g784) & (!sk[49]) & (!g786)) + ((!g122) & (g648) & (g783) & (!g784) & (!sk[49]) & (g786)) + ((!g122) & (g648) & (g783) & (g784) & (!sk[49]) & (!g786)) + ((!g122) & (g648) & (g783) & (g784) & (!sk[49]) & (g786)) + ((g122) & (!g648) & (!g783) & (!g784) & (sk[49]) & (g786)) + ((g122) & (!g648) & (g783) & (!g784) & (!sk[49]) & (g786)) + ((g122) & (!g648) & (g783) & (g784) & (!sk[49]) & (!g786)) + ((g122) & (!g648) & (g783) & (g784) & (!sk[49]) & (g786)) + ((g122) & (g648) & (!g783) & (!g784) & (!sk[49]) & (!g786)) + ((g122) & (g648) & (!g783) & (!g784) & (!sk[49]) & (g786)) + ((g122) & (g648) & (!g783) & (g784) & (!sk[49]) & (!g786)) + ((g122) & (g648) & (!g783) & (g784) & (!sk[49]) & (g786)) + ((g122) & (g648) & (g783) & (!g784) & (!sk[49]) & (!g786)) + ((g122) & (g648) & (g783) & (!g784) & (!sk[49]) & (g786)) + ((g122) & (g648) & (g783) & (g784) & (!sk[49]) & (!g786)) + ((g122) & (g648) & (g783) & (g784) & (!sk[49]) & (g786)));
	assign g788 = (((!sk[50]) & (!g23) & (!g102) & (g684) & (!g703)) + ((!sk[50]) & (!g23) & (!g102) & (g684) & (g703)) + ((!sk[50]) & (!g23) & (g102) & (g684) & (!g703)) + ((!sk[50]) & (!g23) & (g102) & (g684) & (g703)) + ((!sk[50]) & (g23) & (!g102) & (g684) & (!g703)) + ((!sk[50]) & (g23) & (!g102) & (g684) & (g703)) + ((!sk[50]) & (g23) & (g102) & (g684) & (!g703)) + ((!sk[50]) & (g23) & (g102) & (g684) & (g703)) + ((sk[50]) & (!g23) & (g102) & (!g684) & (!g703)) + ((sk[50]) & (!g23) & (g102) & (!g684) & (g703)) + ((sk[50]) & (!g23) & (g102) & (g684) & (!g703)) + ((sk[50]) & (!g23) & (g102) & (g684) & (g703)) + ((sk[50]) & (g23) & (g102) & (!g684) & (!g703)) + ((sk[50]) & (g23) & (g102) & (!g684) & (g703)) + ((sk[50]) & (g23) & (g102) & (g684) & (!g703)));
	assign g789 = (((!g37) & (!g102) & (g105) & (!sk[51]) & (!g699) & (g700)) + ((!g37) & (!g102) & (g105) & (!sk[51]) & (g699) & (!g700)) + ((!g37) & (!g102) & (g105) & (!sk[51]) & (g699) & (g700)) + ((!g37) & (!g102) & (g105) & (sk[51]) & (!g699) & (!g700)) + ((!g37) & (!g102) & (g105) & (sk[51]) & (!g699) & (g700)) + ((!g37) & (!g102) & (g105) & (sk[51]) & (g699) & (!g700)) + ((!g37) & (!g102) & (g105) & (sk[51]) & (g699) & (g700)) + ((!g37) & (g102) & (!g105) & (!sk[51]) & (!g699) & (!g700)) + ((!g37) & (g102) & (!g105) & (!sk[51]) & (!g699) & (g700)) + ((!g37) & (g102) & (!g105) & (!sk[51]) & (g699) & (!g700)) + ((!g37) & (g102) & (!g105) & (!sk[51]) & (g699) & (g700)) + ((!g37) & (g102) & (g105) & (!sk[51]) & (!g699) & (!g700)) + ((!g37) & (g102) & (g105) & (!sk[51]) & (!g699) & (g700)) + ((!g37) & (g102) & (g105) & (!sk[51]) & (g699) & (!g700)) + ((!g37) & (g102) & (g105) & (!sk[51]) & (g699) & (g700)) + ((g37) & (!g102) & (!g105) & (sk[51]) & (g699) & (!g700)) + ((g37) & (!g102) & (!g105) & (sk[51]) & (g699) & (g700)) + ((g37) & (!g102) & (g105) & (!sk[51]) & (!g699) & (g700)) + ((g37) & (!g102) & (g105) & (!sk[51]) & (g699) & (!g700)) + ((g37) & (!g102) & (g105) & (!sk[51]) & (g699) & (g700)) + ((g37) & (!g102) & (g105) & (sk[51]) & (!g699) & (!g700)) + ((g37) & (!g102) & (g105) & (sk[51]) & (!g699) & (g700)) + ((g37) & (!g102) & (g105) & (sk[51]) & (g699) & (!g700)) + ((g37) & (!g102) & (g105) & (sk[51]) & (g699) & (g700)) + ((g37) & (g102) & (!g105) & (!sk[51]) & (!g699) & (!g700)) + ((g37) & (g102) & (!g105) & (!sk[51]) & (!g699) & (g700)) + ((g37) & (g102) & (!g105) & (!sk[51]) & (g699) & (!g700)) + ((g37) & (g102) & (!g105) & (!sk[51]) & (g699) & (g700)) + ((g37) & (g102) & (!g105) & (sk[51]) & (g699) & (g700)) + ((g37) & (g102) & (g105) & (!sk[51]) & (!g699) & (!g700)) + ((g37) & (g102) & (g105) & (!sk[51]) & (!g699) & (g700)) + ((g37) & (g102) & (g105) & (!sk[51]) & (g699) & (!g700)) + ((g37) & (g102) & (g105) & (!sk[51]) & (g699) & (g700)) + ((g37) & (g102) & (g105) & (sk[51]) & (g699) & (g700)));
	assign g790 = (((!g4) & (!g102) & (!sk[52]) & (g91) & (!g788) & (g789)) + ((!g4) & (!g102) & (!sk[52]) & (g91) & (g788) & (!g789)) + ((!g4) & (!g102) & (!sk[52]) & (g91) & (g788) & (g789)) + ((!g4) & (!g102) & (sk[52]) & (!g91) & (!g788) & (g789)) + ((!g4) & (!g102) & (sk[52]) & (g91) & (!g788) & (g789)) + ((!g4) & (g102) & (!sk[52]) & (!g91) & (!g788) & (!g789)) + ((!g4) & (g102) & (!sk[52]) & (!g91) & (!g788) & (g789)) + ((!g4) & (g102) & (!sk[52]) & (!g91) & (g788) & (!g789)) + ((!g4) & (g102) & (!sk[52]) & (!g91) & (g788) & (g789)) + ((!g4) & (g102) & (!sk[52]) & (g91) & (!g788) & (!g789)) + ((!g4) & (g102) & (!sk[52]) & (g91) & (!g788) & (g789)) + ((!g4) & (g102) & (!sk[52]) & (g91) & (g788) & (!g789)) + ((!g4) & (g102) & (!sk[52]) & (g91) & (g788) & (g789)) + ((!g4) & (g102) & (sk[52]) & (!g91) & (!g788) & (g789)) + ((!g4) & (g102) & (sk[52]) & (g91) & (!g788) & (g789)) + ((g4) & (!g102) & (!sk[52]) & (g91) & (!g788) & (g789)) + ((g4) & (!g102) & (!sk[52]) & (g91) & (g788) & (!g789)) + ((g4) & (!g102) & (!sk[52]) & (g91) & (g788) & (g789)) + ((g4) & (!g102) & (sk[52]) & (!g91) & (!g788) & (g789)) + ((g4) & (!g102) & (sk[52]) & (g91) & (!g788) & (g789)) + ((g4) & (g102) & (!sk[52]) & (!g91) & (!g788) & (!g789)) + ((g4) & (g102) & (!sk[52]) & (!g91) & (!g788) & (g789)) + ((g4) & (g102) & (!sk[52]) & (!g91) & (g788) & (!g789)) + ((g4) & (g102) & (!sk[52]) & (!g91) & (g788) & (g789)) + ((g4) & (g102) & (!sk[52]) & (g91) & (!g788) & (!g789)) + ((g4) & (g102) & (!sk[52]) & (g91) & (!g788) & (g789)) + ((g4) & (g102) & (!sk[52]) & (g91) & (g788) & (!g789)) + ((g4) & (g102) & (!sk[52]) & (g91) & (g788) & (g789)) + ((g4) & (g102) & (sk[52]) & (g91) & (!g788) & (g789)));
	assign g791 = (((!g144) & (!g164) & (!sk[53]) & (g684) & (!g703)) + ((!g144) & (!g164) & (!sk[53]) & (g684) & (g703)) + ((!g144) & (g164) & (!sk[53]) & (g684) & (!g703)) + ((!g144) & (g164) & (!sk[53]) & (g684) & (g703)) + ((!g144) & (g164) & (sk[53]) & (!g684) & (!g703)) + ((!g144) & (g164) & (sk[53]) & (!g684) & (g703)) + ((g144) & (!g164) & (!sk[53]) & (g684) & (!g703)) + ((g144) & (!g164) & (!sk[53]) & (g684) & (g703)) + ((g144) & (!g164) & (sk[53]) & (!g684) & (!g703)) + ((g144) & (!g164) & (sk[53]) & (g684) & (!g703)) + ((g144) & (g164) & (!sk[53]) & (g684) & (!g703)) + ((g144) & (g164) & (!sk[53]) & (g684) & (g703)) + ((g144) & (g164) & (sk[53]) & (!g684) & (!g703)) + ((g144) & (g164) & (sk[53]) & (!g684) & (g703)) + ((g144) & (g164) & (sk[53]) & (g684) & (!g703)));
	assign g792 = (((!sk[54]) & (!g19) & (!g126) & (g254) & (!g790) & (g791)) + ((!sk[54]) & (!g19) & (!g126) & (g254) & (g790) & (!g791)) + ((!sk[54]) & (!g19) & (!g126) & (g254) & (g790) & (g791)) + ((!sk[54]) & (!g19) & (g126) & (!g254) & (!g790) & (!g791)) + ((!sk[54]) & (!g19) & (g126) & (!g254) & (!g790) & (g791)) + ((!sk[54]) & (!g19) & (g126) & (!g254) & (g790) & (!g791)) + ((!sk[54]) & (!g19) & (g126) & (!g254) & (g790) & (g791)) + ((!sk[54]) & (!g19) & (g126) & (g254) & (!g790) & (!g791)) + ((!sk[54]) & (!g19) & (g126) & (g254) & (!g790) & (g791)) + ((!sk[54]) & (!g19) & (g126) & (g254) & (g790) & (!g791)) + ((!sk[54]) & (!g19) & (g126) & (g254) & (g790) & (g791)) + ((!sk[54]) & (g19) & (!g126) & (g254) & (!g790) & (g791)) + ((!sk[54]) & (g19) & (!g126) & (g254) & (g790) & (!g791)) + ((!sk[54]) & (g19) & (!g126) & (g254) & (g790) & (g791)) + ((!sk[54]) & (g19) & (g126) & (!g254) & (!g790) & (!g791)) + ((!sk[54]) & (g19) & (g126) & (!g254) & (!g790) & (g791)) + ((!sk[54]) & (g19) & (g126) & (!g254) & (g790) & (!g791)) + ((!sk[54]) & (g19) & (g126) & (!g254) & (g790) & (g791)) + ((!sk[54]) & (g19) & (g126) & (g254) & (!g790) & (!g791)) + ((!sk[54]) & (g19) & (g126) & (g254) & (!g790) & (g791)) + ((!sk[54]) & (g19) & (g126) & (g254) & (g790) & (!g791)) + ((!sk[54]) & (g19) & (g126) & (g254) & (g790) & (g791)) + ((sk[54]) & (!g19) & (!g126) & (!g254) & (g790) & (!g791)) + ((sk[54]) & (!g19) & (!g126) & (g254) & (g790) & (!g791)) + ((sk[54]) & (!g19) & (g126) & (!g254) & (g790) & (!g791)) + ((sk[54]) & (!g19) & (g126) & (g254) & (g790) & (!g791)) + ((sk[54]) & (g19) & (!g126) & (g254) & (g790) & (!g791)) + ((sk[54]) & (g19) & (g126) & (!g254) & (g790) & (!g791)) + ((sk[54]) & (g19) & (g126) & (g254) & (g790) & (!g791)));
	assign g793 = (((!g19) & (!sk[55]) & (!g126) & (g74) & (!g684)) + ((!g19) & (!sk[55]) & (!g126) & (g74) & (g684)) + ((!g19) & (!sk[55]) & (g126) & (g74) & (!g684)) + ((!g19) & (!sk[55]) & (g126) & (g74) & (g684)) + ((!g19) & (sk[55]) & (!g126) & (g74) & (!g684)) + ((!g19) & (sk[55]) & (g126) & (g74) & (!g684)) + ((g19) & (!sk[55]) & (!g126) & (g74) & (!g684)) + ((g19) & (!sk[55]) & (!g126) & (g74) & (g684)) + ((g19) & (!sk[55]) & (g126) & (g74) & (!g684)) + ((g19) & (!sk[55]) & (g126) & (g74) & (g684)) + ((g19) & (sk[55]) & (!g126) & (g74) & (!g684)) + ((g19) & (sk[55]) & (!g126) & (g74) & (g684)) + ((g19) & (sk[55]) & (g126) & (g74) & (!g684)));
	assign g794 = (((!sk[56]) & (!g4) & (!g75) & (g91) & (!g651)) + ((!sk[56]) & (!g4) & (!g75) & (g91) & (g651)) + ((!sk[56]) & (!g4) & (g75) & (g91) & (!g651)) + ((!sk[56]) & (!g4) & (g75) & (g91) & (g651)) + ((!sk[56]) & (g4) & (!g75) & (g91) & (!g651)) + ((!sk[56]) & (g4) & (!g75) & (g91) & (g651)) + ((!sk[56]) & (g4) & (g75) & (g91) & (!g651)) + ((!sk[56]) & (g4) & (g75) & (g91) & (g651)) + ((sk[56]) & (!g4) & (!g75) & (!g91) & (g651)) + ((sk[56]) & (!g4) & (!g75) & (g91) & (g651)) + ((sk[56]) & (g4) & (!g75) & (!g91) & (!g651)) + ((sk[56]) & (g4) & (!g75) & (!g91) & (g651)) + ((sk[56]) & (g4) & (!g75) & (g91) & (g651)));
	assign g795 = (((!sk[57]) & (!g21) & (!g49) & (g33) & (!g120) & (g648)) + ((!sk[57]) & (!g21) & (!g49) & (g33) & (g120) & (!g648)) + ((!sk[57]) & (!g21) & (!g49) & (g33) & (g120) & (g648)) + ((!sk[57]) & (!g21) & (g49) & (!g33) & (!g120) & (!g648)) + ((!sk[57]) & (!g21) & (g49) & (!g33) & (!g120) & (g648)) + ((!sk[57]) & (!g21) & (g49) & (!g33) & (g120) & (!g648)) + ((!sk[57]) & (!g21) & (g49) & (!g33) & (g120) & (g648)) + ((!sk[57]) & (!g21) & (g49) & (g33) & (!g120) & (!g648)) + ((!sk[57]) & (!g21) & (g49) & (g33) & (!g120) & (g648)) + ((!sk[57]) & (!g21) & (g49) & (g33) & (g120) & (!g648)) + ((!sk[57]) & (!g21) & (g49) & (g33) & (g120) & (g648)) + ((!sk[57]) & (g21) & (!g49) & (g33) & (!g120) & (g648)) + ((!sk[57]) & (g21) & (!g49) & (g33) & (g120) & (!g648)) + ((!sk[57]) & (g21) & (!g49) & (g33) & (g120) & (g648)) + ((!sk[57]) & (g21) & (g49) & (!g33) & (!g120) & (!g648)) + ((!sk[57]) & (g21) & (g49) & (!g33) & (!g120) & (g648)) + ((!sk[57]) & (g21) & (g49) & (!g33) & (g120) & (!g648)) + ((!sk[57]) & (g21) & (g49) & (!g33) & (g120) & (g648)) + ((!sk[57]) & (g21) & (g49) & (g33) & (!g120) & (!g648)) + ((!sk[57]) & (g21) & (g49) & (g33) & (!g120) & (g648)) + ((!sk[57]) & (g21) & (g49) & (g33) & (g120) & (!g648)) + ((!sk[57]) & (g21) & (g49) & (g33) & (g120) & (g648)) + ((sk[57]) & (!g21) & (g49) & (!g33) & (g120) & (g648)) + ((sk[57]) & (!g21) & (g49) & (g33) & (g120) & (!g648)) + ((sk[57]) & (!g21) & (g49) & (g33) & (g120) & (g648)) + ((sk[57]) & (g21) & (g49) & (!g33) & (g120) & (!g648)) + ((sk[57]) & (g21) & (g49) & (!g33) & (g120) & (g648)) + ((sk[57]) & (g21) & (g49) & (g33) & (g120) & (!g648)) + ((sk[57]) & (g21) & (g49) & (g33) & (g120) & (g648)));
	assign g796 = (((!sk[58]) & (!g634) & (!g131) & (g648) & (!g700) & (g795)) + ((!sk[58]) & (!g634) & (!g131) & (g648) & (g700) & (!g795)) + ((!sk[58]) & (!g634) & (!g131) & (g648) & (g700) & (g795)) + ((!sk[58]) & (!g634) & (g131) & (!g648) & (!g700) & (!g795)) + ((!sk[58]) & (!g634) & (g131) & (!g648) & (!g700) & (g795)) + ((!sk[58]) & (!g634) & (g131) & (!g648) & (g700) & (!g795)) + ((!sk[58]) & (!g634) & (g131) & (!g648) & (g700) & (g795)) + ((!sk[58]) & (!g634) & (g131) & (g648) & (!g700) & (!g795)) + ((!sk[58]) & (!g634) & (g131) & (g648) & (!g700) & (g795)) + ((!sk[58]) & (!g634) & (g131) & (g648) & (g700) & (!g795)) + ((!sk[58]) & (!g634) & (g131) & (g648) & (g700) & (g795)) + ((!sk[58]) & (g634) & (!g131) & (g648) & (!g700) & (g795)) + ((!sk[58]) & (g634) & (!g131) & (g648) & (g700) & (!g795)) + ((!sk[58]) & (g634) & (!g131) & (g648) & (g700) & (g795)) + ((!sk[58]) & (g634) & (g131) & (!g648) & (!g700) & (!g795)) + ((!sk[58]) & (g634) & (g131) & (!g648) & (!g700) & (g795)) + ((!sk[58]) & (g634) & (g131) & (!g648) & (g700) & (!g795)) + ((!sk[58]) & (g634) & (g131) & (!g648) & (g700) & (g795)) + ((!sk[58]) & (g634) & (g131) & (g648) & (!g700) & (!g795)) + ((!sk[58]) & (g634) & (g131) & (g648) & (!g700) & (g795)) + ((!sk[58]) & (g634) & (g131) & (g648) & (g700) & (!g795)) + ((!sk[58]) & (g634) & (g131) & (g648) & (g700) & (g795)) + ((sk[58]) & (!g634) & (g131) & (!g648) & (!g700) & (!g795)) + ((sk[58]) & (!g634) & (g131) & (!g648) & (g700) & (!g795)) + ((sk[58]) & (!g634) & (g131) & (g648) & (!g700) & (!g795)) + ((sk[58]) & (!g634) & (g131) & (g648) & (g700) & (!g795)) + ((sk[58]) & (g634) & (!g131) & (!g648) & (g700) & (!g795)) + ((sk[58]) & (g634) & (g131) & (!g648) & (!g700) & (!g795)) + ((sk[58]) & (g634) & (g131) & (!g648) & (g700) & (!g795)) + ((sk[58]) & (g634) & (g131) & (g648) & (!g700) & (!g795)) + ((sk[58]) & (g634) & (g131) & (g648) & (g700) & (!g795)));
	assign g797 = (((!g634) & (!g125) & (!g131) & (!g651) & (sk[59]) & (g796)) + ((!g634) & (!g125) & (g131) & (!g651) & (!sk[59]) & (g796)) + ((!g634) & (!g125) & (g131) & (!g651) & (sk[59]) & (g796)) + ((!g634) & (!g125) & (g131) & (g651) & (!sk[59]) & (!g796)) + ((!g634) & (!g125) & (g131) & (g651) & (!sk[59]) & (g796)) + ((!g634) & (!g125) & (g131) & (g651) & (sk[59]) & (g796)) + ((!g634) & (g125) & (!g131) & (!g651) & (!sk[59]) & (!g796)) + ((!g634) & (g125) & (!g131) & (!g651) & (!sk[59]) & (g796)) + ((!g634) & (g125) & (!g131) & (g651) & (!sk[59]) & (!g796)) + ((!g634) & (g125) & (!g131) & (g651) & (!sk[59]) & (g796)) + ((!g634) & (g125) & (g131) & (!g651) & (!sk[59]) & (!g796)) + ((!g634) & (g125) & (g131) & (!g651) & (!sk[59]) & (g796)) + ((!g634) & (g125) & (g131) & (g651) & (!sk[59]) & (!g796)) + ((!g634) & (g125) & (g131) & (g651) & (!sk[59]) & (g796)) + ((g634) & (!g125) & (!g131) & (!g651) & (sk[59]) & (g796)) + ((g634) & (!g125) & (g131) & (!g651) & (!sk[59]) & (g796)) + ((g634) & (!g125) & (g131) & (!g651) & (sk[59]) & (g796)) + ((g634) & (!g125) & (g131) & (g651) & (!sk[59]) & (!g796)) + ((g634) & (!g125) & (g131) & (g651) & (!sk[59]) & (g796)) + ((g634) & (!g125) & (g131) & (g651) & (sk[59]) & (g796)) + ((g634) & (g125) & (!g131) & (!g651) & (!sk[59]) & (!g796)) + ((g634) & (g125) & (!g131) & (!g651) & (!sk[59]) & (g796)) + ((g634) & (g125) & (!g131) & (!g651) & (sk[59]) & (g796)) + ((g634) & (g125) & (!g131) & (g651) & (!sk[59]) & (!g796)) + ((g634) & (g125) & (!g131) & (g651) & (!sk[59]) & (g796)) + ((g634) & (g125) & (g131) & (!g651) & (!sk[59]) & (!g796)) + ((g634) & (g125) & (g131) & (!g651) & (!sk[59]) & (g796)) + ((g634) & (g125) & (g131) & (!g651) & (sk[59]) & (g796)) + ((g634) & (g125) & (g131) & (g651) & (!sk[59]) & (!g796)) + ((g634) & (g125) & (g131) & (g651) & (!sk[59]) & (g796)) + ((g634) & (g125) & (g131) & (g651) & (sk[59]) & (g796)));
	assign g798 = (((!g21) & (!sk[60]) & (!g142) & (g227) & (!g668)) + ((!g21) & (!sk[60]) & (!g142) & (g227) & (g668)) + ((!g21) & (!sk[60]) & (g142) & (g227) & (!g668)) + ((!g21) & (!sk[60]) & (g142) & (g227) & (g668)) + ((!g21) & (sk[60]) & (!g142) & (g227) & (g668)) + ((!g21) & (sk[60]) & (g142) & (g227) & (g668)) + ((g21) & (!sk[60]) & (!g142) & (g227) & (!g668)) + ((g21) & (!sk[60]) & (!g142) & (g227) & (g668)) + ((g21) & (!sk[60]) & (g142) & (g227) & (!g668)) + ((g21) & (!sk[60]) & (g142) & (g227) & (g668)) + ((g21) & (sk[60]) & (!g142) & (!g227) & (!g668)) + ((g21) & (sk[60]) & (!g142) & (!g227) & (g668)) + ((g21) & (sk[60]) & (!g142) & (g227) & (!g668)) + ((g21) & (sk[60]) & (!g142) & (g227) & (g668)) + ((g21) & (sk[60]) & (g142) & (g227) & (g668)));
	assign g799 = (((!g23) & (!g123) & (!sk[61]) & (g684) & (!g703)) + ((!g23) & (!g123) & (!sk[61]) & (g684) & (g703)) + ((!g23) & (!g123) & (sk[61]) & (!g684) & (!g703)) + ((!g23) & (!g123) & (sk[61]) & (!g684) & (g703)) + ((!g23) & (!g123) & (sk[61]) & (g684) & (!g703)) + ((!g23) & (!g123) & (sk[61]) & (g684) & (g703)) + ((!g23) & (g123) & (!sk[61]) & (g684) & (!g703)) + ((!g23) & (g123) & (!sk[61]) & (g684) & (g703)) + ((g23) & (!g123) & (!sk[61]) & (g684) & (!g703)) + ((g23) & (!g123) & (!sk[61]) & (g684) & (g703)) + ((g23) & (!g123) & (sk[61]) & (!g684) & (!g703)) + ((g23) & (!g123) & (sk[61]) & (!g684) & (g703)) + ((g23) & (!g123) & (sk[61]) & (g684) & (!g703)) + ((g23) & (g123) & (!sk[61]) & (g684) & (!g703)) + ((g23) & (g123) & (!sk[61]) & (g684) & (g703)));
	assign g800 = (((!g18) & (!g23) & (!sk[62]) & (g105) & (!g684)) + ((!g18) & (!g23) & (!sk[62]) & (g105) & (g684)) + ((!g18) & (!g23) & (sk[62]) & (!g105) & (!g684)) + ((!g18) & (!g23) & (sk[62]) & (!g105) & (g684)) + ((!g18) & (g23) & (!sk[62]) & (g105) & (!g684)) + ((!g18) & (g23) & (!sk[62]) & (g105) & (g684)) + ((!g18) & (g23) & (sk[62]) & (!g105) & (!g684)) + ((g18) & (!g23) & (!sk[62]) & (g105) & (!g684)) + ((g18) & (!g23) & (!sk[62]) & (g105) & (g684)) + ((g18) & (!g23) & (sk[62]) & (!g105) & (!g684)) + ((g18) & (!g23) & (sk[62]) & (!g105) & (g684)) + ((g18) & (g23) & (!sk[62]) & (g105) & (!g684)) + ((g18) & (g23) & (!sk[62]) & (g105) & (g684)) + ((g18) & (g23) & (sk[62]) & (!g105) & (!g684)) + ((g18) & (g23) & (sk[62]) & (!g105) & (g684)));
	assign g801 = (((!g33) & (!g131) & (g225) & (!sk[63]) & (!g227)) + ((!g33) & (!g131) & (g225) & (!sk[63]) & (g227)) + ((!g33) & (g131) & (g225) & (!sk[63]) & (!g227)) + ((!g33) & (g131) & (g225) & (!sk[63]) & (g227)) + ((g33) & (!g131) & (!g225) & (sk[63]) & (!g227)) + ((g33) & (!g131) & (!g225) & (sk[63]) & (g227)) + ((g33) & (!g131) & (g225) & (!sk[63]) & (!g227)) + ((g33) & (!g131) & (g225) & (!sk[63]) & (g227)) + ((g33) & (!g131) & (g225) & (sk[63]) & (!g227)) + ((g33) & (!g131) & (g225) & (sk[63]) & (g227)) + ((g33) & (g131) & (!g225) & (sk[63]) & (g227)) + ((g33) & (g131) & (g225) & (!sk[63]) & (!g227)) + ((g33) & (g131) & (g225) & (!sk[63]) & (g227)) + ((g33) & (g131) & (g225) & (sk[63]) & (!g227)) + ((g33) & (g131) & (g225) & (sk[63]) & (g227)));
	assign g802 = (((!i_8_) & (!g73) & (g684) & (!sk[64]) & (!g703)) + ((!i_8_) & (!g73) & (g684) & (!sk[64]) & (g703)) + ((!i_8_) & (g73) & (g684) & (!sk[64]) & (!g703)) + ((!i_8_) & (g73) & (g684) & (!sk[64]) & (g703)) + ((i_8_) & (!g73) & (g684) & (!sk[64]) & (!g703)) + ((i_8_) & (!g73) & (g684) & (!sk[64]) & (g703)) + ((i_8_) & (g73) & (!g684) & (sk[64]) & (!g703)) + ((i_8_) & (g73) & (!g684) & (sk[64]) & (g703)) + ((i_8_) & (g73) & (g684) & (!sk[64]) & (!g703)) + ((i_8_) & (g73) & (g684) & (!sk[64]) & (g703)) + ((i_8_) & (g73) & (g684) & (sk[64]) & (!g703)));
	assign g803 = (((!g18) & (!sk[65]) & (!g102) & (g654)) + ((!g18) & (!sk[65]) & (g102) & (!g654)) + ((!g18) & (!sk[65]) & (g102) & (g654)) + ((!g18) & (sk[65]) & (g102) & (g654)) + ((g18) & (!sk[65]) & (!g102) & (g654)) + ((g18) & (!sk[65]) & (g102) & (!g654)) + ((g18) & (!sk[65]) & (g102) & (g654)) + ((g18) & (sk[65]) & (g102) & (!g654)) + ((g18) & (sk[65]) & (g102) & (g654)));
	assign g804 = (((!g23) & (!g130) & (!sk[66]) & (g699) & (!g703)) + ((!g23) & (!g130) & (!sk[66]) & (g699) & (g703)) + ((!g23) & (!g130) & (sk[66]) & (!g699) & (!g703)) + ((!g23) & (!g130) & (sk[66]) & (!g699) & (g703)) + ((!g23) & (!g130) & (sk[66]) & (g699) & (!g703)) + ((!g23) & (!g130) & (sk[66]) & (g699) & (g703)) + ((!g23) & (g130) & (!sk[66]) & (g699) & (!g703)) + ((!g23) & (g130) & (!sk[66]) & (g699) & (g703)) + ((g23) & (!g130) & (!sk[66]) & (g699) & (!g703)) + ((g23) & (!g130) & (!sk[66]) & (g699) & (g703)) + ((g23) & (!g130) & (sk[66]) & (!g699) & (!g703)) + ((g23) & (!g130) & (sk[66]) & (!g699) & (g703)) + ((g23) & (!g130) & (sk[66]) & (g699) & (!g703)) + ((g23) & (g130) & (!sk[66]) & (g699) & (!g703)) + ((g23) & (g130) & (!sk[66]) & (g699) & (g703)));
	assign g805 = (((!g799) & (!g800) & (!g801) & (!g802) & (!g803) & (!g804)));
	assign g806 = (((!sk[68]) & (!g18) & (!g33) & (g142)) + ((!sk[68]) & (!g18) & (g33) & (!g142)) + ((!sk[68]) & (!g18) & (g33) & (g142)) + ((!sk[68]) & (g18) & (!g33) & (g142)) + ((!sk[68]) & (g18) & (g33) & (!g142)) + ((!sk[68]) & (g18) & (g33) & (g142)) + ((sk[68]) & (!g18) & (g33) & (!g142)) + ((sk[68]) & (g18) & (!g33) & (!g142)) + ((sk[68]) & (g18) & (g33) & (!g142)));
	assign g807 = (((!g4) & (!g36) & (g91) & (!sk[69]) & (!g123) & (g130)) + ((!g4) & (!g36) & (g91) & (!sk[69]) & (g123) & (!g130)) + ((!g4) & (!g36) & (g91) & (!sk[69]) & (g123) & (g130)) + ((!g4) & (g36) & (!g91) & (!sk[69]) & (!g123) & (!g130)) + ((!g4) & (g36) & (!g91) & (!sk[69]) & (!g123) & (g130)) + ((!g4) & (g36) & (!g91) & (!sk[69]) & (g123) & (!g130)) + ((!g4) & (g36) & (!g91) & (!sk[69]) & (g123) & (g130)) + ((!g4) & (g36) & (g91) & (!sk[69]) & (!g123) & (!g130)) + ((!g4) & (g36) & (g91) & (!sk[69]) & (!g123) & (g130)) + ((!g4) & (g36) & (g91) & (!sk[69]) & (g123) & (!g130)) + ((!g4) & (g36) & (g91) & (!sk[69]) & (g123) & (g130)) + ((g4) & (!g36) & (!g91) & (sk[69]) & (!g123) & (!g130)) + ((g4) & (!g36) & (!g91) & (sk[69]) & (!g123) & (g130)) + ((g4) & (!g36) & (!g91) & (sk[69]) & (g123) & (!g130)) + ((g4) & (!g36) & (g91) & (!sk[69]) & (!g123) & (g130)) + ((g4) & (!g36) & (g91) & (!sk[69]) & (g123) & (!g130)) + ((g4) & (!g36) & (g91) & (!sk[69]) & (g123) & (g130)) + ((g4) & (g36) & (!g91) & (!sk[69]) & (!g123) & (!g130)) + ((g4) & (g36) & (!g91) & (!sk[69]) & (!g123) & (g130)) + ((g4) & (g36) & (!g91) & (!sk[69]) & (g123) & (!g130)) + ((g4) & (g36) & (!g91) & (!sk[69]) & (g123) & (g130)) + ((g4) & (g36) & (!g91) & (sk[69]) & (!g123) & (!g130)) + ((g4) & (g36) & (!g91) & (sk[69]) & (!g123) & (g130)) + ((g4) & (g36) & (!g91) & (sk[69]) & (g123) & (!g130)) + ((g4) & (g36) & (g91) & (!sk[69]) & (!g123) & (!g130)) + ((g4) & (g36) & (g91) & (!sk[69]) & (!g123) & (g130)) + ((g4) & (g36) & (g91) & (!sk[69]) & (g123) & (!g130)) + ((g4) & (g36) & (g91) & (!sk[69]) & (g123) & (g130)) + ((g4) & (g36) & (g91) & (sk[69]) & (!g123) & (!g130)) + ((g4) & (g36) & (g91) & (sk[69]) & (!g123) & (g130)) + ((g4) & (g36) & (g91) & (sk[69]) & (g123) & (!g130)));
	assign g808 = (((!g125) & (!g122) & (!g105) & (!g651) & (!g700) & (g703)) + ((!g125) & (!g122) & (!g105) & (!g651) & (g700) & (g703)) + ((!g125) & (!g122) & (!g105) & (g651) & (!g700) & (g703)) + ((!g125) & (!g122) & (!g105) & (g651) & (g700) & (g703)) + ((!g125) & (!g122) & (g105) & (!g651) & (!g700) & (!g703)) + ((!g125) & (!g122) & (g105) & (!g651) & (!g700) & (g703)) + ((!g125) & (!g122) & (g105) & (!g651) & (g700) & (!g703)) + ((!g125) & (!g122) & (g105) & (!g651) & (g700) & (g703)) + ((!g125) & (!g122) & (g105) & (g651) & (!g700) & (!g703)) + ((!g125) & (!g122) & (g105) & (g651) & (!g700) & (g703)) + ((!g125) & (!g122) & (g105) & (g651) & (g700) & (!g703)) + ((!g125) & (!g122) & (g105) & (g651) & (g700) & (g703)) + ((!g125) & (g122) & (!g105) & (!g651) & (!g700) & (g703)) + ((!g125) & (g122) & (!g105) & (!g651) & (g700) & (g703)) + ((!g125) & (g122) & (g105) & (!g651) & (!g700) & (g703)) + ((!g125) & (g122) & (g105) & (!g651) & (g700) & (g703)) + ((g125) & (!g122) & (!g105) & (!g651) & (g700) & (g703)) + ((g125) & (!g122) & (g105) & (!g651) & (g700) & (!g703)) + ((g125) & (!g122) & (g105) & (!g651) & (g700) & (g703)) + ((g125) & (g122) & (!g105) & (!g651) & (g700) & (g703)) + ((g125) & (g122) & (g105) & (!g651) & (g700) & (g703)));
	assign g809 = (((!g142) & (g699) & (g700) & (!g806) & (!g807) & (g808)) + ((g142) & (!g699) & (!g700) & (!g806) & (!g807) & (g808)) + ((g142) & (!g699) & (g700) & (!g806) & (!g807) & (g808)) + ((g142) & (g699) & (!g700) & (!g806) & (!g807) & (g808)) + ((g142) & (g699) & (g700) & (!g806) & (!g807) & (g808)));
	assign g810 = (((!g793) & (!g794) & (g797) & (!g798) & (g805) & (g809)));
	assign g811 = (((g211) & (g216) & (g252) & (g787) & (g792) & (g810)));
	assign g812 = (((g623) & (g697) & (g711) & (g781) & (g782) & (g811)));
	assign g813 = (((!g581) & (!g589) & (!sk[75]) & (g596)) + ((!g581) & (g589) & (!sk[75]) & (!g596)) + ((!g581) & (g589) & (!sk[75]) & (g596)) + ((g581) & (!g589) & (!sk[75]) & (g596)) + ((g581) & (g589) & (!sk[75]) & (!g596)) + ((g581) & (g589) & (!sk[75]) & (g596)) + ((g581) & (g589) & (sk[75]) & (g596)));
	assign g814 = (((!g712) & (!sk[76]) & (!g713) & (g714) & (!g717) & (g718)) + ((!g712) & (!sk[76]) & (!g713) & (g714) & (g717) & (!g718)) + ((!g712) & (!sk[76]) & (!g713) & (g714) & (g717) & (g718)) + ((!g712) & (!sk[76]) & (g713) & (!g714) & (!g717) & (!g718)) + ((!g712) & (!sk[76]) & (g713) & (!g714) & (!g717) & (g718)) + ((!g712) & (!sk[76]) & (g713) & (!g714) & (g717) & (!g718)) + ((!g712) & (!sk[76]) & (g713) & (!g714) & (g717) & (g718)) + ((!g712) & (!sk[76]) & (g713) & (g714) & (!g717) & (!g718)) + ((!g712) & (!sk[76]) & (g713) & (g714) & (!g717) & (g718)) + ((!g712) & (!sk[76]) & (g713) & (g714) & (g717) & (!g718)) + ((!g712) & (!sk[76]) & (g713) & (g714) & (g717) & (g718)) + ((!g712) & (sk[76]) & (!g713) & (!g714) & (g717) & (!g718)) + ((g712) & (!sk[76]) & (!g713) & (g714) & (!g717) & (g718)) + ((g712) & (!sk[76]) & (!g713) & (g714) & (g717) & (!g718)) + ((g712) & (!sk[76]) & (!g713) & (g714) & (g717) & (g718)) + ((g712) & (!sk[76]) & (g713) & (!g714) & (!g717) & (!g718)) + ((g712) & (!sk[76]) & (g713) & (!g714) & (!g717) & (g718)) + ((g712) & (!sk[76]) & (g713) & (!g714) & (g717) & (!g718)) + ((g712) & (!sk[76]) & (g713) & (!g714) & (g717) & (g718)) + ((g712) & (!sk[76]) & (g713) & (g714) & (!g717) & (!g718)) + ((g712) & (!sk[76]) & (g713) & (g714) & (!g717) & (g718)) + ((g712) & (!sk[76]) & (g713) & (g714) & (g717) & (!g718)) + ((g712) & (!sk[76]) & (g713) & (g714) & (g717) & (g718)));
	assign g815 = (((!i_11_) & (!i_15_) & (g19) & (!sk[77]) & (!g53) & (g105)) + ((!i_11_) & (!i_15_) & (g19) & (!sk[77]) & (g53) & (!g105)) + ((!i_11_) & (!i_15_) & (g19) & (!sk[77]) & (g53) & (g105)) + ((!i_11_) & (i_15_) & (!g19) & (!sk[77]) & (!g53) & (!g105)) + ((!i_11_) & (i_15_) & (!g19) & (!sk[77]) & (!g53) & (g105)) + ((!i_11_) & (i_15_) & (!g19) & (!sk[77]) & (g53) & (!g105)) + ((!i_11_) & (i_15_) & (!g19) & (!sk[77]) & (g53) & (g105)) + ((!i_11_) & (i_15_) & (g19) & (!sk[77]) & (!g53) & (!g105)) + ((!i_11_) & (i_15_) & (g19) & (!sk[77]) & (!g53) & (g105)) + ((!i_11_) & (i_15_) & (g19) & (!sk[77]) & (g53) & (!g105)) + ((!i_11_) & (i_15_) & (g19) & (!sk[77]) & (g53) & (g105)) + ((i_11_) & (!i_15_) & (g19) & (!sk[77]) & (!g53) & (g105)) + ((i_11_) & (!i_15_) & (g19) & (!sk[77]) & (g53) & (!g105)) + ((i_11_) & (!i_15_) & (g19) & (!sk[77]) & (g53) & (g105)) + ((i_11_) & (!i_15_) & (g19) & (sk[77]) & (g53) & (!g105)) + ((i_11_) & (i_15_) & (!g19) & (!sk[77]) & (!g53) & (!g105)) + ((i_11_) & (i_15_) & (!g19) & (!sk[77]) & (!g53) & (g105)) + ((i_11_) & (i_15_) & (!g19) & (!sk[77]) & (g53) & (!g105)) + ((i_11_) & (i_15_) & (!g19) & (!sk[77]) & (g53) & (g105)) + ((i_11_) & (i_15_) & (g19) & (!sk[77]) & (!g53) & (!g105)) + ((i_11_) & (i_15_) & (g19) & (!sk[77]) & (!g53) & (g105)) + ((i_11_) & (i_15_) & (g19) & (!sk[77]) & (g53) & (!g105)) + ((i_11_) & (i_15_) & (g19) & (!sk[77]) & (g53) & (g105)));
	assign g816 = (((!sk[78]) & (!g112) & (!g154) & (g130)) + ((!sk[78]) & (!g112) & (g154) & (!g130)) + ((!sk[78]) & (!g112) & (g154) & (g130)) + ((!sk[78]) & (g112) & (!g154) & (g130)) + ((!sk[78]) & (g112) & (g154) & (!g130)) + ((!sk[78]) & (g112) & (g154) & (g130)) + ((sk[78]) & (g112) & (!g154) & (!g130)) + ((sk[78]) & (g112) & (!g154) & (g130)) + ((sk[78]) & (g112) & (g154) & (!g130)));
	assign g817 = (((!i_15_) & (!sk[79]) & (!g4) & (g34) & (!g155) & (g816)) + ((!i_15_) & (!sk[79]) & (!g4) & (g34) & (g155) & (!g816)) + ((!i_15_) & (!sk[79]) & (!g4) & (g34) & (g155) & (g816)) + ((!i_15_) & (!sk[79]) & (g4) & (!g34) & (!g155) & (!g816)) + ((!i_15_) & (!sk[79]) & (g4) & (!g34) & (!g155) & (g816)) + ((!i_15_) & (!sk[79]) & (g4) & (!g34) & (g155) & (!g816)) + ((!i_15_) & (!sk[79]) & (g4) & (!g34) & (g155) & (g816)) + ((!i_15_) & (!sk[79]) & (g4) & (g34) & (!g155) & (!g816)) + ((!i_15_) & (!sk[79]) & (g4) & (g34) & (!g155) & (g816)) + ((!i_15_) & (!sk[79]) & (g4) & (g34) & (g155) & (!g816)) + ((!i_15_) & (!sk[79]) & (g4) & (g34) & (g155) & (g816)) + ((i_15_) & (!sk[79]) & (!g4) & (g34) & (!g155) & (g816)) + ((i_15_) & (!sk[79]) & (!g4) & (g34) & (g155) & (!g816)) + ((i_15_) & (!sk[79]) & (!g4) & (g34) & (g155) & (g816)) + ((i_15_) & (!sk[79]) & (g4) & (!g34) & (!g155) & (!g816)) + ((i_15_) & (!sk[79]) & (g4) & (!g34) & (!g155) & (g816)) + ((i_15_) & (!sk[79]) & (g4) & (!g34) & (g155) & (!g816)) + ((i_15_) & (!sk[79]) & (g4) & (!g34) & (g155) & (g816)) + ((i_15_) & (!sk[79]) & (g4) & (g34) & (!g155) & (!g816)) + ((i_15_) & (!sk[79]) & (g4) & (g34) & (!g155) & (g816)) + ((i_15_) & (!sk[79]) & (g4) & (g34) & (g155) & (!g816)) + ((i_15_) & (!sk[79]) & (g4) & (g34) & (g155) & (g816)) + ((i_15_) & (sk[79]) & (g4) & (!g34) & (!g155) & (g816)) + ((i_15_) & (sk[79]) & (g4) & (!g34) & (g155) & (g816)) + ((i_15_) & (sk[79]) & (g4) & (g34) & (!g155) & (!g816)) + ((i_15_) & (sk[79]) & (g4) & (g34) & (!g155) & (g816)) + ((i_15_) & (sk[79]) & (g4) & (g34) & (g155) & (g816)));
	assign g818 = (((!sk[80]) & (!i_9_) & (!i_11_) & (i_15_) & (!g4)) + ((!sk[80]) & (!i_9_) & (!i_11_) & (i_15_) & (g4)) + ((!sk[80]) & (!i_9_) & (i_11_) & (i_15_) & (!g4)) + ((!sk[80]) & (!i_9_) & (i_11_) & (i_15_) & (g4)) + ((!sk[80]) & (i_9_) & (!i_11_) & (i_15_) & (!g4)) + ((!sk[80]) & (i_9_) & (!i_11_) & (i_15_) & (g4)) + ((!sk[80]) & (i_9_) & (i_11_) & (i_15_) & (!g4)) + ((!sk[80]) & (i_9_) & (i_11_) & (i_15_) & (g4)) + ((sk[80]) & (!i_9_) & (!i_11_) & (i_15_) & (g4)));
	assign g819 = (((!sk[81]) & (!g125) & (!g159) & (g703) & (!g818)) + ((!sk[81]) & (!g125) & (!g159) & (g703) & (g818)) + ((!sk[81]) & (!g125) & (g159) & (g703) & (!g818)) + ((!sk[81]) & (!g125) & (g159) & (g703) & (g818)) + ((!sk[81]) & (g125) & (!g159) & (g703) & (!g818)) + ((!sk[81]) & (g125) & (!g159) & (g703) & (g818)) + ((!sk[81]) & (g125) & (g159) & (g703) & (!g818)) + ((!sk[81]) & (g125) & (g159) & (g703) & (g818)) + ((sk[81]) & (!g125) & (!g159) & (!g703) & (!g818)) + ((sk[81]) & (!g125) & (!g159) & (!g703) & (g818)) + ((sk[81]) & (g125) & (!g159) & (!g703) & (!g818)) + ((sk[81]) & (g125) & (!g159) & (!g703) & (g818)) + ((sk[81]) & (g125) & (!g159) & (g703) & (g818)) + ((sk[81]) & (g125) & (g159) & (!g703) & (g818)) + ((sk[81]) & (g125) & (g159) & (g703) & (g818)));
	assign g820 = (((!g19) & (!g27) & (g102) & (!sk[82]) & (!g165) & (g324)) + ((!g19) & (!g27) & (g102) & (!sk[82]) & (g165) & (!g324)) + ((!g19) & (!g27) & (g102) & (!sk[82]) & (g165) & (g324)) + ((!g19) & (g27) & (!g102) & (!sk[82]) & (!g165) & (!g324)) + ((!g19) & (g27) & (!g102) & (!sk[82]) & (!g165) & (g324)) + ((!g19) & (g27) & (!g102) & (!sk[82]) & (g165) & (!g324)) + ((!g19) & (g27) & (!g102) & (!sk[82]) & (g165) & (g324)) + ((!g19) & (g27) & (g102) & (!sk[82]) & (!g165) & (!g324)) + ((!g19) & (g27) & (g102) & (!sk[82]) & (!g165) & (g324)) + ((!g19) & (g27) & (g102) & (!sk[82]) & (g165) & (!g324)) + ((!g19) & (g27) & (g102) & (!sk[82]) & (g165) & (g324)) + ((g19) & (!g27) & (!g102) & (sk[82]) & (g165) & (g324)) + ((g19) & (!g27) & (g102) & (!sk[82]) & (!g165) & (g324)) + ((g19) & (!g27) & (g102) & (!sk[82]) & (g165) & (!g324)) + ((g19) & (!g27) & (g102) & (!sk[82]) & (g165) & (g324)) + ((g19) & (!g27) & (g102) & (sk[82]) & (g165) & (g324)) + ((g19) & (g27) & (!g102) & (!sk[82]) & (!g165) & (!g324)) + ((g19) & (g27) & (!g102) & (!sk[82]) & (!g165) & (g324)) + ((g19) & (g27) & (!g102) & (!sk[82]) & (g165) & (!g324)) + ((g19) & (g27) & (!g102) & (!sk[82]) & (g165) & (g324)) + ((g19) & (g27) & (!g102) & (sk[82]) & (g165) & (g324)) + ((g19) & (g27) & (g102) & (!sk[82]) & (!g165) & (!g324)) + ((g19) & (g27) & (g102) & (!sk[82]) & (!g165) & (g324)) + ((g19) & (g27) & (g102) & (!sk[82]) & (g165) & (!g324)) + ((g19) & (g27) & (g102) & (!sk[82]) & (g165) & (g324)) + ((g19) & (g27) & (g102) & (sk[82]) & (!g165) & (!g324)) + ((g19) & (g27) & (g102) & (sk[82]) & (!g165) & (g324)) + ((g19) & (g27) & (g102) & (sk[82]) & (g165) & (!g324)) + ((g19) & (g27) & (g102) & (sk[82]) & (g165) & (g324)));
	assign g821 = (((!g21) & (!sk[83]) & (!g164) & (g105) & (!g819) & (g820)) + ((!g21) & (!sk[83]) & (!g164) & (g105) & (g819) & (!g820)) + ((!g21) & (!sk[83]) & (!g164) & (g105) & (g819) & (g820)) + ((!g21) & (!sk[83]) & (g164) & (!g105) & (!g819) & (!g820)) + ((!g21) & (!sk[83]) & (g164) & (!g105) & (!g819) & (g820)) + ((!g21) & (!sk[83]) & (g164) & (!g105) & (g819) & (!g820)) + ((!g21) & (!sk[83]) & (g164) & (!g105) & (g819) & (g820)) + ((!g21) & (!sk[83]) & (g164) & (g105) & (!g819) & (!g820)) + ((!g21) & (!sk[83]) & (g164) & (g105) & (!g819) & (g820)) + ((!g21) & (!sk[83]) & (g164) & (g105) & (g819) & (!g820)) + ((!g21) & (!sk[83]) & (g164) & (g105) & (g819) & (g820)) + ((!g21) & (sk[83]) & (!g164) & (!g105) & (!g819) & (!g820)) + ((!g21) & (sk[83]) & (!g164) & (g105) & (!g819) & (!g820)) + ((!g21) & (sk[83]) & (g164) & (!g105) & (!g819) & (!g820)) + ((!g21) & (sk[83]) & (g164) & (g105) & (!g819) & (!g820)) + ((g21) & (!sk[83]) & (!g164) & (g105) & (!g819) & (g820)) + ((g21) & (!sk[83]) & (!g164) & (g105) & (g819) & (!g820)) + ((g21) & (!sk[83]) & (!g164) & (g105) & (g819) & (g820)) + ((g21) & (!sk[83]) & (g164) & (!g105) & (!g819) & (!g820)) + ((g21) & (!sk[83]) & (g164) & (!g105) & (!g819) & (g820)) + ((g21) & (!sk[83]) & (g164) & (!g105) & (g819) & (!g820)) + ((g21) & (!sk[83]) & (g164) & (!g105) & (g819) & (g820)) + ((g21) & (!sk[83]) & (g164) & (g105) & (!g819) & (!g820)) + ((g21) & (!sk[83]) & (g164) & (g105) & (!g819) & (g820)) + ((g21) & (!sk[83]) & (g164) & (g105) & (g819) & (!g820)) + ((g21) & (!sk[83]) & (g164) & (g105) & (g819) & (g820)) + ((g21) & (sk[83]) & (!g164) & (g105) & (!g819) & (!g820)));
	assign g822 = (((!g18) & (!g167) & (!g815) & (!g817) & (sk[84]) & (g821)) + ((!g18) & (!g167) & (g815) & (!g817) & (!sk[84]) & (g821)) + ((!g18) & (!g167) & (g815) & (g817) & (!sk[84]) & (!g821)) + ((!g18) & (!g167) & (g815) & (g817) & (!sk[84]) & (g821)) + ((!g18) & (g167) & (!g815) & (!g817) & (!sk[84]) & (!g821)) + ((!g18) & (g167) & (!g815) & (!g817) & (!sk[84]) & (g821)) + ((!g18) & (g167) & (!g815) & (!g817) & (sk[84]) & (g821)) + ((!g18) & (g167) & (!g815) & (g817) & (!sk[84]) & (!g821)) + ((!g18) & (g167) & (!g815) & (g817) & (!sk[84]) & (g821)) + ((!g18) & (g167) & (g815) & (!g817) & (!sk[84]) & (!g821)) + ((!g18) & (g167) & (g815) & (!g817) & (!sk[84]) & (g821)) + ((!g18) & (g167) & (g815) & (g817) & (!sk[84]) & (!g821)) + ((!g18) & (g167) & (g815) & (g817) & (!sk[84]) & (g821)) + ((g18) & (!g167) & (!g815) & (!g817) & (sk[84]) & (g821)) + ((g18) & (!g167) & (g815) & (!g817) & (!sk[84]) & (g821)) + ((g18) & (!g167) & (g815) & (g817) & (!sk[84]) & (!g821)) + ((g18) & (!g167) & (g815) & (g817) & (!sk[84]) & (g821)) + ((g18) & (g167) & (!g815) & (!g817) & (!sk[84]) & (!g821)) + ((g18) & (g167) & (!g815) & (!g817) & (!sk[84]) & (g821)) + ((g18) & (g167) & (!g815) & (g817) & (!sk[84]) & (!g821)) + ((g18) & (g167) & (!g815) & (g817) & (!sk[84]) & (g821)) + ((g18) & (g167) & (g815) & (!g817) & (!sk[84]) & (!g821)) + ((g18) & (g167) & (g815) & (!g817) & (!sk[84]) & (g821)) + ((g18) & (g167) & (g815) & (g817) & (!sk[84]) & (!g821)) + ((g18) & (g167) & (g815) & (g817) & (!sk[84]) & (g821)));
	assign g823 = (((g814) & (g707) & (g787) & (g792) & (g810) & (g822)));
	assign g824 = (((g80) & (!i_11_) & (i_15_) & (!g76) & (!g414) & (!g447)) + ((g80) & (!i_11_) & (i_15_) & (!g76) & (!g414) & (g447)) + ((g80) & (i_11_) & (i_15_) & (!g76) & (!g414) & (!g447)) + ((g80) & (i_11_) & (i_15_) & (!g76) & (g414) & (!g447)));
	assign g825 = (((!g164) & (!sk[87]) & (!g105) & (g562)) + ((!g164) & (!sk[87]) & (g105) & (!g562)) + ((!g164) & (!sk[87]) & (g105) & (g562)) + ((!g164) & (sk[87]) & (!g105) & (g562)) + ((g164) & (!sk[87]) & (!g105) & (g562)) + ((g164) & (!sk[87]) & (g105) & (!g562)) + ((g164) & (!sk[87]) & (g105) & (g562)) + ((g164) & (sk[87]) & (!g105) & (g562)) + ((g164) & (sk[87]) & (g105) & (g562)));
	assign g826 = (((!sk[88]) & (!g87) & (!g154) & (g557) & (!g518)) + ((!sk[88]) & (!g87) & (!g154) & (g557) & (g518)) + ((!sk[88]) & (!g87) & (g154) & (g557) & (!g518)) + ((!sk[88]) & (!g87) & (g154) & (g557) & (g518)) + ((!sk[88]) & (g87) & (!g154) & (g557) & (!g518)) + ((!sk[88]) & (g87) & (!g154) & (g557) & (g518)) + ((!sk[88]) & (g87) & (g154) & (g557) & (!g518)) + ((!sk[88]) & (g87) & (g154) & (g557) & (g518)) + ((sk[88]) & (!g87) & (!g154) & (!g557) & (g518)) + ((sk[88]) & (!g87) & (!g154) & (g557) & (!g518)) + ((sk[88]) & (!g87) & (!g154) & (g557) & (g518)) + ((sk[88]) & (!g87) & (g154) & (!g557) & (g518)) + ((sk[88]) & (!g87) & (g154) & (g557) & (g518)) + ((sk[88]) & (g87) & (!g154) & (g557) & (!g518)) + ((sk[88]) & (g87) & (!g154) & (g557) & (g518)));
	assign g827 = (((!g17) & (!g76) & (!g107) & (!g168) & (sk[89]) & (!g105)) + ((!g17) & (!g76) & (!g107) & (g168) & (sk[89]) & (!g105)) + ((!g17) & (!g76) & (g107) & (!g168) & (!sk[89]) & (g105)) + ((!g17) & (!g76) & (g107) & (g168) & (!sk[89]) & (!g105)) + ((!g17) & (!g76) & (g107) & (g168) & (!sk[89]) & (g105)) + ((!g17) & (g76) & (!g107) & (!g168) & (!sk[89]) & (!g105)) + ((!g17) & (g76) & (!g107) & (!g168) & (!sk[89]) & (g105)) + ((!g17) & (g76) & (!g107) & (g168) & (!sk[89]) & (!g105)) + ((!g17) & (g76) & (!g107) & (g168) & (!sk[89]) & (g105)) + ((!g17) & (g76) & (g107) & (!g168) & (!sk[89]) & (!g105)) + ((!g17) & (g76) & (g107) & (!g168) & (!sk[89]) & (g105)) + ((!g17) & (g76) & (g107) & (g168) & (!sk[89]) & (!g105)) + ((!g17) & (g76) & (g107) & (g168) & (!sk[89]) & (g105)) + ((g17) & (!g76) & (!g107) & (!g168) & (sk[89]) & (!g105)) + ((g17) & (!g76) & (!g107) & (g168) & (sk[89]) & (!g105)) + ((g17) & (!g76) & (!g107) & (g168) & (sk[89]) & (g105)) + ((g17) & (!g76) & (g107) & (!g168) & (!sk[89]) & (g105)) + ((g17) & (!g76) & (g107) & (g168) & (!sk[89]) & (!g105)) + ((g17) & (!g76) & (g107) & (g168) & (!sk[89]) & (g105)) + ((g17) & (!g76) & (g107) & (g168) & (sk[89]) & (!g105)) + ((g17) & (!g76) & (g107) & (g168) & (sk[89]) & (g105)) + ((g17) & (g76) & (!g107) & (!g168) & (!sk[89]) & (!g105)) + ((g17) & (g76) & (!g107) & (!g168) & (!sk[89]) & (g105)) + ((g17) & (g76) & (!g107) & (g168) & (!sk[89]) & (!g105)) + ((g17) & (g76) & (!g107) & (g168) & (!sk[89]) & (g105)) + ((g17) & (g76) & (g107) & (!g168) & (!sk[89]) & (!g105)) + ((g17) & (g76) & (g107) & (!g168) & (!sk[89]) & (g105)) + ((g17) & (g76) & (g107) & (g168) & (!sk[89]) & (!g105)) + ((g17) & (g76) & (g107) & (g168) & (!sk[89]) & (g105)));
	assign g828 = (((!i_6_) & (!g120) & (!sk[90]) & (g159) & (!g562) & (g751)) + ((!i_6_) & (!g120) & (!sk[90]) & (g159) & (g562) & (!g751)) + ((!i_6_) & (!g120) & (!sk[90]) & (g159) & (g562) & (g751)) + ((!i_6_) & (!g120) & (sk[90]) & (!g159) & (g562) & (!g751)) + ((!i_6_) & (!g120) & (sk[90]) & (!g159) & (g562) & (g751)) + ((!i_6_) & (g120) & (!sk[90]) & (!g159) & (!g562) & (!g751)) + ((!i_6_) & (g120) & (!sk[90]) & (!g159) & (!g562) & (g751)) + ((!i_6_) & (g120) & (!sk[90]) & (!g159) & (g562) & (!g751)) + ((!i_6_) & (g120) & (!sk[90]) & (!g159) & (g562) & (g751)) + ((!i_6_) & (g120) & (!sk[90]) & (g159) & (!g562) & (!g751)) + ((!i_6_) & (g120) & (!sk[90]) & (g159) & (!g562) & (g751)) + ((!i_6_) & (g120) & (!sk[90]) & (g159) & (g562) & (!g751)) + ((!i_6_) & (g120) & (!sk[90]) & (g159) & (g562) & (g751)) + ((!i_6_) & (g120) & (sk[90]) & (!g159) & (!g562) & (g751)) + ((!i_6_) & (g120) & (sk[90]) & (!g159) & (g562) & (!g751)) + ((!i_6_) & (g120) & (sk[90]) & (!g159) & (g562) & (g751)) + ((!i_6_) & (g120) & (sk[90]) & (g159) & (!g562) & (g751)) + ((!i_6_) & (g120) & (sk[90]) & (g159) & (g562) & (g751)) + ((i_6_) & (!g120) & (!sk[90]) & (g159) & (!g562) & (g751)) + ((i_6_) & (!g120) & (!sk[90]) & (g159) & (g562) & (!g751)) + ((i_6_) & (!g120) & (!sk[90]) & (g159) & (g562) & (g751)) + ((i_6_) & (!g120) & (sk[90]) & (!g159) & (g562) & (!g751)) + ((i_6_) & (!g120) & (sk[90]) & (!g159) & (g562) & (g751)) + ((i_6_) & (g120) & (!sk[90]) & (!g159) & (!g562) & (!g751)) + ((i_6_) & (g120) & (!sk[90]) & (!g159) & (!g562) & (g751)) + ((i_6_) & (g120) & (!sk[90]) & (!g159) & (g562) & (!g751)) + ((i_6_) & (g120) & (!sk[90]) & (!g159) & (g562) & (g751)) + ((i_6_) & (g120) & (!sk[90]) & (g159) & (!g562) & (!g751)) + ((i_6_) & (g120) & (!sk[90]) & (g159) & (!g562) & (g751)) + ((i_6_) & (g120) & (!sk[90]) & (g159) & (g562) & (!g751)) + ((i_6_) & (g120) & (!sk[90]) & (g159) & (g562) & (g751)) + ((i_6_) & (g120) & (sk[90]) & (!g159) & (g562) & (!g751)) + ((i_6_) & (g120) & (sk[90]) & (!g159) & (g562) & (g751)));
	assign g829 = (((!g159) & (g89) & (g684) & (!g826) & (!g827) & (!g828)) + ((g159) & (!g89) & (!g684) & (!g826) & (!g827) & (!g828)) + ((g159) & (!g89) & (g684) & (!g826) & (!g827) & (!g828)) + ((g159) & (g89) & (!g684) & (!g826) & (!g827) & (!g828)) + ((g159) & (g89) & (g684) & (!g826) & (!g827) & (!g828)));
	assign g830 = (((!g125) & (!sk[92]) & (!g165) & (g495) & (!g825) & (g829)) + ((!g125) & (!sk[92]) & (!g165) & (g495) & (g825) & (!g829)) + ((!g125) & (!sk[92]) & (!g165) & (g495) & (g825) & (g829)) + ((!g125) & (!sk[92]) & (g165) & (!g495) & (!g825) & (!g829)) + ((!g125) & (!sk[92]) & (g165) & (!g495) & (!g825) & (g829)) + ((!g125) & (!sk[92]) & (g165) & (!g495) & (g825) & (!g829)) + ((!g125) & (!sk[92]) & (g165) & (!g495) & (g825) & (g829)) + ((!g125) & (!sk[92]) & (g165) & (g495) & (!g825) & (!g829)) + ((!g125) & (!sk[92]) & (g165) & (g495) & (!g825) & (g829)) + ((!g125) & (!sk[92]) & (g165) & (g495) & (g825) & (!g829)) + ((!g125) & (!sk[92]) & (g165) & (g495) & (g825) & (g829)) + ((!g125) & (sk[92]) & (!g165) & (!g495) & (!g825) & (g829)) + ((!g125) & (sk[92]) & (!g165) & (g495) & (!g825) & (g829)) + ((!g125) & (sk[92]) & (g165) & (!g495) & (!g825) & (g829)) + ((g125) & (!sk[92]) & (!g165) & (g495) & (!g825) & (g829)) + ((g125) & (!sk[92]) & (!g165) & (g495) & (g825) & (!g829)) + ((g125) & (!sk[92]) & (!g165) & (g495) & (g825) & (g829)) + ((g125) & (!sk[92]) & (g165) & (!g495) & (!g825) & (!g829)) + ((g125) & (!sk[92]) & (g165) & (!g495) & (!g825) & (g829)) + ((g125) & (!sk[92]) & (g165) & (!g495) & (g825) & (!g829)) + ((g125) & (!sk[92]) & (g165) & (!g495) & (g825) & (g829)) + ((g125) & (!sk[92]) & (g165) & (g495) & (!g825) & (!g829)) + ((g125) & (!sk[92]) & (g165) & (g495) & (!g825) & (g829)) + ((g125) & (!sk[92]) & (g165) & (g495) & (g825) & (!g829)) + ((g125) & (!sk[92]) & (g165) & (g495) & (g825) & (g829)) + ((g125) & (sk[92]) & (!g165) & (!g495) & (!g825) & (g829)) + ((g125) & (sk[92]) & (g165) & (!g495) & (!g825) & (g829)));
	assign g831 = (((!g161) & (!g90) & (!g413) & (!g217) & (!g501) & (!g736)) + ((!g161) & (!g90) & (!g413) & (!g217) & (g501) & (!g736)) + ((!g161) & (!g90) & (!g413) & (g217) & (!g501) & (!g736)) + ((!g161) & (!g90) & (!g413) & (g217) & (g501) & (!g736)) + ((!g161) & (!g90) & (g413) & (!g217) & (!g501) & (!g736)) + ((!g161) & (!g90) & (g413) & (!g217) & (!g501) & (g736)) + ((!g161) & (!g90) & (g413) & (!g217) & (g501) & (!g736)) + ((!g161) & (!g90) & (g413) & (!g217) & (g501) & (g736)) + ((!g161) & (!g90) & (g413) & (g217) & (!g501) & (!g736)) + ((!g161) & (!g90) & (g413) & (g217) & (g501) & (!g736)) + ((!g161) & (g90) & (!g413) & (!g217) & (!g501) & (!g736)) + ((!g161) & (g90) & (!g413) & (!g217) & (g501) & (!g736)) + ((!g161) & (g90) & (!g413) & (g217) & (!g501) & (!g736)) + ((!g161) & (g90) & (!g413) & (g217) & (g501) & (!g736)) + ((!g161) & (g90) & (g413) & (!g217) & (!g501) & (!g736)) + ((!g161) & (g90) & (g413) & (!g217) & (!g501) & (g736)) + ((!g161) & (g90) & (g413) & (!g217) & (g501) & (!g736)) + ((!g161) & (g90) & (g413) & (!g217) & (g501) & (g736)) + ((!g161) & (g90) & (g413) & (g217) & (!g501) & (!g736)) + ((!g161) & (g90) & (g413) & (g217) & (g501) & (!g736)) + ((g161) & (!g90) & (!g413) & (!g217) & (!g501) & (!g736)) + ((g161) & (!g90) & (!g413) & (g217) & (!g501) & (!g736)) + ((g161) & (!g90) & (g413) & (!g217) & (!g501) & (!g736)) + ((g161) & (!g90) & (g413) & (!g217) & (!g501) & (g736)) + ((g161) & (!g90) & (g413) & (g217) & (!g501) & (!g736)));
	assign g832 = (((!g78) & (!g356) & (!g392) & (!g486) & (!g534) & (g831)) + ((!g78) & (!g356) & (!g392) & (!g486) & (g534) & (g831)) + ((!g78) & (!g356) & (!g392) & (g486) & (!g534) & (g831)) + ((!g78) & (!g356) & (!g392) & (g486) & (g534) & (g831)) + ((!g78) & (g356) & (!g392) & (!g486) & (!g534) & (g831)) + ((g78) & (!g356) & (!g392) & (!g486) & (!g534) & (g831)) + ((g78) & (!g356) & (!g392) & (!g486) & (g534) & (g831)) + ((g78) & (!g356) & (!g392) & (g486) & (!g534) & (g831)) + ((g78) & (!g356) & (!g392) & (g486) & (g534) & (g831)) + ((g78) & (!g356) & (g392) & (!g486) & (!g534) & (g831)) + ((g78) & (!g356) & (g392) & (!g486) & (g534) & (g831)) + ((g78) & (!g356) & (g392) & (g486) & (!g534) & (g831)) + ((g78) & (!g356) & (g392) & (g486) & (g534) & (g831)) + ((g78) & (g356) & (!g392) & (!g486) & (!g534) & (g831)) + ((g78) & (g356) & (g392) & (!g486) & (!g534) & (g831)));
	assign g833 = (((!g127) & (!g402) & (!g443) & (sk[95]) & (!g642) & (g655)) + ((!g127) & (!g402) & (g443) & (!sk[95]) & (!g642) & (g655)) + ((!g127) & (!g402) & (g443) & (!sk[95]) & (g642) & (!g655)) + ((!g127) & (!g402) & (g443) & (!sk[95]) & (g642) & (g655)) + ((!g127) & (!g402) & (g443) & (sk[95]) & (!g642) & (g655)) + ((!g127) & (!g402) & (g443) & (sk[95]) & (g642) & (g655)) + ((!g127) & (g402) & (!g443) & (!sk[95]) & (!g642) & (!g655)) + ((!g127) & (g402) & (!g443) & (!sk[95]) & (!g642) & (g655)) + ((!g127) & (g402) & (!g443) & (!sk[95]) & (g642) & (!g655)) + ((!g127) & (g402) & (!g443) & (!sk[95]) & (g642) & (g655)) + ((!g127) & (g402) & (!g443) & (sk[95]) & (!g642) & (!g655)) + ((!g127) & (g402) & (!g443) & (sk[95]) & (!g642) & (g655)) + ((!g127) & (g402) & (g443) & (!sk[95]) & (!g642) & (!g655)) + ((!g127) & (g402) & (g443) & (!sk[95]) & (!g642) & (g655)) + ((!g127) & (g402) & (g443) & (!sk[95]) & (g642) & (!g655)) + ((!g127) & (g402) & (g443) & (!sk[95]) & (g642) & (g655)) + ((!g127) & (g402) & (g443) & (sk[95]) & (!g642) & (!g655)) + ((!g127) & (g402) & (g443) & (sk[95]) & (!g642) & (g655)) + ((!g127) & (g402) & (g443) & (sk[95]) & (g642) & (!g655)) + ((!g127) & (g402) & (g443) & (sk[95]) & (g642) & (g655)) + ((g127) & (!g402) & (g443) & (!sk[95]) & (!g642) & (g655)) + ((g127) & (!g402) & (g443) & (!sk[95]) & (g642) & (!g655)) + ((g127) & (!g402) & (g443) & (!sk[95]) & (g642) & (g655)) + ((g127) & (g402) & (!g443) & (!sk[95]) & (!g642) & (!g655)) + ((g127) & (g402) & (!g443) & (!sk[95]) & (!g642) & (g655)) + ((g127) & (g402) & (!g443) & (!sk[95]) & (g642) & (!g655)) + ((g127) & (g402) & (!g443) & (!sk[95]) & (g642) & (g655)) + ((g127) & (g402) & (!g443) & (sk[95]) & (!g642) & (!g655)) + ((g127) & (g402) & (!g443) & (sk[95]) & (!g642) & (g655)) + ((g127) & (g402) & (g443) & (!sk[95]) & (!g642) & (!g655)) + ((g127) & (g402) & (g443) & (!sk[95]) & (!g642) & (g655)) + ((g127) & (g402) & (g443) & (!sk[95]) & (g642) & (!g655)) + ((g127) & (g402) & (g443) & (!sk[95]) & (g642) & (g655)) + ((g127) & (g402) & (g443) & (sk[95]) & (!g642) & (!g655)) + ((g127) & (g402) & (g443) & (sk[95]) & (!g642) & (g655)) + ((g127) & (g402) & (g443) & (sk[95]) & (g642) & (!g655)) + ((g127) & (g402) & (g443) & (sk[95]) & (g642) & (g655)));
	assign g834 = (((!g440) & (!g446) & (!sk[96]) & (g626) & (!g628)) + ((!g440) & (!g446) & (!sk[96]) & (g626) & (g628)) + ((!g440) & (!g446) & (sk[96]) & (!g626) & (!g628)) + ((!g440) & (!g446) & (sk[96]) & (g626) & (!g628)) + ((!g440) & (!g446) & (sk[96]) & (g626) & (g628)) + ((!g440) & (g446) & (!sk[96]) & (g626) & (!g628)) + ((!g440) & (g446) & (!sk[96]) & (g626) & (g628)) + ((!g440) & (g446) & (sk[96]) & (!g626) & (!g628)) + ((!g440) & (g446) & (sk[96]) & (g626) & (!g628)) + ((g440) & (!g446) & (!sk[96]) & (g626) & (!g628)) + ((g440) & (!g446) & (!sk[96]) & (g626) & (g628)) + ((g440) & (!g446) & (sk[96]) & (g626) & (!g628)) + ((g440) & (!g446) & (sk[96]) & (g626) & (g628)) + ((g440) & (g446) & (!sk[96]) & (g626) & (!g628)) + ((g440) & (g446) & (!sk[96]) & (g626) & (g628)));
	assign g835 = (((g61) & (!g824) & (g830) & (g832) & (g833) & (!g834)));
	assign g836 = (((!sk[98]) & (!g98) & (!g225) & (g213) & (!g425)) + ((!sk[98]) & (!g98) & (!g225) & (g213) & (g425)) + ((!sk[98]) & (!g98) & (g225) & (g213) & (!g425)) + ((!sk[98]) & (!g98) & (g225) & (g213) & (g425)) + ((!sk[98]) & (g98) & (!g225) & (g213) & (!g425)) + ((!sk[98]) & (g98) & (!g225) & (g213) & (g425)) + ((!sk[98]) & (g98) & (g225) & (g213) & (!g425)) + ((!sk[98]) & (g98) & (g225) & (g213) & (g425)) + ((sk[98]) & (g98) & (!g225) & (!g213) & (!g425)) + ((sk[98]) & (g98) & (!g225) & (g213) & (!g425)) + ((sk[98]) & (g98) & (!g225) & (g213) & (g425)) + ((sk[98]) & (g98) & (g225) & (!g213) & (!g425)) + ((sk[98]) & (g98) & (g225) & (!g213) & (g425)) + ((sk[98]) & (g98) & (g225) & (g213) & (!g425)) + ((sk[98]) & (g98) & (g225) & (g213) & (g425)));
	assign g837 = (((!g164) & (!sk[99]) & (!g79) & (g142) & (!g402) & (g392)) + ((!g164) & (!sk[99]) & (!g79) & (g142) & (g402) & (!g392)) + ((!g164) & (!sk[99]) & (!g79) & (g142) & (g402) & (g392)) + ((!g164) & (!sk[99]) & (g79) & (!g142) & (!g402) & (!g392)) + ((!g164) & (!sk[99]) & (g79) & (!g142) & (!g402) & (g392)) + ((!g164) & (!sk[99]) & (g79) & (!g142) & (g402) & (!g392)) + ((!g164) & (!sk[99]) & (g79) & (!g142) & (g402) & (g392)) + ((!g164) & (!sk[99]) & (g79) & (g142) & (!g402) & (!g392)) + ((!g164) & (!sk[99]) & (g79) & (g142) & (!g402) & (g392)) + ((!g164) & (!sk[99]) & (g79) & (g142) & (g402) & (!g392)) + ((!g164) & (!sk[99]) & (g79) & (g142) & (g402) & (g392)) + ((!g164) & (sk[99]) & (!g79) & (!g142) & (!g402) & (!g392)) + ((!g164) & (sk[99]) & (!g79) & (!g142) & (!g402) & (g392)) + ((!g164) & (sk[99]) & (!g79) & (!g142) & (g402) & (!g392)) + ((!g164) & (sk[99]) & (!g79) & (!g142) & (g402) & (g392)) + ((!g164) & (sk[99]) & (!g79) & (g142) & (!g402) & (!g392)) + ((!g164) & (sk[99]) & (!g79) & (g142) & (!g402) & (g392)) + ((!g164) & (sk[99]) & (!g79) & (g142) & (g402) & (g392)) + ((g164) & (!sk[99]) & (!g79) & (g142) & (!g402) & (g392)) + ((g164) & (!sk[99]) & (!g79) & (g142) & (g402) & (!g392)) + ((g164) & (!sk[99]) & (!g79) & (g142) & (g402) & (g392)) + ((g164) & (!sk[99]) & (g79) & (!g142) & (!g402) & (!g392)) + ((g164) & (!sk[99]) & (g79) & (!g142) & (!g402) & (g392)) + ((g164) & (!sk[99]) & (g79) & (!g142) & (g402) & (!g392)) + ((g164) & (!sk[99]) & (g79) & (!g142) & (g402) & (g392)) + ((g164) & (!sk[99]) & (g79) & (g142) & (!g402) & (!g392)) + ((g164) & (!sk[99]) & (g79) & (g142) & (!g402) & (g392)) + ((g164) & (!sk[99]) & (g79) & (g142) & (g402) & (!g392)) + ((g164) & (!sk[99]) & (g79) & (g142) & (g402) & (g392)) + ((g164) & (sk[99]) & (!g79) & (!g142) & (!g402) & (!g392)) + ((g164) & (sk[99]) & (!g79) & (!g142) & (!g402) & (g392)) + ((g164) & (sk[99]) & (!g79) & (!g142) & (g402) & (!g392)) + ((g164) & (sk[99]) & (!g79) & (!g142) & (g402) & (g392)) + ((g164) & (sk[99]) & (!g79) & (g142) & (!g402) & (!g392)) + ((g164) & (sk[99]) & (!g79) & (g142) & (!g402) & (g392)) + ((g164) & (sk[99]) & (!g79) & (g142) & (g402) & (!g392)) + ((g164) & (sk[99]) & (!g79) & (g142) & (g402) & (g392)));
	assign g838 = (((!g49) & (!g33) & (g166) & (!g401) & (!sk[100]) & (g534)) + ((!g49) & (!g33) & (g166) & (g401) & (!sk[100]) & (!g534)) + ((!g49) & (!g33) & (g166) & (g401) & (!sk[100]) & (g534)) + ((!g49) & (g33) & (!g166) & (!g401) & (!sk[100]) & (!g534)) + ((!g49) & (g33) & (!g166) & (!g401) & (!sk[100]) & (g534)) + ((!g49) & (g33) & (!g166) & (!g401) & (sk[100]) & (!g534)) + ((!g49) & (g33) & (!g166) & (!g401) & (sk[100]) & (g534)) + ((!g49) & (g33) & (!g166) & (g401) & (!sk[100]) & (!g534)) + ((!g49) & (g33) & (!g166) & (g401) & (!sk[100]) & (g534)) + ((!g49) & (g33) & (g166) & (!g401) & (!sk[100]) & (!g534)) + ((!g49) & (g33) & (g166) & (!g401) & (!sk[100]) & (g534)) + ((!g49) & (g33) & (g166) & (!g401) & (sk[100]) & (!g534)) + ((!g49) & (g33) & (g166) & (!g401) & (sk[100]) & (g534)) + ((!g49) & (g33) & (g166) & (g401) & (!sk[100]) & (!g534)) + ((!g49) & (g33) & (g166) & (g401) & (!sk[100]) & (g534)) + ((g49) & (!g33) & (g166) & (!g401) & (!sk[100]) & (g534)) + ((g49) & (!g33) & (g166) & (!g401) & (sk[100]) & (g534)) + ((g49) & (!g33) & (g166) & (g401) & (!sk[100]) & (!g534)) + ((g49) & (!g33) & (g166) & (g401) & (!sk[100]) & (g534)) + ((g49) & (!g33) & (g166) & (g401) & (sk[100]) & (g534)) + ((g49) & (g33) & (!g166) & (!g401) & (!sk[100]) & (!g534)) + ((g49) & (g33) & (!g166) & (!g401) & (!sk[100]) & (g534)) + ((g49) & (g33) & (!g166) & (!g401) & (sk[100]) & (!g534)) + ((g49) & (g33) & (!g166) & (!g401) & (sk[100]) & (g534)) + ((g49) & (g33) & (!g166) & (g401) & (!sk[100]) & (!g534)) + ((g49) & (g33) & (!g166) & (g401) & (!sk[100]) & (g534)) + ((g49) & (g33) & (g166) & (!g401) & (!sk[100]) & (!g534)) + ((g49) & (g33) & (g166) & (!g401) & (!sk[100]) & (g534)) + ((g49) & (g33) & (g166) & (!g401) & (sk[100]) & (!g534)) + ((g49) & (g33) & (g166) & (!g401) & (sk[100]) & (g534)) + ((g49) & (g33) & (g166) & (g401) & (!sk[100]) & (!g534)) + ((g49) & (g33) & (g166) & (g401) & (!sk[100]) & (g534)) + ((g49) & (g33) & (g166) & (g401) & (sk[100]) & (g534)));
	assign g839 = (((!g130) & (!g425) & (!g648) & (!g688) & (sk[101]) & (!g838)) + ((!g130) & (!g425) & (g648) & (!g688) & (!sk[101]) & (g838)) + ((!g130) & (!g425) & (g648) & (g688) & (!sk[101]) & (!g838)) + ((!g130) & (!g425) & (g648) & (g688) & (!sk[101]) & (g838)) + ((!g130) & (g425) & (!g648) & (!g688) & (!sk[101]) & (!g838)) + ((!g130) & (g425) & (!g648) & (!g688) & (!sk[101]) & (g838)) + ((!g130) & (g425) & (!g648) & (!g688) & (sk[101]) & (!g838)) + ((!g130) & (g425) & (!g648) & (g688) & (!sk[101]) & (!g838)) + ((!g130) & (g425) & (!g648) & (g688) & (!sk[101]) & (g838)) + ((!g130) & (g425) & (g648) & (!g688) & (!sk[101]) & (!g838)) + ((!g130) & (g425) & (g648) & (!g688) & (!sk[101]) & (g838)) + ((!g130) & (g425) & (g648) & (!g688) & (sk[101]) & (!g838)) + ((!g130) & (g425) & (g648) & (g688) & (!sk[101]) & (!g838)) + ((!g130) & (g425) & (g648) & (g688) & (!sk[101]) & (g838)) + ((g130) & (!g425) & (!g648) & (!g688) & (sk[101]) & (!g838)) + ((g130) & (!g425) & (!g648) & (g688) & (sk[101]) & (!g838)) + ((g130) & (!g425) & (g648) & (!g688) & (!sk[101]) & (g838)) + ((g130) & (!g425) & (g648) & (g688) & (!sk[101]) & (!g838)) + ((g130) & (!g425) & (g648) & (g688) & (!sk[101]) & (g838)) + ((g130) & (g425) & (!g648) & (!g688) & (!sk[101]) & (!g838)) + ((g130) & (g425) & (!g648) & (!g688) & (!sk[101]) & (g838)) + ((g130) & (g425) & (!g648) & (!g688) & (sk[101]) & (!g838)) + ((g130) & (g425) & (!g648) & (g688) & (!sk[101]) & (!g838)) + ((g130) & (g425) & (!g648) & (g688) & (!sk[101]) & (g838)) + ((g130) & (g425) & (!g648) & (g688) & (sk[101]) & (!g838)) + ((g130) & (g425) & (g648) & (!g688) & (!sk[101]) & (!g838)) + ((g130) & (g425) & (g648) & (!g688) & (!sk[101]) & (g838)) + ((g130) & (g425) & (g648) & (!g688) & (sk[101]) & (!g838)) + ((g130) & (g425) & (g648) & (g688) & (!sk[101]) & (!g838)) + ((g130) & (g425) & (g648) & (g688) & (!sk[101]) & (g838)) + ((g130) & (g425) & (g648) & (g688) & (sk[101]) & (!g838)));
	assign g840 = (((!g22) & (!g76) & (!g83) & (sk[102]) & (!g435) & (!g444)) + ((!g22) & (!g76) & (!g83) & (sk[102]) & (g435) & (!g444)) + ((!g22) & (!g76) & (g83) & (!sk[102]) & (!g435) & (g444)) + ((!g22) & (!g76) & (g83) & (!sk[102]) & (g435) & (!g444)) + ((!g22) & (!g76) & (g83) & (!sk[102]) & (g435) & (g444)) + ((!g22) & (!g76) & (g83) & (sk[102]) & (!g435) & (!g444)) + ((!g22) & (!g76) & (g83) & (sk[102]) & (!g435) & (g444)) + ((!g22) & (!g76) & (g83) & (sk[102]) & (g435) & (!g444)) + ((!g22) & (g76) & (!g83) & (!sk[102]) & (!g435) & (!g444)) + ((!g22) & (g76) & (!g83) & (!sk[102]) & (!g435) & (g444)) + ((!g22) & (g76) & (!g83) & (!sk[102]) & (g435) & (!g444)) + ((!g22) & (g76) & (!g83) & (!sk[102]) & (g435) & (g444)) + ((!g22) & (g76) & (g83) & (!sk[102]) & (!g435) & (!g444)) + ((!g22) & (g76) & (g83) & (!sk[102]) & (!g435) & (g444)) + ((!g22) & (g76) & (g83) & (!sk[102]) & (g435) & (!g444)) + ((!g22) & (g76) & (g83) & (!sk[102]) & (g435) & (g444)) + ((g22) & (!g76) & (g83) & (!sk[102]) & (!g435) & (g444)) + ((g22) & (!g76) & (g83) & (!sk[102]) & (g435) & (!g444)) + ((g22) & (!g76) & (g83) & (!sk[102]) & (g435) & (g444)) + ((g22) & (!g76) & (g83) & (sk[102]) & (!g435) & (!g444)) + ((g22) & (!g76) & (g83) & (sk[102]) & (!g435) & (g444)) + ((g22) & (g76) & (!g83) & (!sk[102]) & (!g435) & (!g444)) + ((g22) & (g76) & (!g83) & (!sk[102]) & (!g435) & (g444)) + ((g22) & (g76) & (!g83) & (!sk[102]) & (g435) & (!g444)) + ((g22) & (g76) & (!g83) & (!sk[102]) & (g435) & (g444)) + ((g22) & (g76) & (g83) & (!sk[102]) & (!g435) & (!g444)) + ((g22) & (g76) & (g83) & (!sk[102]) & (!g435) & (g444)) + ((g22) & (g76) & (g83) & (!sk[102]) & (g435) & (!g444)) + ((g22) & (g76) & (g83) & (!sk[102]) & (g435) & (g444)));
	assign g841 = (((!i_8_) & (i_6_) & (!i_7_) & (!g21) & (!g23) & (g118)) + ((!i_8_) & (i_6_) & (!i_7_) & (g21) & (!g23) & (g118)) + ((i_8_) & (!i_6_) & (!i_7_) & (g21) & (!g23) & (g118)) + ((i_8_) & (!i_6_) & (!i_7_) & (g21) & (g23) & (g118)));
	assign g842 = (((!g17) & (!sk[104]) & (!g19) & (g434) & (!g841)) + ((!g17) & (!sk[104]) & (!g19) & (g434) & (g841)) + ((!g17) & (!sk[104]) & (g19) & (g434) & (!g841)) + ((!g17) & (!sk[104]) & (g19) & (g434) & (g841)) + ((!g17) & (sk[104]) & (!g19) & (!g434) & (!g841)) + ((!g17) & (sk[104]) & (!g19) & (g434) & (!g841)) + ((!g17) & (sk[104]) & (g19) & (!g434) & (!g841)) + ((!g17) & (sk[104]) & (g19) & (g434) & (!g841)) + ((g17) & (!sk[104]) & (!g19) & (g434) & (!g841)) + ((g17) & (!sk[104]) & (!g19) & (g434) & (g841)) + ((g17) & (!sk[104]) & (g19) & (g434) & (!g841)) + ((g17) & (!sk[104]) & (g19) & (g434) & (g841)) + ((g17) & (sk[104]) & (!g19) & (!g434) & (!g841)) + ((g17) & (sk[104]) & (!g19) & (g434) & (!g841)) + ((g17) & (sk[104]) & (g19) & (!g434) & (!g841)));
	assign g843 = (((!g109) & (!g157) & (!g422) & (sk[105]) & (g842)) + ((!g109) & (!g157) & (g422) & (!sk[105]) & (!g842)) + ((!g109) & (!g157) & (g422) & (!sk[105]) & (g842)) + ((!g109) & (!g157) & (g422) & (sk[105]) & (g842)) + ((!g109) & (g157) & (!g422) & (sk[105]) & (g842)) + ((!g109) & (g157) & (g422) & (!sk[105]) & (!g842)) + ((!g109) & (g157) & (g422) & (!sk[105]) & (g842)) + ((!g109) & (g157) & (g422) & (sk[105]) & (g842)) + ((g109) & (!g157) & (!g422) & (sk[105]) & (g842)) + ((g109) & (!g157) & (g422) & (!sk[105]) & (!g842)) + ((g109) & (!g157) & (g422) & (!sk[105]) & (g842)) + ((g109) & (g157) & (g422) & (!sk[105]) & (!g842)) + ((g109) & (g157) & (g422) & (!sk[105]) & (g842)));
	assign g844 = (((!g836) & (!g837) & (g1511) & (g839) & (!g840) & (g843)));
	assign g845 = (((g173) & (g813) & (g697) & (g823) & (g835) & (g844)));
	assign g846 = (((!i_0_) & (!sk[108]) & (!i_1_) & (g15) & (!g32) & (g39)) + ((!i_0_) & (!sk[108]) & (!i_1_) & (g15) & (g32) & (!g39)) + ((!i_0_) & (!sk[108]) & (!i_1_) & (g15) & (g32) & (g39)) + ((!i_0_) & (!sk[108]) & (i_1_) & (!g15) & (!g32) & (!g39)) + ((!i_0_) & (!sk[108]) & (i_1_) & (!g15) & (!g32) & (g39)) + ((!i_0_) & (!sk[108]) & (i_1_) & (!g15) & (g32) & (!g39)) + ((!i_0_) & (!sk[108]) & (i_1_) & (!g15) & (g32) & (g39)) + ((!i_0_) & (!sk[108]) & (i_1_) & (g15) & (!g32) & (!g39)) + ((!i_0_) & (!sk[108]) & (i_1_) & (g15) & (!g32) & (g39)) + ((!i_0_) & (!sk[108]) & (i_1_) & (g15) & (g32) & (!g39)) + ((!i_0_) & (!sk[108]) & (i_1_) & (g15) & (g32) & (g39)) + ((!i_0_) & (sk[108]) & (!i_1_) & (!g15) & (!g32) & (!g39)) + ((!i_0_) & (sk[108]) & (!i_1_) & (g15) & (!g32) & (!g39)) + ((!i_0_) & (sk[108]) & (i_1_) & (!g15) & (!g32) & (!g39)) + ((!i_0_) & (sk[108]) & (i_1_) & (g15) & (!g32) & (!g39)) + ((i_0_) & (!sk[108]) & (!i_1_) & (g15) & (!g32) & (g39)) + ((i_0_) & (!sk[108]) & (!i_1_) & (g15) & (g32) & (!g39)) + ((i_0_) & (!sk[108]) & (!i_1_) & (g15) & (g32) & (g39)) + ((i_0_) & (!sk[108]) & (i_1_) & (!g15) & (!g32) & (!g39)) + ((i_0_) & (!sk[108]) & (i_1_) & (!g15) & (!g32) & (g39)) + ((i_0_) & (!sk[108]) & (i_1_) & (!g15) & (g32) & (!g39)) + ((i_0_) & (!sk[108]) & (i_1_) & (!g15) & (g32) & (g39)) + ((i_0_) & (!sk[108]) & (i_1_) & (g15) & (!g32) & (!g39)) + ((i_0_) & (!sk[108]) & (i_1_) & (g15) & (!g32) & (g39)) + ((i_0_) & (!sk[108]) & (i_1_) & (g15) & (g32) & (!g39)) + ((i_0_) & (!sk[108]) & (i_1_) & (g15) & (g32) & (g39)) + ((i_0_) & (sk[108]) & (!i_1_) & (!g15) & (!g32) & (!g39)) + ((i_0_) & (sk[108]) & (i_1_) & (!g15) & (!g32) & (!g39)) + ((i_0_) & (sk[108]) & (i_1_) & (g15) & (!g32) & (!g39)));
	assign g847 = (((!sk[109]) & (g4) & (!g86)) + ((!sk[109]) & (g4) & (g86)) + ((sk[109]) & (!g4) & (!g86)) + ((sk[109]) & (!g4) & (g86)) + ((sk[109]) & (g4) & (!g86)));
	assign g848 = (((!i_12_) & (!sk[110]) & (!i_13_) & (i_14_) & (!g86)) + ((!i_12_) & (!sk[110]) & (!i_13_) & (i_14_) & (g86)) + ((!i_12_) & (!sk[110]) & (i_13_) & (i_14_) & (!g86)) + ((!i_12_) & (!sk[110]) & (i_13_) & (i_14_) & (g86)) + ((!i_12_) & (sk[110]) & (!i_13_) & (!i_14_) & (!g86)) + ((!i_12_) & (sk[110]) & (!i_13_) & (!i_14_) & (g86)) + ((!i_12_) & (sk[110]) & (!i_13_) & (i_14_) & (!g86)) + ((!i_12_) & (sk[110]) & (!i_13_) & (i_14_) & (g86)) + ((!i_12_) & (sk[110]) & (i_13_) & (!i_14_) & (!g86)) + ((!i_12_) & (sk[110]) & (i_13_) & (i_14_) & (!g86)) + ((!i_12_) & (sk[110]) & (i_13_) & (i_14_) & (g86)) + ((i_12_) & (!sk[110]) & (!i_13_) & (i_14_) & (!g86)) + ((i_12_) & (!sk[110]) & (!i_13_) & (i_14_) & (g86)) + ((i_12_) & (!sk[110]) & (i_13_) & (i_14_) & (!g86)) + ((i_12_) & (!sk[110]) & (i_13_) & (i_14_) & (g86)) + ((i_12_) & (sk[110]) & (!i_13_) & (!i_14_) & (!g86)) + ((i_12_) & (sk[110]) & (!i_13_) & (i_14_) & (!g86)) + ((i_12_) & (sk[110]) & (!i_13_) & (i_14_) & (g86)) + ((i_12_) & (sk[110]) & (i_13_) & (!i_14_) & (!g86)) + ((i_12_) & (sk[110]) & (i_13_) & (i_14_) & (!g86)) + ((i_12_) & (sk[110]) & (i_13_) & (i_14_) & (g86)));
	assign g849 = (((!i_12_) & (!i_13_) & (i_14_) & (!sk[111]) & (!g35)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[111]) & (g35)) + ((!i_12_) & (i_13_) & (!i_14_) & (sk[111]) & (g35)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[111]) & (!g35)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[111]) & (g35)) + ((i_12_) & (!i_13_) & (!i_14_) & (sk[111]) & (g35)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[111]) & (!g35)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[111]) & (g35)) + ((i_12_) & (i_13_) & (!i_14_) & (sk[111]) & (g35)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[111]) & (!g35)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[111]) & (g35)));
	assign g850 = (((!i_12_) & (!i_13_) & (i_14_) & (!sk[112]) & (!g83)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[112]) & (g83)) + ((!i_12_) & (i_13_) & (!i_14_) & (sk[112]) & (g83)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[112]) & (!g83)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[112]) & (g83)) + ((i_12_) & (!i_13_) & (!i_14_) & (sk[112]) & (g83)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[112]) & (!g83)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[112]) & (g83)) + ((i_12_) & (i_13_) & (!i_14_) & (sk[112]) & (g83)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[112]) & (!g83)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[112]) & (g83)));
	assign g851 = (((!g4) & (sk[113]) & (!g35)) + ((!g4) & (sk[113]) & (g35)) + ((g4) & (!sk[113]) & (!g35)) + ((g4) & (!sk[113]) & (g35)) + ((g4) & (sk[113]) & (!g35)));
	assign g852 = (((g4) & (!sk[114]) & (!g107)) + ((g4) & (!sk[114]) & (g107)) + ((g4) & (sk[114]) & (!g107)));
	assign g853 = (((!i_12_) & (!i_13_) & (i_14_) & (!sk[115]) & (!g107)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[115]) & (g107)) + ((!i_12_) & (i_13_) & (!i_14_) & (sk[115]) & (!g107)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[115]) & (!g107)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[115]) & (g107)) + ((i_12_) & (!i_13_) & (!i_14_) & (sk[115]) & (!g107)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[115]) & (!g107)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[115]) & (g107)) + ((i_12_) & (i_13_) & (!i_14_) & (sk[115]) & (!g107)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[115]) & (!g107)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[115]) & (g107)));
	assign g854 = (((!g253) & (!g849) & (!g852) & (sk[116]) & (!g848) & (!g853)) + ((!g253) & (!g849) & (!g852) & (sk[116]) & (!g848) & (g853)) + ((!g253) & (!g849) & (!g852) & (sk[116]) & (g848) & (g853)) + ((!g253) & (!g849) & (g852) & (!sk[116]) & (!g848) & (g853)) + ((!g253) & (!g849) & (g852) & (!sk[116]) & (g848) & (!g853)) + ((!g253) & (!g849) & (g852) & (!sk[116]) & (g848) & (g853)) + ((!g253) & (!g849) & (g852) & (sk[116]) & (!g848) & (!g853)) + ((!g253) & (!g849) & (g852) & (sk[116]) & (!g848) & (g853)) + ((!g253) & (!g849) & (g852) & (sk[116]) & (g848) & (!g853)) + ((!g253) & (!g849) & (g852) & (sk[116]) & (g848) & (g853)) + ((!g253) & (g849) & (!g852) & (!sk[116]) & (!g848) & (!g853)) + ((!g253) & (g849) & (!g852) & (!sk[116]) & (!g848) & (g853)) + ((!g253) & (g849) & (!g852) & (!sk[116]) & (g848) & (!g853)) + ((!g253) & (g849) & (!g852) & (!sk[116]) & (g848) & (g853)) + ((!g253) & (g849) & (!g852) & (sk[116]) & (!g848) & (!g853)) + ((!g253) & (g849) & (!g852) & (sk[116]) & (!g848) & (g853)) + ((!g253) & (g849) & (!g852) & (sk[116]) & (g848) & (!g853)) + ((!g253) & (g849) & (!g852) & (sk[116]) & (g848) & (g853)) + ((!g253) & (g849) & (g852) & (!sk[116]) & (!g848) & (!g853)) + ((!g253) & (g849) & (g852) & (!sk[116]) & (!g848) & (g853)) + ((!g253) & (g849) & (g852) & (!sk[116]) & (g848) & (!g853)) + ((!g253) & (g849) & (g852) & (!sk[116]) & (g848) & (g853)) + ((!g253) & (g849) & (g852) & (sk[116]) & (!g848) & (!g853)) + ((!g253) & (g849) & (g852) & (sk[116]) & (!g848) & (g853)) + ((!g253) & (g849) & (g852) & (sk[116]) & (g848) & (!g853)) + ((!g253) & (g849) & (g852) & (sk[116]) & (g848) & (g853)) + ((g253) & (!g849) & (g852) & (!sk[116]) & (!g848) & (g853)) + ((g253) & (!g849) & (g852) & (!sk[116]) & (g848) & (!g853)) + ((g253) & (!g849) & (g852) & (!sk[116]) & (g848) & (g853)) + ((g253) & (g849) & (!g852) & (!sk[116]) & (!g848) & (!g853)) + ((g253) & (g849) & (!g852) & (!sk[116]) & (!g848) & (g853)) + ((g253) & (g849) & (!g852) & (!sk[116]) & (g848) & (!g853)) + ((g253) & (g849) & (!g852) & (!sk[116]) & (g848) & (g853)) + ((g253) & (g849) & (g852) & (!sk[116]) & (!g848) & (!g853)) + ((g253) & (g849) & (g852) & (!sk[116]) & (!g848) & (g853)) + ((g253) & (g849) & (g852) & (!sk[116]) & (g848) & (!g853)) + ((g253) & (g849) & (g852) & (!sk[116]) & (g848) & (g853)));
	assign g855 = (((!g164) & (!g849) & (!g847) & (!g850) & (!g851) & (!g854)) + ((!g164) & (!g849) & (!g847) & (!g850) & (g851) & (!g854)) + ((!g164) & (!g849) & (!g847) & (g850) & (!g851) & (!g854)) + ((!g164) & (!g849) & (!g847) & (g850) & (g851) & (!g854)) + ((!g164) & (!g849) & (g847) & (!g850) & (!g851) & (!g854)) + ((!g164) & (!g849) & (g847) & (!g850) & (g851) & (!g854)) + ((!g164) & (!g849) & (g847) & (g850) & (!g851) & (!g854)) + ((!g164) & (!g849) & (g847) & (g850) & (g851) & (!g854)) + ((!g164) & (g849) & (!g847) & (!g850) & (!g851) & (!g854)) + ((!g164) & (g849) & (!g847) & (!g850) & (g851) & (!g854)) + ((!g164) & (g849) & (!g847) & (g850) & (!g851) & (!g854)) + ((!g164) & (g849) & (!g847) & (g850) & (g851) & (!g854)) + ((!g164) & (g849) & (g847) & (!g850) & (!g851) & (!g854)) + ((!g164) & (g849) & (g847) & (!g850) & (g851) & (!g854)) + ((!g164) & (g849) & (g847) & (g850) & (!g851) & (!g854)) + ((!g164) & (g849) & (g847) & (g850) & (g851) & (!g854)) + ((g164) & (!g849) & (g847) & (!g850) & (g851) & (!g854)));
	assign g856 = (((!g125) & (!sk[118]) & (!g164) & (g847) & (!g848) & (g855)) + ((!g125) & (!sk[118]) & (!g164) & (g847) & (g848) & (!g855)) + ((!g125) & (!sk[118]) & (!g164) & (g847) & (g848) & (g855)) + ((!g125) & (!sk[118]) & (g164) & (!g847) & (!g848) & (!g855)) + ((!g125) & (!sk[118]) & (g164) & (!g847) & (!g848) & (g855)) + ((!g125) & (!sk[118]) & (g164) & (!g847) & (g848) & (!g855)) + ((!g125) & (!sk[118]) & (g164) & (!g847) & (g848) & (g855)) + ((!g125) & (!sk[118]) & (g164) & (g847) & (!g848) & (!g855)) + ((!g125) & (!sk[118]) & (g164) & (g847) & (!g848) & (g855)) + ((!g125) & (!sk[118]) & (g164) & (g847) & (g848) & (!g855)) + ((!g125) & (!sk[118]) & (g164) & (g847) & (g848) & (g855)) + ((!g125) & (sk[118]) & (!g164) & (!g847) & (!g848) & (g855)) + ((!g125) & (sk[118]) & (!g164) & (!g847) & (g848) & (g855)) + ((!g125) & (sk[118]) & (!g164) & (g847) & (!g848) & (g855)) + ((!g125) & (sk[118]) & (!g164) & (g847) & (g848) & (g855)) + ((!g125) & (sk[118]) & (g164) & (!g847) & (g848) & (g855)) + ((!g125) & (sk[118]) & (g164) & (g847) & (g848) & (g855)) + ((g125) & (!sk[118]) & (!g164) & (g847) & (!g848) & (g855)) + ((g125) & (!sk[118]) & (!g164) & (g847) & (g848) & (!g855)) + ((g125) & (!sk[118]) & (!g164) & (g847) & (g848) & (g855)) + ((g125) & (!sk[118]) & (g164) & (!g847) & (!g848) & (!g855)) + ((g125) & (!sk[118]) & (g164) & (!g847) & (!g848) & (g855)) + ((g125) & (!sk[118]) & (g164) & (!g847) & (g848) & (!g855)) + ((g125) & (!sk[118]) & (g164) & (!g847) & (g848) & (g855)) + ((g125) & (!sk[118]) & (g164) & (g847) & (!g848) & (!g855)) + ((g125) & (!sk[118]) & (g164) & (g847) & (!g848) & (g855)) + ((g125) & (!sk[118]) & (g164) & (g847) & (g848) & (!g855)) + ((g125) & (!sk[118]) & (g164) & (g847) & (g848) & (g855)) + ((g125) & (sk[118]) & (!g164) & (g847) & (!g848) & (g855)) + ((g125) & (sk[118]) & (!g164) & (g847) & (g848) & (g855)) + ((g125) & (sk[118]) & (g164) & (g847) & (g848) & (g855)));
	assign g857 = (((!sk[119]) & (g4) & (!g126)) + ((!sk[119]) & (g4) & (g126)) + ((sk[119]) & (g4) & (!g126)));
	assign g858 = (((!i_8_) & (!g73) & (!sk[120]) & (g102) & (!g851) & (g857)) + ((!i_8_) & (!g73) & (!sk[120]) & (g102) & (g851) & (!g857)) + ((!i_8_) & (!g73) & (!sk[120]) & (g102) & (g851) & (g857)) + ((!i_8_) & (!g73) & (sk[120]) & (g102) & (!g851) & (!g857)) + ((!i_8_) & (!g73) & (sk[120]) & (g102) & (!g851) & (g857)) + ((!i_8_) & (g73) & (!sk[120]) & (!g102) & (!g851) & (!g857)) + ((!i_8_) & (g73) & (!sk[120]) & (!g102) & (!g851) & (g857)) + ((!i_8_) & (g73) & (!sk[120]) & (!g102) & (g851) & (!g857)) + ((!i_8_) & (g73) & (!sk[120]) & (!g102) & (g851) & (g857)) + ((!i_8_) & (g73) & (!sk[120]) & (g102) & (!g851) & (!g857)) + ((!i_8_) & (g73) & (!sk[120]) & (g102) & (!g851) & (g857)) + ((!i_8_) & (g73) & (!sk[120]) & (g102) & (g851) & (!g857)) + ((!i_8_) & (g73) & (!sk[120]) & (g102) & (g851) & (g857)) + ((!i_8_) & (g73) & (sk[120]) & (!g102) & (!g851) & (!g857)) + ((!i_8_) & (g73) & (sk[120]) & (!g102) & (!g851) & (g857)) + ((!i_8_) & (g73) & (sk[120]) & (!g102) & (g851) & (g857)) + ((!i_8_) & (g73) & (sk[120]) & (g102) & (!g851) & (!g857)) + ((!i_8_) & (g73) & (sk[120]) & (g102) & (!g851) & (g857)) + ((!i_8_) & (g73) & (sk[120]) & (g102) & (g851) & (g857)) + ((i_8_) & (!g73) & (!sk[120]) & (g102) & (!g851) & (g857)) + ((i_8_) & (!g73) & (!sk[120]) & (g102) & (g851) & (!g857)) + ((i_8_) & (!g73) & (!sk[120]) & (g102) & (g851) & (g857)) + ((i_8_) & (!g73) & (sk[120]) & (g102) & (!g851) & (!g857)) + ((i_8_) & (!g73) & (sk[120]) & (g102) & (!g851) & (g857)) + ((i_8_) & (g73) & (!sk[120]) & (!g102) & (!g851) & (!g857)) + ((i_8_) & (g73) & (!sk[120]) & (!g102) & (!g851) & (g857)) + ((i_8_) & (g73) & (!sk[120]) & (!g102) & (g851) & (!g857)) + ((i_8_) & (g73) & (!sk[120]) & (!g102) & (g851) & (g857)) + ((i_8_) & (g73) & (!sk[120]) & (g102) & (!g851) & (!g857)) + ((i_8_) & (g73) & (!sk[120]) & (g102) & (!g851) & (g857)) + ((i_8_) & (g73) & (!sk[120]) & (g102) & (g851) & (!g857)) + ((i_8_) & (g73) & (!sk[120]) & (g102) & (g851) & (g857)) + ((i_8_) & (g73) & (sk[120]) & (!g102) & (!g851) & (g857)) + ((i_8_) & (g73) & (sk[120]) & (!g102) & (g851) & (g857)) + ((i_8_) & (g73) & (sk[120]) & (g102) & (!g851) & (!g857)) + ((i_8_) & (g73) & (sk[120]) & (g102) & (!g851) & (g857)) + ((i_8_) & (g73) & (sk[120]) & (g102) & (g851) & (g857)));
	assign g859 = (((!g21) & (!sk[121]) & (!g73) & (g413) & (!g847) & (g858)) + ((!g21) & (!sk[121]) & (!g73) & (g413) & (g847) & (!g858)) + ((!g21) & (!sk[121]) & (!g73) & (g413) & (g847) & (g858)) + ((!g21) & (!sk[121]) & (g73) & (!g413) & (!g847) & (!g858)) + ((!g21) & (!sk[121]) & (g73) & (!g413) & (!g847) & (g858)) + ((!g21) & (!sk[121]) & (g73) & (!g413) & (g847) & (!g858)) + ((!g21) & (!sk[121]) & (g73) & (!g413) & (g847) & (g858)) + ((!g21) & (!sk[121]) & (g73) & (g413) & (!g847) & (!g858)) + ((!g21) & (!sk[121]) & (g73) & (g413) & (!g847) & (g858)) + ((!g21) & (!sk[121]) & (g73) & (g413) & (g847) & (!g858)) + ((!g21) & (!sk[121]) & (g73) & (g413) & (g847) & (g858)) + ((!g21) & (sk[121]) & (!g73) & (!g413) & (g847) & (!g858)) + ((!g21) & (sk[121]) & (!g73) & (g413) & (!g847) & (!g858)) + ((!g21) & (sk[121]) & (!g73) & (g413) & (g847) & (!g858)) + ((!g21) & (sk[121]) & (g73) & (!g413) & (g847) & (!g858)) + ((!g21) & (sk[121]) & (g73) & (g413) & (g847) & (!g858)) + ((g21) & (!sk[121]) & (!g73) & (g413) & (!g847) & (g858)) + ((g21) & (!sk[121]) & (!g73) & (g413) & (g847) & (!g858)) + ((g21) & (!sk[121]) & (!g73) & (g413) & (g847) & (g858)) + ((g21) & (!sk[121]) & (g73) & (!g413) & (!g847) & (!g858)) + ((g21) & (!sk[121]) & (g73) & (!g413) & (!g847) & (g858)) + ((g21) & (!sk[121]) & (g73) & (!g413) & (g847) & (!g858)) + ((g21) & (!sk[121]) & (g73) & (!g413) & (g847) & (g858)) + ((g21) & (!sk[121]) & (g73) & (g413) & (!g847) & (!g858)) + ((g21) & (!sk[121]) & (g73) & (g413) & (!g847) & (g858)) + ((g21) & (!sk[121]) & (g73) & (g413) & (g847) & (!g858)) + ((g21) & (!sk[121]) & (g73) & (g413) & (g847) & (g858)) + ((g21) & (sk[121]) & (!g73) & (g413) & (!g847) & (!g858)) + ((g21) & (sk[121]) & (!g73) & (g413) & (g847) & (!g858)) + ((g21) & (sk[121]) & (g73) & (g413) & (g847) & (!g858)));
	assign g860 = (((!i_9_) & (!i_10_) & (i_11_) & (!sk[122]) & (!i_15_) & (g460)) + ((!i_9_) & (!i_10_) & (i_11_) & (!sk[122]) & (i_15_) & (!g460)) + ((!i_9_) & (!i_10_) & (i_11_) & (!sk[122]) & (i_15_) & (g460)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[122]) & (!i_15_) & (!g460)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[122]) & (!i_15_) & (g460)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[122]) & (i_15_) & (!g460)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[122]) & (i_15_) & (g460)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[122]) & (!i_15_) & (!g460)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[122]) & (!i_15_) & (g460)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[122]) & (i_15_) & (!g460)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[122]) & (i_15_) & (g460)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[122]) & (!i_15_) & (g460)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[122]) & (i_15_) & (!g460)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[122]) & (i_15_) & (g460)) + ((i_9_) & (!i_10_) & (i_11_) & (sk[122]) & (!i_15_) & (!g460)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[122]) & (!i_15_) & (!g460)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[122]) & (!i_15_) & (g460)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[122]) & (i_15_) & (!g460)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[122]) & (i_15_) & (g460)) + ((i_9_) & (i_10_) & (!i_11_) & (sk[122]) & (!i_15_) & (!g460)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[122]) & (!i_15_) & (!g460)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[122]) & (!i_15_) & (g460)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[122]) & (i_15_) & (!g460)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[122]) & (i_15_) & (g460)));
	assign g861 = (((!i_9_) & (!sk[123]) & (!g101) & (g165) & (!g394) & (g860)) + ((!i_9_) & (!sk[123]) & (!g101) & (g165) & (g394) & (!g860)) + ((!i_9_) & (!sk[123]) & (!g101) & (g165) & (g394) & (g860)) + ((!i_9_) & (!sk[123]) & (g101) & (!g165) & (!g394) & (!g860)) + ((!i_9_) & (!sk[123]) & (g101) & (!g165) & (!g394) & (g860)) + ((!i_9_) & (!sk[123]) & (g101) & (!g165) & (g394) & (!g860)) + ((!i_9_) & (!sk[123]) & (g101) & (!g165) & (g394) & (g860)) + ((!i_9_) & (!sk[123]) & (g101) & (g165) & (!g394) & (!g860)) + ((!i_9_) & (!sk[123]) & (g101) & (g165) & (!g394) & (g860)) + ((!i_9_) & (!sk[123]) & (g101) & (g165) & (g394) & (!g860)) + ((!i_9_) & (!sk[123]) & (g101) & (g165) & (g394) & (g860)) + ((!i_9_) & (sk[123]) & (!g101) & (g165) & (!g394) & (g860)) + ((!i_9_) & (sk[123]) & (!g101) & (g165) & (g394) & (g860)) + ((!i_9_) & (sk[123]) & (g101) & (g165) & (!g394) & (g860)) + ((!i_9_) & (sk[123]) & (g101) & (g165) & (g394) & (g860)) + ((i_9_) & (!sk[123]) & (!g101) & (g165) & (!g394) & (g860)) + ((i_9_) & (!sk[123]) & (!g101) & (g165) & (g394) & (!g860)) + ((i_9_) & (!sk[123]) & (!g101) & (g165) & (g394) & (g860)) + ((i_9_) & (!sk[123]) & (g101) & (!g165) & (!g394) & (!g860)) + ((i_9_) & (!sk[123]) & (g101) & (!g165) & (!g394) & (g860)) + ((i_9_) & (!sk[123]) & (g101) & (!g165) & (g394) & (!g860)) + ((i_9_) & (!sk[123]) & (g101) & (!g165) & (g394) & (g860)) + ((i_9_) & (!sk[123]) & (g101) & (g165) & (!g394) & (!g860)) + ((i_9_) & (!sk[123]) & (g101) & (g165) & (!g394) & (g860)) + ((i_9_) & (!sk[123]) & (g101) & (g165) & (g394) & (!g860)) + ((i_9_) & (!sk[123]) & (g101) & (g165) & (g394) & (g860)) + ((i_9_) & (sk[123]) & (!g101) & (g165) & (!g394) & (g860)) + ((i_9_) & (sk[123]) & (!g101) & (g165) & (g394) & (g860)) + ((i_9_) & (sk[123]) & (g101) & (!g165) & (g394) & (!g860)) + ((i_9_) & (sk[123]) & (g101) & (!g165) & (g394) & (g860)) + ((i_9_) & (sk[123]) & (g101) & (g165) & (!g394) & (g860)) + ((i_9_) & (sk[123]) & (g101) & (g165) & (g394) & (!g860)) + ((i_9_) & (sk[123]) & (g101) & (g165) & (g394) & (g860)));
	assign g862 = (((!g122) & (!g847) & (!sk[124]) & (g851) & (!g861)) + ((!g122) & (!g847) & (!sk[124]) & (g851) & (g861)) + ((!g122) & (!g847) & (sk[124]) & (!g851) & (!g861)) + ((!g122) & (!g847) & (sk[124]) & (g851) & (!g861)) + ((!g122) & (g847) & (!sk[124]) & (g851) & (!g861)) + ((!g122) & (g847) & (!sk[124]) & (g851) & (g861)) + ((!g122) & (g847) & (sk[124]) & (!g851) & (!g861)) + ((!g122) & (g847) & (sk[124]) & (g851) & (!g861)) + ((g122) & (!g847) & (!sk[124]) & (g851) & (!g861)) + ((g122) & (!g847) & (!sk[124]) & (g851) & (g861)) + ((g122) & (g847) & (!sk[124]) & (g851) & (!g861)) + ((g122) & (g847) & (!sk[124]) & (g851) & (g861)) + ((g122) & (g847) & (sk[124]) & (g851) & (!g861)));
	assign g863 = (((!sk[125]) & (!g130) & (!g278) & (g421) & (!g392)) + ((!sk[125]) & (!g130) & (!g278) & (g421) & (g392)) + ((!sk[125]) & (!g130) & (g278) & (g421) & (!g392)) + ((!sk[125]) & (!g130) & (g278) & (g421) & (g392)) + ((!sk[125]) & (g130) & (!g278) & (g421) & (!g392)) + ((!sk[125]) & (g130) & (!g278) & (g421) & (g392)) + ((!sk[125]) & (g130) & (g278) & (g421) & (!g392)) + ((!sk[125]) & (g130) & (g278) & (g421) & (g392)) + ((sk[125]) & (!g130) & (g278) & (!g421) & (!g392)) + ((sk[125]) & (!g130) & (g278) & (!g421) & (g392)) + ((sk[125]) & (!g130) & (g278) & (g421) & (!g392)) + ((sk[125]) & (!g130) & (g278) & (g421) & (g392)) + ((sk[125]) & (g130) & (g278) & (!g421) & (g392)) + ((sk[125]) & (g130) & (g278) & (g421) & (!g392)) + ((sk[125]) & (g130) & (g278) & (g421) & (g392)));
	assign g864 = (((!g25) & (!g164) & (g402) & (!sk[126]) & (!g392) & (g863)) + ((!g25) & (!g164) & (g402) & (!sk[126]) & (g392) & (!g863)) + ((!g25) & (!g164) & (g402) & (!sk[126]) & (g392) & (g863)) + ((!g25) & (!g164) & (g402) & (sk[126]) & (!g392) & (!g863)) + ((!g25) & (g164) & (!g402) & (!sk[126]) & (!g392) & (!g863)) + ((!g25) & (g164) & (!g402) & (!sk[126]) & (!g392) & (g863)) + ((!g25) & (g164) & (!g402) & (!sk[126]) & (g392) & (!g863)) + ((!g25) & (g164) & (!g402) & (!sk[126]) & (g392) & (g863)) + ((!g25) & (g164) & (g402) & (!sk[126]) & (!g392) & (!g863)) + ((!g25) & (g164) & (g402) & (!sk[126]) & (!g392) & (g863)) + ((!g25) & (g164) & (g402) & (!sk[126]) & (g392) & (!g863)) + ((!g25) & (g164) & (g402) & (!sk[126]) & (g392) & (g863)) + ((g25) & (!g164) & (!g402) & (sk[126]) & (!g392) & (!g863)) + ((g25) & (!g164) & (!g402) & (sk[126]) & (g392) & (!g863)) + ((g25) & (!g164) & (g402) & (!sk[126]) & (!g392) & (g863)) + ((g25) & (!g164) & (g402) & (!sk[126]) & (g392) & (!g863)) + ((g25) & (!g164) & (g402) & (!sk[126]) & (g392) & (g863)) + ((g25) & (!g164) & (g402) & (sk[126]) & (!g392) & (!g863)) + ((g25) & (!g164) & (g402) & (sk[126]) & (g392) & (!g863)) + ((g25) & (g164) & (!g402) & (!sk[126]) & (!g392) & (!g863)) + ((g25) & (g164) & (!g402) & (!sk[126]) & (!g392) & (g863)) + ((g25) & (g164) & (!g402) & (!sk[126]) & (g392) & (!g863)) + ((g25) & (g164) & (!g402) & (!sk[126]) & (g392) & (g863)) + ((g25) & (g164) & (!g402) & (sk[126]) & (!g392) & (!g863)) + ((g25) & (g164) & (!g402) & (sk[126]) & (g392) & (!g863)) + ((g25) & (g164) & (g402) & (!sk[126]) & (!g392) & (!g863)) + ((g25) & (g164) & (g402) & (!sk[126]) & (!g392) & (g863)) + ((g25) & (g164) & (g402) & (!sk[126]) & (g392) & (!g863)) + ((g25) & (g164) & (g402) & (!sk[126]) & (g392) & (g863)) + ((g25) & (g164) & (g402) & (sk[126]) & (!g392) & (!g863)) + ((g25) & (g164) & (g402) & (sk[126]) & (g392) & (!g863)));
	assign g865 = (((!i_12_) & (!i_13_) & (!sk[127]) & (i_14_) & (!g20)) + ((!i_12_) & (!i_13_) & (!sk[127]) & (i_14_) & (g20)) + ((!i_12_) & (i_13_) & (!sk[127]) & (i_14_) & (!g20)) + ((!i_12_) & (i_13_) & (!sk[127]) & (i_14_) & (g20)) + ((!i_12_) & (i_13_) & (sk[127]) & (!i_14_) & (g20)) + ((i_12_) & (!i_13_) & (!sk[127]) & (i_14_) & (!g20)) + ((i_12_) & (!i_13_) & (!sk[127]) & (i_14_) & (g20)) + ((i_12_) & (!i_13_) & (sk[127]) & (!i_14_) & (g20)) + ((i_12_) & (i_13_) & (!sk[127]) & (i_14_) & (!g20)) + ((i_12_) & (i_13_) & (!sk[127]) & (i_14_) & (g20)) + ((i_12_) & (i_13_) & (sk[127]) & (!i_14_) & (g20)));
	assign g866 = (((!g123) & (!sk[0]) & (!g130) & (g849) & (!g853)) + ((!g123) & (!sk[0]) & (!g130) & (g849) & (g853)) + ((!g123) & (!sk[0]) & (g130) & (g849) & (!g853)) + ((!g123) & (!sk[0]) & (g130) & (g849) & (g853)) + ((!g123) & (sk[0]) & (!g130) & (!g849) & (!g853)) + ((!g123) & (sk[0]) & (g130) & (!g849) & (!g853)) + ((!g123) & (sk[0]) & (g130) & (!g849) & (g853)) + ((g123) & (!sk[0]) & (!g130) & (g849) & (!g853)) + ((g123) & (!sk[0]) & (!g130) & (g849) & (g853)) + ((g123) & (!sk[0]) & (g130) & (g849) & (!g853)) + ((g123) & (!sk[0]) & (g130) & (g849) & (g853)) + ((g123) & (sk[0]) & (!g130) & (!g849) & (!g853)) + ((g123) & (sk[0]) & (g130) & (!g849) & (!g853)) + ((g123) & (sk[0]) & (g130) & (!g849) & (g853)) + ((g123) & (sk[0]) & (g130) & (g849) & (!g853)) + ((g123) & (sk[0]) & (g130) & (g849) & (g853)));
	assign g867 = (((!g4) & (!g126) & (!sk[1]) & (g91) & (!g105) & (g309)) + ((!g4) & (!g126) & (!sk[1]) & (g91) & (g105) & (!g309)) + ((!g4) & (!g126) & (!sk[1]) & (g91) & (g105) & (g309)) + ((!g4) & (!g126) & (sk[1]) & (!g91) & (!g105) & (g309)) + ((!g4) & (!g126) & (sk[1]) & (g91) & (!g105) & (g309)) + ((!g4) & (g126) & (!sk[1]) & (!g91) & (!g105) & (!g309)) + ((!g4) & (g126) & (!sk[1]) & (!g91) & (!g105) & (g309)) + ((!g4) & (g126) & (!sk[1]) & (!g91) & (g105) & (!g309)) + ((!g4) & (g126) & (!sk[1]) & (!g91) & (g105) & (g309)) + ((!g4) & (g126) & (!sk[1]) & (g91) & (!g105) & (!g309)) + ((!g4) & (g126) & (!sk[1]) & (g91) & (!g105) & (g309)) + ((!g4) & (g126) & (!sk[1]) & (g91) & (g105) & (!g309)) + ((!g4) & (g126) & (!sk[1]) & (g91) & (g105) & (g309)) + ((!g4) & (g126) & (sk[1]) & (!g91) & (!g105) & (g309)) + ((!g4) & (g126) & (sk[1]) & (g91) & (!g105) & (g309)) + ((g4) & (!g126) & (!sk[1]) & (g91) & (!g105) & (g309)) + ((g4) & (!g126) & (!sk[1]) & (g91) & (g105) & (!g309)) + ((g4) & (!g126) & (!sk[1]) & (g91) & (g105) & (g309)) + ((g4) & (!g126) & (sk[1]) & (!g91) & (!g105) & (!g309)) + ((g4) & (!g126) & (sk[1]) & (!g91) & (!g105) & (g309)) + ((g4) & (!g126) & (sk[1]) & (g91) & (!g105) & (!g309)) + ((g4) & (!g126) & (sk[1]) & (g91) & (!g105) & (g309)) + ((g4) & (g126) & (!sk[1]) & (!g91) & (!g105) & (!g309)) + ((g4) & (g126) & (!sk[1]) & (!g91) & (!g105) & (g309)) + ((g4) & (g126) & (!sk[1]) & (!g91) & (g105) & (!g309)) + ((g4) & (g126) & (!sk[1]) & (!g91) & (g105) & (g309)) + ((g4) & (g126) & (!sk[1]) & (g91) & (!g105) & (!g309)) + ((g4) & (g126) & (!sk[1]) & (g91) & (!g105) & (g309)) + ((g4) & (g126) & (!sk[1]) & (g91) & (g105) & (!g309)) + ((g4) & (g126) & (!sk[1]) & (g91) & (g105) & (g309)) + ((g4) & (g126) & (sk[1]) & (!g91) & (!g105) & (!g309)) + ((g4) & (g126) & (sk[1]) & (!g91) & (!g105) & (g309)) + ((g4) & (g126) & (sk[1]) & (g91) & (!g105) & (g309)));
	assign g868 = (((!g123) & (!g850) & (!g865) & (sk[2]) & (g866) & (!g867)) + ((!g123) & (!g850) & (g865) & (!sk[2]) & (!g866) & (g867)) + ((!g123) & (!g850) & (g865) & (!sk[2]) & (g866) & (!g867)) + ((!g123) & (!g850) & (g865) & (!sk[2]) & (g866) & (g867)) + ((!g123) & (g850) & (!g865) & (!sk[2]) & (!g866) & (!g867)) + ((!g123) & (g850) & (!g865) & (!sk[2]) & (!g866) & (g867)) + ((!g123) & (g850) & (!g865) & (!sk[2]) & (g866) & (!g867)) + ((!g123) & (g850) & (!g865) & (!sk[2]) & (g866) & (g867)) + ((!g123) & (g850) & (g865) & (!sk[2]) & (!g866) & (!g867)) + ((!g123) & (g850) & (g865) & (!sk[2]) & (!g866) & (g867)) + ((!g123) & (g850) & (g865) & (!sk[2]) & (g866) & (!g867)) + ((!g123) & (g850) & (g865) & (!sk[2]) & (g866) & (g867)) + ((g123) & (!g850) & (!g865) & (sk[2]) & (g866) & (!g867)) + ((g123) & (!g850) & (g865) & (!sk[2]) & (!g866) & (g867)) + ((g123) & (!g850) & (g865) & (!sk[2]) & (g866) & (!g867)) + ((g123) & (!g850) & (g865) & (!sk[2]) & (g866) & (g867)) + ((g123) & (!g850) & (g865) & (sk[2]) & (g866) & (!g867)) + ((g123) & (g850) & (!g865) & (!sk[2]) & (!g866) & (!g867)) + ((g123) & (g850) & (!g865) & (!sk[2]) & (!g866) & (g867)) + ((g123) & (g850) & (!g865) & (!sk[2]) & (g866) & (!g867)) + ((g123) & (g850) & (!g865) & (!sk[2]) & (g866) & (g867)) + ((g123) & (g850) & (!g865) & (sk[2]) & (g866) & (!g867)) + ((g123) & (g850) & (g865) & (!sk[2]) & (!g866) & (!g867)) + ((g123) & (g850) & (g865) & (!sk[2]) & (!g866) & (g867)) + ((g123) & (g850) & (g865) & (!sk[2]) & (g866) & (!g867)) + ((g123) & (g850) & (g865) & (!sk[2]) & (g866) & (g867)) + ((g123) & (g850) & (g865) & (sk[2]) & (g866) & (!g867)));
	assign g869 = (((!i_9_) & (!sk[3]) & (!i_10_) & (i_11_) & (!i_15_) & (g735)) + ((!i_9_) & (!sk[3]) & (!i_10_) & (i_11_) & (i_15_) & (!g735)) + ((!i_9_) & (!sk[3]) & (!i_10_) & (i_11_) & (i_15_) & (g735)) + ((!i_9_) & (!sk[3]) & (i_10_) & (!i_11_) & (!i_15_) & (!g735)) + ((!i_9_) & (!sk[3]) & (i_10_) & (!i_11_) & (!i_15_) & (g735)) + ((!i_9_) & (!sk[3]) & (i_10_) & (!i_11_) & (i_15_) & (!g735)) + ((!i_9_) & (!sk[3]) & (i_10_) & (!i_11_) & (i_15_) & (g735)) + ((!i_9_) & (!sk[3]) & (i_10_) & (i_11_) & (!i_15_) & (!g735)) + ((!i_9_) & (!sk[3]) & (i_10_) & (i_11_) & (!i_15_) & (g735)) + ((!i_9_) & (!sk[3]) & (i_10_) & (i_11_) & (i_15_) & (!g735)) + ((!i_9_) & (!sk[3]) & (i_10_) & (i_11_) & (i_15_) & (g735)) + ((!i_9_) & (sk[3]) & (!i_10_) & (i_11_) & (!i_15_) & (g735)) + ((i_9_) & (!sk[3]) & (!i_10_) & (i_11_) & (!i_15_) & (g735)) + ((i_9_) & (!sk[3]) & (!i_10_) & (i_11_) & (i_15_) & (!g735)) + ((i_9_) & (!sk[3]) & (!i_10_) & (i_11_) & (i_15_) & (g735)) + ((i_9_) & (!sk[3]) & (i_10_) & (!i_11_) & (!i_15_) & (!g735)) + ((i_9_) & (!sk[3]) & (i_10_) & (!i_11_) & (!i_15_) & (g735)) + ((i_9_) & (!sk[3]) & (i_10_) & (!i_11_) & (i_15_) & (!g735)) + ((i_9_) & (!sk[3]) & (i_10_) & (!i_11_) & (i_15_) & (g735)) + ((i_9_) & (!sk[3]) & (i_10_) & (i_11_) & (!i_15_) & (!g735)) + ((i_9_) & (!sk[3]) & (i_10_) & (i_11_) & (!i_15_) & (g735)) + ((i_9_) & (!sk[3]) & (i_10_) & (i_11_) & (i_15_) & (!g735)) + ((i_9_) & (!sk[3]) & (i_10_) & (i_11_) & (i_15_) & (g735)) + ((i_9_) & (sk[3]) & (!i_10_) & (!i_11_) & (!i_15_) & (g735)));
	assign g870 = (((!sk[4]) & (!g24) & (!g113) & (g492)) + ((!sk[4]) & (!g24) & (g113) & (!g492)) + ((!sk[4]) & (!g24) & (g113) & (g492)) + ((!sk[4]) & (g24) & (!g113) & (g492)) + ((!sk[4]) & (g24) & (g113) & (!g492)) + ((!sk[4]) & (g24) & (g113) & (g492)) + ((sk[4]) & (!g24) & (g113) & (!g492)) + ((sk[4]) & (g24) & (!g113) & (!g492)) + ((sk[4]) & (g24) & (g113) & (!g492)));
	assign g871 = (((!g24) & (!sk[5]) & (!g35) & (g161) & (!g68)) + ((!g24) & (!sk[5]) & (!g35) & (g161) & (g68)) + ((!g24) & (!sk[5]) & (g35) & (g161) & (!g68)) + ((!g24) & (!sk[5]) & (g35) & (g161) & (g68)) + ((!g24) & (sk[5]) & (g35) & (g161) & (!g68)) + ((!g24) & (sk[5]) & (g35) & (g161) & (g68)) + ((g24) & (!sk[5]) & (!g35) & (g161) & (!g68)) + ((g24) & (!sk[5]) & (!g35) & (g161) & (g68)) + ((g24) & (!sk[5]) & (g35) & (g161) & (!g68)) + ((g24) & (!sk[5]) & (g35) & (g161) & (g68)) + ((g24) & (sk[5]) & (g35) & (g161) & (!g68)));
	assign g872 = (((!sk[6]) & (!g257) & (!g351) & (g869) & (!g870) & (g871)) + ((!sk[6]) & (!g257) & (!g351) & (g869) & (g870) & (!g871)) + ((!sk[6]) & (!g257) & (!g351) & (g869) & (g870) & (g871)) + ((!sk[6]) & (!g257) & (g351) & (!g869) & (!g870) & (!g871)) + ((!sk[6]) & (!g257) & (g351) & (!g869) & (!g870) & (g871)) + ((!sk[6]) & (!g257) & (g351) & (!g869) & (g870) & (!g871)) + ((!sk[6]) & (!g257) & (g351) & (!g869) & (g870) & (g871)) + ((!sk[6]) & (!g257) & (g351) & (g869) & (!g870) & (!g871)) + ((!sk[6]) & (!g257) & (g351) & (g869) & (!g870) & (g871)) + ((!sk[6]) & (!g257) & (g351) & (g869) & (g870) & (!g871)) + ((!sk[6]) & (!g257) & (g351) & (g869) & (g870) & (g871)) + ((!sk[6]) & (g257) & (!g351) & (g869) & (!g870) & (g871)) + ((!sk[6]) & (g257) & (!g351) & (g869) & (g870) & (!g871)) + ((!sk[6]) & (g257) & (!g351) & (g869) & (g870) & (g871)) + ((!sk[6]) & (g257) & (g351) & (!g869) & (!g870) & (!g871)) + ((!sk[6]) & (g257) & (g351) & (!g869) & (!g870) & (g871)) + ((!sk[6]) & (g257) & (g351) & (!g869) & (g870) & (!g871)) + ((!sk[6]) & (g257) & (g351) & (!g869) & (g870) & (g871)) + ((!sk[6]) & (g257) & (g351) & (g869) & (!g870) & (!g871)) + ((!sk[6]) & (g257) & (g351) & (g869) & (!g870) & (g871)) + ((!sk[6]) & (g257) & (g351) & (g869) & (g870) & (!g871)) + ((!sk[6]) & (g257) & (g351) & (g869) & (g870) & (g871)) + ((sk[6]) & (!g257) & (!g351) & (!g869) & (g870) & (!g871)) + ((sk[6]) & (!g257) & (!g351) & (g869) & (g870) & (!g871)) + ((sk[6]) & (!g257) & (g351) & (!g869) & (!g870) & (!g871)) + ((sk[6]) & (!g257) & (g351) & (!g869) & (g870) & (!g871)) + ((sk[6]) & (!g257) & (g351) & (g869) & (!g870) & (!g871)) + ((sk[6]) & (!g257) & (g351) & (g869) & (g870) & (!g871)) + ((sk[6]) & (g257) & (!g351) & (!g869) & (g870) & (!g871)) + ((sk[6]) & (g257) & (g351) & (!g869) & (!g870) & (!g871)) + ((sk[6]) & (g257) & (g351) & (!g869) & (g870) & (!g871)));
	assign g873 = (((!sk[7]) & (!g856) & (!g859) & (g1501) & (!g864) & (g1488)) + ((!sk[7]) & (!g856) & (!g859) & (g1501) & (g864) & (!g1488)) + ((!sk[7]) & (!g856) & (!g859) & (g1501) & (g864) & (g1488)) + ((!sk[7]) & (!g856) & (g859) & (!g1501) & (!g864) & (!g1488)) + ((!sk[7]) & (!g856) & (g859) & (!g1501) & (!g864) & (g1488)) + ((!sk[7]) & (!g856) & (g859) & (!g1501) & (g864) & (!g1488)) + ((!sk[7]) & (!g856) & (g859) & (!g1501) & (g864) & (g1488)) + ((!sk[7]) & (!g856) & (g859) & (g1501) & (!g864) & (!g1488)) + ((!sk[7]) & (!g856) & (g859) & (g1501) & (!g864) & (g1488)) + ((!sk[7]) & (!g856) & (g859) & (g1501) & (g864) & (!g1488)) + ((!sk[7]) & (!g856) & (g859) & (g1501) & (g864) & (g1488)) + ((!sk[7]) & (g856) & (!g859) & (g1501) & (!g864) & (g1488)) + ((!sk[7]) & (g856) & (!g859) & (g1501) & (g864) & (!g1488)) + ((!sk[7]) & (g856) & (!g859) & (g1501) & (g864) & (g1488)) + ((!sk[7]) & (g856) & (g859) & (!g1501) & (!g864) & (!g1488)) + ((!sk[7]) & (g856) & (g859) & (!g1501) & (!g864) & (g1488)) + ((!sk[7]) & (g856) & (g859) & (!g1501) & (g864) & (!g1488)) + ((!sk[7]) & (g856) & (g859) & (!g1501) & (g864) & (g1488)) + ((!sk[7]) & (g856) & (g859) & (g1501) & (!g864) & (!g1488)) + ((!sk[7]) & (g856) & (g859) & (g1501) & (!g864) & (g1488)) + ((!sk[7]) & (g856) & (g859) & (g1501) & (g864) & (!g1488)) + ((!sk[7]) & (g856) & (g859) & (g1501) & (g864) & (g1488)) + ((sk[7]) & (g856) & (g859) & (g1501) & (g864) & (g1488)));
	assign g874 = (((!g159) & (!sk[8]) & (!g847) & (g850) & (!g865)) + ((!g159) & (!sk[8]) & (!g847) & (g850) & (g865)) + ((!g159) & (!sk[8]) & (g847) & (g850) & (!g865)) + ((!g159) & (!sk[8]) & (g847) & (g850) & (g865)) + ((!g159) & (sk[8]) & (!g847) & (!g850) & (!g865)) + ((!g159) & (sk[8]) & (!g847) & (!g850) & (g865)) + ((!g159) & (sk[8]) & (!g847) & (g850) & (!g865)) + ((!g159) & (sk[8]) & (!g847) & (g850) & (g865)) + ((!g159) & (sk[8]) & (g847) & (!g850) & (g865)) + ((!g159) & (sk[8]) & (g847) & (g850) & (!g865)) + ((!g159) & (sk[8]) & (g847) & (g850) & (g865)) + ((g159) & (!sk[8]) & (!g847) & (g850) & (!g865)) + ((g159) & (!sk[8]) & (!g847) & (g850) & (g865)) + ((g159) & (!sk[8]) & (g847) & (g850) & (!g865)) + ((g159) & (!sk[8]) & (g847) & (g850) & (g865)));
	assign g875 = (((!i_12_) & (!sk[9]) & (!i_13_) & (i_14_) & (!g27)) + ((!i_12_) & (!sk[9]) & (!i_13_) & (i_14_) & (g27)) + ((!i_12_) & (!sk[9]) & (i_13_) & (i_14_) & (!g27)) + ((!i_12_) & (!sk[9]) & (i_13_) & (i_14_) & (g27)) + ((!i_12_) & (sk[9]) & (i_13_) & (!i_14_) & (g27)) + ((i_12_) & (!sk[9]) & (!i_13_) & (i_14_) & (!g27)) + ((i_12_) & (!sk[9]) & (!i_13_) & (i_14_) & (g27)) + ((i_12_) & (!sk[9]) & (i_13_) & (i_14_) & (!g27)) + ((i_12_) & (!sk[9]) & (i_13_) & (i_14_) & (g27)) + ((i_12_) & (sk[9]) & (!i_13_) & (!i_14_) & (g27)) + ((i_12_) & (sk[9]) & (i_13_) & (!i_14_) & (g27)));
	assign g876 = (((!g159) & (!sk[10]) & (!g852) & (g853) & (!g875)) + ((!g159) & (!sk[10]) & (!g852) & (g853) & (g875)) + ((!g159) & (!sk[10]) & (g852) & (g853) & (!g875)) + ((!g159) & (!sk[10]) & (g852) & (g853) & (g875)) + ((!g159) & (sk[10]) & (!g852) & (!g853) & (g875)) + ((!g159) & (sk[10]) & (!g852) & (g853) & (!g875)) + ((!g159) & (sk[10]) & (!g852) & (g853) & (g875)) + ((!g159) & (sk[10]) & (g852) & (!g853) & (!g875)) + ((!g159) & (sk[10]) & (g852) & (!g853) & (g875)) + ((!g159) & (sk[10]) & (g852) & (g853) & (!g875)) + ((!g159) & (sk[10]) & (g852) & (g853) & (g875)) + ((g159) & (!sk[10]) & (!g852) & (g853) & (!g875)) + ((g159) & (!sk[10]) & (!g852) & (g853) & (g875)) + ((g159) & (!sk[10]) & (g852) & (g853) & (!g875)) + ((g159) & (!sk[10]) & (g852) & (g853) & (g875)));
	assign g877 = (((!g3) & (!i_12_) & (i_13_) & (!sk[11]) & (!i_14_)) + ((!g3) & (!i_12_) & (i_13_) & (!sk[11]) & (i_14_)) + ((!g3) & (i_12_) & (i_13_) & (!sk[11]) & (!i_14_)) + ((!g3) & (i_12_) & (i_13_) & (!sk[11]) & (i_14_)) + ((g3) & (!i_12_) & (i_13_) & (!sk[11]) & (!i_14_)) + ((g3) & (!i_12_) & (i_13_) & (!sk[11]) & (i_14_)) + ((g3) & (!i_12_) & (i_13_) & (sk[11]) & (!i_14_)) + ((g3) & (i_12_) & (!i_13_) & (sk[11]) & (!i_14_)) + ((g3) & (i_12_) & (i_13_) & (!sk[11]) & (!i_14_)) + ((g3) & (i_12_) & (i_13_) & (!sk[11]) & (i_14_)) + ((g3) & (i_12_) & (i_13_) & (sk[11]) & (!i_14_)));
	assign g878 = (((!sk[12]) & (!g154) & (!g849) & (g851)) + ((!sk[12]) & (!g154) & (g849) & (!g851)) + ((!sk[12]) & (!g154) & (g849) & (g851)) + ((!sk[12]) & (g154) & (!g849) & (g851)) + ((!sk[12]) & (g154) & (g849) & (!g851)) + ((!sk[12]) & (g154) & (g849) & (g851)) + ((sk[12]) & (!g154) & (!g849) & (!g851)) + ((sk[12]) & (!g154) & (g849) & (!g851)) + ((sk[12]) & (!g154) & (g849) & (g851)));
	assign g879 = (((!g154) & (!g877) & (!g850) & (!g865) & (sk[13]) & (!g878)) + ((!g154) & (!g877) & (g850) & (!g865) & (!sk[13]) & (g878)) + ((!g154) & (!g877) & (g850) & (g865) & (!sk[13]) & (!g878)) + ((!g154) & (!g877) & (g850) & (g865) & (!sk[13]) & (g878)) + ((!g154) & (g877) & (!g850) & (!g865) & (!sk[13]) & (!g878)) + ((!g154) & (g877) & (!g850) & (!g865) & (!sk[13]) & (g878)) + ((!g154) & (g877) & (!g850) & (g865) & (!sk[13]) & (!g878)) + ((!g154) & (g877) & (!g850) & (g865) & (!sk[13]) & (g878)) + ((!g154) & (g877) & (g850) & (!g865) & (!sk[13]) & (!g878)) + ((!g154) & (g877) & (g850) & (!g865) & (!sk[13]) & (g878)) + ((!g154) & (g877) & (g850) & (g865) & (!sk[13]) & (!g878)) + ((!g154) & (g877) & (g850) & (g865) & (!sk[13]) & (g878)) + ((g154) & (!g877) & (!g850) & (!g865) & (sk[13]) & (!g878)) + ((g154) & (!g877) & (!g850) & (g865) & (sk[13]) & (!g878)) + ((g154) & (!g877) & (g850) & (!g865) & (!sk[13]) & (g878)) + ((g154) & (!g877) & (g850) & (!g865) & (sk[13]) & (!g878)) + ((g154) & (!g877) & (g850) & (g865) & (!sk[13]) & (!g878)) + ((g154) & (!g877) & (g850) & (g865) & (!sk[13]) & (g878)) + ((g154) & (!g877) & (g850) & (g865) & (sk[13]) & (!g878)) + ((g154) & (g877) & (!g850) & (!g865) & (!sk[13]) & (!g878)) + ((g154) & (g877) & (!g850) & (!g865) & (!sk[13]) & (g878)) + ((g154) & (g877) & (!g850) & (!g865) & (sk[13]) & (!g878)) + ((g154) & (g877) & (!g850) & (g865) & (!sk[13]) & (!g878)) + ((g154) & (g877) & (!g850) & (g865) & (!sk[13]) & (g878)) + ((g154) & (g877) & (!g850) & (g865) & (sk[13]) & (!g878)) + ((g154) & (g877) & (g850) & (!g865) & (!sk[13]) & (!g878)) + ((g154) & (g877) & (g850) & (!g865) & (!sk[13]) & (g878)) + ((g154) & (g877) & (g850) & (!g865) & (sk[13]) & (!g878)) + ((g154) & (g877) & (g850) & (g865) & (!sk[13]) & (!g878)) + ((g154) & (g877) & (g850) & (g865) & (!sk[13]) & (g878)) + ((g154) & (g877) & (g850) & (g865) & (sk[13]) & (!g878)));
	assign g880 = (((!g154) & (g847) & (g848) & (!g874) & (!g876) & (g879)) + ((g154) & (!g847) & (!g848) & (!g874) & (!g876) & (g879)) + ((g154) & (!g847) & (g848) & (!g874) & (!g876) & (g879)) + ((g154) & (g847) & (!g848) & (!g874) & (!g876) & (g879)) + ((g154) & (g847) & (g848) & (!g874) & (!g876) & (g879)));
	assign g881 = (((!i_12_) & (!i_13_) & (i_14_) & (!sk[15]) & (!g126)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[15]) & (g126)) + ((!i_12_) & (i_13_) & (!i_14_) & (sk[15]) & (!g126)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[15]) & (!g126)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[15]) & (g126)) + ((i_12_) & (!i_13_) & (!i_14_) & (sk[15]) & (!g126)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[15]) & (!g126)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[15]) & (g126)) + ((i_12_) & (i_13_) & (!i_14_) & (sk[15]) & (!g126)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[15]) & (!g126)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[15]) & (g126)));
	assign g882 = (((!i_9_) & (!i_10_) & (i_11_) & (!sk[16]) & (!i_15_) & (g460)) + ((!i_9_) & (!i_10_) & (i_11_) & (!sk[16]) & (i_15_) & (!g460)) + ((!i_9_) & (!i_10_) & (i_11_) & (!sk[16]) & (i_15_) & (g460)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[16]) & (!i_15_) & (!g460)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[16]) & (!i_15_) & (g460)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[16]) & (i_15_) & (!g460)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[16]) & (i_15_) & (g460)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[16]) & (!i_15_) & (!g460)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[16]) & (!i_15_) & (g460)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[16]) & (i_15_) & (!g460)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[16]) & (i_15_) & (g460)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[16]) & (!i_15_) & (g460)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[16]) & (i_15_) & (!g460)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[16]) & (i_15_) & (g460)) + ((i_9_) & (!i_10_) & (i_11_) & (sk[16]) & (!i_15_) & (!g460)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[16]) & (!i_15_) & (!g460)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[16]) & (!i_15_) & (g460)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[16]) & (i_15_) & (!g460)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[16]) & (i_15_) & (g460)) + ((i_9_) & (i_10_) & (!i_11_) & (sk[16]) & (!i_15_) & (!g460)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[16]) & (!i_15_) & (!g460)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[16]) & (!i_15_) & (g460)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[16]) & (i_15_) & (!g460)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[16]) & (i_15_) & (g460)) + ((i_9_) & (i_10_) & (i_11_) & (sk[16]) & (!i_15_) & (!g460)));
	assign g883 = (((!sk[17]) & (!g24) & (!g144) & (g126) & (!g402) & (g882)) + ((!sk[17]) & (!g24) & (!g144) & (g126) & (g402) & (!g882)) + ((!sk[17]) & (!g24) & (!g144) & (g126) & (g402) & (g882)) + ((!sk[17]) & (!g24) & (g144) & (!g126) & (!g402) & (!g882)) + ((!sk[17]) & (!g24) & (g144) & (!g126) & (!g402) & (g882)) + ((!sk[17]) & (!g24) & (g144) & (!g126) & (g402) & (!g882)) + ((!sk[17]) & (!g24) & (g144) & (!g126) & (g402) & (g882)) + ((!sk[17]) & (!g24) & (g144) & (g126) & (!g402) & (!g882)) + ((!sk[17]) & (!g24) & (g144) & (g126) & (!g402) & (g882)) + ((!sk[17]) & (!g24) & (g144) & (g126) & (g402) & (!g882)) + ((!sk[17]) & (!g24) & (g144) & (g126) & (g402) & (g882)) + ((!sk[17]) & (g24) & (!g144) & (g126) & (!g402) & (g882)) + ((!sk[17]) & (g24) & (!g144) & (g126) & (g402) & (!g882)) + ((!sk[17]) & (g24) & (!g144) & (g126) & (g402) & (g882)) + ((!sk[17]) & (g24) & (g144) & (!g126) & (!g402) & (!g882)) + ((!sk[17]) & (g24) & (g144) & (!g126) & (!g402) & (g882)) + ((!sk[17]) & (g24) & (g144) & (!g126) & (g402) & (!g882)) + ((!sk[17]) & (g24) & (g144) & (!g126) & (g402) & (g882)) + ((!sk[17]) & (g24) & (g144) & (g126) & (!g402) & (!g882)) + ((!sk[17]) & (g24) & (g144) & (g126) & (!g402) & (g882)) + ((!sk[17]) & (g24) & (g144) & (g126) & (g402) & (!g882)) + ((!sk[17]) & (g24) & (g144) & (g126) & (g402) & (g882)) + ((sk[17]) & (!g24) & (!g144) & (!g126) & (!g402) & (!g882)) + ((sk[17]) & (!g24) & (!g144) & (!g126) & (!g402) & (g882)) + ((sk[17]) & (!g24) & (g144) & (!g126) & (!g402) & (!g882)) + ((sk[17]) & (!g24) & (g144) & (!g126) & (!g402) & (g882)) + ((sk[17]) & (!g24) & (g144) & (!g126) & (g402) & (g882)) + ((sk[17]) & (!g24) & (g144) & (g126) & (!g402) & (g882)) + ((sk[17]) & (!g24) & (g144) & (g126) & (g402) & (g882)) + ((sk[17]) & (g24) & (g144) & (!g126) & (!g402) & (g882)) + ((sk[17]) & (g24) & (g144) & (!g126) & (g402) & (g882)) + ((sk[17]) & (g24) & (g144) & (g126) & (!g402) & (g882)) + ((sk[17]) & (g24) & (g144) & (g126) & (g402) & (g882)));
	assign g884 = (((!g257) & (!g356) & (!sk[18]) & (g881) & (!g883)) + ((!g257) & (!g356) & (!sk[18]) & (g881) & (g883)) + ((!g257) & (!g356) & (sk[18]) & (!g881) & (!g883)) + ((!g257) & (!g356) & (sk[18]) & (g881) & (!g883)) + ((!g257) & (g356) & (!sk[18]) & (g881) & (!g883)) + ((!g257) & (g356) & (!sk[18]) & (g881) & (g883)) + ((!g257) & (g356) & (sk[18]) & (!g881) & (!g883)) + ((g257) & (!g356) & (!sk[18]) & (g881) & (!g883)) + ((g257) & (!g356) & (!sk[18]) & (g881) & (g883)) + ((g257) & (!g356) & (sk[18]) & (!g881) & (!g883)) + ((g257) & (g356) & (!sk[18]) & (g881) & (!g883)) + ((g257) & (g356) & (!sk[18]) & (g881) & (g883)) + ((g257) & (g356) & (sk[18]) & (!g881) & (!g883)));
	assign g885 = (((!sk[19]) & (!g125) & (!g159) & (g438) & (!g472) & (g877)) + ((!sk[19]) & (!g125) & (!g159) & (g438) & (g472) & (!g877)) + ((!sk[19]) & (!g125) & (!g159) & (g438) & (g472) & (g877)) + ((!sk[19]) & (!g125) & (g159) & (!g438) & (!g472) & (!g877)) + ((!sk[19]) & (!g125) & (g159) & (!g438) & (!g472) & (g877)) + ((!sk[19]) & (!g125) & (g159) & (!g438) & (g472) & (!g877)) + ((!sk[19]) & (!g125) & (g159) & (!g438) & (g472) & (g877)) + ((!sk[19]) & (!g125) & (g159) & (g438) & (!g472) & (!g877)) + ((!sk[19]) & (!g125) & (g159) & (g438) & (!g472) & (g877)) + ((!sk[19]) & (!g125) & (g159) & (g438) & (g472) & (!g877)) + ((!sk[19]) & (!g125) & (g159) & (g438) & (g472) & (g877)) + ((!sk[19]) & (g125) & (!g159) & (g438) & (!g472) & (g877)) + ((!sk[19]) & (g125) & (!g159) & (g438) & (g472) & (!g877)) + ((!sk[19]) & (g125) & (!g159) & (g438) & (g472) & (g877)) + ((!sk[19]) & (g125) & (g159) & (!g438) & (!g472) & (!g877)) + ((!sk[19]) & (g125) & (g159) & (!g438) & (!g472) & (g877)) + ((!sk[19]) & (g125) & (g159) & (!g438) & (g472) & (!g877)) + ((!sk[19]) & (g125) & (g159) & (!g438) & (g472) & (g877)) + ((!sk[19]) & (g125) & (g159) & (g438) & (!g472) & (!g877)) + ((!sk[19]) & (g125) & (g159) & (g438) & (!g472) & (g877)) + ((!sk[19]) & (g125) & (g159) & (g438) & (g472) & (!g877)) + ((!sk[19]) & (g125) & (g159) & (g438) & (g472) & (g877)) + ((sk[19]) & (!g125) & (!g159) & (!g438) & (!g472) & (!g877)) + ((sk[19]) & (!g125) & (!g159) & (g438) & (!g472) & (!g877)) + ((sk[19]) & (!g125) & (!g159) & (g438) & (g472) & (!g877)) + ((sk[19]) & (!g125) & (g159) & (!g438) & (!g472) & (!g877)) + ((sk[19]) & (!g125) & (g159) & (g438) & (!g472) & (!g877)) + ((sk[19]) & (!g125) & (g159) & (g438) & (!g472) & (g877)) + ((sk[19]) & (!g125) & (g159) & (g438) & (g472) & (!g877)) + ((sk[19]) & (!g125) & (g159) & (g438) & (g472) & (g877)) + ((sk[19]) & (g125) & (!g159) & (!g438) & (!g472) & (!g877)) + ((sk[19]) & (g125) & (!g159) & (g438) & (!g472) & (!g877)) + ((sk[19]) & (g125) & (g159) & (!g438) & (!g472) & (!g877)) + ((sk[19]) & (g125) & (g159) & (g438) & (!g472) & (!g877)) + ((sk[19]) & (g125) & (g159) & (g438) & (!g472) & (g877)));
	assign g886 = (((!g480) & (!g880) & (g884) & (!sk[20]) & (!g885)) + ((!g480) & (!g880) & (g884) & (!sk[20]) & (g885)) + ((!g480) & (g880) & (g884) & (!sk[20]) & (!g885)) + ((!g480) & (g880) & (g884) & (!sk[20]) & (g885)) + ((g480) & (!g880) & (g884) & (!sk[20]) & (!g885)) + ((g480) & (!g880) & (g884) & (!sk[20]) & (g885)) + ((g480) & (g880) & (g884) & (!sk[20]) & (!g885)) + ((g480) & (g880) & (g884) & (!sk[20]) & (g885)) + ((g480) & (g880) & (g884) & (sk[20]) & (g885)));
	assign g887 = (((g102) & (!sk[21]) & (!g881)) + ((g102) & (!sk[21]) & (g881)) + ((g102) & (sk[21]) & (g881)));
	assign g888 = (((!i_12_) & (!sk[22]) & (!i_13_) & (i_14_) & (!g35) & (g102)) + ((!i_12_) & (!sk[22]) & (!i_13_) & (i_14_) & (g35) & (!g102)) + ((!i_12_) & (!sk[22]) & (!i_13_) & (i_14_) & (g35) & (g102)) + ((!i_12_) & (!sk[22]) & (i_13_) & (!i_14_) & (!g35) & (!g102)) + ((!i_12_) & (!sk[22]) & (i_13_) & (!i_14_) & (!g35) & (g102)) + ((!i_12_) & (!sk[22]) & (i_13_) & (!i_14_) & (g35) & (!g102)) + ((!i_12_) & (!sk[22]) & (i_13_) & (!i_14_) & (g35) & (g102)) + ((!i_12_) & (!sk[22]) & (i_13_) & (i_14_) & (!g35) & (!g102)) + ((!i_12_) & (!sk[22]) & (i_13_) & (i_14_) & (!g35) & (g102)) + ((!i_12_) & (!sk[22]) & (i_13_) & (i_14_) & (g35) & (!g102)) + ((!i_12_) & (!sk[22]) & (i_13_) & (i_14_) & (g35) & (g102)) + ((!i_12_) & (sk[22]) & (i_13_) & (!i_14_) & (g35) & (g102)) + ((i_12_) & (!sk[22]) & (!i_13_) & (i_14_) & (!g35) & (g102)) + ((i_12_) & (!sk[22]) & (!i_13_) & (i_14_) & (g35) & (!g102)) + ((i_12_) & (!sk[22]) & (!i_13_) & (i_14_) & (g35) & (g102)) + ((i_12_) & (!sk[22]) & (i_13_) & (!i_14_) & (!g35) & (!g102)) + ((i_12_) & (!sk[22]) & (i_13_) & (!i_14_) & (!g35) & (g102)) + ((i_12_) & (!sk[22]) & (i_13_) & (!i_14_) & (g35) & (!g102)) + ((i_12_) & (!sk[22]) & (i_13_) & (!i_14_) & (g35) & (g102)) + ((i_12_) & (!sk[22]) & (i_13_) & (i_14_) & (!g35) & (!g102)) + ((i_12_) & (!sk[22]) & (i_13_) & (i_14_) & (!g35) & (g102)) + ((i_12_) & (!sk[22]) & (i_13_) & (i_14_) & (g35) & (!g102)) + ((i_12_) & (!sk[22]) & (i_13_) & (i_14_) & (g35) & (g102)) + ((i_12_) & (sk[22]) & (!i_13_) & (!i_14_) & (g35) & (g102)) + ((i_12_) & (sk[22]) & (i_13_) & (!i_14_) & (g35) & (g102)));
	assign g889 = (((!i_12_) & (!i_13_) & (i_14_) & (!sk[23]) & (!g86) & (g102)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[23]) & (g86) & (!g102)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[23]) & (g86) & (g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[23]) & (!g86) & (!g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[23]) & (!g86) & (g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[23]) & (g86) & (!g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[23]) & (g86) & (g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (sk[23]) & (g86) & (g102)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[23]) & (!g86) & (!g102)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[23]) & (!g86) & (g102)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[23]) & (g86) & (!g102)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[23]) & (g86) & (g102)) + ((i_12_) & (!i_13_) & (!i_14_) & (sk[23]) & (g86) & (g102)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[23]) & (!g86) & (g102)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[23]) & (g86) & (!g102)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[23]) & (g86) & (g102)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[23]) & (!g86) & (!g102)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[23]) & (!g86) & (g102)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[23]) & (g86) & (!g102)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[23]) & (g86) & (g102)) + ((i_12_) & (i_13_) & (!i_14_) & (sk[23]) & (g86) & (g102)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[23]) & (!g86) & (!g102)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[23]) & (!g86) & (g102)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[23]) & (g86) & (!g102)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[23]) & (g86) & (g102)));
	assign g890 = (((!i_12_) & (!i_13_) & (!sk[24]) & (i_14_) & (!g107) & (g102)) + ((!i_12_) & (!i_13_) & (!sk[24]) & (i_14_) & (g107) & (!g102)) + ((!i_12_) & (!i_13_) & (!sk[24]) & (i_14_) & (g107) & (g102)) + ((!i_12_) & (i_13_) & (!sk[24]) & (!i_14_) & (!g107) & (!g102)) + ((!i_12_) & (i_13_) & (!sk[24]) & (!i_14_) & (!g107) & (g102)) + ((!i_12_) & (i_13_) & (!sk[24]) & (!i_14_) & (g107) & (!g102)) + ((!i_12_) & (i_13_) & (!sk[24]) & (!i_14_) & (g107) & (g102)) + ((!i_12_) & (i_13_) & (!sk[24]) & (i_14_) & (!g107) & (!g102)) + ((!i_12_) & (i_13_) & (!sk[24]) & (i_14_) & (!g107) & (g102)) + ((!i_12_) & (i_13_) & (!sk[24]) & (i_14_) & (g107) & (!g102)) + ((!i_12_) & (i_13_) & (!sk[24]) & (i_14_) & (g107) & (g102)) + ((!i_12_) & (i_13_) & (sk[24]) & (!i_14_) & (!g107) & (g102)) + ((i_12_) & (!i_13_) & (!sk[24]) & (i_14_) & (!g107) & (g102)) + ((i_12_) & (!i_13_) & (!sk[24]) & (i_14_) & (g107) & (!g102)) + ((i_12_) & (!i_13_) & (!sk[24]) & (i_14_) & (g107) & (g102)) + ((i_12_) & (!i_13_) & (sk[24]) & (!i_14_) & (!g107) & (g102)) + ((i_12_) & (i_13_) & (!sk[24]) & (!i_14_) & (!g107) & (!g102)) + ((i_12_) & (i_13_) & (!sk[24]) & (!i_14_) & (!g107) & (g102)) + ((i_12_) & (i_13_) & (!sk[24]) & (!i_14_) & (g107) & (!g102)) + ((i_12_) & (i_13_) & (!sk[24]) & (!i_14_) & (g107) & (g102)) + ((i_12_) & (i_13_) & (!sk[24]) & (i_14_) & (!g107) & (!g102)) + ((i_12_) & (i_13_) & (!sk[24]) & (i_14_) & (!g107) & (g102)) + ((i_12_) & (i_13_) & (!sk[24]) & (i_14_) & (g107) & (!g102)) + ((i_12_) & (i_13_) & (!sk[24]) & (i_14_) & (g107) & (g102)) + ((i_12_) & (i_13_) & (sk[24]) & (!i_14_) & (!g107) & (g102)));
	assign g891 = (((!g3) & (!i_12_) & (i_13_) & (!i_14_) & (g35) & (!g105)) + ((!g3) & (i_12_) & (!i_13_) & (!i_14_) & (g35) & (!g105)) + ((!g3) & (i_12_) & (i_13_) & (!i_14_) & (g35) & (!g105)) + ((g3) & (!i_12_) & (i_13_) & (!i_14_) & (!g35) & (!g105)) + ((g3) & (!i_12_) & (i_13_) & (!i_14_) & (g35) & (!g105)) + ((g3) & (i_12_) & (!i_13_) & (!i_14_) & (!g35) & (!g105)) + ((g3) & (i_12_) & (!i_13_) & (!i_14_) & (g35) & (!g105)) + ((g3) & (i_12_) & (i_13_) & (!i_14_) & (!g35) & (!g105)) + ((g3) & (i_12_) & (i_13_) & (!i_14_) & (g35) & (!g105)));
	assign g892 = (((g83) & (!sk[26]) & (!g460)) + ((g83) & (!sk[26]) & (g460)) + ((g83) & (sk[26]) & (!g460)));
	assign g893 = (((!g105) & (!g295) & (!g892) & (!g700) & (!g847) & (!g852)) + ((!g105) & (!g295) & (!g892) & (!g700) & (!g847) & (g852)) + ((!g105) & (!g295) & (!g892) & (!g700) & (g847) & (!g852)) + ((!g105) & (!g295) & (!g892) & (!g700) & (g847) & (g852)) + ((!g105) & (!g295) & (!g892) & (g700) & (!g847) & (!g852)) + ((!g105) & (!g295) & (!g892) & (g700) & (!g847) & (g852)) + ((!g105) & (!g295) & (!g892) & (g700) & (g847) & (g852)) + ((!g105) & (!g295) & (g892) & (!g700) & (!g847) & (!g852)) + ((!g105) & (!g295) & (g892) & (!g700) & (!g847) & (g852)) + ((!g105) & (!g295) & (g892) & (!g700) & (g847) & (!g852)) + ((!g105) & (!g295) & (g892) & (!g700) & (g847) & (g852)) + ((!g105) & (!g295) & (g892) & (g700) & (!g847) & (!g852)) + ((!g105) & (!g295) & (g892) & (g700) & (!g847) & (g852)) + ((!g105) & (!g295) & (g892) & (g700) & (g847) & (!g852)) + ((!g105) & (!g295) & (g892) & (g700) & (g847) & (g852)) + ((!g105) & (g295) & (!g892) & (!g700) & (!g847) & (!g852)) + ((!g105) & (g295) & (!g892) & (!g700) & (!g847) & (g852)) + ((!g105) & (g295) & (!g892) & (!g700) & (g847) & (!g852)) + ((!g105) & (g295) & (!g892) & (!g700) & (g847) & (g852)) + ((!g105) & (g295) & (!g892) & (g700) & (!g847) & (!g852)) + ((!g105) & (g295) & (!g892) & (g700) & (!g847) & (g852)) + ((!g105) & (g295) & (!g892) & (g700) & (g847) & (!g852)) + ((!g105) & (g295) & (!g892) & (g700) & (g847) & (g852)) + ((!g105) & (g295) & (g892) & (!g700) & (!g847) & (!g852)) + ((!g105) & (g295) & (g892) & (!g700) & (!g847) & (g852)) + ((!g105) & (g295) & (g892) & (!g700) & (g847) & (!g852)) + ((!g105) & (g295) & (g892) & (!g700) & (g847) & (g852)) + ((!g105) & (g295) & (g892) & (g700) & (!g847) & (!g852)) + ((!g105) & (g295) & (g892) & (g700) & (!g847) & (g852)) + ((!g105) & (g295) & (g892) & (g700) & (g847) & (!g852)) + ((!g105) & (g295) & (g892) & (g700) & (g847) & (g852)));
	assign g894 = (((!sk[28]) & (!g888) & (!g889) & (g890) & (!g891) & (g893)) + ((!sk[28]) & (!g888) & (!g889) & (g890) & (g891) & (!g893)) + ((!sk[28]) & (!g888) & (!g889) & (g890) & (g891) & (g893)) + ((!sk[28]) & (!g888) & (g889) & (!g890) & (!g891) & (!g893)) + ((!sk[28]) & (!g888) & (g889) & (!g890) & (!g891) & (g893)) + ((!sk[28]) & (!g888) & (g889) & (!g890) & (g891) & (!g893)) + ((!sk[28]) & (!g888) & (g889) & (!g890) & (g891) & (g893)) + ((!sk[28]) & (!g888) & (g889) & (g890) & (!g891) & (!g893)) + ((!sk[28]) & (!g888) & (g889) & (g890) & (!g891) & (g893)) + ((!sk[28]) & (!g888) & (g889) & (g890) & (g891) & (!g893)) + ((!sk[28]) & (!g888) & (g889) & (g890) & (g891) & (g893)) + ((!sk[28]) & (g888) & (!g889) & (g890) & (!g891) & (g893)) + ((!sk[28]) & (g888) & (!g889) & (g890) & (g891) & (!g893)) + ((!sk[28]) & (g888) & (!g889) & (g890) & (g891) & (g893)) + ((!sk[28]) & (g888) & (g889) & (!g890) & (!g891) & (!g893)) + ((!sk[28]) & (g888) & (g889) & (!g890) & (!g891) & (g893)) + ((!sk[28]) & (g888) & (g889) & (!g890) & (g891) & (!g893)) + ((!sk[28]) & (g888) & (g889) & (!g890) & (g891) & (g893)) + ((!sk[28]) & (g888) & (g889) & (g890) & (!g891) & (!g893)) + ((!sk[28]) & (g888) & (g889) & (g890) & (!g891) & (g893)) + ((!sk[28]) & (g888) & (g889) & (g890) & (g891) & (!g893)) + ((!sk[28]) & (g888) & (g889) & (g890) & (g891) & (g893)) + ((sk[28]) & (!g888) & (!g889) & (!g890) & (!g891) & (!g893)));
	assign g895 = (((!g20) & (!g164) & (!sk[29]) & (g105) & (!g460)) + ((!g20) & (!g164) & (!sk[29]) & (g105) & (g460)) + ((!g20) & (g164) & (!sk[29]) & (g105) & (!g460)) + ((!g20) & (g164) & (!sk[29]) & (g105) & (g460)) + ((g20) & (!g164) & (!sk[29]) & (g105) & (!g460)) + ((g20) & (!g164) & (!sk[29]) & (g105) & (g460)) + ((g20) & (!g164) & (sk[29]) & (!g105) & (!g460)) + ((g20) & (g164) & (!sk[29]) & (g105) & (!g460)) + ((g20) & (g164) & (!sk[29]) & (g105) & (g460)) + ((g20) & (g164) & (sk[29]) & (!g105) & (!g460)) + ((g20) & (g164) & (sk[29]) & (g105) & (!g460)));
	assign g896 = (((!g159) & (!sk[30]) & (!g154) & (g849) & (!g881)) + ((!g159) & (!sk[30]) & (!g154) & (g849) & (g881)) + ((!g159) & (!sk[30]) & (g154) & (g849) & (!g881)) + ((!g159) & (!sk[30]) & (g154) & (g849) & (g881)) + ((!g159) & (sk[30]) & (!g154) & (!g849) & (!g881)) + ((!g159) & (sk[30]) & (g154) & (!g849) & (!g881)) + ((!g159) & (sk[30]) & (g154) & (!g849) & (g881)) + ((g159) & (!sk[30]) & (!g154) & (g849) & (!g881)) + ((g159) & (!sk[30]) & (!g154) & (g849) & (g881)) + ((g159) & (!sk[30]) & (g154) & (g849) & (!g881)) + ((g159) & (!sk[30]) & (g154) & (g849) & (g881)) + ((g159) & (sk[30]) & (!g154) & (!g849) & (!g881)) + ((g159) & (sk[30]) & (!g154) & (g849) & (!g881)) + ((g159) & (sk[30]) & (g154) & (!g849) & (!g881)) + ((g159) & (sk[30]) & (g154) & (!g849) & (g881)) + ((g159) & (sk[30]) & (g154) & (g849) & (!g881)) + ((g159) & (sk[30]) & (g154) & (g849) & (g881)));
	assign g897 = (((!g3) & (!g383) & (!g460) & (!g895) & (sk[31]) & (g1478)) + ((!g3) & (!g383) & (g460) & (!g895) & (!sk[31]) & (g1478)) + ((!g3) & (!g383) & (g460) & (!g895) & (sk[31]) & (g1478)) + ((!g3) & (!g383) & (g460) & (g895) & (!sk[31]) & (!g1478)) + ((!g3) & (!g383) & (g460) & (g895) & (!sk[31]) & (g1478)) + ((!g3) & (g383) & (!g460) & (!g895) & (!sk[31]) & (!g1478)) + ((!g3) & (g383) & (!g460) & (!g895) & (!sk[31]) & (g1478)) + ((!g3) & (g383) & (!g460) & (!g895) & (sk[31]) & (g1478)) + ((!g3) & (g383) & (!g460) & (g895) & (!sk[31]) & (!g1478)) + ((!g3) & (g383) & (!g460) & (g895) & (!sk[31]) & (g1478)) + ((!g3) & (g383) & (g460) & (!g895) & (!sk[31]) & (!g1478)) + ((!g3) & (g383) & (g460) & (!g895) & (!sk[31]) & (g1478)) + ((!g3) & (g383) & (g460) & (!g895) & (sk[31]) & (g1478)) + ((!g3) & (g383) & (g460) & (g895) & (!sk[31]) & (!g1478)) + ((!g3) & (g383) & (g460) & (g895) & (!sk[31]) & (g1478)) + ((g3) & (!g383) & (g460) & (!g895) & (!sk[31]) & (g1478)) + ((g3) & (!g383) & (g460) & (!g895) & (sk[31]) & (g1478)) + ((g3) & (!g383) & (g460) & (g895) & (!sk[31]) & (!g1478)) + ((g3) & (!g383) & (g460) & (g895) & (!sk[31]) & (g1478)) + ((g3) & (g383) & (!g460) & (!g895) & (!sk[31]) & (!g1478)) + ((g3) & (g383) & (!g460) & (!g895) & (!sk[31]) & (g1478)) + ((g3) & (g383) & (!g460) & (!g895) & (sk[31]) & (g1478)) + ((g3) & (g383) & (!g460) & (g895) & (!sk[31]) & (!g1478)) + ((g3) & (g383) & (!g460) & (g895) & (!sk[31]) & (g1478)) + ((g3) & (g383) & (g460) & (!g895) & (!sk[31]) & (!g1478)) + ((g3) & (g383) & (g460) & (!g895) & (!sk[31]) & (g1478)) + ((g3) & (g383) & (g460) & (!g895) & (sk[31]) & (g1478)) + ((g3) & (g383) & (g460) & (g895) & (!sk[31]) & (!g1478)) + ((g3) & (g383) & (g460) & (g895) & (!sk[31]) & (g1478)));
	assign g898 = (((!g4) & (sk[32]) & (!g83)) + ((!g4) & (sk[32]) & (g83)) + ((g4) & (!sk[32]) & (!g83)) + ((g4) & (!sk[32]) & (g83)) + ((g4) & (sk[32]) & (!g83)));
	assign g899 = (((!g31) & (!sk[33]) & (!g528) & (g898)) + ((!g31) & (!sk[33]) & (g528) & (!g898)) + ((!g31) & (!sk[33]) & (g528) & (g898)) + ((!g31) & (sk[33]) & (!g528) & (g898)) + ((g31) & (!sk[33]) & (!g528) & (g898)) + ((g31) & (!sk[33]) & (g528) & (!g898)) + ((g31) & (!sk[33]) & (g528) & (g898)));
	assign g900 = (((!g107) & (!g165) & (!sk[34]) & (g460)) + ((!g107) & (g165) & (!sk[34]) & (!g460)) + ((!g107) & (g165) & (!sk[34]) & (g460)) + ((!g107) & (g165) & (sk[34]) & (!g460)) + ((g107) & (!g165) & (!sk[34]) & (g460)) + ((g107) & (g165) & (!sk[34]) & (!g460)) + ((g107) & (g165) & (!sk[34]) & (g460)));
	assign g901 = (((!g142) & (!g392) & (!g351) & (!g496) & (g899) & (!g900)) + ((!g142) & (!g392) & (!g351) & (g496) & (g899) & (!g900)) + ((!g142) & (!g392) & (g351) & (!g496) & (g899) & (!g900)) + ((!g142) & (!g392) & (g351) & (g496) & (g899) & (!g900)) + ((!g142) & (g392) & (!g351) & (!g496) & (g899) & (!g900)) + ((!g142) & (g392) & (g351) & (!g496) & (g899) & (!g900)) + ((g142) & (!g392) & (!g351) & (!g496) & (g899) & (!g900)) + ((g142) & (!g392) & (!g351) & (g496) & (g899) & (!g900)) + ((g142) & (!g392) & (g351) & (!g496) & (!g899) & (!g900)) + ((g142) & (!g392) & (g351) & (!g496) & (g899) & (!g900)) + ((g142) & (!g392) & (g351) & (g496) & (!g899) & (!g900)) + ((g142) & (!g392) & (g351) & (g496) & (g899) & (!g900)) + ((g142) & (g392) & (!g351) & (!g496) & (g899) & (!g900)) + ((g142) & (g392) & (g351) & (!g496) & (!g899) & (!g900)) + ((g142) & (g392) & (g351) & (!g496) & (g899) & (!g900)));
	assign g902 = (((!sk[36]) & (!g73) & (!g144) & (g102) & (!g165) & (g130)) + ((!sk[36]) & (!g73) & (!g144) & (g102) & (g165) & (!g130)) + ((!sk[36]) & (!g73) & (!g144) & (g102) & (g165) & (g130)) + ((!sk[36]) & (!g73) & (g144) & (!g102) & (!g165) & (!g130)) + ((!sk[36]) & (!g73) & (g144) & (!g102) & (!g165) & (g130)) + ((!sk[36]) & (!g73) & (g144) & (!g102) & (g165) & (!g130)) + ((!sk[36]) & (!g73) & (g144) & (!g102) & (g165) & (g130)) + ((!sk[36]) & (!g73) & (g144) & (g102) & (!g165) & (!g130)) + ((!sk[36]) & (!g73) & (g144) & (g102) & (!g165) & (g130)) + ((!sk[36]) & (!g73) & (g144) & (g102) & (g165) & (!g130)) + ((!sk[36]) & (!g73) & (g144) & (g102) & (g165) & (g130)) + ((!sk[36]) & (g73) & (!g144) & (g102) & (!g165) & (g130)) + ((!sk[36]) & (g73) & (!g144) & (g102) & (g165) & (!g130)) + ((!sk[36]) & (g73) & (!g144) & (g102) & (g165) & (g130)) + ((!sk[36]) & (g73) & (g144) & (!g102) & (!g165) & (!g130)) + ((!sk[36]) & (g73) & (g144) & (!g102) & (!g165) & (g130)) + ((!sk[36]) & (g73) & (g144) & (!g102) & (g165) & (!g130)) + ((!sk[36]) & (g73) & (g144) & (!g102) & (g165) & (g130)) + ((!sk[36]) & (g73) & (g144) & (g102) & (!g165) & (!g130)) + ((!sk[36]) & (g73) & (g144) & (g102) & (!g165) & (g130)) + ((!sk[36]) & (g73) & (g144) & (g102) & (g165) & (!g130)) + ((!sk[36]) & (g73) & (g144) & (g102) & (g165) & (g130)) + ((sk[36]) & (!g73) & (!g144) & (!g102) & (!g165) & (g130)));
	assign g903 = (((!i_9_) & (i_10_) & (!i_11_) & (i_15_) & (g4) & (!g24)) + ((!i_9_) & (i_10_) & (!i_11_) & (i_15_) & (g4) & (g24)) + ((i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (!g4) & (!g24)) + ((i_9_) & (i_10_) & (!i_11_) & (!i_15_) & (g4) & (!g24)) + ((i_9_) & (i_10_) & (!i_11_) & (i_15_) & (g4) & (!g24)) + ((i_9_) & (i_10_) & (!i_11_) & (i_15_) & (g4) & (g24)) + ((i_9_) & (i_10_) & (i_11_) & (!i_15_) & (!g4) & (!g24)) + ((i_9_) & (i_10_) & (i_11_) & (!i_15_) & (g4) & (!g24)) + ((i_9_) & (i_10_) & (i_11_) & (i_15_) & (g4) & (!g24)) + ((i_9_) & (i_10_) & (i_11_) & (i_15_) & (g4) & (g24)));
	assign g904 = (((!g45) & (!g86) & (!sk[38]) & (g460)) + ((!g45) & (g86) & (!sk[38]) & (!g460)) + ((!g45) & (g86) & (!sk[38]) & (g460)) + ((g45) & (!g86) & (!sk[38]) & (g460)) + ((g45) & (g86) & (!sk[38]) & (!g460)) + ((g45) & (g86) & (!sk[38]) & (g460)) + ((g45) & (g86) & (sk[38]) & (!g460)));
	assign g905 = (((!sk[39]) & (!i_8_) & (!g42) & (g72) & (!g473) & (g904)) + ((!sk[39]) & (!i_8_) & (!g42) & (g72) & (g473) & (!g904)) + ((!sk[39]) & (!i_8_) & (!g42) & (g72) & (g473) & (g904)) + ((!sk[39]) & (!i_8_) & (g42) & (!g72) & (!g473) & (!g904)) + ((!sk[39]) & (!i_8_) & (g42) & (!g72) & (!g473) & (g904)) + ((!sk[39]) & (!i_8_) & (g42) & (!g72) & (g473) & (!g904)) + ((!sk[39]) & (!i_8_) & (g42) & (!g72) & (g473) & (g904)) + ((!sk[39]) & (!i_8_) & (g42) & (g72) & (!g473) & (!g904)) + ((!sk[39]) & (!i_8_) & (g42) & (g72) & (!g473) & (g904)) + ((!sk[39]) & (!i_8_) & (g42) & (g72) & (g473) & (!g904)) + ((!sk[39]) & (!i_8_) & (g42) & (g72) & (g473) & (g904)) + ((!sk[39]) & (i_8_) & (!g42) & (g72) & (!g473) & (g904)) + ((!sk[39]) & (i_8_) & (!g42) & (g72) & (g473) & (!g904)) + ((!sk[39]) & (i_8_) & (!g42) & (g72) & (g473) & (g904)) + ((!sk[39]) & (i_8_) & (g42) & (!g72) & (!g473) & (!g904)) + ((!sk[39]) & (i_8_) & (g42) & (!g72) & (!g473) & (g904)) + ((!sk[39]) & (i_8_) & (g42) & (!g72) & (g473) & (!g904)) + ((!sk[39]) & (i_8_) & (g42) & (!g72) & (g473) & (g904)) + ((!sk[39]) & (i_8_) & (g42) & (g72) & (!g473) & (!g904)) + ((!sk[39]) & (i_8_) & (g42) & (g72) & (!g473) & (g904)) + ((!sk[39]) & (i_8_) & (g42) & (g72) & (g473) & (!g904)) + ((!sk[39]) & (i_8_) & (g42) & (g72) & (g473) & (g904)) + ((sk[39]) & (i_8_) & (!g42) & (g72) & (!g473) & (g904)) + ((sk[39]) & (i_8_) & (g42) & (g72) & (!g473) & (g904)) + ((sk[39]) & (i_8_) & (g42) & (g72) & (g473) & (!g904)) + ((sk[39]) & (i_8_) & (g42) & (g72) & (g473) & (g904)));
	assign g906 = (((!g422) & (!sk[40]) & (!g852) & (g902) & (!g903) & (g905)) + ((!g422) & (!sk[40]) & (!g852) & (g902) & (g903) & (!g905)) + ((!g422) & (!sk[40]) & (!g852) & (g902) & (g903) & (g905)) + ((!g422) & (!sk[40]) & (g852) & (!g902) & (!g903) & (!g905)) + ((!g422) & (!sk[40]) & (g852) & (!g902) & (!g903) & (g905)) + ((!g422) & (!sk[40]) & (g852) & (!g902) & (g903) & (!g905)) + ((!g422) & (!sk[40]) & (g852) & (!g902) & (g903) & (g905)) + ((!g422) & (!sk[40]) & (g852) & (g902) & (!g903) & (!g905)) + ((!g422) & (!sk[40]) & (g852) & (g902) & (!g903) & (g905)) + ((!g422) & (!sk[40]) & (g852) & (g902) & (g903) & (!g905)) + ((!g422) & (!sk[40]) & (g852) & (g902) & (g903) & (g905)) + ((!g422) & (sk[40]) & (!g852) & (!g902) & (!g903) & (!g905)) + ((!g422) & (sk[40]) & (!g852) & (!g902) & (g903) & (!g905)) + ((!g422) & (sk[40]) & (!g852) & (g902) & (!g903) & (!g905)) + ((!g422) & (sk[40]) & (!g852) & (g902) & (g903) & (!g905)) + ((!g422) & (sk[40]) & (g852) & (g902) & (!g903) & (!g905)) + ((!g422) & (sk[40]) & (g852) & (g902) & (g903) & (!g905)) + ((g422) & (!sk[40]) & (!g852) & (g902) & (!g903) & (g905)) + ((g422) & (!sk[40]) & (!g852) & (g902) & (g903) & (!g905)) + ((g422) & (!sk[40]) & (!g852) & (g902) & (g903) & (g905)) + ((g422) & (!sk[40]) & (g852) & (!g902) & (!g903) & (!g905)) + ((g422) & (!sk[40]) & (g852) & (!g902) & (!g903) & (g905)) + ((g422) & (!sk[40]) & (g852) & (!g902) & (g903) & (!g905)) + ((g422) & (!sk[40]) & (g852) & (!g902) & (g903) & (g905)) + ((g422) & (!sk[40]) & (g852) & (g902) & (!g903) & (!g905)) + ((g422) & (!sk[40]) & (g852) & (g902) & (!g903) & (g905)) + ((g422) & (!sk[40]) & (g852) & (g902) & (g903) & (!g905)) + ((g422) & (!sk[40]) & (g852) & (g902) & (g903) & (g905)) + ((g422) & (sk[40]) & (!g852) & (!g902) & (!g903) & (!g905)) + ((g422) & (sk[40]) & (!g852) & (g902) & (!g903) & (!g905)) + ((g422) & (sk[40]) & (g852) & (g902) & (!g903) & (!g905)));
	assign g907 = (((!g119) & (!g272) & (!sk[41]) & (g425) & (!g351) & (g468)) + ((!g119) & (!g272) & (!sk[41]) & (g425) & (g351) & (!g468)) + ((!g119) & (!g272) & (!sk[41]) & (g425) & (g351) & (g468)) + ((!g119) & (!g272) & (sk[41]) & (!g425) & (!g351) & (!g468)) + ((!g119) & (!g272) & (sk[41]) & (!g425) & (g351) & (!g468)) + ((!g119) & (!g272) & (sk[41]) & (!g425) & (g351) & (g468)) + ((!g119) & (!g272) & (sk[41]) & (g425) & (!g351) & (!g468)) + ((!g119) & (!g272) & (sk[41]) & (g425) & (g351) & (!g468)) + ((!g119) & (!g272) & (sk[41]) & (g425) & (g351) & (g468)) + ((!g119) & (g272) & (!sk[41]) & (!g425) & (!g351) & (!g468)) + ((!g119) & (g272) & (!sk[41]) & (!g425) & (!g351) & (g468)) + ((!g119) & (g272) & (!sk[41]) & (!g425) & (g351) & (!g468)) + ((!g119) & (g272) & (!sk[41]) & (!g425) & (g351) & (g468)) + ((!g119) & (g272) & (!sk[41]) & (g425) & (!g351) & (!g468)) + ((!g119) & (g272) & (!sk[41]) & (g425) & (!g351) & (g468)) + ((!g119) & (g272) & (!sk[41]) & (g425) & (g351) & (!g468)) + ((!g119) & (g272) & (!sk[41]) & (g425) & (g351) & (g468)) + ((!g119) & (g272) & (sk[41]) & (g425) & (!g351) & (!g468)) + ((!g119) & (g272) & (sk[41]) & (g425) & (g351) & (!g468)) + ((!g119) & (g272) & (sk[41]) & (g425) & (g351) & (g468)) + ((g119) & (!g272) & (!sk[41]) & (g425) & (!g351) & (g468)) + ((g119) & (!g272) & (!sk[41]) & (g425) & (g351) & (!g468)) + ((g119) & (!g272) & (!sk[41]) & (g425) & (g351) & (g468)) + ((g119) & (!g272) & (sk[41]) & (!g425) & (!g351) & (!g468)) + ((g119) & (!g272) & (sk[41]) & (!g425) & (g351) & (!g468)) + ((g119) & (!g272) & (sk[41]) & (g425) & (!g351) & (!g468)) + ((g119) & (!g272) & (sk[41]) & (g425) & (g351) & (!g468)) + ((g119) & (g272) & (!sk[41]) & (!g425) & (!g351) & (!g468)) + ((g119) & (g272) & (!sk[41]) & (!g425) & (!g351) & (g468)) + ((g119) & (g272) & (!sk[41]) & (!g425) & (g351) & (!g468)) + ((g119) & (g272) & (!sk[41]) & (!g425) & (g351) & (g468)) + ((g119) & (g272) & (!sk[41]) & (g425) & (!g351) & (!g468)) + ((g119) & (g272) & (!sk[41]) & (g425) & (!g351) & (g468)) + ((g119) & (g272) & (!sk[41]) & (g425) & (g351) & (!g468)) + ((g119) & (g272) & (!sk[41]) & (g425) & (g351) & (g468)) + ((g119) & (g272) & (sk[41]) & (g425) & (!g351) & (!g468)) + ((g119) & (g272) & (sk[41]) & (g425) & (g351) & (!g468)));
	assign g908 = (((!g887) & (g894) & (g897) & (g901) & (g906) & (g907)));
	assign g909 = (((!i_9_) & (!i_10_) & (i_11_) & (!sk[43]) & (!i_15_) & (g4)) + ((!i_9_) & (!i_10_) & (i_11_) & (!sk[43]) & (i_15_) & (!g4)) + ((!i_9_) & (!i_10_) & (i_11_) & (!sk[43]) & (i_15_) & (g4)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[43]) & (!i_15_) & (!g4)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[43]) & (!i_15_) & (g4)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[43]) & (i_15_) & (!g4)) + ((!i_9_) & (i_10_) & (!i_11_) & (!sk[43]) & (i_15_) & (g4)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[43]) & (!i_15_) & (!g4)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[43]) & (!i_15_) & (g4)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[43]) & (i_15_) & (!g4)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[43]) & (i_15_) & (g4)) + ((!i_9_) & (i_10_) & (i_11_) & (sk[43]) & (!i_15_) & (g4)) + ((i_9_) & (!i_10_) & (!i_11_) & (sk[43]) & (i_15_) & (g4)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[43]) & (!i_15_) & (g4)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[43]) & (i_15_) & (!g4)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[43]) & (i_15_) & (g4)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[43]) & (!i_15_) & (!g4)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[43]) & (!i_15_) & (g4)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[43]) & (i_15_) & (!g4)) + ((i_9_) & (i_10_) & (!i_11_) & (!sk[43]) & (i_15_) & (g4)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[43]) & (!i_15_) & (!g4)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[43]) & (!i_15_) & (g4)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[43]) & (i_15_) & (!g4)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[43]) & (i_15_) & (g4)));
	assign g910 = (((!i_15_) & (!sk[44]) & (!g102) & (g615) & (!g350) & (g909)) + ((!i_15_) & (!sk[44]) & (!g102) & (g615) & (g350) & (!g909)) + ((!i_15_) & (!sk[44]) & (!g102) & (g615) & (g350) & (g909)) + ((!i_15_) & (!sk[44]) & (g102) & (!g615) & (!g350) & (!g909)) + ((!i_15_) & (!sk[44]) & (g102) & (!g615) & (!g350) & (g909)) + ((!i_15_) & (!sk[44]) & (g102) & (!g615) & (g350) & (!g909)) + ((!i_15_) & (!sk[44]) & (g102) & (!g615) & (g350) & (g909)) + ((!i_15_) & (!sk[44]) & (g102) & (g615) & (!g350) & (!g909)) + ((!i_15_) & (!sk[44]) & (g102) & (g615) & (!g350) & (g909)) + ((!i_15_) & (!sk[44]) & (g102) & (g615) & (g350) & (!g909)) + ((!i_15_) & (!sk[44]) & (g102) & (g615) & (g350) & (g909)) + ((!i_15_) & (sk[44]) & (!g102) & (!g615) & (g350) & (g909)) + ((!i_15_) & (sk[44]) & (!g102) & (g615) & (g350) & (g909)) + ((!i_15_) & (sk[44]) & (g102) & (!g615) & (!g350) & (g909)) + ((!i_15_) & (sk[44]) & (g102) & (!g615) & (g350) & (g909)) + ((!i_15_) & (sk[44]) & (g102) & (g615) & (!g350) & (g909)) + ((!i_15_) & (sk[44]) & (g102) & (g615) & (g350) & (g909)) + ((i_15_) & (!sk[44]) & (!g102) & (g615) & (!g350) & (g909)) + ((i_15_) & (!sk[44]) & (!g102) & (g615) & (g350) & (!g909)) + ((i_15_) & (!sk[44]) & (!g102) & (g615) & (g350) & (g909)) + ((i_15_) & (!sk[44]) & (g102) & (!g615) & (!g350) & (!g909)) + ((i_15_) & (!sk[44]) & (g102) & (!g615) & (!g350) & (g909)) + ((i_15_) & (!sk[44]) & (g102) & (!g615) & (g350) & (!g909)) + ((i_15_) & (!sk[44]) & (g102) & (!g615) & (g350) & (g909)) + ((i_15_) & (!sk[44]) & (g102) & (g615) & (!g350) & (!g909)) + ((i_15_) & (!sk[44]) & (g102) & (g615) & (!g350) & (g909)) + ((i_15_) & (!sk[44]) & (g102) & (g615) & (g350) & (!g909)) + ((i_15_) & (!sk[44]) & (g102) & (g615) & (g350) & (g909)) + ((i_15_) & (sk[44]) & (!g102) & (!g615) & (!g350) & (g909)) + ((i_15_) & (sk[44]) & (!g102) & (!g615) & (g350) & (g909)) + ((i_15_) & (sk[44]) & (g102) & (!g615) & (!g350) & (g909)) + ((i_15_) & (sk[44]) & (g102) & (!g615) & (g350) & (g909)));
	assign g911 = (((!i_11_) & (!i_15_) & (g4) & (g34) & (g125) & (!g218)) + ((!i_11_) & (!i_15_) & (g4) & (g34) & (g125) & (g218)) + ((i_11_) & (!i_15_) & (g4) & (g34) & (!g125) & (g218)) + ((i_11_) & (!i_15_) & (g4) & (g34) & (g125) & (g218)));
	assign g912 = (((!i_14_) & (!sk[46]) & (!g27) & (g226)) + ((!i_14_) & (!sk[46]) & (g27) & (!g226)) + ((!i_14_) & (!sk[46]) & (g27) & (g226)) + ((!i_14_) & (sk[46]) & (g27) & (!g226)) + ((i_14_) & (!sk[46]) & (!g27) & (g226)) + ((i_14_) & (!sk[46]) & (g27) & (!g226)) + ((i_14_) & (!sk[46]) & (g27) & (g226)));
	assign g913 = (((!g123) & (!g105) & (!g852) & (sk[47]) & (!g853) & (!g875)) + ((!g123) & (!g105) & (g852) & (!sk[47]) & (!g853) & (g875)) + ((!g123) & (!g105) & (g852) & (!sk[47]) & (g853) & (!g875)) + ((!g123) & (!g105) & (g852) & (!sk[47]) & (g853) & (g875)) + ((!g123) & (g105) & (!g852) & (!sk[47]) & (!g853) & (!g875)) + ((!g123) & (g105) & (!g852) & (!sk[47]) & (!g853) & (g875)) + ((!g123) & (g105) & (!g852) & (!sk[47]) & (g853) & (!g875)) + ((!g123) & (g105) & (!g852) & (!sk[47]) & (g853) & (g875)) + ((!g123) & (g105) & (!g852) & (sk[47]) & (!g853) & (!g875)) + ((!g123) & (g105) & (g852) & (!sk[47]) & (!g853) & (!g875)) + ((!g123) & (g105) & (g852) & (!sk[47]) & (!g853) & (g875)) + ((!g123) & (g105) & (g852) & (!sk[47]) & (g853) & (!g875)) + ((!g123) & (g105) & (g852) & (!sk[47]) & (g853) & (g875)) + ((g123) & (!g105) & (!g852) & (sk[47]) & (!g853) & (!g875)) + ((g123) & (!g105) & (g852) & (!sk[47]) & (!g853) & (g875)) + ((g123) & (!g105) & (g852) & (!sk[47]) & (g853) & (!g875)) + ((g123) & (!g105) & (g852) & (!sk[47]) & (g853) & (g875)) + ((g123) & (!g105) & (g852) & (sk[47]) & (!g853) & (!g875)) + ((g123) & (g105) & (!g852) & (!sk[47]) & (!g853) & (!g875)) + ((g123) & (g105) & (!g852) & (!sk[47]) & (!g853) & (g875)) + ((g123) & (g105) & (!g852) & (!sk[47]) & (g853) & (!g875)) + ((g123) & (g105) & (!g852) & (!sk[47]) & (g853) & (g875)) + ((g123) & (g105) & (!g852) & (sk[47]) & (!g853) & (!g875)) + ((g123) & (g105) & (!g852) & (sk[47]) & (!g853) & (g875)) + ((g123) & (g105) & (!g852) & (sk[47]) & (g853) & (!g875)) + ((g123) & (g105) & (!g852) & (sk[47]) & (g853) & (g875)) + ((g123) & (g105) & (g852) & (!sk[47]) & (!g853) & (!g875)) + ((g123) & (g105) & (g852) & (!sk[47]) & (!g853) & (g875)) + ((g123) & (g105) & (g852) & (!sk[47]) & (g853) & (!g875)) + ((g123) & (g105) & (g852) & (!sk[47]) & (g853) & (g875)) + ((g123) & (g105) & (g852) & (sk[47]) & (!g853) & (!g875)) + ((g123) & (g105) & (g852) & (sk[47]) & (!g853) & (g875)) + ((g123) & (g105) & (g852) & (sk[47]) & (g853) & (!g875)) + ((g123) & (g105) & (g852) & (sk[47]) & (g853) & (g875)));
	assign g914 = (((!g164) & (!g154) & (!sk[48]) & (g853) & (!g875) & (g913)) + ((!g164) & (!g154) & (!sk[48]) & (g853) & (g875) & (!g913)) + ((!g164) & (!g154) & (!sk[48]) & (g853) & (g875) & (g913)) + ((!g164) & (!g154) & (sk[48]) & (!g853) & (!g875) & (g913)) + ((!g164) & (g154) & (!sk[48]) & (!g853) & (!g875) & (!g913)) + ((!g164) & (g154) & (!sk[48]) & (!g853) & (!g875) & (g913)) + ((!g164) & (g154) & (!sk[48]) & (!g853) & (g875) & (!g913)) + ((!g164) & (g154) & (!sk[48]) & (!g853) & (g875) & (g913)) + ((!g164) & (g154) & (!sk[48]) & (g853) & (!g875) & (!g913)) + ((!g164) & (g154) & (!sk[48]) & (g853) & (!g875) & (g913)) + ((!g164) & (g154) & (!sk[48]) & (g853) & (g875) & (!g913)) + ((!g164) & (g154) & (!sk[48]) & (g853) & (g875) & (g913)) + ((!g164) & (g154) & (sk[48]) & (!g853) & (!g875) & (g913)) + ((!g164) & (g154) & (sk[48]) & (!g853) & (g875) & (g913)) + ((!g164) & (g154) & (sk[48]) & (g853) & (!g875) & (g913)) + ((!g164) & (g154) & (sk[48]) & (g853) & (g875) & (g913)) + ((g164) & (!g154) & (!sk[48]) & (g853) & (!g875) & (g913)) + ((g164) & (!g154) & (!sk[48]) & (g853) & (g875) & (!g913)) + ((g164) & (!g154) & (!sk[48]) & (g853) & (g875) & (g913)) + ((g164) & (!g154) & (sk[48]) & (!g853) & (!g875) & (g913)) + ((g164) & (g154) & (!sk[48]) & (!g853) & (!g875) & (!g913)) + ((g164) & (g154) & (!sk[48]) & (!g853) & (!g875) & (g913)) + ((g164) & (g154) & (!sk[48]) & (!g853) & (g875) & (!g913)) + ((g164) & (g154) & (!sk[48]) & (!g853) & (g875) & (g913)) + ((g164) & (g154) & (!sk[48]) & (g853) & (!g875) & (!g913)) + ((g164) & (g154) & (!sk[48]) & (g853) & (!g875) & (g913)) + ((g164) & (g154) & (!sk[48]) & (g853) & (g875) & (!g913)) + ((g164) & (g154) & (!sk[48]) & (g853) & (g875) & (g913)) + ((g164) & (g154) & (sk[48]) & (!g853) & (!g875) & (g913)));
	assign g915 = (((!sk[49]) & (!g105) & (!g851) & (g911) & (!g912) & (g914)) + ((!sk[49]) & (!g105) & (!g851) & (g911) & (g912) & (!g914)) + ((!sk[49]) & (!g105) & (!g851) & (g911) & (g912) & (g914)) + ((!sk[49]) & (!g105) & (g851) & (!g911) & (!g912) & (!g914)) + ((!sk[49]) & (!g105) & (g851) & (!g911) & (!g912) & (g914)) + ((!sk[49]) & (!g105) & (g851) & (!g911) & (g912) & (!g914)) + ((!sk[49]) & (!g105) & (g851) & (!g911) & (g912) & (g914)) + ((!sk[49]) & (!g105) & (g851) & (g911) & (!g912) & (!g914)) + ((!sk[49]) & (!g105) & (g851) & (g911) & (!g912) & (g914)) + ((!sk[49]) & (!g105) & (g851) & (g911) & (g912) & (!g914)) + ((!sk[49]) & (!g105) & (g851) & (g911) & (g912) & (g914)) + ((!sk[49]) & (g105) & (!g851) & (g911) & (!g912) & (g914)) + ((!sk[49]) & (g105) & (!g851) & (g911) & (g912) & (!g914)) + ((!sk[49]) & (g105) & (!g851) & (g911) & (g912) & (g914)) + ((!sk[49]) & (g105) & (g851) & (!g911) & (!g912) & (!g914)) + ((!sk[49]) & (g105) & (g851) & (!g911) & (!g912) & (g914)) + ((!sk[49]) & (g105) & (g851) & (!g911) & (g912) & (!g914)) + ((!sk[49]) & (g105) & (g851) & (!g911) & (g912) & (g914)) + ((!sk[49]) & (g105) & (g851) & (g911) & (!g912) & (!g914)) + ((!sk[49]) & (g105) & (g851) & (g911) & (!g912) & (g914)) + ((!sk[49]) & (g105) & (g851) & (g911) & (g912) & (!g914)) + ((!sk[49]) & (g105) & (g851) & (g911) & (g912) & (g914)) + ((sk[49]) & (!g105) & (g851) & (!g911) & (!g912) & (g914)) + ((sk[49]) & (g105) & (!g851) & (!g911) & (!g912) & (g914)) + ((sk[49]) & (g105) & (g851) & (!g911) & (!g912) & (g914)));
	assign g916 = (((!g126) & (!g122) & (!g105) & (sk[50]) & (!g383) & (!g460)) + ((!g126) & (!g122) & (!g105) & (sk[50]) & (g383) & (!g460)) + ((!g126) & (!g122) & (g105) & (!sk[50]) & (!g383) & (g460)) + ((!g126) & (!g122) & (g105) & (!sk[50]) & (g383) & (!g460)) + ((!g126) & (!g122) & (g105) & (!sk[50]) & (g383) & (g460)) + ((!g126) & (!g122) & (g105) & (sk[50]) & (!g383) & (!g460)) + ((!g126) & (g122) & (!g105) & (!sk[50]) & (!g383) & (!g460)) + ((!g126) & (g122) & (!g105) & (!sk[50]) & (!g383) & (g460)) + ((!g126) & (g122) & (!g105) & (!sk[50]) & (g383) & (!g460)) + ((!g126) & (g122) & (!g105) & (!sk[50]) & (g383) & (g460)) + ((!g126) & (g122) & (!g105) & (sk[50]) & (!g383) & (!g460)) + ((!g126) & (g122) & (!g105) & (sk[50]) & (g383) & (!g460)) + ((!g126) & (g122) & (g105) & (!sk[50]) & (!g383) & (!g460)) + ((!g126) & (g122) & (g105) & (!sk[50]) & (!g383) & (g460)) + ((!g126) & (g122) & (g105) & (!sk[50]) & (g383) & (!g460)) + ((!g126) & (g122) & (g105) & (!sk[50]) & (g383) & (g460)) + ((!g126) & (g122) & (g105) & (sk[50]) & (!g383) & (!g460)) + ((!g126) & (g122) & (g105) & (sk[50]) & (g383) & (!g460)) + ((g126) & (!g122) & (g105) & (!sk[50]) & (!g383) & (g460)) + ((g126) & (!g122) & (g105) & (!sk[50]) & (g383) & (!g460)) + ((g126) & (!g122) & (g105) & (!sk[50]) & (g383) & (g460)) + ((g126) & (g122) & (!g105) & (!sk[50]) & (!g383) & (!g460)) + ((g126) & (g122) & (!g105) & (!sk[50]) & (!g383) & (g460)) + ((g126) & (g122) & (!g105) & (!sk[50]) & (g383) & (!g460)) + ((g126) & (g122) & (!g105) & (!sk[50]) & (g383) & (g460)) + ((g126) & (g122) & (g105) & (!sk[50]) & (!g383) & (!g460)) + ((g126) & (g122) & (g105) & (!sk[50]) & (!g383) & (g460)) + ((g126) & (g122) & (g105) & (!sk[50]) & (g383) & (!g460)) + ((g126) & (g122) & (g105) & (!sk[50]) & (g383) & (g460)));
	assign g917 = (((!g24) & (!sk[51]) & (!g83) & (g699)) + ((!g24) & (!sk[51]) & (g83) & (!g699)) + ((!g24) & (!sk[51]) & (g83) & (g699)) + ((!g24) & (sk[51]) & (!g83) & (g699)) + ((g24) & (!sk[51]) & (!g83) & (g699)) + ((g24) & (!sk[51]) & (g83) & (!g699)) + ((g24) & (!sk[51]) & (g83) & (g699)) + ((g24) & (sk[51]) & (!g83) & (g699)) + ((g24) & (sk[51]) & (g83) & (g699)));
	assign g918 = (((!g164) & (!sk[52]) & (!g213) & (g270) & (!g402) & (g654)) + ((!g164) & (!sk[52]) & (!g213) & (g270) & (g402) & (!g654)) + ((!g164) & (!sk[52]) & (!g213) & (g270) & (g402) & (g654)) + ((!g164) & (!sk[52]) & (g213) & (!g270) & (!g402) & (!g654)) + ((!g164) & (!sk[52]) & (g213) & (!g270) & (!g402) & (g654)) + ((!g164) & (!sk[52]) & (g213) & (!g270) & (g402) & (!g654)) + ((!g164) & (!sk[52]) & (g213) & (!g270) & (g402) & (g654)) + ((!g164) & (!sk[52]) & (g213) & (g270) & (!g402) & (!g654)) + ((!g164) & (!sk[52]) & (g213) & (g270) & (!g402) & (g654)) + ((!g164) & (!sk[52]) & (g213) & (g270) & (g402) & (!g654)) + ((!g164) & (!sk[52]) & (g213) & (g270) & (g402) & (g654)) + ((!g164) & (sk[52]) & (!g213) & (!g270) & (!g402) & (!g654)) + ((!g164) & (sk[52]) & (!g213) & (!g270) & (g402) & (!g654)) + ((!g164) & (sk[52]) & (!g213) & (!g270) & (g402) & (g654)) + ((!g164) & (sk[52]) & (!g213) & (g270) & (g402) & (!g654)) + ((!g164) & (sk[52]) & (!g213) & (g270) & (g402) & (g654)) + ((!g164) & (sk[52]) & (g213) & (!g270) & (!g402) & (!g654)) + ((!g164) & (sk[52]) & (g213) & (!g270) & (g402) & (!g654)) + ((g164) & (!sk[52]) & (!g213) & (g270) & (!g402) & (g654)) + ((g164) & (!sk[52]) & (!g213) & (g270) & (g402) & (!g654)) + ((g164) & (!sk[52]) & (!g213) & (g270) & (g402) & (g654)) + ((g164) & (!sk[52]) & (g213) & (!g270) & (!g402) & (!g654)) + ((g164) & (!sk[52]) & (g213) & (!g270) & (!g402) & (g654)) + ((g164) & (!sk[52]) & (g213) & (!g270) & (g402) & (!g654)) + ((g164) & (!sk[52]) & (g213) & (!g270) & (g402) & (g654)) + ((g164) & (!sk[52]) & (g213) & (g270) & (!g402) & (!g654)) + ((g164) & (!sk[52]) & (g213) & (g270) & (!g402) & (g654)) + ((g164) & (!sk[52]) & (g213) & (g270) & (g402) & (!g654)) + ((g164) & (!sk[52]) & (g213) & (g270) & (g402) & (g654)) + ((g164) & (sk[52]) & (!g213) & (!g270) & (!g402) & (!g654)) + ((g164) & (sk[52]) & (!g213) & (!g270) & (g402) & (!g654)) + ((g164) & (sk[52]) & (g213) & (!g270) & (!g402) & (!g654)) + ((g164) & (sk[52]) & (g213) & (!g270) & (g402) & (!g654)));
	assign g919 = (((!i_12_) & (!sk[53]) & (!i_13_) & (i_14_) & (!g27) & (g167)) + ((!i_12_) & (!sk[53]) & (!i_13_) & (i_14_) & (g27) & (!g167)) + ((!i_12_) & (!sk[53]) & (!i_13_) & (i_14_) & (g27) & (g167)) + ((!i_12_) & (!sk[53]) & (i_13_) & (!i_14_) & (!g27) & (!g167)) + ((!i_12_) & (!sk[53]) & (i_13_) & (!i_14_) & (!g27) & (g167)) + ((!i_12_) & (!sk[53]) & (i_13_) & (!i_14_) & (g27) & (!g167)) + ((!i_12_) & (!sk[53]) & (i_13_) & (!i_14_) & (g27) & (g167)) + ((!i_12_) & (!sk[53]) & (i_13_) & (i_14_) & (!g27) & (!g167)) + ((!i_12_) & (!sk[53]) & (i_13_) & (i_14_) & (!g27) & (g167)) + ((!i_12_) & (!sk[53]) & (i_13_) & (i_14_) & (g27) & (!g167)) + ((!i_12_) & (!sk[53]) & (i_13_) & (i_14_) & (g27) & (g167)) + ((!i_12_) & (sk[53]) & (!i_13_) & (!i_14_) & (g27) & (g167)) + ((!i_12_) & (sk[53]) & (!i_13_) & (i_14_) & (g27) & (!g167)) + ((!i_12_) & (sk[53]) & (!i_13_) & (i_14_) & (g27) & (g167)) + ((i_12_) & (!sk[53]) & (!i_13_) & (i_14_) & (!g27) & (g167)) + ((i_12_) & (!sk[53]) & (!i_13_) & (i_14_) & (g27) & (!g167)) + ((i_12_) & (!sk[53]) & (!i_13_) & (i_14_) & (g27) & (g167)) + ((i_12_) & (!sk[53]) & (i_13_) & (!i_14_) & (!g27) & (!g167)) + ((i_12_) & (!sk[53]) & (i_13_) & (!i_14_) & (!g27) & (g167)) + ((i_12_) & (!sk[53]) & (i_13_) & (!i_14_) & (g27) & (!g167)) + ((i_12_) & (!sk[53]) & (i_13_) & (!i_14_) & (g27) & (g167)) + ((i_12_) & (!sk[53]) & (i_13_) & (i_14_) & (!g27) & (!g167)) + ((i_12_) & (!sk[53]) & (i_13_) & (i_14_) & (!g27) & (g167)) + ((i_12_) & (!sk[53]) & (i_13_) & (i_14_) & (g27) & (!g167)) + ((i_12_) & (!sk[53]) & (i_13_) & (i_14_) & (g27) & (g167)));
	assign g920 = (((!i_14_) & (!g225) & (!g213) & (sk[54]) & (!g425) & (g919)) + ((!i_14_) & (!g225) & (!g213) & (sk[54]) & (g425) & (g919)) + ((!i_14_) & (!g225) & (g213) & (!sk[54]) & (!g425) & (g919)) + ((!i_14_) & (!g225) & (g213) & (!sk[54]) & (g425) & (!g919)) + ((!i_14_) & (!g225) & (g213) & (!sk[54]) & (g425) & (g919)) + ((!i_14_) & (!g225) & (g213) & (sk[54]) & (!g425) & (g919)) + ((!i_14_) & (!g225) & (g213) & (sk[54]) & (g425) & (g919)) + ((!i_14_) & (g225) & (!g213) & (!sk[54]) & (!g425) & (!g919)) + ((!i_14_) & (g225) & (!g213) & (!sk[54]) & (!g425) & (g919)) + ((!i_14_) & (g225) & (!g213) & (!sk[54]) & (g425) & (!g919)) + ((!i_14_) & (g225) & (!g213) & (!sk[54]) & (g425) & (g919)) + ((!i_14_) & (g225) & (!g213) & (sk[54]) & (!g425) & (g919)) + ((!i_14_) & (g225) & (!g213) & (sk[54]) & (g425) & (g919)) + ((!i_14_) & (g225) & (g213) & (!sk[54]) & (!g425) & (!g919)) + ((!i_14_) & (g225) & (g213) & (!sk[54]) & (!g425) & (g919)) + ((!i_14_) & (g225) & (g213) & (!sk[54]) & (g425) & (!g919)) + ((!i_14_) & (g225) & (g213) & (!sk[54]) & (g425) & (g919)) + ((!i_14_) & (g225) & (g213) & (sk[54]) & (!g425) & (g919)) + ((!i_14_) & (g225) & (g213) & (sk[54]) & (g425) & (g919)) + ((i_14_) & (!g225) & (!g213) & (sk[54]) & (!g425) & (g919)) + ((i_14_) & (!g225) & (g213) & (!sk[54]) & (!g425) & (g919)) + ((i_14_) & (!g225) & (g213) & (!sk[54]) & (g425) & (!g919)) + ((i_14_) & (!g225) & (g213) & (!sk[54]) & (g425) & (g919)) + ((i_14_) & (!g225) & (g213) & (sk[54]) & (!g425) & (g919)) + ((i_14_) & (!g225) & (g213) & (sk[54]) & (g425) & (g919)) + ((i_14_) & (g225) & (!g213) & (!sk[54]) & (!g425) & (!g919)) + ((i_14_) & (g225) & (!g213) & (!sk[54]) & (!g425) & (g919)) + ((i_14_) & (g225) & (!g213) & (!sk[54]) & (g425) & (!g919)) + ((i_14_) & (g225) & (!g213) & (!sk[54]) & (g425) & (g919)) + ((i_14_) & (g225) & (!g213) & (sk[54]) & (!g425) & (g919)) + ((i_14_) & (g225) & (!g213) & (sk[54]) & (g425) & (g919)) + ((i_14_) & (g225) & (g213) & (!sk[54]) & (!g425) & (!g919)) + ((i_14_) & (g225) & (g213) & (!sk[54]) & (!g425) & (g919)) + ((i_14_) & (g225) & (g213) & (!sk[54]) & (g425) & (!g919)) + ((i_14_) & (g225) & (g213) & (!sk[54]) & (g425) & (g919)) + ((i_14_) & (g225) & (g213) & (sk[54]) & (!g425) & (g919)) + ((i_14_) & (g225) & (g213) & (sk[54]) & (g425) & (g919)));
	assign g921 = (((!g435) & (!g916) & (!sk[55]) & (g917) & (!g918) & (g920)) + ((!g435) & (!g916) & (!sk[55]) & (g917) & (g918) & (!g920)) + ((!g435) & (!g916) & (!sk[55]) & (g917) & (g918) & (g920)) + ((!g435) & (!g916) & (sk[55]) & (g917) & (g918) & (!g920)) + ((!g435) & (g916) & (!sk[55]) & (!g917) & (!g918) & (!g920)) + ((!g435) & (g916) & (!sk[55]) & (!g917) & (!g918) & (g920)) + ((!g435) & (g916) & (!sk[55]) & (!g917) & (g918) & (!g920)) + ((!g435) & (g916) & (!sk[55]) & (!g917) & (g918) & (g920)) + ((!g435) & (g916) & (!sk[55]) & (g917) & (!g918) & (!g920)) + ((!g435) & (g916) & (!sk[55]) & (g917) & (!g918) & (g920)) + ((!g435) & (g916) & (!sk[55]) & (g917) & (g918) & (!g920)) + ((!g435) & (g916) & (!sk[55]) & (g917) & (g918) & (g920)) + ((g435) & (!g916) & (!sk[55]) & (g917) & (!g918) & (g920)) + ((g435) & (!g916) & (!sk[55]) & (g917) & (g918) & (!g920)) + ((g435) & (!g916) & (!sk[55]) & (g917) & (g918) & (g920)) + ((g435) & (!g916) & (sk[55]) & (!g917) & (g918) & (!g920)) + ((g435) & (!g916) & (sk[55]) & (g917) & (g918) & (!g920)) + ((g435) & (g916) & (!sk[55]) & (!g917) & (!g918) & (!g920)) + ((g435) & (g916) & (!sk[55]) & (!g917) & (!g918) & (g920)) + ((g435) & (g916) & (!sk[55]) & (!g917) & (g918) & (!g920)) + ((g435) & (g916) & (!sk[55]) & (!g917) & (g918) & (g920)) + ((g435) & (g916) & (!sk[55]) & (g917) & (!g918) & (!g920)) + ((g435) & (g916) & (!sk[55]) & (g917) & (!g918) & (g920)) + ((g435) & (g916) & (!sk[55]) & (g917) & (g918) & (!g920)) + ((g435) & (g916) & (!sk[55]) & (g917) & (g918) & (g920)));
	assign g922 = (((!g5) & (!g539) & (!g910) & (g915) & (sk[56]) & (g921)) + ((!g5) & (!g539) & (g910) & (!g915) & (!sk[56]) & (g921)) + ((!g5) & (!g539) & (g910) & (g915) & (!sk[56]) & (!g921)) + ((!g5) & (!g539) & (g910) & (g915) & (!sk[56]) & (g921)) + ((!g5) & (g539) & (!g910) & (!g915) & (!sk[56]) & (!g921)) + ((!g5) & (g539) & (!g910) & (!g915) & (!sk[56]) & (g921)) + ((!g5) & (g539) & (!g910) & (g915) & (!sk[56]) & (!g921)) + ((!g5) & (g539) & (!g910) & (g915) & (!sk[56]) & (g921)) + ((!g5) & (g539) & (!g910) & (g915) & (sk[56]) & (g921)) + ((!g5) & (g539) & (g910) & (!g915) & (!sk[56]) & (!g921)) + ((!g5) & (g539) & (g910) & (!g915) & (!sk[56]) & (g921)) + ((!g5) & (g539) & (g910) & (g915) & (!sk[56]) & (!g921)) + ((!g5) & (g539) & (g910) & (g915) & (!sk[56]) & (g921)) + ((g5) & (!g539) & (g910) & (!g915) & (!sk[56]) & (g921)) + ((g5) & (!g539) & (g910) & (g915) & (!sk[56]) & (!g921)) + ((g5) & (!g539) & (g910) & (g915) & (!sk[56]) & (g921)) + ((g5) & (g539) & (!g910) & (!g915) & (!sk[56]) & (!g921)) + ((g5) & (g539) & (!g910) & (!g915) & (!sk[56]) & (g921)) + ((g5) & (g539) & (!g910) & (g915) & (!sk[56]) & (!g921)) + ((g5) & (g539) & (!g910) & (g915) & (!sk[56]) & (g921)) + ((g5) & (g539) & (!g910) & (g915) & (sk[56]) & (g921)) + ((g5) & (g539) & (g910) & (!g915) & (!sk[56]) & (!g921)) + ((g5) & (g539) & (g910) & (!g915) & (!sk[56]) & (g921)) + ((g5) & (g539) & (g910) & (g915) & (!sk[56]) & (!g921)) + ((g5) & (g539) & (g910) & (g915) & (!sk[56]) & (g921)));
	assign g923 = (((g332) & (g823) & (g873) & (g886) & (g908) & (g922)));
	assign g924 = (((!sk[58]) & (i_11_) & (!g34)) + ((!sk[58]) & (i_11_) & (g34)) + ((sk[58]) & (!i_11_) & (g34)));
	assign g925 = (((!sk[59]) & (!g102) & (!g337) & (g605) & (!g635) & (g851)) + ((!sk[59]) & (!g102) & (!g337) & (g605) & (g635) & (!g851)) + ((!sk[59]) & (!g102) & (!g337) & (g605) & (g635) & (g851)) + ((!sk[59]) & (!g102) & (g337) & (!g605) & (!g635) & (!g851)) + ((!sk[59]) & (!g102) & (g337) & (!g605) & (!g635) & (g851)) + ((!sk[59]) & (!g102) & (g337) & (!g605) & (g635) & (!g851)) + ((!sk[59]) & (!g102) & (g337) & (!g605) & (g635) & (g851)) + ((!sk[59]) & (!g102) & (g337) & (g605) & (!g635) & (!g851)) + ((!sk[59]) & (!g102) & (g337) & (g605) & (!g635) & (g851)) + ((!sk[59]) & (!g102) & (g337) & (g605) & (g635) & (!g851)) + ((!sk[59]) & (!g102) & (g337) & (g605) & (g635) & (g851)) + ((!sk[59]) & (g102) & (!g337) & (g605) & (!g635) & (g851)) + ((!sk[59]) & (g102) & (!g337) & (g605) & (g635) & (!g851)) + ((!sk[59]) & (g102) & (!g337) & (g605) & (g635) & (g851)) + ((!sk[59]) & (g102) & (g337) & (!g605) & (!g635) & (!g851)) + ((!sk[59]) & (g102) & (g337) & (!g605) & (!g635) & (g851)) + ((!sk[59]) & (g102) & (g337) & (!g605) & (g635) & (!g851)) + ((!sk[59]) & (g102) & (g337) & (!g605) & (g635) & (g851)) + ((!sk[59]) & (g102) & (g337) & (g605) & (!g635) & (!g851)) + ((!sk[59]) & (g102) & (g337) & (g605) & (!g635) & (g851)) + ((!sk[59]) & (g102) & (g337) & (g605) & (g635) & (!g851)) + ((!sk[59]) & (g102) & (g337) & (g605) & (g635) & (g851)) + ((sk[59]) & (g102) & (!g337) & (!g605) & (!g635) & (!g851)) + ((sk[59]) & (g102) & (!g337) & (!g605) & (g635) & (!g851)) + ((sk[59]) & (g102) & (!g337) & (!g605) & (g635) & (g851)) + ((sk[59]) & (g102) & (!g337) & (g605) & (!g635) & (!g851)) + ((sk[59]) & (g102) & (!g337) & (g605) & (!g635) & (g851)) + ((sk[59]) & (g102) & (!g337) & (g605) & (g635) & (!g851)) + ((sk[59]) & (g102) & (!g337) & (g605) & (g635) & (g851)) + ((sk[59]) & (g102) & (g337) & (!g605) & (!g635) & (!g851)) + ((sk[59]) & (g102) & (g337) & (!g605) & (!g635) & (g851)) + ((sk[59]) & (g102) & (g337) & (!g605) & (g635) & (!g851)) + ((sk[59]) & (g102) & (g337) & (!g605) & (g635) & (g851)) + ((sk[59]) & (g102) & (g337) & (g605) & (!g635) & (!g851)) + ((sk[59]) & (g102) & (g337) & (g605) & (!g635) & (g851)) + ((sk[59]) & (g102) & (g337) & (g605) & (g635) & (!g851)) + ((sk[59]) & (g102) & (g337) & (g605) & (g635) & (g851)));
	assign g926 = (((!g43) & (!g924) & (!g394) & (sk[60]) & (!g925)) + ((!g43) & (!g924) & (g394) & (!sk[60]) & (!g925)) + ((!g43) & (!g924) & (g394) & (!sk[60]) & (g925)) + ((!g43) & (!g924) & (g394) & (sk[60]) & (!g925)) + ((!g43) & (g924) & (!g394) & (sk[60]) & (!g925)) + ((!g43) & (g924) & (g394) & (!sk[60]) & (!g925)) + ((!g43) & (g924) & (g394) & (!sk[60]) & (g925)) + ((!g43) & (g924) & (g394) & (sk[60]) & (!g925)) + ((g43) & (!g924) & (!g394) & (sk[60]) & (!g925)) + ((g43) & (!g924) & (g394) & (!sk[60]) & (!g925)) + ((g43) & (!g924) & (g394) & (!sk[60]) & (g925)) + ((g43) & (!g924) & (g394) & (sk[60]) & (!g925)) + ((g43) & (g924) & (!g394) & (sk[60]) & (!g925)) + ((g43) & (g924) & (g394) & (!sk[60]) & (!g925)) + ((g43) & (g924) & (g394) & (!sk[60]) & (g925)));
	assign g927 = (((!g3) & (!i_12_) & (i_13_) & (!i_14_) & (!sk[61]) & (g69)) + ((!g3) & (!i_12_) & (i_13_) & (!i_14_) & (sk[61]) & (g69)) + ((!g3) & (!i_12_) & (i_13_) & (i_14_) & (!sk[61]) & (!g69)) + ((!g3) & (!i_12_) & (i_13_) & (i_14_) & (!sk[61]) & (g69)) + ((!g3) & (i_12_) & (!i_13_) & (!i_14_) & (!sk[61]) & (!g69)) + ((!g3) & (i_12_) & (!i_13_) & (!i_14_) & (!sk[61]) & (g69)) + ((!g3) & (i_12_) & (!i_13_) & (i_14_) & (!sk[61]) & (!g69)) + ((!g3) & (i_12_) & (!i_13_) & (i_14_) & (!sk[61]) & (g69)) + ((!g3) & (i_12_) & (i_13_) & (!i_14_) & (!sk[61]) & (!g69)) + ((!g3) & (i_12_) & (i_13_) & (!i_14_) & (!sk[61]) & (g69)) + ((!g3) & (i_12_) & (i_13_) & (i_14_) & (!sk[61]) & (!g69)) + ((!g3) & (i_12_) & (i_13_) & (i_14_) & (!sk[61]) & (g69)) + ((!g3) & (i_12_) & (i_13_) & (i_14_) & (sk[61]) & (g69)) + ((g3) & (!i_12_) & (!i_13_) & (!i_14_) & (sk[61]) & (!g69)) + ((g3) & (!i_12_) & (!i_13_) & (!i_14_) & (sk[61]) & (g69)) + ((g3) & (!i_12_) & (i_13_) & (!i_14_) & (!sk[61]) & (g69)) + ((g3) & (!i_12_) & (i_13_) & (!i_14_) & (sk[61]) & (g69)) + ((g3) & (!i_12_) & (i_13_) & (i_14_) & (!sk[61]) & (!g69)) + ((g3) & (!i_12_) & (i_13_) & (i_14_) & (!sk[61]) & (g69)) + ((g3) & (i_12_) & (!i_13_) & (!i_14_) & (!sk[61]) & (!g69)) + ((g3) & (i_12_) & (!i_13_) & (!i_14_) & (!sk[61]) & (g69)) + ((g3) & (i_12_) & (!i_13_) & (i_14_) & (!sk[61]) & (!g69)) + ((g3) & (i_12_) & (!i_13_) & (i_14_) & (!sk[61]) & (g69)) + ((g3) & (i_12_) & (!i_13_) & (i_14_) & (sk[61]) & (!g69)) + ((g3) & (i_12_) & (!i_13_) & (i_14_) & (sk[61]) & (g69)) + ((g3) & (i_12_) & (i_13_) & (!i_14_) & (!sk[61]) & (!g69)) + ((g3) & (i_12_) & (i_13_) & (!i_14_) & (!sk[61]) & (g69)) + ((g3) & (i_12_) & (i_13_) & (i_14_) & (!sk[61]) & (!g69)) + ((g3) & (i_12_) & (i_13_) & (i_14_) & (!sk[61]) & (g69)) + ((g3) & (i_12_) & (i_13_) & (i_14_) & (sk[61]) & (g69)));
	assign g928 = (((!sk[62]) & (!g17) & (!g81) & (g174) & (!g927)) + ((!sk[62]) & (!g17) & (!g81) & (g174) & (g927)) + ((!sk[62]) & (!g17) & (g81) & (g174) & (!g927)) + ((!sk[62]) & (!g17) & (g81) & (g174) & (g927)) + ((!sk[62]) & (g17) & (!g81) & (g174) & (!g927)) + ((!sk[62]) & (g17) & (!g81) & (g174) & (g927)) + ((!sk[62]) & (g17) & (g81) & (g174) & (!g927)) + ((!sk[62]) & (g17) & (g81) & (g174) & (g927)) + ((sk[62]) & (!g17) & (!g81) & (!g174) & (!g927)) + ((sk[62]) & (!g17) & (!g81) & (g174) & (!g927)) + ((sk[62]) & (!g17) & (g81) & (g174) & (!g927)) + ((sk[62]) & (g17) & (!g81) & (g174) & (!g927)) + ((sk[62]) & (g17) & (g81) & (g174) & (!g927)));
	assign g929 = (((!g4) & (!g27) & (!sk[63]) & (g928)) + ((!g4) & (!g27) & (sk[63]) & (g928)) + ((!g4) & (g27) & (!sk[63]) & (!g928)) + ((!g4) & (g27) & (!sk[63]) & (g928)) + ((!g4) & (g27) & (sk[63]) & (g928)) + ((g4) & (!g27) & (!sk[63]) & (g928)) + ((g4) & (!g27) & (sk[63]) & (g928)) + ((g4) & (g27) & (!sk[63]) & (!g928)) + ((g4) & (g27) & (!sk[63]) & (g928)));
	assign g930 = (((!g892) & (sk[64]) & (!g473)) + ((g892) & (!sk[64]) & (!g473)) + ((g892) & (!sk[64]) & (g473)));
	assign g931 = (((!sk[65]) & (!i_15_) & (!g428) & (g24) & (!g460)) + ((!sk[65]) & (!i_15_) & (!g428) & (g24) & (g460)) + ((!sk[65]) & (!i_15_) & (g428) & (g24) & (!g460)) + ((!sk[65]) & (!i_15_) & (g428) & (g24) & (g460)) + ((!sk[65]) & (i_15_) & (!g428) & (g24) & (!g460)) + ((!sk[65]) & (i_15_) & (!g428) & (g24) & (g460)) + ((!sk[65]) & (i_15_) & (g428) & (g24) & (!g460)) + ((!sk[65]) & (i_15_) & (g428) & (g24) & (g460)) + ((sk[65]) & (!i_15_) & (!g428) & (!g24) & (!g460)) + ((sk[65]) & (!i_15_) & (!g428) & (g24) & (!g460)) + ((sk[65]) & (i_15_) & (!g428) & (!g24) & (!g460)) + ((sk[65]) & (i_15_) & (!g428) & (!g24) & (g460)));
	assign g932 = (((!g468) & (!g743) & (!sk[66]) & (g770) & (!g877)) + ((!g468) & (!g743) & (!sk[66]) & (g770) & (g877)) + ((!g468) & (!g743) & (sk[66]) & (!g770) & (!g877)) + ((!g468) & (g743) & (!sk[66]) & (g770) & (!g877)) + ((!g468) & (g743) & (!sk[66]) & (g770) & (g877)) + ((g468) & (!g743) & (!sk[66]) & (g770) & (!g877)) + ((g468) & (!g743) & (!sk[66]) & (g770) & (g877)) + ((g468) & (g743) & (!sk[66]) & (g770) & (!g877)) + ((g468) & (g743) & (!sk[66]) & (g770) & (g877)));
	assign g933 = (((!sk[67]) & (!g929) & (!g930) & (g931) & (!g932)) + ((!sk[67]) & (!g929) & (!g930) & (g931) & (g932)) + ((!sk[67]) & (!g929) & (g930) & (g931) & (!g932)) + ((!sk[67]) & (!g929) & (g930) & (g931) & (g932)) + ((!sk[67]) & (g929) & (!g930) & (g931) & (!g932)) + ((!sk[67]) & (g929) & (!g930) & (g931) & (g932)) + ((!sk[67]) & (g929) & (g930) & (g931) & (!g932)) + ((!sk[67]) & (g929) & (g930) & (g931) & (g932)) + ((sk[67]) & (g929) & (g930) & (!g931) & (g932)));
	assign g934 = (((!g342) & (!g522) & (!sk[68]) & (g630)) + ((!g342) & (!g522) & (sk[68]) & (!g630)) + ((!g342) & (g522) & (!sk[68]) & (!g630)) + ((!g342) & (g522) & (!sk[68]) & (g630)) + ((g342) & (!g522) & (!sk[68]) & (g630)) + ((g342) & (g522) & (!sk[68]) & (!g630)) + ((g342) & (g522) & (!sk[68]) & (g630)));
	assign g935 = (((!g21) & (!g397) & (!g508) & (sk[69]) & (g934)) + ((!g21) & (!g397) & (g508) & (!sk[69]) & (!g934)) + ((!g21) & (!g397) & (g508) & (!sk[69]) & (g934)) + ((!g21) & (g397) & (g508) & (!sk[69]) & (!g934)) + ((!g21) & (g397) & (g508) & (!sk[69]) & (g934)) + ((g21) & (!g397) & (g508) & (!sk[69]) & (!g934)) + ((g21) & (!g397) & (g508) & (!sk[69]) & (g934)) + ((g21) & (g397) & (g508) & (!sk[69]) & (!g934)) + ((g21) & (g397) & (g508) & (!sk[69]) & (g934)));
	assign g936 = (((!i_8_) & (g168) & (!g898) & (!g928) & (!g933) & (!g935)) + ((!i_8_) & (g168) & (!g898) & (!g928) & (!g933) & (g935)) + ((!i_8_) & (g168) & (!g898) & (!g928) & (g933) & (!g935)) + ((!i_8_) & (g168) & (!g898) & (!g928) & (g933) & (g935)) + ((!i_8_) & (g168) & (!g898) & (g928) & (!g933) & (!g935)) + ((!i_8_) & (g168) & (!g898) & (g928) & (!g933) & (g935)) + ((!i_8_) & (g168) & (!g898) & (g928) & (g933) & (!g935)) + ((!i_8_) & (g168) & (!g898) & (g928) & (g933) & (g935)) + ((!i_8_) & (g168) & (g898) & (!g928) & (!g933) & (!g935)) + ((!i_8_) & (g168) & (g898) & (!g928) & (!g933) & (g935)) + ((!i_8_) & (g168) & (g898) & (!g928) & (g933) & (!g935)) + ((!i_8_) & (g168) & (g898) & (g928) & (!g933) & (!g935)) + ((!i_8_) & (g168) & (g898) & (g928) & (!g933) & (g935)) + ((!i_8_) & (g168) & (g898) & (g928) & (g933) & (!g935)) + ((i_8_) & (g168) & (!g898) & (!g928) & (!g933) & (!g935)) + ((i_8_) & (g168) & (!g898) & (!g928) & (!g933) & (g935)) + ((i_8_) & (g168) & (!g898) & (!g928) & (g933) & (!g935)) + ((i_8_) & (g168) & (!g898) & (!g928) & (g933) & (g935)) + ((i_8_) & (g168) & (g898) & (!g928) & (!g933) & (!g935)) + ((i_8_) & (g168) & (g898) & (!g928) & (!g933) & (g935)) + ((i_8_) & (g168) & (g898) & (!g928) & (g933) & (!g935)) + ((i_8_) & (g168) & (g898) & (!g928) & (g933) & (g935)));
	assign g937 = (((!g102) & (!sk[71]) & (!g358) & (g487) & (!g652) & (g852)) + ((!g102) & (!sk[71]) & (!g358) & (g487) & (g652) & (!g852)) + ((!g102) & (!sk[71]) & (!g358) & (g487) & (g652) & (g852)) + ((!g102) & (!sk[71]) & (g358) & (!g487) & (!g652) & (!g852)) + ((!g102) & (!sk[71]) & (g358) & (!g487) & (!g652) & (g852)) + ((!g102) & (!sk[71]) & (g358) & (!g487) & (g652) & (!g852)) + ((!g102) & (!sk[71]) & (g358) & (!g487) & (g652) & (g852)) + ((!g102) & (!sk[71]) & (g358) & (g487) & (!g652) & (!g852)) + ((!g102) & (!sk[71]) & (g358) & (g487) & (!g652) & (g852)) + ((!g102) & (!sk[71]) & (g358) & (g487) & (g652) & (!g852)) + ((!g102) & (!sk[71]) & (g358) & (g487) & (g652) & (g852)) + ((g102) & (!sk[71]) & (!g358) & (g487) & (!g652) & (g852)) + ((g102) & (!sk[71]) & (!g358) & (g487) & (g652) & (!g852)) + ((g102) & (!sk[71]) & (!g358) & (g487) & (g652) & (g852)) + ((g102) & (!sk[71]) & (g358) & (!g487) & (!g652) & (!g852)) + ((g102) & (!sk[71]) & (g358) & (!g487) & (!g652) & (g852)) + ((g102) & (!sk[71]) & (g358) & (!g487) & (g652) & (!g852)) + ((g102) & (!sk[71]) & (g358) & (!g487) & (g652) & (g852)) + ((g102) & (!sk[71]) & (g358) & (g487) & (!g652) & (!g852)) + ((g102) & (!sk[71]) & (g358) & (g487) & (!g652) & (g852)) + ((g102) & (!sk[71]) & (g358) & (g487) & (g652) & (!g852)) + ((g102) & (!sk[71]) & (g358) & (g487) & (g652) & (g852)) + ((g102) & (sk[71]) & (!g358) & (!g487) & (!g652) & (g852)) + ((g102) & (sk[71]) & (!g358) & (!g487) & (g652) & (!g852)) + ((g102) & (sk[71]) & (!g358) & (!g487) & (g652) & (g852)) + ((g102) & (sk[71]) & (!g358) & (g487) & (!g652) & (!g852)) + ((g102) & (sk[71]) & (!g358) & (g487) & (!g652) & (g852)) + ((g102) & (sk[71]) & (!g358) & (g487) & (g652) & (!g852)) + ((g102) & (sk[71]) & (!g358) & (g487) & (g652) & (g852)) + ((g102) & (sk[71]) & (g358) & (!g487) & (!g652) & (!g852)) + ((g102) & (sk[71]) & (g358) & (!g487) & (!g652) & (g852)) + ((g102) & (sk[71]) & (g358) & (!g487) & (g652) & (!g852)) + ((g102) & (sk[71]) & (g358) & (!g487) & (g652) & (g852)) + ((g102) & (sk[71]) & (g358) & (g487) & (!g652) & (!g852)) + ((g102) & (sk[71]) & (g358) & (g487) & (!g652) & (g852)) + ((g102) & (sk[71]) & (g358) & (g487) & (g652) & (!g852)) + ((g102) & (sk[71]) & (g358) & (g487) & (g652) & (g852)));
	assign g938 = (((!g19) & (!g102) & (!sk[72]) & (g113) & (!g105) & (g174)) + ((!g19) & (!g102) & (!sk[72]) & (g113) & (g105) & (!g174)) + ((!g19) & (!g102) & (!sk[72]) & (g113) & (g105) & (g174)) + ((!g19) & (!g102) & (sk[72]) & (!g113) & (!g105) & (!g174)) + ((!g19) & (g102) & (!sk[72]) & (!g113) & (!g105) & (!g174)) + ((!g19) & (g102) & (!sk[72]) & (!g113) & (!g105) & (g174)) + ((!g19) & (g102) & (!sk[72]) & (!g113) & (g105) & (!g174)) + ((!g19) & (g102) & (!sk[72]) & (!g113) & (g105) & (g174)) + ((!g19) & (g102) & (!sk[72]) & (g113) & (!g105) & (!g174)) + ((!g19) & (g102) & (!sk[72]) & (g113) & (!g105) & (g174)) + ((!g19) & (g102) & (!sk[72]) & (g113) & (g105) & (!g174)) + ((!g19) & (g102) & (!sk[72]) & (g113) & (g105) & (g174)) + ((!g19) & (g102) & (sk[72]) & (!g113) & (!g105) & (!g174)) + ((g19) & (!g102) & (!sk[72]) & (g113) & (!g105) & (g174)) + ((g19) & (!g102) & (!sk[72]) & (g113) & (g105) & (!g174)) + ((g19) & (!g102) & (!sk[72]) & (g113) & (g105) & (g174)) + ((g19) & (!g102) & (sk[72]) & (!g113) & (!g105) & (!g174)) + ((g19) & (!g102) & (sk[72]) & (!g113) & (!g105) & (g174)) + ((g19) & (g102) & (!sk[72]) & (!g113) & (!g105) & (!g174)) + ((g19) & (g102) & (!sk[72]) & (!g113) & (!g105) & (g174)) + ((g19) & (g102) & (!sk[72]) & (!g113) & (g105) & (!g174)) + ((g19) & (g102) & (!sk[72]) & (!g113) & (g105) & (g174)) + ((g19) & (g102) & (!sk[72]) & (g113) & (!g105) & (!g174)) + ((g19) & (g102) & (!sk[72]) & (g113) & (!g105) & (g174)) + ((g19) & (g102) & (!sk[72]) & (g113) & (g105) & (!g174)) + ((g19) & (g102) & (!sk[72]) & (g113) & (g105) & (g174)) + ((g19) & (g102) & (sk[72]) & (!g113) & (!g105) & (!g174)) + ((g19) & (g102) & (sk[72]) & (!g113) & (!g105) & (g174)) + ((g19) & (g102) & (sk[72]) & (!g113) & (g105) & (!g174)) + ((g19) & (g102) & (sk[72]) & (!g113) & (g105) & (g174)));
	assign g939 = (((!g4) & (!g126) & (!g102) & (sk[73]) & (!g105) & (!g176)) + ((!g4) & (!g126) & (g102) & (!sk[73]) & (!g105) & (g176)) + ((!g4) & (!g126) & (g102) & (!sk[73]) & (g105) & (!g176)) + ((!g4) & (!g126) & (g102) & (!sk[73]) & (g105) & (g176)) + ((!g4) & (!g126) & (g102) & (sk[73]) & (!g105) & (!g176)) + ((!g4) & (g126) & (!g102) & (!sk[73]) & (!g105) & (!g176)) + ((!g4) & (g126) & (!g102) & (!sk[73]) & (!g105) & (g176)) + ((!g4) & (g126) & (!g102) & (!sk[73]) & (g105) & (!g176)) + ((!g4) & (g126) & (!g102) & (!sk[73]) & (g105) & (g176)) + ((!g4) & (g126) & (g102) & (!sk[73]) & (!g105) & (!g176)) + ((!g4) & (g126) & (g102) & (!sk[73]) & (!g105) & (g176)) + ((!g4) & (g126) & (g102) & (!sk[73]) & (g105) & (!g176)) + ((!g4) & (g126) & (g102) & (!sk[73]) & (g105) & (g176)) + ((g4) & (!g126) & (!g102) & (sk[73]) & (!g105) & (!g176)) + ((g4) & (!g126) & (!g102) & (sk[73]) & (!g105) & (g176)) + ((g4) & (!g126) & (g102) & (!sk[73]) & (!g105) & (g176)) + ((g4) & (!g126) & (g102) & (!sk[73]) & (g105) & (!g176)) + ((g4) & (!g126) & (g102) & (!sk[73]) & (g105) & (g176)) + ((g4) & (!g126) & (g102) & (sk[73]) & (!g105) & (!g176)) + ((g4) & (!g126) & (g102) & (sk[73]) & (!g105) & (g176)) + ((g4) & (!g126) & (g102) & (sk[73]) & (g105) & (!g176)) + ((g4) & (!g126) & (g102) & (sk[73]) & (g105) & (g176)) + ((g4) & (g126) & (!g102) & (!sk[73]) & (!g105) & (!g176)) + ((g4) & (g126) & (!g102) & (!sk[73]) & (!g105) & (g176)) + ((g4) & (g126) & (!g102) & (!sk[73]) & (g105) & (!g176)) + ((g4) & (g126) & (!g102) & (!sk[73]) & (g105) & (g176)) + ((g4) & (g126) & (g102) & (!sk[73]) & (!g105) & (!g176)) + ((g4) & (g126) & (g102) & (!sk[73]) & (!g105) & (g176)) + ((g4) & (g126) & (g102) & (!sk[73]) & (g105) & (!g176)) + ((g4) & (g126) & (g102) & (!sk[73]) & (g105) & (g176)));
	assign g940 = (((!g105) & (!g853) & (!sk[74]) & (g937) & (!g938) & (g939)) + ((!g105) & (!g853) & (!sk[74]) & (g937) & (g938) & (!g939)) + ((!g105) & (!g853) & (!sk[74]) & (g937) & (g938) & (g939)) + ((!g105) & (!g853) & (sk[74]) & (!g937) & (!g938) & (!g939)) + ((!g105) & (g853) & (!sk[74]) & (!g937) & (!g938) & (!g939)) + ((!g105) & (g853) & (!sk[74]) & (!g937) & (!g938) & (g939)) + ((!g105) & (g853) & (!sk[74]) & (!g937) & (g938) & (!g939)) + ((!g105) & (g853) & (!sk[74]) & (!g937) & (g938) & (g939)) + ((!g105) & (g853) & (!sk[74]) & (g937) & (!g938) & (!g939)) + ((!g105) & (g853) & (!sk[74]) & (g937) & (!g938) & (g939)) + ((!g105) & (g853) & (!sk[74]) & (g937) & (g938) & (!g939)) + ((!g105) & (g853) & (!sk[74]) & (g937) & (g938) & (g939)) + ((g105) & (!g853) & (!sk[74]) & (g937) & (!g938) & (g939)) + ((g105) & (!g853) & (!sk[74]) & (g937) & (g938) & (!g939)) + ((g105) & (!g853) & (!sk[74]) & (g937) & (g938) & (g939)) + ((g105) & (!g853) & (sk[74]) & (!g937) & (!g938) & (!g939)) + ((g105) & (g853) & (!sk[74]) & (!g937) & (!g938) & (!g939)) + ((g105) & (g853) & (!sk[74]) & (!g937) & (!g938) & (g939)) + ((g105) & (g853) & (!sk[74]) & (!g937) & (g938) & (!g939)) + ((g105) & (g853) & (!sk[74]) & (!g937) & (g938) & (g939)) + ((g105) & (g853) & (!sk[74]) & (g937) & (!g938) & (!g939)) + ((g105) & (g853) & (!sk[74]) & (g937) & (!g938) & (g939)) + ((g105) & (g853) & (!sk[74]) & (g937) & (g938) & (!g939)) + ((g105) & (g853) & (!sk[74]) & (g937) & (g938) & (g939)) + ((g105) & (g853) & (sk[74]) & (!g937) & (!g938) & (!g939)));
	assign g941 = (((!g102) & (!g105) & (!sk[75]) & (g654) & (!g847)) + ((!g102) & (!g105) & (!sk[75]) & (g654) & (g847)) + ((!g102) & (!g105) & (sk[75]) & (g654) & (!g847)) + ((!g102) & (!g105) & (sk[75]) & (g654) & (g847)) + ((!g102) & (g105) & (!sk[75]) & (g654) & (!g847)) + ((!g102) & (g105) & (!sk[75]) & (g654) & (g847)) + ((g102) & (!g105) & (!sk[75]) & (g654) & (!g847)) + ((g102) & (!g105) & (!sk[75]) & (g654) & (g847)) + ((g102) & (!g105) & (sk[75]) & (!g654) & (!g847)) + ((g102) & (!g105) & (sk[75]) & (g654) & (!g847)) + ((g102) & (!g105) & (sk[75]) & (g654) & (g847)) + ((g102) & (g105) & (!sk[75]) & (g654) & (!g847)) + ((g102) & (g105) & (!sk[75]) & (g654) & (g847)) + ((g102) & (g105) & (sk[75]) & (!g654) & (!g847)) + ((g102) & (g105) & (sk[75]) & (g654) & (!g847)));
	assign g942 = (((!g305) & (!sk[76]) & (!g307) & (g308) & (!g310) & (g941)) + ((!g305) & (!sk[76]) & (!g307) & (g308) & (g310) & (!g941)) + ((!g305) & (!sk[76]) & (!g307) & (g308) & (g310) & (g941)) + ((!g305) & (!sk[76]) & (g307) & (!g308) & (!g310) & (!g941)) + ((!g305) & (!sk[76]) & (g307) & (!g308) & (!g310) & (g941)) + ((!g305) & (!sk[76]) & (g307) & (!g308) & (g310) & (!g941)) + ((!g305) & (!sk[76]) & (g307) & (!g308) & (g310) & (g941)) + ((!g305) & (!sk[76]) & (g307) & (g308) & (!g310) & (!g941)) + ((!g305) & (!sk[76]) & (g307) & (g308) & (!g310) & (g941)) + ((!g305) & (!sk[76]) & (g307) & (g308) & (g310) & (!g941)) + ((!g305) & (!sk[76]) & (g307) & (g308) & (g310) & (g941)) + ((!g305) & (sk[76]) & (!g307) & (!g308) & (!g310) & (!g941)) + ((g305) & (!sk[76]) & (!g307) & (g308) & (!g310) & (g941)) + ((g305) & (!sk[76]) & (!g307) & (g308) & (g310) & (!g941)) + ((g305) & (!sk[76]) & (!g307) & (g308) & (g310) & (g941)) + ((g305) & (!sk[76]) & (g307) & (!g308) & (!g310) & (!g941)) + ((g305) & (!sk[76]) & (g307) & (!g308) & (!g310) & (g941)) + ((g305) & (!sk[76]) & (g307) & (!g308) & (g310) & (!g941)) + ((g305) & (!sk[76]) & (g307) & (!g308) & (g310) & (g941)) + ((g305) & (!sk[76]) & (g307) & (g308) & (!g310) & (!g941)) + ((g305) & (!sk[76]) & (g307) & (g308) & (!g310) & (g941)) + ((g305) & (!sk[76]) & (g307) & (g308) & (g310) & (!g941)) + ((g305) & (!sk[76]) & (g307) & (g308) & (g310) & (g941)));
	assign g943 = (((!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g112) & (!g105)) + ((!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g112) & (!g105)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g112) & (!g105)) + ((!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112) & (!g105)) + ((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112) & (!g105)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g112) & (!g105)) + ((i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (g112) & (!g105)) + ((i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112) & (!g105)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112) & (!g105)));
	assign g944 = (((!g105) & (!g719) & (!sk[78]) & (g943)) + ((!g105) & (g719) & (!sk[78]) & (!g943)) + ((!g105) & (g719) & (!sk[78]) & (g943)) + ((!g105) & (g719) & (sk[78]) & (!g943)) + ((g105) & (!g719) & (!sk[78]) & (g943)) + ((g105) & (!g719) & (sk[78]) & (!g943)) + ((g105) & (g719) & (!sk[78]) & (!g943)) + ((g105) & (g719) & (!sk[78]) & (g943)) + ((g105) & (g719) & (sk[78]) & (!g943)));
	assign g945 = (((!g22) & (!sk[79]) & (!g48) & (g174)) + ((!g22) & (!sk[79]) & (g48) & (!g174)) + ((!g22) & (!sk[79]) & (g48) & (g174)) + ((!g22) & (sk[79]) & (!g48) & (g174)) + ((g22) & (!sk[79]) & (!g48) & (g174)) + ((g22) & (!sk[79]) & (g48) & (!g174)) + ((g22) & (!sk[79]) & (g48) & (g174)) + ((g22) & (sk[79]) & (!g48) & (!g174)) + ((g22) & (sk[79]) & (!g48) & (g174)));
	assign g946 = (((!sk[80]) & (!g105) & (!g188) & (g875)) + ((!sk[80]) & (!g105) & (g188) & (!g875)) + ((!sk[80]) & (!g105) & (g188) & (g875)) + ((!sk[80]) & (g105) & (!g188) & (g875)) + ((!sk[80]) & (g105) & (g188) & (!g875)) + ((!sk[80]) & (g105) & (g188) & (g875)) + ((sk[80]) & (!g105) & (!g188) & (g875)) + ((sk[80]) & (!g105) & (g188) & (!g875)) + ((sk[80]) & (!g105) & (g188) & (g875)));
	assign g947 = (((!g236) & (!g237) & (!g238) & (g240) & (!g241) & (!g946)));
	assign g948 = (((!sk[82]) & (!g337) & (!g605) & (g635)) + ((!sk[82]) & (!g337) & (g605) & (!g635)) + ((!sk[82]) & (!g337) & (g605) & (g635)) + ((!sk[82]) & (g337) & (!g605) & (g635)) + ((!sk[82]) & (g337) & (g605) & (!g635)) + ((!sk[82]) & (g337) & (g605) & (g635)) + ((sk[82]) & (!g337) & (!g605) & (!g635)));
	assign g949 = (((!sk[83]) & (g770) & (!g898)) + ((!sk[83]) & (g770) & (g898)) + ((sk[83]) & (!g770) & (g898)));
	assign g950 = (((!g105) & (!g948) & (!sk[84]) & (g949) & (!g638)) + ((!g105) & (!g948) & (!sk[84]) & (g949) & (g638)) + ((!g105) & (g948) & (!sk[84]) & (g949) & (!g638)) + ((!g105) & (g948) & (!sk[84]) & (g949) & (g638)) + ((!g105) & (g948) & (sk[84]) & (g949) & (!g638)) + ((g105) & (!g948) & (!sk[84]) & (g949) & (!g638)) + ((g105) & (!g948) & (!sk[84]) & (g949) & (g638)) + ((g105) & (!g948) & (sk[84]) & (!g949) & (!g638)) + ((g105) & (!g948) & (sk[84]) & (g949) & (!g638)) + ((g105) & (g948) & (!sk[84]) & (g949) & (!g638)) + ((g105) & (g948) & (!sk[84]) & (g949) & (g638)) + ((g105) & (g948) & (sk[84]) & (!g949) & (!g638)) + ((g105) & (g948) & (sk[84]) & (g949) & (!g638)));
	assign g951 = (((g944) & (g360) & (g1543) & (g1467) & (g947) & (g950)));
	assign g952 = (((!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g429) & (!g105)) + ((!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g429) & (!g105)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g429) & (!g105)) + ((!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g429) & (!g105)) + ((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g429) & (!g105)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g429) & (!g105)) + ((i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (g429) & (!g105)) + ((i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g429) & (!g105)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g429) & (!g105)));
	assign g953 = (((!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (!g428) & (!g105)) + ((!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (!g428) & (!g105)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g428) & (!g105)) + ((!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g428) & (!g105)) + ((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g428) & (!g105)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g428) & (!g105)) + ((i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (!g428) & (!g105)) + ((i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g428) & (!g105)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g428) & (!g105)));
	assign g954 = (((!sk[88]) & (!g18) & (!g97) & (g102) & (!g578) & (g875)) + ((!sk[88]) & (!g18) & (!g97) & (g102) & (g578) & (!g875)) + ((!sk[88]) & (!g18) & (!g97) & (g102) & (g578) & (g875)) + ((!sk[88]) & (!g18) & (g97) & (!g102) & (!g578) & (!g875)) + ((!sk[88]) & (!g18) & (g97) & (!g102) & (!g578) & (g875)) + ((!sk[88]) & (!g18) & (g97) & (!g102) & (g578) & (!g875)) + ((!sk[88]) & (!g18) & (g97) & (!g102) & (g578) & (g875)) + ((!sk[88]) & (!g18) & (g97) & (g102) & (!g578) & (!g875)) + ((!sk[88]) & (!g18) & (g97) & (g102) & (!g578) & (g875)) + ((!sk[88]) & (!g18) & (g97) & (g102) & (g578) & (!g875)) + ((!sk[88]) & (!g18) & (g97) & (g102) & (g578) & (g875)) + ((!sk[88]) & (g18) & (!g97) & (g102) & (!g578) & (g875)) + ((!sk[88]) & (g18) & (!g97) & (g102) & (g578) & (!g875)) + ((!sk[88]) & (g18) & (!g97) & (g102) & (g578) & (g875)) + ((!sk[88]) & (g18) & (g97) & (!g102) & (!g578) & (!g875)) + ((!sk[88]) & (g18) & (g97) & (!g102) & (!g578) & (g875)) + ((!sk[88]) & (g18) & (g97) & (!g102) & (g578) & (!g875)) + ((!sk[88]) & (g18) & (g97) & (!g102) & (g578) & (g875)) + ((!sk[88]) & (g18) & (g97) & (g102) & (!g578) & (!g875)) + ((!sk[88]) & (g18) & (g97) & (g102) & (!g578) & (g875)) + ((!sk[88]) & (g18) & (g97) & (g102) & (g578) & (!g875)) + ((!sk[88]) & (g18) & (g97) & (g102) & (g578) & (g875)) + ((sk[88]) & (!g18) & (!g97) & (g102) & (!g578) & (!g875)) + ((sk[88]) & (!g18) & (!g97) & (g102) & (!g578) & (g875)) + ((sk[88]) & (!g18) & (!g97) & (g102) & (g578) & (!g875)) + ((sk[88]) & (!g18) & (!g97) & (g102) & (g578) & (g875)) + ((sk[88]) & (!g18) & (g97) & (g102) & (!g578) & (g875)) + ((sk[88]) & (!g18) & (g97) & (g102) & (g578) & (!g875)) + ((sk[88]) & (!g18) & (g97) & (g102) & (g578) & (g875)) + ((sk[88]) & (g18) & (!g97) & (g102) & (!g578) & (!g875)) + ((sk[88]) & (g18) & (!g97) & (g102) & (!g578) & (g875)) + ((sk[88]) & (g18) & (!g97) & (g102) & (g578) & (!g875)) + ((sk[88]) & (g18) & (!g97) & (g102) & (g578) & (g875)) + ((sk[88]) & (g18) & (g97) & (g102) & (!g578) & (!g875)) + ((sk[88]) & (g18) & (g97) & (g102) & (!g578) & (g875)) + ((sk[88]) & (g18) & (g97) & (g102) & (g578) & (!g875)) + ((sk[88]) & (g18) & (g97) & (g102) & (g578) & (g875)));
	assign g955 = (((!sk[89]) & (!g105) & (!g500) & (g954)) + ((!sk[89]) & (!g105) & (g500) & (!g954)) + ((!sk[89]) & (!g105) & (g500) & (g954)) + ((!sk[89]) & (g105) & (!g500) & (g954)) + ((!sk[89]) & (g105) & (g500) & (!g954)) + ((!sk[89]) & (g105) & (g500) & (g954)) + ((sk[89]) & (!g105) & (!g500) & (!g954)) + ((sk[89]) & (g105) & (!g500) & (!g954)) + ((sk[89]) & (g105) & (g500) & (!g954)));
	assign g956 = (((!g887) & (g790) & (g894) & (!g952) & (!g953) & (g955)));
	assign g957 = (((!i_12_) & (!i_13_) & (!i_14_) & (!g107) & (!g91) & (!g105)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g107) & (!g91) & (!g105)) + ((!i_12_) & (!i_13_) & (i_14_) & (!g107) & (!g91) & (!g105)) + ((!i_12_) & (!i_13_) & (i_14_) & (!g107) & (g91) & (!g105)) + ((!i_12_) & (i_13_) & (i_14_) & (!g107) & (!g91) & (!g105)) + ((!i_12_) & (i_13_) & (i_14_) & (!g107) & (g91) & (!g105)) + ((i_12_) & (!i_13_) & (!i_14_) & (!g107) & (!g91) & (!g105)) + ((i_12_) & (!i_13_) & (!i_14_) & (g107) & (!g91) & (!g105)) + ((i_12_) & (i_13_) & (!i_14_) & (!g107) & (!g91) & (!g105)) + ((i_12_) & (i_13_) & (!i_14_) & (g107) & (!g91) & (!g105)) + ((i_12_) & (i_13_) & (i_14_) & (!g107) & (!g91) & (!g105)) + ((i_12_) & (i_13_) & (i_14_) & (!g107) & (g91) & (!g105)));
	assign g958 = (((!i_12_) & (!i_13_) & (!i_14_) & (!g17) & (g27) & (!g105)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g17) & (!g27) & (!g105)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g17) & (g27) & (!g105)) + ((!i_12_) & (!i_13_) & (i_14_) & (!g17) & (g27) & (!g105)) + ((!i_12_) & (!i_13_) & (i_14_) & (g17) & (!g27) & (!g105)) + ((!i_12_) & (!i_13_) & (i_14_) & (g17) & (g27) & (!g105)) + ((!i_12_) & (i_13_) & (!i_14_) & (g17) & (!g27) & (!g105)) + ((!i_12_) & (i_13_) & (!i_14_) & (g17) & (g27) & (!g105)) + ((!i_12_) & (i_13_) & (i_14_) & (!g17) & (g27) & (!g105)) + ((!i_12_) & (i_13_) & (i_14_) & (g17) & (!g27) & (!g105)) + ((!i_12_) & (i_13_) & (i_14_) & (g17) & (g27) & (!g105)) + ((i_12_) & (!i_13_) & (!i_14_) & (g17) & (!g27) & (!g105)) + ((i_12_) & (!i_13_) & (!i_14_) & (g17) & (g27) & (!g105)) + ((i_12_) & (!i_13_) & (i_14_) & (!g17) & (g27) & (!g105)) + ((i_12_) & (!i_13_) & (i_14_) & (g17) & (!g27) & (!g105)) + ((i_12_) & (!i_13_) & (i_14_) & (g17) & (g27) & (!g105)) + ((i_12_) & (i_13_) & (!i_14_) & (g17) & (!g27) & (!g105)) + ((i_12_) & (i_13_) & (!i_14_) & (g17) & (g27) & (!g105)) + ((i_12_) & (i_13_) & (i_14_) & (!g17) & (g27) & (!g105)) + ((i_12_) & (i_13_) & (i_14_) & (g17) & (g27) & (!g105)));
	assign g959 = (((!sk[93]) & (g957) & (!g958)) + ((!sk[93]) & (g957) & (g958)) + ((sk[93]) & (!g957) & (!g958)));
	assign g960 = (((!sk[94]) & (!g538) & (!g111) & (g116) & (!g548) & (g959)) + ((!sk[94]) & (!g538) & (!g111) & (g116) & (g548) & (!g959)) + ((!sk[94]) & (!g538) & (!g111) & (g116) & (g548) & (g959)) + ((!sk[94]) & (!g538) & (g111) & (!g116) & (!g548) & (!g959)) + ((!sk[94]) & (!g538) & (g111) & (!g116) & (!g548) & (g959)) + ((!sk[94]) & (!g538) & (g111) & (!g116) & (g548) & (!g959)) + ((!sk[94]) & (!g538) & (g111) & (!g116) & (g548) & (g959)) + ((!sk[94]) & (!g538) & (g111) & (g116) & (!g548) & (!g959)) + ((!sk[94]) & (!g538) & (g111) & (g116) & (!g548) & (g959)) + ((!sk[94]) & (!g538) & (g111) & (g116) & (g548) & (!g959)) + ((!sk[94]) & (!g538) & (g111) & (g116) & (g548) & (g959)) + ((!sk[94]) & (g538) & (!g111) & (g116) & (!g548) & (g959)) + ((!sk[94]) & (g538) & (!g111) & (g116) & (g548) & (!g959)) + ((!sk[94]) & (g538) & (!g111) & (g116) & (g548) & (g959)) + ((!sk[94]) & (g538) & (g111) & (!g116) & (!g548) & (!g959)) + ((!sk[94]) & (g538) & (g111) & (!g116) & (!g548) & (g959)) + ((!sk[94]) & (g538) & (g111) & (!g116) & (g548) & (!g959)) + ((!sk[94]) & (g538) & (g111) & (!g116) & (g548) & (g959)) + ((!sk[94]) & (g538) & (g111) & (g116) & (!g548) & (!g959)) + ((!sk[94]) & (g538) & (g111) & (g116) & (!g548) & (g959)) + ((!sk[94]) & (g538) & (g111) & (g116) & (g548) & (!g959)) + ((!sk[94]) & (g538) & (g111) & (g116) & (g548) & (g959)) + ((sk[94]) & (!g538) & (g111) & (g116) & (g548) & (g959)));
	assign g961 = (((!g936) & (g940) & (g942) & (g951) & (g956) & (g960)));
	assign g962 = (((!i_8_) & (!i_9_) & (!i_10_) & (i_11_) & (g42) & (g394)) + ((!i_8_) & (!i_9_) & (i_10_) & (!i_11_) & (g42) & (g394)) + ((!i_8_) & (i_9_) & (!i_10_) & (i_11_) & (g42) & (g394)) + ((i_8_) & (!i_9_) & (!i_10_) & (i_11_) & (g42) & (g394)) + ((i_8_) & (!i_9_) & (i_10_) & (!i_11_) & (g42) & (g394)) + ((i_8_) & (i_9_) & (!i_10_) & (i_11_) & (g42) & (g394)) + ((i_8_) & (i_9_) & (i_10_) & (!i_11_) & (g42) & (g394)));
	assign g963 = (((!sk[97]) & (!g926) & (!g961) & (g962)) + ((!sk[97]) & (!g926) & (g961) & (!g962)) + ((!sk[97]) & (!g926) & (g961) & (g962)) + ((!sk[97]) & (g926) & (!g961) & (g962)) + ((!sk[97]) & (g926) & (g961) & (!g962)) + ((!sk[97]) & (g926) & (g961) & (g962)) + ((sk[97]) & (g926) & (g961) & (!g962)));
	assign g964 = (((!g107) & (!sk[98]) & (!g176) & (g487) & (!g652)) + ((!g107) & (!sk[98]) & (!g176) & (g487) & (g652)) + ((!g107) & (!sk[98]) & (g176) & (g487) & (!g652)) + ((!g107) & (!sk[98]) & (g176) & (g487) & (g652)) + ((!g107) & (sk[98]) & (g176) & (!g487) & (!g652)) + ((g107) & (!sk[98]) & (!g176) & (g487) & (!g652)) + ((g107) & (!sk[98]) & (!g176) & (g487) & (g652)) + ((g107) & (!sk[98]) & (g176) & (g487) & (!g652)) + ((g107) & (!sk[98]) & (g176) & (g487) & (g652)) + ((g107) & (sk[98]) & (!g176) & (!g487) & (!g652)) + ((g107) & (sk[98]) & (g176) & (!g487) & (!g652)));
	assign g965 = (((!g83) & (!g735) & (!g738) & (sk[99]) & (g933)) + ((!g83) & (!g735) & (g738) & (!sk[99]) & (!g933)) + ((!g83) & (!g735) & (g738) & (!sk[99]) & (g933)) + ((!g83) & (g735) & (!g738) & (sk[99]) & (g933)) + ((!g83) & (g735) & (g738) & (!sk[99]) & (!g933)) + ((!g83) & (g735) & (g738) & (!sk[99]) & (g933)) + ((g83) & (!g735) & (!g738) & (sk[99]) & (g933)) + ((g83) & (!g735) & (g738) & (!sk[99]) & (!g933)) + ((g83) & (!g735) & (g738) & (!sk[99]) & (g933)) + ((g83) & (g735) & (g738) & (!sk[99]) & (!g933)) + ((g83) & (g735) & (g738) & (!sk[99]) & (g933)));
	assign g966 = (((!sk[100]) & (!g605) & (!g761) & (g934)) + ((!sk[100]) & (!g605) & (g761) & (!g934)) + ((!sk[100]) & (!g605) & (g761) & (g934)) + ((!sk[100]) & (g605) & (!g761) & (g934)) + ((!sk[100]) & (g605) & (g761) & (!g934)) + ((!sk[100]) & (g605) & (g761) & (g934)) + ((sk[100]) & (!g605) & (g761) & (g934)));
	assign g967 = (((!g489) & (!g723) & (g851) & (!sk[101]) & (!g964)) + ((!g489) & (!g723) & (g851) & (!sk[101]) & (g964)) + ((!g489) & (!g723) & (g851) & (sk[101]) & (g964)) + ((!g489) & (g723) & (g851) & (!sk[101]) & (!g964)) + ((!g489) & (g723) & (g851) & (!sk[101]) & (g964)) + ((g489) & (!g723) & (g851) & (!sk[101]) & (!g964)) + ((g489) & (!g723) & (g851) & (!sk[101]) & (g964)) + ((g489) & (g723) & (g851) & (!sk[101]) & (!g964)) + ((g489) & (g723) & (g851) & (!sk[101]) & (g964)));
	assign g968 = (((!sk[102]) & (!g20) & (!g735) & (g847) & (!g966) & (g967)) + ((!sk[102]) & (!g20) & (!g735) & (g847) & (g966) & (!g967)) + ((!sk[102]) & (!g20) & (!g735) & (g847) & (g966) & (g967)) + ((!sk[102]) & (!g20) & (g735) & (!g847) & (!g966) & (!g967)) + ((!sk[102]) & (!g20) & (g735) & (!g847) & (!g966) & (g967)) + ((!sk[102]) & (!g20) & (g735) & (!g847) & (g966) & (!g967)) + ((!sk[102]) & (!g20) & (g735) & (!g847) & (g966) & (g967)) + ((!sk[102]) & (!g20) & (g735) & (g847) & (!g966) & (!g967)) + ((!sk[102]) & (!g20) & (g735) & (g847) & (!g966) & (g967)) + ((!sk[102]) & (!g20) & (g735) & (g847) & (g966) & (!g967)) + ((!sk[102]) & (!g20) & (g735) & (g847) & (g966) & (g967)) + ((!sk[102]) & (g20) & (!g735) & (g847) & (!g966) & (g967)) + ((!sk[102]) & (g20) & (!g735) & (g847) & (g966) & (!g967)) + ((!sk[102]) & (g20) & (!g735) & (g847) & (g966) & (g967)) + ((!sk[102]) & (g20) & (g735) & (!g847) & (!g966) & (!g967)) + ((!sk[102]) & (g20) & (g735) & (!g847) & (!g966) & (g967)) + ((!sk[102]) & (g20) & (g735) & (!g847) & (g966) & (!g967)) + ((!sk[102]) & (g20) & (g735) & (!g847) & (g966) & (g967)) + ((!sk[102]) & (g20) & (g735) & (g847) & (!g966) & (!g967)) + ((!sk[102]) & (g20) & (g735) & (g847) & (!g966) & (g967)) + ((!sk[102]) & (g20) & (g735) & (g847) & (g966) & (!g967)) + ((!sk[102]) & (g20) & (g735) & (g847) & (g966) & (g967)) + ((sk[102]) & (!g20) & (!g735) & (g847) & (g966) & (g967)) + ((sk[102]) & (!g20) & (g735) & (g847) & (g966) & (g967)) + ((sk[102]) & (g20) & (!g735) & (g847) & (g966) & (g967)));
	assign g969 = (((!i_8_) & (!g421) & (g964) & (!sk[103]) & (!g965) & (g968)) + ((!i_8_) & (!g421) & (g964) & (!sk[103]) & (g965) & (!g968)) + ((!i_8_) & (!g421) & (g964) & (!sk[103]) & (g965) & (g968)) + ((!i_8_) & (g421) & (!g964) & (!sk[103]) & (!g965) & (!g968)) + ((!i_8_) & (g421) & (!g964) & (!sk[103]) & (!g965) & (g968)) + ((!i_8_) & (g421) & (!g964) & (!sk[103]) & (g965) & (!g968)) + ((!i_8_) & (g421) & (!g964) & (!sk[103]) & (g965) & (g968)) + ((!i_8_) & (g421) & (!g964) & (sk[103]) & (!g965) & (!g968)) + ((!i_8_) & (g421) & (!g964) & (sk[103]) & (!g965) & (g968)) + ((!i_8_) & (g421) & (!g964) & (sk[103]) & (g965) & (!g968)) + ((!i_8_) & (g421) & (g964) & (!sk[103]) & (!g965) & (!g968)) + ((!i_8_) & (g421) & (g964) & (!sk[103]) & (!g965) & (g968)) + ((!i_8_) & (g421) & (g964) & (!sk[103]) & (g965) & (!g968)) + ((!i_8_) & (g421) & (g964) & (!sk[103]) & (g965) & (g968)) + ((!i_8_) & (g421) & (g964) & (sk[103]) & (!g965) & (!g968)) + ((!i_8_) & (g421) & (g964) & (sk[103]) & (!g965) & (g968)) + ((!i_8_) & (g421) & (g964) & (sk[103]) & (g965) & (!g968)) + ((i_8_) & (!g421) & (g964) & (!sk[103]) & (!g965) & (g968)) + ((i_8_) & (!g421) & (g964) & (!sk[103]) & (g965) & (!g968)) + ((i_8_) & (!g421) & (g964) & (!sk[103]) & (g965) & (g968)) + ((i_8_) & (g421) & (!g964) & (!sk[103]) & (!g965) & (!g968)) + ((i_8_) & (g421) & (!g964) & (!sk[103]) & (!g965) & (g968)) + ((i_8_) & (g421) & (!g964) & (!sk[103]) & (g965) & (!g968)) + ((i_8_) & (g421) & (!g964) & (!sk[103]) & (g965) & (g968)) + ((i_8_) & (g421) & (!g964) & (sk[103]) & (!g965) & (!g968)) + ((i_8_) & (g421) & (!g964) & (sk[103]) & (!g965) & (g968)) + ((i_8_) & (g421) & (!g964) & (sk[103]) & (g965) & (!g968)) + ((i_8_) & (g421) & (g964) & (!sk[103]) & (!g965) & (!g968)) + ((i_8_) & (g421) & (g964) & (!sk[103]) & (!g965) & (g968)) + ((i_8_) & (g421) & (g964) & (!sk[103]) & (g965) & (!g968)) + ((i_8_) & (g421) & (g964) & (!sk[103]) & (g965) & (g968)));
	assign g970 = (((!g164) & (!g253) & (!sk[104]) & (g468) & (!g483) & (g855)) + ((!g164) & (!g253) & (!sk[104]) & (g468) & (g483) & (!g855)) + ((!g164) & (!g253) & (!sk[104]) & (g468) & (g483) & (g855)) + ((!g164) & (!g253) & (sk[104]) & (!g468) & (!g483) & (g855)) + ((!g164) & (!g253) & (sk[104]) & (g468) & (!g483) & (g855)) + ((!g164) & (g253) & (!sk[104]) & (!g468) & (!g483) & (!g855)) + ((!g164) & (g253) & (!sk[104]) & (!g468) & (!g483) & (g855)) + ((!g164) & (g253) & (!sk[104]) & (!g468) & (g483) & (!g855)) + ((!g164) & (g253) & (!sk[104]) & (!g468) & (g483) & (g855)) + ((!g164) & (g253) & (!sk[104]) & (g468) & (!g483) & (!g855)) + ((!g164) & (g253) & (!sk[104]) & (g468) & (!g483) & (g855)) + ((!g164) & (g253) & (!sk[104]) & (g468) & (g483) & (!g855)) + ((!g164) & (g253) & (!sk[104]) & (g468) & (g483) & (g855)) + ((!g164) & (g253) & (sk[104]) & (!g468) & (!g483) & (g855)) + ((!g164) & (g253) & (sk[104]) & (!g468) & (g483) & (g855)) + ((!g164) & (g253) & (sk[104]) & (g468) & (!g483) & (g855)) + ((!g164) & (g253) & (sk[104]) & (g468) & (g483) & (g855)) + ((g164) & (!g253) & (!sk[104]) & (g468) & (!g483) & (g855)) + ((g164) & (!g253) & (!sk[104]) & (g468) & (g483) & (!g855)) + ((g164) & (!g253) & (!sk[104]) & (g468) & (g483) & (g855)) + ((g164) & (!g253) & (sk[104]) & (!g468) & (!g483) & (g855)) + ((g164) & (g253) & (!sk[104]) & (!g468) & (!g483) & (!g855)) + ((g164) & (g253) & (!sk[104]) & (!g468) & (!g483) & (g855)) + ((g164) & (g253) & (!sk[104]) & (!g468) & (g483) & (!g855)) + ((g164) & (g253) & (!sk[104]) & (!g468) & (g483) & (g855)) + ((g164) & (g253) & (!sk[104]) & (g468) & (!g483) & (!g855)) + ((g164) & (g253) & (!sk[104]) & (g468) & (!g483) & (g855)) + ((g164) & (g253) & (!sk[104]) & (g468) & (g483) & (!g855)) + ((g164) & (g253) & (!sk[104]) & (g468) & (g483) & (g855)) + ((g164) & (g253) & (sk[104]) & (!g468) & (!g483) & (g855)) + ((g164) & (g253) & (sk[104]) & (!g468) & (g483) & (g855)));
	assign g971 = (((g898) & (!sk[105]) & (!g945)) + ((g898) & (!sk[105]) & (g945)) + ((g898) & (sk[105]) & (g945)));
	assign g972 = (((!sk[106]) & (!g421) & (!g508) & (g725) & (!g971)) + ((!sk[106]) & (!g421) & (!g508) & (g725) & (g971)) + ((!sk[106]) & (!g421) & (g508) & (g725) & (!g971)) + ((!sk[106]) & (!g421) & (g508) & (g725) & (g971)) + ((!sk[106]) & (g421) & (!g508) & (g725) & (!g971)) + ((!sk[106]) & (g421) & (!g508) & (g725) & (g971)) + ((!sk[106]) & (g421) & (g508) & (g725) & (!g971)) + ((!sk[106]) & (g421) & (g508) & (g725) & (g971)) + ((sk[106]) & (g421) & (!g508) & (!g725) & (!g971)) + ((sk[106]) & (g421) & (!g508) & (!g725) & (g971)) + ((sk[106]) & (g421) & (!g508) & (g725) & (!g971)) + ((sk[106]) & (g421) & (g508) & (!g725) & (!g971)) + ((sk[106]) & (g421) & (g508) & (!g725) & (g971)) + ((sk[106]) & (g421) & (g508) & (g725) & (!g971)) + ((sk[106]) & (g421) & (g508) & (g725) & (g971)));
	assign g973 = (((!g253) & (!g338) & (!g484) & (sk[107]) & (g665)) + ((!g253) & (!g338) & (g484) & (!sk[107]) & (!g665)) + ((!g253) & (!g338) & (g484) & (!sk[107]) & (g665)) + ((!g253) & (!g338) & (g484) & (sk[107]) & (!g665)) + ((!g253) & (!g338) & (g484) & (sk[107]) & (g665)) + ((!g253) & (g338) & (!g484) & (sk[107]) & (!g665)) + ((!g253) & (g338) & (!g484) & (sk[107]) & (g665)) + ((!g253) & (g338) & (g484) & (!sk[107]) & (!g665)) + ((!g253) & (g338) & (g484) & (!sk[107]) & (g665)) + ((!g253) & (g338) & (g484) & (sk[107]) & (!g665)) + ((!g253) & (g338) & (g484) & (sk[107]) & (g665)) + ((g253) & (!g338) & (g484) & (!sk[107]) & (!g665)) + ((g253) & (!g338) & (g484) & (!sk[107]) & (g665)) + ((g253) & (g338) & (g484) & (!sk[107]) & (!g665)) + ((g253) & (g338) & (g484) & (!sk[107]) & (g665)));
	assign g974 = (((!sk[108]) & (!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[108]) & (!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[108]) & (!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g112)) + ((!sk[108]) & (!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g112)) + ((!sk[108]) & (!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((!sk[108]) & (!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g112)) + ((!sk[108]) & (!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g112)) + ((!sk[108]) & (!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g112)) + ((!sk[108]) & (!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[108]) & (!i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[108]) & (!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g112)) + ((!sk[108]) & (i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[108]) & (i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[108]) & (i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g112)) + ((!sk[108]) & (i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g112)) + ((!sk[108]) & (i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((!sk[108]) & (i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g112)) + ((!sk[108]) & (i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g112)) + ((!sk[108]) & (i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g112)) + ((!sk[108]) & (i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[108]) & (i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[108]) & (i_15_) & (i_12_) & (i_13_) & (i_14_) & (g112)) + ((sk[108]) & (!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g112)) + ((sk[108]) & (!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g112)) + ((sk[108]) & (!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g112)) + ((sk[108]) & (!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((sk[108]) & (!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112)) + ((sk[108]) & (!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g112)) + ((sk[108]) & (i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((sk[108]) & (i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((sk[108]) & (i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112)));
	assign g975 = (((!g336) & (!sk[109]) & (!g627) & (g848)) + ((!g336) & (!sk[109]) & (g627) & (!g848)) + ((!g336) & (!sk[109]) & (g627) & (g848)) + ((g336) & (!sk[109]) & (!g627) & (g848)) + ((g336) & (!sk[109]) & (g627) & (!g848)) + ((g336) & (!sk[109]) & (g627) & (g848)) + ((g336) & (sk[109]) & (!g627) & (g848)));
	assign g976 = (((!g164) & (!sk[110]) & (!g335) & (g597) & (!g629)) + ((!g164) & (!sk[110]) & (!g335) & (g597) & (g629)) + ((!g164) & (!sk[110]) & (g335) & (g597) & (!g629)) + ((!g164) & (!sk[110]) & (g335) & (g597) & (g629)) + ((g164) & (!sk[110]) & (!g335) & (g597) & (!g629)) + ((g164) & (!sk[110]) & (!g335) & (g597) & (g629)) + ((g164) & (!sk[110]) & (g335) & (g597) & (!g629)) + ((g164) & (!sk[110]) & (g335) & (g597) & (g629)) + ((g164) & (sk[110]) & (!g335) & (!g597) & (g629)) + ((g164) & (sk[110]) & (!g335) & (g597) & (!g629)) + ((g164) & (sk[110]) & (!g335) & (g597) & (g629)) + ((g164) & (sk[110]) & (g335) & (!g597) & (!g629)) + ((g164) & (sk[110]) & (g335) & (!g597) & (g629)) + ((g164) & (sk[110]) & (g335) & (g597) & (!g629)) + ((g164) & (sk[110]) & (g335) & (g597) & (g629)));
	assign g977 = (((!sk[111]) & (!g164) & (!g974) & (g975) & (!g976)) + ((!sk[111]) & (!g164) & (!g974) & (g975) & (g976)) + ((!sk[111]) & (!g164) & (g974) & (g975) & (!g976)) + ((!sk[111]) & (!g164) & (g974) & (g975) & (g976)) + ((!sk[111]) & (g164) & (!g974) & (g975) & (!g976)) + ((!sk[111]) & (g164) & (!g974) & (g975) & (g976)) + ((!sk[111]) & (g164) & (g974) & (g975) & (!g976)) + ((!sk[111]) & (g164) & (g974) & (g975) & (g976)) + ((sk[111]) & (!g164) & (!g974) & (!g975) & (!g976)) + ((sk[111]) & (!g164) & (!g974) & (g975) & (!g976)) + ((sk[111]) & (!g164) & (g974) & (!g975) & (!g976)) + ((sk[111]) & (!g164) & (g974) & (g975) & (!g976)) + ((sk[111]) & (g164) & (!g974) & (g975) & (!g976)));
	assign g978 = (((!sk[112]) & (!g333) & (!g625) & (g865)) + ((!sk[112]) & (!g333) & (g625) & (!g865)) + ((!sk[112]) & (!g333) & (g625) & (g865)) + ((!sk[112]) & (g333) & (!g625) & (g865)) + ((!sk[112]) & (g333) & (g625) & (!g865)) + ((!sk[112]) & (g333) & (g625) & (g865)) + ((sk[112]) & (!g333) & (!g625) & (!g865)));
	assign g979 = (((g164) & (!g334) & (!g489) & (!g624) & (!g877) & (!g875)) + ((g164) & (!g334) & (!g489) & (!g624) & (!g877) & (g875)) + ((g164) & (!g334) & (!g489) & (!g624) & (g877) & (!g875)) + ((g164) & (!g334) & (!g489) & (!g624) & (g877) & (g875)) + ((g164) & (!g334) & (!g489) & (g624) & (!g877) & (!g875)) + ((g164) & (!g334) & (!g489) & (g624) & (!g877) & (g875)) + ((g164) & (!g334) & (!g489) & (g624) & (g877) & (!g875)) + ((g164) & (!g334) & (!g489) & (g624) & (g877) & (g875)) + ((g164) & (!g334) & (g489) & (!g624) & (!g877) & (!g875)) + ((g164) & (!g334) & (g489) & (!g624) & (!g877) & (g875)) + ((g164) & (!g334) & (g489) & (!g624) & (g877) & (!g875)) + ((g164) & (!g334) & (g489) & (!g624) & (g877) & (g875)) + ((g164) & (!g334) & (g489) & (g624) & (!g877) & (!g875)) + ((g164) & (!g334) & (g489) & (g624) & (!g877) & (g875)) + ((g164) & (!g334) & (g489) & (g624) & (g877) & (!g875)) + ((g164) & (!g334) & (g489) & (g624) & (g877) & (g875)) + ((g164) & (g334) & (!g489) & (!g624) & (!g877) & (!g875)) + ((g164) & (g334) & (!g489) & (!g624) & (!g877) & (g875)) + ((g164) & (g334) & (!g489) & (!g624) & (g877) & (!g875)) + ((g164) & (g334) & (!g489) & (!g624) & (g877) & (g875)) + ((g164) & (g334) & (!g489) & (g624) & (!g877) & (g875)) + ((g164) & (g334) & (!g489) & (g624) & (g877) & (!g875)) + ((g164) & (g334) & (!g489) & (g624) & (g877) & (g875)) + ((g164) & (g334) & (g489) & (!g624) & (!g877) & (!g875)) + ((g164) & (g334) & (g489) & (!g624) & (!g877) & (g875)) + ((g164) & (g334) & (g489) & (!g624) & (g877) & (!g875)) + ((g164) & (g334) & (g489) & (!g624) & (g877) & (g875)) + ((g164) & (g334) & (g489) & (g624) & (!g877) & (!g875)) + ((g164) & (g334) & (g489) & (g624) & (!g877) & (g875)) + ((g164) & (g334) & (g489) & (g624) & (g877) & (!g875)) + ((g164) & (g334) & (g489) & (g624) & (g877) & (g875)));
	assign g980 = (((!g164) & (!g948) & (!g929) & (sk[114]) & (!g978) & (!g979)) + ((!g164) & (!g948) & (!g929) & (sk[114]) & (g978) & (!g979)) + ((!g164) & (!g948) & (g929) & (!sk[114]) & (!g978) & (g979)) + ((!g164) & (!g948) & (g929) & (!sk[114]) & (g978) & (!g979)) + ((!g164) & (!g948) & (g929) & (!sk[114]) & (g978) & (g979)) + ((!g164) & (!g948) & (g929) & (sk[114]) & (!g978) & (!g979)) + ((!g164) & (!g948) & (g929) & (sk[114]) & (g978) & (!g979)) + ((!g164) & (g948) & (!g929) & (!sk[114]) & (!g978) & (!g979)) + ((!g164) & (g948) & (!g929) & (!sk[114]) & (!g978) & (g979)) + ((!g164) & (g948) & (!g929) & (!sk[114]) & (g978) & (!g979)) + ((!g164) & (g948) & (!g929) & (!sk[114]) & (g978) & (g979)) + ((!g164) & (g948) & (!g929) & (sk[114]) & (!g978) & (!g979)) + ((!g164) & (g948) & (!g929) & (sk[114]) & (g978) & (!g979)) + ((!g164) & (g948) & (g929) & (!sk[114]) & (!g978) & (!g979)) + ((!g164) & (g948) & (g929) & (!sk[114]) & (!g978) & (g979)) + ((!g164) & (g948) & (g929) & (!sk[114]) & (g978) & (!g979)) + ((!g164) & (g948) & (g929) & (!sk[114]) & (g978) & (g979)) + ((!g164) & (g948) & (g929) & (sk[114]) & (!g978) & (!g979)) + ((!g164) & (g948) & (g929) & (sk[114]) & (g978) & (!g979)) + ((g164) & (!g948) & (g929) & (!sk[114]) & (!g978) & (g979)) + ((g164) & (!g948) & (g929) & (!sk[114]) & (g978) & (!g979)) + ((g164) & (!g948) & (g929) & (!sk[114]) & (g978) & (g979)) + ((g164) & (g948) & (!g929) & (!sk[114]) & (!g978) & (!g979)) + ((g164) & (g948) & (!g929) & (!sk[114]) & (!g978) & (g979)) + ((g164) & (g948) & (!g929) & (!sk[114]) & (g978) & (!g979)) + ((g164) & (g948) & (!g929) & (!sk[114]) & (g978) & (g979)) + ((g164) & (g948) & (g929) & (!sk[114]) & (!g978) & (!g979)) + ((g164) & (g948) & (g929) & (!sk[114]) & (!g978) & (g979)) + ((g164) & (g948) & (g929) & (!sk[114]) & (g978) & (!g979)) + ((g164) & (g948) & (g929) & (!sk[114]) & (g978) & (g979)) + ((g164) & (g948) & (g929) & (sk[114]) & (g978) & (!g979)));
	assign g981 = (((!g972) & (!g973) & (g676) & (!g977) & (!sk[115]) & (g980)) + ((!g972) & (!g973) & (g676) & (g977) & (!sk[115]) & (!g980)) + ((!g972) & (!g973) & (g676) & (g977) & (!sk[115]) & (g980)) + ((!g972) & (!g973) & (g676) & (g977) & (sk[115]) & (g980)) + ((!g972) & (g973) & (!g676) & (!g977) & (!sk[115]) & (!g980)) + ((!g972) & (g973) & (!g676) & (!g977) & (!sk[115]) & (g980)) + ((!g972) & (g973) & (!g676) & (g977) & (!sk[115]) & (!g980)) + ((!g972) & (g973) & (!g676) & (g977) & (!sk[115]) & (g980)) + ((!g972) & (g973) & (g676) & (!g977) & (!sk[115]) & (!g980)) + ((!g972) & (g973) & (g676) & (!g977) & (!sk[115]) & (g980)) + ((!g972) & (g973) & (g676) & (g977) & (!sk[115]) & (!g980)) + ((!g972) & (g973) & (g676) & (g977) & (!sk[115]) & (g980)) + ((g972) & (!g973) & (g676) & (!g977) & (!sk[115]) & (g980)) + ((g972) & (!g973) & (g676) & (g977) & (!sk[115]) & (!g980)) + ((g972) & (!g973) & (g676) & (g977) & (!sk[115]) & (g980)) + ((g972) & (g973) & (!g676) & (!g977) & (!sk[115]) & (!g980)) + ((g972) & (g973) & (!g676) & (!g977) & (!sk[115]) & (g980)) + ((g972) & (g973) & (!g676) & (g977) & (!sk[115]) & (!g980)) + ((g972) & (g973) & (!g676) & (g977) & (!sk[115]) & (g980)) + ((g972) & (g973) & (g676) & (!g977) & (!sk[115]) & (!g980)) + ((g972) & (g973) & (g676) & (!g977) & (!sk[115]) & (g980)) + ((g972) & (g973) & (g676) & (g977) & (!sk[115]) & (!g980)) + ((g972) & (g973) & (g676) & (g977) & (!sk[115]) & (g980)));
	assign g982 = (((!g164) & (!sk[116]) & (!g253) & (g500) & (!g624) & (g875)) + ((!g164) & (!sk[116]) & (!g253) & (g500) & (g624) & (!g875)) + ((!g164) & (!sk[116]) & (!g253) & (g500) & (g624) & (g875)) + ((!g164) & (!sk[116]) & (g253) & (!g500) & (!g624) & (!g875)) + ((!g164) & (!sk[116]) & (g253) & (!g500) & (!g624) & (g875)) + ((!g164) & (!sk[116]) & (g253) & (!g500) & (g624) & (!g875)) + ((!g164) & (!sk[116]) & (g253) & (!g500) & (g624) & (g875)) + ((!g164) & (!sk[116]) & (g253) & (g500) & (!g624) & (!g875)) + ((!g164) & (!sk[116]) & (g253) & (g500) & (!g624) & (g875)) + ((!g164) & (!sk[116]) & (g253) & (g500) & (g624) & (!g875)) + ((!g164) & (!sk[116]) & (g253) & (g500) & (g624) & (g875)) + ((!g164) & (sk[116]) & (!g253) & (!g500) & (g624) & (!g875)) + ((!g164) & (sk[116]) & (!g253) & (g500) & (g624) & (!g875)) + ((!g164) & (sk[116]) & (g253) & (!g500) & (!g624) & (!g875)) + ((!g164) & (sk[116]) & (g253) & (!g500) & (!g624) & (g875)) + ((!g164) & (sk[116]) & (g253) & (!g500) & (g624) & (!g875)) + ((!g164) & (sk[116]) & (g253) & (!g500) & (g624) & (g875)) + ((!g164) & (sk[116]) & (g253) & (g500) & (!g624) & (!g875)) + ((!g164) & (sk[116]) & (g253) & (g500) & (!g624) & (g875)) + ((!g164) & (sk[116]) & (g253) & (g500) & (g624) & (!g875)) + ((!g164) & (sk[116]) & (g253) & (g500) & (g624) & (g875)) + ((g164) & (!sk[116]) & (!g253) & (g500) & (!g624) & (g875)) + ((g164) & (!sk[116]) & (!g253) & (g500) & (g624) & (!g875)) + ((g164) & (!sk[116]) & (!g253) & (g500) & (g624) & (g875)) + ((g164) & (!sk[116]) & (g253) & (!g500) & (!g624) & (!g875)) + ((g164) & (!sk[116]) & (g253) & (!g500) & (!g624) & (g875)) + ((g164) & (!sk[116]) & (g253) & (!g500) & (g624) & (!g875)) + ((g164) & (!sk[116]) & (g253) & (!g500) & (g624) & (g875)) + ((g164) & (!sk[116]) & (g253) & (g500) & (!g624) & (!g875)) + ((g164) & (!sk[116]) & (g253) & (g500) & (!g624) & (g875)) + ((g164) & (!sk[116]) & (g253) & (g500) & (g624) & (!g875)) + ((g164) & (!sk[116]) & (g253) & (g500) & (g624) & (g875)) + ((g164) & (sk[116]) & (!g253) & (!g500) & (g624) & (!g875)) + ((g164) & (sk[116]) & (g253) & (!g500) & (!g624) & (!g875)) + ((g164) & (sk[116]) & (g253) & (!g500) & (!g624) & (g875)) + ((g164) & (sk[116]) & (g253) & (!g500) & (g624) & (!g875)) + ((g164) & (sk[116]) & (g253) & (!g500) & (g624) & (g875)));
	assign g983 = (((!i_15_) & (!i_12_) & (!i_13_) & (sk[117]) & (!i_14_) & (g112)) + ((!i_15_) & (!i_12_) & (i_13_) & (!sk[117]) & (!i_14_) & (g112)) + ((!i_15_) & (!i_12_) & (i_13_) & (!sk[117]) & (i_14_) & (!g112)) + ((!i_15_) & (!i_12_) & (i_13_) & (!sk[117]) & (i_14_) & (g112)) + ((!i_15_) & (i_12_) & (!i_13_) & (!sk[117]) & (!i_14_) & (!g112)) + ((!i_15_) & (i_12_) & (!i_13_) & (!sk[117]) & (!i_14_) & (g112)) + ((!i_15_) & (i_12_) & (!i_13_) & (!sk[117]) & (i_14_) & (!g112)) + ((!i_15_) & (i_12_) & (!i_13_) & (!sk[117]) & (i_14_) & (g112)) + ((!i_15_) & (i_12_) & (!i_13_) & (sk[117]) & (i_14_) & (g112)) + ((!i_15_) & (i_12_) & (i_13_) & (!sk[117]) & (!i_14_) & (!g112)) + ((!i_15_) & (i_12_) & (i_13_) & (!sk[117]) & (!i_14_) & (g112)) + ((!i_15_) & (i_12_) & (i_13_) & (!sk[117]) & (i_14_) & (!g112)) + ((!i_15_) & (i_12_) & (i_13_) & (!sk[117]) & (i_14_) & (g112)) + ((i_15_) & (!i_12_) & (i_13_) & (!sk[117]) & (!i_14_) & (g112)) + ((i_15_) & (!i_12_) & (i_13_) & (!sk[117]) & (i_14_) & (!g112)) + ((i_15_) & (!i_12_) & (i_13_) & (!sk[117]) & (i_14_) & (g112)) + ((i_15_) & (!i_12_) & (i_13_) & (sk[117]) & (!i_14_) & (g112)) + ((i_15_) & (i_12_) & (!i_13_) & (!sk[117]) & (!i_14_) & (!g112)) + ((i_15_) & (i_12_) & (!i_13_) & (!sk[117]) & (!i_14_) & (g112)) + ((i_15_) & (i_12_) & (!i_13_) & (!sk[117]) & (i_14_) & (!g112)) + ((i_15_) & (i_12_) & (!i_13_) & (!sk[117]) & (i_14_) & (g112)) + ((i_15_) & (i_12_) & (i_13_) & (!sk[117]) & (!i_14_) & (!g112)) + ((i_15_) & (i_12_) & (i_13_) & (!sk[117]) & (!i_14_) & (g112)) + ((i_15_) & (i_12_) & (i_13_) & (!sk[117]) & (i_14_) & (!g112)) + ((i_15_) & (i_12_) & (i_13_) & (!sk[117]) & (i_14_) & (g112)) + ((i_15_) & (i_12_) & (i_13_) & (sk[117]) & (i_14_) & (g112)));
	assign g984 = (((!g113) & (sk[118]) & (g482)) + ((g113) & (!sk[118]) & (!g482)) + ((g113) & (!sk[118]) & (g482)));
	assign g985 = (((!g164) & (!g253) & (!g369) & (!g664) & (sk[119]) & (!g853)) + ((!g164) & (!g253) & (!g369) & (!g664) & (sk[119]) & (g853)) + ((!g164) & (!g253) & (g369) & (!g664) & (!sk[119]) & (g853)) + ((!g164) & (!g253) & (g369) & (g664) & (!sk[119]) & (!g853)) + ((!g164) & (!g253) & (g369) & (g664) & (!sk[119]) & (g853)) + ((!g164) & (g253) & (!g369) & (!g664) & (!sk[119]) & (!g853)) + ((!g164) & (g253) & (!g369) & (!g664) & (!sk[119]) & (g853)) + ((!g164) & (g253) & (!g369) & (!g664) & (sk[119]) & (!g853)) + ((!g164) & (g253) & (!g369) & (!g664) & (sk[119]) & (g853)) + ((!g164) & (g253) & (!g369) & (g664) & (!sk[119]) & (!g853)) + ((!g164) & (g253) & (!g369) & (g664) & (!sk[119]) & (g853)) + ((!g164) & (g253) & (!g369) & (g664) & (sk[119]) & (!g853)) + ((!g164) & (g253) & (!g369) & (g664) & (sk[119]) & (g853)) + ((!g164) & (g253) & (g369) & (!g664) & (!sk[119]) & (!g853)) + ((!g164) & (g253) & (g369) & (!g664) & (!sk[119]) & (g853)) + ((!g164) & (g253) & (g369) & (!g664) & (sk[119]) & (!g853)) + ((!g164) & (g253) & (g369) & (!g664) & (sk[119]) & (g853)) + ((!g164) & (g253) & (g369) & (g664) & (!sk[119]) & (!g853)) + ((!g164) & (g253) & (g369) & (g664) & (!sk[119]) & (g853)) + ((!g164) & (g253) & (g369) & (g664) & (sk[119]) & (!g853)) + ((!g164) & (g253) & (g369) & (g664) & (sk[119]) & (g853)) + ((g164) & (!g253) & (!g369) & (!g664) & (sk[119]) & (!g853)) + ((g164) & (!g253) & (g369) & (!g664) & (!sk[119]) & (g853)) + ((g164) & (!g253) & (g369) & (g664) & (!sk[119]) & (!g853)) + ((g164) & (!g253) & (g369) & (g664) & (!sk[119]) & (g853)) + ((g164) & (g253) & (!g369) & (!g664) & (!sk[119]) & (!g853)) + ((g164) & (g253) & (!g369) & (!g664) & (!sk[119]) & (g853)) + ((g164) & (g253) & (!g369) & (!g664) & (sk[119]) & (!g853)) + ((g164) & (g253) & (!g369) & (g664) & (!sk[119]) & (!g853)) + ((g164) & (g253) & (!g369) & (g664) & (!sk[119]) & (g853)) + ((g164) & (g253) & (!g369) & (g664) & (sk[119]) & (!g853)) + ((g164) & (g253) & (g369) & (!g664) & (!sk[119]) & (!g853)) + ((g164) & (g253) & (g369) & (!g664) & (!sk[119]) & (g853)) + ((g164) & (g253) & (g369) & (!g664) & (sk[119]) & (!g853)) + ((g164) & (g253) & (g369) & (g664) & (!sk[119]) & (!g853)) + ((g164) & (g253) & (g369) & (g664) & (!sk[119]) & (g853)) + ((g164) & (g253) & (g369) & (g664) & (sk[119]) & (!g853)));
	assign g986 = (((!g164) & (!g253) & (!g984) & (!g881) & (!g852) & (g985)) + ((!g164) & (!g253) & (!g984) & (!g881) & (g852) & (g985)) + ((!g164) & (g253) & (!g984) & (!g881) & (!g852) & (g985)) + ((!g164) & (g253) & (!g984) & (!g881) & (g852) & (g985)) + ((!g164) & (g253) & (!g984) & (g881) & (!g852) & (g985)) + ((!g164) & (g253) & (!g984) & (g881) & (g852) & (g985)) + ((!g164) & (g253) & (g984) & (!g881) & (!g852) & (g985)) + ((!g164) & (g253) & (g984) & (!g881) & (g852) & (g985)) + ((!g164) & (g253) & (g984) & (g881) & (!g852) & (g985)) + ((!g164) & (g253) & (g984) & (g881) & (g852) & (g985)) + ((g164) & (!g253) & (!g984) & (!g881) & (!g852) & (g985)) + ((g164) & (g253) & (!g984) & (!g881) & (!g852) & (g985)) + ((g164) & (g253) & (!g984) & (g881) & (!g852) & (g985)));
	assign g987 = (((!g421) & (!g983) & (!sk[121]) & (g986)) + ((!g421) & (!g983) & (sk[121]) & (g986)) + ((!g421) & (g983) & (!sk[121]) & (!g986)) + ((!g421) & (g983) & (!sk[121]) & (g986)) + ((!g421) & (g983) & (sk[121]) & (g986)) + ((g421) & (!g983) & (!sk[121]) & (g986)) + ((g421) & (!g983) & (sk[121]) & (g986)) + ((g421) & (g983) & (!sk[121]) & (!g986)) + ((g421) & (g983) & (!sk[121]) & (g986)));
	assign g988 = (((!sk[122]) & (!g346) & (!g524) & (g982) & (!g987)) + ((!sk[122]) & (!g346) & (!g524) & (g982) & (g987)) + ((!sk[122]) & (!g346) & (g524) & (g982) & (!g987)) + ((!sk[122]) & (!g346) & (g524) & (g982) & (g987)) + ((!sk[122]) & (g346) & (!g524) & (g982) & (!g987)) + ((!sk[122]) & (g346) & (!g524) & (g982) & (g987)) + ((!sk[122]) & (g346) & (g524) & (g982) & (!g987)) + ((!sk[122]) & (g346) & (g524) & (g982) & (g987)) + ((sk[122]) & (g346) & (g524) & (g982) & (g987)));
	assign g989 = (((!g969) & (!g970) & (g981) & (!sk[123]) & (!g988)) + ((!g969) & (!g970) & (g981) & (!sk[123]) & (g988)) + ((!g969) & (g970) & (g981) & (!sk[123]) & (!g988)) + ((!g969) & (g970) & (g981) & (!sk[123]) & (g988)) + ((!g969) & (g970) & (g981) & (sk[123]) & (g988)) + ((g969) & (!g970) & (g981) & (!sk[123]) & (!g988)) + ((g969) & (!g970) & (g981) & (!sk[123]) & (g988)) + ((g969) & (g970) & (g981) & (!sk[123]) & (!g988)) + ((g969) & (g970) & (g981) & (!sk[123]) & (g988)));
	assign g990 = (((!i_9_) & (!i_10_) & (i_11_) & (!sk[124]) & (!g225)) + ((!i_9_) & (!i_10_) & (i_11_) & (!sk[124]) & (g225)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[124]) & (!g225)) + ((!i_9_) & (i_10_) & (i_11_) & (!sk[124]) & (g225)) + ((i_9_) & (!i_10_) & (!i_11_) & (sk[124]) & (g225)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[124]) & (!g225)) + ((i_9_) & (!i_10_) & (i_11_) & (!sk[124]) & (g225)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[124]) & (!g225)) + ((i_9_) & (i_10_) & (i_11_) & (!sk[124]) & (g225)));
	assign g991 = (((!g3) & (!i_12_) & (!i_13_) & (sk[125]) & (!i_14_) & (!g69)) + ((!g3) & (!i_12_) & (!i_13_) & (sk[125]) & (i_14_) & (!g69)) + ((!g3) & (!i_12_) & (!i_13_) & (sk[125]) & (i_14_) & (g69)) + ((!g3) & (!i_12_) & (i_13_) & (!sk[125]) & (!i_14_) & (g69)) + ((!g3) & (!i_12_) & (i_13_) & (!sk[125]) & (i_14_) & (!g69)) + ((!g3) & (!i_12_) & (i_13_) & (!sk[125]) & (i_14_) & (g69)) + ((!g3) & (!i_12_) & (i_13_) & (sk[125]) & (!i_14_) & (!g69)) + ((!g3) & (!i_12_) & (i_13_) & (sk[125]) & (!i_14_) & (g69)) + ((!g3) & (!i_12_) & (i_13_) & (sk[125]) & (i_14_) & (!g69)) + ((!g3) & (!i_12_) & (i_13_) & (sk[125]) & (i_14_) & (g69)) + ((!g3) & (i_12_) & (!i_13_) & (!sk[125]) & (!i_14_) & (!g69)) + ((!g3) & (i_12_) & (!i_13_) & (!sk[125]) & (!i_14_) & (g69)) + ((!g3) & (i_12_) & (!i_13_) & (!sk[125]) & (i_14_) & (!g69)) + ((!g3) & (i_12_) & (!i_13_) & (!sk[125]) & (i_14_) & (g69)) + ((!g3) & (i_12_) & (!i_13_) & (sk[125]) & (!i_14_) & (!g69)) + ((!g3) & (i_12_) & (!i_13_) & (sk[125]) & (i_14_) & (!g69)) + ((!g3) & (i_12_) & (!i_13_) & (sk[125]) & (i_14_) & (g69)) + ((!g3) & (i_12_) & (i_13_) & (!sk[125]) & (!i_14_) & (!g69)) + ((!g3) & (i_12_) & (i_13_) & (!sk[125]) & (!i_14_) & (g69)) + ((!g3) & (i_12_) & (i_13_) & (!sk[125]) & (i_14_) & (!g69)) + ((!g3) & (i_12_) & (i_13_) & (!sk[125]) & (i_14_) & (g69)) + ((!g3) & (i_12_) & (i_13_) & (sk[125]) & (!i_14_) & (!g69)) + ((!g3) & (i_12_) & (i_13_) & (sk[125]) & (i_14_) & (!g69)) + ((g3) & (!i_12_) & (i_13_) & (!sk[125]) & (!i_14_) & (g69)) + ((g3) & (!i_12_) & (i_13_) & (!sk[125]) & (i_14_) & (!g69)) + ((g3) & (!i_12_) & (i_13_) & (!sk[125]) & (i_14_) & (g69)) + ((g3) & (!i_12_) & (i_13_) & (sk[125]) & (!i_14_) & (!g69)) + ((g3) & (!i_12_) & (i_13_) & (sk[125]) & (!i_14_) & (g69)) + ((g3) & (i_12_) & (!i_13_) & (!sk[125]) & (!i_14_) & (!g69)) + ((g3) & (i_12_) & (!i_13_) & (!sk[125]) & (!i_14_) & (g69)) + ((g3) & (i_12_) & (!i_13_) & (!sk[125]) & (i_14_) & (!g69)) + ((g3) & (i_12_) & (!i_13_) & (!sk[125]) & (i_14_) & (g69)) + ((g3) & (i_12_) & (!i_13_) & (sk[125]) & (!i_14_) & (!g69)) + ((g3) & (i_12_) & (i_13_) & (!sk[125]) & (!i_14_) & (!g69)) + ((g3) & (i_12_) & (i_13_) & (!sk[125]) & (!i_14_) & (g69)) + ((g3) & (i_12_) & (i_13_) & (!sk[125]) & (i_14_) & (!g69)) + ((g3) & (i_12_) & (i_13_) & (!sk[125]) & (i_14_) & (g69)) + ((g3) & (i_12_) & (i_13_) & (sk[125]) & (!i_14_) & (!g69)));
	assign g992 = (((!g3) & (!g227) & (g735) & (!sk[126]) & (!g927)) + ((!g3) & (!g227) & (g735) & (!sk[126]) & (g927)) + ((!g3) & (g227) & (!g735) & (sk[126]) & (g927)) + ((!g3) & (g227) & (g735) & (!sk[126]) & (!g927)) + ((!g3) & (g227) & (g735) & (!sk[126]) & (g927)) + ((!g3) & (g227) & (g735) & (sk[126]) & (g927)) + ((g3) & (!g227) & (g735) & (!sk[126]) & (!g927)) + ((g3) & (!g227) & (g735) & (!sk[126]) & (g927)) + ((g3) & (g227) & (!g735) & (sk[126]) & (g927)) + ((g3) & (g227) & (g735) & (!sk[126]) & (!g927)) + ((g3) & (g227) & (g735) & (!sk[126]) & (g927)) + ((g3) & (g227) & (g735) & (sk[126]) & (!g927)) + ((g3) & (g227) & (g735) & (sk[126]) & (g927)));
	assign g993 = (((g17) & (!sk[127]) & (!g174)) + ((g17) & (!sk[127]) & (g174)) + ((g17) & (sk[127]) & (!g174)));
	assign g994 = (((!g17) & (!sk[0]) & (!g27) & (g227)) + ((!g17) & (!sk[0]) & (g27) & (!g227)) + ((!g17) & (!sk[0]) & (g27) & (g227)) + ((!g17) & (sk[0]) & (g27) & (g227)) + ((g17) & (!sk[0]) & (!g27) & (g227)) + ((g17) & (!sk[0]) & (g27) & (!g227)) + ((g17) & (!sk[0]) & (g27) & (g227)) + ((g17) & (sk[0]) & (!g27) & (g227)) + ((g17) & (sk[0]) & (g27) & (g227)));
	assign g995 = (((!g226) & (!g993) & (!sk[1]) & (g725) & (!g994)) + ((!g226) & (!g993) & (!sk[1]) & (g725) & (g994)) + ((!g226) & (!g993) & (sk[1]) & (g725) & (!g994)) + ((!g226) & (g993) & (!sk[1]) & (g725) & (!g994)) + ((!g226) & (g993) & (!sk[1]) & (g725) & (g994)) + ((g226) & (!g993) & (!sk[1]) & (g725) & (!g994)) + ((g226) & (!g993) & (!sk[1]) & (g725) & (g994)) + ((g226) & (!g993) & (sk[1]) & (!g725) & (!g994)) + ((g226) & (!g993) & (sk[1]) & (g725) & (!g994)) + ((g226) & (g993) & (!sk[1]) & (g725) & (!g994)) + ((g226) & (g993) & (!sk[1]) & (g725) & (g994)) + ((g226) & (g993) & (sk[1]) & (!g725) & (!g994)) + ((g226) & (g993) & (sk[1]) & (g725) & (!g994)));
	assign g996 = (((!g3) & (!g19) & (g68) & (!g69) & (!sk[2]) & (g226)) + ((!g3) & (!g19) & (g68) & (g69) & (!sk[2]) & (!g226)) + ((!g3) & (!g19) & (g68) & (g69) & (!sk[2]) & (g226)) + ((!g3) & (g19) & (!g68) & (!g69) & (!sk[2]) & (!g226)) + ((!g3) & (g19) & (!g68) & (!g69) & (!sk[2]) & (g226)) + ((!g3) & (g19) & (!g68) & (g69) & (!sk[2]) & (!g226)) + ((!g3) & (g19) & (!g68) & (g69) & (!sk[2]) & (g226)) + ((!g3) & (g19) & (!g68) & (g69) & (sk[2]) & (!g226)) + ((!g3) & (g19) & (g68) & (!g69) & (!sk[2]) & (!g226)) + ((!g3) & (g19) & (g68) & (!g69) & (!sk[2]) & (g226)) + ((!g3) & (g19) & (g68) & (g69) & (!sk[2]) & (!g226)) + ((!g3) & (g19) & (g68) & (g69) & (!sk[2]) & (g226)) + ((!g3) & (g19) & (g68) & (g69) & (sk[2]) & (!g226)) + ((g3) & (!g19) & (!g68) & (!g69) & (sk[2]) & (!g226)) + ((g3) & (!g19) & (!g68) & (g69) & (sk[2]) & (!g226)) + ((g3) & (!g19) & (g68) & (!g69) & (!sk[2]) & (g226)) + ((g3) & (!g19) & (g68) & (g69) & (!sk[2]) & (!g226)) + ((g3) & (!g19) & (g68) & (g69) & (!sk[2]) & (g226)) + ((g3) & (g19) & (!g68) & (!g69) & (!sk[2]) & (!g226)) + ((g3) & (g19) & (!g68) & (!g69) & (!sk[2]) & (g226)) + ((g3) & (g19) & (!g68) & (!g69) & (sk[2]) & (!g226)) + ((g3) & (g19) & (!g68) & (g69) & (!sk[2]) & (!g226)) + ((g3) & (g19) & (!g68) & (g69) & (!sk[2]) & (g226)) + ((g3) & (g19) & (!g68) & (g69) & (sk[2]) & (!g226)) + ((g3) & (g19) & (g68) & (!g69) & (!sk[2]) & (!g226)) + ((g3) & (g19) & (g68) & (!g69) & (!sk[2]) & (g226)) + ((g3) & (g19) & (g68) & (!g69) & (sk[2]) & (!g226)) + ((g3) & (g19) & (g68) & (g69) & (!sk[2]) & (!g226)) + ((g3) & (g19) & (g68) & (g69) & (!sk[2]) & (g226)) + ((g3) & (g19) & (g68) & (g69) & (sk[2]) & (!g226)));
	assign g997 = (((!g227) & (!g341) & (!g655) & (sk[3]) & (!g996)) + ((!g227) & (!g341) & (g655) & (!sk[3]) & (!g996)) + ((!g227) & (!g341) & (g655) & (!sk[3]) & (g996)) + ((!g227) & (!g341) & (g655) & (sk[3]) & (!g996)) + ((!g227) & (g341) & (!g655) & (sk[3]) & (!g996)) + ((!g227) & (g341) & (g655) & (!sk[3]) & (!g996)) + ((!g227) & (g341) & (g655) & (!sk[3]) & (g996)) + ((!g227) & (g341) & (g655) & (sk[3]) & (!g996)) + ((g227) & (!g341) & (g655) & (!sk[3]) & (!g996)) + ((g227) & (!g341) & (g655) & (!sk[3]) & (g996)) + ((g227) & (g341) & (g655) & (!sk[3]) & (!g996)) + ((g227) & (g341) & (g655) & (!sk[3]) & (g996)) + ((g227) & (g341) & (g655) & (sk[3]) & (!g996)));
	assign g998 = (((!g194) & (!g213) & (!g912) & (sk[4]) & (g997)) + ((!g194) & (!g213) & (g912) & (!sk[4]) & (!g997)) + ((!g194) & (!g213) & (g912) & (!sk[4]) & (g997)) + ((!g194) & (g213) & (!g912) & (sk[4]) & (g997)) + ((!g194) & (g213) & (g912) & (!sk[4]) & (!g997)) + ((!g194) & (g213) & (g912) & (!sk[4]) & (g997)) + ((g194) & (!g213) & (!g912) & (sk[4]) & (g997)) + ((g194) & (!g213) & (g912) & (!sk[4]) & (!g997)) + ((g194) & (!g213) & (g912) & (!sk[4]) & (g997)) + ((g194) & (g213) & (g912) & (!sk[4]) & (!g997)) + ((g194) & (g213) & (g912) & (!sk[4]) & (g997)));
	assign g999 = (((!i_12_) & (!i_13_) & (!i_14_) & (g17) & (!g27) & (!g226)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g17) & (g27) & (!g226)) + ((!i_12_) & (!i_13_) & (i_14_) & (!g17) & (g27) & (!g226)) + ((!i_12_) & (!i_13_) & (i_14_) & (g17) & (!g27) & (!g226)) + ((!i_12_) & (!i_13_) & (i_14_) & (g17) & (g27) & (!g226)) + ((!i_12_) & (i_13_) & (i_14_) & (!g17) & (g27) & (!g226)) + ((!i_12_) & (i_13_) & (i_14_) & (g17) & (!g27) & (!g226)) + ((!i_12_) & (i_13_) & (i_14_) & (g17) & (g27) & (!g226)) + ((i_12_) & (!i_13_) & (!i_14_) & (g17) & (!g27) & (!g226)) + ((i_12_) & (!i_13_) & (!i_14_) & (g17) & (g27) & (!g226)) + ((i_12_) & (!i_13_) & (i_14_) & (g17) & (!g27) & (!g226)) + ((i_12_) & (!i_13_) & (i_14_) & (g17) & (g27) & (!g226)) + ((i_12_) & (i_13_) & (!i_14_) & (g17) & (!g27) & (!g226)) + ((i_12_) & (i_13_) & (!i_14_) & (g17) & (g27) & (!g226)) + ((i_12_) & (i_13_) & (i_14_) & (!g17) & (g27) & (!g226)) + ((i_12_) & (i_13_) & (i_14_) & (g17) & (g27) & (!g226)));
	assign g1000 = (((!sk[6]) & (!g213) & (!g552) & (g469) & (!g999)) + ((!sk[6]) & (!g213) & (!g552) & (g469) & (g999)) + ((!sk[6]) & (!g213) & (g552) & (g469) & (!g999)) + ((!sk[6]) & (!g213) & (g552) & (g469) & (g999)) + ((!sk[6]) & (g213) & (!g552) & (g469) & (!g999)) + ((!sk[6]) & (g213) & (!g552) & (g469) & (g999)) + ((!sk[6]) & (g213) & (g552) & (g469) & (!g999)) + ((!sk[6]) & (g213) & (g552) & (g469) & (g999)) + ((sk[6]) & (!g213) & (!g552) & (!g469) & (!g999)) + ((sk[6]) & (!g213) & (!g552) & (g469) & (!g999)) + ((sk[6]) & (!g213) & (g552) & (!g469) & (!g999)) + ((sk[6]) & (!g213) & (g552) & (g469) & (!g999)) + ((sk[6]) & (g213) & (g552) & (g469) & (!g999)));
	assign g1001 = (((!g226) & (g991) & (!g992) & (g995) & (g998) & (g1000)) + ((g226) & (!g991) & (!g992) & (g995) & (g998) & (g1000)) + ((g226) & (g991) & (!g992) & (g995) & (g998) & (g1000)));
	assign g1002 = (((!i_9_) & (!i_10_) & (!i_11_) & (!i_15_) & (!i_13_) & (!i_14_)) + ((!i_9_) & (!i_10_) & (!i_11_) & (!i_15_) & (!i_13_) & (i_14_)) + ((!i_9_) & (!i_10_) & (!i_11_) & (!i_15_) & (i_13_) & (!i_14_)) + ((!i_9_) & (!i_10_) & (!i_11_) & (!i_15_) & (i_13_) & (i_14_)) + ((!i_9_) & (!i_10_) & (!i_11_) & (i_15_) & (!i_13_) & (i_14_)) + ((!i_9_) & (!i_10_) & (!i_11_) & (i_15_) & (i_13_) & (!i_14_)) + ((!i_9_) & (!i_10_) & (!i_11_) & (i_15_) & (i_13_) & (i_14_)));
	assign g1003 = (((!g70) & (!g121) & (!g654) & (!g990) & (g1001) & (!g1002)) + ((!g70) & (!g121) & (!g654) & (!g990) & (g1001) & (g1002)) + ((!g70) & (!g121) & (g654) & (!g990) & (g1001) & (!g1002)) + ((!g70) & (!g121) & (g654) & (!g990) & (g1001) & (g1002)) + ((!g70) & (g121) & (!g654) & (!g990) & (g1001) & (!g1002)) + ((g70) & (!g121) & (!g654) & (!g990) & (g1001) & (!g1002)) + ((g70) & (!g121) & (!g654) & (!g990) & (g1001) & (g1002)) + ((g70) & (!g121) & (g654) & (!g990) & (g1001) & (!g1002)) + ((g70) & (!g121) & (g654) & (!g990) & (g1001) & (g1002)));
	assign g1004 = (((!sk[10]) & (g445) & (!g142)) + ((!sk[10]) & (g445) & (g142)) + ((sk[10]) & (g445) & (!g142)));
	assign g1005 = (((!sk[11]) & (!g17) & (!g27) & (g142)) + ((!sk[11]) & (!g17) & (g27) & (!g142)) + ((!sk[11]) & (!g17) & (g27) & (g142)) + ((!sk[11]) & (g17) & (!g27) & (g142)) + ((!sk[11]) & (g17) & (g27) & (!g142)) + ((!sk[11]) & (g17) & (g27) & (g142)) + ((sk[11]) & (!g17) & (g27) & (!g142)) + ((sk[11]) & (g17) & (!g27) & (!g142)) + ((sk[11]) & (g17) & (g27) & (!g142)));
	assign g1006 = (((!g428) & (sk[12]) & (!g142)) + ((g428) & (!sk[12]) & (!g142)) + ((g428) & (!sk[12]) & (g142)));
	assign g1007 = (((!i_12_) & (!i_13_) & (!i_14_) & (!g107) & (sk[13]) & (g91)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g107) & (sk[13]) & (g91)) + ((!i_12_) & (!i_13_) & (i_14_) & (!g107) & (!sk[13]) & (g91)) + ((!i_12_) & (!i_13_) & (i_14_) & (g107) & (!sk[13]) & (!g91)) + ((!i_12_) & (!i_13_) & (i_14_) & (g107) & (!sk[13]) & (g91)) + ((!i_12_) & (!i_13_) & (i_14_) & (g107) & (sk[13]) & (g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g107) & (!sk[13]) & (!g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g107) & (!sk[13]) & (g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g107) & (sk[13]) & (!g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g107) & (sk[13]) & (g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (g107) & (!sk[13]) & (!g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (g107) & (!sk[13]) & (g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (g107) & (sk[13]) & (!g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (g107) & (sk[13]) & (g91)) + ((!i_12_) & (i_13_) & (i_14_) & (!g107) & (!sk[13]) & (!g91)) + ((!i_12_) & (i_13_) & (i_14_) & (!g107) & (!sk[13]) & (g91)) + ((!i_12_) & (i_13_) & (i_14_) & (g107) & (!sk[13]) & (!g91)) + ((!i_12_) & (i_13_) & (i_14_) & (g107) & (!sk[13]) & (g91)) + ((!i_12_) & (i_13_) & (i_14_) & (g107) & (sk[13]) & (g91)) + ((i_12_) & (!i_13_) & (!i_14_) & (!g107) & (sk[13]) & (g91)) + ((i_12_) & (!i_13_) & (!i_14_) & (g107) & (sk[13]) & (g91)) + ((i_12_) & (!i_13_) & (i_14_) & (!g107) & (!sk[13]) & (g91)) + ((i_12_) & (!i_13_) & (i_14_) & (!g107) & (sk[13]) & (g91)) + ((i_12_) & (!i_13_) & (i_14_) & (g107) & (!sk[13]) & (!g91)) + ((i_12_) & (!i_13_) & (i_14_) & (g107) & (!sk[13]) & (g91)) + ((i_12_) & (!i_13_) & (i_14_) & (g107) & (sk[13]) & (g91)) + ((i_12_) & (i_13_) & (!i_14_) & (!g107) & (!sk[13]) & (!g91)) + ((i_12_) & (i_13_) & (!i_14_) & (!g107) & (!sk[13]) & (g91)) + ((i_12_) & (i_13_) & (!i_14_) & (!g107) & (sk[13]) & (g91)) + ((i_12_) & (i_13_) & (!i_14_) & (g107) & (!sk[13]) & (!g91)) + ((i_12_) & (i_13_) & (!i_14_) & (g107) & (!sk[13]) & (g91)) + ((i_12_) & (i_13_) & (!i_14_) & (g107) & (sk[13]) & (g91)) + ((i_12_) & (i_13_) & (i_14_) & (!g107) & (!sk[13]) & (!g91)) + ((i_12_) & (i_13_) & (i_14_) & (!g107) & (!sk[13]) & (g91)) + ((i_12_) & (i_13_) & (i_14_) & (g107) & (!sk[13]) & (!g91)) + ((i_12_) & (i_13_) & (i_14_) & (g107) & (!sk[13]) & (g91)) + ((i_12_) & (i_13_) & (i_14_) & (g107) & (sk[13]) & (!g91)) + ((i_12_) & (i_13_) & (i_14_) & (g107) & (sk[13]) & (g91)));
	assign g1008 = (((!sk[14]) & (!g154) & (!g984) & (g852) & (!g853) & (g1007)) + ((!sk[14]) & (!g154) & (!g984) & (g852) & (g853) & (!g1007)) + ((!sk[14]) & (!g154) & (!g984) & (g852) & (g853) & (g1007)) + ((!sk[14]) & (!g154) & (g984) & (!g852) & (!g853) & (!g1007)) + ((!sk[14]) & (!g154) & (g984) & (!g852) & (!g853) & (g1007)) + ((!sk[14]) & (!g154) & (g984) & (!g852) & (g853) & (!g1007)) + ((!sk[14]) & (!g154) & (g984) & (!g852) & (g853) & (g1007)) + ((!sk[14]) & (!g154) & (g984) & (g852) & (!g853) & (!g1007)) + ((!sk[14]) & (!g154) & (g984) & (g852) & (!g853) & (g1007)) + ((!sk[14]) & (!g154) & (g984) & (g852) & (g853) & (!g1007)) + ((!sk[14]) & (!g154) & (g984) & (g852) & (g853) & (g1007)) + ((!sk[14]) & (g154) & (!g984) & (g852) & (!g853) & (g1007)) + ((!sk[14]) & (g154) & (!g984) & (g852) & (g853) & (!g1007)) + ((!sk[14]) & (g154) & (!g984) & (g852) & (g853) & (g1007)) + ((!sk[14]) & (g154) & (g984) & (!g852) & (!g853) & (!g1007)) + ((!sk[14]) & (g154) & (g984) & (!g852) & (!g853) & (g1007)) + ((!sk[14]) & (g154) & (g984) & (!g852) & (g853) & (!g1007)) + ((!sk[14]) & (g154) & (g984) & (!g852) & (g853) & (g1007)) + ((!sk[14]) & (g154) & (g984) & (g852) & (!g853) & (!g1007)) + ((!sk[14]) & (g154) & (g984) & (g852) & (!g853) & (g1007)) + ((!sk[14]) & (g154) & (g984) & (g852) & (g853) & (!g1007)) + ((!sk[14]) & (g154) & (g984) & (g852) & (g853) & (g1007)) + ((sk[14]) & (!g154) & (!g984) & (!g852) & (!g853) & (!g1007)) + ((sk[14]) & (!g154) & (!g984) & (!g852) & (g853) & (!g1007)) + ((sk[14]) & (!g154) & (!g984) & (!g852) & (g853) & (g1007)) + ((sk[14]) & (!g154) & (!g984) & (g852) & (!g853) & (!g1007)) + ((sk[14]) & (!g154) & (!g984) & (g852) & (!g853) & (g1007)) + ((sk[14]) & (!g154) & (!g984) & (g852) & (g853) & (!g1007)) + ((sk[14]) & (!g154) & (!g984) & (g852) & (g853) & (g1007)) + ((sk[14]) & (!g154) & (g984) & (!g852) & (!g853) & (!g1007)) + ((sk[14]) & (!g154) & (g984) & (!g852) & (!g853) & (g1007)) + ((sk[14]) & (!g154) & (g984) & (!g852) & (g853) & (!g1007)) + ((sk[14]) & (!g154) & (g984) & (!g852) & (g853) & (g1007)) + ((sk[14]) & (!g154) & (g984) & (g852) & (!g853) & (!g1007)) + ((sk[14]) & (!g154) & (g984) & (g852) & (!g853) & (g1007)) + ((sk[14]) & (!g154) & (g984) & (g852) & (g853) & (!g1007)) + ((sk[14]) & (!g154) & (g984) & (g852) & (g853) & (g1007)));
	assign g1009 = (((!g159) & (!g217) & (!g984) & (!g974) & (!g983) & (!g1008)) + ((!g159) & (!g217) & (!g984) & (!g974) & (g983) & (!g1008)) + ((!g159) & (g217) & (!g984) & (!g974) & (!g983) & (!g1008)) + ((g159) & (!g217) & (!g984) & (!g974) & (!g983) & (!g1008)) + ((g159) & (!g217) & (!g984) & (!g974) & (g983) & (!g1008)) + ((g159) & (!g217) & (!g984) & (g974) & (!g983) & (!g1008)) + ((g159) & (!g217) & (!g984) & (g974) & (g983) & (!g1008)) + ((g159) & (!g217) & (g984) & (!g974) & (!g983) & (!g1008)) + ((g159) & (!g217) & (g984) & (!g974) & (g983) & (!g1008)) + ((g159) & (!g217) & (g984) & (g974) & (!g983) & (!g1008)) + ((g159) & (!g217) & (g984) & (g974) & (g983) & (!g1008)) + ((g159) & (g217) & (!g984) & (!g974) & (!g983) & (!g1008)) + ((g159) & (g217) & (!g984) & (g974) & (!g983) & (!g1008)) + ((g159) & (g217) & (g984) & (!g974) & (!g983) & (!g1008)) + ((g159) & (g217) & (g984) & (g974) & (!g983) & (!g1008)));
	assign g1010 = (((!g159) & (!g154) & (!g641) & (!g849) & (sk[16]) & (g964)) + ((!g159) & (!g154) & (g641) & (!g849) & (!sk[16]) & (g964)) + ((!g159) & (!g154) & (g641) & (g849) & (!sk[16]) & (!g964)) + ((!g159) & (!g154) & (g641) & (g849) & (!sk[16]) & (g964)) + ((!g159) & (g154) & (!g641) & (!g849) & (!sk[16]) & (!g964)) + ((!g159) & (g154) & (!g641) & (!g849) & (!sk[16]) & (g964)) + ((!g159) & (g154) & (!g641) & (!g849) & (sk[16]) & (!g964)) + ((!g159) & (g154) & (!g641) & (!g849) & (sk[16]) & (g964)) + ((!g159) & (g154) & (!g641) & (g849) & (!sk[16]) & (!g964)) + ((!g159) & (g154) & (!g641) & (g849) & (!sk[16]) & (g964)) + ((!g159) & (g154) & (g641) & (!g849) & (!sk[16]) & (!g964)) + ((!g159) & (g154) & (g641) & (!g849) & (!sk[16]) & (g964)) + ((!g159) & (g154) & (g641) & (g849) & (!sk[16]) & (!g964)) + ((!g159) & (g154) & (g641) & (g849) & (!sk[16]) & (g964)) + ((g159) & (!g154) & (!g641) & (!g849) & (sk[16]) & (g964)) + ((g159) & (!g154) & (!g641) & (g849) & (sk[16]) & (g964)) + ((g159) & (!g154) & (g641) & (!g849) & (!sk[16]) & (g964)) + ((g159) & (!g154) & (g641) & (!g849) & (sk[16]) & (g964)) + ((g159) & (!g154) & (g641) & (g849) & (!sk[16]) & (!g964)) + ((g159) & (!g154) & (g641) & (g849) & (!sk[16]) & (g964)) + ((g159) & (!g154) & (g641) & (g849) & (sk[16]) & (g964)) + ((g159) & (g154) & (!g641) & (!g849) & (!sk[16]) & (!g964)) + ((g159) & (g154) & (!g641) & (!g849) & (!sk[16]) & (g964)) + ((g159) & (g154) & (!g641) & (!g849) & (sk[16]) & (!g964)) + ((g159) & (g154) & (!g641) & (!g849) & (sk[16]) & (g964)) + ((g159) & (g154) & (!g641) & (g849) & (!sk[16]) & (!g964)) + ((g159) & (g154) & (!g641) & (g849) & (!sk[16]) & (g964)) + ((g159) & (g154) & (!g641) & (g849) & (sk[16]) & (!g964)) + ((g159) & (g154) & (!g641) & (g849) & (sk[16]) & (g964)) + ((g159) & (g154) & (g641) & (!g849) & (!sk[16]) & (!g964)) + ((g159) & (g154) & (g641) & (!g849) & (!sk[16]) & (g964)) + ((g159) & (g154) & (g641) & (!g849) & (sk[16]) & (!g964)) + ((g159) & (g154) & (g641) & (!g849) & (sk[16]) & (g964)) + ((g159) & (g154) & (g641) & (g849) & (!sk[16]) & (!g964)) + ((g159) & (g154) & (g641) & (g849) & (!sk[16]) & (g964)) + ((g159) & (g154) & (g641) & (g849) & (sk[16]) & (!g964)) + ((g159) & (g154) & (g641) & (g849) & (sk[16]) & (g964)));
	assign g1011 = (((!g159) & (!sk[17]) & (!g975) & (g964) & (!g1010) & (g1007)) + ((!g159) & (!sk[17]) & (!g975) & (g964) & (g1010) & (!g1007)) + ((!g159) & (!sk[17]) & (!g975) & (g964) & (g1010) & (g1007)) + ((!g159) & (!sk[17]) & (g975) & (!g964) & (!g1010) & (!g1007)) + ((!g159) & (!sk[17]) & (g975) & (!g964) & (!g1010) & (g1007)) + ((!g159) & (!sk[17]) & (g975) & (!g964) & (g1010) & (!g1007)) + ((!g159) & (!sk[17]) & (g975) & (!g964) & (g1010) & (g1007)) + ((!g159) & (!sk[17]) & (g975) & (g964) & (!g1010) & (!g1007)) + ((!g159) & (!sk[17]) & (g975) & (g964) & (!g1010) & (g1007)) + ((!g159) & (!sk[17]) & (g975) & (g964) & (g1010) & (!g1007)) + ((!g159) & (!sk[17]) & (g975) & (g964) & (g1010) & (g1007)) + ((!g159) & (sk[17]) & (g975) & (g964) & (g1010) & (g1007)) + ((g159) & (!sk[17]) & (!g975) & (g964) & (!g1010) & (g1007)) + ((g159) & (!sk[17]) & (!g975) & (g964) & (g1010) & (!g1007)) + ((g159) & (!sk[17]) & (!g975) & (g964) & (g1010) & (g1007)) + ((g159) & (!sk[17]) & (g975) & (!g964) & (!g1010) & (!g1007)) + ((g159) & (!sk[17]) & (g975) & (!g964) & (!g1010) & (g1007)) + ((g159) & (!sk[17]) & (g975) & (!g964) & (g1010) & (!g1007)) + ((g159) & (!sk[17]) & (g975) & (!g964) & (g1010) & (g1007)) + ((g159) & (!sk[17]) & (g975) & (g964) & (!g1010) & (!g1007)) + ((g159) & (!sk[17]) & (g975) & (g964) & (!g1010) & (g1007)) + ((g159) & (!sk[17]) & (g975) & (g964) & (g1010) & (!g1007)) + ((g159) & (!sk[17]) & (g975) & (g964) & (g1010) & (g1007)) + ((g159) & (sk[17]) & (!g975) & (!g964) & (g1010) & (!g1007)) + ((g159) & (sk[17]) & (!g975) & (!g964) & (g1010) & (g1007)) + ((g159) & (sk[17]) & (!g975) & (g964) & (g1010) & (!g1007)) + ((g159) & (sk[17]) & (!g975) & (g964) & (g1010) & (g1007)) + ((g159) & (sk[17]) & (g975) & (!g964) & (g1010) & (!g1007)) + ((g159) & (sk[17]) & (g975) & (!g964) & (g1010) & (g1007)) + ((g159) & (sk[17]) & (g975) & (g964) & (g1010) & (!g1007)) + ((g159) & (sk[17]) & (g975) & (g964) & (g1010) & (g1007)));
	assign g1012 = (((!g69) & (!g154) & (!sk[18]) & (g482) & (!g743)) + ((!g69) & (!g154) & (!sk[18]) & (g482) & (g743)) + ((!g69) & (!g154) & (sk[18]) & (!g482) & (g743)) + ((!g69) & (!g154) & (sk[18]) & (g482) & (g743)) + ((!g69) & (g154) & (!sk[18]) & (g482) & (!g743)) + ((!g69) & (g154) & (!sk[18]) & (g482) & (g743)) + ((g69) & (!g154) & (!sk[18]) & (g482) & (!g743)) + ((g69) & (!g154) & (!sk[18]) & (g482) & (g743)) + ((g69) & (!g154) & (sk[18]) & (!g482) & (g743)) + ((g69) & (!g154) & (sk[18]) & (g482) & (!g743)) + ((g69) & (!g154) & (sk[18]) & (g482) & (g743)) + ((g69) & (g154) & (!sk[18]) & (g482) & (!g743)) + ((g69) & (g154) & (!sk[18]) & (g482) & (g743)));
	assign g1013 = (((!g725) & (!g929) & (!sk[19]) & (g971) & (!g1012)) + ((!g725) & (!g929) & (!sk[19]) & (g971) & (g1012)) + ((!g725) & (g929) & (!sk[19]) & (g971) & (!g1012)) + ((!g725) & (g929) & (!sk[19]) & (g971) & (g1012)) + ((g725) & (!g929) & (!sk[19]) & (g971) & (!g1012)) + ((g725) & (!g929) & (!sk[19]) & (g971) & (g1012)) + ((g725) & (g929) & (!sk[19]) & (g971) & (!g1012)) + ((g725) & (g929) & (!sk[19]) & (g971) & (g1012)) + ((g725) & (g929) & (sk[19]) & (g971) & (!g1012)));
	assign g1014 = (((!g154) & (!sk[20]) & (!g217) & (g974) & (!g1013) & (g1455)) + ((!g154) & (!sk[20]) & (!g217) & (g974) & (g1013) & (!g1455)) + ((!g154) & (!sk[20]) & (!g217) & (g974) & (g1013) & (g1455)) + ((!g154) & (!sk[20]) & (g217) & (!g974) & (!g1013) & (!g1455)) + ((!g154) & (!sk[20]) & (g217) & (!g974) & (!g1013) & (g1455)) + ((!g154) & (!sk[20]) & (g217) & (!g974) & (g1013) & (!g1455)) + ((!g154) & (!sk[20]) & (g217) & (!g974) & (g1013) & (g1455)) + ((!g154) & (!sk[20]) & (g217) & (g974) & (!g1013) & (!g1455)) + ((!g154) & (!sk[20]) & (g217) & (g974) & (!g1013) & (g1455)) + ((!g154) & (!sk[20]) & (g217) & (g974) & (g1013) & (!g1455)) + ((!g154) & (!sk[20]) & (g217) & (g974) & (g1013) & (g1455)) + ((!g154) & (sk[20]) & (!g217) & (!g974) & (!g1013) & (!g1455)) + ((!g154) & (sk[20]) & (!g217) & (!g974) & (g1013) & (!g1455)) + ((!g154) & (sk[20]) & (g217) & (!g974) & (g1013) & (!g1455)) + ((g154) & (!sk[20]) & (!g217) & (g974) & (!g1013) & (g1455)) + ((g154) & (!sk[20]) & (!g217) & (g974) & (g1013) & (!g1455)) + ((g154) & (!sk[20]) & (!g217) & (g974) & (g1013) & (g1455)) + ((g154) & (!sk[20]) & (g217) & (!g974) & (!g1013) & (!g1455)) + ((g154) & (!sk[20]) & (g217) & (!g974) & (!g1013) & (g1455)) + ((g154) & (!sk[20]) & (g217) & (!g974) & (g1013) & (!g1455)) + ((g154) & (!sk[20]) & (g217) & (!g974) & (g1013) & (g1455)) + ((g154) & (!sk[20]) & (g217) & (g974) & (!g1013) & (!g1455)) + ((g154) & (!sk[20]) & (g217) & (g974) & (!g1013) & (g1455)) + ((g154) & (!sk[20]) & (g217) & (g974) & (g1013) & (!g1455)) + ((g154) & (!sk[20]) & (g217) & (g974) & (g1013) & (g1455)) + ((g154) & (sk[20]) & (!g217) & (!g974) & (!g1013) & (!g1455)) + ((g154) & (sk[20]) & (!g217) & (!g974) & (g1013) & (!g1455)) + ((g154) & (sk[20]) & (!g217) & (g974) & (!g1013) & (!g1455)) + ((g154) & (sk[20]) & (!g217) & (g974) & (g1013) & (!g1455)) + ((g154) & (sk[20]) & (g217) & (!g974) & (g1013) & (!g1455)) + ((g154) & (sk[20]) & (g217) & (g974) & (g1013) & (!g1455)));
	assign g1015 = (((!g335) & (!g508) & (!sk[21]) & (g629) & (!g851)) + ((!g335) & (!g508) & (!sk[21]) & (g629) & (g851)) + ((!g335) & (!g508) & (sk[21]) & (!g629) & (g851)) + ((!g335) & (g508) & (!sk[21]) & (g629) & (!g851)) + ((!g335) & (g508) & (!sk[21]) & (g629) & (g851)) + ((g335) & (!g508) & (!sk[21]) & (g629) & (!g851)) + ((g335) & (!g508) & (!sk[21]) & (g629) & (g851)) + ((g335) & (g508) & (!sk[21]) & (g629) & (!g851)) + ((g335) & (g508) & (!sk[21]) & (g629) & (g851)));
	assign g1016 = (((!g159) & (!sk[22]) & (!g635) & (g932) & (!g966) & (g1015)) + ((!g159) & (!sk[22]) & (!g635) & (g932) & (g966) & (!g1015)) + ((!g159) & (!sk[22]) & (!g635) & (g932) & (g966) & (g1015)) + ((!g159) & (!sk[22]) & (g635) & (!g932) & (!g966) & (!g1015)) + ((!g159) & (!sk[22]) & (g635) & (!g932) & (!g966) & (g1015)) + ((!g159) & (!sk[22]) & (g635) & (!g932) & (g966) & (!g1015)) + ((!g159) & (!sk[22]) & (g635) & (!g932) & (g966) & (g1015)) + ((!g159) & (!sk[22]) & (g635) & (g932) & (!g966) & (!g1015)) + ((!g159) & (!sk[22]) & (g635) & (g932) & (!g966) & (g1015)) + ((!g159) & (!sk[22]) & (g635) & (g932) & (g966) & (!g1015)) + ((!g159) & (!sk[22]) & (g635) & (g932) & (g966) & (g1015)) + ((!g159) & (sk[22]) & (!g635) & (!g932) & (!g966) & (!g1015)) + ((!g159) & (sk[22]) & (!g635) & (!g932) & (!g966) & (g1015)) + ((!g159) & (sk[22]) & (!g635) & (!g932) & (g966) & (!g1015)) + ((!g159) & (sk[22]) & (!g635) & (!g932) & (g966) & (g1015)) + ((!g159) & (sk[22]) & (!g635) & (g932) & (!g966) & (!g1015)) + ((!g159) & (sk[22]) & (!g635) & (g932) & (!g966) & (g1015)) + ((!g159) & (sk[22]) & (!g635) & (g932) & (g966) & (!g1015)) + ((!g159) & (sk[22]) & (g635) & (!g932) & (!g966) & (!g1015)) + ((!g159) & (sk[22]) & (g635) & (!g932) & (!g966) & (g1015)) + ((!g159) & (sk[22]) & (g635) & (!g932) & (g966) & (!g1015)) + ((!g159) & (sk[22]) & (g635) & (!g932) & (g966) & (g1015)) + ((!g159) & (sk[22]) & (g635) & (g932) & (!g966) & (!g1015)) + ((!g159) & (sk[22]) & (g635) & (g932) & (!g966) & (g1015)) + ((!g159) & (sk[22]) & (g635) & (g932) & (g966) & (!g1015)) + ((!g159) & (sk[22]) & (g635) & (g932) & (g966) & (g1015)) + ((g159) & (!sk[22]) & (!g635) & (g932) & (!g966) & (g1015)) + ((g159) & (!sk[22]) & (!g635) & (g932) & (g966) & (!g1015)) + ((g159) & (!sk[22]) & (!g635) & (g932) & (g966) & (g1015)) + ((g159) & (!sk[22]) & (g635) & (!g932) & (!g966) & (!g1015)) + ((g159) & (!sk[22]) & (g635) & (!g932) & (!g966) & (g1015)) + ((g159) & (!sk[22]) & (g635) & (!g932) & (g966) & (!g1015)) + ((g159) & (!sk[22]) & (g635) & (!g932) & (g966) & (g1015)) + ((g159) & (!sk[22]) & (g635) & (g932) & (!g966) & (!g1015)) + ((g159) & (!sk[22]) & (g635) & (g932) & (!g966) & (g1015)) + ((g159) & (!sk[22]) & (g635) & (g932) & (g966) & (!g1015)) + ((g159) & (!sk[22]) & (g635) & (g932) & (g966) & (g1015)));
	assign g1017 = (((!g154) & (!g875) & (!g1016) & (g365) & (g632) & (g880)) + ((g154) & (!g875) & (!g1016) & (g365) & (g632) & (g880)) + ((g154) & (g875) & (!g1016) & (g365) & (g632) & (g880)));
	assign g1018 = (((!g600) & (!g1009) & (g1011) & (!g1014) & (!sk[24]) & (g1017)) + ((!g600) & (!g1009) & (g1011) & (g1014) & (!sk[24]) & (!g1017)) + ((!g600) & (!g1009) & (g1011) & (g1014) & (!sk[24]) & (g1017)) + ((!g600) & (g1009) & (!g1011) & (!g1014) & (!sk[24]) & (!g1017)) + ((!g600) & (g1009) & (!g1011) & (!g1014) & (!sk[24]) & (g1017)) + ((!g600) & (g1009) & (!g1011) & (g1014) & (!sk[24]) & (!g1017)) + ((!g600) & (g1009) & (!g1011) & (g1014) & (!sk[24]) & (g1017)) + ((!g600) & (g1009) & (g1011) & (!g1014) & (!sk[24]) & (!g1017)) + ((!g600) & (g1009) & (g1011) & (!g1014) & (!sk[24]) & (g1017)) + ((!g600) & (g1009) & (g1011) & (g1014) & (!sk[24]) & (!g1017)) + ((!g600) & (g1009) & (g1011) & (g1014) & (!sk[24]) & (g1017)) + ((g600) & (!g1009) & (g1011) & (!g1014) & (!sk[24]) & (g1017)) + ((g600) & (!g1009) & (g1011) & (g1014) & (!sk[24]) & (!g1017)) + ((g600) & (!g1009) & (g1011) & (g1014) & (!sk[24]) & (g1017)) + ((g600) & (g1009) & (!g1011) & (!g1014) & (!sk[24]) & (!g1017)) + ((g600) & (g1009) & (!g1011) & (!g1014) & (!sk[24]) & (g1017)) + ((g600) & (g1009) & (!g1011) & (g1014) & (!sk[24]) & (!g1017)) + ((g600) & (g1009) & (!g1011) & (g1014) & (!sk[24]) & (g1017)) + ((g600) & (g1009) & (g1011) & (!g1014) & (!sk[24]) & (!g1017)) + ((g600) & (g1009) & (g1011) & (!g1014) & (!sk[24]) & (g1017)) + ((g600) & (g1009) & (g1011) & (g1014) & (!sk[24]) & (!g1017)) + ((g600) & (g1009) & (g1011) & (g1014) & (!sk[24]) & (g1017)) + ((g600) & (g1009) & (g1011) & (g1014) & (sk[24]) & (g1017)));
	assign g1019 = (((!sk[25]) & (!g357) & (!g857) & (g948)) + ((!sk[25]) & (!g357) & (g857) & (!g948)) + ((!sk[25]) & (!g357) & (g857) & (g948)) + ((!sk[25]) & (g357) & (!g857) & (g948)) + ((!sk[25]) & (g357) & (g857) & (!g948)) + ((!sk[25]) & (g357) & (g857) & (g948)) + ((sk[25]) & (!g357) & (!g857) & (g948)));
	assign g1020 = (((!g125) & (!g469) & (g720) & (!g929) & (!sk[26]) & (g1019)) + ((!g125) & (!g469) & (g720) & (g929) & (!sk[26]) & (!g1019)) + ((!g125) & (!g469) & (g720) & (g929) & (!sk[26]) & (g1019)) + ((!g125) & (g469) & (!g720) & (!g929) & (!sk[26]) & (!g1019)) + ((!g125) & (g469) & (!g720) & (!g929) & (!sk[26]) & (g1019)) + ((!g125) & (g469) & (!g720) & (g929) & (!sk[26]) & (!g1019)) + ((!g125) & (g469) & (!g720) & (g929) & (!sk[26]) & (g1019)) + ((!g125) & (g469) & (g720) & (!g929) & (!sk[26]) & (!g1019)) + ((!g125) & (g469) & (g720) & (!g929) & (!sk[26]) & (g1019)) + ((!g125) & (g469) & (g720) & (g929) & (!sk[26]) & (!g1019)) + ((!g125) & (g469) & (g720) & (g929) & (!sk[26]) & (g1019)) + ((g125) & (!g469) & (!g720) & (!g929) & (sk[26]) & (!g1019)) + ((g125) & (!g469) & (!g720) & (!g929) & (sk[26]) & (g1019)) + ((g125) & (!g469) & (!g720) & (g929) & (sk[26]) & (!g1019)) + ((g125) & (!g469) & (!g720) & (g929) & (sk[26]) & (g1019)) + ((g125) & (!g469) & (g720) & (!g929) & (!sk[26]) & (g1019)) + ((g125) & (!g469) & (g720) & (!g929) & (sk[26]) & (!g1019)) + ((g125) & (!g469) & (g720) & (!g929) & (sk[26]) & (g1019)) + ((g125) & (!g469) & (g720) & (g929) & (!sk[26]) & (!g1019)) + ((g125) & (!g469) & (g720) & (g929) & (!sk[26]) & (g1019)) + ((g125) & (!g469) & (g720) & (g929) & (sk[26]) & (!g1019)) + ((g125) & (!g469) & (g720) & (g929) & (sk[26]) & (g1019)) + ((g125) & (g469) & (!g720) & (!g929) & (!sk[26]) & (!g1019)) + ((g125) & (g469) & (!g720) & (!g929) & (!sk[26]) & (g1019)) + ((g125) & (g469) & (!g720) & (!g929) & (sk[26]) & (!g1019)) + ((g125) & (g469) & (!g720) & (!g929) & (sk[26]) & (g1019)) + ((g125) & (g469) & (!g720) & (g929) & (!sk[26]) & (!g1019)) + ((g125) & (g469) & (!g720) & (g929) & (!sk[26]) & (g1019)) + ((g125) & (g469) & (!g720) & (g929) & (sk[26]) & (!g1019)) + ((g125) & (g469) & (!g720) & (g929) & (sk[26]) & (g1019)) + ((g125) & (g469) & (g720) & (!g929) & (!sk[26]) & (!g1019)) + ((g125) & (g469) & (g720) & (!g929) & (!sk[26]) & (g1019)) + ((g125) & (g469) & (g720) & (!g929) & (sk[26]) & (!g1019)) + ((g125) & (g469) & (g720) & (!g929) & (sk[26]) & (g1019)) + ((g125) & (g469) & (g720) & (g929) & (!sk[26]) & (!g1019)) + ((g125) & (g469) & (g720) & (g929) & (!sk[26]) & (g1019)) + ((g125) & (g469) & (g720) & (g929) & (sk[26]) & (!g1019)));
	assign g1021 = (((!i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (sk[27]) & (g112)) + ((!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (sk[27]) & (g112)) + ((!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (!sk[27]) & (g112)) + ((!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (sk[27]) & (g112)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!sk[27]) & (!g112)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!sk[27]) & (g112)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (sk[27]) & (g112)) + ((!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!sk[27]) & (!g112)) + ((!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!sk[27]) & (g112)) + ((!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (sk[27]) & (g112)) + ((!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!sk[27]) & (!g112)) + ((!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!sk[27]) & (g112)) + ((!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (sk[27]) & (g112)) + ((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!sk[27]) & (!g112)) + ((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!sk[27]) & (g112)) + ((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (sk[27]) & (g112)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (!sk[27]) & (!g112)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (!sk[27]) & (g112)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (sk[27]) & (g112)) + ((i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (!sk[27]) & (g112)) + ((i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (sk[27]) & (g112)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!sk[27]) & (!g112)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!sk[27]) & (g112)) + ((i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!sk[27]) & (!g112)) + ((i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!sk[27]) & (g112)) + ((i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!sk[27]) & (!g112)) + ((i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!sk[27]) & (g112)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!sk[27]) & (!g112)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!sk[27]) & (g112)) + ((i_15_) & (i_12_) & (i_13_) & (i_14_) & (!sk[27]) & (!g112)) + ((i_15_) & (i_12_) & (i_13_) & (i_14_) & (!sk[27]) & (g112)));
	assign g1022 = (((!i_12_) & (!sk[28]) & (!i_13_) & (i_14_) & (!g144) & (g113)) + ((!i_12_) & (!sk[28]) & (!i_13_) & (i_14_) & (g144) & (!g113)) + ((!i_12_) & (!sk[28]) & (!i_13_) & (i_14_) & (g144) & (g113)) + ((!i_12_) & (!sk[28]) & (i_13_) & (!i_14_) & (!g144) & (!g113)) + ((!i_12_) & (!sk[28]) & (i_13_) & (!i_14_) & (!g144) & (g113)) + ((!i_12_) & (!sk[28]) & (i_13_) & (!i_14_) & (g144) & (!g113)) + ((!i_12_) & (!sk[28]) & (i_13_) & (!i_14_) & (g144) & (g113)) + ((!i_12_) & (!sk[28]) & (i_13_) & (i_14_) & (!g144) & (!g113)) + ((!i_12_) & (!sk[28]) & (i_13_) & (i_14_) & (!g144) & (g113)) + ((!i_12_) & (!sk[28]) & (i_13_) & (i_14_) & (g144) & (!g113)) + ((!i_12_) & (!sk[28]) & (i_13_) & (i_14_) & (g144) & (g113)) + ((!i_12_) & (sk[28]) & (!i_13_) & (i_14_) & (g144) & (!g113)) + ((i_12_) & (!sk[28]) & (!i_13_) & (i_14_) & (!g144) & (g113)) + ((i_12_) & (!sk[28]) & (!i_13_) & (i_14_) & (g144) & (!g113)) + ((i_12_) & (!sk[28]) & (!i_13_) & (i_14_) & (g144) & (g113)) + ((i_12_) & (!sk[28]) & (i_13_) & (!i_14_) & (!g144) & (!g113)) + ((i_12_) & (!sk[28]) & (i_13_) & (!i_14_) & (!g144) & (g113)) + ((i_12_) & (!sk[28]) & (i_13_) & (!i_14_) & (g144) & (!g113)) + ((i_12_) & (!sk[28]) & (i_13_) & (!i_14_) & (g144) & (g113)) + ((i_12_) & (!sk[28]) & (i_13_) & (i_14_) & (!g144) & (!g113)) + ((i_12_) & (!sk[28]) & (i_13_) & (i_14_) & (!g144) & (g113)) + ((i_12_) & (!sk[28]) & (i_13_) & (i_14_) & (g144) & (!g113)) + ((i_12_) & (!sk[28]) & (i_13_) & (i_14_) & (g144) & (g113)) + ((i_12_) & (sk[28]) & (i_13_) & (i_14_) & (g144) & (!g113)));
	assign g1023 = (((!g131) & (!g197) & (!g557) & (sk[29]) & (g664)) + ((!g131) & (!g197) & (g557) & (!sk[29]) & (!g664)) + ((!g131) & (!g197) & (g557) & (!sk[29]) & (g664)) + ((!g131) & (!g197) & (g557) & (sk[29]) & (!g664)) + ((!g131) & (!g197) & (g557) & (sk[29]) & (g664)) + ((!g131) & (g197) & (!g557) & (sk[29]) & (!g664)) + ((!g131) & (g197) & (!g557) & (sk[29]) & (g664)) + ((!g131) & (g197) & (g557) & (!sk[29]) & (!g664)) + ((!g131) & (g197) & (g557) & (!sk[29]) & (g664)) + ((!g131) & (g197) & (g557) & (sk[29]) & (!g664)) + ((!g131) & (g197) & (g557) & (sk[29]) & (g664)) + ((g131) & (!g197) & (g557) & (!sk[29]) & (!g664)) + ((g131) & (!g197) & (g557) & (!sk[29]) & (g664)) + ((g131) & (g197) & (g557) & (!sk[29]) & (!g664)) + ((g131) & (g197) & (g557) & (!sk[29]) & (g664)));
	assign g1024 = (((!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g125) & (g112)) + ((!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g125) & (g112)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g125) & (g112)) + ((!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g125) & (g112)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g125) & (g112)) + ((i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g125) & (g112)));
	assign g1025 = (((!g131) & (!g1021) & (!sk[31]) & (g1022) & (!g1023) & (g1024)) + ((!g131) & (!g1021) & (!sk[31]) & (g1022) & (g1023) & (!g1024)) + ((!g131) & (!g1021) & (!sk[31]) & (g1022) & (g1023) & (g1024)) + ((!g131) & (!g1021) & (sk[31]) & (!g1022) & (!g1023) & (!g1024)) + ((!g131) & (g1021) & (!sk[31]) & (!g1022) & (!g1023) & (!g1024)) + ((!g131) & (g1021) & (!sk[31]) & (!g1022) & (!g1023) & (g1024)) + ((!g131) & (g1021) & (!sk[31]) & (!g1022) & (g1023) & (!g1024)) + ((!g131) & (g1021) & (!sk[31]) & (!g1022) & (g1023) & (g1024)) + ((!g131) & (g1021) & (!sk[31]) & (g1022) & (!g1023) & (!g1024)) + ((!g131) & (g1021) & (!sk[31]) & (g1022) & (!g1023) & (g1024)) + ((!g131) & (g1021) & (!sk[31]) & (g1022) & (g1023) & (!g1024)) + ((!g131) & (g1021) & (!sk[31]) & (g1022) & (g1023) & (g1024)) + ((g131) & (!g1021) & (!sk[31]) & (g1022) & (!g1023) & (g1024)) + ((g131) & (!g1021) & (!sk[31]) & (g1022) & (g1023) & (!g1024)) + ((g131) & (!g1021) & (!sk[31]) & (g1022) & (g1023) & (g1024)) + ((g131) & (!g1021) & (sk[31]) & (!g1022) & (!g1023) & (!g1024)) + ((g131) & (g1021) & (!sk[31]) & (!g1022) & (!g1023) & (!g1024)) + ((g131) & (g1021) & (!sk[31]) & (!g1022) & (!g1023) & (g1024)) + ((g131) & (g1021) & (!sk[31]) & (!g1022) & (g1023) & (!g1024)) + ((g131) & (g1021) & (!sk[31]) & (!g1022) & (g1023) & (g1024)) + ((g131) & (g1021) & (!sk[31]) & (g1022) & (!g1023) & (!g1024)) + ((g131) & (g1021) & (!sk[31]) & (g1022) & (!g1023) & (g1024)) + ((g131) & (g1021) & (!sk[31]) & (g1022) & (g1023) & (!g1024)) + ((g131) & (g1021) & (!sk[31]) & (g1022) & (g1023) & (g1024)) + ((g131) & (g1021) & (sk[31]) & (!g1022) & (!g1023) & (!g1024)));
	assign g1026 = (((!sk[32]) & (!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[32]) & (!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[32]) & (!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g112)) + ((!sk[32]) & (!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g112)) + ((!sk[32]) & (!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((!sk[32]) & (!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g112)) + ((!sk[32]) & (!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g112)) + ((!sk[32]) & (!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g112)) + ((!sk[32]) & (!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[32]) & (!i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[32]) & (!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g112)) + ((!sk[32]) & (i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[32]) & (i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[32]) & (i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g112)) + ((!sk[32]) & (i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g112)) + ((!sk[32]) & (i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((!sk[32]) & (i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g112)) + ((!sk[32]) & (i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g112)) + ((!sk[32]) & (i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g112)) + ((!sk[32]) & (i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[32]) & (i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[32]) & (i_15_) & (i_12_) & (i_13_) & (i_14_) & (g112)) + ((sk[32]) & (!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((sk[32]) & (!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112)) + ((sk[32]) & (!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g112)) + ((sk[32]) & (i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((sk[32]) & (i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((sk[32]) & (i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112)));
	assign g1027 = (((!i_12_) & (!i_13_) & (i_14_) & (!g107) & (!g91) & (!g131)) + ((!i_12_) & (!i_13_) & (i_14_) & (!g107) & (g91) & (!g131)) + ((!i_12_) & (!i_13_) & (i_14_) & (g107) & (!g91) & (!g131)) + ((!i_12_) & (i_13_) & (i_14_) & (!g107) & (!g91) & (!g131)) + ((!i_12_) & (i_13_) & (i_14_) & (!g107) & (g91) & (!g131)) + ((!i_12_) & (i_13_) & (i_14_) & (g107) & (!g91) & (!g131)) + ((i_12_) & (!i_13_) & (i_14_) & (!g107) & (!g91) & (!g131)) + ((i_12_) & (!i_13_) & (i_14_) & (g107) & (!g91) & (!g131)) + ((i_12_) & (i_13_) & (!i_14_) & (!g107) & (!g91) & (!g131)) + ((i_12_) & (i_13_) & (!i_14_) & (g107) & (!g91) & (!g131)) + ((i_12_) & (i_13_) & (i_14_) & (!g107) & (!g91) & (!g131)) + ((i_12_) & (i_13_) & (i_14_) & (!g107) & (g91) & (!g131)));
	assign g1028 = (((!sk[34]) & (!g107) & (!g460) & (g640)) + ((!sk[34]) & (!g107) & (g460) & (!g640)) + ((!sk[34]) & (!g107) & (g460) & (g640)) + ((!sk[34]) & (g107) & (!g460) & (g640)) + ((!sk[34]) & (g107) & (g460) & (!g640)) + ((!sk[34]) & (g107) & (g460) & (g640)) + ((sk[34]) & (!g107) & (g460) & (!g640)) + ((sk[34]) & (g107) & (!g460) & (!g640)) + ((sk[34]) & (g107) & (g460) & (!g640)));
	assign g1029 = (((!g4) & (!g107) & (!sk[35]) & (g176) & (!g652)) + ((!g4) & (!g107) & (!sk[35]) & (g176) & (g652)) + ((!g4) & (!g107) & (sk[35]) & (g176) & (!g652)) + ((!g4) & (g107) & (!sk[35]) & (g176) & (!g652)) + ((!g4) & (g107) & (!sk[35]) & (g176) & (g652)) + ((!g4) & (g107) & (sk[35]) & (!g176) & (!g652)) + ((!g4) & (g107) & (sk[35]) & (g176) & (!g652)) + ((g4) & (!g107) & (!sk[35]) & (g176) & (!g652)) + ((g4) & (!g107) & (!sk[35]) & (g176) & (g652)) + ((g4) & (g107) & (!sk[35]) & (g176) & (!g652)) + ((g4) & (g107) & (!sk[35]) & (g176) & (g652)) + ((g4) & (g107) & (sk[35]) & (!g176) & (!g652)) + ((g4) & (g107) & (sk[35]) & (g176) & (!g652)));
	assign g1030 = (((!g125) & (!g296) & (g651) & (!g1028) & (!sk[36]) & (g1029)) + ((!g125) & (!g296) & (g651) & (g1028) & (!sk[36]) & (!g1029)) + ((!g125) & (!g296) & (g651) & (g1028) & (!sk[36]) & (g1029)) + ((!g125) & (g296) & (!g651) & (!g1028) & (!sk[36]) & (!g1029)) + ((!g125) & (g296) & (!g651) & (!g1028) & (!sk[36]) & (g1029)) + ((!g125) & (g296) & (!g651) & (g1028) & (!sk[36]) & (!g1029)) + ((!g125) & (g296) & (!g651) & (g1028) & (!sk[36]) & (g1029)) + ((!g125) & (g296) & (g651) & (!g1028) & (!sk[36]) & (!g1029)) + ((!g125) & (g296) & (g651) & (!g1028) & (!sk[36]) & (g1029)) + ((!g125) & (g296) & (g651) & (g1028) & (!sk[36]) & (!g1029)) + ((!g125) & (g296) & (g651) & (g1028) & (!sk[36]) & (g1029)) + ((g125) & (!g296) & (!g651) & (!g1028) & (sk[36]) & (!g1029)) + ((g125) & (!g296) & (!g651) & (!g1028) & (sk[36]) & (g1029)) + ((g125) & (!g296) & (!g651) & (g1028) & (sk[36]) & (!g1029)) + ((g125) & (!g296) & (g651) & (!g1028) & (!sk[36]) & (g1029)) + ((g125) & (!g296) & (g651) & (!g1028) & (sk[36]) & (!g1029)) + ((g125) & (!g296) & (g651) & (!g1028) & (sk[36]) & (g1029)) + ((g125) & (!g296) & (g651) & (g1028) & (!sk[36]) & (!g1029)) + ((g125) & (!g296) & (g651) & (g1028) & (!sk[36]) & (g1029)) + ((g125) & (!g296) & (g651) & (g1028) & (sk[36]) & (!g1029)) + ((g125) & (!g296) & (g651) & (g1028) & (sk[36]) & (g1029)) + ((g125) & (g296) & (!g651) & (!g1028) & (!sk[36]) & (!g1029)) + ((g125) & (g296) & (!g651) & (!g1028) & (!sk[36]) & (g1029)) + ((g125) & (g296) & (!g651) & (!g1028) & (sk[36]) & (!g1029)) + ((g125) & (g296) & (!g651) & (!g1028) & (sk[36]) & (g1029)) + ((g125) & (g296) & (!g651) & (g1028) & (!sk[36]) & (!g1029)) + ((g125) & (g296) & (!g651) & (g1028) & (!sk[36]) & (g1029)) + ((g125) & (g296) & (!g651) & (g1028) & (sk[36]) & (!g1029)) + ((g125) & (g296) & (!g651) & (g1028) & (sk[36]) & (g1029)) + ((g125) & (g296) & (g651) & (!g1028) & (!sk[36]) & (!g1029)) + ((g125) & (g296) & (g651) & (!g1028) & (!sk[36]) & (g1029)) + ((g125) & (g296) & (g651) & (!g1028) & (sk[36]) & (!g1029)) + ((g125) & (g296) & (g651) & (!g1028) & (sk[36]) & (g1029)) + ((g125) & (g296) & (g651) & (g1028) & (!sk[36]) & (!g1029)) + ((g125) & (g296) & (g651) & (g1028) & (!sk[36]) & (g1029)) + ((g125) & (g296) & (g651) & (g1028) & (sk[36]) & (!g1029)) + ((g125) & (g296) & (g651) & (g1028) & (sk[36]) & (g1029)));
	assign g1031 = (((!sk[37]) & (!g125) & (!g1026) & (g1027) & (!g1030)) + ((!sk[37]) & (!g125) & (!g1026) & (g1027) & (g1030)) + ((!sk[37]) & (!g125) & (g1026) & (g1027) & (!g1030)) + ((!sk[37]) & (!g125) & (g1026) & (g1027) & (g1030)) + ((!sk[37]) & (g125) & (!g1026) & (g1027) & (!g1030)) + ((!sk[37]) & (g125) & (!g1026) & (g1027) & (g1030)) + ((!sk[37]) & (g125) & (g1026) & (g1027) & (!g1030)) + ((!sk[37]) & (g125) & (g1026) & (g1027) & (g1030)) + ((sk[37]) & (!g125) & (!g1026) & (!g1027) & (!g1030)) + ((sk[37]) & (!g125) & (g1026) & (!g1027) & (!g1030)) + ((sk[37]) & (g125) & (!g1026) & (!g1027) & (!g1030)));
	assign g1032 = (((!sk[38]) & (!g20) & (!g496) & (g522) & (!g735) & (g847)) + ((!sk[38]) & (!g20) & (!g496) & (g522) & (g735) & (!g847)) + ((!sk[38]) & (!g20) & (!g496) & (g522) & (g735) & (g847)) + ((!sk[38]) & (!g20) & (g496) & (!g522) & (!g735) & (!g847)) + ((!sk[38]) & (!g20) & (g496) & (!g522) & (!g735) & (g847)) + ((!sk[38]) & (!g20) & (g496) & (!g522) & (g735) & (!g847)) + ((!sk[38]) & (!g20) & (g496) & (!g522) & (g735) & (g847)) + ((!sk[38]) & (!g20) & (g496) & (g522) & (!g735) & (!g847)) + ((!sk[38]) & (!g20) & (g496) & (g522) & (!g735) & (g847)) + ((!sk[38]) & (!g20) & (g496) & (g522) & (g735) & (!g847)) + ((!sk[38]) & (!g20) & (g496) & (g522) & (g735) & (g847)) + ((!sk[38]) & (g20) & (!g496) & (g522) & (!g735) & (g847)) + ((!sk[38]) & (g20) & (!g496) & (g522) & (g735) & (!g847)) + ((!sk[38]) & (g20) & (!g496) & (g522) & (g735) & (g847)) + ((!sk[38]) & (g20) & (g496) & (!g522) & (!g735) & (!g847)) + ((!sk[38]) & (g20) & (g496) & (!g522) & (!g735) & (g847)) + ((!sk[38]) & (g20) & (g496) & (!g522) & (g735) & (!g847)) + ((!sk[38]) & (g20) & (g496) & (!g522) & (g735) & (g847)) + ((!sk[38]) & (g20) & (g496) & (g522) & (!g735) & (!g847)) + ((!sk[38]) & (g20) & (g496) & (g522) & (!g735) & (g847)) + ((!sk[38]) & (g20) & (g496) & (g522) & (g735) & (!g847)) + ((!sk[38]) & (g20) & (g496) & (g522) & (g735) & (g847)) + ((sk[38]) & (!g20) & (!g496) & (!g522) & (!g735) & (g847)) + ((sk[38]) & (!g20) & (!g496) & (!g522) & (g735) & (g847)) + ((sk[38]) & (g20) & (!g496) & (!g522) & (!g735) & (g847)));
	assign g1033 = (((!sk[39]) & (!g508) & (!g514) & (g852)) + ((!sk[39]) & (!g508) & (g514) & (!g852)) + ((!sk[39]) & (!g508) & (g514) & (g852)) + ((!sk[39]) & (g508) & (!g514) & (g852)) + ((!sk[39]) & (g508) & (g514) & (!g852)) + ((!sk[39]) & (g508) & (g514) & (g852)) + ((sk[39]) & (!g508) & (!g514) & (!g852)));
	assign g1034 = (((!i_12_) & (!i_14_) & (!g88) & (sk[40]) & (!g477)) + ((!i_12_) & (!i_14_) & (g88) & (!sk[40]) & (!g477)) + ((!i_12_) & (!i_14_) & (g88) & (!sk[40]) & (g477)) + ((!i_12_) & (!i_14_) & (g88) & (sk[40]) & (!g477)) + ((!i_12_) & (i_14_) & (!g88) & (sk[40]) & (!g477)) + ((!i_12_) & (i_14_) & (g88) & (!sk[40]) & (!g477)) + ((!i_12_) & (i_14_) & (g88) & (!sk[40]) & (g477)) + ((!i_12_) & (i_14_) & (g88) & (sk[40]) & (!g477)) + ((i_12_) & (!i_14_) & (!g88) & (sk[40]) & (!g477)) + ((i_12_) & (!i_14_) & (g88) & (!sk[40]) & (!g477)) + ((i_12_) & (!i_14_) & (g88) & (!sk[40]) & (g477)) + ((i_12_) & (i_14_) & (!g88) & (sk[40]) & (!g477)) + ((i_12_) & (i_14_) & (g88) & (!sk[40]) & (!g477)) + ((i_12_) & (i_14_) & (g88) & (!sk[40]) & (g477)) + ((i_12_) & (i_14_) & (g88) & (sk[40]) & (!g477)));
	assign g1035 = (((!i_12_) & (!i_13_) & (i_14_) & (!g20) & (g27) & (!g91)) + ((!i_12_) & (!i_13_) & (i_14_) & (!g20) & (g27) & (g91)) + ((!i_12_) & (!i_13_) & (i_14_) & (g20) & (g27) & (!g91)) + ((!i_12_) & (!i_13_) & (i_14_) & (g20) & (g27) & (g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g20) & (!g27) & (!g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g20) & (g27) & (!g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g20) & (g27) & (g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (g20) & (!g27) & (!g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (g20) & (g27) & (!g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (g20) & (g27) & (g91)) + ((!i_12_) & (i_13_) & (i_14_) & (!g20) & (g27) & (!g91)) + ((!i_12_) & (i_13_) & (i_14_) & (!g20) & (g27) & (g91)) + ((!i_12_) & (i_13_) & (i_14_) & (g20) & (!g27) & (!g91)) + ((!i_12_) & (i_13_) & (i_14_) & (g20) & (!g27) & (g91)) + ((!i_12_) & (i_13_) & (i_14_) & (g20) & (g27) & (!g91)) + ((!i_12_) & (i_13_) & (i_14_) & (g20) & (g27) & (g91)) + ((i_12_) & (!i_13_) & (!i_14_) & (!g20) & (g27) & (!g91)) + ((i_12_) & (!i_13_) & (!i_14_) & (!g20) & (g27) & (g91)) + ((i_12_) & (!i_13_) & (!i_14_) & (g20) & (g27) & (!g91)) + ((i_12_) & (!i_13_) & (!i_14_) & (g20) & (g27) & (g91)) + ((i_12_) & (i_13_) & (!i_14_) & (!g20) & (g27) & (!g91)) + ((i_12_) & (i_13_) & (!i_14_) & (!g20) & (g27) & (g91)) + ((i_12_) & (i_13_) & (!i_14_) & (g20) & (g27) & (!g91)) + ((i_12_) & (i_13_) & (!i_14_) & (g20) & (g27) & (g91)) + ((i_12_) & (i_13_) & (i_14_) & (!g20) & (!g27) & (!g91)) + ((i_12_) & (i_13_) & (i_14_) & (!g20) & (g27) & (!g91)) + ((i_12_) & (i_13_) & (i_14_) & (!g20) & (g27) & (g91)) + ((i_12_) & (i_13_) & (i_14_) & (g20) & (!g27) & (!g91)) + ((i_12_) & (i_13_) & (i_14_) & (g20) & (!g27) & (g91)) + ((i_12_) & (i_13_) & (i_14_) & (g20) & (g27) & (!g91)) + ((i_12_) & (i_13_) & (i_14_) & (g20) & (g27) & (g91)));
	assign g1036 = (((!g725) & (!g1032) & (!sk[42]) & (g1033) & (!g1034) & (g1035)) + ((!g725) & (!g1032) & (!sk[42]) & (g1033) & (g1034) & (!g1035)) + ((!g725) & (!g1032) & (!sk[42]) & (g1033) & (g1034) & (g1035)) + ((!g725) & (g1032) & (!sk[42]) & (!g1033) & (!g1034) & (!g1035)) + ((!g725) & (g1032) & (!sk[42]) & (!g1033) & (!g1034) & (g1035)) + ((!g725) & (g1032) & (!sk[42]) & (!g1033) & (g1034) & (!g1035)) + ((!g725) & (g1032) & (!sk[42]) & (!g1033) & (g1034) & (g1035)) + ((!g725) & (g1032) & (!sk[42]) & (g1033) & (!g1034) & (!g1035)) + ((!g725) & (g1032) & (!sk[42]) & (g1033) & (!g1034) & (g1035)) + ((!g725) & (g1032) & (!sk[42]) & (g1033) & (g1034) & (!g1035)) + ((!g725) & (g1032) & (!sk[42]) & (g1033) & (g1034) & (g1035)) + ((g725) & (!g1032) & (!sk[42]) & (g1033) & (!g1034) & (g1035)) + ((g725) & (!g1032) & (!sk[42]) & (g1033) & (g1034) & (!g1035)) + ((g725) & (!g1032) & (!sk[42]) & (g1033) & (g1034) & (g1035)) + ((g725) & (g1032) & (!sk[42]) & (!g1033) & (!g1034) & (!g1035)) + ((g725) & (g1032) & (!sk[42]) & (!g1033) & (!g1034) & (g1035)) + ((g725) & (g1032) & (!sk[42]) & (!g1033) & (g1034) & (!g1035)) + ((g725) & (g1032) & (!sk[42]) & (!g1033) & (g1034) & (g1035)) + ((g725) & (g1032) & (!sk[42]) & (g1033) & (!g1034) & (!g1035)) + ((g725) & (g1032) & (!sk[42]) & (g1033) & (!g1034) & (g1035)) + ((g725) & (g1032) & (!sk[42]) & (g1033) & (g1034) & (!g1035)) + ((g725) & (g1032) & (!sk[42]) & (g1033) & (g1034) & (g1035)) + ((g725) & (g1032) & (sk[42]) & (g1033) & (g1034) & (!g1035)));
	assign g1037 = (((!i_12_) & (!i_13_) & (!sk[43]) & (i_14_) & (!g86) & (g83)) + ((!i_12_) & (!i_13_) & (!sk[43]) & (i_14_) & (g86) & (!g83)) + ((!i_12_) & (!i_13_) & (!sk[43]) & (i_14_) & (g86) & (g83)) + ((!i_12_) & (!i_13_) & (sk[43]) & (!i_14_) & (!g86) & (g83)) + ((!i_12_) & (!i_13_) & (sk[43]) & (!i_14_) & (g86) & (g83)) + ((!i_12_) & (!i_13_) & (sk[43]) & (i_14_) & (!g86) & (g83)) + ((!i_12_) & (!i_13_) & (sk[43]) & (i_14_) & (g86) & (g83)) + ((!i_12_) & (i_13_) & (!sk[43]) & (!i_14_) & (!g86) & (!g83)) + ((!i_12_) & (i_13_) & (!sk[43]) & (!i_14_) & (!g86) & (g83)) + ((!i_12_) & (i_13_) & (!sk[43]) & (!i_14_) & (g86) & (!g83)) + ((!i_12_) & (i_13_) & (!sk[43]) & (!i_14_) & (g86) & (g83)) + ((!i_12_) & (i_13_) & (!sk[43]) & (i_14_) & (!g86) & (!g83)) + ((!i_12_) & (i_13_) & (!sk[43]) & (i_14_) & (!g86) & (g83)) + ((!i_12_) & (i_13_) & (!sk[43]) & (i_14_) & (g86) & (!g83)) + ((!i_12_) & (i_13_) & (!sk[43]) & (i_14_) & (g86) & (g83)) + ((!i_12_) & (i_13_) & (sk[43]) & (i_14_) & (!g86) & (g83)) + ((!i_12_) & (i_13_) & (sk[43]) & (i_14_) & (g86) & (g83)) + ((i_12_) & (!i_13_) & (!sk[43]) & (i_14_) & (!g86) & (g83)) + ((i_12_) & (!i_13_) & (!sk[43]) & (i_14_) & (g86) & (!g83)) + ((i_12_) & (!i_13_) & (!sk[43]) & (i_14_) & (g86) & (g83)) + ((i_12_) & (i_13_) & (!sk[43]) & (!i_14_) & (!g86) & (!g83)) + ((i_12_) & (i_13_) & (!sk[43]) & (!i_14_) & (!g86) & (g83)) + ((i_12_) & (i_13_) & (!sk[43]) & (!i_14_) & (g86) & (!g83)) + ((i_12_) & (i_13_) & (!sk[43]) & (!i_14_) & (g86) & (g83)) + ((i_12_) & (i_13_) & (!sk[43]) & (i_14_) & (!g86) & (!g83)) + ((i_12_) & (i_13_) & (!sk[43]) & (i_14_) & (!g86) & (g83)) + ((i_12_) & (i_13_) & (!sk[43]) & (i_14_) & (g86) & (!g83)) + ((i_12_) & (i_13_) & (!sk[43]) & (i_14_) & (g86) & (g83)) + ((i_12_) & (i_13_) & (sk[43]) & (!i_14_) & (g86) & (!g83)) + ((i_12_) & (i_13_) & (sk[43]) & (!i_14_) & (g86) & (g83)));
	assign g1038 = (((!g629) & (!sk[44]) & (!g703) & (g851) & (!g1037)) + ((!g629) & (!sk[44]) & (!g703) & (g851) & (g1037)) + ((!g629) & (!sk[44]) & (g703) & (g851) & (!g1037)) + ((!g629) & (!sk[44]) & (g703) & (g851) & (g1037)) + ((!g629) & (sk[44]) & (g703) & (g851) & (!g1037)) + ((g629) & (!sk[44]) & (!g703) & (g851) & (!g1037)) + ((g629) & (!sk[44]) & (!g703) & (g851) & (g1037)) + ((g629) & (!sk[44]) & (g703) & (g851) & (!g1037)) + ((g629) & (!sk[44]) & (g703) & (g851) & (g1037)));
	assign g1039 = (((!g25) & (!g358) & (g933) & (!sk[45]) & (!g1038)) + ((!g25) & (!g358) & (g933) & (!sk[45]) & (g1038)) + ((!g25) & (g358) & (g933) & (!sk[45]) & (!g1038)) + ((!g25) & (g358) & (g933) & (!sk[45]) & (g1038)) + ((g25) & (!g358) & (g933) & (!sk[45]) & (!g1038)) + ((g25) & (!g358) & (g933) & (!sk[45]) & (g1038)) + ((g25) & (!g358) & (g933) & (sk[45]) & (g1038)) + ((g25) & (g358) & (g933) & (!sk[45]) & (!g1038)) + ((g25) & (g358) & (g933) & (!sk[45]) & (g1038)));
	assign g1040 = (((!i_8_) & (!sk[46]) & (!g144) & (g898) & (!g1036) & (g1039)) + ((!i_8_) & (!sk[46]) & (!g144) & (g898) & (g1036) & (!g1039)) + ((!i_8_) & (!sk[46]) & (!g144) & (g898) & (g1036) & (g1039)) + ((!i_8_) & (!sk[46]) & (g144) & (!g898) & (!g1036) & (!g1039)) + ((!i_8_) & (!sk[46]) & (g144) & (!g898) & (!g1036) & (g1039)) + ((!i_8_) & (!sk[46]) & (g144) & (!g898) & (g1036) & (!g1039)) + ((!i_8_) & (!sk[46]) & (g144) & (!g898) & (g1036) & (g1039)) + ((!i_8_) & (!sk[46]) & (g144) & (g898) & (!g1036) & (!g1039)) + ((!i_8_) & (!sk[46]) & (g144) & (g898) & (!g1036) & (g1039)) + ((!i_8_) & (!sk[46]) & (g144) & (g898) & (g1036) & (!g1039)) + ((!i_8_) & (!sk[46]) & (g144) & (g898) & (g1036) & (g1039)) + ((!i_8_) & (sk[46]) & (g144) & (!g898) & (!g1036) & (!g1039)) + ((!i_8_) & (sk[46]) & (g144) & (!g898) & (!g1036) & (g1039)) + ((!i_8_) & (sk[46]) & (g144) & (!g898) & (g1036) & (!g1039)) + ((!i_8_) & (sk[46]) & (g144) & (g898) & (!g1036) & (!g1039)) + ((!i_8_) & (sk[46]) & (g144) & (g898) & (!g1036) & (g1039)) + ((!i_8_) & (sk[46]) & (g144) & (g898) & (g1036) & (!g1039)) + ((i_8_) & (!sk[46]) & (!g144) & (g898) & (!g1036) & (g1039)) + ((i_8_) & (!sk[46]) & (!g144) & (g898) & (g1036) & (!g1039)) + ((i_8_) & (!sk[46]) & (!g144) & (g898) & (g1036) & (g1039)) + ((i_8_) & (!sk[46]) & (g144) & (!g898) & (!g1036) & (!g1039)) + ((i_8_) & (!sk[46]) & (g144) & (!g898) & (!g1036) & (g1039)) + ((i_8_) & (!sk[46]) & (g144) & (!g898) & (g1036) & (!g1039)) + ((i_8_) & (!sk[46]) & (g144) & (!g898) & (g1036) & (g1039)) + ((i_8_) & (!sk[46]) & (g144) & (g898) & (!g1036) & (!g1039)) + ((i_8_) & (!sk[46]) & (g144) & (g898) & (!g1036) & (g1039)) + ((i_8_) & (!sk[46]) & (g144) & (g898) & (g1036) & (!g1039)) + ((i_8_) & (!sk[46]) & (g144) & (g898) & (g1036) & (g1039)) + ((i_8_) & (sk[46]) & (g144) & (!g898) & (!g1036) & (!g1039)) + ((i_8_) & (sk[46]) & (g144) & (!g898) & (!g1036) & (g1039)) + ((i_8_) & (sk[46]) & (g144) & (!g898) & (g1036) & (!g1039)));
	assign g1041 = (((g761) & (!sk[47]) & (!g945)) + ((g761) & (!sk[47]) & (g945)) + ((g761) & (sk[47]) & (g945)));
	assign g1042 = (((!sk[48]) & (!g125) & (!g144) & (g851) & (!g1041)) + ((!sk[48]) & (!g125) & (!g144) & (g851) & (g1041)) + ((!sk[48]) & (!g125) & (g144) & (g851) & (!g1041)) + ((!sk[48]) & (!g125) & (g144) & (g851) & (g1041)) + ((!sk[48]) & (g125) & (!g144) & (g851) & (!g1041)) + ((!sk[48]) & (g125) & (!g144) & (g851) & (g1041)) + ((!sk[48]) & (g125) & (g144) & (g851) & (!g1041)) + ((!sk[48]) & (g125) & (g144) & (g851) & (g1041)) + ((sk[48]) & (!g125) & (g144) & (!g851) & (!g1041)) + ((sk[48]) & (!g125) & (g144) & (g851) & (!g1041)) + ((sk[48]) & (g125) & (!g144) & (!g851) & (!g1041)) + ((sk[48]) & (g125) & (!g144) & (!g851) & (g1041)) + ((sk[48]) & (g125) & (g144) & (!g851) & (!g1041)) + ((sk[48]) & (g125) & (g144) & (!g851) & (g1041)) + ((sk[48]) & (g125) & (g144) & (g851) & (!g1041)));
	assign g1043 = (((!sk[49]) & (!g317) & (!g318) & (g319) & (!g320)) + ((!sk[49]) & (!g317) & (!g318) & (g319) & (g320)) + ((!sk[49]) & (!g317) & (g318) & (g319) & (!g320)) + ((!sk[49]) & (!g317) & (g318) & (g319) & (g320)) + ((!sk[49]) & (g317) & (!g318) & (g319) & (!g320)) + ((!sk[49]) & (g317) & (!g318) & (g319) & (g320)) + ((!sk[49]) & (g317) & (g318) & (g319) & (!g320)) + ((!sk[49]) & (g317) & (g318) & (g319) & (g320)) + ((sk[49]) & (!g317) & (!g318) & (!g319) & (!g320)));
	assign g1044 = (((!sk[50]) & (!g355) & (!g35) & (g460) & (!g641)) + ((!sk[50]) & (!g355) & (!g35) & (g460) & (g641)) + ((!sk[50]) & (!g355) & (g35) & (g460) & (!g641)) + ((!sk[50]) & (!g355) & (g35) & (g460) & (g641)) + ((!sk[50]) & (g355) & (!g35) & (g460) & (!g641)) + ((!sk[50]) & (g355) & (!g35) & (g460) & (g641)) + ((!sk[50]) & (g355) & (g35) & (g460) & (!g641)) + ((!sk[50]) & (g355) & (g35) & (g460) & (g641)) + ((sk[50]) & (!g355) & (!g35) & (!g460) & (!g641)) + ((sk[50]) & (!g355) & (!g35) & (g460) & (!g641)) + ((sk[50]) & (!g355) & (g35) & (g460) & (!g641)) + ((sk[50]) & (g355) & (!g35) & (!g460) & (!g641)) + ((sk[50]) & (g355) & (!g35) & (g460) & (!g641)));
	assign g1045 = (((!sk[51]) & (!g125) & (!g131) & (g487) & (!g948) & (g1044)) + ((!sk[51]) & (!g125) & (!g131) & (g487) & (g948) & (!g1044)) + ((!sk[51]) & (!g125) & (!g131) & (g487) & (g948) & (g1044)) + ((!sk[51]) & (!g125) & (g131) & (!g487) & (!g948) & (!g1044)) + ((!sk[51]) & (!g125) & (g131) & (!g487) & (!g948) & (g1044)) + ((!sk[51]) & (!g125) & (g131) & (!g487) & (g948) & (!g1044)) + ((!sk[51]) & (!g125) & (g131) & (!g487) & (g948) & (g1044)) + ((!sk[51]) & (!g125) & (g131) & (g487) & (!g948) & (!g1044)) + ((!sk[51]) & (!g125) & (g131) & (g487) & (!g948) & (g1044)) + ((!sk[51]) & (!g125) & (g131) & (g487) & (g948) & (!g1044)) + ((!sk[51]) & (!g125) & (g131) & (g487) & (g948) & (g1044)) + ((!sk[51]) & (g125) & (!g131) & (g487) & (!g948) & (g1044)) + ((!sk[51]) & (g125) & (!g131) & (g487) & (g948) & (!g1044)) + ((!sk[51]) & (g125) & (!g131) & (g487) & (g948) & (g1044)) + ((!sk[51]) & (g125) & (g131) & (!g487) & (!g948) & (!g1044)) + ((!sk[51]) & (g125) & (g131) & (!g487) & (!g948) & (g1044)) + ((!sk[51]) & (g125) & (g131) & (!g487) & (g948) & (!g1044)) + ((!sk[51]) & (g125) & (g131) & (!g487) & (g948) & (g1044)) + ((!sk[51]) & (g125) & (g131) & (g487) & (!g948) & (!g1044)) + ((!sk[51]) & (g125) & (g131) & (g487) & (!g948) & (g1044)) + ((!sk[51]) & (g125) & (g131) & (g487) & (g948) & (!g1044)) + ((!sk[51]) & (g125) & (g131) & (g487) & (g948) & (g1044)) + ((sk[51]) & (!g125) & (!g131) & (!g487) & (g948) & (g1044)) + ((sk[51]) & (!g125) & (!g131) & (g487) & (g948) & (g1044)) + ((sk[51]) & (!g125) & (g131) & (!g487) & (!g948) & (!g1044)) + ((sk[51]) & (!g125) & (g131) & (!g487) & (!g948) & (g1044)) + ((sk[51]) & (!g125) & (g131) & (!g487) & (g948) & (!g1044)) + ((sk[51]) & (!g125) & (g131) & (!g487) & (g948) & (g1044)) + ((sk[51]) & (!g125) & (g131) & (g487) & (!g948) & (!g1044)) + ((sk[51]) & (!g125) & (g131) & (g487) & (!g948) & (g1044)) + ((sk[51]) & (!g125) & (g131) & (g487) & (g948) & (!g1044)) + ((sk[51]) & (!g125) & (g131) & (g487) & (g948) & (g1044)) + ((sk[51]) & (g125) & (!g131) & (!g487) & (g948) & (g1044)) + ((sk[51]) & (g125) & (g131) & (!g487) & (!g948) & (!g1044)) + ((sk[51]) & (g125) & (g131) & (!g487) & (!g948) & (g1044)) + ((sk[51]) & (g125) & (g131) & (!g487) & (g948) & (!g1044)) + ((sk[51]) & (g125) & (g131) & (!g487) & (g948) & (g1044)));
	assign g1046 = (((!i_12_) & (!i_13_) & (!i_14_) & (g17) & (!g27) & (g125)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g17) & (g27) & (g125)) + ((!i_12_) & (!i_13_) & (i_14_) & (!g17) & (g27) & (g125)) + ((!i_12_) & (!i_13_) & (i_14_) & (g17) & (!g27) & (g125)) + ((!i_12_) & (!i_13_) & (i_14_) & (g17) & (g27) & (g125)) + ((!i_12_) & (i_13_) & (i_14_) & (!g17) & (g27) & (g125)) + ((!i_12_) & (i_13_) & (i_14_) & (g17) & (!g27) & (g125)) + ((!i_12_) & (i_13_) & (i_14_) & (g17) & (g27) & (g125)) + ((i_12_) & (!i_13_) & (!i_14_) & (g17) & (!g27) & (g125)) + ((i_12_) & (!i_13_) & (!i_14_) & (g17) & (g27) & (g125)) + ((i_12_) & (i_13_) & (!i_14_) & (!g17) & (g27) & (g125)) + ((i_12_) & (i_13_) & (!i_14_) & (g17) & (!g27) & (g125)) + ((i_12_) & (i_13_) & (!i_14_) & (g17) & (g27) & (g125)) + ((i_12_) & (i_13_) & (i_14_) & (!g17) & (g27) & (g125)) + ((i_12_) & (i_13_) & (i_14_) & (g17) & (g27) & (g125)));
	assign g1047 = (((!g125) & (!g79) & (g625) & (!sk[53]) & (!g931)) + ((!g125) & (!g79) & (g625) & (!sk[53]) & (g931)) + ((!g125) & (g79) & (g625) & (!sk[53]) & (!g931)) + ((!g125) & (g79) & (g625) & (!sk[53]) & (g931)) + ((g125) & (!g79) & (!g625) & (sk[53]) & (!g931)) + ((g125) & (!g79) & (!g625) & (sk[53]) & (g931)) + ((g125) & (!g79) & (g625) & (!sk[53]) & (!g931)) + ((g125) & (!g79) & (g625) & (!sk[53]) & (g931)) + ((g125) & (!g79) & (g625) & (sk[53]) & (!g931)) + ((g125) & (!g79) & (g625) & (sk[53]) & (g931)) + ((g125) & (g79) & (!g625) & (sk[53]) & (g931)) + ((g125) & (g79) & (g625) & (!sk[53]) & (!g931)) + ((g125) & (g79) & (g625) & (!sk[53]) & (g931)) + ((g125) & (g79) & (g625) & (sk[53]) & (!g931)) + ((g125) & (g79) & (g625) & (sk[53]) & (g931)));
	assign g1048 = (((!i_12_) & (!i_13_) & (!i_14_) & (!g35) & (g36) & (g125)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g35) & (g36) & (g125)) + ((!i_12_) & (!i_13_) & (i_14_) & (!g35) & (g36) & (g125)) + ((!i_12_) & (!i_13_) & (i_14_) & (g35) & (g36) & (g125)) + ((!i_12_) & (i_13_) & (i_14_) & (!g35) & (g36) & (g125)) + ((!i_12_) & (i_13_) & (i_14_) & (g35) & (g36) & (g125)) + ((i_12_) & (!i_13_) & (!i_14_) & (!g35) & (g36) & (g125)) + ((i_12_) & (!i_13_) & (!i_14_) & (g35) & (g36) & (g125)) + ((i_12_) & (i_13_) & (!i_14_) & (g35) & (!g36) & (g125)) + ((i_12_) & (i_13_) & (!i_14_) & (g35) & (g36) & (g125)) + ((i_12_) & (i_13_) & (i_14_) & (g35) & (!g36) & (g125)) + ((i_12_) & (i_13_) & (i_14_) & (g35) & (g36) & (g125)));
	assign g1049 = (((!i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (g429) & (g125)) + ((!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g429) & (g125)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g429) & (g125)) + ((!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g429) & (g125)) + ((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g429) & (g125)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g429) & (g125)) + ((i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (g429) & (g125)) + ((i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g429) & (g125)) + ((i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g429) & (g125)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g429) & (g125)) + ((i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g429) & (g125)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g429) & (g125)) + ((i_15_) & (i_12_) & (i_13_) & (i_14_) & (g429) & (g125)));
	assign g1050 = (((!sk[56]) & (!g125) & (!g282) & (g552) & (!g668) & (g698)) + ((!sk[56]) & (!g125) & (!g282) & (g552) & (g668) & (!g698)) + ((!sk[56]) & (!g125) & (!g282) & (g552) & (g668) & (g698)) + ((!sk[56]) & (!g125) & (g282) & (!g552) & (!g668) & (!g698)) + ((!sk[56]) & (!g125) & (g282) & (!g552) & (!g668) & (g698)) + ((!sk[56]) & (!g125) & (g282) & (!g552) & (g668) & (!g698)) + ((!sk[56]) & (!g125) & (g282) & (!g552) & (g668) & (g698)) + ((!sk[56]) & (!g125) & (g282) & (g552) & (!g668) & (!g698)) + ((!sk[56]) & (!g125) & (g282) & (g552) & (!g668) & (g698)) + ((!sk[56]) & (!g125) & (g282) & (g552) & (g668) & (!g698)) + ((!sk[56]) & (!g125) & (g282) & (g552) & (g668) & (g698)) + ((!sk[56]) & (g125) & (!g282) & (g552) & (!g668) & (g698)) + ((!sk[56]) & (g125) & (!g282) & (g552) & (g668) & (!g698)) + ((!sk[56]) & (g125) & (!g282) & (g552) & (g668) & (g698)) + ((!sk[56]) & (g125) & (g282) & (!g552) & (!g668) & (!g698)) + ((!sk[56]) & (g125) & (g282) & (!g552) & (!g668) & (g698)) + ((!sk[56]) & (g125) & (g282) & (!g552) & (g668) & (!g698)) + ((!sk[56]) & (g125) & (g282) & (!g552) & (g668) & (g698)) + ((!sk[56]) & (g125) & (g282) & (g552) & (!g668) & (!g698)) + ((!sk[56]) & (g125) & (g282) & (g552) & (!g668) & (g698)) + ((!sk[56]) & (g125) & (g282) & (g552) & (g668) & (!g698)) + ((!sk[56]) & (g125) & (g282) & (g552) & (g668) & (g698)) + ((sk[56]) & (g125) & (!g282) & (!g552) & (!g668) & (!g698)) + ((sk[56]) & (g125) & (!g282) & (!g552) & (!g668) & (g698)) + ((sk[56]) & (g125) & (!g282) & (!g552) & (g668) & (!g698)) + ((sk[56]) & (g125) & (!g282) & (!g552) & (g668) & (g698)) + ((sk[56]) & (g125) & (!g282) & (g552) & (!g668) & (!g698)) + ((sk[56]) & (g125) & (!g282) & (g552) & (g668) & (!g698)) + ((sk[56]) & (g125) & (!g282) & (g552) & (g668) & (g698)) + ((sk[56]) & (g125) & (g282) & (!g552) & (!g668) & (!g698)) + ((sk[56]) & (g125) & (g282) & (!g552) & (!g668) & (g698)) + ((sk[56]) & (g125) & (g282) & (!g552) & (g668) & (!g698)) + ((sk[56]) & (g125) & (g282) & (!g552) & (g668) & (g698)) + ((sk[56]) & (g125) & (g282) & (g552) & (!g668) & (!g698)) + ((sk[56]) & (g125) & (g282) & (g552) & (!g668) & (g698)) + ((sk[56]) & (g125) & (g282) & (g552) & (g668) & (!g698)) + ((sk[56]) & (g125) & (g282) & (g552) & (g668) & (g698)));
	assign g1051 = (((!g87) & (!g131) & (g342) & (!sk[57]) & (!g1028) & (g1050)) + ((!g87) & (!g131) & (g342) & (!sk[57]) & (g1028) & (!g1050)) + ((!g87) & (!g131) & (g342) & (!sk[57]) & (g1028) & (g1050)) + ((!g87) & (g131) & (!g342) & (!sk[57]) & (!g1028) & (!g1050)) + ((!g87) & (g131) & (!g342) & (!sk[57]) & (!g1028) & (g1050)) + ((!g87) & (g131) & (!g342) & (!sk[57]) & (g1028) & (!g1050)) + ((!g87) & (g131) & (!g342) & (!sk[57]) & (g1028) & (g1050)) + ((!g87) & (g131) & (!g342) & (sk[57]) & (!g1028) & (!g1050)) + ((!g87) & (g131) & (!g342) & (sk[57]) & (g1028) & (!g1050)) + ((!g87) & (g131) & (g342) & (!sk[57]) & (!g1028) & (!g1050)) + ((!g87) & (g131) & (g342) & (!sk[57]) & (!g1028) & (g1050)) + ((!g87) & (g131) & (g342) & (!sk[57]) & (g1028) & (!g1050)) + ((!g87) & (g131) & (g342) & (!sk[57]) & (g1028) & (g1050)) + ((!g87) & (g131) & (g342) & (sk[57]) & (!g1028) & (!g1050)) + ((!g87) & (g131) & (g342) & (sk[57]) & (g1028) & (!g1050)) + ((g87) & (!g131) & (!g342) & (sk[57]) & (g1028) & (!g1050)) + ((g87) & (!g131) & (g342) & (!sk[57]) & (!g1028) & (g1050)) + ((g87) & (!g131) & (g342) & (!sk[57]) & (g1028) & (!g1050)) + ((g87) & (!g131) & (g342) & (!sk[57]) & (g1028) & (g1050)) + ((g87) & (g131) & (!g342) & (!sk[57]) & (!g1028) & (!g1050)) + ((g87) & (g131) & (!g342) & (!sk[57]) & (!g1028) & (g1050)) + ((g87) & (g131) & (!g342) & (!sk[57]) & (g1028) & (!g1050)) + ((g87) & (g131) & (!g342) & (!sk[57]) & (g1028) & (g1050)) + ((g87) & (g131) & (!g342) & (sk[57]) & (!g1028) & (!g1050)) + ((g87) & (g131) & (!g342) & (sk[57]) & (g1028) & (!g1050)) + ((g87) & (g131) & (g342) & (!sk[57]) & (!g1028) & (!g1050)) + ((g87) & (g131) & (g342) & (!sk[57]) & (!g1028) & (g1050)) + ((g87) & (g131) & (g342) & (!sk[57]) & (g1028) & (!g1050)) + ((g87) & (g131) & (g342) & (!sk[57]) & (g1028) & (g1050)) + ((g87) & (g131) & (g342) & (sk[57]) & (!g1028) & (!g1050)) + ((g87) & (g131) & (g342) & (sk[57]) & (g1028) & (!g1050)));
	assign g1052 = (((!g1046) & (!g1047) & (!sk[58]) & (g1048) & (!g1049) & (g1051)) + ((!g1046) & (!g1047) & (!sk[58]) & (g1048) & (g1049) & (!g1051)) + ((!g1046) & (!g1047) & (!sk[58]) & (g1048) & (g1049) & (g1051)) + ((!g1046) & (!g1047) & (sk[58]) & (!g1048) & (!g1049) & (g1051)) + ((!g1046) & (g1047) & (!sk[58]) & (!g1048) & (!g1049) & (!g1051)) + ((!g1046) & (g1047) & (!sk[58]) & (!g1048) & (!g1049) & (g1051)) + ((!g1046) & (g1047) & (!sk[58]) & (!g1048) & (g1049) & (!g1051)) + ((!g1046) & (g1047) & (!sk[58]) & (!g1048) & (g1049) & (g1051)) + ((!g1046) & (g1047) & (!sk[58]) & (g1048) & (!g1049) & (!g1051)) + ((!g1046) & (g1047) & (!sk[58]) & (g1048) & (!g1049) & (g1051)) + ((!g1046) & (g1047) & (!sk[58]) & (g1048) & (g1049) & (!g1051)) + ((!g1046) & (g1047) & (!sk[58]) & (g1048) & (g1049) & (g1051)) + ((g1046) & (!g1047) & (!sk[58]) & (g1048) & (!g1049) & (g1051)) + ((g1046) & (!g1047) & (!sk[58]) & (g1048) & (g1049) & (!g1051)) + ((g1046) & (!g1047) & (!sk[58]) & (g1048) & (g1049) & (g1051)) + ((g1046) & (g1047) & (!sk[58]) & (!g1048) & (!g1049) & (!g1051)) + ((g1046) & (g1047) & (!sk[58]) & (!g1048) & (!g1049) & (g1051)) + ((g1046) & (g1047) & (!sk[58]) & (!g1048) & (g1049) & (!g1051)) + ((g1046) & (g1047) & (!sk[58]) & (!g1048) & (g1049) & (g1051)) + ((g1046) & (g1047) & (!sk[58]) & (g1048) & (!g1049) & (!g1051)) + ((g1046) & (g1047) & (!sk[58]) & (g1048) & (!g1049) & (g1051)) + ((g1046) & (g1047) & (!sk[58]) & (g1048) & (g1049) & (!g1051)) + ((g1046) & (g1047) & (!sk[58]) & (g1048) & (g1049) & (g1051)));
	assign g1053 = (((!g1042) & (g1043) & (!g576) & (g577) & (g1045) & (g1052)));
	assign g1054 = (((!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g125) & (g445)) + ((!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g125) & (g445)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g125) & (g445)) + ((!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g125) & (g445)) + ((!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g125) & (g445)) + ((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g125) & (g445)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g125) & (g445)) + ((i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g125) & (g445)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g125) & (g445)));
	assign g1055 = (((!g125) & (!sk[61]) & (!g504) & (g729) & (!g643) & (g1054)) + ((!g125) & (!sk[61]) & (!g504) & (g729) & (g643) & (!g1054)) + ((!g125) & (!sk[61]) & (!g504) & (g729) & (g643) & (g1054)) + ((!g125) & (!sk[61]) & (g504) & (!g729) & (!g643) & (!g1054)) + ((!g125) & (!sk[61]) & (g504) & (!g729) & (!g643) & (g1054)) + ((!g125) & (!sk[61]) & (g504) & (!g729) & (g643) & (!g1054)) + ((!g125) & (!sk[61]) & (g504) & (!g729) & (g643) & (g1054)) + ((!g125) & (!sk[61]) & (g504) & (g729) & (!g643) & (!g1054)) + ((!g125) & (!sk[61]) & (g504) & (g729) & (!g643) & (g1054)) + ((!g125) & (!sk[61]) & (g504) & (g729) & (g643) & (!g1054)) + ((!g125) & (!sk[61]) & (g504) & (g729) & (g643) & (g1054)) + ((!g125) & (sk[61]) & (!g504) & (!g729) & (!g643) & (!g1054)) + ((!g125) & (sk[61]) & (!g504) & (g729) & (!g643) & (!g1054)) + ((!g125) & (sk[61]) & (g504) & (!g729) & (!g643) & (!g1054)) + ((!g125) & (sk[61]) & (g504) & (g729) & (!g643) & (!g1054)) + ((g125) & (!sk[61]) & (!g504) & (g729) & (!g643) & (g1054)) + ((g125) & (!sk[61]) & (!g504) & (g729) & (g643) & (!g1054)) + ((g125) & (!sk[61]) & (!g504) & (g729) & (g643) & (g1054)) + ((g125) & (!sk[61]) & (g504) & (!g729) & (!g643) & (!g1054)) + ((g125) & (!sk[61]) & (g504) & (!g729) & (!g643) & (g1054)) + ((g125) & (!sk[61]) & (g504) & (!g729) & (g643) & (!g1054)) + ((g125) & (!sk[61]) & (g504) & (!g729) & (g643) & (g1054)) + ((g125) & (!sk[61]) & (g504) & (g729) & (!g643) & (!g1054)) + ((g125) & (!sk[61]) & (g504) & (g729) & (!g643) & (g1054)) + ((g125) & (!sk[61]) & (g504) & (g729) & (g643) & (!g1054)) + ((g125) & (!sk[61]) & (g504) & (g729) & (g643) & (g1054)) + ((g125) & (sk[61]) & (g504) & (g729) & (!g643) & (!g1054)));
	assign g1056 = (((!sk[62]) & (!g211) & (!g695) & (g797) & (!g1055)) + ((!sk[62]) & (!g211) & (!g695) & (g797) & (g1055)) + ((!sk[62]) & (!g211) & (g695) & (g797) & (!g1055)) + ((!sk[62]) & (!g211) & (g695) & (g797) & (g1055)) + ((!sk[62]) & (g211) & (!g695) & (g797) & (!g1055)) + ((!sk[62]) & (g211) & (!g695) & (g797) & (g1055)) + ((!sk[62]) & (g211) & (g695) & (g797) & (!g1055)) + ((!sk[62]) & (g211) & (g695) & (g797) & (g1055)) + ((sk[62]) & (g211) & (g695) & (g797) & (g1055)));
	assign g1057 = (((!g1020) & (g1025) & (g1031) & (!g1040) & (g1053) & (g1056)));
	assign g1058 = (((g2) & (!sk[64]) & (!g12)) + ((g2) & (!sk[64]) & (g12)) + ((g2) & (sk[64]) & (g12)));
	assign o_19_ = (((!i_4_) & (!sk[65]) & (!i_3_) & (i_5_) & (!g1058)) + ((!i_4_) & (!sk[65]) & (!i_3_) & (i_5_) & (g1058)) + ((!i_4_) & (!sk[65]) & (i_3_) & (i_5_) & (!g1058)) + ((!i_4_) & (!sk[65]) & (i_3_) & (i_5_) & (g1058)) + ((!i_4_) & (sk[65]) & (i_3_) & (i_5_) & (g1058)) + ((i_4_) & (!sk[65]) & (!i_3_) & (i_5_) & (!g1058)) + ((i_4_) & (!sk[65]) & (!i_3_) & (i_5_) & (g1058)) + ((i_4_) & (!sk[65]) & (i_3_) & (i_5_) & (!g1058)) + ((i_4_) & (!sk[65]) & (i_3_) & (i_5_) & (g1058)));
	assign g1060 = (((!i_4_) & (!sk[66]) & (!i_3_) & (i_5_)) + ((!i_4_) & (!sk[66]) & (i_3_) & (!i_5_)) + ((!i_4_) & (!sk[66]) & (i_3_) & (i_5_)) + ((i_4_) & (!sk[66]) & (!i_3_) & (i_5_)) + ((i_4_) & (!sk[66]) & (i_3_) & (!i_5_)) + ((i_4_) & (!sk[66]) & (i_3_) & (i_5_)) + ((i_4_) & (sk[66]) & (i_3_) & (!i_5_)));
	assign o_20_ = (((g1058) & (!sk[67]) & (!g1060)) + ((g1058) & (!sk[67]) & (g1060)) + ((g1058) & (sk[67]) & (g1060)));
	assign g1062 = (((!g6) & (!g14) & (!sk[68]) & (g101)) + ((!g6) & (g14) & (!sk[68]) & (!g101)) + ((!g6) & (g14) & (!sk[68]) & (g101)) + ((g6) & (!g14) & (!sk[68]) & (g101)) + ((g6) & (g14) & (!sk[68]) & (!g101)) + ((g6) & (g14) & (!sk[68]) & (g101)) + ((g6) & (g14) & (sk[68]) & (g101)));
	assign g1063 = (((!g18) & (!g23) & (g28) & (!sk[69]) & (!g33)) + ((!g18) & (!g23) & (g28) & (!sk[69]) & (g33)) + ((!g18) & (g23) & (!g28) & (sk[69]) & (!g33)) + ((!g18) & (g23) & (g28) & (!sk[69]) & (!g33)) + ((!g18) & (g23) & (g28) & (!sk[69]) & (g33)) + ((g18) & (!g23) & (g28) & (!sk[69]) & (!g33)) + ((g18) & (!g23) & (g28) & (!sk[69]) & (g33)) + ((g18) & (g23) & (g28) & (!sk[69]) & (!g33)) + ((g18) & (g23) & (g28) & (!sk[69]) & (g33)));
	assign g1064 = (((!g20) & (!sk[70]) & (!g56) & (g1062) & (!g1063)) + ((!g20) & (!sk[70]) & (!g56) & (g1062) & (g1063)) + ((!g20) & (!sk[70]) & (g56) & (g1062) & (!g1063)) + ((!g20) & (!sk[70]) & (g56) & (g1062) & (g1063)) + ((!g20) & (sk[70]) & (!g56) & (g1062) & (!g1063)) + ((!g20) & (sk[70]) & (g56) & (g1062) & (!g1063)) + ((g20) & (!sk[70]) & (!g56) & (g1062) & (!g1063)) + ((g20) & (!sk[70]) & (!g56) & (g1062) & (g1063)) + ((g20) & (!sk[70]) & (g56) & (g1062) & (!g1063)) + ((g20) & (!sk[70]) & (g56) & (g1062) & (g1063)) + ((g20) & (sk[70]) & (!g56) & (g1062) & (!g1063)) + ((g20) & (sk[70]) & (g56) & (g1062) & (!g1063)) + ((g20) & (sk[70]) & (g56) & (g1062) & (g1063)));
	assign g1065 = (((!i_8_) & (!sk[71]) & (!i_7_) & (g48)) + ((!i_8_) & (!sk[71]) & (i_7_) & (!g48)) + ((!i_8_) & (!sk[71]) & (i_7_) & (g48)) + ((i_8_) & (!sk[71]) & (!i_7_) & (g48)) + ((i_8_) & (!sk[71]) & (i_7_) & (!g48)) + ((i_8_) & (!sk[71]) & (i_7_) & (g48)) + ((i_8_) & (sk[71]) & (!i_7_) & (g48)));
	assign o_21_ = (((!sk[72]) & (!g55) & (!g1064) & (g1065)) + ((!sk[72]) & (!g55) & (g1064) & (!g1065)) + ((!sk[72]) & (!g55) & (g1064) & (g1065)) + ((!sk[72]) & (g55) & (!g1064) & (g1065)) + ((!sk[72]) & (g55) & (g1064) & (!g1065)) + ((!sk[72]) & (g55) & (g1064) & (g1065)) + ((sk[72]) & (!g55) & (g1064) & (!g1065)) + ((sk[72]) & (!g55) & (g1064) & (g1065)) + ((sk[72]) & (g55) & (!g1064) & (g1065)) + ((sk[72]) & (g55) & (g1064) & (!g1065)) + ((sk[72]) & (g55) & (g1064) & (g1065)));
	assign g1067 = (((!sk[73]) & (!g26) & (!g28) & (g33)) + ((!sk[73]) & (!g26) & (g28) & (!g33)) + ((!sk[73]) & (!g26) & (g28) & (g33)) + ((!sk[73]) & (g26) & (!g28) & (g33)) + ((!sk[73]) & (g26) & (g28) & (!g33)) + ((!sk[73]) & (g26) & (g28) & (g33)) + ((sk[73]) & (g26) & (!g28) & (!g33)));
	assign g1068 = (((!g14) & (!sk[74]) & (!g62) & (g101)) + ((!g14) & (!sk[74]) & (g62) & (!g101)) + ((!g14) & (!sk[74]) & (g62) & (g101)) + ((g14) & (!sk[74]) & (!g62) & (g101)) + ((g14) & (!sk[74]) & (g62) & (!g101)) + ((g14) & (!sk[74]) & (g62) & (g101)) + ((g14) & (sk[74]) & (g62) & (g101)));
	assign g1069 = (((!i_8_) & (!i_7_) & (g14) & (!sk[75]) & (!g62)) + ((!i_8_) & (!i_7_) & (g14) & (!sk[75]) & (g62)) + ((!i_8_) & (!i_7_) & (g14) & (sk[75]) & (g62)) + ((!i_8_) & (i_7_) & (g14) & (!sk[75]) & (!g62)) + ((!i_8_) & (i_7_) & (g14) & (!sk[75]) & (g62)) + ((i_8_) & (!i_7_) & (g14) & (!sk[75]) & (!g62)) + ((i_8_) & (!i_7_) & (g14) & (!sk[75]) & (g62)) + ((i_8_) & (i_7_) & (g14) & (!sk[75]) & (!g62)) + ((i_8_) & (i_7_) & (g14) & (!sk[75]) & (g62)));
	assign g1070 = (((!g6) & (!g14) & (!sk[76]) & (g43) & (!g1069)) + ((!g6) & (!g14) & (!sk[76]) & (g43) & (g1069)) + ((!g6) & (!g14) & (sk[76]) & (!g43) & (!g1069)) + ((!g6) & (!g14) & (sk[76]) & (g43) & (!g1069)) + ((!g6) & (g14) & (!sk[76]) & (g43) & (!g1069)) + ((!g6) & (g14) & (!sk[76]) & (g43) & (g1069)) + ((!g6) & (g14) & (sk[76]) & (!g43) & (!g1069)) + ((!g6) & (g14) & (sk[76]) & (g43) & (!g1069)) + ((g6) & (!g14) & (!sk[76]) & (g43) & (!g1069)) + ((g6) & (!g14) & (!sk[76]) & (g43) & (g1069)) + ((g6) & (!g14) & (sk[76]) & (!g43) & (!g1069)) + ((g6) & (!g14) & (sk[76]) & (g43) & (!g1069)) + ((g6) & (g14) & (!sk[76]) & (g43) & (!g1069)) + ((g6) & (g14) & (!sk[76]) & (g43) & (g1069)) + ((g6) & (g14) & (sk[76]) & (!g43) & (!g1069)));
	assign g1071 = (((!g2) & (!sk[77]) & (!g16) & (g43) & (!g1070)) + ((!g2) & (!sk[77]) & (!g16) & (g43) & (g1070)) + ((!g2) & (!sk[77]) & (g16) & (g43) & (!g1070)) + ((!g2) & (!sk[77]) & (g16) & (g43) & (g1070)) + ((!g2) & (sk[77]) & (!g16) & (!g43) & (g1070)) + ((!g2) & (sk[77]) & (!g16) & (g43) & (g1070)) + ((!g2) & (sk[77]) & (g16) & (!g43) & (g1070)) + ((g2) & (!sk[77]) & (!g16) & (g43) & (!g1070)) + ((g2) & (!sk[77]) & (!g16) & (g43) & (g1070)) + ((g2) & (!sk[77]) & (g16) & (g43) & (!g1070)) + ((g2) & (!sk[77]) & (g16) & (g43) & (g1070)) + ((g2) & (sk[77]) & (!g16) & (!g43) & (g1070)) + ((g2) & (sk[77]) & (!g16) & (g43) & (g1070)));
	assign g1072 = (((!sk[78]) & (g1068) & (!g1071)) + ((!sk[78]) & (g1068) & (g1071)) + ((sk[78]) & (!g1068) & (g1071)));
	assign g1073 = (((!g26) & (!g28) & (!g1068) & (sk[79]) & (g1070)) + ((!g26) & (!g28) & (g1068) & (!sk[79]) & (!g1070)) + ((!g26) & (!g28) & (g1068) & (!sk[79]) & (g1070)) + ((!g26) & (g28) & (!g1068) & (sk[79]) & (g1070)) + ((!g26) & (g28) & (g1068) & (!sk[79]) & (!g1070)) + ((!g26) & (g28) & (g1068) & (!sk[79]) & (g1070)) + ((g26) & (!g28) & (!g1068) & (sk[79]) & (!g1070)) + ((g26) & (!g28) & (!g1068) & (sk[79]) & (g1070)) + ((g26) & (!g28) & (g1068) & (!sk[79]) & (!g1070)) + ((g26) & (!g28) & (g1068) & (!sk[79]) & (g1070)) + ((g26) & (!g28) & (g1068) & (sk[79]) & (!g1070)) + ((g26) & (!g28) & (g1068) & (sk[79]) & (g1070)) + ((g26) & (g28) & (!g1068) & (sk[79]) & (g1070)) + ((g26) & (g28) & (g1068) & (!sk[79]) & (!g1070)) + ((g26) & (g28) & (g1068) & (!sk[79]) & (g1070)));
	assign g1074 = (((g59) & (!sk[80]) & (!g65)) + ((g59) & (!sk[80]) & (g65)) + ((g59) & (sk[80]) & (g65)));
	assign g1075 = (((!sk[81]) & (!i_0_) & (!i_1_) & (g6) & (!g15)) + ((!sk[81]) & (!i_0_) & (!i_1_) & (g6) & (g15)) + ((!sk[81]) & (!i_0_) & (i_1_) & (g6) & (!g15)) + ((!sk[81]) & (!i_0_) & (i_1_) & (g6) & (g15)) + ((!sk[81]) & (i_0_) & (!i_1_) & (g6) & (!g15)) + ((!sk[81]) & (i_0_) & (!i_1_) & (g6) & (g15)) + ((!sk[81]) & (i_0_) & (i_1_) & (g6) & (!g15)) + ((!sk[81]) & (i_0_) & (i_1_) & (g6) & (g15)) + ((sk[81]) & (i_0_) & (!i_1_) & (!g6) & (g15)) + ((sk[81]) & (i_0_) & (!i_1_) & (g6) & (!g15)) + ((sk[81]) & (i_0_) & (!i_1_) & (g6) & (g15)));
	assign g1076 = (((!g16) & (!g28) & (!g29) & (!g43) & (!g46) & (!g1064)) + ((!g16) & (!g28) & (!g29) & (g43) & (!g46) & (!g1064)) + ((!g16) & (!g28) & (g29) & (!g43) & (!g46) & (!g1064)) + ((!g16) & (!g28) & (g29) & (g43) & (!g46) & (!g1064)) + ((!g16) & (g28) & (!g29) & (!g43) & (!g46) & (!g1064)) + ((!g16) & (g28) & (!g29) & (g43) & (!g46) & (!g1064)) + ((!g16) & (g28) & (g29) & (!g43) & (!g46) & (!g1064)) + ((!g16) & (g28) & (g29) & (g43) & (!g46) & (!g1064)) + ((g16) & (!g28) & (g29) & (!g43) & (!g46) & (!g1064)) + ((g16) & (!g28) & (g29) & (g43) & (!g46) & (!g1064)) + ((g16) & (g28) & (g29) & (!g43) & (!g46) & (!g1064)));
	assign g1077 = (((!g33) & (!g1072) & (g1073) & (g1074) & (!g1075) & (g1076)) + ((!g33) & (g1072) & (g1073) & (g1074) & (!g1075) & (g1076)) + ((g33) & (g1072) & (g1073) & (g1074) & (!g1075) & (g1076)));
	assign o_24_ = (((!i_4_) & (!i_3_) & (g14) & (!sk[84]) & (!g42)) + ((!i_4_) & (!i_3_) & (g14) & (!sk[84]) & (g42)) + ((!i_4_) & (i_3_) & (g14) & (!sk[84]) & (!g42)) + ((!i_4_) & (i_3_) & (g14) & (!sk[84]) & (g42)) + ((i_4_) & (!i_3_) & (g14) & (!sk[84]) & (!g42)) + ((i_4_) & (!i_3_) & (g14) & (!sk[84]) & (g42)) + ((i_4_) & (i_3_) & (g14) & (!sk[84]) & (!g42)) + ((i_4_) & (i_3_) & (g14) & (!sk[84]) & (g42)) + ((i_4_) & (i_3_) & (g14) & (sk[84]) & (g42)));
	assign o_25_ = (((!sk[85]) & (!i_4_) & (!i_3_) & (g10) & (!g14)) + ((!sk[85]) & (!i_4_) & (!i_3_) & (g10) & (g14)) + ((!sk[85]) & (!i_4_) & (i_3_) & (g10) & (!g14)) + ((!sk[85]) & (!i_4_) & (i_3_) & (g10) & (g14)) + ((!sk[85]) & (i_4_) & (!i_3_) & (g10) & (!g14)) + ((!sk[85]) & (i_4_) & (!i_3_) & (g10) & (g14)) + ((!sk[85]) & (i_4_) & (i_3_) & (g10) & (!g14)) + ((!sk[85]) & (i_4_) & (i_3_) & (g10) & (g14)) + ((sk[85]) & (i_4_) & (i_3_) & (g10) & (g14)));
	assign g1080 = (((!sk[86]) & (!g2) & (!g43) & (g55)) + ((!sk[86]) & (!g2) & (g43) & (!g55)) + ((!sk[86]) & (!g2) & (g43) & (g55)) + ((!sk[86]) & (g2) & (!g43) & (g55)) + ((!sk[86]) & (g2) & (g43) & (!g55)) + ((!sk[86]) & (g2) & (g43) & (g55)) + ((sk[86]) & (!g2) & (g43) & (g55)) + ((sk[86]) & (g2) & (!g43) & (g55)) + ((sk[86]) & (g2) & (g43) & (g55)));
	assign g1081 = (((!g1062) & (!sk[87]) & (!g1072) & (g1080)) + ((!g1062) & (!sk[87]) & (g1072) & (!g1080)) + ((!g1062) & (!sk[87]) & (g1072) & (g1080)) + ((!g1062) & (sk[87]) & (g1072) & (!g1080)) + ((g1062) & (!sk[87]) & (!g1072) & (g1080)) + ((g1062) & (!sk[87]) & (g1072) & (!g1080)) + ((g1062) & (!sk[87]) & (g1072) & (g1080)));
	assign g1082 = (((!i_6_) & (!sk[88]) & (!i_7_) & (g14) & (!g40) & (g1060)) + ((!i_6_) & (!sk[88]) & (!i_7_) & (g14) & (g40) & (!g1060)) + ((!i_6_) & (!sk[88]) & (!i_7_) & (g14) & (g40) & (g1060)) + ((!i_6_) & (!sk[88]) & (i_7_) & (!g14) & (!g40) & (!g1060)) + ((!i_6_) & (!sk[88]) & (i_7_) & (!g14) & (!g40) & (g1060)) + ((!i_6_) & (!sk[88]) & (i_7_) & (!g14) & (g40) & (!g1060)) + ((!i_6_) & (!sk[88]) & (i_7_) & (!g14) & (g40) & (g1060)) + ((!i_6_) & (!sk[88]) & (i_7_) & (g14) & (!g40) & (!g1060)) + ((!i_6_) & (!sk[88]) & (i_7_) & (g14) & (!g40) & (g1060)) + ((!i_6_) & (!sk[88]) & (i_7_) & (g14) & (g40) & (!g1060)) + ((!i_6_) & (!sk[88]) & (i_7_) & (g14) & (g40) & (g1060)) + ((!i_6_) & (sk[88]) & (!i_7_) & (!g14) & (g40) & (!g1060)) + ((!i_6_) & (sk[88]) & (!i_7_) & (!g14) & (g40) & (g1060)) + ((!i_6_) & (sk[88]) & (!i_7_) & (g14) & (g40) & (!g1060)) + ((!i_6_) & (sk[88]) & (!i_7_) & (g14) & (g40) & (g1060)) + ((!i_6_) & (sk[88]) & (i_7_) & (g14) & (!g40) & (g1060)) + ((!i_6_) & (sk[88]) & (i_7_) & (g14) & (g40) & (g1060)) + ((i_6_) & (!sk[88]) & (!i_7_) & (g14) & (!g40) & (g1060)) + ((i_6_) & (!sk[88]) & (!i_7_) & (g14) & (g40) & (!g1060)) + ((i_6_) & (!sk[88]) & (!i_7_) & (g14) & (g40) & (g1060)) + ((i_6_) & (!sk[88]) & (i_7_) & (!g14) & (!g40) & (!g1060)) + ((i_6_) & (!sk[88]) & (i_7_) & (!g14) & (!g40) & (g1060)) + ((i_6_) & (!sk[88]) & (i_7_) & (!g14) & (g40) & (!g1060)) + ((i_6_) & (!sk[88]) & (i_7_) & (!g14) & (g40) & (g1060)) + ((i_6_) & (!sk[88]) & (i_7_) & (g14) & (!g40) & (!g1060)) + ((i_6_) & (!sk[88]) & (i_7_) & (g14) & (!g40) & (g1060)) + ((i_6_) & (!sk[88]) & (i_7_) & (g14) & (g40) & (!g1060)) + ((i_6_) & (!sk[88]) & (i_7_) & (g14) & (g40) & (g1060)) + ((i_6_) & (sk[88]) & (!i_7_) & (!g14) & (g40) & (!g1060)) + ((i_6_) & (sk[88]) & (!i_7_) & (!g14) & (g40) & (g1060)) + ((i_6_) & (sk[88]) & (!i_7_) & (g14) & (!g40) & (g1060)) + ((i_6_) & (sk[88]) & (!i_7_) & (g14) & (g40) & (!g1060)) + ((i_6_) & (sk[88]) & (!i_7_) & (g14) & (g40) & (g1060)) + ((i_6_) & (sk[88]) & (i_7_) & (g14) & (!g40) & (g1060)) + ((i_6_) & (sk[88]) & (i_7_) & (g14) & (g40) & (g1060)));
	assign o_26_ = (((!g21) & (!g23) & (!g25) & (sk[89]) & (!g1081) & (!g1082)) + ((!g21) & (!g23) & (!g25) & (sk[89]) & (!g1081) & (g1082)) + ((!g21) & (!g23) & (!g25) & (sk[89]) & (g1081) & (g1082)) + ((!g21) & (!g23) & (g25) & (!sk[89]) & (!g1081) & (g1082)) + ((!g21) & (!g23) & (g25) & (!sk[89]) & (g1081) & (!g1082)) + ((!g21) & (!g23) & (g25) & (!sk[89]) & (g1081) & (g1082)) + ((!g21) & (!g23) & (g25) & (sk[89]) & (!g1081) & (!g1082)) + ((!g21) & (!g23) & (g25) & (sk[89]) & (!g1081) & (g1082)) + ((!g21) & (!g23) & (g25) & (sk[89]) & (g1081) & (g1082)) + ((!g21) & (g23) & (!g25) & (!sk[89]) & (!g1081) & (!g1082)) + ((!g21) & (g23) & (!g25) & (!sk[89]) & (!g1081) & (g1082)) + ((!g21) & (g23) & (!g25) & (!sk[89]) & (g1081) & (!g1082)) + ((!g21) & (g23) & (!g25) & (!sk[89]) & (g1081) & (g1082)) + ((!g21) & (g23) & (!g25) & (sk[89]) & (!g1081) & (!g1082)) + ((!g21) & (g23) & (!g25) & (sk[89]) & (!g1081) & (g1082)) + ((!g21) & (g23) & (!g25) & (sk[89]) & (g1081) & (g1082)) + ((!g21) & (g23) & (g25) & (!sk[89]) & (!g1081) & (!g1082)) + ((!g21) & (g23) & (g25) & (!sk[89]) & (!g1081) & (g1082)) + ((!g21) & (g23) & (g25) & (!sk[89]) & (g1081) & (!g1082)) + ((!g21) & (g23) & (g25) & (!sk[89]) & (g1081) & (g1082)) + ((!g21) & (g23) & (g25) & (sk[89]) & (!g1081) & (g1082)) + ((!g21) & (g23) & (g25) & (sk[89]) & (g1081) & (g1082)) + ((g21) & (!g23) & (!g25) & (sk[89]) & (!g1081) & (!g1082)) + ((g21) & (!g23) & (!g25) & (sk[89]) & (!g1081) & (g1082)) + ((g21) & (!g23) & (!g25) & (sk[89]) & (g1081) & (g1082)) + ((g21) & (!g23) & (g25) & (!sk[89]) & (!g1081) & (g1082)) + ((g21) & (!g23) & (g25) & (!sk[89]) & (g1081) & (!g1082)) + ((g21) & (!g23) & (g25) & (!sk[89]) & (g1081) & (g1082)) + ((g21) & (!g23) & (g25) & (sk[89]) & (!g1081) & (!g1082)) + ((g21) & (!g23) & (g25) & (sk[89]) & (!g1081) & (g1082)) + ((g21) & (!g23) & (g25) & (sk[89]) & (g1081) & (g1082)) + ((g21) & (g23) & (!g25) & (!sk[89]) & (!g1081) & (!g1082)) + ((g21) & (g23) & (!g25) & (!sk[89]) & (!g1081) & (g1082)) + ((g21) & (g23) & (!g25) & (!sk[89]) & (g1081) & (!g1082)) + ((g21) & (g23) & (!g25) & (!sk[89]) & (g1081) & (g1082)) + ((g21) & (g23) & (!g25) & (sk[89]) & (!g1081) & (!g1082)) + ((g21) & (g23) & (!g25) & (sk[89]) & (!g1081) & (g1082)) + ((g21) & (g23) & (!g25) & (sk[89]) & (g1081) & (g1082)) + ((g21) & (g23) & (g25) & (!sk[89]) & (!g1081) & (!g1082)) + ((g21) & (g23) & (g25) & (!sk[89]) & (!g1081) & (g1082)) + ((g21) & (g23) & (g25) & (!sk[89]) & (g1081) & (!g1082)) + ((g21) & (g23) & (g25) & (!sk[89]) & (g1081) & (g1082)) + ((g21) & (g23) & (g25) & (sk[89]) & (!g1081) & (!g1082)) + ((g21) & (g23) & (g25) & (sk[89]) & (!g1081) & (g1082)) + ((g21) & (g23) & (g25) & (sk[89]) & (g1081) & (g1082)));
	assign g1084 = (((!g1) & (!i_4_) & (!sk[90]) & (i_3_) & (!i_5_) & (g14)) + ((!g1) & (!i_4_) & (!sk[90]) & (i_3_) & (i_5_) & (!g14)) + ((!g1) & (!i_4_) & (!sk[90]) & (i_3_) & (i_5_) & (g14)) + ((!g1) & (i_4_) & (!sk[90]) & (!i_3_) & (!i_5_) & (!g14)) + ((!g1) & (i_4_) & (!sk[90]) & (!i_3_) & (!i_5_) & (g14)) + ((!g1) & (i_4_) & (!sk[90]) & (!i_3_) & (i_5_) & (!g14)) + ((!g1) & (i_4_) & (!sk[90]) & (!i_3_) & (i_5_) & (g14)) + ((!g1) & (i_4_) & (!sk[90]) & (i_3_) & (!i_5_) & (!g14)) + ((!g1) & (i_4_) & (!sk[90]) & (i_3_) & (!i_5_) & (g14)) + ((!g1) & (i_4_) & (!sk[90]) & (i_3_) & (i_5_) & (!g14)) + ((!g1) & (i_4_) & (!sk[90]) & (i_3_) & (i_5_) & (g14)) + ((!g1) & (i_4_) & (sk[90]) & (i_3_) & (i_5_) & (g14)) + ((g1) & (!i_4_) & (!sk[90]) & (i_3_) & (!i_5_) & (g14)) + ((g1) & (!i_4_) & (!sk[90]) & (i_3_) & (i_5_) & (!g14)) + ((g1) & (!i_4_) & (!sk[90]) & (i_3_) & (i_5_) & (g14)) + ((g1) & (i_4_) & (!sk[90]) & (!i_3_) & (!i_5_) & (!g14)) + ((g1) & (i_4_) & (!sk[90]) & (!i_3_) & (!i_5_) & (g14)) + ((g1) & (i_4_) & (!sk[90]) & (!i_3_) & (i_5_) & (!g14)) + ((g1) & (i_4_) & (!sk[90]) & (!i_3_) & (i_5_) & (g14)) + ((g1) & (i_4_) & (!sk[90]) & (i_3_) & (!i_5_) & (!g14)) + ((g1) & (i_4_) & (!sk[90]) & (i_3_) & (!i_5_) & (g14)) + ((g1) & (i_4_) & (!sk[90]) & (i_3_) & (i_5_) & (!g14)) + ((g1) & (i_4_) & (!sk[90]) & (i_3_) & (i_5_) & (g14)));
	assign g1085 = (((!sk[91]) & (!g10) & (!g18) & (g40) & (!g457) & (g1081)) + ((!sk[91]) & (!g10) & (!g18) & (g40) & (g457) & (!g1081)) + ((!sk[91]) & (!g10) & (!g18) & (g40) & (g457) & (g1081)) + ((!sk[91]) & (!g10) & (g18) & (!g40) & (!g457) & (!g1081)) + ((!sk[91]) & (!g10) & (g18) & (!g40) & (!g457) & (g1081)) + ((!sk[91]) & (!g10) & (g18) & (!g40) & (g457) & (!g1081)) + ((!sk[91]) & (!g10) & (g18) & (!g40) & (g457) & (g1081)) + ((!sk[91]) & (!g10) & (g18) & (g40) & (!g457) & (!g1081)) + ((!sk[91]) & (!g10) & (g18) & (g40) & (!g457) & (g1081)) + ((!sk[91]) & (!g10) & (g18) & (g40) & (g457) & (!g1081)) + ((!sk[91]) & (!g10) & (g18) & (g40) & (g457) & (g1081)) + ((!sk[91]) & (g10) & (!g18) & (g40) & (!g457) & (g1081)) + ((!sk[91]) & (g10) & (!g18) & (g40) & (g457) & (!g1081)) + ((!sk[91]) & (g10) & (!g18) & (g40) & (g457) & (g1081)) + ((!sk[91]) & (g10) & (g18) & (!g40) & (!g457) & (!g1081)) + ((!sk[91]) & (g10) & (g18) & (!g40) & (!g457) & (g1081)) + ((!sk[91]) & (g10) & (g18) & (!g40) & (g457) & (!g1081)) + ((!sk[91]) & (g10) & (g18) & (!g40) & (g457) & (g1081)) + ((!sk[91]) & (g10) & (g18) & (g40) & (!g457) & (!g1081)) + ((!sk[91]) & (g10) & (g18) & (g40) & (!g457) & (g1081)) + ((!sk[91]) & (g10) & (g18) & (g40) & (g457) & (!g1081)) + ((!sk[91]) & (g10) & (g18) & (g40) & (g457) & (g1081)) + ((sk[91]) & (!g10) & (g18) & (!g40) & (!g457) & (!g1081)) + ((sk[91]) & (!g10) & (g18) & (!g40) & (g457) & (!g1081)) + ((sk[91]) & (!g10) & (g18) & (g40) & (!g457) & (!g1081)) + ((sk[91]) & (!g10) & (g18) & (g40) & (g457) & (!g1081)) + ((sk[91]) & (g10) & (!g18) & (g40) & (!g457) & (!g1081)) + ((sk[91]) & (g10) & (!g18) & (g40) & (!g457) & (g1081)) + ((sk[91]) & (g10) & (!g18) & (g40) & (g457) & (!g1081)) + ((sk[91]) & (g10) & (!g18) & (g40) & (g457) & (g1081)) + ((sk[91]) & (g10) & (g18) & (!g40) & (!g457) & (!g1081)) + ((sk[91]) & (g10) & (g18) & (!g40) & (g457) & (!g1081)) + ((sk[91]) & (g10) & (g18) & (!g40) & (g457) & (g1081)) + ((sk[91]) & (g10) & (g18) & (g40) & (!g457) & (!g1081)) + ((sk[91]) & (g10) & (g18) & (g40) & (!g457) & (g1081)) + ((sk[91]) & (g10) & (g18) & (g40) & (g457) & (!g1081)) + ((sk[91]) & (g10) & (g18) & (g40) & (g457) & (g1081)));
	assign g1086 = (((!g33) & (!g1062) & (g1072) & (!sk[92]) & (!g1080)) + ((!g33) & (!g1062) & (g1072) & (!sk[92]) & (g1080)) + ((!g33) & (g1062) & (g1072) & (!sk[92]) & (!g1080)) + ((!g33) & (g1062) & (g1072) & (!sk[92]) & (g1080)) + ((g33) & (!g1062) & (!g1072) & (sk[92]) & (!g1080)) + ((g33) & (!g1062) & (!g1072) & (sk[92]) & (g1080)) + ((g33) & (!g1062) & (g1072) & (!sk[92]) & (!g1080)) + ((g33) & (!g1062) & (g1072) & (!sk[92]) & (g1080)) + ((g33) & (!g1062) & (g1072) & (sk[92]) & (g1080)) + ((g33) & (g1062) & (!g1072) & (sk[92]) & (!g1080)) + ((g33) & (g1062) & (!g1072) & (sk[92]) & (g1080)) + ((g33) & (g1062) & (g1072) & (!sk[92]) & (!g1080)) + ((g33) & (g1062) & (g1072) & (!sk[92]) & (g1080)) + ((g33) & (g1062) & (g1072) & (sk[92]) & (!g1080)) + ((g33) & (g1062) & (g1072) & (sk[92]) & (g1080)));
	assign g1087 = (((!i_4_) & (!g40) & (!sk[93]) & (g1075)) + ((!i_4_) & (!g40) & (sk[93]) & (!g1075)) + ((!i_4_) & (g40) & (!sk[93]) & (!g1075)) + ((!i_4_) & (g40) & (!sk[93]) & (g1075)) + ((!i_4_) & (g40) & (sk[93]) & (!g1075)) + ((i_4_) & (!g40) & (!sk[93]) & (g1075)) + ((i_4_) & (!g40) & (sk[93]) & (!g1075)) + ((i_4_) & (g40) & (!sk[93]) & (!g1075)) + ((i_4_) & (g40) & (!sk[93]) & (g1075)));
	assign g1088 = (((!g28) & (!g45) & (!g1062) & (!g1072) & (!g1080) & (!g1087)) + ((!g28) & (!g45) & (!g1062) & (!g1072) & (!g1080) & (g1087)) + ((!g28) & (!g45) & (!g1062) & (!g1072) & (g1080) & (!g1087)) + ((!g28) & (!g45) & (!g1062) & (!g1072) & (g1080) & (g1087)) + ((!g28) & (!g45) & (!g1062) & (g1072) & (!g1080) & (!g1087)) + ((!g28) & (!g45) & (!g1062) & (g1072) & (!g1080) & (g1087)) + ((!g28) & (!g45) & (!g1062) & (g1072) & (g1080) & (!g1087)) + ((!g28) & (!g45) & (!g1062) & (g1072) & (g1080) & (g1087)) + ((!g28) & (!g45) & (g1062) & (!g1072) & (!g1080) & (!g1087)) + ((!g28) & (!g45) & (g1062) & (!g1072) & (!g1080) & (g1087)) + ((!g28) & (!g45) & (g1062) & (!g1072) & (g1080) & (!g1087)) + ((!g28) & (!g45) & (g1062) & (!g1072) & (g1080) & (g1087)) + ((!g28) & (!g45) & (g1062) & (g1072) & (!g1080) & (!g1087)) + ((!g28) & (!g45) & (g1062) & (g1072) & (!g1080) & (g1087)) + ((!g28) & (!g45) & (g1062) & (g1072) & (g1080) & (!g1087)) + ((!g28) & (!g45) & (g1062) & (g1072) & (g1080) & (g1087)) + ((!g28) & (g45) & (!g1062) & (!g1072) & (!g1080) & (g1087)) + ((!g28) & (g45) & (!g1062) & (!g1072) & (g1080) & (g1087)) + ((!g28) & (g45) & (!g1062) & (g1072) & (!g1080) & (g1087)) + ((!g28) & (g45) & (!g1062) & (g1072) & (g1080) & (g1087)) + ((!g28) & (g45) & (g1062) & (!g1072) & (!g1080) & (g1087)) + ((!g28) & (g45) & (g1062) & (!g1072) & (g1080) & (g1087)) + ((!g28) & (g45) & (g1062) & (g1072) & (!g1080) & (g1087)) + ((!g28) & (g45) & (g1062) & (g1072) & (g1080) & (g1087)) + ((g28) & (!g45) & (!g1062) & (g1072) & (!g1080) & (!g1087)) + ((g28) & (!g45) & (!g1062) & (g1072) & (!g1080) & (g1087)) + ((g28) & (g45) & (!g1062) & (g1072) & (!g1080) & (g1087)));
	assign o_27_ = (((!g1084) & (!sk[95]) & (!g1085) & (g1086) & (!g1088)) + ((!g1084) & (!sk[95]) & (!g1085) & (g1086) & (g1088)) + ((!g1084) & (!sk[95]) & (g1085) & (g1086) & (!g1088)) + ((!g1084) & (!sk[95]) & (g1085) & (g1086) & (g1088)) + ((!g1084) & (sk[95]) & (!g1085) & (!g1086) & (!g1088)) + ((!g1084) & (sk[95]) & (!g1085) & (g1086) & (!g1088)) + ((!g1084) & (sk[95]) & (!g1085) & (g1086) & (g1088)) + ((!g1084) & (sk[95]) & (g1085) & (!g1086) & (!g1088)) + ((!g1084) & (sk[95]) & (g1085) & (!g1086) & (g1088)) + ((!g1084) & (sk[95]) & (g1085) & (g1086) & (!g1088)) + ((!g1084) & (sk[95]) & (g1085) & (g1086) & (g1088)) + ((g1084) & (!sk[95]) & (!g1085) & (g1086) & (!g1088)) + ((g1084) & (!sk[95]) & (!g1085) & (g1086) & (g1088)) + ((g1084) & (!sk[95]) & (g1085) & (g1086) & (!g1088)) + ((g1084) & (!sk[95]) & (g1085) & (g1086) & (g1088)) + ((g1084) & (sk[95]) & (!g1085) & (!g1086) & (!g1088)) + ((g1084) & (sk[95]) & (!g1085) & (!g1086) & (g1088)) + ((g1084) & (sk[95]) & (!g1085) & (g1086) & (!g1088)) + ((g1084) & (sk[95]) & (!g1085) & (g1086) & (g1088)) + ((g1084) & (sk[95]) & (g1085) & (!g1086) & (!g1088)) + ((g1084) & (sk[95]) & (g1085) & (!g1086) & (g1088)) + ((g1084) & (sk[95]) & (g1085) & (g1086) & (!g1088)) + ((g1084) & (sk[95]) & (g1085) & (g1086) & (g1088)));
	assign g1090 = (((g1071) & (!sk[96]) & (!g1080)) + ((g1071) & (!sk[96]) & (g1080)) + ((g1071) & (sk[96]) & (!g1080)));
	assign g1091 = (((g1) & (!sk[97]) & (!g40)) + ((g1) & (!sk[97]) & (g40)) + ((g1) & (sk[97]) & (g40)));
	assign o_28_ = (((!g23) & (!g37) & (!g1081) & (!g1085) & (!g1090) & (!g1091)) + ((!g23) & (!g37) & (!g1081) & (!g1085) & (!g1090) & (g1091)) + ((!g23) & (!g37) & (!g1081) & (!g1085) & (g1090) & (!g1091)) + ((!g23) & (!g37) & (!g1081) & (!g1085) & (g1090) & (g1091)) + ((!g23) & (!g37) & (!g1081) & (g1085) & (!g1090) & (!g1091)) + ((!g23) & (!g37) & (!g1081) & (g1085) & (!g1090) & (g1091)) + ((!g23) & (!g37) & (!g1081) & (g1085) & (g1090) & (!g1091)) + ((!g23) & (!g37) & (!g1081) & (g1085) & (g1090) & (g1091)) + ((!g23) & (!g37) & (g1081) & (!g1085) & (!g1090) & (!g1091)) + ((!g23) & (!g37) & (g1081) & (!g1085) & (!g1090) & (g1091)) + ((!g23) & (!g37) & (g1081) & (!g1085) & (g1090) & (g1091)) + ((!g23) & (!g37) & (g1081) & (g1085) & (!g1090) & (!g1091)) + ((!g23) & (!g37) & (g1081) & (g1085) & (!g1090) & (g1091)) + ((!g23) & (!g37) & (g1081) & (g1085) & (g1090) & (!g1091)) + ((!g23) & (!g37) & (g1081) & (g1085) & (g1090) & (g1091)) + ((!g23) & (g37) & (!g1081) & (!g1085) & (!g1090) & (!g1091)) + ((!g23) & (g37) & (!g1081) & (!g1085) & (!g1090) & (g1091)) + ((!g23) & (g37) & (!g1081) & (!g1085) & (g1090) & (!g1091)) + ((!g23) & (g37) & (!g1081) & (!g1085) & (g1090) & (g1091)) + ((!g23) & (g37) & (!g1081) & (g1085) & (!g1090) & (!g1091)) + ((!g23) & (g37) & (!g1081) & (g1085) & (!g1090) & (g1091)) + ((!g23) & (g37) & (!g1081) & (g1085) & (g1090) & (!g1091)) + ((!g23) & (g37) & (!g1081) & (g1085) & (g1090) & (g1091)) + ((!g23) & (g37) & (g1081) & (!g1085) & (!g1090) & (g1091)) + ((!g23) & (g37) & (g1081) & (!g1085) & (g1090) & (g1091)) + ((!g23) & (g37) & (g1081) & (g1085) & (!g1090) & (!g1091)) + ((!g23) & (g37) & (g1081) & (g1085) & (!g1090) & (g1091)) + ((!g23) & (g37) & (g1081) & (g1085) & (g1090) & (!g1091)) + ((!g23) & (g37) & (g1081) & (g1085) & (g1090) & (g1091)) + ((g23) & (!g37) & (!g1081) & (!g1085) & (!g1090) & (!g1091)) + ((g23) & (!g37) & (!g1081) & (!g1085) & (!g1090) & (g1091)) + ((g23) & (!g37) & (!g1081) & (!g1085) & (g1090) & (g1091)) + ((g23) & (!g37) & (!g1081) & (g1085) & (!g1090) & (!g1091)) + ((g23) & (!g37) & (!g1081) & (g1085) & (!g1090) & (g1091)) + ((g23) & (!g37) & (!g1081) & (g1085) & (g1090) & (!g1091)) + ((g23) & (!g37) & (!g1081) & (g1085) & (g1090) & (g1091)) + ((g23) & (!g37) & (g1081) & (!g1085) & (!g1090) & (!g1091)) + ((g23) & (!g37) & (g1081) & (!g1085) & (!g1090) & (g1091)) + ((g23) & (!g37) & (g1081) & (!g1085) & (g1090) & (g1091)) + ((g23) & (!g37) & (g1081) & (g1085) & (!g1090) & (!g1091)) + ((g23) & (!g37) & (g1081) & (g1085) & (!g1090) & (g1091)) + ((g23) & (!g37) & (g1081) & (g1085) & (g1090) & (!g1091)) + ((g23) & (!g37) & (g1081) & (g1085) & (g1090) & (g1091)) + ((g23) & (g37) & (!g1081) & (!g1085) & (!g1090) & (g1091)) + ((g23) & (g37) & (!g1081) & (!g1085) & (g1090) & (g1091)) + ((g23) & (g37) & (!g1081) & (g1085) & (!g1090) & (!g1091)) + ((g23) & (g37) & (!g1081) & (g1085) & (!g1090) & (g1091)) + ((g23) & (g37) & (!g1081) & (g1085) & (g1090) & (!g1091)) + ((g23) & (g37) & (!g1081) & (g1085) & (g1090) & (g1091)) + ((g23) & (g37) & (g1081) & (!g1085) & (!g1090) & (g1091)) + ((g23) & (g37) & (g1081) & (!g1085) & (g1090) & (g1091)) + ((g23) & (g37) & (g1081) & (g1085) & (!g1090) & (!g1091)) + ((g23) & (g37) & (g1081) & (g1085) & (!g1090) & (g1091)) + ((g23) & (g37) & (g1081) & (g1085) & (g1090) & (!g1091)) + ((g23) & (g37) & (g1081) & (g1085) & (g1090) & (g1091)));
	assign o_29_ = (((!g21) & (!g634) & (!g1081) & (sk[99]) & (!g1086) & (!g1090)) + ((!g21) & (!g634) & (!g1081) & (sk[99]) & (g1086) & (!g1090)) + ((!g21) & (!g634) & (!g1081) & (sk[99]) & (g1086) & (g1090)) + ((!g21) & (!g634) & (g1081) & (!sk[99]) & (!g1086) & (g1090)) + ((!g21) & (!g634) & (g1081) & (!sk[99]) & (g1086) & (!g1090)) + ((!g21) & (!g634) & (g1081) & (!sk[99]) & (g1086) & (g1090)) + ((!g21) & (!g634) & (g1081) & (sk[99]) & (!g1086) & (!g1090)) + ((!g21) & (!g634) & (g1081) & (sk[99]) & (g1086) & (!g1090)) + ((!g21) & (!g634) & (g1081) & (sk[99]) & (g1086) & (g1090)) + ((!g21) & (g634) & (!g1081) & (!sk[99]) & (!g1086) & (!g1090)) + ((!g21) & (g634) & (!g1081) & (!sk[99]) & (!g1086) & (g1090)) + ((!g21) & (g634) & (!g1081) & (!sk[99]) & (g1086) & (!g1090)) + ((!g21) & (g634) & (!g1081) & (!sk[99]) & (g1086) & (g1090)) + ((!g21) & (g634) & (!g1081) & (sk[99]) & (g1086) & (!g1090)) + ((!g21) & (g634) & (!g1081) & (sk[99]) & (g1086) & (g1090)) + ((!g21) & (g634) & (g1081) & (!sk[99]) & (!g1086) & (!g1090)) + ((!g21) & (g634) & (g1081) & (!sk[99]) & (!g1086) & (g1090)) + ((!g21) & (g634) & (g1081) & (!sk[99]) & (g1086) & (!g1090)) + ((!g21) & (g634) & (g1081) & (!sk[99]) & (g1086) & (g1090)) + ((!g21) & (g634) & (g1081) & (sk[99]) & (g1086) & (!g1090)) + ((!g21) & (g634) & (g1081) & (sk[99]) & (g1086) & (g1090)) + ((g21) & (!g634) & (!g1081) & (sk[99]) & (!g1086) & (!g1090)) + ((g21) & (!g634) & (!g1081) & (sk[99]) & (!g1086) & (g1090)) + ((g21) & (!g634) & (!g1081) & (sk[99]) & (g1086) & (!g1090)) + ((g21) & (!g634) & (!g1081) & (sk[99]) & (g1086) & (g1090)) + ((g21) & (!g634) & (g1081) & (!sk[99]) & (!g1086) & (g1090)) + ((g21) & (!g634) & (g1081) & (!sk[99]) & (g1086) & (!g1090)) + ((g21) & (!g634) & (g1081) & (!sk[99]) & (g1086) & (g1090)) + ((g21) & (!g634) & (g1081) & (sk[99]) & (!g1086) & (!g1090)) + ((g21) & (!g634) & (g1081) & (sk[99]) & (g1086) & (!g1090)) + ((g21) & (!g634) & (g1081) & (sk[99]) & (g1086) & (g1090)) + ((g21) & (g634) & (!g1081) & (!sk[99]) & (!g1086) & (!g1090)) + ((g21) & (g634) & (!g1081) & (!sk[99]) & (!g1086) & (g1090)) + ((g21) & (g634) & (!g1081) & (!sk[99]) & (g1086) & (!g1090)) + ((g21) & (g634) & (!g1081) & (!sk[99]) & (g1086) & (g1090)) + ((g21) & (g634) & (!g1081) & (sk[99]) & (!g1086) & (!g1090)) + ((g21) & (g634) & (!g1081) & (sk[99]) & (!g1086) & (g1090)) + ((g21) & (g634) & (!g1081) & (sk[99]) & (g1086) & (!g1090)) + ((g21) & (g634) & (!g1081) & (sk[99]) & (g1086) & (g1090)) + ((g21) & (g634) & (g1081) & (!sk[99]) & (!g1086) & (!g1090)) + ((g21) & (g634) & (g1081) & (!sk[99]) & (!g1086) & (g1090)) + ((g21) & (g634) & (g1081) & (!sk[99]) & (g1086) & (!g1090)) + ((g21) & (g634) & (g1081) & (!sk[99]) & (g1086) & (g1090)) + ((g21) & (g634) & (g1081) & (sk[99]) & (g1086) & (!g1090)) + ((g21) & (g634) & (g1081) & (sk[99]) & (g1086) & (g1090)));
	assign g1094 = (((!sk[100]) & (!g127) & (!g74) & (g114)) + ((!sk[100]) & (!g127) & (g74) & (!g114)) + ((!sk[100]) & (!g127) & (g74) & (g114)) + ((!sk[100]) & (g127) & (!g74) & (g114)) + ((!sk[100]) & (g127) & (g74) & (!g114)) + ((!sk[100]) & (g127) & (g74) & (g114)) + ((sk[100]) & (!g127) & (g74) & (!g114)) + ((sk[100]) & (g127) & (g74) & (!g114)) + ((sk[100]) & (g127) & (g74) & (g114)));
	assign g1095 = (((!i_12_) & (!i_13_) & (i_14_) & (!g107) & (g74) & (!g91)) + ((!i_12_) & (!i_13_) & (i_14_) & (!g107) & (g74) & (g91)) + ((!i_12_) & (!i_13_) & (i_14_) & (g107) & (g74) & (!g91)) + ((!i_12_) & (i_13_) & (i_14_) & (!g107) & (g74) & (!g91)) + ((!i_12_) & (i_13_) & (i_14_) & (!g107) & (g74) & (g91)) + ((!i_12_) & (i_13_) & (i_14_) & (g107) & (g74) & (!g91)) + ((i_12_) & (!i_13_) & (i_14_) & (!g107) & (g74) & (!g91)) + ((i_12_) & (!i_13_) & (i_14_) & (g107) & (g74) & (!g91)) + ((i_12_) & (i_13_) & (!i_14_) & (!g107) & (g74) & (!g91)) + ((i_12_) & (i_13_) & (!i_14_) & (g107) & (g74) & (!g91)) + ((i_12_) & (i_13_) & (i_14_) & (!g107) & (g74) & (!g91)) + ((i_12_) & (i_13_) & (i_14_) & (!g107) & (g74) & (g91)));
	assign g1096 = (((!i_12_) & (!i_13_) & (!i_14_) & (!g75) & (!g107) & (!g91)) + ((!i_12_) & (!i_13_) & (!i_14_) & (!g75) & (g107) & (!g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g75) & (!g107) & (!g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g75) & (!g107) & (g91)) + ((i_12_) & (!i_13_) & (!i_14_) & (!g75) & (!g107) & (!g91)) + ((i_12_) & (!i_13_) & (!i_14_) & (!g75) & (!g107) & (g91)) + ((i_12_) & (!i_13_) & (!i_14_) & (!g75) & (g107) & (!g91)) + ((i_12_) & (i_13_) & (!i_14_) & (!g75) & (!g107) & (!g91)) + ((i_12_) & (i_13_) & (!i_14_) & (!g75) & (!g107) & (g91)));
	assign g1097 = (((!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (!g75) & (g112)) + ((!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (!g75) & (g112)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g75) & (g112)) + ((!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g75) & (g112)) + ((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g75) & (g112)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g75) & (g112)) + ((i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (!g75) & (g112)) + ((i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (!g75) & (g112)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g75) & (g112)) + ((i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g75) & (g112)) + ((i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g75) & (g112)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g75) & (g112)));
	assign g1098 = (((!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g112) & (g74)) + ((!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112) & (g74)) + ((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112) & (g74)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g112) & (g74)) + ((i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g112) & (g74)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g112) & (g74)) + ((i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g112) & (g74)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112) & (g74)));
	assign g1099 = (((!g1094) & (!g793) & (!g1095) & (!g1096) & (!g1097) & (!g1098)));
	assign g1100 = (((!i_8_) & (!sk[106]) & (!g73) & (g358)) + ((!i_8_) & (!sk[106]) & (g73) & (!g358)) + ((!i_8_) & (!sk[106]) & (g73) & (g358)) + ((!i_8_) & (sk[106]) & (g73) & (g358)) + ((i_8_) & (!sk[106]) & (!g73) & (g358)) + ((i_8_) & (!sk[106]) & (g73) & (!g358)) + ((i_8_) & (!sk[106]) & (g73) & (g358)));
	assign g1101 = (((!g1100) & (!g670) & (!g463) & (!g464) & (!g465) & (!g466)));
	assign g1102 = (((!sk[108]) & (!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[108]) & (!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[108]) & (!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g112)) + ((!sk[108]) & (!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g112)) + ((!sk[108]) & (!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((!sk[108]) & (!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g112)) + ((!sk[108]) & (!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g112)) + ((!sk[108]) & (!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g112)) + ((!sk[108]) & (!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[108]) & (!i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[108]) & (!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g112)) + ((!sk[108]) & (i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[108]) & (i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[108]) & (i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g112)) + ((!sk[108]) & (i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g112)) + ((!sk[108]) & (i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((!sk[108]) & (i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g112)) + ((!sk[108]) & (i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g112)) + ((!sk[108]) & (i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g112)) + ((!sk[108]) & (i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[108]) & (i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[108]) & (i_15_) & (i_12_) & (i_13_) & (i_14_) & (g112)) + ((sk[108]) & (!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g112)) + ((sk[108]) & (i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g112)) + ((sk[108]) & (i_15_) & (i_12_) & (i_13_) & (i_14_) & (g112)));
	assign g1103 = (((!g22) & (!g174) & (!sk[109]) & (g761)) + ((!g22) & (g174) & (!sk[109]) & (!g761)) + ((!g22) & (g174) & (!sk[109]) & (g761)) + ((!g22) & (g174) & (sk[109]) & (g761)) + ((g22) & (!g174) & (!sk[109]) & (g761)) + ((g22) & (!g174) & (sk[109]) & (g761)) + ((g22) & (g174) & (!sk[109]) & (!g761)) + ((g22) & (g174) & (!sk[109]) & (g761)) + ((g22) & (g174) & (sk[109]) & (g761)));
	assign g1104 = (((!i_8_) & (!g73) & (!sk[110]) & (g605) & (!g635)) + ((!i_8_) & (!g73) & (!sk[110]) & (g605) & (g635)) + ((!i_8_) & (g73) & (!sk[110]) & (g605) & (!g635)) + ((!i_8_) & (g73) & (!sk[110]) & (g605) & (g635)) + ((i_8_) & (!g73) & (!sk[110]) & (g605) & (!g635)) + ((i_8_) & (!g73) & (!sk[110]) & (g605) & (g635)) + ((i_8_) & (g73) & (!sk[110]) & (g605) & (!g635)) + ((i_8_) & (g73) & (!sk[110]) & (g605) & (g635)) + ((i_8_) & (g73) & (sk[110]) & (!g605) & (g635)) + ((i_8_) & (g73) & (sk[110]) & (g605) & (!g635)) + ((i_8_) & (g73) & (sk[110]) & (g605) & (g635)));
	assign g1105 = (((!i_8_) & (!sk[111]) & (!g73) & (g337) & (!g851)) + ((!i_8_) & (!sk[111]) & (!g73) & (g337) & (g851)) + ((!i_8_) & (!sk[111]) & (g73) & (g337) & (!g851)) + ((!i_8_) & (!sk[111]) & (g73) & (g337) & (g851)) + ((i_8_) & (!sk[111]) & (!g73) & (g337) & (!g851)) + ((i_8_) & (!sk[111]) & (!g73) & (g337) & (g851)) + ((i_8_) & (!sk[111]) & (g73) & (g337) & (!g851)) + ((i_8_) & (!sk[111]) & (g73) & (g337) & (g851)) + ((i_8_) & (sk[111]) & (g73) & (!g337) & (!g851)) + ((i_8_) & (sk[111]) & (g73) & (g337) & (!g851)) + ((i_8_) & (sk[111]) & (g73) & (g337) & (g851)));
	assign g1106 = (((!g75) & (g949) & (!g1102) & (g1103) & (!g1104) & (!g1105)) + ((g75) & (!g949) & (!g1102) & (!g1103) & (!g1104) & (!g1105)) + ((g75) & (!g949) & (!g1102) & (g1103) & (!g1104) & (!g1105)) + ((g75) & (!g949) & (g1102) & (!g1103) & (!g1104) & (!g1105)) + ((g75) & (!g949) & (g1102) & (g1103) & (!g1104) & (!g1105)) + ((g75) & (g949) & (!g1102) & (!g1103) & (!g1104) & (!g1105)) + ((g75) & (g949) & (!g1102) & (g1103) & (!g1104) & (!g1105)) + ((g75) & (g949) & (g1102) & (!g1103) & (!g1104) & (!g1105)) + ((g75) & (g949) & (g1102) & (g1103) & (!g1104) & (!g1105)));
	assign g1107 = (((!sk[113]) & (!g4) & (!g27) & (g725)) + ((!sk[113]) & (!g4) & (g27) & (!g725)) + ((!sk[113]) & (!g4) & (g27) & (g725)) + ((!sk[113]) & (g4) & (!g27) & (g725)) + ((!sk[113]) & (g4) & (g27) & (!g725)) + ((!sk[113]) & (g4) & (g27) & (g725)) + ((sk[113]) & (!g4) & (!g27) & (g725)) + ((sk[113]) & (!g4) & (g27) & (g725)) + ((sk[113]) & (g4) & (!g27) & (g725)));
	assign g1108 = (((!i_8_) & (!g4) & (!sk[114]) & (g27) & (!g73)) + ((!i_8_) & (!g4) & (!sk[114]) & (g27) & (g73)) + ((!i_8_) & (g4) & (!sk[114]) & (g27) & (!g73)) + ((!i_8_) & (g4) & (!sk[114]) & (g27) & (g73)) + ((i_8_) & (!g4) & (!sk[114]) & (g27) & (!g73)) + ((i_8_) & (!g4) & (!sk[114]) & (g27) & (g73)) + ((i_8_) & (g4) & (!sk[114]) & (g27) & (!g73)) + ((i_8_) & (g4) & (!sk[114]) & (g27) & (g73)) + ((i_8_) & (g4) & (sk[114]) & (g27) & (g73)));
	assign g1109 = (((!g74) & (!g847) & (!g934) & (!g1107) & (!g1041) & (!g1108)) + ((!g74) & (!g847) & (!g934) & (!g1107) & (g1041) & (!g1108)) + ((!g74) & (!g847) & (!g934) & (g1107) & (!g1041) & (!g1108)) + ((!g74) & (!g847) & (!g934) & (g1107) & (g1041) & (!g1108)) + ((!g74) & (!g847) & (g934) & (!g1107) & (!g1041) & (!g1108)) + ((!g74) & (!g847) & (g934) & (!g1107) & (g1041) & (!g1108)) + ((!g74) & (!g847) & (g934) & (g1107) & (!g1041) & (!g1108)) + ((!g74) & (!g847) & (g934) & (g1107) & (g1041) & (!g1108)) + ((!g74) & (g847) & (!g934) & (!g1107) & (!g1041) & (!g1108)) + ((!g74) & (g847) & (!g934) & (!g1107) & (g1041) & (!g1108)) + ((!g74) & (g847) & (!g934) & (g1107) & (!g1041) & (!g1108)) + ((!g74) & (g847) & (!g934) & (g1107) & (g1041) & (!g1108)) + ((!g74) & (g847) & (g934) & (!g1107) & (!g1041) & (!g1108)) + ((!g74) & (g847) & (g934) & (!g1107) & (g1041) & (!g1108)) + ((!g74) & (g847) & (g934) & (g1107) & (!g1041) & (!g1108)) + ((!g74) & (g847) & (g934) & (g1107) & (g1041) & (!g1108)) + ((g74) & (g847) & (g934) & (g1107) & (g1041) & (!g1108)));
	assign g1110 = (((!sk[116]) & (!g102) & (!g337) & (g605) & (!g635) & (g858)) + ((!sk[116]) & (!g102) & (!g337) & (g605) & (g635) & (!g858)) + ((!sk[116]) & (!g102) & (!g337) & (g605) & (g635) & (g858)) + ((!sk[116]) & (!g102) & (g337) & (!g605) & (!g635) & (!g858)) + ((!sk[116]) & (!g102) & (g337) & (!g605) & (!g635) & (g858)) + ((!sk[116]) & (!g102) & (g337) & (!g605) & (g635) & (!g858)) + ((!sk[116]) & (!g102) & (g337) & (!g605) & (g635) & (g858)) + ((!sk[116]) & (!g102) & (g337) & (g605) & (!g635) & (!g858)) + ((!sk[116]) & (!g102) & (g337) & (g605) & (!g635) & (g858)) + ((!sk[116]) & (!g102) & (g337) & (g605) & (g635) & (!g858)) + ((!sk[116]) & (!g102) & (g337) & (g605) & (g635) & (g858)) + ((!sk[116]) & (g102) & (!g337) & (g605) & (!g635) & (g858)) + ((!sk[116]) & (g102) & (!g337) & (g605) & (g635) & (!g858)) + ((!sk[116]) & (g102) & (!g337) & (g605) & (g635) & (g858)) + ((!sk[116]) & (g102) & (g337) & (!g605) & (!g635) & (!g858)) + ((!sk[116]) & (g102) & (g337) & (!g605) & (!g635) & (g858)) + ((!sk[116]) & (g102) & (g337) & (!g605) & (g635) & (!g858)) + ((!sk[116]) & (g102) & (g337) & (!g605) & (g635) & (g858)) + ((!sk[116]) & (g102) & (g337) & (g605) & (!g635) & (!g858)) + ((!sk[116]) & (g102) & (g337) & (g605) & (!g635) & (g858)) + ((!sk[116]) & (g102) & (g337) & (g605) & (g635) & (!g858)) + ((!sk[116]) & (g102) & (g337) & (g605) & (g635) & (g858)) + ((sk[116]) & (!g102) & (!g337) & (!g605) & (!g635) & (!g858)) + ((sk[116]) & (!g102) & (!g337) & (!g605) & (g635) & (!g858)) + ((sk[116]) & (!g102) & (!g337) & (g605) & (!g635) & (!g858)) + ((sk[116]) & (!g102) & (!g337) & (g605) & (g635) & (!g858)) + ((sk[116]) & (!g102) & (g337) & (!g605) & (!g635) & (!g858)) + ((sk[116]) & (!g102) & (g337) & (!g605) & (g635) & (!g858)) + ((sk[116]) & (!g102) & (g337) & (g605) & (!g635) & (!g858)) + ((sk[116]) & (!g102) & (g337) & (g605) & (g635) & (!g858)) + ((sk[116]) & (g102) & (!g337) & (!g605) & (!g635) & (!g858)));
	assign g1111 = (((!sk[117]) & (!i_8_) & (!g48) & (g73) & (!g337) & (g605)) + ((!sk[117]) & (!i_8_) & (!g48) & (g73) & (g337) & (!g605)) + ((!sk[117]) & (!i_8_) & (!g48) & (g73) & (g337) & (g605)) + ((!sk[117]) & (!i_8_) & (g48) & (!g73) & (!g337) & (!g605)) + ((!sk[117]) & (!i_8_) & (g48) & (!g73) & (!g337) & (g605)) + ((!sk[117]) & (!i_8_) & (g48) & (!g73) & (g337) & (!g605)) + ((!sk[117]) & (!i_8_) & (g48) & (!g73) & (g337) & (g605)) + ((!sk[117]) & (!i_8_) & (g48) & (g73) & (!g337) & (!g605)) + ((!sk[117]) & (!i_8_) & (g48) & (g73) & (!g337) & (g605)) + ((!sk[117]) & (!i_8_) & (g48) & (g73) & (g337) & (!g605)) + ((!sk[117]) & (!i_8_) & (g48) & (g73) & (g337) & (g605)) + ((!sk[117]) & (i_8_) & (!g48) & (g73) & (!g337) & (g605)) + ((!sk[117]) & (i_8_) & (!g48) & (g73) & (g337) & (!g605)) + ((!sk[117]) & (i_8_) & (!g48) & (g73) & (g337) & (g605)) + ((!sk[117]) & (i_8_) & (g48) & (!g73) & (!g337) & (!g605)) + ((!sk[117]) & (i_8_) & (g48) & (!g73) & (!g337) & (g605)) + ((!sk[117]) & (i_8_) & (g48) & (!g73) & (g337) & (!g605)) + ((!sk[117]) & (i_8_) & (g48) & (!g73) & (g337) & (g605)) + ((!sk[117]) & (i_8_) & (g48) & (g73) & (!g337) & (!g605)) + ((!sk[117]) & (i_8_) & (g48) & (g73) & (!g337) & (g605)) + ((!sk[117]) & (i_8_) & (g48) & (g73) & (g337) & (!g605)) + ((!sk[117]) & (i_8_) & (g48) & (g73) & (g337) & (g605)) + ((sk[117]) & (!i_8_) & (!g48) & (g73) & (!g337) & (g605)) + ((sk[117]) & (!i_8_) & (!g48) & (g73) & (g337) & (!g605)) + ((sk[117]) & (!i_8_) & (!g48) & (g73) & (g337) & (g605)) + ((sk[117]) & (!i_8_) & (g48) & (g73) & (!g337) & (g605)) + ((sk[117]) & (!i_8_) & (g48) & (g73) & (g337) & (!g605)) + ((sk[117]) & (!i_8_) & (g48) & (g73) & (g337) & (g605)) + ((sk[117]) & (i_8_) & (g48) & (g73) & (!g337) & (!g605)) + ((sk[117]) & (i_8_) & (g48) & (g73) & (!g337) & (g605)) + ((sk[117]) & (i_8_) & (g48) & (g73) & (g337) & (!g605)) + ((sk[117]) & (i_8_) & (g48) & (g73) & (g337) & (g605)));
	assign g1112 = (((!g75) & (!g725) & (g1029) & (!sk[118]) & (!g1111)) + ((!g75) & (!g725) & (g1029) & (!sk[118]) & (g1111)) + ((!g75) & (g725) & (g1029) & (!sk[118]) & (!g1111)) + ((!g75) & (g725) & (g1029) & (!sk[118]) & (g1111)) + ((!g75) & (g725) & (g1029) & (sk[118]) & (!g1111)) + ((g75) & (!g725) & (!g1029) & (sk[118]) & (!g1111)) + ((g75) & (!g725) & (g1029) & (!sk[118]) & (!g1111)) + ((g75) & (!g725) & (g1029) & (!sk[118]) & (g1111)) + ((g75) & (!g725) & (g1029) & (sk[118]) & (!g1111)) + ((g75) & (g725) & (!g1029) & (sk[118]) & (!g1111)) + ((g75) & (g725) & (g1029) & (!sk[118]) & (!g1111)) + ((g75) & (g725) & (g1029) & (!sk[118]) & (g1111)) + ((g75) & (g725) & (g1029) & (sk[118]) & (!g1111)));
	assign g1113 = (((g1460) & (g1101) & (g1106) & (g1109) & (g1110) & (g1112)));
	assign g1114 = (((!sk[120]) & (!g496) & (!g738) & (g1102) & (!g1033)) + ((!sk[120]) & (!g496) & (!g738) & (g1102) & (g1033)) + ((!sk[120]) & (!g496) & (g738) & (g1102) & (!g1033)) + ((!sk[120]) & (!g496) & (g738) & (g1102) & (g1033)) + ((!sk[120]) & (g496) & (!g738) & (g1102) & (!g1033)) + ((!sk[120]) & (g496) & (!g738) & (g1102) & (g1033)) + ((!sk[120]) & (g496) & (g738) & (g1102) & (!g1033)) + ((!sk[120]) & (g496) & (g738) & (g1102) & (g1033)) + ((sk[120]) & (!g496) & (!g738) & (!g1102) & (g1033)));
	assign g1115 = (((!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (!g75) & (g429)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g75) & (g429)) + ((!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g75) & (g429)) + ((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g75) & (g429)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g75) & (g429)) + ((i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (!g75) & (g429)) + ((i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (!g75) & (g429)) + ((i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (!g75) & (g429)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g75) & (g429)) + ((i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g75) & (g429)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g75) & (g429)) + ((i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g75) & (g429)));
	assign g1116 = (((!i_8_) & (!g73) & (!g993) & (!g927) & (!g1114) & (!g1115)) + ((!i_8_) & (!g73) & (!g993) & (!g927) & (g1114) & (!g1115)) + ((!i_8_) & (!g73) & (!g993) & (g927) & (!g1114) & (!g1115)) + ((!i_8_) & (!g73) & (!g993) & (g927) & (g1114) & (!g1115)) + ((!i_8_) & (!g73) & (g993) & (!g927) & (!g1114) & (!g1115)) + ((!i_8_) & (!g73) & (g993) & (!g927) & (g1114) & (!g1115)) + ((!i_8_) & (!g73) & (g993) & (g927) & (!g1114) & (!g1115)) + ((!i_8_) & (!g73) & (g993) & (g927) & (g1114) & (!g1115)) + ((!i_8_) & (g73) & (!g993) & (!g927) & (g1114) & (!g1115)) + ((i_8_) & (!g73) & (!g993) & (!g927) & (!g1114) & (!g1115)) + ((i_8_) & (!g73) & (!g993) & (!g927) & (g1114) & (!g1115)) + ((i_8_) & (!g73) & (!g993) & (g927) & (!g1114) & (!g1115)) + ((i_8_) & (!g73) & (!g993) & (g927) & (g1114) & (!g1115)) + ((i_8_) & (!g73) & (g993) & (!g927) & (!g1114) & (!g1115)) + ((i_8_) & (!g73) & (g993) & (!g927) & (g1114) & (!g1115)) + ((i_8_) & (!g73) & (g993) & (g927) & (!g1114) & (!g1115)) + ((i_8_) & (!g73) & (g993) & (g927) & (g1114) & (!g1115)) + ((i_8_) & (g73) & (!g993) & (!g927) & (!g1114) & (!g1115)) + ((i_8_) & (g73) & (!g993) & (!g927) & (g1114) & (!g1115)));
	assign g1117 = (((g285) & (g589) & (g530) & (g1099) & (g1113) & (g1116)));
	assign g1118 = (((!g24) & (!g35) & (!sk[124]) & (g1090)) + ((!g24) & (g35) & (!sk[124]) & (!g1090)) + ((!g24) & (g35) & (!sk[124]) & (g1090)) + ((!g24) & (g35) & (sk[124]) & (!g1090)) + ((g24) & (!g35) & (!sk[124]) & (g1090)) + ((g24) & (g35) & (!sk[124]) & (!g1090)) + ((g24) & (g35) & (!sk[124]) & (g1090)));
	assign g1119 = (((!g25) & (!g42) & (!g40) & (g1081) & (!g1118) & (g1088)) + ((!g25) & (!g42) & (g40) & (g1081) & (!g1118) & (g1088)) + ((!g25) & (g42) & (!g40) & (g1081) & (!g1118) & (g1088)) + ((g25) & (!g42) & (!g40) & (!g1081) & (!g1118) & (g1088)) + ((g25) & (!g42) & (!g40) & (g1081) & (!g1118) & (g1088)) + ((g25) & (!g42) & (g40) & (!g1081) & (!g1118) & (g1088)) + ((g25) & (!g42) & (g40) & (g1081) & (!g1118) & (g1088)) + ((g25) & (g42) & (!g40) & (!g1081) & (!g1118) & (g1088)) + ((g25) & (g42) & (!g40) & (g1081) & (!g1118) & (g1088)));
	assign o_30_ = (((!g100) & (!sk[126]) & (!g711) & (g961) & (!g1117) & (g1119)) + ((!g100) & (!sk[126]) & (!g711) & (g961) & (g1117) & (!g1119)) + ((!g100) & (!sk[126]) & (!g711) & (g961) & (g1117) & (g1119)) + ((!g100) & (!sk[126]) & (g711) & (!g961) & (!g1117) & (!g1119)) + ((!g100) & (!sk[126]) & (g711) & (!g961) & (!g1117) & (g1119)) + ((!g100) & (!sk[126]) & (g711) & (!g961) & (g1117) & (!g1119)) + ((!g100) & (!sk[126]) & (g711) & (!g961) & (g1117) & (g1119)) + ((!g100) & (!sk[126]) & (g711) & (g961) & (!g1117) & (!g1119)) + ((!g100) & (!sk[126]) & (g711) & (g961) & (!g1117) & (g1119)) + ((!g100) & (!sk[126]) & (g711) & (g961) & (g1117) & (!g1119)) + ((!g100) & (!sk[126]) & (g711) & (g961) & (g1117) & (g1119)) + ((!g100) & (sk[126]) & (!g711) & (!g961) & (!g1117) & (!g1119)) + ((!g100) & (sk[126]) & (!g711) & (!g961) & (!g1117) & (g1119)) + ((!g100) & (sk[126]) & (!g711) & (!g961) & (g1117) & (!g1119)) + ((!g100) & (sk[126]) & (!g711) & (!g961) & (g1117) & (g1119)) + ((!g100) & (sk[126]) & (!g711) & (g961) & (!g1117) & (!g1119)) + ((!g100) & (sk[126]) & (!g711) & (g961) & (!g1117) & (g1119)) + ((!g100) & (sk[126]) & (!g711) & (g961) & (g1117) & (!g1119)) + ((!g100) & (sk[126]) & (!g711) & (g961) & (g1117) & (g1119)) + ((!g100) & (sk[126]) & (g711) & (!g961) & (!g1117) & (!g1119)) + ((!g100) & (sk[126]) & (g711) & (!g961) & (!g1117) & (g1119)) + ((!g100) & (sk[126]) & (g711) & (!g961) & (g1117) & (!g1119)) + ((!g100) & (sk[126]) & (g711) & (!g961) & (g1117) & (g1119)) + ((!g100) & (sk[126]) & (g711) & (g961) & (!g1117) & (!g1119)) + ((!g100) & (sk[126]) & (g711) & (g961) & (!g1117) & (g1119)) + ((!g100) & (sk[126]) & (g711) & (g961) & (g1117) & (!g1119)) + ((!g100) & (sk[126]) & (g711) & (g961) & (g1117) & (g1119)) + ((g100) & (!sk[126]) & (!g711) & (g961) & (!g1117) & (g1119)) + ((g100) & (!sk[126]) & (!g711) & (g961) & (g1117) & (!g1119)) + ((g100) & (!sk[126]) & (!g711) & (g961) & (g1117) & (g1119)) + ((g100) & (!sk[126]) & (g711) & (!g961) & (!g1117) & (!g1119)) + ((g100) & (!sk[126]) & (g711) & (!g961) & (!g1117) & (g1119)) + ((g100) & (!sk[126]) & (g711) & (!g961) & (g1117) & (!g1119)) + ((g100) & (!sk[126]) & (g711) & (!g961) & (g1117) & (g1119)) + ((g100) & (!sk[126]) & (g711) & (g961) & (!g1117) & (!g1119)) + ((g100) & (!sk[126]) & (g711) & (g961) & (!g1117) & (g1119)) + ((g100) & (!sk[126]) & (g711) & (g961) & (g1117) & (!g1119)) + ((g100) & (!sk[126]) & (g711) & (g961) & (g1117) & (g1119)) + ((g100) & (sk[126]) & (!g711) & (!g961) & (!g1117) & (!g1119)) + ((g100) & (sk[126]) & (!g711) & (!g961) & (!g1117) & (g1119)) + ((g100) & (sk[126]) & (!g711) & (!g961) & (g1117) & (!g1119)) + ((g100) & (sk[126]) & (!g711) & (!g961) & (g1117) & (g1119)) + ((g100) & (sk[126]) & (!g711) & (g961) & (!g1117) & (!g1119)) + ((g100) & (sk[126]) & (!g711) & (g961) & (!g1117) & (g1119)) + ((g100) & (sk[126]) & (!g711) & (g961) & (g1117) & (!g1119)) + ((g100) & (sk[126]) & (!g711) & (g961) & (g1117) & (g1119)) + ((g100) & (sk[126]) & (g711) & (!g961) & (!g1117) & (!g1119)) + ((g100) & (sk[126]) & (g711) & (!g961) & (!g1117) & (g1119)) + ((g100) & (sk[126]) & (g711) & (!g961) & (g1117) & (!g1119)) + ((g100) & (sk[126]) & (g711) & (!g961) & (g1117) & (g1119)) + ((g100) & (sk[126]) & (g711) & (g961) & (!g1117) & (!g1119)) + ((g100) & (sk[126]) & (g711) & (g961) & (!g1117) & (g1119)) + ((g100) & (sk[126]) & (g711) & (g961) & (g1117) & (!g1119)));
	assign o_31_ = (((!i_6_) & (!i_7_) & (i_4_) & (i_3_) & (i_5_) & (g14)) + ((!i_6_) & (i_7_) & (!i_4_) & (!i_3_) & (!i_5_) & (g14)) + ((!i_6_) & (i_7_) & (i_4_) & (!i_3_) & (!i_5_) & (g14)) + ((i_6_) & (i_7_) & (!i_4_) & (!i_3_) & (!i_5_) & (g14)) + ((i_6_) & (i_7_) & (i_4_) & (!i_3_) & (!i_5_) & (g14)) + ((i_6_) & (i_7_) & (i_4_) & (i_3_) & (!i_5_) & (g14)) + ((i_6_) & (i_7_) & (i_4_) & (i_3_) & (i_5_) & (g14)));
	assign g1122 = (((!g1) & (!i_4_) & (!sk[0]) & (i_3_) & (!i_5_) & (g14)) + ((!g1) & (!i_4_) & (!sk[0]) & (i_3_) & (i_5_) & (!g14)) + ((!g1) & (!i_4_) & (!sk[0]) & (i_3_) & (i_5_) & (g14)) + ((!g1) & (i_4_) & (!sk[0]) & (!i_3_) & (!i_5_) & (!g14)) + ((!g1) & (i_4_) & (!sk[0]) & (!i_3_) & (!i_5_) & (g14)) + ((!g1) & (i_4_) & (!sk[0]) & (!i_3_) & (i_5_) & (!g14)) + ((!g1) & (i_4_) & (!sk[0]) & (!i_3_) & (i_5_) & (g14)) + ((!g1) & (i_4_) & (!sk[0]) & (i_3_) & (!i_5_) & (!g14)) + ((!g1) & (i_4_) & (!sk[0]) & (i_3_) & (!i_5_) & (g14)) + ((!g1) & (i_4_) & (!sk[0]) & (i_3_) & (i_5_) & (!g14)) + ((!g1) & (i_4_) & (!sk[0]) & (i_3_) & (i_5_) & (g14)) + ((g1) & (!i_4_) & (!sk[0]) & (i_3_) & (!i_5_) & (g14)) + ((g1) & (!i_4_) & (!sk[0]) & (i_3_) & (i_5_) & (!g14)) + ((g1) & (!i_4_) & (!sk[0]) & (i_3_) & (i_5_) & (g14)) + ((g1) & (i_4_) & (!sk[0]) & (!i_3_) & (!i_5_) & (!g14)) + ((g1) & (i_4_) & (!sk[0]) & (!i_3_) & (!i_5_) & (g14)) + ((g1) & (i_4_) & (!sk[0]) & (!i_3_) & (i_5_) & (!g14)) + ((g1) & (i_4_) & (!sk[0]) & (!i_3_) & (i_5_) & (g14)) + ((g1) & (i_4_) & (!sk[0]) & (i_3_) & (!i_5_) & (!g14)) + ((g1) & (i_4_) & (!sk[0]) & (i_3_) & (!i_5_) & (g14)) + ((g1) & (i_4_) & (!sk[0]) & (i_3_) & (i_5_) & (!g14)) + ((g1) & (i_4_) & (!sk[0]) & (i_3_) & (i_5_) & (g14)) + ((g1) & (i_4_) & (sk[0]) & (i_3_) & (i_5_) & (g14)));
	assign g1123 = (((!g43) & (!g38) & (!g55) & (sk[1]) & (!g57) & (!g1122)) + ((!g43) & (!g38) & (g55) & (!sk[1]) & (!g57) & (g1122)) + ((!g43) & (!g38) & (g55) & (!sk[1]) & (g57) & (!g1122)) + ((!g43) & (!g38) & (g55) & (!sk[1]) & (g57) & (g1122)) + ((!g43) & (!g38) & (g55) & (sk[1]) & (!g57) & (!g1122)) + ((!g43) & (g38) & (!g55) & (!sk[1]) & (!g57) & (!g1122)) + ((!g43) & (g38) & (!g55) & (!sk[1]) & (!g57) & (g1122)) + ((!g43) & (g38) & (!g55) & (!sk[1]) & (g57) & (!g1122)) + ((!g43) & (g38) & (!g55) & (!sk[1]) & (g57) & (g1122)) + ((!g43) & (g38) & (!g55) & (sk[1]) & (!g57) & (!g1122)) + ((!g43) & (g38) & (g55) & (!sk[1]) & (!g57) & (!g1122)) + ((!g43) & (g38) & (g55) & (!sk[1]) & (!g57) & (g1122)) + ((!g43) & (g38) & (g55) & (!sk[1]) & (g57) & (!g1122)) + ((!g43) & (g38) & (g55) & (!sk[1]) & (g57) & (g1122)) + ((!g43) & (g38) & (g55) & (sk[1]) & (!g57) & (!g1122)) + ((g43) & (!g38) & (!g55) & (sk[1]) & (!g57) & (!g1122)) + ((g43) & (!g38) & (g55) & (!sk[1]) & (!g57) & (g1122)) + ((g43) & (!g38) & (g55) & (!sk[1]) & (g57) & (!g1122)) + ((g43) & (!g38) & (g55) & (!sk[1]) & (g57) & (g1122)) + ((g43) & (g38) & (!g55) & (!sk[1]) & (!g57) & (!g1122)) + ((g43) & (g38) & (!g55) & (!sk[1]) & (!g57) & (g1122)) + ((g43) & (g38) & (!g55) & (!sk[1]) & (g57) & (!g1122)) + ((g43) & (g38) & (!g55) & (!sk[1]) & (g57) & (g1122)) + ((g43) & (g38) & (!g55) & (sk[1]) & (!g57) & (!g1122)) + ((g43) & (g38) & (g55) & (!sk[1]) & (!g57) & (!g1122)) + ((g43) & (g38) & (g55) & (!sk[1]) & (!g57) & (g1122)) + ((g43) & (g38) & (g55) & (!sk[1]) & (g57) & (!g1122)) + ((g43) & (g38) & (g55) & (!sk[1]) & (g57) & (g1122)) + ((g43) & (g38) & (g55) & (sk[1]) & (!g57) & (!g1122)));
	assign g1124 = (((!g38) & (!g1067) & (!sk[2]) & (g1068) & (!g1069) & (g1074)) + ((!g38) & (!g1067) & (!sk[2]) & (g1068) & (g1069) & (!g1074)) + ((!g38) & (!g1067) & (!sk[2]) & (g1068) & (g1069) & (g1074)) + ((!g38) & (!g1067) & (sk[2]) & (!g1068) & (!g1069) & (g1074)) + ((!g38) & (g1067) & (!sk[2]) & (!g1068) & (!g1069) & (!g1074)) + ((!g38) & (g1067) & (!sk[2]) & (!g1068) & (!g1069) & (g1074)) + ((!g38) & (g1067) & (!sk[2]) & (!g1068) & (g1069) & (!g1074)) + ((!g38) & (g1067) & (!sk[2]) & (!g1068) & (g1069) & (g1074)) + ((!g38) & (g1067) & (!sk[2]) & (g1068) & (!g1069) & (!g1074)) + ((!g38) & (g1067) & (!sk[2]) & (g1068) & (!g1069) & (g1074)) + ((!g38) & (g1067) & (!sk[2]) & (g1068) & (g1069) & (!g1074)) + ((!g38) & (g1067) & (!sk[2]) & (g1068) & (g1069) & (g1074)) + ((!g38) & (g1067) & (sk[2]) & (!g1068) & (!g1069) & (g1074)) + ((!g38) & (g1067) & (sk[2]) & (g1068) & (!g1069) & (g1074)) + ((g38) & (!g1067) & (!sk[2]) & (g1068) & (!g1069) & (g1074)) + ((g38) & (!g1067) & (!sk[2]) & (g1068) & (g1069) & (!g1074)) + ((g38) & (!g1067) & (!sk[2]) & (g1068) & (g1069) & (g1074)) + ((g38) & (!g1067) & (sk[2]) & (!g1068) & (!g1069) & (g1074)) + ((g38) & (g1067) & (!sk[2]) & (!g1068) & (!g1069) & (!g1074)) + ((g38) & (g1067) & (!sk[2]) & (!g1068) & (!g1069) & (g1074)) + ((g38) & (g1067) & (!sk[2]) & (!g1068) & (g1069) & (!g1074)) + ((g38) & (g1067) & (!sk[2]) & (!g1068) & (g1069) & (g1074)) + ((g38) & (g1067) & (!sk[2]) & (g1068) & (!g1069) & (!g1074)) + ((g38) & (g1067) & (!sk[2]) & (g1068) & (!g1069) & (g1074)) + ((g38) & (g1067) & (!sk[2]) & (g1068) & (g1069) & (!g1074)) + ((g38) & (g1067) & (!sk[2]) & (g1068) & (g1069) & (g1074)) + ((g38) & (g1067) & (sk[2]) & (!g1068) & (!g1069) & (g1074)) + ((g38) & (g1067) & (sk[2]) & (!g1068) & (g1069) & (g1074)) + ((g38) & (g1067) & (sk[2]) & (g1068) & (!g1069) & (g1074)) + ((g38) & (g1067) & (sk[2]) & (g1068) & (g1069) & (g1074)));
	assign g1125 = (((g100) & (g711) & (g961) & (g1117) & (g1123) & (g1124)));
	assign g1126 = (((!sk[4]) & (g38) & (!g1067)) + ((!sk[4]) & (g38) & (g1067)) + ((sk[4]) & (g38) & (g1067)));
	assign g1127 = (((!g6) & (!sk[5]) & (!g14) & (g43) & (!g1126)) + ((!g6) & (!sk[5]) & (!g14) & (g43) & (g1126)) + ((!g6) & (!sk[5]) & (g14) & (g43) & (!g1126)) + ((!g6) & (!sk[5]) & (g14) & (g43) & (g1126)) + ((g6) & (!sk[5]) & (!g14) & (g43) & (!g1126)) + ((g6) & (!sk[5]) & (!g14) & (g43) & (g1126)) + ((g6) & (!sk[5]) & (g14) & (g43) & (!g1126)) + ((g6) & (!sk[5]) & (g14) & (g43) & (g1126)) + ((g6) & (sk[5]) & (g14) & (g43) & (!g1126)));
	assign g1128 = (((!g44) & (!g41) & (g1127) & (!sk[6]) & (!g1076)) + ((!g44) & (!g41) & (g1127) & (!sk[6]) & (g1076)) + ((!g44) & (g41) & (!g1127) & (sk[6]) & (g1076)) + ((!g44) & (g41) & (g1127) & (!sk[6]) & (!g1076)) + ((!g44) & (g41) & (g1127) & (!sk[6]) & (g1076)) + ((g44) & (!g41) & (g1127) & (!sk[6]) & (!g1076)) + ((g44) & (!g41) & (g1127) & (!sk[6]) & (g1076)) + ((g44) & (g41) & (g1127) & (!sk[6]) & (!g1076)) + ((g44) & (g41) & (g1127) & (!sk[6]) & (g1076)));
	assign g1129 = (((!g100) & (!g711) & (!sk[7]) & (g961) & (!g1117)) + ((!g100) & (!g711) & (!sk[7]) & (g961) & (g1117)) + ((!g100) & (g711) & (!sk[7]) & (g961) & (!g1117)) + ((!g100) & (g711) & (!sk[7]) & (g961) & (g1117)) + ((g100) & (!g711) & (!sk[7]) & (g961) & (!g1117)) + ((g100) & (!g711) & (!sk[7]) & (g961) & (g1117)) + ((g100) & (g711) & (!sk[7]) & (g961) & (!g1117)) + ((g100) & (g711) & (!sk[7]) & (g961) & (g1117)) + ((g100) & (g711) & (sk[7]) & (g961) & (g1117)));
	assign g1130 = (((!i_8_) & (!g73) & (g112) & (!g636) & (!sk[8]) & (g857)) + ((!i_8_) & (!g73) & (g112) & (g636) & (!sk[8]) & (!g857)) + ((!i_8_) & (!g73) & (g112) & (g636) & (!sk[8]) & (g857)) + ((!i_8_) & (!g73) & (g112) & (g636) & (sk[8]) & (!g857)) + ((!i_8_) & (!g73) & (g112) & (g636) & (sk[8]) & (g857)) + ((!i_8_) & (g73) & (!g112) & (!g636) & (!sk[8]) & (!g857)) + ((!i_8_) & (g73) & (!g112) & (!g636) & (!sk[8]) & (g857)) + ((!i_8_) & (g73) & (!g112) & (g636) & (!sk[8]) & (!g857)) + ((!i_8_) & (g73) & (!g112) & (g636) & (!sk[8]) & (g857)) + ((!i_8_) & (g73) & (g112) & (!g636) & (!sk[8]) & (!g857)) + ((!i_8_) & (g73) & (g112) & (!g636) & (!sk[8]) & (g857)) + ((!i_8_) & (g73) & (g112) & (g636) & (!sk[8]) & (!g857)) + ((!i_8_) & (g73) & (g112) & (g636) & (!sk[8]) & (g857)) + ((!i_8_) & (g73) & (g112) & (g636) & (sk[8]) & (!g857)) + ((!i_8_) & (g73) & (g112) & (g636) & (sk[8]) & (g857)) + ((i_8_) & (!g73) & (g112) & (!g636) & (!sk[8]) & (g857)) + ((i_8_) & (!g73) & (g112) & (g636) & (!sk[8]) & (!g857)) + ((i_8_) & (!g73) & (g112) & (g636) & (!sk[8]) & (g857)) + ((i_8_) & (!g73) & (g112) & (g636) & (sk[8]) & (!g857)) + ((i_8_) & (!g73) & (g112) & (g636) & (sk[8]) & (g857)) + ((i_8_) & (g73) & (!g112) & (!g636) & (!sk[8]) & (!g857)) + ((i_8_) & (g73) & (!g112) & (!g636) & (!sk[8]) & (g857)) + ((i_8_) & (g73) & (!g112) & (!g636) & (sk[8]) & (g857)) + ((i_8_) & (g73) & (!g112) & (g636) & (!sk[8]) & (!g857)) + ((i_8_) & (g73) & (!g112) & (g636) & (!sk[8]) & (g857)) + ((i_8_) & (g73) & (!g112) & (g636) & (sk[8]) & (g857)) + ((i_8_) & (g73) & (g112) & (!g636) & (!sk[8]) & (!g857)) + ((i_8_) & (g73) & (g112) & (!g636) & (!sk[8]) & (g857)) + ((i_8_) & (g73) & (g112) & (!g636) & (sk[8]) & (g857)) + ((i_8_) & (g73) & (g112) & (g636) & (!sk[8]) & (!g857)) + ((i_8_) & (g73) & (g112) & (g636) & (!sk[8]) & (g857)) + ((i_8_) & (g73) & (g112) & (g636) & (sk[8]) & (!g857)) + ((i_8_) & (g73) & (g112) & (g636) & (sk[8]) & (g857)));
	assign g1131 = (((!sk[9]) & (!g164) & (!g154) & (g974) & (!g1130)) + ((!sk[9]) & (!g164) & (!g154) & (g974) & (g1130)) + ((!sk[9]) & (!g164) & (g154) & (g974) & (!g1130)) + ((!sk[9]) & (!g164) & (g154) & (g974) & (g1130)) + ((!sk[9]) & (g164) & (!g154) & (g974) & (!g1130)) + ((!sk[9]) & (g164) & (!g154) & (g974) & (g1130)) + ((!sk[9]) & (g164) & (g154) & (g974) & (!g1130)) + ((!sk[9]) & (g164) & (g154) & (g974) & (g1130)) + ((sk[9]) & (!g164) & (!g154) & (!g974) & (!g1130)) + ((sk[9]) & (!g164) & (g154) & (!g974) & (!g1130)) + ((sk[9]) & (!g164) & (g154) & (g974) & (!g1130)) + ((sk[9]) & (g164) & (!g154) & (!g974) & (!g1130)) + ((sk[9]) & (g164) & (g154) & (!g974) & (!g1130)));
	assign g1132 = (((!g154) & (!sk[10]) & (!g106) & (g784) & (!g964)) + ((!g154) & (!sk[10]) & (!g106) & (g784) & (g964)) + ((!g154) & (!sk[10]) & (g106) & (g784) & (!g964)) + ((!g154) & (!sk[10]) & (g106) & (g784) & (g964)) + ((!g154) & (sk[10]) & (!g106) & (!g784) & (g964)) + ((g154) & (!sk[10]) & (!g106) & (g784) & (!g964)) + ((g154) & (!sk[10]) & (!g106) & (g784) & (g964)) + ((g154) & (!sk[10]) & (g106) & (g784) & (!g964)) + ((g154) & (!sk[10]) & (g106) & (g784) & (g964)) + ((g154) & (sk[10]) & (!g106) & (!g784) & (!g964)) + ((g154) & (sk[10]) & (!g106) & (!g784) & (g964)));
	assign g1133 = (((!sk[11]) & (!g123) & (!g770) & (g629) & (!g1132)) + ((!sk[11]) & (!g123) & (!g770) & (g629) & (g1132)) + ((!sk[11]) & (!g123) & (g770) & (g629) & (!g1132)) + ((!sk[11]) & (!g123) & (g770) & (g629) & (g1132)) + ((!sk[11]) & (g123) & (!g770) & (g629) & (!g1132)) + ((!sk[11]) & (g123) & (!g770) & (g629) & (g1132)) + ((!sk[11]) & (g123) & (g770) & (g629) & (!g1132)) + ((!sk[11]) & (g123) & (g770) & (g629) & (g1132)) + ((sk[11]) & (!g123) & (!g770) & (!g629) & (g1132)) + ((sk[11]) & (g123) & (!g770) & (!g629) & (g1132)) + ((sk[11]) & (g123) & (!g770) & (g629) & (g1132)) + ((sk[11]) & (g123) & (g770) & (!g629) & (g1132)) + ((sk[11]) & (g123) & (g770) & (g629) & (g1132)));
	assign g1134 = (((!g164) & (!g123) & (g597) & (!sk[12]) & (!g628)) + ((!g164) & (!g123) & (g597) & (!sk[12]) & (g628)) + ((!g164) & (!g123) & (g597) & (sk[12]) & (!g628)) + ((!g164) & (!g123) & (g597) & (sk[12]) & (g628)) + ((!g164) & (g123) & (g597) & (!sk[12]) & (!g628)) + ((!g164) & (g123) & (g597) & (!sk[12]) & (g628)) + ((g164) & (!g123) & (!g597) & (sk[12]) & (!g628)) + ((g164) & (!g123) & (g597) & (!sk[12]) & (!g628)) + ((g164) & (!g123) & (g597) & (!sk[12]) & (g628)) + ((g164) & (!g123) & (g597) & (sk[12]) & (!g628)) + ((g164) & (!g123) & (g597) & (sk[12]) & (g628)) + ((g164) & (g123) & (!g597) & (sk[12]) & (!g628)) + ((g164) & (g123) & (g597) & (!sk[12]) & (!g628)) + ((g164) & (g123) & (g597) & (!sk[12]) & (g628)) + ((g164) & (g123) & (g597) & (sk[12]) & (!g628)));
	assign g1135 = (((!g75) & (!g182) & (!g183) & (!g582) & (!g976) & (!g1134)) + ((g75) & (!g182) & (!g183) & (!g582) & (!g976) & (!g1134)) + ((g75) & (!g182) & (g183) & (!g582) & (!g976) & (!g1134)) + ((g75) & (g182) & (!g183) & (!g582) & (!g976) & (!g1134)) + ((g75) & (g182) & (g183) & (!g582) & (!g976) & (!g1134)));
	assign g1136 = (((!g24) & (!sk[14]) & (!g75) & (g68) & (!g83)) + ((!g24) & (!sk[14]) & (!g75) & (g68) & (g83)) + ((!g24) & (!sk[14]) & (g75) & (g68) & (!g83)) + ((!g24) & (!sk[14]) & (g75) & (g68) & (g83)) + ((!g24) & (sk[14]) & (!g75) & (!g68) & (g83)) + ((!g24) & (sk[14]) & (!g75) & (g68) & (g83)) + ((g24) & (!sk[14]) & (!g75) & (g68) & (!g83)) + ((g24) & (!sk[14]) & (!g75) & (g68) & (g83)) + ((g24) & (!sk[14]) & (g75) & (g68) & (!g83)) + ((g24) & (!sk[14]) & (g75) & (g68) & (g83)) + ((g24) & (sk[14]) & (!g75) & (!g68) & (g83)));
	assign g1137 = (((!i_8_) & (!i_6_) & (i_7_) & (!sk[15]) & (!g445) & (g394)) + ((!i_8_) & (!i_6_) & (i_7_) & (!sk[15]) & (g445) & (!g394)) + ((!i_8_) & (!i_6_) & (i_7_) & (!sk[15]) & (g445) & (g394)) + ((!i_8_) & (i_6_) & (!i_7_) & (!sk[15]) & (!g445) & (!g394)) + ((!i_8_) & (i_6_) & (!i_7_) & (!sk[15]) & (!g445) & (g394)) + ((!i_8_) & (i_6_) & (!i_7_) & (!sk[15]) & (g445) & (!g394)) + ((!i_8_) & (i_6_) & (!i_7_) & (!sk[15]) & (g445) & (g394)) + ((!i_8_) & (i_6_) & (i_7_) & (!sk[15]) & (!g445) & (!g394)) + ((!i_8_) & (i_6_) & (i_7_) & (!sk[15]) & (!g445) & (g394)) + ((!i_8_) & (i_6_) & (i_7_) & (!sk[15]) & (g445) & (!g394)) + ((!i_8_) & (i_6_) & (i_7_) & (!sk[15]) & (g445) & (g394)) + ((i_8_) & (!i_6_) & (i_7_) & (!sk[15]) & (!g445) & (g394)) + ((i_8_) & (!i_6_) & (i_7_) & (!sk[15]) & (g445) & (!g394)) + ((i_8_) & (!i_6_) & (i_7_) & (!sk[15]) & (g445) & (g394)) + ((i_8_) & (!i_6_) & (i_7_) & (sk[15]) & (g445) & (g394)) + ((i_8_) & (i_6_) & (!i_7_) & (!sk[15]) & (!g445) & (!g394)) + ((i_8_) & (i_6_) & (!i_7_) & (!sk[15]) & (!g445) & (g394)) + ((i_8_) & (i_6_) & (!i_7_) & (!sk[15]) & (g445) & (!g394)) + ((i_8_) & (i_6_) & (!i_7_) & (!sk[15]) & (g445) & (g394)) + ((i_8_) & (i_6_) & (!i_7_) & (sk[15]) & (g445) & (g394)) + ((i_8_) & (i_6_) & (i_7_) & (!sk[15]) & (!g445) & (!g394)) + ((i_8_) & (i_6_) & (i_7_) & (!sk[15]) & (!g445) & (g394)) + ((i_8_) & (i_6_) & (i_7_) & (!sk[15]) & (g445) & (!g394)) + ((i_8_) & (i_6_) & (i_7_) & (!sk[15]) & (g445) & (g394)) + ((i_8_) & (i_6_) & (i_7_) & (sk[15]) & (g445) & (g394)));
	assign g1138 = (((!sk[16]) & (!g154) & (!g597) & (g628) & (!g629)) + ((!sk[16]) & (!g154) & (!g597) & (g628) & (g629)) + ((!sk[16]) & (!g154) & (g597) & (g628) & (!g629)) + ((!sk[16]) & (!g154) & (g597) & (g628) & (g629)) + ((!sk[16]) & (g154) & (!g597) & (g628) & (!g629)) + ((!sk[16]) & (g154) & (!g597) & (g628) & (g629)) + ((!sk[16]) & (g154) & (g597) & (g628) & (!g629)) + ((!sk[16]) & (g154) & (g597) & (g628) & (g629)) + ((sk[16]) & (!g154) & (!g597) & (!g628) & (!g629)) + ((sk[16]) & (!g154) & (!g597) & (!g628) & (g629)) + ((sk[16]) & (!g154) & (!g597) & (g628) & (g629)) + ((sk[16]) & (!g154) & (g597) & (!g628) & (!g629)) + ((sk[16]) & (!g154) & (g597) & (!g628) & (g629)) + ((sk[16]) & (!g154) & (g597) & (g628) & (!g629)) + ((sk[16]) & (!g154) & (g597) & (g628) & (g629)));
	assign g1139 = (((!i_12_) & (!i_13_) & (!sk[17]) & (i_14_) & (!g122) & (g83)) + ((!i_12_) & (!i_13_) & (!sk[17]) & (i_14_) & (g122) & (!g83)) + ((!i_12_) & (!i_13_) & (!sk[17]) & (i_14_) & (g122) & (g83)) + ((!i_12_) & (!i_13_) & (sk[17]) & (i_14_) & (g122) & (g83)) + ((!i_12_) & (i_13_) & (!sk[17]) & (!i_14_) & (!g122) & (!g83)) + ((!i_12_) & (i_13_) & (!sk[17]) & (!i_14_) & (!g122) & (g83)) + ((!i_12_) & (i_13_) & (!sk[17]) & (!i_14_) & (g122) & (!g83)) + ((!i_12_) & (i_13_) & (!sk[17]) & (!i_14_) & (g122) & (g83)) + ((!i_12_) & (i_13_) & (!sk[17]) & (i_14_) & (!g122) & (!g83)) + ((!i_12_) & (i_13_) & (!sk[17]) & (i_14_) & (!g122) & (g83)) + ((!i_12_) & (i_13_) & (!sk[17]) & (i_14_) & (g122) & (!g83)) + ((!i_12_) & (i_13_) & (!sk[17]) & (i_14_) & (g122) & (g83)) + ((i_12_) & (!i_13_) & (!sk[17]) & (i_14_) & (!g122) & (g83)) + ((i_12_) & (!i_13_) & (!sk[17]) & (i_14_) & (g122) & (!g83)) + ((i_12_) & (!i_13_) & (!sk[17]) & (i_14_) & (g122) & (g83)) + ((i_12_) & (!i_13_) & (sk[17]) & (!i_14_) & (g122) & (g83)) + ((i_12_) & (i_13_) & (!sk[17]) & (!i_14_) & (!g122) & (!g83)) + ((i_12_) & (i_13_) & (!sk[17]) & (!i_14_) & (!g122) & (g83)) + ((i_12_) & (i_13_) & (!sk[17]) & (!i_14_) & (g122) & (!g83)) + ((i_12_) & (i_13_) & (!sk[17]) & (!i_14_) & (g122) & (g83)) + ((i_12_) & (i_13_) & (!sk[17]) & (i_14_) & (!g122) & (!g83)) + ((i_12_) & (i_13_) & (!sk[17]) & (i_14_) & (!g122) & (g83)) + ((i_12_) & (i_13_) & (!sk[17]) & (i_14_) & (g122) & (!g83)) + ((i_12_) & (i_13_) & (!sk[17]) & (i_14_) & (g122) & (g83)) + ((i_12_) & (i_13_) & (sk[17]) & (i_14_) & (g122) & (g83)));
	assign g1140 = (((!sk[18]) & (!g123) & (!g335) & (g850)) + ((!sk[18]) & (!g123) & (g335) & (!g850)) + ((!sk[18]) & (!g123) & (g335) & (g850)) + ((!sk[18]) & (g123) & (!g335) & (g850)) + ((!sk[18]) & (g123) & (g335) & (!g850)) + ((!sk[18]) & (g123) & (g335) & (g850)) + ((sk[18]) & (!g123) & (!g335) & (g850)) + ((sk[18]) & (!g123) & (g335) & (!g850)) + ((sk[18]) & (!g123) & (g335) & (g850)));
	assign g1141 = (((!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g445) & (!g105)) + ((!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g445) & (!g105)) + ((!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g445) & (!g105)) + ((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g445) & (!g105)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g445) & (!g105)) + ((i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (g445) & (!g105)) + ((i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g445) & (!g105)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g445) & (!g105)) + ((i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g445) & (!g105)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g445) & (!g105)) + ((i_15_) & (i_12_) & (i_13_) & (i_14_) & (g445) & (!g105)));
	assign g1142 = (((!g1137) & (!sk[20]) & (!g1138) & (g1139) & (!g1140) & (g1141)) + ((!g1137) & (!sk[20]) & (!g1138) & (g1139) & (g1140) & (!g1141)) + ((!g1137) & (!sk[20]) & (!g1138) & (g1139) & (g1140) & (g1141)) + ((!g1137) & (!sk[20]) & (g1138) & (!g1139) & (!g1140) & (!g1141)) + ((!g1137) & (!sk[20]) & (g1138) & (!g1139) & (!g1140) & (g1141)) + ((!g1137) & (!sk[20]) & (g1138) & (!g1139) & (g1140) & (!g1141)) + ((!g1137) & (!sk[20]) & (g1138) & (!g1139) & (g1140) & (g1141)) + ((!g1137) & (!sk[20]) & (g1138) & (g1139) & (!g1140) & (!g1141)) + ((!g1137) & (!sk[20]) & (g1138) & (g1139) & (!g1140) & (g1141)) + ((!g1137) & (!sk[20]) & (g1138) & (g1139) & (g1140) & (!g1141)) + ((!g1137) & (!sk[20]) & (g1138) & (g1139) & (g1140) & (g1141)) + ((!g1137) & (sk[20]) & (!g1138) & (!g1139) & (!g1140) & (!g1141)) + ((g1137) & (!sk[20]) & (!g1138) & (g1139) & (!g1140) & (g1141)) + ((g1137) & (!sk[20]) & (!g1138) & (g1139) & (g1140) & (!g1141)) + ((g1137) & (!sk[20]) & (!g1138) & (g1139) & (g1140) & (g1141)) + ((g1137) & (!sk[20]) & (g1138) & (!g1139) & (!g1140) & (!g1141)) + ((g1137) & (!sk[20]) & (g1138) & (!g1139) & (!g1140) & (g1141)) + ((g1137) & (!sk[20]) & (g1138) & (!g1139) & (g1140) & (!g1141)) + ((g1137) & (!sk[20]) & (g1138) & (!g1139) & (g1140) & (g1141)) + ((g1137) & (!sk[20]) & (g1138) & (g1139) & (!g1140) & (!g1141)) + ((g1137) & (!sk[20]) & (g1138) & (g1139) & (!g1140) & (g1141)) + ((g1137) & (!sk[20]) & (g1138) & (g1139) & (g1140) & (!g1141)) + ((g1137) & (!sk[20]) & (g1138) & (g1139) & (g1140) & (g1141)));
	assign g1143 = (((!g161) & (!sk[21]) & (!g125) & (g185) & (!g182)) + ((!g161) & (!sk[21]) & (!g125) & (g185) & (g182)) + ((!g161) & (!sk[21]) & (g125) & (g185) & (!g182)) + ((!g161) & (!sk[21]) & (g125) & (g185) & (g182)) + ((!g161) & (sk[21]) & (!g125) & (!g185) & (!g182)) + ((!g161) & (sk[21]) & (!g125) & (!g185) & (g182)) + ((!g161) & (sk[21]) & (!g125) & (g185) & (!g182)) + ((!g161) & (sk[21]) & (!g125) & (g185) & (g182)) + ((!g161) & (sk[21]) & (g125) & (!g185) & (!g182)) + ((g161) & (!sk[21]) & (!g125) & (g185) & (!g182)) + ((g161) & (!sk[21]) & (!g125) & (g185) & (g182)) + ((g161) & (!sk[21]) & (g125) & (g185) & (!g182)) + ((g161) & (!sk[21]) & (g125) & (g185) & (g182)) + ((g161) & (sk[21]) & (!g125) & (!g185) & (!g182)) + ((g161) & (sk[21]) & (!g125) & (g185) & (!g182)) + ((g161) & (sk[21]) & (g125) & (!g185) & (!g182)));
	assign g1144 = (((!g164) & (!g154) & (!g340) & (sk[22]) & (!g850)) + ((!g164) & (!g154) & (g340) & (!sk[22]) & (!g850)) + ((!g164) & (!g154) & (g340) & (!sk[22]) & (g850)) + ((!g164) & (!g154) & (g340) & (sk[22]) & (!g850)) + ((!g164) & (g154) & (!g340) & (sk[22]) & (!g850)) + ((!g164) & (g154) & (!g340) & (sk[22]) & (g850)) + ((!g164) & (g154) & (g340) & (!sk[22]) & (!g850)) + ((!g164) & (g154) & (g340) & (!sk[22]) & (g850)) + ((!g164) & (g154) & (g340) & (sk[22]) & (!g850)) + ((!g164) & (g154) & (g340) & (sk[22]) & (g850)) + ((g164) & (!g154) & (g340) & (!sk[22]) & (!g850)) + ((g164) & (!g154) & (g340) & (!sk[22]) & (g850)) + ((g164) & (!g154) & (g340) & (sk[22]) & (!g850)) + ((g164) & (g154) & (g340) & (!sk[22]) & (!g850)) + ((g164) & (g154) & (g340) & (!sk[22]) & (g850)) + ((g164) & (g154) & (g340) & (sk[22]) & (!g850)));
	assign g1145 = (((!g161) & (!g122) & (!g501) & (sk[23]) & (!g543)) + ((!g161) & (!g122) & (!g501) & (sk[23]) & (g543)) + ((!g161) & (!g122) & (g501) & (!sk[23]) & (!g543)) + ((!g161) & (!g122) & (g501) & (!sk[23]) & (g543)) + ((!g161) & (!g122) & (g501) & (sk[23]) & (!g543)) + ((!g161) & (!g122) & (g501) & (sk[23]) & (g543)) + ((!g161) & (g122) & (!g501) & (sk[23]) & (!g543)) + ((!g161) & (g122) & (g501) & (!sk[23]) & (!g543)) + ((!g161) & (g122) & (g501) & (!sk[23]) & (g543)) + ((g161) & (!g122) & (!g501) & (sk[23]) & (!g543)) + ((g161) & (!g122) & (g501) & (!sk[23]) & (!g543)) + ((g161) & (!g122) & (g501) & (!sk[23]) & (g543)) + ((g161) & (!g122) & (g501) & (sk[23]) & (!g543)) + ((g161) & (g122) & (!g501) & (sk[23]) & (!g543)) + ((g161) & (g122) & (g501) & (!sk[23]) & (!g543)) + ((g161) & (g122) & (g501) & (!sk[23]) & (g543)));
	assign g1146 = (((!sk[24]) & (!g362) & (!g1143) & (g1144) & (!g1145)) + ((!sk[24]) & (!g362) & (!g1143) & (g1144) & (g1145)) + ((!sk[24]) & (!g362) & (g1143) & (g1144) & (!g1145)) + ((!sk[24]) & (!g362) & (g1143) & (g1144) & (g1145)) + ((!sk[24]) & (g362) & (!g1143) & (g1144) & (!g1145)) + ((!sk[24]) & (g362) & (!g1143) & (g1144) & (g1145)) + ((!sk[24]) & (g362) & (g1143) & (g1144) & (!g1145)) + ((!sk[24]) & (g362) & (g1143) & (g1144) & (g1145)) + ((sk[24]) & (!g362) & (g1143) & (g1144) & (g1145)));
	assign g1147 = (((!g75) & (!sk[25]) & (!g84) & (g699) & (!g700)) + ((!g75) & (!sk[25]) & (!g84) & (g699) & (g700)) + ((!g75) & (!sk[25]) & (g84) & (g699) & (!g700)) + ((!g75) & (!sk[25]) & (g84) & (g699) & (g700)) + ((!g75) & (sk[25]) & (!g84) & (g699) & (g700)) + ((g75) & (!sk[25]) & (!g84) & (g699) & (!g700)) + ((g75) & (!sk[25]) & (!g84) & (g699) & (g700)) + ((g75) & (!sk[25]) & (g84) & (g699) & (!g700)) + ((g75) & (!sk[25]) & (g84) & (g699) & (g700)) + ((g75) & (sk[25]) & (!g84) & (!g699) & (!g700)) + ((g75) & (sk[25]) & (!g84) & (!g699) & (g700)) + ((g75) & (sk[25]) & (!g84) & (g699) & (!g700)) + ((g75) & (sk[25]) & (!g84) & (g699) & (g700)));
	assign g1148 = (((!g136) & (!g1136) & (!sk[26]) & (g1142) & (!g1146) & (g1147)) + ((!g136) & (!g1136) & (!sk[26]) & (g1142) & (g1146) & (!g1147)) + ((!g136) & (!g1136) & (!sk[26]) & (g1142) & (g1146) & (g1147)) + ((!g136) & (!g1136) & (sk[26]) & (g1142) & (g1146) & (g1147)) + ((!g136) & (g1136) & (!sk[26]) & (!g1142) & (!g1146) & (!g1147)) + ((!g136) & (g1136) & (!sk[26]) & (!g1142) & (!g1146) & (g1147)) + ((!g136) & (g1136) & (!sk[26]) & (!g1142) & (g1146) & (!g1147)) + ((!g136) & (g1136) & (!sk[26]) & (!g1142) & (g1146) & (g1147)) + ((!g136) & (g1136) & (!sk[26]) & (g1142) & (!g1146) & (!g1147)) + ((!g136) & (g1136) & (!sk[26]) & (g1142) & (!g1146) & (g1147)) + ((!g136) & (g1136) & (!sk[26]) & (g1142) & (g1146) & (!g1147)) + ((!g136) & (g1136) & (!sk[26]) & (g1142) & (g1146) & (g1147)) + ((g136) & (!g1136) & (!sk[26]) & (g1142) & (!g1146) & (g1147)) + ((g136) & (!g1136) & (!sk[26]) & (g1142) & (g1146) & (!g1147)) + ((g136) & (!g1136) & (!sk[26]) & (g1142) & (g1146) & (g1147)) + ((g136) & (g1136) & (!sk[26]) & (!g1142) & (!g1146) & (!g1147)) + ((g136) & (g1136) & (!sk[26]) & (!g1142) & (!g1146) & (g1147)) + ((g136) & (g1136) & (!sk[26]) & (!g1142) & (g1146) & (!g1147)) + ((g136) & (g1136) & (!sk[26]) & (!g1142) & (g1146) & (g1147)) + ((g136) & (g1136) & (!sk[26]) & (g1142) & (!g1146) & (!g1147)) + ((g136) & (g1136) & (!sk[26]) & (g1142) & (!g1146) & (g1147)) + ((g136) & (g1136) & (!sk[26]) & (g1142) & (g1146) & (!g1147)) + ((g136) & (g1136) & (!sk[26]) & (g1142) & (g1146) & (g1147)));
	assign g1149 = (((!sk[27]) & (g892) & (!g608)) + ((!sk[27]) & (g892) & (g608)) + ((sk[27]) & (!g892) & (g608)));
	assign g1150 = (((!g75) & (!sk[28]) & (!g105) & (g892) & (!g473) & (g949)) + ((!g75) & (!sk[28]) & (!g105) & (g892) & (g473) & (!g949)) + ((!g75) & (!sk[28]) & (!g105) & (g892) & (g473) & (g949)) + ((!g75) & (!sk[28]) & (g105) & (!g892) & (!g473) & (!g949)) + ((!g75) & (!sk[28]) & (g105) & (!g892) & (!g473) & (g949)) + ((!g75) & (!sk[28]) & (g105) & (!g892) & (g473) & (!g949)) + ((!g75) & (!sk[28]) & (g105) & (!g892) & (g473) & (g949)) + ((!g75) & (!sk[28]) & (g105) & (g892) & (!g473) & (!g949)) + ((!g75) & (!sk[28]) & (g105) & (g892) & (!g473) & (g949)) + ((!g75) & (!sk[28]) & (g105) & (g892) & (g473) & (!g949)) + ((!g75) & (!sk[28]) & (g105) & (g892) & (g473) & (g949)) + ((!g75) & (sk[28]) & (!g105) & (!g892) & (!g473) & (g949)) + ((!g75) & (sk[28]) & (g105) & (!g892) & (!g473) & (g949)) + ((g75) & (!sk[28]) & (!g105) & (g892) & (!g473) & (g949)) + ((g75) & (!sk[28]) & (!g105) & (g892) & (g473) & (!g949)) + ((g75) & (!sk[28]) & (!g105) & (g892) & (g473) & (g949)) + ((g75) & (!sk[28]) & (g105) & (!g892) & (!g473) & (!g949)) + ((g75) & (!sk[28]) & (g105) & (!g892) & (!g473) & (g949)) + ((g75) & (!sk[28]) & (g105) & (!g892) & (g473) & (!g949)) + ((g75) & (!sk[28]) & (g105) & (!g892) & (g473) & (g949)) + ((g75) & (!sk[28]) & (g105) & (g892) & (!g473) & (!g949)) + ((g75) & (!sk[28]) & (g105) & (g892) & (!g473) & (g949)) + ((g75) & (!sk[28]) & (g105) & (g892) & (g473) & (!g949)) + ((g75) & (!sk[28]) & (g105) & (g892) & (g473) & (g949)) + ((g75) & (sk[28]) & (!g105) & (!g892) & (!g473) & (g949)) + ((g75) & (sk[28]) & (!g105) & (!g892) & (g473) & (g949)) + ((g75) & (sk[28]) & (!g105) & (g892) & (!g473) & (g949)) + ((g75) & (sk[28]) & (!g105) & (g892) & (g473) & (g949)) + ((g75) & (sk[28]) & (g105) & (!g892) & (!g473) & (!g949)) + ((g75) & (sk[28]) & (g105) & (!g892) & (!g473) & (g949)) + ((g75) & (sk[28]) & (g105) & (!g892) & (g473) & (!g949)) + ((g75) & (sk[28]) & (g105) & (!g892) & (g473) & (g949)) + ((g75) & (sk[28]) & (g105) & (g892) & (!g473) & (!g949)) + ((g75) & (sk[28]) & (g105) & (g892) & (!g473) & (g949)) + ((g75) & (sk[28]) & (g105) & (g892) & (g473) & (!g949)) + ((g75) & (sk[28]) & (g105) & (g892) & (g473) & (g949)));
	assign g1151 = (((!g161) & (!g1149) & (g503) & (!g1055) & (!sk[29]) & (g1150)) + ((!g161) & (!g1149) & (g503) & (g1055) & (!sk[29]) & (!g1150)) + ((!g161) & (!g1149) & (g503) & (g1055) & (!sk[29]) & (g1150)) + ((!g161) & (!g1149) & (g503) & (g1055) & (sk[29]) & (g1150)) + ((!g161) & (g1149) & (!g503) & (!g1055) & (!sk[29]) & (!g1150)) + ((!g161) & (g1149) & (!g503) & (!g1055) & (!sk[29]) & (g1150)) + ((!g161) & (g1149) & (!g503) & (g1055) & (!sk[29]) & (!g1150)) + ((!g161) & (g1149) & (!g503) & (g1055) & (!sk[29]) & (g1150)) + ((!g161) & (g1149) & (g503) & (!g1055) & (!sk[29]) & (!g1150)) + ((!g161) & (g1149) & (g503) & (!g1055) & (!sk[29]) & (g1150)) + ((!g161) & (g1149) & (g503) & (g1055) & (!sk[29]) & (!g1150)) + ((!g161) & (g1149) & (g503) & (g1055) & (!sk[29]) & (g1150)) + ((!g161) & (g1149) & (g503) & (g1055) & (sk[29]) & (g1150)) + ((g161) & (!g1149) & (g503) & (!g1055) & (!sk[29]) & (g1150)) + ((g161) & (!g1149) & (g503) & (g1055) & (!sk[29]) & (!g1150)) + ((g161) & (!g1149) & (g503) & (g1055) & (!sk[29]) & (g1150)) + ((g161) & (g1149) & (!g503) & (!g1055) & (!sk[29]) & (!g1150)) + ((g161) & (g1149) & (!g503) & (!g1055) & (!sk[29]) & (g1150)) + ((g161) & (g1149) & (!g503) & (g1055) & (!sk[29]) & (!g1150)) + ((g161) & (g1149) & (!g503) & (g1055) & (!sk[29]) & (g1150)) + ((g161) & (g1149) & (g503) & (!g1055) & (!sk[29]) & (!g1150)) + ((g161) & (g1149) & (g503) & (!g1055) & (!sk[29]) & (g1150)) + ((g161) & (g1149) & (g503) & (g1055) & (!sk[29]) & (!g1150)) + ((g161) & (g1149) & (g503) & (g1055) & (!sk[29]) & (g1150)) + ((g161) & (g1149) & (g503) & (g1055) & (sk[29]) & (g1150)));
	assign g1152 = (((!sk[30]) & (!g1131) & (!g1133) & (g1135) & (!g1148) & (g1151)) + ((!sk[30]) & (!g1131) & (!g1133) & (g1135) & (g1148) & (!g1151)) + ((!sk[30]) & (!g1131) & (!g1133) & (g1135) & (g1148) & (g1151)) + ((!sk[30]) & (!g1131) & (g1133) & (!g1135) & (!g1148) & (!g1151)) + ((!sk[30]) & (!g1131) & (g1133) & (!g1135) & (!g1148) & (g1151)) + ((!sk[30]) & (!g1131) & (g1133) & (!g1135) & (g1148) & (!g1151)) + ((!sk[30]) & (!g1131) & (g1133) & (!g1135) & (g1148) & (g1151)) + ((!sk[30]) & (!g1131) & (g1133) & (g1135) & (!g1148) & (!g1151)) + ((!sk[30]) & (!g1131) & (g1133) & (g1135) & (!g1148) & (g1151)) + ((!sk[30]) & (!g1131) & (g1133) & (g1135) & (g1148) & (!g1151)) + ((!sk[30]) & (!g1131) & (g1133) & (g1135) & (g1148) & (g1151)) + ((!sk[30]) & (g1131) & (!g1133) & (g1135) & (!g1148) & (g1151)) + ((!sk[30]) & (g1131) & (!g1133) & (g1135) & (g1148) & (!g1151)) + ((!sk[30]) & (g1131) & (!g1133) & (g1135) & (g1148) & (g1151)) + ((!sk[30]) & (g1131) & (g1133) & (!g1135) & (!g1148) & (!g1151)) + ((!sk[30]) & (g1131) & (g1133) & (!g1135) & (!g1148) & (g1151)) + ((!sk[30]) & (g1131) & (g1133) & (!g1135) & (g1148) & (!g1151)) + ((!sk[30]) & (g1131) & (g1133) & (!g1135) & (g1148) & (g1151)) + ((!sk[30]) & (g1131) & (g1133) & (g1135) & (!g1148) & (!g1151)) + ((!sk[30]) & (g1131) & (g1133) & (g1135) & (!g1148) & (g1151)) + ((!sk[30]) & (g1131) & (g1133) & (g1135) & (g1148) & (!g1151)) + ((!sk[30]) & (g1131) & (g1133) & (g1135) & (g1148) & (g1151)) + ((sk[30]) & (g1131) & (g1133) & (g1135) & (g1148) & (g1151)));
	assign g1153 = (((!sk[31]) & (g1104) & (!g1105)) + ((!sk[31]) & (g1104) & (g1105)) + ((sk[31]) & (!g1104) & (!g1105)));
	assign g1154 = (((!i_12_) & (!i_13_) & (!i_14_) & (!g35) & (g36) & (!g123)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g35) & (!g36) & (!g123)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g35) & (g36) & (!g123)) + ((!i_12_) & (!i_13_) & (i_14_) & (!g35) & (g36) & (!g123)) + ((!i_12_) & (!i_13_) & (i_14_) & (g35) & (!g36) & (!g123)) + ((!i_12_) & (!i_13_) & (i_14_) & (g35) & (g36) & (!g123)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g35) & (g36) & (!g123)) + ((!i_12_) & (i_13_) & (!i_14_) & (g35) & (!g36) & (!g123)) + ((!i_12_) & (i_13_) & (!i_14_) & (g35) & (g36) & (!g123)) + ((!i_12_) & (i_13_) & (i_14_) & (!g35) & (g36) & (!g123)) + ((!i_12_) & (i_13_) & (i_14_) & (g35) & (!g36) & (!g123)) + ((!i_12_) & (i_13_) & (i_14_) & (g35) & (g36) & (!g123)) + ((i_12_) & (!i_13_) & (!i_14_) & (!g35) & (g36) & (!g123)) + ((i_12_) & (!i_13_) & (!i_14_) & (g35) & (!g36) & (!g123)) + ((i_12_) & (!i_13_) & (!i_14_) & (g35) & (g36) & (!g123)) + ((i_12_) & (!i_13_) & (i_14_) & (!g35) & (g36) & (!g123)) + ((i_12_) & (!i_13_) & (i_14_) & (g35) & (!g36) & (!g123)) + ((i_12_) & (!i_13_) & (i_14_) & (g35) & (g36) & (!g123)) + ((i_12_) & (i_13_) & (!i_14_) & (!g35) & (g36) & (!g123)) + ((i_12_) & (i_13_) & (!i_14_) & (g35) & (!g36) & (!g123)) + ((i_12_) & (i_13_) & (!i_14_) & (g35) & (g36) & (!g123)) + ((i_12_) & (i_13_) & (i_14_) & (g35) & (!g36) & (!g123)) + ((i_12_) & (i_13_) & (i_14_) & (g35) & (g36) & (!g123)));
	assign g1155 = (((!sk[33]) & (!g125) & (!g122) & (g186) & (!g513)) + ((!sk[33]) & (!g125) & (!g122) & (g186) & (g513)) + ((!sk[33]) & (!g125) & (g122) & (g186) & (!g513)) + ((!sk[33]) & (!g125) & (g122) & (g186) & (g513)) + ((!sk[33]) & (g125) & (!g122) & (g186) & (!g513)) + ((!sk[33]) & (g125) & (!g122) & (g186) & (g513)) + ((!sk[33]) & (g125) & (g122) & (g186) & (!g513)) + ((!sk[33]) & (g125) & (g122) & (g186) & (g513)) + ((sk[33]) & (!g125) & (!g122) & (!g186) & (!g513)) + ((sk[33]) & (!g125) & (!g122) & (!g186) & (g513)) + ((sk[33]) & (!g125) & (!g122) & (g186) & (!g513)) + ((sk[33]) & (!g125) & (!g122) & (g186) & (g513)) + ((sk[33]) & (!g125) & (g122) & (!g186) & (g513)) + ((sk[33]) & (g125) & (!g122) & (!g186) & (!g513)) + ((sk[33]) & (g125) & (!g122) & (!g186) & (g513)) + ((sk[33]) & (g125) & (g122) & (!g186) & (g513)));
	assign g1156 = (((!i_8_) & (!i_6_) & (!sk[34]) & (i_7_) & (!g924) & (g394)) + ((!i_8_) & (!i_6_) & (!sk[34]) & (i_7_) & (g924) & (!g394)) + ((!i_8_) & (!i_6_) & (!sk[34]) & (i_7_) & (g924) & (g394)) + ((!i_8_) & (i_6_) & (!sk[34]) & (!i_7_) & (!g924) & (!g394)) + ((!i_8_) & (i_6_) & (!sk[34]) & (!i_7_) & (!g924) & (g394)) + ((!i_8_) & (i_6_) & (!sk[34]) & (!i_7_) & (g924) & (!g394)) + ((!i_8_) & (i_6_) & (!sk[34]) & (!i_7_) & (g924) & (g394)) + ((!i_8_) & (i_6_) & (!sk[34]) & (i_7_) & (!g924) & (!g394)) + ((!i_8_) & (i_6_) & (!sk[34]) & (i_7_) & (!g924) & (g394)) + ((!i_8_) & (i_6_) & (!sk[34]) & (i_7_) & (g924) & (!g394)) + ((!i_8_) & (i_6_) & (!sk[34]) & (i_7_) & (g924) & (g394)) + ((i_8_) & (!i_6_) & (!sk[34]) & (i_7_) & (!g924) & (g394)) + ((i_8_) & (!i_6_) & (!sk[34]) & (i_7_) & (g924) & (!g394)) + ((i_8_) & (!i_6_) & (!sk[34]) & (i_7_) & (g924) & (g394)) + ((i_8_) & (!i_6_) & (sk[34]) & (i_7_) & (g924) & (g394)) + ((i_8_) & (i_6_) & (!sk[34]) & (!i_7_) & (!g924) & (!g394)) + ((i_8_) & (i_6_) & (!sk[34]) & (!i_7_) & (!g924) & (g394)) + ((i_8_) & (i_6_) & (!sk[34]) & (!i_7_) & (g924) & (!g394)) + ((i_8_) & (i_6_) & (!sk[34]) & (!i_7_) & (g924) & (g394)) + ((i_8_) & (i_6_) & (!sk[34]) & (i_7_) & (!g924) & (!g394)) + ((i_8_) & (i_6_) & (!sk[34]) & (i_7_) & (!g924) & (g394)) + ((i_8_) & (i_6_) & (!sk[34]) & (i_7_) & (g924) & (!g394)) + ((i_8_) & (i_6_) & (!sk[34]) & (i_7_) & (g924) & (g394)) + ((i_8_) & (i_6_) & (sk[34]) & (!i_7_) & (g924) & (g394)));
	assign g1157 = (((!sk[35]) & (!i_12_) & (!i_13_) & (i_14_) & (!g35) & (g105)) + ((!sk[35]) & (!i_12_) & (!i_13_) & (i_14_) & (g35) & (!g105)) + ((!sk[35]) & (!i_12_) & (!i_13_) & (i_14_) & (g35) & (g105)) + ((!sk[35]) & (!i_12_) & (i_13_) & (!i_14_) & (!g35) & (!g105)) + ((!sk[35]) & (!i_12_) & (i_13_) & (!i_14_) & (!g35) & (g105)) + ((!sk[35]) & (!i_12_) & (i_13_) & (!i_14_) & (g35) & (!g105)) + ((!sk[35]) & (!i_12_) & (i_13_) & (!i_14_) & (g35) & (g105)) + ((!sk[35]) & (!i_12_) & (i_13_) & (i_14_) & (!g35) & (!g105)) + ((!sk[35]) & (!i_12_) & (i_13_) & (i_14_) & (!g35) & (g105)) + ((!sk[35]) & (!i_12_) & (i_13_) & (i_14_) & (g35) & (!g105)) + ((!sk[35]) & (!i_12_) & (i_13_) & (i_14_) & (g35) & (g105)) + ((!sk[35]) & (i_12_) & (!i_13_) & (i_14_) & (!g35) & (g105)) + ((!sk[35]) & (i_12_) & (!i_13_) & (i_14_) & (g35) & (!g105)) + ((!sk[35]) & (i_12_) & (!i_13_) & (i_14_) & (g35) & (g105)) + ((!sk[35]) & (i_12_) & (i_13_) & (!i_14_) & (!g35) & (!g105)) + ((!sk[35]) & (i_12_) & (i_13_) & (!i_14_) & (!g35) & (g105)) + ((!sk[35]) & (i_12_) & (i_13_) & (!i_14_) & (g35) & (!g105)) + ((!sk[35]) & (i_12_) & (i_13_) & (!i_14_) & (g35) & (g105)) + ((!sk[35]) & (i_12_) & (i_13_) & (i_14_) & (!g35) & (!g105)) + ((!sk[35]) & (i_12_) & (i_13_) & (i_14_) & (!g35) & (g105)) + ((!sk[35]) & (i_12_) & (i_13_) & (i_14_) & (g35) & (!g105)) + ((!sk[35]) & (i_12_) & (i_13_) & (i_14_) & (g35) & (g105)) + ((sk[35]) & (!i_12_) & (!i_13_) & (i_14_) & (g35) & (!g105)) + ((sk[35]) & (!i_12_) & (i_13_) & (!i_14_) & (g35) & (!g105)) + ((sk[35]) & (i_12_) & (!i_13_) & (!i_14_) & (g35) & (!g105)) + ((sk[35]) & (i_12_) & (i_13_) & (!i_14_) & (g35) & (!g105)) + ((sk[35]) & (i_12_) & (i_13_) & (i_14_) & (g35) & (!g105)));
	assign g1158 = (((!g164) & (!g483) & (!g641) & (!g1156) & (sk[36]) & (!g1157)) + ((!g164) & (!g483) & (g641) & (!g1156) & (!sk[36]) & (g1157)) + ((!g164) & (!g483) & (g641) & (!g1156) & (sk[36]) & (!g1157)) + ((!g164) & (!g483) & (g641) & (g1156) & (!sk[36]) & (!g1157)) + ((!g164) & (!g483) & (g641) & (g1156) & (!sk[36]) & (g1157)) + ((!g164) & (g483) & (!g641) & (!g1156) & (!sk[36]) & (!g1157)) + ((!g164) & (g483) & (!g641) & (!g1156) & (!sk[36]) & (g1157)) + ((!g164) & (g483) & (!g641) & (!g1156) & (sk[36]) & (!g1157)) + ((!g164) & (g483) & (!g641) & (g1156) & (!sk[36]) & (!g1157)) + ((!g164) & (g483) & (!g641) & (g1156) & (!sk[36]) & (g1157)) + ((!g164) & (g483) & (g641) & (!g1156) & (!sk[36]) & (!g1157)) + ((!g164) & (g483) & (g641) & (!g1156) & (!sk[36]) & (g1157)) + ((!g164) & (g483) & (g641) & (!g1156) & (sk[36]) & (!g1157)) + ((!g164) & (g483) & (g641) & (g1156) & (!sk[36]) & (!g1157)) + ((!g164) & (g483) & (g641) & (g1156) & (!sk[36]) & (g1157)) + ((g164) & (!g483) & (!g641) & (!g1156) & (sk[36]) & (!g1157)) + ((g164) & (!g483) & (g641) & (!g1156) & (!sk[36]) & (g1157)) + ((g164) & (!g483) & (g641) & (g1156) & (!sk[36]) & (!g1157)) + ((g164) & (!g483) & (g641) & (g1156) & (!sk[36]) & (g1157)) + ((g164) & (g483) & (!g641) & (!g1156) & (!sk[36]) & (!g1157)) + ((g164) & (g483) & (!g641) & (!g1156) & (!sk[36]) & (g1157)) + ((g164) & (g483) & (!g641) & (g1156) & (!sk[36]) & (!g1157)) + ((g164) & (g483) & (!g641) & (g1156) & (!sk[36]) & (g1157)) + ((g164) & (g483) & (g641) & (!g1156) & (!sk[36]) & (!g1157)) + ((g164) & (g483) & (g641) & (!g1156) & (!sk[36]) & (g1157)) + ((g164) & (g483) & (g641) & (g1156) & (!sk[36]) & (!g1157)) + ((g164) & (g483) & (g641) & (g1156) & (!sk[36]) & (g1157)));
	assign g1159 = (((!g161) & (!g186) & (!g192) & (!g878) & (g1155) & (g1158)) + ((!g161) & (!g186) & (g192) & (!g878) & (g1155) & (g1158)) + ((!g161) & (g186) & (!g192) & (!g878) & (g1155) & (g1158)) + ((!g161) & (g186) & (g192) & (!g878) & (g1155) & (g1158)) + ((g161) & (!g186) & (!g192) & (!g878) & (g1155) & (g1158)));
	assign g1160 = (((!i_12_) & (!i_13_) & (!i_14_) & (!g35) & (g36) & (!g105)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g35) & (g36) & (!g105)) + ((!i_12_) & (!i_13_) & (i_14_) & (!g35) & (g36) & (!g105)) + ((!i_12_) & (!i_13_) & (i_14_) & (g35) & (g36) & (!g105)) + ((!i_12_) & (i_13_) & (i_14_) & (!g35) & (g36) & (!g105)) + ((!i_12_) & (i_13_) & (i_14_) & (g35) & (!g36) & (!g105)) + ((!i_12_) & (i_13_) & (i_14_) & (g35) & (g36) & (!g105)) + ((i_12_) & (!i_13_) & (!i_14_) & (!g35) & (g36) & (!g105)) + ((i_12_) & (!i_13_) & (!i_14_) & (g35) & (g36) & (!g105)) + ((i_12_) & (!i_13_) & (i_14_) & (!g35) & (g36) & (!g105)) + ((i_12_) & (!i_13_) & (i_14_) & (g35) & (g36) & (!g105)) + ((i_12_) & (i_13_) & (!i_14_) & (!g35) & (g36) & (!g105)) + ((i_12_) & (i_13_) & (!i_14_) & (g35) & (g36) & (!g105)));
	assign g1161 = (((!g161) & (!sk[39]) & (!g122) & (g337) & (!g851) & (g1160)) + ((!g161) & (!sk[39]) & (!g122) & (g337) & (g851) & (!g1160)) + ((!g161) & (!sk[39]) & (!g122) & (g337) & (g851) & (g1160)) + ((!g161) & (!sk[39]) & (g122) & (!g337) & (!g851) & (!g1160)) + ((!g161) & (!sk[39]) & (g122) & (!g337) & (!g851) & (g1160)) + ((!g161) & (!sk[39]) & (g122) & (!g337) & (g851) & (!g1160)) + ((!g161) & (!sk[39]) & (g122) & (!g337) & (g851) & (g1160)) + ((!g161) & (!sk[39]) & (g122) & (g337) & (!g851) & (!g1160)) + ((!g161) & (!sk[39]) & (g122) & (g337) & (!g851) & (g1160)) + ((!g161) & (!sk[39]) & (g122) & (g337) & (g851) & (!g1160)) + ((!g161) & (!sk[39]) & (g122) & (g337) & (g851) & (g1160)) + ((!g161) & (sk[39]) & (!g122) & (!g337) & (!g851) & (!g1160)) + ((!g161) & (sk[39]) & (!g122) & (!g337) & (g851) & (!g1160)) + ((!g161) & (sk[39]) & (!g122) & (g337) & (!g851) & (!g1160)) + ((!g161) & (sk[39]) & (!g122) & (g337) & (g851) & (!g1160)) + ((!g161) & (sk[39]) & (g122) & (!g337) & (g851) & (!g1160)) + ((!g161) & (sk[39]) & (g122) & (g337) & (g851) & (!g1160)) + ((g161) & (!sk[39]) & (!g122) & (g337) & (!g851) & (g1160)) + ((g161) & (!sk[39]) & (!g122) & (g337) & (g851) & (!g1160)) + ((g161) & (!sk[39]) & (!g122) & (g337) & (g851) & (g1160)) + ((g161) & (!sk[39]) & (g122) & (!g337) & (!g851) & (!g1160)) + ((g161) & (!sk[39]) & (g122) & (!g337) & (!g851) & (g1160)) + ((g161) & (!sk[39]) & (g122) & (!g337) & (g851) & (!g1160)) + ((g161) & (!sk[39]) & (g122) & (!g337) & (g851) & (g1160)) + ((g161) & (!sk[39]) & (g122) & (g337) & (!g851) & (!g1160)) + ((g161) & (!sk[39]) & (g122) & (g337) & (!g851) & (g1160)) + ((g161) & (!sk[39]) & (g122) & (g337) & (g851) & (!g1160)) + ((g161) & (!sk[39]) & (g122) & (g337) & (g851) & (g1160)) + ((g161) & (sk[39]) & (!g122) & (!g337) & (!g851) & (!g1160)) + ((g161) & (sk[39]) & (!g122) & (!g337) & (g851) & (!g1160)) + ((g161) & (sk[39]) & (g122) & (!g337) & (g851) & (!g1160)));
	assign g1162 = (((!g75) & (!g192) & (!sk[40]) & (g513) & (!g514) & (g1161)) + ((!g75) & (!g192) & (!sk[40]) & (g513) & (g514) & (!g1161)) + ((!g75) & (!g192) & (!sk[40]) & (g513) & (g514) & (g1161)) + ((!g75) & (!g192) & (sk[40]) & (g513) & (!g514) & (g1161)) + ((!g75) & (g192) & (!sk[40]) & (!g513) & (!g514) & (!g1161)) + ((!g75) & (g192) & (!sk[40]) & (!g513) & (!g514) & (g1161)) + ((!g75) & (g192) & (!sk[40]) & (!g513) & (g514) & (!g1161)) + ((!g75) & (g192) & (!sk[40]) & (!g513) & (g514) & (g1161)) + ((!g75) & (g192) & (!sk[40]) & (g513) & (!g514) & (!g1161)) + ((!g75) & (g192) & (!sk[40]) & (g513) & (!g514) & (g1161)) + ((!g75) & (g192) & (!sk[40]) & (g513) & (g514) & (!g1161)) + ((!g75) & (g192) & (!sk[40]) & (g513) & (g514) & (g1161)) + ((g75) & (!g192) & (!sk[40]) & (g513) & (!g514) & (g1161)) + ((g75) & (!g192) & (!sk[40]) & (g513) & (g514) & (!g1161)) + ((g75) & (!g192) & (!sk[40]) & (g513) & (g514) & (g1161)) + ((g75) & (!g192) & (sk[40]) & (!g513) & (!g514) & (g1161)) + ((g75) & (!g192) & (sk[40]) & (!g513) & (g514) & (g1161)) + ((g75) & (!g192) & (sk[40]) & (g513) & (!g514) & (g1161)) + ((g75) & (!g192) & (sk[40]) & (g513) & (g514) & (g1161)) + ((g75) & (g192) & (!sk[40]) & (!g513) & (!g514) & (!g1161)) + ((g75) & (g192) & (!sk[40]) & (!g513) & (!g514) & (g1161)) + ((g75) & (g192) & (!sk[40]) & (!g513) & (g514) & (!g1161)) + ((g75) & (g192) & (!sk[40]) & (!g513) & (g514) & (g1161)) + ((g75) & (g192) & (!sk[40]) & (g513) & (!g514) & (!g1161)) + ((g75) & (g192) & (!sk[40]) & (g513) & (!g514) & (g1161)) + ((g75) & (g192) & (!sk[40]) & (g513) & (g514) & (!g1161)) + ((g75) & (g192) & (!sk[40]) & (g513) & (g514) & (g1161)) + ((g75) & (g192) & (sk[40]) & (!g513) & (!g514) & (g1161)) + ((g75) & (g192) & (sk[40]) & (!g513) & (g514) & (g1161)) + ((g75) & (g192) & (sk[40]) & (g513) & (!g514) & (g1161)) + ((g75) & (g192) & (sk[40]) & (g513) & (g514) & (g1161)));
	assign g1163 = (((!sk[41]) & (!g634) & (!g37) & (g75) & (!g759) & (g710)) + ((!sk[41]) & (!g634) & (!g37) & (g75) & (g759) & (!g710)) + ((!sk[41]) & (!g634) & (!g37) & (g75) & (g759) & (g710)) + ((!sk[41]) & (!g634) & (g37) & (!g75) & (!g759) & (!g710)) + ((!sk[41]) & (!g634) & (g37) & (!g75) & (!g759) & (g710)) + ((!sk[41]) & (!g634) & (g37) & (!g75) & (g759) & (!g710)) + ((!sk[41]) & (!g634) & (g37) & (!g75) & (g759) & (g710)) + ((!sk[41]) & (!g634) & (g37) & (g75) & (!g759) & (!g710)) + ((!sk[41]) & (!g634) & (g37) & (g75) & (!g759) & (g710)) + ((!sk[41]) & (!g634) & (g37) & (g75) & (g759) & (!g710)) + ((!sk[41]) & (!g634) & (g37) & (g75) & (g759) & (g710)) + ((!sk[41]) & (g634) & (!g37) & (g75) & (!g759) & (g710)) + ((!sk[41]) & (g634) & (!g37) & (g75) & (g759) & (!g710)) + ((!sk[41]) & (g634) & (!g37) & (g75) & (g759) & (g710)) + ((!sk[41]) & (g634) & (g37) & (!g75) & (!g759) & (!g710)) + ((!sk[41]) & (g634) & (g37) & (!g75) & (!g759) & (g710)) + ((!sk[41]) & (g634) & (g37) & (!g75) & (g759) & (!g710)) + ((!sk[41]) & (g634) & (g37) & (!g75) & (g759) & (g710)) + ((!sk[41]) & (g634) & (g37) & (g75) & (!g759) & (!g710)) + ((!sk[41]) & (g634) & (g37) & (g75) & (!g759) & (g710)) + ((!sk[41]) & (g634) & (g37) & (g75) & (g759) & (!g710)) + ((!sk[41]) & (g634) & (g37) & (g75) & (g759) & (g710)) + ((sk[41]) & (!g634) & (!g37) & (g75) & (g759) & (!g710)) + ((sk[41]) & (!g634) & (g37) & (g75) & (g759) & (!g710)) + ((sk[41]) & (g634) & (!g37) & (g75) & (g759) & (!g710)) + ((sk[41]) & (g634) & (g37) & (!g75) & (g759) & (!g710)) + ((sk[41]) & (g634) & (g37) & (g75) & (g759) & (!g710)));
	assign g1164 = (((!g164) & (!sk[42]) & (!g339) & (g849) & (!g851)) + ((!g164) & (!sk[42]) & (!g339) & (g849) & (g851)) + ((!g164) & (!sk[42]) & (g339) & (g849) & (!g851)) + ((!g164) & (!sk[42]) & (g339) & (g849) & (g851)) + ((g164) & (!sk[42]) & (!g339) & (g849) & (!g851)) + ((g164) & (!sk[42]) & (!g339) & (g849) & (g851)) + ((g164) & (!sk[42]) & (g339) & (g849) & (!g851)) + ((g164) & (!sk[42]) & (g339) & (g849) & (g851)) + ((g164) & (sk[42]) & (!g339) & (!g849) & (!g851)) + ((g164) & (sk[42]) & (!g339) & (g849) & (!g851)) + ((g164) & (sk[42]) & (!g339) & (g849) & (g851)) + ((g164) & (sk[42]) & (g339) & (!g849) & (!g851)) + ((g164) & (sk[42]) & (g339) & (!g849) & (g851)) + ((g164) & (sk[42]) & (g339) & (g849) & (!g851)) + ((g164) & (sk[42]) & (g339) & (g849) & (g851)));
	assign g1165 = (((!sk[43]) & (!i_8_) & (!g35) & (g73) & (!g68) & (g460)) + ((!sk[43]) & (!i_8_) & (!g35) & (g73) & (g68) & (!g460)) + ((!sk[43]) & (!i_8_) & (!g35) & (g73) & (g68) & (g460)) + ((!sk[43]) & (!i_8_) & (g35) & (!g73) & (!g68) & (!g460)) + ((!sk[43]) & (!i_8_) & (g35) & (!g73) & (!g68) & (g460)) + ((!sk[43]) & (!i_8_) & (g35) & (!g73) & (g68) & (!g460)) + ((!sk[43]) & (!i_8_) & (g35) & (!g73) & (g68) & (g460)) + ((!sk[43]) & (!i_8_) & (g35) & (g73) & (!g68) & (!g460)) + ((!sk[43]) & (!i_8_) & (g35) & (g73) & (!g68) & (g460)) + ((!sk[43]) & (!i_8_) & (g35) & (g73) & (g68) & (!g460)) + ((!sk[43]) & (!i_8_) & (g35) & (g73) & (g68) & (g460)) + ((!sk[43]) & (i_8_) & (!g35) & (g73) & (!g68) & (g460)) + ((!sk[43]) & (i_8_) & (!g35) & (g73) & (g68) & (!g460)) + ((!sk[43]) & (i_8_) & (!g35) & (g73) & (g68) & (g460)) + ((!sk[43]) & (i_8_) & (g35) & (!g73) & (!g68) & (!g460)) + ((!sk[43]) & (i_8_) & (g35) & (!g73) & (!g68) & (g460)) + ((!sk[43]) & (i_8_) & (g35) & (!g73) & (g68) & (!g460)) + ((!sk[43]) & (i_8_) & (g35) & (!g73) & (g68) & (g460)) + ((!sk[43]) & (i_8_) & (g35) & (g73) & (!g68) & (!g460)) + ((!sk[43]) & (i_8_) & (g35) & (g73) & (!g68) & (g460)) + ((!sk[43]) & (i_8_) & (g35) & (g73) & (g68) & (!g460)) + ((!sk[43]) & (i_8_) & (g35) & (g73) & (g68) & (g460)) + ((sk[43]) & (i_8_) & (g35) & (g73) & (!g68) & (!g460)) + ((sk[43]) & (i_8_) & (g35) & (g73) & (!g68) & (g460)) + ((sk[43]) & (i_8_) & (g35) & (g73) & (g68) & (!g460)));
	assign g1166 = (((!g30) & (!sk[44]) & (!g49) & (g118) & (!g605) & (g514)) + ((!g30) & (!sk[44]) & (!g49) & (g118) & (g605) & (!g514)) + ((!g30) & (!sk[44]) & (!g49) & (g118) & (g605) & (g514)) + ((!g30) & (!sk[44]) & (g49) & (!g118) & (!g605) & (!g514)) + ((!g30) & (!sk[44]) & (g49) & (!g118) & (!g605) & (g514)) + ((!g30) & (!sk[44]) & (g49) & (!g118) & (g605) & (!g514)) + ((!g30) & (!sk[44]) & (g49) & (!g118) & (g605) & (g514)) + ((!g30) & (!sk[44]) & (g49) & (g118) & (!g605) & (!g514)) + ((!g30) & (!sk[44]) & (g49) & (g118) & (!g605) & (g514)) + ((!g30) & (!sk[44]) & (g49) & (g118) & (g605) & (!g514)) + ((!g30) & (!sk[44]) & (g49) & (g118) & (g605) & (g514)) + ((!g30) & (sk[44]) & (!g49) & (g118) & (g605) & (g514)) + ((!g30) & (sk[44]) & (g49) & (g118) & (!g605) & (g514)) + ((!g30) & (sk[44]) & (g49) & (g118) & (g605) & (g514)) + ((g30) & (!sk[44]) & (!g49) & (g118) & (!g605) & (g514)) + ((g30) & (!sk[44]) & (!g49) & (g118) & (g605) & (!g514)) + ((g30) & (!sk[44]) & (!g49) & (g118) & (g605) & (g514)) + ((g30) & (!sk[44]) & (g49) & (!g118) & (!g605) & (!g514)) + ((g30) & (!sk[44]) & (g49) & (!g118) & (!g605) & (g514)) + ((g30) & (!sk[44]) & (g49) & (!g118) & (g605) & (!g514)) + ((g30) & (!sk[44]) & (g49) & (!g118) & (g605) & (g514)) + ((g30) & (!sk[44]) & (g49) & (g118) & (!g605) & (!g514)) + ((g30) & (!sk[44]) & (g49) & (g118) & (!g605) & (g514)) + ((g30) & (!sk[44]) & (g49) & (g118) & (g605) & (!g514)) + ((g30) & (!sk[44]) & (g49) & (g118) & (g605) & (g514)) + ((g30) & (sk[44]) & (!g49) & (g118) & (g605) & (!g514)) + ((g30) & (sk[44]) & (!g49) & (g118) & (g605) & (g514)) + ((g30) & (sk[44]) & (g49) & (g118) & (!g605) & (!g514)) + ((g30) & (sk[44]) & (g49) & (g118) & (!g605) & (g514)) + ((g30) & (sk[44]) & (g49) & (g118) & (g605) & (!g514)) + ((g30) & (sk[44]) & (g49) & (g118) & (g605) & (g514)));
	assign g1167 = (((i_8_) & (!i_7_) & (!i_12_) & (!i_13_) & (i_14_) & (g36)) + ((i_8_) & (!i_7_) & (i_12_) & (i_13_) & (i_14_) & (g36)));
	assign g1168 = (((!i_8_) & (!g73) & (!g90) & (!g186) & (g1166) & (g1167)) + ((!i_8_) & (!g73) & (!g90) & (g186) & (g1166) & (g1167)) + ((!i_8_) & (!g73) & (g90) & (!g186) & (g1166) & (g1167)) + ((!i_8_) & (!g73) & (g90) & (g186) & (g1166) & (g1167)) + ((!i_8_) & (g73) & (!g90) & (!g186) & (g1166) & (g1167)) + ((!i_8_) & (g73) & (!g90) & (g186) & (g1166) & (g1167)) + ((!i_8_) & (g73) & (g90) & (!g186) & (g1166) & (g1167)) + ((!i_8_) & (g73) & (g90) & (g186) & (g1166) & (g1167)) + ((i_8_) & (!g73) & (!g90) & (!g186) & (g1166) & (g1167)) + ((i_8_) & (!g73) & (!g90) & (g186) & (g1166) & (g1167)) + ((i_8_) & (!g73) & (g90) & (!g186) & (g1166) & (g1167)) + ((i_8_) & (!g73) & (g90) & (g186) & (g1166) & (g1167)) + ((i_8_) & (g73) & (!g90) & (!g186) & (g1166) & (g1167)) + ((i_8_) & (g73) & (!g90) & (g186) & (!g1166) & (!g1167)) + ((i_8_) & (g73) & (!g90) & (g186) & (!g1166) & (g1167)) + ((i_8_) & (g73) & (!g90) & (g186) & (g1166) & (!g1167)) + ((i_8_) & (g73) & (!g90) & (g186) & (g1166) & (g1167)) + ((i_8_) & (g73) & (g90) & (!g186) & (!g1166) & (!g1167)) + ((i_8_) & (g73) & (g90) & (!g186) & (!g1166) & (g1167)) + ((i_8_) & (g73) & (g90) & (!g186) & (g1166) & (!g1167)) + ((i_8_) & (g73) & (g90) & (!g186) & (g1166) & (g1167)) + ((i_8_) & (g73) & (g90) & (g186) & (!g1166) & (!g1167)) + ((i_8_) & (g73) & (g90) & (g186) & (!g1166) & (g1167)) + ((i_8_) & (g73) & (g90) & (g186) & (g1166) & (!g1167)) + ((i_8_) & (g73) & (g90) & (g186) & (g1166) & (g1167)));
	assign g1169 = (((!g634) & (!g125) & (!g281) & (!g1165) & (sk[47]) & (!g1168)) + ((!g634) & (!g125) & (g281) & (!g1165) & (!sk[47]) & (g1168)) + ((!g634) & (!g125) & (g281) & (!g1165) & (sk[47]) & (!g1168)) + ((!g634) & (!g125) & (g281) & (g1165) & (!sk[47]) & (!g1168)) + ((!g634) & (!g125) & (g281) & (g1165) & (!sk[47]) & (g1168)) + ((!g634) & (g125) & (!g281) & (!g1165) & (!sk[47]) & (!g1168)) + ((!g634) & (g125) & (!g281) & (!g1165) & (!sk[47]) & (g1168)) + ((!g634) & (g125) & (!g281) & (g1165) & (!sk[47]) & (!g1168)) + ((!g634) & (g125) & (!g281) & (g1165) & (!sk[47]) & (g1168)) + ((!g634) & (g125) & (g281) & (!g1165) & (!sk[47]) & (!g1168)) + ((!g634) & (g125) & (g281) & (!g1165) & (!sk[47]) & (g1168)) + ((!g634) & (g125) & (g281) & (g1165) & (!sk[47]) & (!g1168)) + ((!g634) & (g125) & (g281) & (g1165) & (!sk[47]) & (g1168)) + ((g634) & (!g125) & (!g281) & (!g1165) & (sk[47]) & (!g1168)) + ((g634) & (!g125) & (g281) & (!g1165) & (!sk[47]) & (g1168)) + ((g634) & (!g125) & (g281) & (!g1165) & (sk[47]) & (!g1168)) + ((g634) & (!g125) & (g281) & (g1165) & (!sk[47]) & (!g1168)) + ((g634) & (!g125) & (g281) & (g1165) & (!sk[47]) & (g1168)) + ((g634) & (g125) & (!g281) & (!g1165) & (!sk[47]) & (!g1168)) + ((g634) & (g125) & (!g281) & (!g1165) & (!sk[47]) & (g1168)) + ((g634) & (g125) & (!g281) & (!g1165) & (sk[47]) & (!g1168)) + ((g634) & (g125) & (!g281) & (g1165) & (!sk[47]) & (!g1168)) + ((g634) & (g125) & (!g281) & (g1165) & (!sk[47]) & (g1168)) + ((g634) & (g125) & (g281) & (!g1165) & (!sk[47]) & (!g1168)) + ((g634) & (g125) & (g281) & (!g1165) & (!sk[47]) & (g1168)) + ((g634) & (g125) & (g281) & (g1165) & (!sk[47]) & (!g1168)) + ((g634) & (g125) & (g281) & (g1165) & (!sk[47]) & (g1168)));
	assign g1170 = (((!g125) & (!g164) & (!g122) & (!g105) & (sk[48]) & (!g948)) + ((!g125) & (!g164) & (g122) & (!g105) & (!sk[48]) & (g948)) + ((!g125) & (!g164) & (g122) & (!g105) & (sk[48]) & (!g948)) + ((!g125) & (!g164) & (g122) & (g105) & (!sk[48]) & (!g948)) + ((!g125) & (!g164) & (g122) & (g105) & (!sk[48]) & (g948)) + ((!g125) & (!g164) & (g122) & (g105) & (sk[48]) & (!g948)) + ((!g125) & (g164) & (!g122) & (!g105) & (!sk[48]) & (!g948)) + ((!g125) & (g164) & (!g122) & (!g105) & (!sk[48]) & (g948)) + ((!g125) & (g164) & (!g122) & (!g105) & (sk[48]) & (!g948)) + ((!g125) & (g164) & (!g122) & (g105) & (!sk[48]) & (!g948)) + ((!g125) & (g164) & (!g122) & (g105) & (!sk[48]) & (g948)) + ((!g125) & (g164) & (!g122) & (g105) & (sk[48]) & (!g948)) + ((!g125) & (g164) & (g122) & (!g105) & (!sk[48]) & (!g948)) + ((!g125) & (g164) & (g122) & (!g105) & (!sk[48]) & (g948)) + ((!g125) & (g164) & (g122) & (!g105) & (sk[48]) & (!g948)) + ((!g125) & (g164) & (g122) & (g105) & (!sk[48]) & (!g948)) + ((!g125) & (g164) & (g122) & (g105) & (!sk[48]) & (g948)) + ((!g125) & (g164) & (g122) & (g105) & (sk[48]) & (!g948)) + ((g125) & (!g164) & (!g122) & (!g105) & (sk[48]) & (!g948)) + ((g125) & (!g164) & (!g122) & (g105) & (sk[48]) & (!g948)) + ((g125) & (!g164) & (g122) & (!g105) & (!sk[48]) & (g948)) + ((g125) & (!g164) & (g122) & (!g105) & (sk[48]) & (!g948)) + ((g125) & (!g164) & (g122) & (g105) & (!sk[48]) & (!g948)) + ((g125) & (!g164) & (g122) & (g105) & (!sk[48]) & (g948)) + ((g125) & (!g164) & (g122) & (g105) & (sk[48]) & (!g948)) + ((g125) & (g164) & (!g122) & (!g105) & (!sk[48]) & (!g948)) + ((g125) & (g164) & (!g122) & (!g105) & (!sk[48]) & (g948)) + ((g125) & (g164) & (!g122) & (!g105) & (sk[48]) & (!g948)) + ((g125) & (g164) & (!g122) & (g105) & (!sk[48]) & (!g948)) + ((g125) & (g164) & (!g122) & (g105) & (!sk[48]) & (g948)) + ((g125) & (g164) & (!g122) & (g105) & (sk[48]) & (!g948)) + ((g125) & (g164) & (g122) & (!g105) & (!sk[48]) & (!g948)) + ((g125) & (g164) & (g122) & (!g105) & (!sk[48]) & (g948)) + ((g125) & (g164) & (g122) & (!g105) & (sk[48]) & (!g948)) + ((g125) & (g164) & (g122) & (g105) & (!sk[48]) & (!g948)) + ((g125) & (g164) & (g122) & (g105) & (!sk[48]) & (g948)) + ((g125) & (g164) & (g122) & (g105) & (sk[48]) & (!g948)));
	assign g1171 = (((!sk[49]) & (!g1455) & (!g1048) & (g1164) & (!g1169) & (g1170)) + ((!sk[49]) & (!g1455) & (!g1048) & (g1164) & (g1169) & (!g1170)) + ((!sk[49]) & (!g1455) & (!g1048) & (g1164) & (g1169) & (g1170)) + ((!sk[49]) & (!g1455) & (g1048) & (!g1164) & (!g1169) & (!g1170)) + ((!sk[49]) & (!g1455) & (g1048) & (!g1164) & (!g1169) & (g1170)) + ((!sk[49]) & (!g1455) & (g1048) & (!g1164) & (g1169) & (!g1170)) + ((!sk[49]) & (!g1455) & (g1048) & (!g1164) & (g1169) & (g1170)) + ((!sk[49]) & (!g1455) & (g1048) & (g1164) & (!g1169) & (!g1170)) + ((!sk[49]) & (!g1455) & (g1048) & (g1164) & (!g1169) & (g1170)) + ((!sk[49]) & (!g1455) & (g1048) & (g1164) & (g1169) & (!g1170)) + ((!sk[49]) & (!g1455) & (g1048) & (g1164) & (g1169) & (g1170)) + ((!sk[49]) & (g1455) & (!g1048) & (g1164) & (!g1169) & (g1170)) + ((!sk[49]) & (g1455) & (!g1048) & (g1164) & (g1169) & (!g1170)) + ((!sk[49]) & (g1455) & (!g1048) & (g1164) & (g1169) & (g1170)) + ((!sk[49]) & (g1455) & (g1048) & (!g1164) & (!g1169) & (!g1170)) + ((!sk[49]) & (g1455) & (g1048) & (!g1164) & (!g1169) & (g1170)) + ((!sk[49]) & (g1455) & (g1048) & (!g1164) & (g1169) & (!g1170)) + ((!sk[49]) & (g1455) & (g1048) & (!g1164) & (g1169) & (g1170)) + ((!sk[49]) & (g1455) & (g1048) & (g1164) & (!g1169) & (!g1170)) + ((!sk[49]) & (g1455) & (g1048) & (g1164) & (!g1169) & (g1170)) + ((!sk[49]) & (g1455) & (g1048) & (g1164) & (g1169) & (!g1170)) + ((!sk[49]) & (g1455) & (g1048) & (g1164) & (g1169) & (g1170)) + ((sk[49]) & (!g1455) & (!g1048) & (!g1164) & (g1169) & (!g1170)));
	assign g1172 = (((g1153) & (!g1154) & (g1159) & (g1162) & (g1163) & (g1171)));
	assign g1173 = (((!g125) & (!sk[51]) & (!g122) & (g648) & (!g847)) + ((!g125) & (!sk[51]) & (!g122) & (g648) & (g847)) + ((!g125) & (!sk[51]) & (g122) & (g648) & (!g847)) + ((!g125) & (!sk[51]) & (g122) & (g648) & (g847)) + ((!g125) & (sk[51]) & (!g122) & (!g648) & (!g847)) + ((!g125) & (sk[51]) & (!g122) & (!g648) & (g847)) + ((!g125) & (sk[51]) & (!g122) & (g648) & (!g847)) + ((!g125) & (sk[51]) & (!g122) & (g648) & (g847)) + ((!g125) & (sk[51]) & (g122) & (!g648) & (g847)) + ((g125) & (!sk[51]) & (!g122) & (g648) & (!g847)) + ((g125) & (!sk[51]) & (!g122) & (g648) & (g847)) + ((g125) & (!sk[51]) & (g122) & (g648) & (!g847)) + ((g125) & (!sk[51]) & (g122) & (g648) & (g847)) + ((g125) & (sk[51]) & (!g122) & (!g648) & (!g847)) + ((g125) & (sk[51]) & (!g122) & (!g648) & (g847)) + ((g125) & (sk[51]) & (g122) & (!g648) & (g847)));
	assign g1174 = (((!i_8_) & (!i_6_) & (i_7_) & (!sk[52]) & (!g429) & (g394)) + ((!i_8_) & (!i_6_) & (i_7_) & (!sk[52]) & (g429) & (!g394)) + ((!i_8_) & (!i_6_) & (i_7_) & (!sk[52]) & (g429) & (g394)) + ((!i_8_) & (i_6_) & (!i_7_) & (!sk[52]) & (!g429) & (!g394)) + ((!i_8_) & (i_6_) & (!i_7_) & (!sk[52]) & (!g429) & (g394)) + ((!i_8_) & (i_6_) & (!i_7_) & (!sk[52]) & (g429) & (!g394)) + ((!i_8_) & (i_6_) & (!i_7_) & (!sk[52]) & (g429) & (g394)) + ((!i_8_) & (i_6_) & (i_7_) & (!sk[52]) & (!g429) & (!g394)) + ((!i_8_) & (i_6_) & (i_7_) & (!sk[52]) & (!g429) & (g394)) + ((!i_8_) & (i_6_) & (i_7_) & (!sk[52]) & (g429) & (!g394)) + ((!i_8_) & (i_6_) & (i_7_) & (!sk[52]) & (g429) & (g394)) + ((i_8_) & (!i_6_) & (i_7_) & (!sk[52]) & (!g429) & (g394)) + ((i_8_) & (!i_6_) & (i_7_) & (!sk[52]) & (g429) & (!g394)) + ((i_8_) & (!i_6_) & (i_7_) & (!sk[52]) & (g429) & (g394)) + ((i_8_) & (!i_6_) & (i_7_) & (sk[52]) & (g429) & (g394)) + ((i_8_) & (i_6_) & (!i_7_) & (!sk[52]) & (!g429) & (!g394)) + ((i_8_) & (i_6_) & (!i_7_) & (!sk[52]) & (!g429) & (g394)) + ((i_8_) & (i_6_) & (!i_7_) & (!sk[52]) & (g429) & (!g394)) + ((i_8_) & (i_6_) & (!i_7_) & (!sk[52]) & (g429) & (g394)) + ((i_8_) & (i_6_) & (!i_7_) & (sk[52]) & (g429) & (g394)) + ((i_8_) & (i_6_) & (i_7_) & (!sk[52]) & (!g429) & (!g394)) + ((i_8_) & (i_6_) & (i_7_) & (!sk[52]) & (!g429) & (g394)) + ((i_8_) & (i_6_) & (i_7_) & (!sk[52]) & (g429) & (!g394)) + ((i_8_) & (i_6_) & (i_7_) & (!sk[52]) & (g429) & (g394)));
	assign g1175 = (((!g68) & (!g86) & (g125) & (!g122) & (!sk[53]) & (g460)) + ((!g68) & (!g86) & (g125) & (g122) & (!sk[53]) & (!g460)) + ((!g68) & (!g86) & (g125) & (g122) & (!sk[53]) & (g460)) + ((!g68) & (g86) & (!g125) & (!g122) & (!sk[53]) & (!g460)) + ((!g68) & (g86) & (!g125) & (!g122) & (!sk[53]) & (g460)) + ((!g68) & (g86) & (!g125) & (g122) & (!sk[53]) & (!g460)) + ((!g68) & (g86) & (!g125) & (g122) & (!sk[53]) & (g460)) + ((!g68) & (g86) & (!g125) & (g122) & (sk[53]) & (!g460)) + ((!g68) & (g86) & (!g125) & (g122) & (sk[53]) & (g460)) + ((!g68) & (g86) & (g125) & (!g122) & (!sk[53]) & (!g460)) + ((!g68) & (g86) & (g125) & (!g122) & (!sk[53]) & (g460)) + ((!g68) & (g86) & (g125) & (!g122) & (sk[53]) & (!g460)) + ((!g68) & (g86) & (g125) & (!g122) & (sk[53]) & (g460)) + ((!g68) & (g86) & (g125) & (g122) & (!sk[53]) & (!g460)) + ((!g68) & (g86) & (g125) & (g122) & (!sk[53]) & (g460)) + ((!g68) & (g86) & (g125) & (g122) & (sk[53]) & (!g460)) + ((!g68) & (g86) & (g125) & (g122) & (sk[53]) & (g460)) + ((g68) & (!g86) & (g125) & (!g122) & (!sk[53]) & (g460)) + ((g68) & (!g86) & (g125) & (g122) & (!sk[53]) & (!g460)) + ((g68) & (!g86) & (g125) & (g122) & (!sk[53]) & (g460)) + ((g68) & (g86) & (!g125) & (!g122) & (!sk[53]) & (!g460)) + ((g68) & (g86) & (!g125) & (!g122) & (!sk[53]) & (g460)) + ((g68) & (g86) & (!g125) & (g122) & (!sk[53]) & (!g460)) + ((g68) & (g86) & (!g125) & (g122) & (!sk[53]) & (g460)) + ((g68) & (g86) & (!g125) & (g122) & (sk[53]) & (!g460)) + ((g68) & (g86) & (g125) & (!g122) & (!sk[53]) & (!g460)) + ((g68) & (g86) & (g125) & (!g122) & (!sk[53]) & (g460)) + ((g68) & (g86) & (g125) & (g122) & (!sk[53]) & (!g460)) + ((g68) & (g86) & (g125) & (g122) & (!sk[53]) & (g460)) + ((g68) & (g86) & (g125) & (g122) & (sk[53]) & (!g460)));
	assign g1176 = (((!g75) & (!g273) & (!g648) & (sk[54]) & (!g1174) & (!g1175)) + ((!g75) & (!g273) & (g648) & (!sk[54]) & (!g1174) & (g1175)) + ((!g75) & (!g273) & (g648) & (!sk[54]) & (g1174) & (!g1175)) + ((!g75) & (!g273) & (g648) & (!sk[54]) & (g1174) & (g1175)) + ((!g75) & (g273) & (!g648) & (!sk[54]) & (!g1174) & (!g1175)) + ((!g75) & (g273) & (!g648) & (!sk[54]) & (!g1174) & (g1175)) + ((!g75) & (g273) & (!g648) & (!sk[54]) & (g1174) & (!g1175)) + ((!g75) & (g273) & (!g648) & (!sk[54]) & (g1174) & (g1175)) + ((!g75) & (g273) & (g648) & (!sk[54]) & (!g1174) & (!g1175)) + ((!g75) & (g273) & (g648) & (!sk[54]) & (!g1174) & (g1175)) + ((!g75) & (g273) & (g648) & (!sk[54]) & (g1174) & (!g1175)) + ((!g75) & (g273) & (g648) & (!sk[54]) & (g1174) & (g1175)) + ((g75) & (!g273) & (!g648) & (sk[54]) & (!g1174) & (!g1175)) + ((g75) & (!g273) & (g648) & (!sk[54]) & (!g1174) & (g1175)) + ((g75) & (!g273) & (g648) & (!sk[54]) & (g1174) & (!g1175)) + ((g75) & (!g273) & (g648) & (!sk[54]) & (g1174) & (g1175)) + ((g75) & (!g273) & (g648) & (sk[54]) & (!g1174) & (!g1175)) + ((g75) & (g273) & (!g648) & (!sk[54]) & (!g1174) & (!g1175)) + ((g75) & (g273) & (!g648) & (!sk[54]) & (!g1174) & (g1175)) + ((g75) & (g273) & (!g648) & (!sk[54]) & (g1174) & (!g1175)) + ((g75) & (g273) & (!g648) & (!sk[54]) & (g1174) & (g1175)) + ((g75) & (g273) & (!g648) & (sk[54]) & (!g1174) & (!g1175)) + ((g75) & (g273) & (g648) & (!sk[54]) & (!g1174) & (!g1175)) + ((g75) & (g273) & (g648) & (!sk[54]) & (!g1174) & (g1175)) + ((g75) & (g273) & (g648) & (!sk[54]) & (g1174) & (!g1175)) + ((g75) & (g273) & (g648) & (!sk[54]) & (g1174) & (g1175)) + ((g75) & (g273) & (g648) & (sk[54]) & (!g1174) & (!g1175)));
	assign g1177 = (((!sk[55]) & (!g75) & (!g125) & (g187) & (!g1173) & (g1176)) + ((!sk[55]) & (!g75) & (!g125) & (g187) & (g1173) & (!g1176)) + ((!sk[55]) & (!g75) & (!g125) & (g187) & (g1173) & (g1176)) + ((!sk[55]) & (!g75) & (g125) & (!g187) & (!g1173) & (!g1176)) + ((!sk[55]) & (!g75) & (g125) & (!g187) & (!g1173) & (g1176)) + ((!sk[55]) & (!g75) & (g125) & (!g187) & (g1173) & (!g1176)) + ((!sk[55]) & (!g75) & (g125) & (!g187) & (g1173) & (g1176)) + ((!sk[55]) & (!g75) & (g125) & (g187) & (!g1173) & (!g1176)) + ((!sk[55]) & (!g75) & (g125) & (g187) & (!g1173) & (g1176)) + ((!sk[55]) & (!g75) & (g125) & (g187) & (g1173) & (!g1176)) + ((!sk[55]) & (!g75) & (g125) & (g187) & (g1173) & (g1176)) + ((!sk[55]) & (g75) & (!g125) & (g187) & (!g1173) & (g1176)) + ((!sk[55]) & (g75) & (!g125) & (g187) & (g1173) & (!g1176)) + ((!sk[55]) & (g75) & (!g125) & (g187) & (g1173) & (g1176)) + ((!sk[55]) & (g75) & (g125) & (!g187) & (!g1173) & (!g1176)) + ((!sk[55]) & (g75) & (g125) & (!g187) & (!g1173) & (g1176)) + ((!sk[55]) & (g75) & (g125) & (!g187) & (g1173) & (!g1176)) + ((!sk[55]) & (g75) & (g125) & (!g187) & (g1173) & (g1176)) + ((!sk[55]) & (g75) & (g125) & (g187) & (!g1173) & (!g1176)) + ((!sk[55]) & (g75) & (g125) & (g187) & (!g1173) & (g1176)) + ((!sk[55]) & (g75) & (g125) & (g187) & (g1173) & (!g1176)) + ((!sk[55]) & (g75) & (g125) & (g187) & (g1173) & (g1176)) + ((sk[55]) & (!g75) & (!g125) & (!g187) & (g1173) & (g1176)) + ((sk[55]) & (!g75) & (g125) & (!g187) & (g1173) & (g1176)) + ((sk[55]) & (g75) & (!g125) & (!g187) & (g1173) & (g1176)) + ((sk[55]) & (g75) & (!g125) & (g187) & (g1173) & (g1176)) + ((sk[55]) & (g75) & (g125) & (!g187) & (g1173) & (g1176)));
	assign g1178 = (((!sk[56]) & (!i_15_) & (!i_14_) & (g429) & (!g122)) + ((!sk[56]) & (!i_15_) & (!i_14_) & (g429) & (g122)) + ((!sk[56]) & (!i_15_) & (i_14_) & (g429) & (!g122)) + ((!sk[56]) & (!i_15_) & (i_14_) & (g429) & (g122)) + ((!sk[56]) & (i_15_) & (!i_14_) & (g429) & (!g122)) + ((!sk[56]) & (i_15_) & (!i_14_) & (g429) & (g122)) + ((!sk[56]) & (i_15_) & (i_14_) & (g429) & (!g122)) + ((!sk[56]) & (i_15_) & (i_14_) & (g429) & (g122)) + ((sk[56]) & (!i_15_) & (i_14_) & (g429) & (g122)) + ((sk[56]) & (i_15_) & (!i_14_) & (g429) & (g122)) + ((sk[56]) & (i_15_) & (i_14_) & (g429) & (g122)));
	assign g1179 = (((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g161) & (g429)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g161) & (g429)) + ((i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g161) & (g429)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g161) & (g429)) + ((i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g161) & (g429)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g161) & (g429)) + ((i_15_) & (i_12_) & (i_13_) & (i_14_) & (g161) & (g429)));
	assign g1180 = (((!g164) & (!g105) & (!g342) & (!g522) & (!g630) & (g847)) + ((!g164) & (g105) & (!g342) & (!g522) & (!g630) & (!g847)) + ((!g164) & (g105) & (!g342) & (!g522) & (!g630) & (g847)) + ((!g164) & (g105) & (!g342) & (!g522) & (g630) & (!g847)) + ((!g164) & (g105) & (!g342) & (!g522) & (g630) & (g847)) + ((!g164) & (g105) & (!g342) & (g522) & (!g630) & (!g847)) + ((!g164) & (g105) & (!g342) & (g522) & (!g630) & (g847)) + ((!g164) & (g105) & (!g342) & (g522) & (g630) & (!g847)) + ((!g164) & (g105) & (!g342) & (g522) & (g630) & (g847)) + ((!g164) & (g105) & (g342) & (!g522) & (!g630) & (!g847)) + ((!g164) & (g105) & (g342) & (!g522) & (!g630) & (g847)) + ((!g164) & (g105) & (g342) & (!g522) & (g630) & (!g847)) + ((!g164) & (g105) & (g342) & (!g522) & (g630) & (g847)) + ((!g164) & (g105) & (g342) & (g522) & (!g630) & (!g847)) + ((!g164) & (g105) & (g342) & (g522) & (!g630) & (g847)) + ((!g164) & (g105) & (g342) & (g522) & (g630) & (!g847)) + ((!g164) & (g105) & (g342) & (g522) & (g630) & (g847)) + ((g164) & (!g105) & (!g342) & (!g522) & (!g630) & (g847)) + ((g164) & (g105) & (!g342) & (!g522) & (!g630) & (g847)));
	assign g1181 = (((!sk[59]) & (g429) & (!g123)) + ((!sk[59]) & (g429) & (g123)) + ((sk[59]) & (g429) & (!g123)));
	assign g1182 = (((!g164) & (!g975) & (!sk[60]) & (g952) & (!g1181)) + ((!g164) & (!g975) & (!sk[60]) & (g952) & (g1181)) + ((!g164) & (!g975) & (sk[60]) & (!g952) & (!g1181)) + ((!g164) & (g975) & (!sk[60]) & (g952) & (!g1181)) + ((!g164) & (g975) & (!sk[60]) & (g952) & (g1181)) + ((!g164) & (g975) & (sk[60]) & (!g952) & (!g1181)) + ((g164) & (!g975) & (!sk[60]) & (g952) & (!g1181)) + ((g164) & (!g975) & (!sk[60]) & (g952) & (g1181)) + ((g164) & (g975) & (!sk[60]) & (g952) & (!g1181)) + ((g164) & (g975) & (!sk[60]) & (g952) & (g1181)) + ((g164) & (g975) & (sk[60]) & (!g952) & (!g1181)));
	assign g1183 = (((!sk[61]) & (!g1049) & (!g1115) & (g1177) & (!g1453) & (g1182)) + ((!sk[61]) & (!g1049) & (!g1115) & (g1177) & (g1453) & (!g1182)) + ((!sk[61]) & (!g1049) & (!g1115) & (g1177) & (g1453) & (g1182)) + ((!sk[61]) & (!g1049) & (g1115) & (!g1177) & (!g1453) & (!g1182)) + ((!sk[61]) & (!g1049) & (g1115) & (!g1177) & (!g1453) & (g1182)) + ((!sk[61]) & (!g1049) & (g1115) & (!g1177) & (g1453) & (!g1182)) + ((!sk[61]) & (!g1049) & (g1115) & (!g1177) & (g1453) & (g1182)) + ((!sk[61]) & (!g1049) & (g1115) & (g1177) & (!g1453) & (!g1182)) + ((!sk[61]) & (!g1049) & (g1115) & (g1177) & (!g1453) & (g1182)) + ((!sk[61]) & (!g1049) & (g1115) & (g1177) & (g1453) & (!g1182)) + ((!sk[61]) & (!g1049) & (g1115) & (g1177) & (g1453) & (g1182)) + ((!sk[61]) & (g1049) & (!g1115) & (g1177) & (!g1453) & (g1182)) + ((!sk[61]) & (g1049) & (!g1115) & (g1177) & (g1453) & (!g1182)) + ((!sk[61]) & (g1049) & (!g1115) & (g1177) & (g1453) & (g1182)) + ((!sk[61]) & (g1049) & (g1115) & (!g1177) & (!g1453) & (!g1182)) + ((!sk[61]) & (g1049) & (g1115) & (!g1177) & (!g1453) & (g1182)) + ((!sk[61]) & (g1049) & (g1115) & (!g1177) & (g1453) & (!g1182)) + ((!sk[61]) & (g1049) & (g1115) & (!g1177) & (g1453) & (g1182)) + ((!sk[61]) & (g1049) & (g1115) & (g1177) & (!g1453) & (!g1182)) + ((!sk[61]) & (g1049) & (g1115) & (g1177) & (!g1453) & (g1182)) + ((!sk[61]) & (g1049) & (g1115) & (g1177) & (g1453) & (!g1182)) + ((!sk[61]) & (g1049) & (g1115) & (g1177) & (g1453) & (g1182)) + ((sk[61]) & (!g1049) & (!g1115) & (g1177) & (g1453) & (g1182)));
	assign g1184 = (((!g122) & (!sk[62]) & (!g487) & (g1029)) + ((!g122) & (!sk[62]) & (g487) & (!g1029)) + ((!g122) & (!sk[62]) & (g487) & (g1029)) + ((g122) & (!sk[62]) & (!g487) & (g1029)) + ((g122) & (!sk[62]) & (g487) & (!g1029)) + ((g122) & (!sk[62]) & (g487) & (g1029)) + ((g122) & (sk[62]) & (!g487) & (!g1029)) + ((g122) & (sk[62]) & (g487) & (!g1029)) + ((g122) & (sk[62]) & (g487) & (g1029)));
	assign g1185 = (((!i_14_) & (!g107) & (!sk[63]) & (g91) & (!g123)) + ((!i_14_) & (!g107) & (!sk[63]) & (g91) & (g123)) + ((!i_14_) & (!g107) & (sk[63]) & (!g91) & (!g123)) + ((!i_14_) & (g107) & (!sk[63]) & (g91) & (!g123)) + ((!i_14_) & (g107) & (!sk[63]) & (g91) & (g123)) + ((!i_14_) & (g107) & (sk[63]) & (!g91) & (!g123)) + ((i_14_) & (!g107) & (!sk[63]) & (g91) & (!g123)) + ((i_14_) & (!g107) & (!sk[63]) & (g91) & (g123)) + ((i_14_) & (!g107) & (sk[63]) & (!g91) & (!g123)) + ((i_14_) & (!g107) & (sk[63]) & (g91) & (!g123)) + ((i_14_) & (g107) & (!sk[63]) & (g91) & (!g123)) + ((i_14_) & (g107) & (!sk[63]) & (g91) & (g123)) + ((i_14_) & (g107) & (sk[63]) & (!g91) & (!g123)));
	assign g1186 = (((!g105) & (!g487) & (!g484) & (sk[64]) & (g652)) + ((!g105) & (!g487) & (g484) & (!sk[64]) & (!g652)) + ((!g105) & (!g487) & (g484) & (!sk[64]) & (g652)) + ((!g105) & (!g487) & (g484) & (sk[64]) & (!g652)) + ((!g105) & (!g487) & (g484) & (sk[64]) & (g652)) + ((!g105) & (g487) & (!g484) & (sk[64]) & (!g652)) + ((!g105) & (g487) & (!g484) & (sk[64]) & (g652)) + ((!g105) & (g487) & (g484) & (!sk[64]) & (!g652)) + ((!g105) & (g487) & (g484) & (!sk[64]) & (g652)) + ((!g105) & (g487) & (g484) & (sk[64]) & (!g652)) + ((!g105) & (g487) & (g484) & (sk[64]) & (g652)) + ((g105) & (!g487) & (g484) & (!sk[64]) & (!g652)) + ((g105) & (!g487) & (g484) & (!sk[64]) & (g652)) + ((g105) & (g487) & (g484) & (!sk[64]) & (!g652)) + ((g105) & (g487) & (g484) & (!sk[64]) & (g652)));
	assign g1187 = (((!g105) & (!g358) & (!sk[65]) & (g852) & (!g1186) & (g1452)) + ((!g105) & (!g358) & (!sk[65]) & (g852) & (g1186) & (!g1452)) + ((!g105) & (!g358) & (!sk[65]) & (g852) & (g1186) & (g1452)) + ((!g105) & (!g358) & (sk[65]) & (!g852) & (!g1186) & (!g1452)) + ((!g105) & (g358) & (!sk[65]) & (!g852) & (!g1186) & (!g1452)) + ((!g105) & (g358) & (!sk[65]) & (!g852) & (!g1186) & (g1452)) + ((!g105) & (g358) & (!sk[65]) & (!g852) & (g1186) & (!g1452)) + ((!g105) & (g358) & (!sk[65]) & (!g852) & (g1186) & (g1452)) + ((!g105) & (g358) & (!sk[65]) & (g852) & (!g1186) & (!g1452)) + ((!g105) & (g358) & (!sk[65]) & (g852) & (!g1186) & (g1452)) + ((!g105) & (g358) & (!sk[65]) & (g852) & (g1186) & (!g1452)) + ((!g105) & (g358) & (!sk[65]) & (g852) & (g1186) & (g1452)) + ((g105) & (!g358) & (!sk[65]) & (g852) & (!g1186) & (g1452)) + ((g105) & (!g358) & (!sk[65]) & (g852) & (g1186) & (!g1452)) + ((g105) & (!g358) & (!sk[65]) & (g852) & (g1186) & (g1452)) + ((g105) & (!g358) & (sk[65]) & (!g852) & (!g1186) & (!g1452)) + ((g105) & (!g358) & (sk[65]) & (g852) & (!g1186) & (!g1452)) + ((g105) & (g358) & (!sk[65]) & (!g852) & (!g1186) & (!g1452)) + ((g105) & (g358) & (!sk[65]) & (!g852) & (!g1186) & (g1452)) + ((g105) & (g358) & (!sk[65]) & (!g852) & (g1186) & (!g1452)) + ((g105) & (g358) & (!sk[65]) & (!g852) & (g1186) & (g1452)) + ((g105) & (g358) & (!sk[65]) & (g852) & (!g1186) & (!g1452)) + ((g105) & (g358) & (!sk[65]) & (g852) & (!g1186) & (g1452)) + ((g105) & (g358) & (!sk[65]) & (g852) & (g1186) & (!g1452)) + ((g105) & (g358) & (!sk[65]) & (g852) & (g1186) & (g1452)) + ((g105) & (g358) & (sk[65]) & (!g852) & (!g1186) & (!g1452)) + ((g105) & (g358) & (sk[65]) & (g852) & (!g1186) & (!g1452)));
	assign g1188 = (((!g75) & (!g122) & (!g185) & (!g486) & (!g487) & (!g708)) + ((!g75) & (g122) & (!g185) & (!g486) & (!g487) & (!g708)) + ((g75) & (!g122) & (!g185) & (!g486) & (!g487) & (!g708)) + ((g75) & (!g122) & (!g185) & (!g486) & (g487) & (!g708)) + ((g75) & (!g122) & (!g185) & (g486) & (!g487) & (!g708)) + ((g75) & (!g122) & (!g185) & (g486) & (g487) & (!g708)) + ((g75) & (!g122) & (g185) & (!g486) & (!g487) & (!g708)) + ((g75) & (!g122) & (g185) & (!g486) & (g487) & (!g708)) + ((g75) & (!g122) & (g185) & (g486) & (!g487) & (!g708)) + ((g75) & (!g122) & (g185) & (g486) & (g487) & (!g708)) + ((g75) & (g122) & (!g185) & (!g486) & (!g487) & (!g708)) + ((g75) & (g122) & (!g185) & (!g486) & (g487) & (!g708)) + ((g75) & (g122) & (!g185) & (g486) & (!g487) & (!g708)) + ((g75) & (g122) & (!g185) & (g486) & (g487) & (!g708)));
	assign g1189 = (((!g1184) & (!g527) & (!sk[67]) & (g1185) & (!g1187) & (g1188)) + ((!g1184) & (!g527) & (!sk[67]) & (g1185) & (g1187) & (!g1188)) + ((!g1184) & (!g527) & (!sk[67]) & (g1185) & (g1187) & (g1188)) + ((!g1184) & (!g527) & (sk[67]) & (!g1185) & (g1187) & (g1188)) + ((!g1184) & (g527) & (!sk[67]) & (!g1185) & (!g1187) & (!g1188)) + ((!g1184) & (g527) & (!sk[67]) & (!g1185) & (!g1187) & (g1188)) + ((!g1184) & (g527) & (!sk[67]) & (!g1185) & (g1187) & (!g1188)) + ((!g1184) & (g527) & (!sk[67]) & (!g1185) & (g1187) & (g1188)) + ((!g1184) & (g527) & (!sk[67]) & (g1185) & (!g1187) & (!g1188)) + ((!g1184) & (g527) & (!sk[67]) & (g1185) & (!g1187) & (g1188)) + ((!g1184) & (g527) & (!sk[67]) & (g1185) & (g1187) & (!g1188)) + ((!g1184) & (g527) & (!sk[67]) & (g1185) & (g1187) & (g1188)) + ((g1184) & (!g527) & (!sk[67]) & (g1185) & (!g1187) & (g1188)) + ((g1184) & (!g527) & (!sk[67]) & (g1185) & (g1187) & (!g1188)) + ((g1184) & (!g527) & (!sk[67]) & (g1185) & (g1187) & (g1188)) + ((g1184) & (g527) & (!sk[67]) & (!g1185) & (!g1187) & (!g1188)) + ((g1184) & (g527) & (!sk[67]) & (!g1185) & (!g1187) & (g1188)) + ((g1184) & (g527) & (!sk[67]) & (!g1185) & (g1187) & (!g1188)) + ((g1184) & (g527) & (!sk[67]) & (!g1185) & (g1187) & (g1188)) + ((g1184) & (g527) & (!sk[67]) & (g1185) & (!g1187) & (!g1188)) + ((g1184) & (g527) & (!sk[67]) & (g1185) & (!g1187) & (g1188)) + ((g1184) & (g527) & (!sk[67]) & (g1185) & (g1187) & (!g1188)) + ((g1184) & (g527) & (!sk[67]) & (g1185) & (g1187) & (g1188)));
	assign g1190 = (((!g154) & (!sk[68]) & (!g334) & (g489) & (!g624)) + ((!g154) & (!sk[68]) & (!g334) & (g489) & (g624)) + ((!g154) & (!sk[68]) & (g334) & (g489) & (!g624)) + ((!g154) & (!sk[68]) & (g334) & (g489) & (g624)) + ((!g154) & (sk[68]) & (!g334) & (!g489) & (!g624)) + ((!g154) & (sk[68]) & (!g334) & (!g489) & (g624)) + ((!g154) & (sk[68]) & (!g334) & (g489) & (!g624)) + ((!g154) & (sk[68]) & (!g334) & (g489) & (g624)) + ((!g154) & (sk[68]) & (g334) & (!g489) & (!g624)) + ((!g154) & (sk[68]) & (g334) & (g489) & (!g624)) + ((!g154) & (sk[68]) & (g334) & (g489) & (g624)) + ((g154) & (!sk[68]) & (!g334) & (g489) & (!g624)) + ((g154) & (!sk[68]) & (!g334) & (g489) & (g624)) + ((g154) & (!sk[68]) & (g334) & (g489) & (!g624)) + ((g154) & (!sk[68]) & (g334) & (g489) & (g624)));
	assign g1191 = (((!g18) & (!g33) & (!g97) & (!g98) & (!g122) & (!g1190)) + ((!g18) & (!g33) & (!g97) & (g98) & (!g122) & (!g1190)) + ((!g18) & (!g33) & (g97) & (!g98) & (!g122) & (!g1190)) + ((!g18) & (!g33) & (g97) & (!g98) & (g122) & (!g1190)) + ((!g18) & (!g33) & (g97) & (g98) & (!g122) & (!g1190)) + ((!g18) & (g33) & (!g97) & (!g98) & (!g122) & (!g1190)) + ((!g18) & (g33) & (!g97) & (g98) & (!g122) & (!g1190)) + ((!g18) & (g33) & (g97) & (!g98) & (!g122) & (!g1190)) + ((!g18) & (g33) & (g97) & (g98) & (!g122) & (!g1190)) + ((g18) & (!g33) & (!g97) & (!g98) & (!g122) & (!g1190)) + ((g18) & (!g33) & (!g97) & (g98) & (!g122) & (!g1190)) + ((g18) & (!g33) & (g97) & (!g98) & (!g122) & (!g1190)) + ((g18) & (!g33) & (g97) & (g98) & (!g122) & (!g1190)) + ((g18) & (g33) & (!g97) & (!g98) & (!g122) & (!g1190)) + ((g18) & (g33) & (!g97) & (g98) & (!g122) & (!g1190)) + ((g18) & (g33) & (g97) & (!g98) & (!g122) & (!g1190)) + ((g18) & (g33) & (g97) & (g98) & (!g122) & (!g1190)));
	assign g1192 = (((!sk[70]) & (!g105) & (!g993) & (g1191)) + ((!sk[70]) & (!g105) & (g993) & (!g1191)) + ((!sk[70]) & (!g105) & (g993) & (g1191)) + ((!sk[70]) & (g105) & (!g993) & (g1191)) + ((!sk[70]) & (g105) & (g993) & (!g1191)) + ((!sk[70]) & (g105) & (g993) & (g1191)) + ((sk[70]) & (!g105) & (!g993) & (g1191)) + ((sk[70]) & (g105) & (!g993) & (g1191)) + ((sk[70]) & (g105) & (g993) & (g1191)));
	assign g1193 = (((!sk[71]) & (!i_8_) & (!g73) & (g578) & (!g461)) + ((!sk[71]) & (!i_8_) & (!g73) & (g578) & (g461)) + ((!sk[71]) & (!i_8_) & (g73) & (g578) & (!g461)) + ((!sk[71]) & (!i_8_) & (g73) & (g578) & (g461)) + ((!sk[71]) & (i_8_) & (!g73) & (g578) & (!g461)) + ((!sk[71]) & (i_8_) & (!g73) & (g578) & (g461)) + ((!sk[71]) & (i_8_) & (g73) & (g578) & (!g461)) + ((!sk[71]) & (i_8_) & (g73) & (g578) & (g461)) + ((sk[71]) & (i_8_) & (g73) & (!g578) & (g461)) + ((sk[71]) & (i_8_) & (g73) & (g578) & (!g461)) + ((sk[71]) & (i_8_) & (g73) & (g578) & (g461)));
	assign g1194 = (((!g17) & (!g76) & (g122) & (!g91) & (!sk[72]) & (g460)) + ((!g17) & (!g76) & (g122) & (!g91) & (sk[72]) & (!g460)) + ((!g17) & (!g76) & (g122) & (!g91) & (sk[72]) & (g460)) + ((!g17) & (!g76) & (g122) & (g91) & (!sk[72]) & (!g460)) + ((!g17) & (!g76) & (g122) & (g91) & (!sk[72]) & (g460)) + ((!g17) & (g76) & (!g122) & (!g91) & (!sk[72]) & (!g460)) + ((!g17) & (g76) & (!g122) & (!g91) & (!sk[72]) & (g460)) + ((!g17) & (g76) & (!g122) & (g91) & (!sk[72]) & (!g460)) + ((!g17) & (g76) & (!g122) & (g91) & (!sk[72]) & (g460)) + ((!g17) & (g76) & (g122) & (!g91) & (!sk[72]) & (!g460)) + ((!g17) & (g76) & (g122) & (!g91) & (!sk[72]) & (g460)) + ((!g17) & (g76) & (g122) & (g91) & (!sk[72]) & (!g460)) + ((!g17) & (g76) & (g122) & (g91) & (!sk[72]) & (g460)) + ((g17) & (!g76) & (g122) & (!g91) & (!sk[72]) & (g460)) + ((g17) & (!g76) & (g122) & (!g91) & (sk[72]) & (!g460)) + ((g17) & (!g76) & (g122) & (!g91) & (sk[72]) & (g460)) + ((g17) & (!g76) & (g122) & (g91) & (!sk[72]) & (!g460)) + ((g17) & (!g76) & (g122) & (g91) & (!sk[72]) & (g460)) + ((g17) & (!g76) & (g122) & (g91) & (sk[72]) & (!g460)) + ((g17) & (!g76) & (g122) & (g91) & (sk[72]) & (g460)) + ((g17) & (g76) & (!g122) & (!g91) & (!sk[72]) & (!g460)) + ((g17) & (g76) & (!g122) & (!g91) & (!sk[72]) & (g460)) + ((g17) & (g76) & (!g122) & (g91) & (!sk[72]) & (!g460)) + ((g17) & (g76) & (!g122) & (g91) & (!sk[72]) & (g460)) + ((g17) & (g76) & (g122) & (!g91) & (!sk[72]) & (!g460)) + ((g17) & (g76) & (g122) & (!g91) & (!sk[72]) & (g460)) + ((g17) & (g76) & (g122) & (!g91) & (sk[72]) & (!g460)) + ((g17) & (g76) & (g122) & (g91) & (!sk[72]) & (!g460)) + ((g17) & (g76) & (g122) & (g91) & (!sk[72]) & (g460)) + ((g17) & (g76) & (g122) & (g91) & (sk[72]) & (!g460)));
	assign g1195 = (((!g28) & (!g122) & (g180) & (!sk[73]) & (!g275)) + ((!g28) & (!g122) & (g180) & (!sk[73]) & (g275)) + ((!g28) & (g122) & (!g180) & (sk[73]) & (g275)) + ((!g28) & (g122) & (g180) & (!sk[73]) & (!g275)) + ((!g28) & (g122) & (g180) & (!sk[73]) & (g275)) + ((!g28) & (g122) & (g180) & (sk[73]) & (!g275)) + ((!g28) & (g122) & (g180) & (sk[73]) & (g275)) + ((g28) & (!g122) & (g180) & (!sk[73]) & (!g275)) + ((g28) & (!g122) & (g180) & (!sk[73]) & (g275)) + ((g28) & (g122) & (!g180) & (sk[73]) & (!g275)) + ((g28) & (g122) & (!g180) & (sk[73]) & (g275)) + ((g28) & (g122) & (g180) & (!sk[73]) & (!g275)) + ((g28) & (g122) & (g180) & (!sk[73]) & (g275)) + ((g28) & (g122) & (g180) & (sk[73]) & (!g275)) + ((g28) & (g122) & (g180) & (sk[73]) & (g275)));
	assign g1196 = (((!i_12_) & (!i_13_) & (!i_14_) & (!g17) & (g27) & (g125)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g17) & (g27) & (g125)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g17) & (g27) & (g125)) + ((!i_12_) & (i_13_) & (!i_14_) & (g17) & (!g27) & (g125)) + ((!i_12_) & (i_13_) & (!i_14_) & (g17) & (g27) & (g125)) + ((i_12_) & (!i_13_) & (!i_14_) & (!g17) & (g27) & (g125)) + ((i_12_) & (!i_13_) & (!i_14_) & (g17) & (g27) & (g125)) + ((i_12_) & (!i_13_) & (i_14_) & (!g17) & (g27) & (g125)) + ((i_12_) & (!i_13_) & (i_14_) & (g17) & (!g27) & (g125)) + ((i_12_) & (!i_13_) & (i_14_) & (g17) & (g27) & (g125)));
	assign g1197 = (((!g276) & (!g1193) & (!sk[75]) & (g1194) & (!g1195) & (g1196)) + ((!g276) & (!g1193) & (!sk[75]) & (g1194) & (g1195) & (!g1196)) + ((!g276) & (!g1193) & (!sk[75]) & (g1194) & (g1195) & (g1196)) + ((!g276) & (!g1193) & (sk[75]) & (!g1194) & (!g1195) & (!g1196)) + ((!g276) & (g1193) & (!sk[75]) & (!g1194) & (!g1195) & (!g1196)) + ((!g276) & (g1193) & (!sk[75]) & (!g1194) & (!g1195) & (g1196)) + ((!g276) & (g1193) & (!sk[75]) & (!g1194) & (g1195) & (!g1196)) + ((!g276) & (g1193) & (!sk[75]) & (!g1194) & (g1195) & (g1196)) + ((!g276) & (g1193) & (!sk[75]) & (g1194) & (!g1195) & (!g1196)) + ((!g276) & (g1193) & (!sk[75]) & (g1194) & (!g1195) & (g1196)) + ((!g276) & (g1193) & (!sk[75]) & (g1194) & (g1195) & (!g1196)) + ((!g276) & (g1193) & (!sk[75]) & (g1194) & (g1195) & (g1196)) + ((g276) & (!g1193) & (!sk[75]) & (g1194) & (!g1195) & (g1196)) + ((g276) & (!g1193) & (!sk[75]) & (g1194) & (g1195) & (!g1196)) + ((g276) & (!g1193) & (!sk[75]) & (g1194) & (g1195) & (g1196)) + ((g276) & (g1193) & (!sk[75]) & (!g1194) & (!g1195) & (!g1196)) + ((g276) & (g1193) & (!sk[75]) & (!g1194) & (!g1195) & (g1196)) + ((g276) & (g1193) & (!sk[75]) & (!g1194) & (g1195) & (!g1196)) + ((g276) & (g1193) & (!sk[75]) & (!g1194) & (g1195) & (g1196)) + ((g276) & (g1193) & (!sk[75]) & (g1194) & (!g1195) & (!g1196)) + ((g276) & (g1193) & (!sk[75]) & (g1194) & (!g1195) & (g1196)) + ((g276) & (g1193) & (!sk[75]) & (g1194) & (g1195) & (!g1196)) + ((g276) & (g1193) & (!sk[75]) & (g1194) & (g1195) & (g1196)));
	assign g1198 = (((!g164) & (!g123) & (g334) & (!g489) & (g624) & (g1107)) + ((!g164) & (g123) & (!g334) & (!g489) & (!g624) & (!g1107)) + ((!g164) & (g123) & (!g334) & (!g489) & (!g624) & (g1107)) + ((!g164) & (g123) & (!g334) & (!g489) & (g624) & (!g1107)) + ((!g164) & (g123) & (!g334) & (!g489) & (g624) & (g1107)) + ((!g164) & (g123) & (!g334) & (g489) & (!g624) & (!g1107)) + ((!g164) & (g123) & (!g334) & (g489) & (!g624) & (g1107)) + ((!g164) & (g123) & (!g334) & (g489) & (g624) & (!g1107)) + ((!g164) & (g123) & (!g334) & (g489) & (g624) & (g1107)) + ((!g164) & (g123) & (g334) & (!g489) & (!g624) & (!g1107)) + ((!g164) & (g123) & (g334) & (!g489) & (!g624) & (g1107)) + ((!g164) & (g123) & (g334) & (!g489) & (g624) & (!g1107)) + ((!g164) & (g123) & (g334) & (!g489) & (g624) & (g1107)) + ((!g164) & (g123) & (g334) & (g489) & (!g624) & (!g1107)) + ((!g164) & (g123) & (g334) & (g489) & (!g624) & (g1107)) + ((!g164) & (g123) & (g334) & (g489) & (g624) & (!g1107)) + ((!g164) & (g123) & (g334) & (g489) & (g624) & (g1107)) + ((g164) & (!g123) & (g334) & (!g489) & (g624) & (g1107)) + ((g164) & (g123) & (g334) & (!g489) & (g624) & (g1107)));
	assign g1199 = (((!i_12_) & (!i_13_) & (!i_14_) & (!g17) & (!g27) & (g86)) + ((!i_12_) & (!i_13_) & (!i_14_) & (!g17) & (g27) & (!g86)) + ((!i_12_) & (!i_13_) & (!i_14_) & (!g17) & (g27) & (g86)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g17) & (!g27) & (g86)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g17) & (g27) & (!g86)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g17) & (g27) & (g86)) + ((!i_12_) & (!i_13_) & (i_14_) & (g17) & (!g27) & (!g86)) + ((!i_12_) & (!i_13_) & (i_14_) & (g17) & (!g27) & (g86)) + ((!i_12_) & (!i_13_) & (i_14_) & (g17) & (g27) & (!g86)) + ((!i_12_) & (!i_13_) & (i_14_) & (g17) & (g27) & (g86)) + ((!i_12_) & (i_13_) & (i_14_) & (g17) & (!g27) & (!g86)) + ((!i_12_) & (i_13_) & (i_14_) & (g17) & (!g27) & (g86)) + ((!i_12_) & (i_13_) & (i_14_) & (g17) & (g27) & (!g86)) + ((!i_12_) & (i_13_) & (i_14_) & (g17) & (g27) & (g86)) + ((i_12_) & (i_13_) & (i_14_) & (g17) & (!g27) & (!g86)) + ((i_12_) & (i_13_) & (i_14_) & (g17) & (!g27) & (g86)) + ((i_12_) & (i_13_) & (i_14_) & (g17) & (g27) & (!g86)) + ((i_12_) & (i_13_) & (i_14_) & (g17) & (g27) & (g86)));
	assign g1200 = (((!g75) & (!g97) & (!g98) & (!g725) & (!g1029) & (!g1199)) + ((!g75) & (!g97) & (!g98) & (!g725) & (!g1029) & (g1199)) + ((!g75) & (!g97) & (!g98) & (!g725) & (g1029) & (!g1199)) + ((!g75) & (!g97) & (!g98) & (!g725) & (g1029) & (g1199)) + ((!g75) & (!g97) & (!g98) & (g725) & (!g1029) & (!g1199)) + ((!g75) & (!g97) & (!g98) & (g725) & (!g1029) & (g1199)) + ((!g75) & (!g97) & (!g98) & (g725) & (g1029) & (!g1199)) + ((!g75) & (!g97) & (!g98) & (g725) & (g1029) & (g1199)) + ((!g75) & (!g97) & (g98) & (!g725) & (!g1029) & (!g1199)) + ((!g75) & (!g97) & (g98) & (!g725) & (!g1029) & (g1199)) + ((!g75) & (!g97) & (g98) & (!g725) & (g1029) & (!g1199)) + ((!g75) & (!g97) & (g98) & (!g725) & (g1029) & (g1199)) + ((!g75) & (!g97) & (g98) & (g725) & (!g1029) & (!g1199)) + ((!g75) & (!g97) & (g98) & (g725) & (!g1029) & (g1199)) + ((!g75) & (!g97) & (g98) & (g725) & (g1029) & (!g1199)) + ((!g75) & (!g97) & (g98) & (g725) & (g1029) & (g1199)) + ((!g75) & (g97) & (!g98) & (!g725) & (!g1029) & (!g1199)) + ((!g75) & (g97) & (!g98) & (!g725) & (!g1029) & (g1199)) + ((!g75) & (g97) & (!g98) & (!g725) & (g1029) & (!g1199)) + ((!g75) & (g97) & (!g98) & (!g725) & (g1029) & (g1199)) + ((!g75) & (g97) & (!g98) & (g725) & (!g1029) & (!g1199)) + ((!g75) & (g97) & (!g98) & (g725) & (!g1029) & (g1199)) + ((!g75) & (g97) & (!g98) & (g725) & (g1029) & (g1199)) + ((!g75) & (g97) & (g98) & (!g725) & (!g1029) & (!g1199)) + ((!g75) & (g97) & (g98) & (!g725) & (!g1029) & (g1199)) + ((!g75) & (g97) & (g98) & (!g725) & (g1029) & (!g1199)) + ((!g75) & (g97) & (g98) & (!g725) & (g1029) & (g1199)) + ((!g75) & (g97) & (g98) & (g725) & (!g1029) & (!g1199)) + ((!g75) & (g97) & (g98) & (g725) & (!g1029) & (g1199)) + ((!g75) & (g97) & (g98) & (g725) & (g1029) & (!g1199)) + ((!g75) & (g97) & (g98) & (g725) & (g1029) & (g1199)));
	assign g1201 = (((!g18) & (!g33) & (!g75) & (!g1030) & (sk[79]) & (!g1046)) + ((!g18) & (!g33) & (g75) & (!g1030) & (!sk[79]) & (g1046)) + ((!g18) & (!g33) & (g75) & (!g1030) & (sk[79]) & (!g1046)) + ((!g18) & (!g33) & (g75) & (g1030) & (!sk[79]) & (!g1046)) + ((!g18) & (!g33) & (g75) & (g1030) & (!sk[79]) & (g1046)) + ((!g18) & (g33) & (!g75) & (!g1030) & (!sk[79]) & (!g1046)) + ((!g18) & (g33) & (!g75) & (!g1030) & (!sk[79]) & (g1046)) + ((!g18) & (g33) & (!g75) & (g1030) & (!sk[79]) & (!g1046)) + ((!g18) & (g33) & (!g75) & (g1030) & (!sk[79]) & (g1046)) + ((!g18) & (g33) & (g75) & (!g1030) & (!sk[79]) & (!g1046)) + ((!g18) & (g33) & (g75) & (!g1030) & (!sk[79]) & (g1046)) + ((!g18) & (g33) & (g75) & (!g1030) & (sk[79]) & (!g1046)) + ((!g18) & (g33) & (g75) & (g1030) & (!sk[79]) & (!g1046)) + ((!g18) & (g33) & (g75) & (g1030) & (!sk[79]) & (g1046)) + ((g18) & (!g33) & (g75) & (!g1030) & (!sk[79]) & (g1046)) + ((g18) & (!g33) & (g75) & (!g1030) & (sk[79]) & (!g1046)) + ((g18) & (!g33) & (g75) & (g1030) & (!sk[79]) & (!g1046)) + ((g18) & (!g33) & (g75) & (g1030) & (!sk[79]) & (g1046)) + ((g18) & (g33) & (!g75) & (!g1030) & (!sk[79]) & (!g1046)) + ((g18) & (g33) & (!g75) & (!g1030) & (!sk[79]) & (g1046)) + ((g18) & (g33) & (!g75) & (g1030) & (!sk[79]) & (!g1046)) + ((g18) & (g33) & (!g75) & (g1030) & (!sk[79]) & (g1046)) + ((g18) & (g33) & (g75) & (!g1030) & (!sk[79]) & (!g1046)) + ((g18) & (g33) & (g75) & (!g1030) & (!sk[79]) & (g1046)) + ((g18) & (g33) & (g75) & (!g1030) & (sk[79]) & (!g1046)) + ((g18) & (g33) & (g75) & (g1030) & (!sk[79]) & (!g1046)) + ((g18) & (g33) & (g75) & (g1030) & (!sk[79]) & (g1046)));
	assign g1202 = (((!g181) & (!g1096) & (g1197) & (g1198) & (!g1200) & (g1201)));
	assign g1203 = (((!sk[81]) & (g461) & (!g477)) + ((!sk[81]) & (g461) & (g477)) + ((sk[81]) & (!g461) & (!g477)));
	assign g1204 = (((!i_11_) & (!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g34)) + ((!i_11_) & (!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g34)) + ((!i_11_) & (!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g34)) + ((!i_11_) & (!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g34)) + ((!i_11_) & (!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g34)) + ((!i_11_) & (!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g34)) + ((!i_11_) & (i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (g34)) + ((!i_11_) & (i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g34)) + ((!i_11_) & (i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g34)) + ((i_11_) & (!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g34)) + ((i_11_) & (!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g34)) + ((i_11_) & (!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g34)) + ((i_11_) & (i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (g34)) + ((i_11_) & (i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g34)) + ((i_11_) & (i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g34)) + ((i_11_) & (i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g34)));
	assign g1205 = (((!g179) & (!g853) & (g1203) & (!sk[83]) & (!g1204)) + ((!g179) & (!g853) & (g1203) & (!sk[83]) & (g1204)) + ((!g179) & (!g853) & (g1203) & (sk[83]) & (!g1204)) + ((!g179) & (g853) & (g1203) & (!sk[83]) & (!g1204)) + ((!g179) & (g853) & (g1203) & (!sk[83]) & (g1204)) + ((g179) & (!g853) & (g1203) & (!sk[83]) & (!g1204)) + ((g179) & (!g853) & (g1203) & (!sk[83]) & (g1204)) + ((g179) & (g853) & (g1203) & (!sk[83]) & (!g1204)) + ((g179) & (g853) & (g1203) & (!sk[83]) & (g1204)));
	assign g1206 = (((!sk[84]) & (!g154) & (!g122) & (g1007) & (!g1205) & (g999)) + ((!sk[84]) & (!g154) & (!g122) & (g1007) & (g1205) & (!g999)) + ((!sk[84]) & (!g154) & (!g122) & (g1007) & (g1205) & (g999)) + ((!sk[84]) & (!g154) & (g122) & (!g1007) & (!g1205) & (!g999)) + ((!sk[84]) & (!g154) & (g122) & (!g1007) & (!g1205) & (g999)) + ((!sk[84]) & (!g154) & (g122) & (!g1007) & (g1205) & (!g999)) + ((!sk[84]) & (!g154) & (g122) & (!g1007) & (g1205) & (g999)) + ((!sk[84]) & (!g154) & (g122) & (g1007) & (!g1205) & (!g999)) + ((!sk[84]) & (!g154) & (g122) & (g1007) & (!g1205) & (g999)) + ((!sk[84]) & (!g154) & (g122) & (g1007) & (g1205) & (!g999)) + ((!sk[84]) & (!g154) & (g122) & (g1007) & (g1205) & (g999)) + ((!sk[84]) & (g154) & (!g122) & (g1007) & (!g1205) & (g999)) + ((!sk[84]) & (g154) & (!g122) & (g1007) & (g1205) & (!g999)) + ((!sk[84]) & (g154) & (!g122) & (g1007) & (g1205) & (g999)) + ((!sk[84]) & (g154) & (g122) & (!g1007) & (!g1205) & (!g999)) + ((!sk[84]) & (g154) & (g122) & (!g1007) & (!g1205) & (g999)) + ((!sk[84]) & (g154) & (g122) & (!g1007) & (g1205) & (!g999)) + ((!sk[84]) & (g154) & (g122) & (!g1007) & (g1205) & (g999)) + ((!sk[84]) & (g154) & (g122) & (g1007) & (!g1205) & (!g999)) + ((!sk[84]) & (g154) & (g122) & (g1007) & (!g1205) & (g999)) + ((!sk[84]) & (g154) & (g122) & (g1007) & (g1205) & (!g999)) + ((!sk[84]) & (g154) & (g122) & (g1007) & (g1205) & (g999)) + ((sk[84]) & (!g154) & (!g122) & (g1007) & (!g1205) & (!g999)) + ((sk[84]) & (!g154) & (!g122) & (g1007) & (g1205) & (!g999)) + ((sk[84]) & (!g154) & (g122) & (g1007) & (g1205) & (!g999)) + ((sk[84]) & (g154) & (!g122) & (!g1007) & (!g1205) & (!g999)) + ((sk[84]) & (g154) & (!g122) & (!g1007) & (g1205) & (!g999)) + ((sk[84]) & (g154) & (!g122) & (g1007) & (!g1205) & (!g999)) + ((sk[84]) & (g154) & (!g122) & (g1007) & (g1205) & (!g999)) + ((sk[84]) & (g154) & (g122) & (!g1007) & (g1205) & (!g999)) + ((sk[84]) & (g154) & (g122) & (g1007) & (g1205) & (!g999)));
	assign g1207 = (((g915) & (g959) & (g1189) & (g1192) & (g1202) & (g1206)));
	assign g1208 = (((g722) & (!sk[86]) & (!g203)) + ((g722) & (!sk[86]) & (g203)) + ((g722) & (sk[86]) & (g203)));
	assign g1209 = (((!sk[87]) & (!i_8_) & (!g73) & (g551) & (!g495)) + ((!sk[87]) & (!i_8_) & (!g73) & (g551) & (g495)) + ((!sk[87]) & (!i_8_) & (g73) & (g551) & (!g495)) + ((!sk[87]) & (!i_8_) & (g73) & (g551) & (g495)) + ((!sk[87]) & (i_8_) & (!g73) & (g551) & (!g495)) + ((!sk[87]) & (i_8_) & (!g73) & (g551) & (g495)) + ((!sk[87]) & (i_8_) & (g73) & (g551) & (!g495)) + ((!sk[87]) & (i_8_) & (g73) & (g551) & (g495)) + ((sk[87]) & (i_8_) & (g73) & (!g551) & (!g495)) + ((sk[87]) & (i_8_) & (g73) & (!g551) & (g495)) + ((sk[87]) & (i_8_) & (g73) & (g551) & (g495)));
	assign g1210 = (((!g78) & (!sk[88]) & (!g122) & (g278) & (!g551)) + ((!g78) & (!sk[88]) & (!g122) & (g278) & (g551)) + ((!g78) & (!sk[88]) & (g122) & (g278) & (!g551)) + ((!g78) & (!sk[88]) & (g122) & (g278) & (g551)) + ((!g78) & (sk[88]) & (g122) & (!g278) & (!g551)) + ((!g78) & (sk[88]) & (g122) & (!g278) & (g551)) + ((!g78) & (sk[88]) & (g122) & (g278) & (!g551)) + ((!g78) & (sk[88]) & (g122) & (g278) & (g551)) + ((g78) & (!sk[88]) & (!g122) & (g278) & (!g551)) + ((g78) & (!sk[88]) & (!g122) & (g278) & (g551)) + ((g78) & (!sk[88]) & (g122) & (g278) & (!g551)) + ((g78) & (!sk[88]) & (g122) & (g278) & (g551)) + ((g78) & (sk[88]) & (g122) & (!g278) & (!g551)) + ((g78) & (sk[88]) & (g122) & (g278) & (!g551)) + ((g78) & (sk[88]) & (g122) & (g278) & (g551)));
	assign g1211 = (((!sk[89]) & (!g164) & (!g154) & (g333) & (!g343)) + ((!sk[89]) & (!g164) & (!g154) & (g333) & (g343)) + ((!sk[89]) & (!g164) & (g154) & (g333) & (!g343)) + ((!sk[89]) & (!g164) & (g154) & (g333) & (g343)) + ((!sk[89]) & (g164) & (!g154) & (g333) & (!g343)) + ((!sk[89]) & (g164) & (!g154) & (g333) & (g343)) + ((!sk[89]) & (g164) & (g154) & (g333) & (!g343)) + ((!sk[89]) & (g164) & (g154) & (g333) & (g343)) + ((sk[89]) & (!g164) & (!g154) & (!g333) & (g343)) + ((sk[89]) & (!g164) & (g154) & (!g333) & (!g343)) + ((sk[89]) & (!g164) & (g154) & (!g333) & (g343)) + ((sk[89]) & (!g164) & (g154) & (g333) & (!g343)) + ((sk[89]) & (!g164) & (g154) & (g333) & (g343)) + ((sk[89]) & (g164) & (!g154) & (!g333) & (g343)) + ((sk[89]) & (g164) & (g154) & (!g333) & (g343)) + ((sk[89]) & (g164) & (g154) & (g333) & (g343)));
	assign g1212 = (((!sk[90]) & (!g21) & (!g25) & (g125) & (!g278)) + ((!sk[90]) & (!g21) & (!g25) & (g125) & (g278)) + ((!sk[90]) & (!g21) & (g25) & (g125) & (!g278)) + ((!sk[90]) & (!g21) & (g25) & (g125) & (g278)) + ((!sk[90]) & (g21) & (!g25) & (g125) & (!g278)) + ((!sk[90]) & (g21) & (!g25) & (g125) & (g278)) + ((!sk[90]) & (g21) & (g25) & (g125) & (!g278)) + ((!sk[90]) & (g21) & (g25) & (g125) & (g278)) + ((sk[90]) & (!g21) & (!g25) & (g125) & (!g278)) + ((sk[90]) & (!g21) & (!g25) & (g125) & (g278)) + ((sk[90]) & (!g21) & (g25) & (g125) & (g278)) + ((sk[90]) & (g21) & (!g25) & (g125) & (!g278)) + ((sk[90]) & (g21) & (!g25) & (g125) & (g278)) + ((sk[90]) & (g21) & (g25) & (g125) & (!g278)) + ((sk[90]) & (g21) & (g25) & (g125) & (g278)));
	assign g1213 = (((!g154) & (!g105) & (!g521) & (!g625) & (sk[91]) & (!g626)) + ((!g154) & (!g105) & (g521) & (!g625) & (!sk[91]) & (g626)) + ((!g154) & (!g105) & (g521) & (g625) & (!sk[91]) & (!g626)) + ((!g154) & (!g105) & (g521) & (g625) & (!sk[91]) & (g626)) + ((!g154) & (g105) & (!g521) & (!g625) & (!sk[91]) & (!g626)) + ((!g154) & (g105) & (!g521) & (!g625) & (!sk[91]) & (g626)) + ((!g154) & (g105) & (!g521) & (!g625) & (sk[91]) & (!g626)) + ((!g154) & (g105) & (!g521) & (g625) & (!sk[91]) & (!g626)) + ((!g154) & (g105) & (!g521) & (g625) & (!sk[91]) & (g626)) + ((!g154) & (g105) & (g521) & (!g625) & (!sk[91]) & (!g626)) + ((!g154) & (g105) & (g521) & (!g625) & (!sk[91]) & (g626)) + ((!g154) & (g105) & (g521) & (g625) & (!sk[91]) & (!g626)) + ((!g154) & (g105) & (g521) & (g625) & (!sk[91]) & (g626)) + ((g154) & (!g105) & (!g521) & (!g625) & (sk[91]) & (!g626)) + ((g154) & (!g105) & (!g521) & (!g625) & (sk[91]) & (g626)) + ((g154) & (!g105) & (!g521) & (g625) & (sk[91]) & (!g626)) + ((g154) & (!g105) & (!g521) & (g625) & (sk[91]) & (g626)) + ((g154) & (!g105) & (g521) & (!g625) & (!sk[91]) & (g626)) + ((g154) & (!g105) & (g521) & (g625) & (!sk[91]) & (!g626)) + ((g154) & (!g105) & (g521) & (g625) & (!sk[91]) & (g626)) + ((g154) & (g105) & (!g521) & (!g625) & (!sk[91]) & (!g626)) + ((g154) & (g105) & (!g521) & (!g625) & (!sk[91]) & (g626)) + ((g154) & (g105) & (!g521) & (!g625) & (sk[91]) & (!g626)) + ((g154) & (g105) & (!g521) & (!g625) & (sk[91]) & (g626)) + ((g154) & (g105) & (!g521) & (g625) & (!sk[91]) & (!g626)) + ((g154) & (g105) & (!g521) & (g625) & (!sk[91]) & (g626)) + ((g154) & (g105) & (!g521) & (g625) & (sk[91]) & (!g626)) + ((g154) & (g105) & (!g521) & (g625) & (sk[91]) & (g626)) + ((g154) & (g105) & (g521) & (!g625) & (!sk[91]) & (!g626)) + ((g154) & (g105) & (g521) & (!g625) & (!sk[91]) & (g626)) + ((g154) & (g105) & (g521) & (!g625) & (sk[91]) & (!g626)) + ((g154) & (g105) & (g521) & (!g625) & (sk[91]) & (g626)) + ((g154) & (g105) & (g521) & (g625) & (!sk[91]) & (!g626)) + ((g154) & (g105) & (g521) & (g625) & (!sk[91]) & (g626)) + ((g154) & (g105) & (g521) & (g625) & (sk[91]) & (!g626)) + ((g154) & (g105) & (g521) & (g625) & (sk[91]) & (g626)));
	assign g1214 = (((!g1209) & (!g1210) & (g1211) & (!g1212) & (!sk[92]) & (g1213)) + ((!g1209) & (!g1210) & (g1211) & (!g1212) & (sk[92]) & (g1213)) + ((!g1209) & (!g1210) & (g1211) & (g1212) & (!sk[92]) & (!g1213)) + ((!g1209) & (!g1210) & (g1211) & (g1212) & (!sk[92]) & (g1213)) + ((!g1209) & (g1210) & (!g1211) & (!g1212) & (!sk[92]) & (!g1213)) + ((!g1209) & (g1210) & (!g1211) & (!g1212) & (!sk[92]) & (g1213)) + ((!g1209) & (g1210) & (!g1211) & (g1212) & (!sk[92]) & (!g1213)) + ((!g1209) & (g1210) & (!g1211) & (g1212) & (!sk[92]) & (g1213)) + ((!g1209) & (g1210) & (g1211) & (!g1212) & (!sk[92]) & (!g1213)) + ((!g1209) & (g1210) & (g1211) & (!g1212) & (!sk[92]) & (g1213)) + ((!g1209) & (g1210) & (g1211) & (g1212) & (!sk[92]) & (!g1213)) + ((!g1209) & (g1210) & (g1211) & (g1212) & (!sk[92]) & (g1213)) + ((g1209) & (!g1210) & (g1211) & (!g1212) & (!sk[92]) & (g1213)) + ((g1209) & (!g1210) & (g1211) & (g1212) & (!sk[92]) & (!g1213)) + ((g1209) & (!g1210) & (g1211) & (g1212) & (!sk[92]) & (g1213)) + ((g1209) & (g1210) & (!g1211) & (!g1212) & (!sk[92]) & (!g1213)) + ((g1209) & (g1210) & (!g1211) & (!g1212) & (!sk[92]) & (g1213)) + ((g1209) & (g1210) & (!g1211) & (g1212) & (!sk[92]) & (!g1213)) + ((g1209) & (g1210) & (!g1211) & (g1212) & (!sk[92]) & (g1213)) + ((g1209) & (g1210) & (g1211) & (!g1212) & (!sk[92]) & (!g1213)) + ((g1209) & (g1210) & (g1211) & (!g1212) & (!sk[92]) & (g1213)) + ((g1209) & (g1210) & (g1211) & (g1212) & (!sk[92]) & (!g1213)) + ((g1209) & (g1210) & (g1211) & (g1212) & (!sk[92]) & (g1213)));
	assign g1215 = (((!i_8_) & (!i_6_) & (!sk[93]) & (i_7_) & (!g428) & (g394)) + ((!i_8_) & (!i_6_) & (!sk[93]) & (i_7_) & (g428) & (!g394)) + ((!i_8_) & (!i_6_) & (!sk[93]) & (i_7_) & (g428) & (g394)) + ((!i_8_) & (i_6_) & (!sk[93]) & (!i_7_) & (!g428) & (!g394)) + ((!i_8_) & (i_6_) & (!sk[93]) & (!i_7_) & (!g428) & (g394)) + ((!i_8_) & (i_6_) & (!sk[93]) & (!i_7_) & (g428) & (!g394)) + ((!i_8_) & (i_6_) & (!sk[93]) & (!i_7_) & (g428) & (g394)) + ((!i_8_) & (i_6_) & (!sk[93]) & (i_7_) & (!g428) & (!g394)) + ((!i_8_) & (i_6_) & (!sk[93]) & (i_7_) & (!g428) & (g394)) + ((!i_8_) & (i_6_) & (!sk[93]) & (i_7_) & (g428) & (!g394)) + ((!i_8_) & (i_6_) & (!sk[93]) & (i_7_) & (g428) & (g394)) + ((i_8_) & (!i_6_) & (!sk[93]) & (i_7_) & (!g428) & (g394)) + ((i_8_) & (!i_6_) & (!sk[93]) & (i_7_) & (g428) & (!g394)) + ((i_8_) & (!i_6_) & (!sk[93]) & (i_7_) & (g428) & (g394)) + ((i_8_) & (!i_6_) & (sk[93]) & (i_7_) & (!g428) & (g394)) + ((i_8_) & (i_6_) & (!sk[93]) & (!i_7_) & (!g428) & (!g394)) + ((i_8_) & (i_6_) & (!sk[93]) & (!i_7_) & (!g428) & (g394)) + ((i_8_) & (i_6_) & (!sk[93]) & (!i_7_) & (g428) & (!g394)) + ((i_8_) & (i_6_) & (!sk[93]) & (!i_7_) & (g428) & (g394)) + ((i_8_) & (i_6_) & (!sk[93]) & (i_7_) & (!g428) & (!g394)) + ((i_8_) & (i_6_) & (!sk[93]) & (i_7_) & (!g428) & (g394)) + ((i_8_) & (i_6_) & (!sk[93]) & (i_7_) & (g428) & (!g394)) + ((i_8_) & (i_6_) & (!sk[93]) & (i_7_) & (g428) & (g394)) + ((i_8_) & (i_6_) & (sk[93]) & (!i_7_) & (!g428) & (g394)) + ((i_8_) & (i_6_) & (sk[93]) & (i_7_) & (!g428) & (g394)));
	assign g1216 = (((!sk[94]) & (!i_8_) & (!g25) & (g73) & (!g278) & (g1215)) + ((!sk[94]) & (!i_8_) & (!g25) & (g73) & (g278) & (!g1215)) + ((!sk[94]) & (!i_8_) & (!g25) & (g73) & (g278) & (g1215)) + ((!sk[94]) & (!i_8_) & (g25) & (!g73) & (!g278) & (!g1215)) + ((!sk[94]) & (!i_8_) & (g25) & (!g73) & (!g278) & (g1215)) + ((!sk[94]) & (!i_8_) & (g25) & (!g73) & (g278) & (!g1215)) + ((!sk[94]) & (!i_8_) & (g25) & (!g73) & (g278) & (g1215)) + ((!sk[94]) & (!i_8_) & (g25) & (g73) & (!g278) & (!g1215)) + ((!sk[94]) & (!i_8_) & (g25) & (g73) & (!g278) & (g1215)) + ((!sk[94]) & (!i_8_) & (g25) & (g73) & (g278) & (!g1215)) + ((!sk[94]) & (!i_8_) & (g25) & (g73) & (g278) & (g1215)) + ((!sk[94]) & (i_8_) & (!g25) & (g73) & (!g278) & (g1215)) + ((!sk[94]) & (i_8_) & (!g25) & (g73) & (g278) & (!g1215)) + ((!sk[94]) & (i_8_) & (!g25) & (g73) & (g278) & (g1215)) + ((!sk[94]) & (i_8_) & (g25) & (!g73) & (!g278) & (!g1215)) + ((!sk[94]) & (i_8_) & (g25) & (!g73) & (!g278) & (g1215)) + ((!sk[94]) & (i_8_) & (g25) & (!g73) & (g278) & (!g1215)) + ((!sk[94]) & (i_8_) & (g25) & (!g73) & (g278) & (g1215)) + ((!sk[94]) & (i_8_) & (g25) & (g73) & (!g278) & (!g1215)) + ((!sk[94]) & (i_8_) & (g25) & (g73) & (!g278) & (g1215)) + ((!sk[94]) & (i_8_) & (g25) & (g73) & (g278) & (!g1215)) + ((!sk[94]) & (i_8_) & (g25) & (g73) & (g278) & (g1215)) + ((sk[94]) & (!i_8_) & (!g25) & (!g73) & (!g278) & (!g1215)) + ((sk[94]) & (!i_8_) & (!g25) & (!g73) & (g278) & (!g1215)) + ((sk[94]) & (!i_8_) & (!g25) & (g73) & (!g278) & (!g1215)) + ((sk[94]) & (!i_8_) & (!g25) & (g73) & (g278) & (!g1215)) + ((sk[94]) & (!i_8_) & (g25) & (!g73) & (!g278) & (!g1215)) + ((sk[94]) & (!i_8_) & (g25) & (!g73) & (g278) & (!g1215)) + ((sk[94]) & (!i_8_) & (g25) & (g73) & (!g278) & (!g1215)) + ((sk[94]) & (!i_8_) & (g25) & (g73) & (g278) & (!g1215)) + ((sk[94]) & (i_8_) & (!g25) & (!g73) & (!g278) & (!g1215)) + ((sk[94]) & (i_8_) & (!g25) & (!g73) & (g278) & (!g1215)) + ((sk[94]) & (i_8_) & (g25) & (!g73) & (!g278) & (!g1215)) + ((sk[94]) & (i_8_) & (g25) & (!g73) & (g278) & (!g1215)) + ((sk[94]) & (i_8_) & (g25) & (g73) & (!g278) & (!g1215)));
	assign g1217 = (((!g222) & (!g207) & (!g776) & (sk[95]) & (!g783) & (g1216)) + ((!g222) & (!g207) & (g776) & (!sk[95]) & (!g783) & (g1216)) + ((!g222) & (!g207) & (g776) & (!sk[95]) & (g783) & (!g1216)) + ((!g222) & (!g207) & (g776) & (!sk[95]) & (g783) & (g1216)) + ((!g222) & (g207) & (!g776) & (!sk[95]) & (!g783) & (!g1216)) + ((!g222) & (g207) & (!g776) & (!sk[95]) & (!g783) & (g1216)) + ((!g222) & (g207) & (!g776) & (!sk[95]) & (g783) & (!g1216)) + ((!g222) & (g207) & (!g776) & (!sk[95]) & (g783) & (g1216)) + ((!g222) & (g207) & (g776) & (!sk[95]) & (!g783) & (!g1216)) + ((!g222) & (g207) & (g776) & (!sk[95]) & (!g783) & (g1216)) + ((!g222) & (g207) & (g776) & (!sk[95]) & (g783) & (!g1216)) + ((!g222) & (g207) & (g776) & (!sk[95]) & (g783) & (g1216)) + ((g222) & (!g207) & (g776) & (!sk[95]) & (!g783) & (g1216)) + ((g222) & (!g207) & (g776) & (!sk[95]) & (g783) & (!g1216)) + ((g222) & (!g207) & (g776) & (!sk[95]) & (g783) & (g1216)) + ((g222) & (g207) & (!g776) & (!sk[95]) & (!g783) & (!g1216)) + ((g222) & (g207) & (!g776) & (!sk[95]) & (!g783) & (g1216)) + ((g222) & (g207) & (!g776) & (!sk[95]) & (g783) & (!g1216)) + ((g222) & (g207) & (!g776) & (!sk[95]) & (g783) & (g1216)) + ((g222) & (g207) & (g776) & (!sk[95]) & (!g783) & (!g1216)) + ((g222) & (g207) & (g776) & (!sk[95]) & (!g783) & (g1216)) + ((g222) & (g207) & (g776) & (!sk[95]) & (g783) & (!g1216)) + ((g222) & (g207) & (g776) & (!sk[95]) & (g783) & (g1216)));
	assign g1218 = (((!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (!g428) & (!g75)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g428) & (!g75)) + ((!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g428) & (!g75)) + ((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g428) & (!g75)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g428) & (!g75)) + ((i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (!g428) & (!g75)) + ((i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (!g428) & (!g75)) + ((i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (!g428) & (!g75)) + ((i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g428) & (!g75)) + ((i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g428) & (!g75)) + ((i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g428) & (!g75)));
	assign g1219 = (((!g125) & (!g164) & (!sk[97]) & (g551) & (!g626)) + ((!g125) & (!g164) & (!sk[97]) & (g551) & (g626)) + ((!g125) & (g164) & (!sk[97]) & (g551) & (!g626)) + ((!g125) & (g164) & (!sk[97]) & (g551) & (g626)) + ((!g125) & (g164) & (sk[97]) & (!g551) & (g626)) + ((!g125) & (g164) & (sk[97]) & (g551) & (g626)) + ((g125) & (!g164) & (!sk[97]) & (g551) & (!g626)) + ((g125) & (!g164) & (!sk[97]) & (g551) & (g626)) + ((g125) & (!g164) & (sk[97]) & (!g551) & (!g626)) + ((g125) & (!g164) & (sk[97]) & (!g551) & (g626)) + ((g125) & (g164) & (!sk[97]) & (g551) & (!g626)) + ((g125) & (g164) & (!sk[97]) & (g551) & (g626)) + ((g125) & (g164) & (sk[97]) & (!g551) & (!g626)) + ((g125) & (g164) & (sk[97]) & (!g551) & (g626)) + ((g125) & (g164) & (sk[97]) & (g551) & (g626)));
	assign g1220 = (((!g161) & (!g164) & (!g343) & (!g452) & (!g521) & (!g1219)) + ((!g161) & (!g164) & (!g343) & (!g452) & (g521) & (!g1219)) + ((!g161) & (!g164) & (g343) & (!g452) & (!g521) & (!g1219)) + ((!g161) & (!g164) & (g343) & (!g452) & (g521) & (!g1219)) + ((!g161) & (g164) & (!g343) & (!g452) & (!g521) & (!g1219)) + ((!g161) & (g164) & (g343) & (!g452) & (!g521) & (!g1219)) + ((g161) & (!g164) & (g343) & (!g452) & (!g521) & (!g1219)) + ((g161) & (!g164) & (g343) & (!g452) & (g521) & (!g1219)) + ((g161) & (g164) & (g343) & (!g452) & (!g521) & (!g1219)));
	assign g1221 = (((!g164) & (!g154) & (!sk[99]) & (g865) & (!g978) & (g1047)) + ((!g164) & (!g154) & (!sk[99]) & (g865) & (g978) & (!g1047)) + ((!g164) & (!g154) & (!sk[99]) & (g865) & (g978) & (g1047)) + ((!g164) & (!g154) & (sk[99]) & (!g865) & (!g978) & (!g1047)) + ((!g164) & (!g154) & (sk[99]) & (!g865) & (g978) & (!g1047)) + ((!g164) & (g154) & (!sk[99]) & (!g865) & (!g978) & (!g1047)) + ((!g164) & (g154) & (!sk[99]) & (!g865) & (!g978) & (g1047)) + ((!g164) & (g154) & (!sk[99]) & (!g865) & (g978) & (!g1047)) + ((!g164) & (g154) & (!sk[99]) & (!g865) & (g978) & (g1047)) + ((!g164) & (g154) & (!sk[99]) & (g865) & (!g978) & (!g1047)) + ((!g164) & (g154) & (!sk[99]) & (g865) & (!g978) & (g1047)) + ((!g164) & (g154) & (!sk[99]) & (g865) & (g978) & (!g1047)) + ((!g164) & (g154) & (!sk[99]) & (g865) & (g978) & (g1047)) + ((!g164) & (g154) & (sk[99]) & (!g865) & (!g978) & (!g1047)) + ((!g164) & (g154) & (sk[99]) & (!g865) & (g978) & (!g1047)) + ((!g164) & (g154) & (sk[99]) & (g865) & (!g978) & (!g1047)) + ((!g164) & (g154) & (sk[99]) & (g865) & (g978) & (!g1047)) + ((g164) & (!g154) & (!sk[99]) & (g865) & (!g978) & (g1047)) + ((g164) & (!g154) & (!sk[99]) & (g865) & (g978) & (!g1047)) + ((g164) & (!g154) & (!sk[99]) & (g865) & (g978) & (g1047)) + ((g164) & (!g154) & (sk[99]) & (!g865) & (g978) & (!g1047)) + ((g164) & (g154) & (!sk[99]) & (!g865) & (!g978) & (!g1047)) + ((g164) & (g154) & (!sk[99]) & (!g865) & (!g978) & (g1047)) + ((g164) & (g154) & (!sk[99]) & (!g865) & (g978) & (!g1047)) + ((g164) & (g154) & (!sk[99]) & (!g865) & (g978) & (g1047)) + ((g164) & (g154) & (!sk[99]) & (g865) & (!g978) & (!g1047)) + ((g164) & (g154) & (!sk[99]) & (g865) & (!g978) & (g1047)) + ((g164) & (g154) & (!sk[99]) & (g865) & (g978) & (!g1047)) + ((g164) & (g154) & (!sk[99]) & (g865) & (g978) & (g1047)) + ((g164) & (g154) & (sk[99]) & (!g865) & (g978) & (!g1047)) + ((g164) & (g154) & (sk[99]) & (g865) & (g978) & (!g1047)));
	assign g1222 = (((!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (!g428) & (!g123)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g428) & (!g123)) + ((!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g428) & (!g123)) + ((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g428) & (!g123)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g428) & (!g123)) + ((i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (!g428) & (!g123)) + ((i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (!g428) & (!g123)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g428) & (!g123)) + ((i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g428) & (!g123)));
	assign g1223 = (((!g953) & (sk[101]) & (!g1222)) + ((g953) & (!sk[101]) & (!g1222)) + ((g953) & (!sk[101]) & (g1222)));
	assign g1224 = (((g1214) & (g1217) & (!g1218) & (g1220) & (g1221) & (g1223)));
	assign g1225 = (((!g3) & (!sk[103]) & (!g48) & (g119) & (!g460)) + ((!g3) & (!sk[103]) & (!g48) & (g119) & (g460)) + ((!g3) & (!sk[103]) & (g48) & (g119) & (!g460)) + ((!g3) & (!sk[103]) & (g48) & (g119) & (g460)) + ((!g3) & (sk[103]) & (!g48) & (!g119) & (!g460)) + ((!g3) & (sk[103]) & (!g48) & (!g119) & (g460)) + ((!g3) & (sk[103]) & (!g48) & (g119) & (!g460)) + ((!g3) & (sk[103]) & (!g48) & (g119) & (g460)) + ((g3) & (!sk[103]) & (!g48) & (g119) & (!g460)) + ((g3) & (!sk[103]) & (!g48) & (g119) & (g460)) + ((g3) & (!sk[103]) & (g48) & (g119) & (!g460)) + ((g3) & (!sk[103]) & (g48) & (g119) & (g460)) + ((g3) & (sk[103]) & (!g48) & (!g119) & (!g460)) + ((g3) & (sk[103]) & (!g48) & (!g119) & (g460)) + ((g3) & (sk[103]) & (!g48) & (g119) & (g460)));
	assign g1226 = (((!i_8_) & (!sk[104]) & (!i_3_) & (i_5_) & (!g10) & (g71)) + ((!i_8_) & (!sk[104]) & (!i_3_) & (i_5_) & (g10) & (!g71)) + ((!i_8_) & (!sk[104]) & (!i_3_) & (i_5_) & (g10) & (g71)) + ((!i_8_) & (!sk[104]) & (i_3_) & (!i_5_) & (!g10) & (!g71)) + ((!i_8_) & (!sk[104]) & (i_3_) & (!i_5_) & (!g10) & (g71)) + ((!i_8_) & (!sk[104]) & (i_3_) & (!i_5_) & (g10) & (!g71)) + ((!i_8_) & (!sk[104]) & (i_3_) & (!i_5_) & (g10) & (g71)) + ((!i_8_) & (!sk[104]) & (i_3_) & (i_5_) & (!g10) & (!g71)) + ((!i_8_) & (!sk[104]) & (i_3_) & (i_5_) & (!g10) & (g71)) + ((!i_8_) & (!sk[104]) & (i_3_) & (i_5_) & (g10) & (!g71)) + ((!i_8_) & (!sk[104]) & (i_3_) & (i_5_) & (g10) & (g71)) + ((i_8_) & (!sk[104]) & (!i_3_) & (i_5_) & (!g10) & (g71)) + ((i_8_) & (!sk[104]) & (!i_3_) & (i_5_) & (g10) & (!g71)) + ((i_8_) & (!sk[104]) & (!i_3_) & (i_5_) & (g10) & (g71)) + ((i_8_) & (!sk[104]) & (i_3_) & (!i_5_) & (!g10) & (!g71)) + ((i_8_) & (!sk[104]) & (i_3_) & (!i_5_) & (!g10) & (g71)) + ((i_8_) & (!sk[104]) & (i_3_) & (!i_5_) & (g10) & (!g71)) + ((i_8_) & (!sk[104]) & (i_3_) & (!i_5_) & (g10) & (g71)) + ((i_8_) & (!sk[104]) & (i_3_) & (i_5_) & (!g10) & (!g71)) + ((i_8_) & (!sk[104]) & (i_3_) & (i_5_) & (!g10) & (g71)) + ((i_8_) & (!sk[104]) & (i_3_) & (i_5_) & (g10) & (!g71)) + ((i_8_) & (!sk[104]) & (i_3_) & (i_5_) & (g10) & (g71)) + ((i_8_) & (sk[104]) & (!i_3_) & (i_5_) & (g10) & (g71)));
	assign g1227 = (((!g3) & (!g75) & (!g460) & (sk[105]) & (!g927) & (g1226)) + ((!g3) & (!g75) & (!g460) & (sk[105]) & (g927) & (g1226)) + ((!g3) & (!g75) & (g460) & (!sk[105]) & (!g927) & (g1226)) + ((!g3) & (!g75) & (g460) & (!sk[105]) & (g927) & (!g1226)) + ((!g3) & (!g75) & (g460) & (!sk[105]) & (g927) & (g1226)) + ((!g3) & (!g75) & (g460) & (sk[105]) & (!g927) & (g1226)) + ((!g3) & (!g75) & (g460) & (sk[105]) & (g927) & (g1226)) + ((!g3) & (g75) & (!g460) & (!sk[105]) & (!g927) & (!g1226)) + ((!g3) & (g75) & (!g460) & (!sk[105]) & (!g927) & (g1226)) + ((!g3) & (g75) & (!g460) & (!sk[105]) & (g927) & (!g1226)) + ((!g3) & (g75) & (!g460) & (!sk[105]) & (g927) & (g1226)) + ((!g3) & (g75) & (!g460) & (sk[105]) & (g927) & (g1226)) + ((!g3) & (g75) & (g460) & (!sk[105]) & (!g927) & (!g1226)) + ((!g3) & (g75) & (g460) & (!sk[105]) & (!g927) & (g1226)) + ((!g3) & (g75) & (g460) & (!sk[105]) & (g927) & (!g1226)) + ((!g3) & (g75) & (g460) & (!sk[105]) & (g927) & (g1226)) + ((!g3) & (g75) & (g460) & (sk[105]) & (g927) & (g1226)) + ((g3) & (!g75) & (!g460) & (sk[105]) & (!g927) & (g1226)) + ((g3) & (!g75) & (!g460) & (sk[105]) & (g927) & (g1226)) + ((g3) & (!g75) & (g460) & (!sk[105]) & (!g927) & (g1226)) + ((g3) & (!g75) & (g460) & (!sk[105]) & (g927) & (!g1226)) + ((g3) & (!g75) & (g460) & (!sk[105]) & (g927) & (g1226)) + ((g3) & (!g75) & (g460) & (sk[105]) & (!g927) & (g1226)) + ((g3) & (!g75) & (g460) & (sk[105]) & (g927) & (g1226)) + ((g3) & (g75) & (!g460) & (!sk[105]) & (!g927) & (!g1226)) + ((g3) & (g75) & (!g460) & (!sk[105]) & (!g927) & (g1226)) + ((g3) & (g75) & (!g460) & (!sk[105]) & (g927) & (!g1226)) + ((g3) & (g75) & (!g460) & (!sk[105]) & (g927) & (g1226)) + ((g3) & (g75) & (!g460) & (sk[105]) & (!g927) & (g1226)) + ((g3) & (g75) & (!g460) & (sk[105]) & (g927) & (g1226)) + ((g3) & (g75) & (g460) & (!sk[105]) & (!g927) & (!g1226)) + ((g3) & (g75) & (g460) & (!sk[105]) & (!g927) & (g1226)) + ((g3) & (g75) & (g460) & (!sk[105]) & (g927) & (!g1226)) + ((g3) & (g75) & (g460) & (!sk[105]) & (g927) & (g1226)) + ((g3) & (g75) & (g460) & (sk[105]) & (g927) & (g1226)));
	assign g1228 = (((!g468) & (!g608) & (!g927) & (sk[106]) & (!g1225) & (g1227)) + ((!g468) & (!g608) & (!g927) & (sk[106]) & (g1225) & (g1227)) + ((!g468) & (!g608) & (g927) & (!sk[106]) & (!g1225) & (g1227)) + ((!g468) & (!g608) & (g927) & (!sk[106]) & (g1225) & (!g1227)) + ((!g468) & (!g608) & (g927) & (!sk[106]) & (g1225) & (g1227)) + ((!g468) & (!g608) & (g927) & (sk[106]) & (!g1225) & (g1227)) + ((!g468) & (!g608) & (g927) & (sk[106]) & (g1225) & (g1227)) + ((!g468) & (g608) & (!g927) & (!sk[106]) & (!g1225) & (!g1227)) + ((!g468) & (g608) & (!g927) & (!sk[106]) & (!g1225) & (g1227)) + ((!g468) & (g608) & (!g927) & (!sk[106]) & (g1225) & (!g1227)) + ((!g468) & (g608) & (!g927) & (!sk[106]) & (g1225) & (g1227)) + ((!g468) & (g608) & (!g927) & (sk[106]) & (!g1225) & (g1227)) + ((!g468) & (g608) & (g927) & (!sk[106]) & (!g1225) & (!g1227)) + ((!g468) & (g608) & (g927) & (!sk[106]) & (!g1225) & (g1227)) + ((!g468) & (g608) & (g927) & (!sk[106]) & (g1225) & (!g1227)) + ((!g468) & (g608) & (g927) & (!sk[106]) & (g1225) & (g1227)) + ((!g468) & (g608) & (g927) & (sk[106]) & (!g1225) & (g1227)) + ((!g468) & (g608) & (g927) & (sk[106]) & (g1225) & (g1227)) + ((g468) & (!g608) & (!g927) & (sk[106]) & (!g1225) & (g1227)) + ((g468) & (!g608) & (!g927) & (sk[106]) & (g1225) & (g1227)) + ((g468) & (!g608) & (g927) & (!sk[106]) & (!g1225) & (g1227)) + ((g468) & (!g608) & (g927) & (!sk[106]) & (g1225) & (!g1227)) + ((g468) & (!g608) & (g927) & (!sk[106]) & (g1225) & (g1227)) + ((g468) & (!g608) & (g927) & (sk[106]) & (!g1225) & (g1227)) + ((g468) & (!g608) & (g927) & (sk[106]) & (g1225) & (g1227)) + ((g468) & (g608) & (!g927) & (!sk[106]) & (!g1225) & (!g1227)) + ((g468) & (g608) & (!g927) & (!sk[106]) & (!g1225) & (g1227)) + ((g468) & (g608) & (!g927) & (!sk[106]) & (g1225) & (!g1227)) + ((g468) & (g608) & (!g927) & (!sk[106]) & (g1225) & (g1227)) + ((g468) & (g608) & (!g927) & (sk[106]) & (!g1225) & (g1227)) + ((g468) & (g608) & (!g927) & (sk[106]) & (g1225) & (g1227)) + ((g468) & (g608) & (g927) & (!sk[106]) & (!g1225) & (!g1227)) + ((g468) & (g608) & (g927) & (!sk[106]) & (!g1225) & (g1227)) + ((g468) & (g608) & (g927) & (!sk[106]) & (g1225) & (!g1227)) + ((g468) & (g608) & (g927) & (!sk[106]) & (g1225) & (g1227)) + ((g468) & (g608) & (g927) & (sk[106]) & (!g1225) & (g1227)) + ((g468) & (g608) & (g927) & (sk[106]) & (g1225) & (g1227)));
	assign g1229 = (((!g69) & (!g113) & (!sk[107]) & (g105) & (!g482)) + ((!g69) & (!g113) & (!sk[107]) & (g105) & (g482)) + ((!g69) & (!g113) & (sk[107]) & (!g105) & (g482)) + ((!g69) & (g113) & (!sk[107]) & (g105) & (!g482)) + ((!g69) & (g113) & (!sk[107]) & (g105) & (g482)) + ((g69) & (!g113) & (!sk[107]) & (g105) & (!g482)) + ((g69) & (!g113) & (!sk[107]) & (g105) & (g482)) + ((g69) & (!g113) & (sk[107]) & (!g105) & (g482)) + ((g69) & (g113) & (!sk[107]) & (g105) & (!g482)) + ((g69) & (g113) & (!sk[107]) & (g105) & (g482)) + ((g69) & (g113) & (sk[107]) & (!g105) & (g482)));
	assign g1230 = (((!g355) & (!g126) & (g122) & (!g182) & (!g460) & (!g552)) + ((!g355) & (!g126) & (g122) & (!g182) & (!g460) & (g552)) + ((!g355) & (!g126) & (g122) & (!g182) & (g460) & (!g552)) + ((!g355) & (!g126) & (g122) & (g182) & (!g460) & (!g552)) + ((!g355) & (!g126) & (g122) & (g182) & (!g460) & (g552)) + ((!g355) & (!g126) & (g122) & (g182) & (g460) & (!g552)) + ((!g355) & (!g126) & (g122) & (g182) & (g460) & (g552)) + ((!g355) & (g126) & (g122) & (!g182) & (!g460) & (!g552)) + ((!g355) & (g126) & (g122) & (!g182) & (g460) & (!g552)) + ((!g355) & (g126) & (g122) & (g182) & (!g460) & (!g552)) + ((!g355) & (g126) & (g122) & (g182) & (!g460) & (g552)) + ((!g355) & (g126) & (g122) & (g182) & (g460) & (!g552)) + ((!g355) & (g126) & (g122) & (g182) & (g460) & (g552)) + ((g355) & (!g126) & (g122) & (!g182) & (!g460) & (!g552)) + ((g355) & (!g126) & (g122) & (!g182) & (!g460) & (g552)) + ((g355) & (!g126) & (g122) & (!g182) & (g460) & (!g552)) + ((g355) & (!g126) & (g122) & (!g182) & (g460) & (g552)) + ((g355) & (!g126) & (g122) & (g182) & (!g460) & (!g552)) + ((g355) & (!g126) & (g122) & (g182) & (!g460) & (g552)) + ((g355) & (!g126) & (g122) & (g182) & (g460) & (!g552)) + ((g355) & (!g126) & (g122) & (g182) & (g460) & (g552)) + ((g355) & (g126) & (g122) & (!g182) & (!g460) & (!g552)) + ((g355) & (g126) & (g122) & (!g182) & (g460) & (!g552)) + ((g355) & (g126) & (g122) & (g182) & (!g460) & (!g552)) + ((g355) & (g126) & (g122) & (g182) & (!g460) & (g552)) + ((g355) & (g126) & (g122) & (g182) & (g460) & (!g552)) + ((g355) & (g126) & (g122) & (g182) & (g460) & (g552)));
	assign g1231 = (((!g75) & (!g282) & (!g270) & (!g585) & (sk[109]) & (!g1230)) + ((!g75) & (!g282) & (g270) & (!g585) & (!sk[109]) & (g1230)) + ((!g75) & (!g282) & (g270) & (g585) & (!sk[109]) & (!g1230)) + ((!g75) & (!g282) & (g270) & (g585) & (!sk[109]) & (g1230)) + ((!g75) & (g282) & (!g270) & (!g585) & (!sk[109]) & (!g1230)) + ((!g75) & (g282) & (!g270) & (!g585) & (!sk[109]) & (g1230)) + ((!g75) & (g282) & (!g270) & (g585) & (!sk[109]) & (!g1230)) + ((!g75) & (g282) & (!g270) & (g585) & (!sk[109]) & (g1230)) + ((!g75) & (g282) & (g270) & (!g585) & (!sk[109]) & (!g1230)) + ((!g75) & (g282) & (g270) & (!g585) & (!sk[109]) & (g1230)) + ((!g75) & (g282) & (g270) & (g585) & (!sk[109]) & (!g1230)) + ((!g75) & (g282) & (g270) & (g585) & (!sk[109]) & (g1230)) + ((g75) & (!g282) & (!g270) & (!g585) & (sk[109]) & (!g1230)) + ((g75) & (!g282) & (g270) & (!g585) & (!sk[109]) & (g1230)) + ((g75) & (!g282) & (g270) & (!g585) & (sk[109]) & (!g1230)) + ((g75) & (!g282) & (g270) & (g585) & (!sk[109]) & (!g1230)) + ((g75) & (!g282) & (g270) & (g585) & (!sk[109]) & (g1230)) + ((g75) & (g282) & (!g270) & (!g585) & (!sk[109]) & (!g1230)) + ((g75) & (g282) & (!g270) & (!g585) & (!sk[109]) & (g1230)) + ((g75) & (g282) & (!g270) & (!g585) & (sk[109]) & (!g1230)) + ((g75) & (g282) & (!g270) & (g585) & (!sk[109]) & (!g1230)) + ((g75) & (g282) & (!g270) & (g585) & (!sk[109]) & (g1230)) + ((g75) & (g282) & (g270) & (!g585) & (!sk[109]) & (!g1230)) + ((g75) & (g282) & (g270) & (!g585) & (!sk[109]) & (g1230)) + ((g75) & (g282) & (g270) & (!g585) & (sk[109]) & (!g1230)) + ((g75) & (g282) & (g270) & (g585) & (!sk[109]) & (!g1230)) + ((g75) & (g282) & (g270) & (g585) & (!sk[109]) & (g1230)));
	assign g1232 = (((!sk[110]) & (!g105) & (!g1229) & (g877) & (!g857) & (g1231)) + ((!sk[110]) & (!g105) & (!g1229) & (g877) & (g857) & (!g1231)) + ((!sk[110]) & (!g105) & (!g1229) & (g877) & (g857) & (g1231)) + ((!sk[110]) & (!g105) & (g1229) & (!g877) & (!g857) & (!g1231)) + ((!sk[110]) & (!g105) & (g1229) & (!g877) & (!g857) & (g1231)) + ((!sk[110]) & (!g105) & (g1229) & (!g877) & (g857) & (!g1231)) + ((!sk[110]) & (!g105) & (g1229) & (!g877) & (g857) & (g1231)) + ((!sk[110]) & (!g105) & (g1229) & (g877) & (!g857) & (!g1231)) + ((!sk[110]) & (!g105) & (g1229) & (g877) & (!g857) & (g1231)) + ((!sk[110]) & (!g105) & (g1229) & (g877) & (g857) & (!g1231)) + ((!sk[110]) & (!g105) & (g1229) & (g877) & (g857) & (g1231)) + ((!sk[110]) & (g105) & (!g1229) & (g877) & (!g857) & (g1231)) + ((!sk[110]) & (g105) & (!g1229) & (g877) & (g857) & (!g1231)) + ((!sk[110]) & (g105) & (!g1229) & (g877) & (g857) & (g1231)) + ((!sk[110]) & (g105) & (g1229) & (!g877) & (!g857) & (!g1231)) + ((!sk[110]) & (g105) & (g1229) & (!g877) & (!g857) & (g1231)) + ((!sk[110]) & (g105) & (g1229) & (!g877) & (g857) & (!g1231)) + ((!sk[110]) & (g105) & (g1229) & (!g877) & (g857) & (g1231)) + ((!sk[110]) & (g105) & (g1229) & (g877) & (!g857) & (!g1231)) + ((!sk[110]) & (g105) & (g1229) & (g877) & (!g857) & (g1231)) + ((!sk[110]) & (g105) & (g1229) & (g877) & (g857) & (!g1231)) + ((!sk[110]) & (g105) & (g1229) & (g877) & (g857) & (g1231)) + ((sk[110]) & (!g105) & (!g1229) & (!g877) & (!g857) & (g1231)) + ((sk[110]) & (g105) & (!g1229) & (!g877) & (!g857) & (g1231)) + ((sk[110]) & (g105) & (!g1229) & (!g877) & (g857) & (g1231)) + ((sk[110]) & (g105) & (!g1229) & (g877) & (!g857) & (g1231)) + ((sk[110]) & (g105) & (!g1229) & (g877) & (g857) & (g1231)));
	assign g1233 = (((!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (!g75) & (g112)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g75) & (g112)) + ((!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g75) & (g112)) + ((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g75) & (g112)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g75) & (g112)) + ((i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (!g75) & (g112)) + ((i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (!g75) & (g112)) + ((i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (!g75) & (g112)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g75) & (g112)) + ((i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g75) & (g112)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g75) & (g112)) + ((i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g75) & (g112)));
	assign g1234 = (((!g125) & (!g154) & (!g688) & (!g877) & (g929) & (!g1012)) + ((!g125) & (!g154) & (g688) & (!g877) & (g929) & (!g1012)) + ((!g125) & (g154) & (!g688) & (!g877) & (!g929) & (!g1012)) + ((!g125) & (g154) & (!g688) & (!g877) & (g929) & (!g1012)) + ((!g125) & (g154) & (!g688) & (g877) & (!g929) & (!g1012)) + ((!g125) & (g154) & (!g688) & (g877) & (g929) & (!g1012)) + ((!g125) & (g154) & (g688) & (!g877) & (!g929) & (!g1012)) + ((!g125) & (g154) & (g688) & (!g877) & (g929) & (!g1012)) + ((!g125) & (g154) & (g688) & (g877) & (!g929) & (!g1012)) + ((!g125) & (g154) & (g688) & (g877) & (g929) & (!g1012)) + ((g125) & (!g154) & (!g688) & (!g877) & (g929) & (!g1012)) + ((g125) & (g154) & (!g688) & (!g877) & (!g929) & (!g1012)) + ((g125) & (g154) & (!g688) & (!g877) & (g929) & (!g1012)) + ((g125) & (g154) & (!g688) & (g877) & (!g929) & (!g1012)) + ((g125) & (g154) & (!g688) & (g877) & (g929) & (!g1012)));
	assign g1235 = (((!g5) & (!sk[113]) & (!g17) & (g69) & (!g174)) + ((!g5) & (!sk[113]) & (!g17) & (g69) & (g174)) + ((!g5) & (!sk[113]) & (g17) & (g69) & (!g174)) + ((!g5) & (!sk[113]) & (g17) & (g69) & (g174)) + ((!g5) & (sk[113]) & (!g17) & (!g69) & (!g174)) + ((!g5) & (sk[113]) & (!g17) & (!g69) & (g174)) + ((!g5) & (sk[113]) & (!g17) & (g69) & (g174)) + ((!g5) & (sk[113]) & (g17) & (!g69) & (g174)) + ((!g5) & (sk[113]) & (g17) & (g69) & (g174)) + ((g5) & (!sk[113]) & (!g17) & (g69) & (!g174)) + ((g5) & (!sk[113]) & (!g17) & (g69) & (g174)) + ((g5) & (!sk[113]) & (g17) & (g69) & (!g174)) + ((g5) & (!sk[113]) & (g17) & (g69) & (g174)));
	assign g1236 = (((!g226) & (!g469) & (!g508) & (!g725) & (sk[114]) & (!g1235)) + ((!g226) & (!g469) & (!g508) & (!g725) & (sk[114]) & (g1235)) + ((!g226) & (!g469) & (!g508) & (g725) & (sk[114]) & (!g1235)) + ((!g226) & (!g469) & (!g508) & (g725) & (sk[114]) & (g1235)) + ((!g226) & (!g469) & (g508) & (!g725) & (!sk[114]) & (g1235)) + ((!g226) & (!g469) & (g508) & (!g725) & (sk[114]) & (!g1235)) + ((!g226) & (!g469) & (g508) & (!g725) & (sk[114]) & (g1235)) + ((!g226) & (!g469) & (g508) & (g725) & (!sk[114]) & (!g1235)) + ((!g226) & (!g469) & (g508) & (g725) & (!sk[114]) & (g1235)) + ((!g226) & (!g469) & (g508) & (g725) & (sk[114]) & (!g1235)) + ((!g226) & (!g469) & (g508) & (g725) & (sk[114]) & (g1235)) + ((!g226) & (g469) & (!g508) & (!g725) & (!sk[114]) & (!g1235)) + ((!g226) & (g469) & (!g508) & (!g725) & (!sk[114]) & (g1235)) + ((!g226) & (g469) & (!g508) & (!g725) & (sk[114]) & (!g1235)) + ((!g226) & (g469) & (!g508) & (!g725) & (sk[114]) & (g1235)) + ((!g226) & (g469) & (!g508) & (g725) & (!sk[114]) & (!g1235)) + ((!g226) & (g469) & (!g508) & (g725) & (!sk[114]) & (g1235)) + ((!g226) & (g469) & (!g508) & (g725) & (sk[114]) & (!g1235)) + ((!g226) & (g469) & (g508) & (!g725) & (!sk[114]) & (!g1235)) + ((!g226) & (g469) & (g508) & (!g725) & (!sk[114]) & (g1235)) + ((!g226) & (g469) & (g508) & (!g725) & (sk[114]) & (!g1235)) + ((!g226) & (g469) & (g508) & (!g725) & (sk[114]) & (g1235)) + ((!g226) & (g469) & (g508) & (g725) & (!sk[114]) & (!g1235)) + ((!g226) & (g469) & (g508) & (g725) & (!sk[114]) & (g1235)) + ((!g226) & (g469) & (g508) & (g725) & (sk[114]) & (!g1235)) + ((!g226) & (g469) & (g508) & (g725) & (sk[114]) & (g1235)) + ((g226) & (!g469) & (g508) & (!g725) & (!sk[114]) & (g1235)) + ((g226) & (!g469) & (g508) & (g725) & (!sk[114]) & (!g1235)) + ((g226) & (!g469) & (g508) & (g725) & (!sk[114]) & (g1235)) + ((g226) & (g469) & (!g508) & (!g725) & (!sk[114]) & (!g1235)) + ((g226) & (g469) & (!g508) & (!g725) & (!sk[114]) & (g1235)) + ((g226) & (g469) & (!g508) & (g725) & (!sk[114]) & (!g1235)) + ((g226) & (g469) & (!g508) & (g725) & (!sk[114]) & (g1235)) + ((g226) & (g469) & (g508) & (!g725) & (!sk[114]) & (!g1235)) + ((g226) & (g469) & (g508) & (!g725) & (!sk[114]) & (g1235)) + ((g226) & (g469) & (g508) & (g725) & (!sk[114]) & (!g1235)) + ((g226) & (g469) & (g508) & (g725) & (!sk[114]) & (g1235)));
	assign g1237 = (((!g164) & (!g341) & (!g742) & (sk[115]) & (!g655) & (!g1236)) + ((!g164) & (!g341) & (!g742) & (sk[115]) & (g655) & (!g1236)) + ((!g164) & (!g341) & (g742) & (!sk[115]) & (!g655) & (g1236)) + ((!g164) & (!g341) & (g742) & (!sk[115]) & (g655) & (!g1236)) + ((!g164) & (!g341) & (g742) & (!sk[115]) & (g655) & (g1236)) + ((!g164) & (!g341) & (g742) & (sk[115]) & (!g655) & (!g1236)) + ((!g164) & (!g341) & (g742) & (sk[115]) & (g655) & (!g1236)) + ((!g164) & (g341) & (!g742) & (!sk[115]) & (!g655) & (!g1236)) + ((!g164) & (g341) & (!g742) & (!sk[115]) & (!g655) & (g1236)) + ((!g164) & (g341) & (!g742) & (!sk[115]) & (g655) & (!g1236)) + ((!g164) & (g341) & (!g742) & (!sk[115]) & (g655) & (g1236)) + ((!g164) & (g341) & (!g742) & (sk[115]) & (!g655) & (!g1236)) + ((!g164) & (g341) & (!g742) & (sk[115]) & (g655) & (!g1236)) + ((!g164) & (g341) & (g742) & (!sk[115]) & (!g655) & (!g1236)) + ((!g164) & (g341) & (g742) & (!sk[115]) & (!g655) & (g1236)) + ((!g164) & (g341) & (g742) & (!sk[115]) & (g655) & (!g1236)) + ((!g164) & (g341) & (g742) & (!sk[115]) & (g655) & (g1236)) + ((!g164) & (g341) & (g742) & (sk[115]) & (!g655) & (!g1236)) + ((!g164) & (g341) & (g742) & (sk[115]) & (g655) & (!g1236)) + ((g164) & (!g341) & (g742) & (!sk[115]) & (!g655) & (g1236)) + ((g164) & (!g341) & (g742) & (!sk[115]) & (g655) & (!g1236)) + ((g164) & (!g341) & (g742) & (!sk[115]) & (g655) & (g1236)) + ((g164) & (g341) & (!g742) & (!sk[115]) & (!g655) & (!g1236)) + ((g164) & (g341) & (!g742) & (!sk[115]) & (!g655) & (g1236)) + ((g164) & (g341) & (!g742) & (!sk[115]) & (g655) & (!g1236)) + ((g164) & (g341) & (!g742) & (!sk[115]) & (g655) & (g1236)) + ((g164) & (g341) & (g742) & (!sk[115]) & (!g655) & (!g1236)) + ((g164) & (g341) & (g742) & (!sk[115]) & (!g655) & (g1236)) + ((g164) & (g341) & (g742) & (!sk[115]) & (g655) & (!g1236)) + ((g164) & (g341) & (g742) & (!sk[115]) & (g655) & (g1236)) + ((g164) & (g341) & (g742) & (sk[115]) & (g655) & (!g1236)));
	assign g1238 = (((!g341) & (!g469) & (!sk[116]) & (g927)) + ((!g341) & (g469) & (!sk[116]) & (!g927)) + ((!g341) & (g469) & (!sk[116]) & (g927)) + ((g341) & (!g469) & (!sk[116]) & (g927)) + ((g341) & (g469) & (!sk[116]) & (!g927)) + ((g341) & (g469) & (!sk[116]) & (g927)) + ((g341) & (g469) & (sk[116]) & (!g927)));
	assign g1239 = (((!g347) & (!g121) & (g725) & (g945) & (!g983) & (!g1238)) + ((!g347) & (!g121) & (g725) & (g945) & (!g983) & (g1238)) + ((!g347) & (g121) & (g725) & (g945) & (!g983) & (g1238)) + ((g347) & (!g121) & (!g725) & (!g945) & (!g983) & (!g1238)) + ((g347) & (!g121) & (!g725) & (!g945) & (!g983) & (g1238)) + ((g347) & (!g121) & (!g725) & (!g945) & (g983) & (!g1238)) + ((g347) & (!g121) & (!g725) & (!g945) & (g983) & (g1238)) + ((g347) & (!g121) & (!g725) & (g945) & (!g983) & (!g1238)) + ((g347) & (!g121) & (!g725) & (g945) & (!g983) & (g1238)) + ((g347) & (!g121) & (!g725) & (g945) & (g983) & (!g1238)) + ((g347) & (!g121) & (!g725) & (g945) & (g983) & (g1238)) + ((g347) & (!g121) & (g725) & (!g945) & (!g983) & (!g1238)) + ((g347) & (!g121) & (g725) & (!g945) & (!g983) & (g1238)) + ((g347) & (!g121) & (g725) & (!g945) & (g983) & (!g1238)) + ((g347) & (!g121) & (g725) & (!g945) & (g983) & (g1238)) + ((g347) & (!g121) & (g725) & (g945) & (!g983) & (!g1238)) + ((g347) & (!g121) & (g725) & (g945) & (!g983) & (g1238)) + ((g347) & (!g121) & (g725) & (g945) & (g983) & (!g1238)) + ((g347) & (!g121) & (g725) & (g945) & (g983) & (g1238)) + ((g347) & (g121) & (!g725) & (!g945) & (!g983) & (g1238)) + ((g347) & (g121) & (!g725) & (!g945) & (g983) & (g1238)) + ((g347) & (g121) & (!g725) & (g945) & (!g983) & (g1238)) + ((g347) & (g121) & (!g725) & (g945) & (g983) & (g1238)) + ((g347) & (g121) & (g725) & (!g945) & (!g983) & (g1238)) + ((g347) & (g121) & (g725) & (!g945) & (g983) & (g1238)) + ((g347) & (g121) & (g725) & (g945) & (!g983) & (g1238)) + ((g347) & (g121) & (g725) & (g945) & (g983) & (g1238)));
	assign g1240 = (((!g290) & (!g1233) & (!sk[118]) & (g1234) & (!g1237) & (g1239)) + ((!g290) & (!g1233) & (!sk[118]) & (g1234) & (g1237) & (!g1239)) + ((!g290) & (!g1233) & (!sk[118]) & (g1234) & (g1237) & (g1239)) + ((!g290) & (g1233) & (!sk[118]) & (!g1234) & (!g1237) & (!g1239)) + ((!g290) & (g1233) & (!sk[118]) & (!g1234) & (!g1237) & (g1239)) + ((!g290) & (g1233) & (!sk[118]) & (!g1234) & (g1237) & (!g1239)) + ((!g290) & (g1233) & (!sk[118]) & (!g1234) & (g1237) & (g1239)) + ((!g290) & (g1233) & (!sk[118]) & (g1234) & (!g1237) & (!g1239)) + ((!g290) & (g1233) & (!sk[118]) & (g1234) & (!g1237) & (g1239)) + ((!g290) & (g1233) & (!sk[118]) & (g1234) & (g1237) & (!g1239)) + ((!g290) & (g1233) & (!sk[118]) & (g1234) & (g1237) & (g1239)) + ((g290) & (!g1233) & (!sk[118]) & (g1234) & (!g1237) & (g1239)) + ((g290) & (!g1233) & (!sk[118]) & (g1234) & (g1237) & (!g1239)) + ((g290) & (!g1233) & (!sk[118]) & (g1234) & (g1237) & (g1239)) + ((g290) & (!g1233) & (sk[118]) & (g1234) & (g1237) & (g1239)) + ((g290) & (g1233) & (!sk[118]) & (!g1234) & (!g1237) & (!g1239)) + ((g290) & (g1233) & (!sk[118]) & (!g1234) & (!g1237) & (g1239)) + ((g290) & (g1233) & (!sk[118]) & (!g1234) & (g1237) & (!g1239)) + ((g290) & (g1233) & (!sk[118]) & (!g1234) & (g1237) & (g1239)) + ((g290) & (g1233) & (!sk[118]) & (g1234) & (!g1237) & (!g1239)) + ((g290) & (g1233) & (!sk[118]) & (g1234) & (!g1237) & (g1239)) + ((g290) & (g1233) & (!sk[118]) & (g1234) & (g1237) & (!g1239)) + ((g290) & (g1233) & (!sk[118]) & (g1234) & (g1237) & (g1239)));
	assign g1241 = (((!g24) & (!sk[119]) & (!g113) & (g174) & (!g857)) + ((!g24) & (!sk[119]) & (!g113) & (g174) & (g857)) + ((!g24) & (!sk[119]) & (g113) & (g174) & (!g857)) + ((!g24) & (!sk[119]) & (g113) & (g174) & (g857)) + ((!g24) & (sk[119]) & (g113) & (!g174) & (!g857)) + ((!g24) & (sk[119]) & (g113) & (g174) & (!g857)) + ((g24) & (!sk[119]) & (!g113) & (g174) & (!g857)) + ((g24) & (!sk[119]) & (!g113) & (g174) & (g857)) + ((g24) & (!sk[119]) & (g113) & (g174) & (!g857)) + ((g24) & (!sk[119]) & (g113) & (g174) & (g857)) + ((g24) & (sk[119]) & (!g113) & (g174) & (!g857)) + ((g24) & (sk[119]) & (g113) & (!g174) & (!g857)) + ((g24) & (sk[119]) & (g113) & (g174) & (!g857)));
	assign g1242 = (((!sk[120]) & (!g383) & (!g469) & (g928) & (!g971) & (g1241)) + ((!sk[120]) & (!g383) & (!g469) & (g928) & (g971) & (!g1241)) + ((!sk[120]) & (!g383) & (!g469) & (g928) & (g971) & (g1241)) + ((!sk[120]) & (!g383) & (g469) & (!g928) & (!g971) & (!g1241)) + ((!sk[120]) & (!g383) & (g469) & (!g928) & (!g971) & (g1241)) + ((!sk[120]) & (!g383) & (g469) & (!g928) & (g971) & (!g1241)) + ((!sk[120]) & (!g383) & (g469) & (!g928) & (g971) & (g1241)) + ((!sk[120]) & (!g383) & (g469) & (g928) & (!g971) & (!g1241)) + ((!sk[120]) & (!g383) & (g469) & (g928) & (!g971) & (g1241)) + ((!sk[120]) & (!g383) & (g469) & (g928) & (g971) & (!g1241)) + ((!sk[120]) & (!g383) & (g469) & (g928) & (g971) & (g1241)) + ((!sk[120]) & (g383) & (!g469) & (g928) & (!g971) & (g1241)) + ((!sk[120]) & (g383) & (!g469) & (g928) & (g971) & (!g1241)) + ((!sk[120]) & (g383) & (!g469) & (g928) & (g971) & (g1241)) + ((!sk[120]) & (g383) & (g469) & (!g928) & (!g971) & (!g1241)) + ((!sk[120]) & (g383) & (g469) & (!g928) & (!g971) & (g1241)) + ((!sk[120]) & (g383) & (g469) & (!g928) & (g971) & (!g1241)) + ((!sk[120]) & (g383) & (g469) & (!g928) & (g971) & (g1241)) + ((!sk[120]) & (g383) & (g469) & (g928) & (!g971) & (!g1241)) + ((!sk[120]) & (g383) & (g469) & (g928) & (!g971) & (g1241)) + ((!sk[120]) & (g383) & (g469) & (g928) & (g971) & (!g1241)) + ((!sk[120]) & (g383) & (g469) & (g928) & (g971) & (g1241)) + ((sk[120]) & (!g383) & (!g469) & (!g928) & (!g971) & (!g1241)) + ((sk[120]) & (!g383) & (!g469) & (!g928) & (!g971) & (g1241)) + ((sk[120]) & (!g383) & (!g469) & (!g928) & (g971) & (!g1241)) + ((sk[120]) & (!g383) & (!g469) & (!g928) & (g971) & (g1241)) + ((sk[120]) & (!g383) & (!g469) & (g928) & (!g971) & (!g1241)) + ((sk[120]) & (!g383) & (!g469) & (g928) & (!g971) & (g1241)) + ((sk[120]) & (!g383) & (!g469) & (g928) & (g971) & (!g1241)) + ((sk[120]) & (!g383) & (!g469) & (g928) & (g971) & (g1241)) + ((sk[120]) & (!g383) & (g469) & (!g928) & (!g971) & (!g1241)) + ((sk[120]) & (!g383) & (g469) & (!g928) & (!g971) & (g1241)) + ((sk[120]) & (!g383) & (g469) & (!g928) & (g971) & (!g1241)) + ((sk[120]) & (!g383) & (g469) & (!g928) & (g971) & (g1241)) + ((sk[120]) & (!g383) & (g469) & (g928) & (!g971) & (!g1241)) + ((sk[120]) & (!g383) & (g469) & (g928) & (!g971) & (g1241)) + ((sk[120]) & (!g383) & (g469) & (g928) & (g971) & (!g1241)));
	assign g1243 = (((!g77) & (!sk[121]) & (!g105) & (g927) & (!g945)) + ((!g77) & (!sk[121]) & (!g105) & (g927) & (g945)) + ((!g77) & (!sk[121]) & (g105) & (g927) & (!g945)) + ((!g77) & (!sk[121]) & (g105) & (g927) & (g945)) + ((!g77) & (sk[121]) & (!g105) & (!g927) & (!g945)) + ((!g77) & (sk[121]) & (!g105) & (g927) & (!g945)) + ((!g77) & (sk[121]) & (!g105) & (g927) & (g945)) + ((g77) & (!sk[121]) & (!g105) & (g927) & (!g945)) + ((g77) & (!sk[121]) & (!g105) & (g927) & (g945)) + ((g77) & (!sk[121]) & (g105) & (g927) & (!g945)) + ((g77) & (!sk[121]) & (g105) & (g927) & (g945)) + ((g77) & (sk[121]) & (!g105) & (!g927) & (!g945)) + ((g77) & (sk[121]) & (!g105) & (!g927) & (g945)) + ((g77) & (sk[121]) & (!g105) & (g927) & (!g945)) + ((g77) & (sk[121]) & (!g105) & (g927) & (g945)));
	assign g1244 = (((!sk[122]) & (!g125) & (!g205) & (g761) & (!g1243)) + ((!sk[122]) & (!g125) & (!g205) & (g761) & (g1243)) + ((!sk[122]) & (!g125) & (g205) & (g761) & (!g1243)) + ((!sk[122]) & (!g125) & (g205) & (g761) & (g1243)) + ((!sk[122]) & (g125) & (!g205) & (g761) & (!g1243)) + ((!sk[122]) & (g125) & (!g205) & (g761) & (g1243)) + ((!sk[122]) & (g125) & (g205) & (g761) & (!g1243)) + ((!sk[122]) & (g125) & (g205) & (g761) & (g1243)) + ((sk[122]) & (!g125) & (!g205) & (!g761) & (!g1243)) + ((sk[122]) & (!g125) & (!g205) & (g761) & (!g1243)) + ((sk[122]) & (g125) & (!g205) & (g761) & (!g1243)));
	assign g1245 = (((!g3) & (!i_12_) & (!i_13_) & (!i_14_) & (!g75) & (g69)) + ((!g3) & (i_12_) & (!i_13_) & (!i_14_) & (!g75) & (g69)) + ((!g3) & (i_12_) & (!i_13_) & (i_14_) & (!g75) & (g69)) + ((g3) & (!i_12_) & (!i_13_) & (!i_14_) & (!g75) & (g69)) + ((g3) & (!i_12_) & (i_13_) & (!i_14_) & (!g75) & (!g69)) + ((g3) & (!i_12_) & (i_13_) & (!i_14_) & (!g75) & (g69)) + ((g3) & (!i_12_) & (i_13_) & (i_14_) & (!g75) & (!g69)) + ((g3) & (!i_12_) & (i_13_) & (i_14_) & (!g75) & (g69)) + ((g3) & (i_12_) & (!i_13_) & (!i_14_) & (!g75) & (g69)) + ((g3) & (i_12_) & (!i_13_) & (i_14_) & (!g75) & (g69)) + ((g3) & (i_12_) & (i_13_) & (!i_14_) & (!g75) & (!g69)) + ((g3) & (i_12_) & (i_13_) & (!i_14_) & (!g75) & (g69)) + ((g3) & (i_12_) & (i_13_) & (i_14_) & (!g75) & (!g69)) + ((g3) & (i_12_) & (i_13_) & (i_14_) & (!g75) & (g69)));
	assign g1246 = (((g944) & (!g1242) & (g129) & (g391) & (g1244) & (!g1245)));
	assign g1247 = (((!i_15_) & (!sk[125]) & (!g125) & (g112) & (!g122) & (g460)) + ((!i_15_) & (!sk[125]) & (!g125) & (g112) & (g122) & (!g460)) + ((!i_15_) & (!sk[125]) & (!g125) & (g112) & (g122) & (g460)) + ((!i_15_) & (!sk[125]) & (g125) & (!g112) & (!g122) & (!g460)) + ((!i_15_) & (!sk[125]) & (g125) & (!g112) & (!g122) & (g460)) + ((!i_15_) & (!sk[125]) & (g125) & (!g112) & (g122) & (!g460)) + ((!i_15_) & (!sk[125]) & (g125) & (!g112) & (g122) & (g460)) + ((!i_15_) & (!sk[125]) & (g125) & (g112) & (!g122) & (!g460)) + ((!i_15_) & (!sk[125]) & (g125) & (g112) & (!g122) & (g460)) + ((!i_15_) & (!sk[125]) & (g125) & (g112) & (g122) & (!g460)) + ((!i_15_) & (!sk[125]) & (g125) & (g112) & (g122) & (g460)) + ((!i_15_) & (sk[125]) & (g125) & (g112) & (!g122) & (!g460)) + ((!i_15_) & (sk[125]) & (g125) & (g112) & (g122) & (!g460)) + ((i_15_) & (!sk[125]) & (!g125) & (g112) & (!g122) & (g460)) + ((i_15_) & (!sk[125]) & (!g125) & (g112) & (g122) & (!g460)) + ((i_15_) & (!sk[125]) & (!g125) & (g112) & (g122) & (g460)) + ((i_15_) & (!sk[125]) & (g125) & (!g112) & (!g122) & (!g460)) + ((i_15_) & (!sk[125]) & (g125) & (!g112) & (!g122) & (g460)) + ((i_15_) & (!sk[125]) & (g125) & (!g112) & (g122) & (!g460)) + ((i_15_) & (!sk[125]) & (g125) & (!g112) & (g122) & (g460)) + ((i_15_) & (!sk[125]) & (g125) & (g112) & (!g122) & (!g460)) + ((i_15_) & (!sk[125]) & (g125) & (g112) & (!g122) & (g460)) + ((i_15_) & (!sk[125]) & (g125) & (g112) & (g122) & (!g460)) + ((i_15_) & (!sk[125]) & (g125) & (g112) & (g122) & (g460)) + ((i_15_) & (sk[125]) & (!g125) & (g112) & (g122) & (!g460)) + ((i_15_) & (sk[125]) & (g125) & (g112) & (g122) & (!g460)));
	assign g1248 = (((!i_15_) & (!sk[126]) & (!i_12_) & (i_13_) & (!i_14_) & (g428)) + ((!i_15_) & (!sk[126]) & (!i_12_) & (i_13_) & (i_14_) & (!g428)) + ((!i_15_) & (!sk[126]) & (!i_12_) & (i_13_) & (i_14_) & (g428)) + ((!i_15_) & (!sk[126]) & (i_12_) & (!i_13_) & (!i_14_) & (!g428)) + ((!i_15_) & (!sk[126]) & (i_12_) & (!i_13_) & (!i_14_) & (g428)) + ((!i_15_) & (!sk[126]) & (i_12_) & (!i_13_) & (i_14_) & (!g428)) + ((!i_15_) & (!sk[126]) & (i_12_) & (!i_13_) & (i_14_) & (g428)) + ((!i_15_) & (!sk[126]) & (i_12_) & (i_13_) & (!i_14_) & (!g428)) + ((!i_15_) & (!sk[126]) & (i_12_) & (i_13_) & (!i_14_) & (g428)) + ((!i_15_) & (!sk[126]) & (i_12_) & (i_13_) & (i_14_) & (!g428)) + ((!i_15_) & (!sk[126]) & (i_12_) & (i_13_) & (i_14_) & (g428)) + ((!i_15_) & (sk[126]) & (!i_12_) & (!i_13_) & (i_14_) & (!g428)) + ((!i_15_) & (sk[126]) & (i_12_) & (!i_13_) & (i_14_) & (!g428)) + ((i_15_) & (!sk[126]) & (!i_12_) & (i_13_) & (!i_14_) & (g428)) + ((i_15_) & (!sk[126]) & (!i_12_) & (i_13_) & (i_14_) & (!g428)) + ((i_15_) & (!sk[126]) & (!i_12_) & (i_13_) & (i_14_) & (g428)) + ((i_15_) & (!sk[126]) & (i_12_) & (!i_13_) & (!i_14_) & (!g428)) + ((i_15_) & (!sk[126]) & (i_12_) & (!i_13_) & (!i_14_) & (g428)) + ((i_15_) & (!sk[126]) & (i_12_) & (!i_13_) & (i_14_) & (!g428)) + ((i_15_) & (!sk[126]) & (i_12_) & (!i_13_) & (i_14_) & (g428)) + ((i_15_) & (!sk[126]) & (i_12_) & (i_13_) & (!i_14_) & (!g428)) + ((i_15_) & (!sk[126]) & (i_12_) & (i_13_) & (!i_14_) & (g428)) + ((i_15_) & (!sk[126]) & (i_12_) & (i_13_) & (i_14_) & (!g428)) + ((i_15_) & (!sk[126]) & (i_12_) & (i_13_) & (i_14_) & (g428)) + ((i_15_) & (sk[126]) & (!i_12_) & (i_13_) & (!i_14_) & (!g428)) + ((i_15_) & (sk[126]) & (i_12_) & (!i_13_) & (!i_14_) & (!g428)) + ((i_15_) & (sk[126]) & (i_12_) & (i_13_) & (!i_14_) & (!g428)));
	assign g1249 = (((!sk[127]) & (!g123) & (!g1248) & (g974)) + ((!sk[127]) & (!g123) & (g1248) & (!g974)) + ((!sk[127]) & (!g123) & (g1248) & (g974)) + ((!sk[127]) & (g123) & (!g1248) & (g974)) + ((!sk[127]) & (g123) & (g1248) & (!g974)) + ((!sk[127]) & (g123) & (g1248) & (g974)) + ((sk[127]) & (!g123) & (!g1248) & (g974)) + ((sk[127]) & (!g123) & (g1248) & (!g974)) + ((sk[127]) & (!g123) & (g1248) & (g974)));
	assign g1250 = (((!g164) & (!g347) & (!g557) & (g898) & (!g1247) & (!g1249)) + ((!g164) & (!g347) & (g557) & (g898) & (!g1247) & (!g1249)) + ((!g164) & (g347) & (!g557) & (!g898) & (!g1247) & (!g1249)) + ((!g164) & (g347) & (!g557) & (g898) & (!g1247) & (!g1249)) + ((!g164) & (g347) & (g557) & (!g898) & (!g1247) & (!g1249)) + ((!g164) & (g347) & (g557) & (g898) & (!g1247) & (!g1249)) + ((g164) & (!g347) & (!g557) & (g898) & (!g1247) & (!g1249)) + ((g164) & (g347) & (!g557) & (!g898) & (!g1247) & (!g1249)) + ((g164) & (g347) & (!g557) & (g898) & (!g1247) & (!g1249)));
	assign g1251 = (((!g122) & (!g933) & (g559) & (g532) & (g1457) & (g1250)) + ((!g122) & (g933) & (g559) & (g532) & (g1457) & (g1250)) + ((g122) & (g933) & (g559) & (g532) & (g1457) & (g1250)));
	assign g1252 = (((g1224) & (!g1228) & (g1232) & (g1240) & (g1246) & (g1251)));
	assign g1253 = (((g1152) & (g1172) & (g1183) & (g1207) & (g1208) & (g1252)));
	assign g1254 = (((!i_12_) & (!i_13_) & (!i_14_) & (!g107) & (!g91) & (!g130)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g107) & (!g91) & (!g130)) + ((!i_12_) & (!i_13_) & (i_14_) & (!g107) & (!g91) & (!g130)) + ((!i_12_) & (!i_13_) & (i_14_) & (!g107) & (g91) & (!g130)) + ((!i_12_) & (!i_13_) & (i_14_) & (g107) & (!g91) & (!g130)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g107) & (!g91) & (!g130)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g107) & (g91) & (!g130)) + ((!i_12_) & (i_13_) & (i_14_) & (!g107) & (!g91) & (!g130)) + ((!i_12_) & (i_13_) & (i_14_) & (!g107) & (g91) & (!g130)) + ((!i_12_) & (i_13_) & (i_14_) & (g107) & (!g91) & (!g130)) + ((i_12_) & (!i_13_) & (!i_14_) & (!g107) & (!g91) & (!g130)) + ((i_12_) & (!i_13_) & (!i_14_) & (!g107) & (g91) & (!g130)) + ((i_12_) & (!i_13_) & (!i_14_) & (g107) & (!g91) & (!g130)) + ((i_12_) & (!i_13_) & (i_14_) & (!g107) & (!g91) & (!g130)) + ((i_12_) & (!i_13_) & (i_14_) & (!g107) & (g91) & (!g130)) + ((i_12_) & (!i_13_) & (i_14_) & (g107) & (!g91) & (!g130)) + ((i_12_) & (i_13_) & (!i_14_) & (!g107) & (!g91) & (!g130)) + ((i_12_) & (i_13_) & (!i_14_) & (!g107) & (g91) & (!g130)) + ((i_12_) & (i_13_) & (!i_14_) & (g107) & (!g91) & (!g130)) + ((i_12_) & (i_13_) & (i_14_) & (!g107) & (!g91) & (!g130)) + ((i_12_) & (i_13_) & (i_14_) & (!g107) & (g91) & (!g130)));
	assign g1255 = (((!i_12_) & (!i_13_) & (i_14_) & (!g107) & (!sk[5]) & (g102)) + ((!i_12_) & (!i_13_) & (i_14_) & (!g107) & (sk[5]) & (g102)) + ((!i_12_) & (!i_13_) & (i_14_) & (g107) & (!sk[5]) & (!g102)) + ((!i_12_) & (!i_13_) & (i_14_) & (g107) & (!sk[5]) & (g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g107) & (!sk[5]) & (!g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g107) & (!sk[5]) & (g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g107) & (sk[5]) & (g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (g107) & (!sk[5]) & (!g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (g107) & (!sk[5]) & (g102)) + ((!i_12_) & (i_13_) & (i_14_) & (!g107) & (!sk[5]) & (!g102)) + ((!i_12_) & (i_13_) & (i_14_) & (!g107) & (!sk[5]) & (g102)) + ((!i_12_) & (i_13_) & (i_14_) & (!g107) & (sk[5]) & (g102)) + ((!i_12_) & (i_13_) & (i_14_) & (g107) & (!sk[5]) & (!g102)) + ((!i_12_) & (i_13_) & (i_14_) & (g107) & (!sk[5]) & (g102)) + ((i_12_) & (!i_13_) & (!i_14_) & (!g107) & (sk[5]) & (g102)) + ((i_12_) & (!i_13_) & (i_14_) & (!g107) & (!sk[5]) & (g102)) + ((i_12_) & (!i_13_) & (i_14_) & (g107) & (!sk[5]) & (!g102)) + ((i_12_) & (!i_13_) & (i_14_) & (g107) & (!sk[5]) & (g102)) + ((i_12_) & (i_13_) & (!i_14_) & (!g107) & (!sk[5]) & (!g102)) + ((i_12_) & (i_13_) & (!i_14_) & (!g107) & (!sk[5]) & (g102)) + ((i_12_) & (i_13_) & (!i_14_) & (!g107) & (sk[5]) & (g102)) + ((i_12_) & (i_13_) & (!i_14_) & (g107) & (!sk[5]) & (!g102)) + ((i_12_) & (i_13_) & (!i_14_) & (g107) & (!sk[5]) & (g102)) + ((i_12_) & (i_13_) & (i_14_) & (!g107) & (!sk[5]) & (!g102)) + ((i_12_) & (i_13_) & (i_14_) & (!g107) & (!sk[5]) & (g102)) + ((i_12_) & (i_13_) & (i_14_) & (g107) & (!sk[5]) & (!g102)) + ((i_12_) & (i_13_) & (i_14_) & (g107) & (!sk[5]) & (g102)));
	assign g1256 = (((!i_8_) & (!g73) & (g107) & (!g176) & (!sk[6]) & (g460)) + ((!i_8_) & (!g73) & (g107) & (g176) & (!sk[6]) & (!g460)) + ((!i_8_) & (!g73) & (g107) & (g176) & (!sk[6]) & (g460)) + ((!i_8_) & (g73) & (!g107) & (!g176) & (!sk[6]) & (!g460)) + ((!i_8_) & (g73) & (!g107) & (!g176) & (!sk[6]) & (g460)) + ((!i_8_) & (g73) & (!g107) & (!g176) & (sk[6]) & (!g460)) + ((!i_8_) & (g73) & (!g107) & (!g176) & (sk[6]) & (g460)) + ((!i_8_) & (g73) & (!g107) & (g176) & (!sk[6]) & (!g460)) + ((!i_8_) & (g73) & (!g107) & (g176) & (!sk[6]) & (g460)) + ((!i_8_) & (g73) & (!g107) & (g176) & (sk[6]) & (!g460)) + ((!i_8_) & (g73) & (g107) & (!g176) & (!sk[6]) & (!g460)) + ((!i_8_) & (g73) & (g107) & (!g176) & (!sk[6]) & (g460)) + ((!i_8_) & (g73) & (g107) & (g176) & (!sk[6]) & (!g460)) + ((!i_8_) & (g73) & (g107) & (g176) & (!sk[6]) & (g460)) + ((i_8_) & (!g73) & (g107) & (!g176) & (!sk[6]) & (g460)) + ((i_8_) & (!g73) & (g107) & (g176) & (!sk[6]) & (!g460)) + ((i_8_) & (!g73) & (g107) & (g176) & (!sk[6]) & (g460)) + ((i_8_) & (g73) & (!g107) & (!g176) & (!sk[6]) & (!g460)) + ((i_8_) & (g73) & (!g107) & (!g176) & (!sk[6]) & (g460)) + ((i_8_) & (g73) & (!g107) & (g176) & (!sk[6]) & (!g460)) + ((i_8_) & (g73) & (!g107) & (g176) & (!sk[6]) & (g460)) + ((i_8_) & (g73) & (g107) & (!g176) & (!sk[6]) & (!g460)) + ((i_8_) & (g73) & (g107) & (!g176) & (!sk[6]) & (g460)) + ((i_8_) & (g73) & (g107) & (g176) & (!sk[6]) & (!g460)) + ((i_8_) & (g73) & (g107) & (g176) & (!sk[6]) & (g460)));
	assign g1257 = (((!i_12_) & (!i_13_) & (!i_14_) & (sk[7]) & (g102) & (!g91)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[7]) & (!g102) & (g91)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[7]) & (g102) & (!g91)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[7]) & (g102) & (g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[7]) & (!g102) & (!g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[7]) & (!g102) & (g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[7]) & (g102) & (!g91)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[7]) & (g102) & (g91)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[7]) & (!g102) & (!g91)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[7]) & (!g102) & (g91)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[7]) & (g102) & (!g91)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[7]) & (g102) & (g91)) + ((i_12_) & (!i_13_) & (!i_14_) & (sk[7]) & (g102) & (!g91)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[7]) & (!g102) & (g91)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[7]) & (g102) & (!g91)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[7]) & (g102) & (g91)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[7]) & (!g102) & (!g91)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[7]) & (!g102) & (g91)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[7]) & (g102) & (!g91)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[7]) & (g102) & (g91)) + ((i_12_) & (i_13_) & (!i_14_) & (sk[7]) & (g102) & (!g91)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[7]) & (!g102) & (!g91)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[7]) & (!g102) & (g91)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[7]) & (g102) & (!g91)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[7]) & (g102) & (g91)));
	assign g1258 = (((!g159) & (!g253) & (!g852) & (!g853) & (sk[8]) & (g964)) + ((!g159) & (!g253) & (g852) & (!g853) & (!sk[8]) & (g964)) + ((!g159) & (!g253) & (g852) & (g853) & (!sk[8]) & (!g964)) + ((!g159) & (!g253) & (g852) & (g853) & (!sk[8]) & (g964)) + ((!g159) & (g253) & (!g852) & (!g853) & (!sk[8]) & (!g964)) + ((!g159) & (g253) & (!g852) & (!g853) & (!sk[8]) & (g964)) + ((!g159) & (g253) & (!g852) & (!g853) & (sk[8]) & (!g964)) + ((!g159) & (g253) & (!g852) & (!g853) & (sk[8]) & (g964)) + ((!g159) & (g253) & (!g852) & (g853) & (!sk[8]) & (!g964)) + ((!g159) & (g253) & (!g852) & (g853) & (!sk[8]) & (g964)) + ((!g159) & (g253) & (g852) & (!g853) & (!sk[8]) & (!g964)) + ((!g159) & (g253) & (g852) & (!g853) & (!sk[8]) & (g964)) + ((!g159) & (g253) & (g852) & (g853) & (!sk[8]) & (!g964)) + ((!g159) & (g253) & (g852) & (g853) & (!sk[8]) & (g964)) + ((g159) & (!g253) & (!g852) & (!g853) & (sk[8]) & (g964)) + ((g159) & (!g253) & (g852) & (!g853) & (!sk[8]) & (g964)) + ((g159) & (!g253) & (g852) & (g853) & (!sk[8]) & (!g964)) + ((g159) & (!g253) & (g852) & (g853) & (!sk[8]) & (g964)) + ((g159) & (g253) & (!g852) & (!g853) & (!sk[8]) & (!g964)) + ((g159) & (g253) & (!g852) & (!g853) & (!sk[8]) & (g964)) + ((g159) & (g253) & (!g852) & (!g853) & (sk[8]) & (!g964)) + ((g159) & (g253) & (!g852) & (!g853) & (sk[8]) & (g964)) + ((g159) & (g253) & (!g852) & (g853) & (!sk[8]) & (!g964)) + ((g159) & (g253) & (!g852) & (g853) & (!sk[8]) & (g964)) + ((g159) & (g253) & (!g852) & (g853) & (sk[8]) & (!g964)) + ((g159) & (g253) & (!g852) & (g853) & (sk[8]) & (g964)) + ((g159) & (g253) & (g852) & (!g853) & (!sk[8]) & (!g964)) + ((g159) & (g253) & (g852) & (!g853) & (!sk[8]) & (g964)) + ((g159) & (g253) & (g852) & (!g853) & (sk[8]) & (!g964)) + ((g159) & (g253) & (g852) & (!g853) & (sk[8]) & (g964)) + ((g159) & (g253) & (g852) & (g853) & (!sk[8]) & (!g964)) + ((g159) & (g253) & (g852) & (g853) & (!sk[8]) & (g964)) + ((g159) & (g253) & (g852) & (g853) & (sk[8]) & (!g964)) + ((g159) & (g253) & (g852) & (g853) & (sk[8]) & (g964)));
	assign g1259 = (((!g1255) & (!g1256) & (!g1257) & (sk[9]) & (g1258)) + ((!g1255) & (!g1256) & (g1257) & (!sk[9]) & (!g1258)) + ((!g1255) & (!g1256) & (g1257) & (!sk[9]) & (g1258)) + ((!g1255) & (g1256) & (g1257) & (!sk[9]) & (!g1258)) + ((!g1255) & (g1256) & (g1257) & (!sk[9]) & (g1258)) + ((g1255) & (!g1256) & (g1257) & (!sk[9]) & (!g1258)) + ((g1255) & (!g1256) & (g1257) & (!sk[9]) & (g1258)) + ((g1255) & (g1256) & (g1257) & (!sk[9]) & (!g1258)) + ((g1255) & (g1256) & (g1257) & (!sk[9]) & (g1258)));
	assign g1260 = (((!sk[10]) & (g130) & (!g652)) + ((!sk[10]) & (g130) & (g652)) + ((sk[10]) & (!g130) & (g652)));
	assign g1261 = (((!i_8_) & (!sk[11]) & (!g4) & (g73) & (!g91)) + ((!i_8_) & (!sk[11]) & (!g4) & (g73) & (g91)) + ((!i_8_) & (!sk[11]) & (g4) & (g73) & (!g91)) + ((!i_8_) & (!sk[11]) & (g4) & (g73) & (g91)) + ((!i_8_) & (sk[11]) & (g4) & (g73) & (!g91)) + ((i_8_) & (!sk[11]) & (!g4) & (g73) & (!g91)) + ((i_8_) & (!sk[11]) & (!g4) & (g73) & (g91)) + ((i_8_) & (!sk[11]) & (g4) & (g73) & (!g91)) + ((i_8_) & (!sk[11]) & (g4) & (g73) & (g91)));
	assign g1262 = (((!sk[12]) & (!g135) & (!g131) & (g296) & (!g651)) + ((!sk[12]) & (!g135) & (!g131) & (g296) & (g651)) + ((!sk[12]) & (!g135) & (g131) & (g296) & (!g651)) + ((!sk[12]) & (!g135) & (g131) & (g296) & (g651)) + ((!sk[12]) & (g135) & (!g131) & (g296) & (!g651)) + ((!sk[12]) & (g135) & (!g131) & (g296) & (g651)) + ((!sk[12]) & (g135) & (g131) & (g296) & (!g651)) + ((!sk[12]) & (g135) & (g131) & (g296) & (g651)) + ((sk[12]) & (!g135) & (!g131) & (!g296) & (!g651)) + ((sk[12]) & (!g135) & (g131) & (!g296) & (!g651)) + ((sk[12]) & (g135) & (!g131) & (!g296) & (!g651)) + ((sk[12]) & (g135) & (g131) & (!g296) & (!g651)) + ((sk[12]) & (g135) & (g131) & (!g296) & (g651)) + ((sk[12]) & (g135) & (g131) & (g296) & (!g651)) + ((sk[12]) & (g135) & (g131) & (g296) & (g651)));
	assign g1263 = (((!i_8_) & (!g19) & (g73) & (!g107) & (!g68) & (!g91)) + ((!i_8_) & (!g19) & (g73) & (!g107) & (!g68) & (g91)) + ((!i_8_) & (!g19) & (g73) & (g107) & (!g68) & (!g91)) + ((!i_8_) & (g19) & (g73) & (!g107) & (!g68) & (!g91)) + ((!i_8_) & (g19) & (g73) & (!g107) & (!g68) & (g91)) + ((!i_8_) & (g19) & (g73) & (!g107) & (g68) & (!g91)) + ((!i_8_) & (g19) & (g73) & (!g107) & (g68) & (g91)) + ((!i_8_) & (g19) & (g73) & (g107) & (!g68) & (!g91)) + ((!i_8_) & (g19) & (g73) & (g107) & (g68) & (!g91)));
	assign g1264 = (((!g131) & (g1028) & (!g1260) & (!g1261) & (g1262) & (!g1263)) + ((g131) & (!g1028) & (!g1260) & (!g1261) & (g1262) & (!g1263)) + ((g131) & (g1028) & (!g1260) & (!g1261) & (g1262) & (!g1263)));
	assign g1265 = (((!i_11_) & (!sk[15]) & (!g34) & (g101) & (!g394)) + ((!i_11_) & (!sk[15]) & (!g34) & (g101) & (g394)) + ((!i_11_) & (!sk[15]) & (g34) & (g101) & (!g394)) + ((!i_11_) & (!sk[15]) & (g34) & (g101) & (g394)) + ((i_11_) & (!sk[15]) & (!g34) & (g101) & (!g394)) + ((i_11_) & (!sk[15]) & (!g34) & (g101) & (g394)) + ((i_11_) & (!sk[15]) & (g34) & (g101) & (!g394)) + ((i_11_) & (!sk[15]) & (g34) & (g101) & (g394)) + ((i_11_) & (sk[15]) & (g34) & (g101) & (g394)));
	assign g1266 = (((!g131) & (!g348) & (!g487) & (!g852) & (g964) & (!g1265)) + ((!g131) & (g348) & (!g487) & (!g852) & (g964) & (!g1265)) + ((!g131) & (g348) & (g487) & (!g852) & (g964) & (!g1265)) + ((g131) & (!g348) & (!g487) & (!g852) & (!g964) & (!g1265)) + ((g131) & (!g348) & (!g487) & (!g852) & (g964) & (!g1265)) + ((g131) & (g348) & (!g487) & (!g852) & (!g964) & (!g1265)) + ((g131) & (g348) & (!g487) & (!g852) & (g964) & (!g1265)) + ((g131) & (g348) & (!g487) & (g852) & (!g964) & (!g1265)) + ((g131) & (g348) & (!g487) & (g852) & (g964) & (!g1265)) + ((g131) & (g348) & (g487) & (!g852) & (!g964) & (!g1265)) + ((g131) & (g348) & (g487) & (!g852) & (g964) & (!g1265)) + ((g131) & (g348) & (g487) & (g852) & (!g964) & (!g1265)) + ((g131) & (g348) & (g487) & (g852) & (g964) & (!g1265)));
	assign g1267 = (((!i_12_) & (!sk[17]) & (!i_13_) & (i_14_) & (!g107) & (g91)) + ((!i_12_) & (!sk[17]) & (!i_13_) & (i_14_) & (g107) & (!g91)) + ((!i_12_) & (!sk[17]) & (!i_13_) & (i_14_) & (g107) & (g91)) + ((!i_12_) & (!sk[17]) & (i_13_) & (!i_14_) & (!g107) & (!g91)) + ((!i_12_) & (!sk[17]) & (i_13_) & (!i_14_) & (!g107) & (g91)) + ((!i_12_) & (!sk[17]) & (i_13_) & (!i_14_) & (g107) & (!g91)) + ((!i_12_) & (!sk[17]) & (i_13_) & (!i_14_) & (g107) & (g91)) + ((!i_12_) & (!sk[17]) & (i_13_) & (i_14_) & (!g107) & (!g91)) + ((!i_12_) & (!sk[17]) & (i_13_) & (i_14_) & (!g107) & (g91)) + ((!i_12_) & (!sk[17]) & (i_13_) & (i_14_) & (g107) & (!g91)) + ((!i_12_) & (!sk[17]) & (i_13_) & (i_14_) & (g107) & (g91)) + ((!i_12_) & (sk[17]) & (!i_13_) & (!i_14_) & (!g107) & (!g91)) + ((!i_12_) & (sk[17]) & (!i_13_) & (!i_14_) & (g107) & (!g91)) + ((!i_12_) & (sk[17]) & (!i_13_) & (i_14_) & (!g107) & (!g91)) + ((!i_12_) & (sk[17]) & (!i_13_) & (i_14_) & (!g107) & (g91)) + ((!i_12_) & (sk[17]) & (!i_13_) & (i_14_) & (g107) & (!g91)) + ((!i_12_) & (sk[17]) & (i_13_) & (i_14_) & (!g107) & (!g91)) + ((!i_12_) & (sk[17]) & (i_13_) & (i_14_) & (!g107) & (g91)) + ((i_12_) & (!sk[17]) & (!i_13_) & (i_14_) & (!g107) & (g91)) + ((i_12_) & (!sk[17]) & (!i_13_) & (i_14_) & (g107) & (!g91)) + ((i_12_) & (!sk[17]) & (!i_13_) & (i_14_) & (g107) & (g91)) + ((i_12_) & (!sk[17]) & (i_13_) & (!i_14_) & (!g107) & (!g91)) + ((i_12_) & (!sk[17]) & (i_13_) & (!i_14_) & (!g107) & (g91)) + ((i_12_) & (!sk[17]) & (i_13_) & (!i_14_) & (g107) & (!g91)) + ((i_12_) & (!sk[17]) & (i_13_) & (!i_14_) & (g107) & (g91)) + ((i_12_) & (!sk[17]) & (i_13_) & (i_14_) & (!g107) & (!g91)) + ((i_12_) & (!sk[17]) & (i_13_) & (i_14_) & (!g107) & (g91)) + ((i_12_) & (!sk[17]) & (i_13_) & (i_14_) & (g107) & (!g91)) + ((i_12_) & (!sk[17]) & (i_13_) & (i_14_) & (g107) & (g91)) + ((i_12_) & (sk[17]) & (!i_13_) & (!i_14_) & (!g107) & (!g91)) + ((i_12_) & (sk[17]) & (!i_13_) & (!i_14_) & (g107) & (!g91)) + ((i_12_) & (sk[17]) & (i_13_) & (!i_14_) & (!g107) & (!g91)) + ((i_12_) & (sk[17]) & (i_13_) & (!i_14_) & (!g107) & (g91)) + ((i_12_) & (sk[17]) & (i_13_) & (!i_14_) & (g107) & (!g91)) + ((i_12_) & (sk[17]) & (i_13_) & (i_14_) & (!g107) & (!g91)) + ((i_12_) & (sk[17]) & (i_13_) & (i_14_) & (!g107) & (g91)));
	assign g1268 = (((!g135) & (!g562) & (!g1029) & (sk[18]) & (!g1267)) + ((!g135) & (!g562) & (!g1029) & (sk[18]) & (g1267)) + ((!g135) & (!g562) & (g1029) & (!sk[18]) & (!g1267)) + ((!g135) & (!g562) & (g1029) & (!sk[18]) & (g1267)) + ((!g135) & (!g562) & (g1029) & (sk[18]) & (g1267)) + ((!g135) & (g562) & (!g1029) & (sk[18]) & (!g1267)) + ((!g135) & (g562) & (!g1029) & (sk[18]) & (g1267)) + ((!g135) & (g562) & (g1029) & (!sk[18]) & (!g1267)) + ((!g135) & (g562) & (g1029) & (!sk[18]) & (g1267)) + ((!g135) & (g562) & (g1029) & (sk[18]) & (!g1267)) + ((!g135) & (g562) & (g1029) & (sk[18]) & (g1267)) + ((g135) & (!g562) & (g1029) & (!sk[18]) & (!g1267)) + ((g135) & (!g562) & (g1029) & (!sk[18]) & (g1267)) + ((g135) & (g562) & (g1029) & (!sk[18]) & (!g1267)) + ((g135) & (g562) & (g1029) & (!sk[18]) & (g1267)));
	assign g1269 = (((!g159) & (!g964) & (g1007) & (!sk[19]) & (!g1268)) + ((!g159) & (!g964) & (g1007) & (!sk[19]) & (g1268)) + ((!g159) & (g964) & (g1007) & (!sk[19]) & (!g1268)) + ((!g159) & (g964) & (g1007) & (!sk[19]) & (g1268)) + ((!g159) & (g964) & (g1007) & (sk[19]) & (!g1268)) + ((g159) & (!g964) & (!g1007) & (sk[19]) & (!g1268)) + ((g159) & (!g964) & (g1007) & (!sk[19]) & (!g1268)) + ((g159) & (!g964) & (g1007) & (!sk[19]) & (g1268)) + ((g159) & (!g964) & (g1007) & (sk[19]) & (!g1268)) + ((g159) & (g964) & (!g1007) & (sk[19]) & (!g1268)) + ((g159) & (g964) & (g1007) & (!sk[19]) & (!g1268)) + ((g159) & (g964) & (g1007) & (!sk[19]) & (g1268)) + ((g159) & (g964) & (g1007) & (sk[19]) & (!g1268)));
	assign g1270 = (((!g973) & (!g1254) & (g1259) & (g1264) & (g1266) & (g1269)));
	assign g1271 = (((!i_4_) & (!i_3_) & (i_5_) & (!g43) & (!sk[21]) & (g71)) + ((!i_4_) & (!i_3_) & (i_5_) & (g43) & (!sk[21]) & (!g71)) + ((!i_4_) & (!i_3_) & (i_5_) & (g43) & (!sk[21]) & (g71)) + ((!i_4_) & (!i_3_) & (i_5_) & (g43) & (sk[21]) & (g71)) + ((!i_4_) & (i_3_) & (!i_5_) & (!g43) & (!sk[21]) & (!g71)) + ((!i_4_) & (i_3_) & (!i_5_) & (!g43) & (!sk[21]) & (g71)) + ((!i_4_) & (i_3_) & (!i_5_) & (g43) & (!sk[21]) & (!g71)) + ((!i_4_) & (i_3_) & (!i_5_) & (g43) & (!sk[21]) & (g71)) + ((!i_4_) & (i_3_) & (i_5_) & (!g43) & (!sk[21]) & (!g71)) + ((!i_4_) & (i_3_) & (i_5_) & (!g43) & (!sk[21]) & (g71)) + ((!i_4_) & (i_3_) & (i_5_) & (g43) & (!sk[21]) & (!g71)) + ((!i_4_) & (i_3_) & (i_5_) & (g43) & (!sk[21]) & (g71)) + ((i_4_) & (!i_3_) & (!i_5_) & (g43) & (sk[21]) & (g71)) + ((i_4_) & (!i_3_) & (i_5_) & (!g43) & (!sk[21]) & (g71)) + ((i_4_) & (!i_3_) & (i_5_) & (g43) & (!sk[21]) & (!g71)) + ((i_4_) & (!i_3_) & (i_5_) & (g43) & (!sk[21]) & (g71)) + ((i_4_) & (!i_3_) & (i_5_) & (g43) & (sk[21]) & (g71)) + ((i_4_) & (i_3_) & (!i_5_) & (!g43) & (!sk[21]) & (!g71)) + ((i_4_) & (i_3_) & (!i_5_) & (!g43) & (!sk[21]) & (g71)) + ((i_4_) & (i_3_) & (!i_5_) & (g43) & (!sk[21]) & (!g71)) + ((i_4_) & (i_3_) & (!i_5_) & (g43) & (!sk[21]) & (g71)) + ((i_4_) & (i_3_) & (i_5_) & (!g43) & (!sk[21]) & (!g71)) + ((i_4_) & (i_3_) & (i_5_) & (!g43) & (!sk[21]) & (g71)) + ((i_4_) & (i_3_) & (i_5_) & (g43) & (!sk[21]) & (!g71)) + ((i_4_) & (i_3_) & (i_5_) & (g43) & (!sk[21]) & (g71)));
	assign g1272 = (((!i_15_) & (!g429) & (g74) & (!g460) & (!sk[22]) & (g1271)) + ((!i_15_) & (!g429) & (g74) & (g460) & (!sk[22]) & (!g1271)) + ((!i_15_) & (!g429) & (g74) & (g460) & (!sk[22]) & (g1271)) + ((!i_15_) & (g429) & (!g74) & (!g460) & (!sk[22]) & (!g1271)) + ((!i_15_) & (g429) & (!g74) & (!g460) & (!sk[22]) & (g1271)) + ((!i_15_) & (g429) & (!g74) & (!g460) & (sk[22]) & (g1271)) + ((!i_15_) & (g429) & (!g74) & (g460) & (!sk[22]) & (!g1271)) + ((!i_15_) & (g429) & (!g74) & (g460) & (!sk[22]) & (g1271)) + ((!i_15_) & (g429) & (g74) & (!g460) & (!sk[22]) & (!g1271)) + ((!i_15_) & (g429) & (g74) & (!g460) & (!sk[22]) & (g1271)) + ((!i_15_) & (g429) & (g74) & (!g460) & (sk[22]) & (!g1271)) + ((!i_15_) & (g429) & (g74) & (!g460) & (sk[22]) & (g1271)) + ((!i_15_) & (g429) & (g74) & (g460) & (!sk[22]) & (!g1271)) + ((!i_15_) & (g429) & (g74) & (g460) & (!sk[22]) & (g1271)) + ((i_15_) & (!g429) & (g74) & (!g460) & (!sk[22]) & (g1271)) + ((i_15_) & (!g429) & (g74) & (g460) & (!sk[22]) & (!g1271)) + ((i_15_) & (!g429) & (g74) & (g460) & (!sk[22]) & (g1271)) + ((i_15_) & (g429) & (!g74) & (!g460) & (!sk[22]) & (!g1271)) + ((i_15_) & (g429) & (!g74) & (!g460) & (!sk[22]) & (g1271)) + ((i_15_) & (g429) & (!g74) & (g460) & (!sk[22]) & (!g1271)) + ((i_15_) & (g429) & (!g74) & (g460) & (!sk[22]) & (g1271)) + ((i_15_) & (g429) & (g74) & (!g460) & (!sk[22]) & (!g1271)) + ((i_15_) & (g429) & (g74) & (!g460) & (!sk[22]) & (g1271)) + ((i_15_) & (g429) & (g74) & (g460) & (!sk[22]) & (!g1271)) + ((i_15_) & (g429) & (g74) & (g460) & (!sk[22]) & (g1271)));
	assign g1273 = (((!i_12_) & (!sk[23]) & (!i_14_) & (g88) & (!g130)) + ((!i_12_) & (!sk[23]) & (!i_14_) & (g88) & (g130)) + ((!i_12_) & (!sk[23]) & (i_14_) & (g88) & (!g130)) + ((!i_12_) & (!sk[23]) & (i_14_) & (g88) & (g130)) + ((i_12_) & (!sk[23]) & (!i_14_) & (g88) & (!g130)) + ((i_12_) & (!sk[23]) & (!i_14_) & (g88) & (g130)) + ((i_12_) & (!sk[23]) & (i_14_) & (g88) & (!g130)) + ((i_12_) & (!sk[23]) & (i_14_) & (g88) & (g130)) + ((i_12_) & (sk[23]) & (!i_14_) & (g88) & (!g130)));
	assign g1274 = (((!g135) & (!g648) & (!sk[24]) & (g703) & (!g775)) + ((!g135) & (!g648) & (!sk[24]) & (g703) & (g775)) + ((!g135) & (!g648) & (sk[24]) & (g703) & (!g775)) + ((!g135) & (g648) & (!sk[24]) & (g703) & (!g775)) + ((!g135) & (g648) & (!sk[24]) & (g703) & (g775)) + ((g135) & (!g648) & (!sk[24]) & (g703) & (!g775)) + ((g135) & (!g648) & (!sk[24]) & (g703) & (g775)) + ((g135) & (!g648) & (sk[24]) & (!g703) & (!g775)) + ((g135) & (!g648) & (sk[24]) & (g703) & (!g775)) + ((g135) & (g648) & (!sk[24]) & (g703) & (!g775)) + ((g135) & (g648) & (!sk[24]) & (g703) & (g775)) + ((g135) & (g648) & (sk[24]) & (!g703) & (!g775)) + ((g135) & (g648) & (sk[24]) & (g703) & (!g775)));
	assign g1275 = (((!g74) & (!g104) & (!g847) & (sk[25]) & (!g1273) & (g1274)) + ((!g74) & (!g104) & (g847) & (!sk[25]) & (!g1273) & (g1274)) + ((!g74) & (!g104) & (g847) & (!sk[25]) & (g1273) & (!g1274)) + ((!g74) & (!g104) & (g847) & (!sk[25]) & (g1273) & (g1274)) + ((!g74) & (!g104) & (g847) & (sk[25]) & (!g1273) & (g1274)) + ((!g74) & (g104) & (!g847) & (!sk[25]) & (!g1273) & (!g1274)) + ((!g74) & (g104) & (!g847) & (!sk[25]) & (!g1273) & (g1274)) + ((!g74) & (g104) & (!g847) & (!sk[25]) & (g1273) & (!g1274)) + ((!g74) & (g104) & (!g847) & (!sk[25]) & (g1273) & (g1274)) + ((!g74) & (g104) & (g847) & (!sk[25]) & (!g1273) & (!g1274)) + ((!g74) & (g104) & (g847) & (!sk[25]) & (!g1273) & (g1274)) + ((!g74) & (g104) & (g847) & (!sk[25]) & (g1273) & (!g1274)) + ((!g74) & (g104) & (g847) & (!sk[25]) & (g1273) & (g1274)) + ((g74) & (!g104) & (g847) & (!sk[25]) & (!g1273) & (g1274)) + ((g74) & (!g104) & (g847) & (!sk[25]) & (g1273) & (!g1274)) + ((g74) & (!g104) & (g847) & (!sk[25]) & (g1273) & (g1274)) + ((g74) & (!g104) & (g847) & (sk[25]) & (!g1273) & (g1274)) + ((g74) & (g104) & (!g847) & (!sk[25]) & (!g1273) & (!g1274)) + ((g74) & (g104) & (!g847) & (!sk[25]) & (!g1273) & (g1274)) + ((g74) & (g104) & (!g847) & (!sk[25]) & (g1273) & (!g1274)) + ((g74) & (g104) & (!g847) & (!sk[25]) & (g1273) & (g1274)) + ((g74) & (g104) & (g847) & (!sk[25]) & (!g1273) & (!g1274)) + ((g74) & (g104) & (g847) & (!sk[25]) & (!g1273) & (g1274)) + ((g74) & (g104) & (g847) & (!sk[25]) & (g1273) & (!g1274)) + ((g74) & (g104) & (g847) & (!sk[25]) & (g1273) & (g1274)));
	assign g1276 = (((!sk[26]) & (!g313) & (!g348) & (g496) & (!g535)) + ((!sk[26]) & (!g313) & (!g348) & (g496) & (g535)) + ((!sk[26]) & (!g313) & (g348) & (g496) & (!g535)) + ((!sk[26]) & (!g313) & (g348) & (g496) & (g535)) + ((!sk[26]) & (g313) & (!g348) & (g496) & (!g535)) + ((!sk[26]) & (g313) & (!g348) & (g496) & (g535)) + ((!sk[26]) & (g313) & (g348) & (g496) & (!g535)) + ((!sk[26]) & (g313) & (g348) & (g496) & (g535)) + ((sk[26]) & (!g313) & (!g348) & (!g496) & (!g535)) + ((sk[26]) & (!g313) & (g348) & (!g496) & (!g535)) + ((sk[26]) & (!g313) & (g348) & (g496) & (!g535)) + ((sk[26]) & (g313) & (!g348) & (!g496) & (!g535)) + ((sk[26]) & (g313) & (g348) & (!g496) & (!g535)));
	assign g1277 = (((!g413) & (!g522) & (g847) & (!sk[27]) & (!g1276)) + ((!g413) & (!g522) & (g847) & (!sk[27]) & (g1276)) + ((!g413) & (!g522) & (g847) & (sk[27]) & (g1276)) + ((!g413) & (g522) & (g847) & (!sk[27]) & (!g1276)) + ((!g413) & (g522) & (g847) & (!sk[27]) & (g1276)) + ((g413) & (!g522) & (!g847) & (sk[27]) & (g1276)) + ((g413) & (!g522) & (g847) & (!sk[27]) & (!g1276)) + ((g413) & (!g522) & (g847) & (!sk[27]) & (g1276)) + ((g413) & (!g522) & (g847) & (sk[27]) & (g1276)) + ((g413) & (g522) & (!g847) & (sk[27]) & (g1276)) + ((g413) & (g522) & (g847) & (!sk[27]) & (!g1276)) + ((g413) & (g522) & (g847) & (!sk[27]) & (g1276)) + ((g413) & (g522) & (g847) & (sk[27]) & (g1276)));
	assign g1278 = (((!sk[28]) & (!g135) & (!g191) & (g187)) + ((!sk[28]) & (!g135) & (g191) & (!g187)) + ((!sk[28]) & (!g135) & (g191) & (g187)) + ((!sk[28]) & (g135) & (!g191) & (g187)) + ((!sk[28]) & (g135) & (g191) & (!g187)) + ((!sk[28]) & (g135) & (g191) & (g187)) + ((sk[28]) & (!g135) & (!g191) & (g187)) + ((sk[28]) & (!g135) & (g191) & (!g187)) + ((sk[28]) & (!g135) & (g191) & (g187)));
	assign g1279 = (((!sk[29]) & (!g102) & (!g534) & (g500) & (!g703)) + ((!sk[29]) & (!g102) & (!g534) & (g500) & (g703)) + ((!sk[29]) & (!g102) & (g534) & (g500) & (!g703)) + ((!sk[29]) & (!g102) & (g534) & (g500) & (g703)) + ((!sk[29]) & (g102) & (!g534) & (g500) & (!g703)) + ((!sk[29]) & (g102) & (!g534) & (g500) & (g703)) + ((!sk[29]) & (g102) & (g534) & (g500) & (!g703)) + ((!sk[29]) & (g102) & (g534) & (g500) & (g703)) + ((sk[29]) & (g102) & (!g534) & (!g500) & (!g703)) + ((sk[29]) & (g102) & (!g534) & (g500) & (!g703)) + ((sk[29]) & (g102) & (!g534) & (g500) & (g703)) + ((sk[29]) & (g102) & (g534) & (!g500) & (!g703)) + ((sk[29]) & (g102) & (g534) & (!g500) & (g703)) + ((sk[29]) & (g102) & (g534) & (g500) & (!g703)) + ((sk[29]) & (g102) & (g534) & (g500) & (g703)));
	assign g1280 = (((!g135) & (!g89) & (!sk[30]) & (g630)) + ((!g135) & (!g89) & (sk[30]) & (!g630)) + ((!g135) & (!g89) & (sk[30]) & (g630)) + ((!g135) & (g89) & (!sk[30]) & (!g630)) + ((!g135) & (g89) & (!sk[30]) & (g630)) + ((!g135) & (g89) & (sk[30]) & (g630)) + ((g135) & (!g89) & (!sk[30]) & (g630)) + ((g135) & (g89) & (!sk[30]) & (!g630)) + ((g135) & (g89) & (!sk[30]) & (g630)));
	assign g1281 = (((!i_12_) & (!i_13_) & (i_14_) & (!sk[31]) & (!g86) & (g102)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[31]) & (g86) & (!g102)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[31]) & (g86) & (g102)) + ((!i_12_) & (!i_13_) & (i_14_) & (sk[31]) & (g86) & (g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[31]) & (!g86) & (!g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[31]) & (!g86) & (g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[31]) & (g86) & (!g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[31]) & (g86) & (g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (sk[31]) & (g86) & (g102)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[31]) & (!g86) & (!g102)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[31]) & (!g86) & (g102)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[31]) & (g86) & (!g102)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[31]) & (g86) & (g102)) + ((i_12_) & (!i_13_) & (!i_14_) & (sk[31]) & (g86) & (g102)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[31]) & (!g86) & (g102)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[31]) & (g86) & (!g102)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[31]) & (g86) & (g102)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[31]) & (!g86) & (!g102)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[31]) & (!g86) & (g102)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[31]) & (g86) & (!g102)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[31]) & (g86) & (g102)) + ((i_12_) & (i_13_) & (!i_14_) & (sk[31]) & (g86) & (g102)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[31]) & (!g86) & (!g102)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[31]) & (!g86) & (g102)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[31]) & (g86) & (!g102)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[31]) & (g86) & (g102)) + ((i_12_) & (i_13_) & (i_14_) & (sk[31]) & (g86) & (g102)));
	assign g1282 = (((!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g429) & (!g131)) + ((!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g429) & (!g131)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g429) & (!g131)) + ((!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g429) & (!g131)) + ((i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (g429) & (!g131)) + ((i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g429) & (!g131)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g429) & (!g131)) + ((i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g429) & (!g131)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g429) & (!g131)));
	assign g1283 = (((!sk[33]) & (!g1278) & (!g1279) & (g1280) & (!g1281) & (g1282)) + ((!sk[33]) & (!g1278) & (!g1279) & (g1280) & (g1281) & (!g1282)) + ((!sk[33]) & (!g1278) & (!g1279) & (g1280) & (g1281) & (g1282)) + ((!sk[33]) & (!g1278) & (g1279) & (!g1280) & (!g1281) & (!g1282)) + ((!sk[33]) & (!g1278) & (g1279) & (!g1280) & (!g1281) & (g1282)) + ((!sk[33]) & (!g1278) & (g1279) & (!g1280) & (g1281) & (!g1282)) + ((!sk[33]) & (!g1278) & (g1279) & (!g1280) & (g1281) & (g1282)) + ((!sk[33]) & (!g1278) & (g1279) & (g1280) & (!g1281) & (!g1282)) + ((!sk[33]) & (!g1278) & (g1279) & (g1280) & (!g1281) & (g1282)) + ((!sk[33]) & (!g1278) & (g1279) & (g1280) & (g1281) & (!g1282)) + ((!sk[33]) & (!g1278) & (g1279) & (g1280) & (g1281) & (g1282)) + ((!sk[33]) & (g1278) & (!g1279) & (g1280) & (!g1281) & (g1282)) + ((!sk[33]) & (g1278) & (!g1279) & (g1280) & (g1281) & (!g1282)) + ((!sk[33]) & (g1278) & (!g1279) & (g1280) & (g1281) & (g1282)) + ((!sk[33]) & (g1278) & (g1279) & (!g1280) & (!g1281) & (!g1282)) + ((!sk[33]) & (g1278) & (g1279) & (!g1280) & (!g1281) & (g1282)) + ((!sk[33]) & (g1278) & (g1279) & (!g1280) & (g1281) & (!g1282)) + ((!sk[33]) & (g1278) & (g1279) & (!g1280) & (g1281) & (g1282)) + ((!sk[33]) & (g1278) & (g1279) & (g1280) & (!g1281) & (!g1282)) + ((!sk[33]) & (g1278) & (g1279) & (g1280) & (!g1281) & (g1282)) + ((!sk[33]) & (g1278) & (g1279) & (g1280) & (g1281) & (!g1282)) + ((!sk[33]) & (g1278) & (g1279) & (g1280) & (g1281) & (g1282)) + ((sk[33]) & (!g1278) & (!g1279) & (!g1280) & (!g1281) & (!g1282)));
	assign g1284 = (((!g135) & (!sk[34]) & (!g131) & (g273) & (!g342)) + ((!g135) & (!sk[34]) & (!g131) & (g273) & (g342)) + ((!g135) & (!sk[34]) & (g131) & (g273) & (!g342)) + ((!g135) & (!sk[34]) & (g131) & (g273) & (g342)) + ((!g135) & (sk[34]) & (!g131) & (!g273) & (!g342)) + ((!g135) & (sk[34]) & (g131) & (!g273) & (!g342)) + ((g135) & (!sk[34]) & (!g131) & (g273) & (!g342)) + ((g135) & (!sk[34]) & (!g131) & (g273) & (g342)) + ((g135) & (!sk[34]) & (g131) & (g273) & (!g342)) + ((g135) & (!sk[34]) & (g131) & (g273) & (g342)) + ((g135) & (sk[34]) & (!g131) & (!g273) & (!g342)) + ((g135) & (sk[34]) & (!g131) & (g273) & (!g342)) + ((g135) & (sk[34]) & (g131) & (!g273) & (!g342)) + ((g135) & (sk[34]) & (g131) & (!g273) & (g342)) + ((g135) & (sk[34]) & (g131) & (g273) & (!g342)) + ((g135) & (sk[34]) & (g131) & (g273) & (g342)));
	assign g1285 = (((!g159) & (!g253) & (g336) & (!g500) & (!g627) & (g848)) + ((!g159) & (g253) & (!g336) & (!g500) & (!g627) & (!g848)) + ((!g159) & (g253) & (!g336) & (!g500) & (!g627) & (g848)) + ((!g159) & (g253) & (!g336) & (!g500) & (g627) & (!g848)) + ((!g159) & (g253) & (!g336) & (!g500) & (g627) & (g848)) + ((!g159) & (g253) & (g336) & (!g500) & (!g627) & (!g848)) + ((!g159) & (g253) & (g336) & (!g500) & (!g627) & (g848)) + ((!g159) & (g253) & (g336) & (!g500) & (g627) & (!g848)) + ((!g159) & (g253) & (g336) & (!g500) & (g627) & (g848)) + ((g159) & (!g253) & (g336) & (!g500) & (!g627) & (g848)) + ((g159) & (g253) & (!g336) & (!g500) & (!g627) & (!g848)) + ((g159) & (g253) & (!g336) & (!g500) & (!g627) & (g848)) + ((g159) & (g253) & (!g336) & (!g500) & (g627) & (!g848)) + ((g159) & (g253) & (!g336) & (!g500) & (g627) & (g848)) + ((g159) & (g253) & (!g336) & (g500) & (!g627) & (!g848)) + ((g159) & (g253) & (!g336) & (g500) & (!g627) & (g848)) + ((g159) & (g253) & (!g336) & (g500) & (g627) & (!g848)) + ((g159) & (g253) & (!g336) & (g500) & (g627) & (g848)) + ((g159) & (g253) & (g336) & (!g500) & (!g627) & (!g848)) + ((g159) & (g253) & (g336) & (!g500) & (!g627) & (g848)) + ((g159) & (g253) & (g336) & (!g500) & (g627) & (!g848)) + ((g159) & (g253) & (g336) & (!g500) & (g627) & (g848)) + ((g159) & (g253) & (g336) & (g500) & (!g627) & (!g848)) + ((g159) & (g253) & (g336) & (g500) & (!g627) & (g848)) + ((g159) & (g253) & (g336) & (g500) & (g627) & (!g848)) + ((g159) & (g253) & (g336) & (g500) & (g627) & (g848)));
	assign g1286 = (((!g274) & (!sk[36]) & (!g584) & (g1284) & (!g1285)) + ((!g274) & (!sk[36]) & (!g584) & (g1284) & (g1285)) + ((!g274) & (!sk[36]) & (g584) & (g1284) & (!g1285)) + ((!g274) & (!sk[36]) & (g584) & (g1284) & (g1285)) + ((!g274) & (sk[36]) & (!g584) & (g1284) & (g1285)) + ((g274) & (!sk[36]) & (!g584) & (g1284) & (!g1285)) + ((g274) & (!sk[36]) & (!g584) & (g1284) & (g1285)) + ((g274) & (!sk[36]) & (g584) & (g1284) & (!g1285)) + ((g274) & (!sk[36]) & (g584) & (g1284) & (g1285)));
	assign g1287 = (((!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g429) & (!g130)) + ((!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g429) & (!g130)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g429) & (!g130)) + ((!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g429) & (!g130)) + ((!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g429) & (!g130)) + ((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g429) & (!g130)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g429) & (!g130)) + ((i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (g429) & (!g130)) + ((i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g429) & (!g130)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g429) & (!g130)) + ((i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g429) & (!g130)));
	assign g1288 = (((!g76) & (!g157) & (!g135) & (sk[38]) & (g88) & (!g176)) + ((!g76) & (!g157) & (!g135) & (sk[38]) & (g88) & (g176)) + ((!g76) & (!g157) & (g135) & (!sk[38]) & (!g88) & (g176)) + ((!g76) & (!g157) & (g135) & (!sk[38]) & (g88) & (!g176)) + ((!g76) & (!g157) & (g135) & (!sk[38]) & (g88) & (g176)) + ((!g76) & (g157) & (!g135) & (!sk[38]) & (!g88) & (!g176)) + ((!g76) & (g157) & (!g135) & (!sk[38]) & (!g88) & (g176)) + ((!g76) & (g157) & (!g135) & (!sk[38]) & (g88) & (!g176)) + ((!g76) & (g157) & (!g135) & (!sk[38]) & (g88) & (g176)) + ((!g76) & (g157) & (!g135) & (sk[38]) & (g88) & (!g176)) + ((!g76) & (g157) & (!g135) & (sk[38]) & (g88) & (g176)) + ((!g76) & (g157) & (g135) & (!sk[38]) & (!g88) & (!g176)) + ((!g76) & (g157) & (g135) & (!sk[38]) & (!g88) & (g176)) + ((!g76) & (g157) & (g135) & (!sk[38]) & (g88) & (!g176)) + ((!g76) & (g157) & (g135) & (!sk[38]) & (g88) & (g176)) + ((!g76) & (g157) & (g135) & (sk[38]) & (g88) & (!g176)) + ((!g76) & (g157) & (g135) & (sk[38]) & (g88) & (g176)) + ((g76) & (!g157) & (g135) & (!sk[38]) & (!g88) & (g176)) + ((g76) & (!g157) & (g135) & (!sk[38]) & (g88) & (!g176)) + ((g76) & (!g157) & (g135) & (!sk[38]) & (g88) & (g176)) + ((g76) & (g157) & (!g135) & (!sk[38]) & (!g88) & (!g176)) + ((g76) & (g157) & (!g135) & (!sk[38]) & (!g88) & (g176)) + ((g76) & (g157) & (!g135) & (!sk[38]) & (g88) & (!g176)) + ((g76) & (g157) & (!g135) & (!sk[38]) & (g88) & (g176)) + ((g76) & (g157) & (!g135) & (sk[38]) & (g88) & (!g176)) + ((g76) & (g157) & (g135) & (!sk[38]) & (!g88) & (!g176)) + ((g76) & (g157) & (g135) & (!sk[38]) & (!g88) & (g176)) + ((g76) & (g157) & (g135) & (!sk[38]) & (g88) & (!g176)) + ((g76) & (g157) & (g135) & (!sk[38]) & (g88) & (g176)) + ((g76) & (g157) & (g135) & (sk[38]) & (g88) & (!g176)));
	assign g1289 = (((!i_8_) & (!i_6_) & (i_7_) & (!g429) & (!sk[39]) & (g394)) + ((!i_8_) & (!i_6_) & (i_7_) & (g429) & (!sk[39]) & (!g394)) + ((!i_8_) & (!i_6_) & (i_7_) & (g429) & (!sk[39]) & (g394)) + ((!i_8_) & (!i_6_) & (i_7_) & (g429) & (sk[39]) & (g394)) + ((!i_8_) & (i_6_) & (!i_7_) & (!g429) & (!sk[39]) & (!g394)) + ((!i_8_) & (i_6_) & (!i_7_) & (!g429) & (!sk[39]) & (g394)) + ((!i_8_) & (i_6_) & (!i_7_) & (g429) & (!sk[39]) & (!g394)) + ((!i_8_) & (i_6_) & (!i_7_) & (g429) & (!sk[39]) & (g394)) + ((!i_8_) & (i_6_) & (!i_7_) & (g429) & (sk[39]) & (g394)) + ((!i_8_) & (i_6_) & (i_7_) & (!g429) & (!sk[39]) & (!g394)) + ((!i_8_) & (i_6_) & (i_7_) & (!g429) & (!sk[39]) & (g394)) + ((!i_8_) & (i_6_) & (i_7_) & (g429) & (!sk[39]) & (!g394)) + ((!i_8_) & (i_6_) & (i_7_) & (g429) & (!sk[39]) & (g394)) + ((!i_8_) & (i_6_) & (i_7_) & (g429) & (sk[39]) & (g394)) + ((i_8_) & (!i_6_) & (i_7_) & (!g429) & (!sk[39]) & (g394)) + ((i_8_) & (!i_6_) & (i_7_) & (g429) & (!sk[39]) & (!g394)) + ((i_8_) & (!i_6_) & (i_7_) & (g429) & (!sk[39]) & (g394)) + ((i_8_) & (i_6_) & (!i_7_) & (!g429) & (!sk[39]) & (!g394)) + ((i_8_) & (i_6_) & (!i_7_) & (!g429) & (!sk[39]) & (g394)) + ((i_8_) & (i_6_) & (!i_7_) & (g429) & (!sk[39]) & (!g394)) + ((i_8_) & (i_6_) & (!i_7_) & (g429) & (!sk[39]) & (g394)) + ((i_8_) & (i_6_) & (i_7_) & (!g429) & (!sk[39]) & (!g394)) + ((i_8_) & (i_6_) & (i_7_) & (!g429) & (!sk[39]) & (g394)) + ((i_8_) & (i_6_) & (i_7_) & (g429) & (!sk[39]) & (!g394)) + ((i_8_) & (i_6_) & (i_7_) & (g429) & (!sk[39]) & (g394)));
	assign g1290 = (((!g206) & (!g1287) & (!g1288) & (sk[40]) & (!g1289)) + ((!g206) & (!g1287) & (g1288) & (!sk[40]) & (!g1289)) + ((!g206) & (!g1287) & (g1288) & (!sk[40]) & (g1289)) + ((!g206) & (g1287) & (g1288) & (!sk[40]) & (!g1289)) + ((!g206) & (g1287) & (g1288) & (!sk[40]) & (g1289)) + ((g206) & (!g1287) & (g1288) & (!sk[40]) & (!g1289)) + ((g206) & (!g1287) & (g1288) & (!sk[40]) & (g1289)) + ((g206) & (g1287) & (g1288) & (!sk[40]) & (!g1289)) + ((g206) & (g1287) & (g1288) & (!sk[40]) & (g1289)));
	assign g1291 = (((!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g429) & (g74)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g429) & (g74)) + ((!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g429) & (g74)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g429) & (g74)) + ((i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (g429) & (g74)) + ((i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g429) & (g74)) + ((i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g429) & (g74)) + ((i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g429) & (g74)) + ((i_15_) & (i_12_) & (i_13_) & (i_14_) & (g429) & (g74)));
	assign g1292 = (((!g102) & (!g253) & (!sk[42]) & (g342) & (!g630)) + ((!g102) & (!g253) & (!sk[42]) & (g342) & (g630)) + ((!g102) & (!g253) & (sk[42]) & (!g342) & (!g630)) + ((!g102) & (g253) & (!sk[42]) & (g342) & (!g630)) + ((!g102) & (g253) & (!sk[42]) & (g342) & (g630)) + ((!g102) & (g253) & (sk[42]) & (!g342) & (!g630)) + ((!g102) & (g253) & (sk[42]) & (!g342) & (g630)) + ((!g102) & (g253) & (sk[42]) & (g342) & (!g630)) + ((!g102) & (g253) & (sk[42]) & (g342) & (g630)) + ((g102) & (!g253) & (!sk[42]) & (g342) & (!g630)) + ((g102) & (!g253) & (!sk[42]) & (g342) & (g630)) + ((g102) & (!g253) & (sk[42]) & (!g342) & (!g630)) + ((g102) & (g253) & (!sk[42]) & (g342) & (!g630)) + ((g102) & (g253) & (!sk[42]) & (g342) & (g630)) + ((g102) & (g253) & (sk[42]) & (!g342) & (!g630)));
	assign g1293 = (((!g159) & (!sk[43]) & (!g847) & (g934) & (!g975) & (g1292)) + ((!g159) & (!sk[43]) & (!g847) & (g934) & (g975) & (!g1292)) + ((!g159) & (!sk[43]) & (!g847) & (g934) & (g975) & (g1292)) + ((!g159) & (!sk[43]) & (g847) & (!g934) & (!g975) & (!g1292)) + ((!g159) & (!sk[43]) & (g847) & (!g934) & (!g975) & (g1292)) + ((!g159) & (!sk[43]) & (g847) & (!g934) & (g975) & (!g1292)) + ((!g159) & (!sk[43]) & (g847) & (!g934) & (g975) & (g1292)) + ((!g159) & (!sk[43]) & (g847) & (g934) & (!g975) & (!g1292)) + ((!g159) & (!sk[43]) & (g847) & (g934) & (!g975) & (g1292)) + ((!g159) & (!sk[43]) & (g847) & (g934) & (g975) & (!g1292)) + ((!g159) & (!sk[43]) & (g847) & (g934) & (g975) & (g1292)) + ((!g159) & (sk[43]) & (g847) & (g934) & (g975) & (g1292)) + ((g159) & (!sk[43]) & (!g847) & (g934) & (!g975) & (g1292)) + ((g159) & (!sk[43]) & (!g847) & (g934) & (g975) & (!g1292)) + ((g159) & (!sk[43]) & (!g847) & (g934) & (g975) & (g1292)) + ((g159) & (!sk[43]) & (g847) & (!g934) & (!g975) & (!g1292)) + ((g159) & (!sk[43]) & (g847) & (!g934) & (!g975) & (g1292)) + ((g159) & (!sk[43]) & (g847) & (!g934) & (g975) & (!g1292)) + ((g159) & (!sk[43]) & (g847) & (!g934) & (g975) & (g1292)) + ((g159) & (!sk[43]) & (g847) & (g934) & (!g975) & (!g1292)) + ((g159) & (!sk[43]) & (g847) & (g934) & (!g975) & (g1292)) + ((g159) & (!sk[43]) & (g847) & (g934) & (g975) & (!g1292)) + ((g159) & (!sk[43]) & (g847) & (g934) & (g975) & (g1292)) + ((g159) & (sk[43]) & (!g847) & (!g934) & (!g975) & (g1292)) + ((g159) & (sk[43]) & (!g847) & (!g934) & (g975) & (g1292)) + ((g159) & (sk[43]) & (!g847) & (g934) & (!g975) & (g1292)) + ((g159) & (sk[43]) & (!g847) & (g934) & (g975) & (g1292)) + ((g159) & (sk[43]) & (g847) & (!g934) & (!g975) & (g1292)) + ((g159) & (sk[43]) & (g847) & (!g934) & (g975) & (g1292)) + ((g159) & (sk[43]) & (g847) & (g934) & (!g975) & (g1292)) + ((g159) & (sk[43]) & (g847) & (g934) & (g975) & (g1292)));
	assign g1294 = (((!g1283) & (!g1286) & (g1290) & (!sk[44]) & (!g1291) & (g1293)) + ((!g1283) & (!g1286) & (g1290) & (!sk[44]) & (g1291) & (!g1293)) + ((!g1283) & (!g1286) & (g1290) & (!sk[44]) & (g1291) & (g1293)) + ((!g1283) & (g1286) & (!g1290) & (!sk[44]) & (!g1291) & (!g1293)) + ((!g1283) & (g1286) & (!g1290) & (!sk[44]) & (!g1291) & (g1293)) + ((!g1283) & (g1286) & (!g1290) & (!sk[44]) & (g1291) & (!g1293)) + ((!g1283) & (g1286) & (!g1290) & (!sk[44]) & (g1291) & (g1293)) + ((!g1283) & (g1286) & (g1290) & (!sk[44]) & (!g1291) & (!g1293)) + ((!g1283) & (g1286) & (g1290) & (!sk[44]) & (!g1291) & (g1293)) + ((!g1283) & (g1286) & (g1290) & (!sk[44]) & (g1291) & (!g1293)) + ((!g1283) & (g1286) & (g1290) & (!sk[44]) & (g1291) & (g1293)) + ((g1283) & (!g1286) & (g1290) & (!sk[44]) & (!g1291) & (g1293)) + ((g1283) & (!g1286) & (g1290) & (!sk[44]) & (g1291) & (!g1293)) + ((g1283) & (!g1286) & (g1290) & (!sk[44]) & (g1291) & (g1293)) + ((g1283) & (g1286) & (!g1290) & (!sk[44]) & (!g1291) & (!g1293)) + ((g1283) & (g1286) & (!g1290) & (!sk[44]) & (!g1291) & (g1293)) + ((g1283) & (g1286) & (!g1290) & (!sk[44]) & (g1291) & (!g1293)) + ((g1283) & (g1286) & (!g1290) & (!sk[44]) & (g1291) & (g1293)) + ((g1283) & (g1286) & (g1290) & (!sk[44]) & (!g1291) & (!g1293)) + ((g1283) & (g1286) & (g1290) & (!sk[44]) & (!g1291) & (g1293)) + ((g1283) & (g1286) & (g1290) & (!sk[44]) & (g1291) & (!g1293)) + ((g1283) & (g1286) & (g1290) & (!sk[44]) & (g1291) & (g1293)) + ((g1283) & (g1286) & (g1290) & (sk[44]) & (!g1291) & (g1293)));
	assign g1295 = (((!g1270) & (!g1272) & (!sk[45]) & (g1275) & (!g1277) & (g1294)) + ((!g1270) & (!g1272) & (!sk[45]) & (g1275) & (g1277) & (!g1294)) + ((!g1270) & (!g1272) & (!sk[45]) & (g1275) & (g1277) & (g1294)) + ((!g1270) & (g1272) & (!sk[45]) & (!g1275) & (!g1277) & (!g1294)) + ((!g1270) & (g1272) & (!sk[45]) & (!g1275) & (!g1277) & (g1294)) + ((!g1270) & (g1272) & (!sk[45]) & (!g1275) & (g1277) & (!g1294)) + ((!g1270) & (g1272) & (!sk[45]) & (!g1275) & (g1277) & (g1294)) + ((!g1270) & (g1272) & (!sk[45]) & (g1275) & (!g1277) & (!g1294)) + ((!g1270) & (g1272) & (!sk[45]) & (g1275) & (!g1277) & (g1294)) + ((!g1270) & (g1272) & (!sk[45]) & (g1275) & (g1277) & (!g1294)) + ((!g1270) & (g1272) & (!sk[45]) & (g1275) & (g1277) & (g1294)) + ((g1270) & (!g1272) & (!sk[45]) & (g1275) & (!g1277) & (g1294)) + ((g1270) & (!g1272) & (!sk[45]) & (g1275) & (g1277) & (!g1294)) + ((g1270) & (!g1272) & (!sk[45]) & (g1275) & (g1277) & (g1294)) + ((g1270) & (!g1272) & (sk[45]) & (g1275) & (g1277) & (g1294)) + ((g1270) & (g1272) & (!sk[45]) & (!g1275) & (!g1277) & (!g1294)) + ((g1270) & (g1272) & (!sk[45]) & (!g1275) & (!g1277) & (g1294)) + ((g1270) & (g1272) & (!sk[45]) & (!g1275) & (g1277) & (!g1294)) + ((g1270) & (g1272) & (!sk[45]) & (!g1275) & (g1277) & (g1294)) + ((g1270) & (g1272) & (!sk[45]) & (g1275) & (!g1277) & (!g1294)) + ((g1270) & (g1272) & (!sk[45]) & (g1275) & (!g1277) & (g1294)) + ((g1270) & (g1272) & (!sk[45]) & (g1275) & (g1277) & (!g1294)) + ((g1270) & (g1272) & (!sk[45]) & (g1275) & (g1277) & (g1294)));
	assign g1296 = (((!i_12_) & (!i_13_) & (!i_14_) & (!g35) & (g36) & (!g130)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g35) & (g36) & (!g130)) + ((!i_12_) & (!i_13_) & (i_14_) & (g35) & (!g36) & (!g130)) + ((!i_12_) & (!i_13_) & (i_14_) & (g35) & (g36) & (!g130)) + ((!i_12_) & (i_13_) & (!i_14_) & (g35) & (!g36) & (!g130)) + ((!i_12_) & (i_13_) & (!i_14_) & (g35) & (g36) & (!g130)) + ((!i_12_) & (i_13_) & (i_14_) & (!g35) & (g36) & (!g130)) + ((!i_12_) & (i_13_) & (i_14_) & (g35) & (!g36) & (!g130)) + ((!i_12_) & (i_13_) & (i_14_) & (g35) & (g36) & (!g130)) + ((i_12_) & (!i_13_) & (!i_14_) & (!g35) & (g36) & (!g130)) + ((i_12_) & (!i_13_) & (!i_14_) & (g35) & (!g36) & (!g130)) + ((i_12_) & (!i_13_) & (!i_14_) & (g35) & (g36) & (!g130)) + ((i_12_) & (!i_13_) & (i_14_) & (!g35) & (g36) & (!g130)) + ((i_12_) & (!i_13_) & (i_14_) & (g35) & (g36) & (!g130)) + ((i_12_) & (i_13_) & (!i_14_) & (!g35) & (g36) & (!g130)) + ((i_12_) & (i_13_) & (!i_14_) & (g35) & (!g36) & (!g130)) + ((i_12_) & (i_13_) & (!i_14_) & (g35) & (g36) & (!g130)) + ((i_12_) & (i_13_) & (i_14_) & (g35) & (!g36) & (!g130)) + ((i_12_) & (i_13_) & (i_14_) & (g35) & (g36) & (!g130)));
	assign g1297 = (((!g135) & (!g130) & (!g337) & (!g635) & (g851) & (!g1296)) + ((!g135) & (g130) & (!g337) & (!g635) & (!g851) & (!g1296)) + ((!g135) & (g130) & (!g337) & (!g635) & (g851) & (!g1296)) + ((g135) & (!g130) & (!g337) & (!g635) & (g851) & (!g1296)) + ((g135) & (g130) & (!g337) & (!g635) & (!g851) & (!g1296)) + ((g135) & (g130) & (!g337) & (!g635) & (g851) & (!g1296)) + ((g135) & (g130) & (!g337) & (g635) & (!g851) & (!g1296)) + ((g135) & (g130) & (!g337) & (g635) & (g851) & (!g1296)) + ((g135) & (g130) & (g337) & (!g635) & (!g851) & (!g1296)) + ((g135) & (g130) & (g337) & (!g635) & (g851) & (!g1296)) + ((g135) & (g130) & (g337) & (g635) & (!g851) & (!g1296)) + ((g135) & (g130) & (g337) & (g635) & (g851) & (!g1296)));
	assign g1298 = (((!g157) & (!sk[48]) & (!g135) & (g186) & (!g337)) + ((!g157) & (!sk[48]) & (!g135) & (g186) & (g337)) + ((!g157) & (!sk[48]) & (g135) & (g186) & (!g337)) + ((!g157) & (!sk[48]) & (g135) & (g186) & (g337)) + ((!g157) & (sk[48]) & (!g135) & (g186) & (!g337)) + ((!g157) & (sk[48]) & (!g135) & (g186) & (g337)) + ((g157) & (!sk[48]) & (!g135) & (g186) & (!g337)) + ((g157) & (!sk[48]) & (!g135) & (g186) & (g337)) + ((g157) & (!sk[48]) & (g135) & (g186) & (!g337)) + ((g157) & (!sk[48]) & (g135) & (g186) & (g337)) + ((g157) & (sk[48]) & (!g135) & (!g186) & (g337)) + ((g157) & (sk[48]) & (!g135) & (g186) & (!g337)) + ((g157) & (sk[48]) & (!g135) & (g186) & (g337)) + ((g157) & (sk[48]) & (g135) & (!g186) & (g337)) + ((g157) & (sk[48]) & (g135) & (g186) & (g337)));
	assign g1299 = (((!g109) & (!sk[49]) & (!g90) & (g102)) + ((!g109) & (!sk[49]) & (g90) & (!g102)) + ((!g109) & (!sk[49]) & (g90) & (g102)) + ((!g109) & (sk[49]) & (g90) & (g102)) + ((g109) & (!sk[49]) & (!g90) & (g102)) + ((g109) & (!sk[49]) & (g90) & (!g102)) + ((g109) & (!sk[49]) & (g90) & (g102)) + ((g109) & (sk[49]) & (!g90) & (g102)) + ((g109) & (sk[49]) & (g90) & (g102)));
	assign g1300 = (((!g35) & (!g157) & (!sk[50]) & (g460)) + ((!g35) & (!g157) & (sk[50]) & (!g460)) + ((!g35) & (!g157) & (sk[50]) & (g460)) + ((!g35) & (g157) & (!sk[50]) & (!g460)) + ((!g35) & (g157) & (!sk[50]) & (g460)) + ((g35) & (!g157) & (!sk[50]) & (g460)) + ((g35) & (!g157) & (sk[50]) & (g460)) + ((g35) & (g157) & (!sk[50]) & (!g460)) + ((g35) & (g157) & (!sk[50]) & (g460)));
	assign g1301 = (((!i_12_) & (!i_14_) & (!sk[51]) & (g35) & (!g72)) + ((!i_12_) & (!i_14_) & (!sk[51]) & (g35) & (g72)) + ((!i_12_) & (i_14_) & (!sk[51]) & (g35) & (!g72)) + ((!i_12_) & (i_14_) & (!sk[51]) & (g35) & (g72)) + ((i_12_) & (!i_14_) & (!sk[51]) & (g35) & (!g72)) + ((i_12_) & (!i_14_) & (!sk[51]) & (g35) & (g72)) + ((i_12_) & (!i_14_) & (sk[51]) & (g35) & (g72)) + ((i_12_) & (i_14_) & (!sk[51]) & (g35) & (!g72)) + ((i_12_) & (i_14_) & (!sk[51]) & (g35) & (g72)));
	assign g1302 = (((!i_8_) & (!sk[52]) & (!i_6_) & (i_7_) & (!g1301)) + ((!i_8_) & (!sk[52]) & (!i_6_) & (i_7_) & (g1301)) + ((!i_8_) & (!sk[52]) & (i_6_) & (i_7_) & (!g1301)) + ((!i_8_) & (!sk[52]) & (i_6_) & (i_7_) & (g1301)) + ((!i_8_) & (sk[52]) & (!i_6_) & (i_7_) & (g1301)) + ((!i_8_) & (sk[52]) & (i_6_) & (!i_7_) & (g1301)) + ((i_8_) & (!sk[52]) & (!i_6_) & (i_7_) & (!g1301)) + ((i_8_) & (!sk[52]) & (!i_6_) & (i_7_) & (g1301)) + ((i_8_) & (!sk[52]) & (i_6_) & (i_7_) & (!g1301)) + ((i_8_) & (!sk[52]) & (i_6_) & (i_7_) & (g1301)));
	assign g1303 = (((!g74) & (!g1299) & (!g281) & (!g1300) & (sk[53]) & (!g1302)) + ((!g74) & (!g1299) & (!g281) & (!g1300) & (sk[53]) & (g1302)) + ((!g74) & (!g1299) & (!g281) & (g1300) & (sk[53]) & (!g1302)) + ((!g74) & (!g1299) & (!g281) & (g1300) & (sk[53]) & (g1302)) + ((!g74) & (!g1299) & (g281) & (!g1300) & (!sk[53]) & (g1302)) + ((!g74) & (!g1299) & (g281) & (!g1300) & (sk[53]) & (!g1302)) + ((!g74) & (!g1299) & (g281) & (g1300) & (!sk[53]) & (!g1302)) + ((!g74) & (!g1299) & (g281) & (g1300) & (!sk[53]) & (g1302)) + ((!g74) & (!g1299) & (g281) & (g1300) & (sk[53]) & (!g1302)) + ((!g74) & (!g1299) & (g281) & (g1300) & (sk[53]) & (g1302)) + ((!g74) & (g1299) & (!g281) & (!g1300) & (!sk[53]) & (!g1302)) + ((!g74) & (g1299) & (!g281) & (!g1300) & (!sk[53]) & (g1302)) + ((!g74) & (g1299) & (!g281) & (g1300) & (!sk[53]) & (!g1302)) + ((!g74) & (g1299) & (!g281) & (g1300) & (!sk[53]) & (g1302)) + ((!g74) & (g1299) & (g281) & (!g1300) & (!sk[53]) & (!g1302)) + ((!g74) & (g1299) & (g281) & (!g1300) & (!sk[53]) & (g1302)) + ((!g74) & (g1299) & (g281) & (g1300) & (!sk[53]) & (!g1302)) + ((!g74) & (g1299) & (g281) & (g1300) & (!sk[53]) & (g1302)) + ((g74) & (!g1299) & (!g281) & (!g1300) & (sk[53]) & (!g1302)) + ((g74) & (!g1299) & (!g281) & (g1300) & (sk[53]) & (!g1302)) + ((g74) & (!g1299) & (!g281) & (g1300) & (sk[53]) & (g1302)) + ((g74) & (!g1299) & (g281) & (!g1300) & (!sk[53]) & (g1302)) + ((g74) & (!g1299) & (g281) & (!g1300) & (sk[53]) & (!g1302)) + ((g74) & (!g1299) & (g281) & (g1300) & (!sk[53]) & (!g1302)) + ((g74) & (!g1299) & (g281) & (g1300) & (!sk[53]) & (g1302)) + ((g74) & (!g1299) & (g281) & (g1300) & (sk[53]) & (!g1302)) + ((g74) & (!g1299) & (g281) & (g1300) & (sk[53]) & (g1302)) + ((g74) & (g1299) & (!g281) & (!g1300) & (!sk[53]) & (!g1302)) + ((g74) & (g1299) & (!g281) & (!g1300) & (!sk[53]) & (g1302)) + ((g74) & (g1299) & (!g281) & (g1300) & (!sk[53]) & (!g1302)) + ((g74) & (g1299) & (!g281) & (g1300) & (!sk[53]) & (g1302)) + ((g74) & (g1299) & (g281) & (!g1300) & (!sk[53]) & (!g1302)) + ((g74) & (g1299) & (g281) & (!g1300) & (!sk[53]) & (g1302)) + ((g74) & (g1299) & (g281) & (g1300) & (!sk[53]) & (!g1302)) + ((g74) & (g1299) & (g281) & (g1300) & (!sk[53]) & (g1302)));
	assign g1304 = (((!g74) & (!g313) & (!g253) & (g851) & (!g1298) & (g1303)) + ((!g74) & (!g313) & (g253) & (!g851) & (!g1298) & (g1303)) + ((!g74) & (!g313) & (g253) & (g851) & (!g1298) & (g1303)) + ((!g74) & (g313) & (!g253) & (g851) & (!g1298) & (g1303)) + ((!g74) & (g313) & (g253) & (g851) & (!g1298) & (g1303)) + ((g74) & (!g313) & (!g253) & (g851) & (!g1298) & (g1303)) + ((g74) & (!g313) & (g253) & (g851) & (!g1298) & (g1303)) + ((g74) & (g313) & (!g253) & (g851) & (!g1298) & (g1303)) + ((g74) & (g313) & (g253) & (g851) & (!g1298) & (g1303)));
	assign g1305 = (((!g253) & (!sk[55]) & (!g337) & (g339) & (!g849)) + ((!g253) & (!sk[55]) & (!g337) & (g339) & (g849)) + ((!g253) & (!sk[55]) & (g337) & (g339) & (!g849)) + ((!g253) & (!sk[55]) & (g337) & (g339) & (g849)) + ((!g253) & (sk[55]) & (!g337) & (!g339) & (g849)) + ((!g253) & (sk[55]) & (!g337) & (g339) & (!g849)) + ((!g253) & (sk[55]) & (!g337) & (g339) & (g849)) + ((!g253) & (sk[55]) & (g337) & (!g339) & (!g849)) + ((!g253) & (sk[55]) & (g337) & (!g339) & (g849)) + ((!g253) & (sk[55]) & (g337) & (g339) & (!g849)) + ((!g253) & (sk[55]) & (g337) & (g339) & (g849)) + ((g253) & (!sk[55]) & (!g337) & (g339) & (!g849)) + ((g253) & (!sk[55]) & (!g337) & (g339) & (g849)) + ((g253) & (!sk[55]) & (g337) & (g339) & (!g849)) + ((g253) & (!sk[55]) & (g337) & (g339) & (g849)));
	assign g1306 = (((!g37) & (!sk[56]) & (!g102) & (g555) & (!g483)) + ((!g37) & (!sk[56]) & (!g102) & (g555) & (g483)) + ((!g37) & (!sk[56]) & (g102) & (g555) & (!g483)) + ((!g37) & (!sk[56]) & (g102) & (g555) & (g483)) + ((!g37) & (sk[56]) & (g102) & (!g555) & (!g483)) + ((!g37) & (sk[56]) & (g102) & (!g555) & (g483)) + ((!g37) & (sk[56]) & (g102) & (g555) & (!g483)) + ((!g37) & (sk[56]) & (g102) & (g555) & (g483)) + ((g37) & (!sk[56]) & (!g102) & (g555) & (!g483)) + ((g37) & (!sk[56]) & (!g102) & (g555) & (g483)) + ((g37) & (!sk[56]) & (g102) & (g555) & (!g483)) + ((g37) & (!sk[56]) & (g102) & (g555) & (g483)) + ((g37) & (sk[56]) & (g102) & (!g555) & (g483)) + ((g37) & (sk[56]) & (g102) & (g555) & (!g483)) + ((g37) & (sk[56]) & (g102) & (g555) & (g483)));
	assign g1307 = (((!i_12_) & (!i_13_) & (i_14_) & (!g35) & (!sk[57]) & (g102)) + ((!i_12_) & (!i_13_) & (i_14_) & (g35) & (!sk[57]) & (!g102)) + ((!i_12_) & (!i_13_) & (i_14_) & (g35) & (!sk[57]) & (g102)) + ((!i_12_) & (!i_13_) & (i_14_) & (g35) & (sk[57]) & (g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g35) & (!sk[57]) & (!g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g35) & (!sk[57]) & (g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (g35) & (!sk[57]) & (!g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (g35) & (!sk[57]) & (g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (g35) & (sk[57]) & (g102)) + ((!i_12_) & (i_13_) & (i_14_) & (!g35) & (!sk[57]) & (!g102)) + ((!i_12_) & (i_13_) & (i_14_) & (!g35) & (!sk[57]) & (g102)) + ((!i_12_) & (i_13_) & (i_14_) & (g35) & (!sk[57]) & (!g102)) + ((!i_12_) & (i_13_) & (i_14_) & (g35) & (!sk[57]) & (g102)) + ((i_12_) & (!i_13_) & (!i_14_) & (g35) & (sk[57]) & (g102)) + ((i_12_) & (!i_13_) & (i_14_) & (!g35) & (!sk[57]) & (g102)) + ((i_12_) & (!i_13_) & (i_14_) & (g35) & (!sk[57]) & (!g102)) + ((i_12_) & (!i_13_) & (i_14_) & (g35) & (!sk[57]) & (g102)) + ((i_12_) & (i_13_) & (!i_14_) & (!g35) & (!sk[57]) & (!g102)) + ((i_12_) & (i_13_) & (!i_14_) & (!g35) & (!sk[57]) & (g102)) + ((i_12_) & (i_13_) & (!i_14_) & (g35) & (!sk[57]) & (!g102)) + ((i_12_) & (i_13_) & (!i_14_) & (g35) & (!sk[57]) & (g102)) + ((i_12_) & (i_13_) & (!i_14_) & (g35) & (sk[57]) & (g102)) + ((i_12_) & (i_13_) & (i_14_) & (!g35) & (!sk[57]) & (!g102)) + ((i_12_) & (i_13_) & (i_14_) & (!g35) & (!sk[57]) & (g102)) + ((i_12_) & (i_13_) & (i_14_) & (g35) & (!sk[57]) & (!g102)) + ((i_12_) & (i_13_) & (i_14_) & (g35) & (!sk[57]) & (g102)) + ((i_12_) & (i_13_) & (i_14_) & (g35) & (sk[57]) & (g102)));
	assign g1308 = (((!g634) & (!g135) & (!sk[58]) & (g131) & (!g281) & (g513)) + ((!g634) & (!g135) & (!sk[58]) & (g131) & (g281) & (!g513)) + ((!g634) & (!g135) & (!sk[58]) & (g131) & (g281) & (g513)) + ((!g634) & (g135) & (!sk[58]) & (!g131) & (!g281) & (!g513)) + ((!g634) & (g135) & (!sk[58]) & (!g131) & (!g281) & (g513)) + ((!g634) & (g135) & (!sk[58]) & (!g131) & (g281) & (!g513)) + ((!g634) & (g135) & (!sk[58]) & (!g131) & (g281) & (g513)) + ((!g634) & (g135) & (!sk[58]) & (g131) & (!g281) & (!g513)) + ((!g634) & (g135) & (!sk[58]) & (g131) & (!g281) & (g513)) + ((!g634) & (g135) & (!sk[58]) & (g131) & (g281) & (!g513)) + ((!g634) & (g135) & (!sk[58]) & (g131) & (g281) & (g513)) + ((!g634) & (g135) & (sk[58]) & (g131) & (!g281) & (!g513)) + ((!g634) & (g135) & (sk[58]) & (g131) & (!g281) & (g513)) + ((!g634) & (g135) & (sk[58]) & (g131) & (g281) & (!g513)) + ((!g634) & (g135) & (sk[58]) & (g131) & (g281) & (g513)) + ((g634) & (!g135) & (!sk[58]) & (g131) & (!g281) & (g513)) + ((g634) & (!g135) & (!sk[58]) & (g131) & (g281) & (!g513)) + ((g634) & (!g135) & (!sk[58]) & (g131) & (g281) & (g513)) + ((g634) & (!g135) & (sk[58]) & (!g131) & (!g281) & (g513)) + ((g634) & (!g135) & (sk[58]) & (g131) & (!g281) & (g513)) + ((g634) & (g135) & (!sk[58]) & (!g131) & (!g281) & (!g513)) + ((g634) & (g135) & (!sk[58]) & (!g131) & (!g281) & (g513)) + ((g634) & (g135) & (!sk[58]) & (!g131) & (g281) & (!g513)) + ((g634) & (g135) & (!sk[58]) & (!g131) & (g281) & (g513)) + ((g634) & (g135) & (!sk[58]) & (g131) & (!g281) & (!g513)) + ((g634) & (g135) & (!sk[58]) & (g131) & (!g281) & (g513)) + ((g634) & (g135) & (!sk[58]) & (g131) & (g281) & (!g513)) + ((g634) & (g135) & (!sk[58]) & (g131) & (g281) & (g513)) + ((g634) & (g135) & (sk[58]) & (!g131) & (!g281) & (g513)) + ((g634) & (g135) & (sk[58]) & (g131) & (!g281) & (!g513)) + ((g634) & (g135) & (sk[58]) & (g131) & (!g281) & (g513)) + ((g634) & (g135) & (sk[58]) & (g131) & (g281) & (!g513)) + ((g634) & (g135) & (sk[58]) & (g131) & (g281) & (g513)));
	assign g1309 = (((!sk[59]) & (!g1305) & (!g1306) & (g1307) & (!g1308)) + ((!sk[59]) & (!g1305) & (!g1306) & (g1307) & (g1308)) + ((!sk[59]) & (!g1305) & (g1306) & (g1307) & (!g1308)) + ((!sk[59]) & (!g1305) & (g1306) & (g1307) & (g1308)) + ((!sk[59]) & (g1305) & (!g1306) & (g1307) & (!g1308)) + ((!sk[59]) & (g1305) & (!g1306) & (g1307) & (g1308)) + ((!sk[59]) & (g1305) & (g1306) & (g1307) & (!g1308)) + ((!sk[59]) & (g1305) & (g1306) & (g1307) & (g1308)) + ((sk[59]) & (!g1305) & (!g1306) & (!g1307) & (g1308)));
	assign g1310 = (((!i_12_) & (!i_13_) & (!i_14_) & (g35) & (!g36) & (!g159)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g35) & (g36) & (!g159)) + ((!i_12_) & (!i_13_) & (i_14_) & (!g35) & (g36) & (!g159)) + ((!i_12_) & (!i_13_) & (i_14_) & (g35) & (!g36) & (!g159)) + ((!i_12_) & (!i_13_) & (i_14_) & (g35) & (g36) & (!g159)) + ((!i_12_) & (i_13_) & (!i_14_) & (!g35) & (g36) & (!g159)) + ((!i_12_) & (i_13_) & (!i_14_) & (g35) & (g36) & (!g159)) + ((!i_12_) & (i_13_) & (i_14_) & (!g35) & (g36) & (!g159)) + ((!i_12_) & (i_13_) & (i_14_) & (g35) & (!g36) & (!g159)) + ((!i_12_) & (i_13_) & (i_14_) & (g35) & (g36) & (!g159)) + ((i_12_) & (!i_13_) & (i_14_) & (!g35) & (g36) & (!g159)) + ((i_12_) & (!i_13_) & (i_14_) & (g35) & (!g36) & (!g159)) + ((i_12_) & (!i_13_) & (i_14_) & (g35) & (g36) & (!g159)) + ((i_12_) & (i_13_) & (i_14_) & (!g35) & (g36) & (!g159)) + ((i_12_) & (i_13_) & (i_14_) & (g35) & (!g36) & (!g159)) + ((i_12_) & (i_13_) & (i_14_) & (g35) & (g36) & (!g159)));
	assign g1311 = (((!g90) & (!g74) & (!g281) & (!g513) & (!g635) & (!g1310)) + ((!g90) & (!g74) & (!g281) & (!g513) & (g635) & (!g1310)) + ((!g90) & (!g74) & (!g281) & (g513) & (!g635) & (!g1310)) + ((!g90) & (!g74) & (!g281) & (g513) & (g635) & (!g1310)) + ((!g90) & (!g74) & (g281) & (!g513) & (!g635) & (!g1310)) + ((!g90) & (!g74) & (g281) & (!g513) & (g635) & (!g1310)) + ((!g90) & (!g74) & (g281) & (g513) & (!g635) & (!g1310)) + ((!g90) & (!g74) & (g281) & (g513) & (g635) & (!g1310)) + ((!g90) & (g74) & (!g281) & (g513) & (!g635) & (!g1310)) + ((g90) & (!g74) & (!g281) & (!g513) & (!g635) & (!g1310)) + ((g90) & (!g74) & (!g281) & (!g513) & (g635) & (!g1310)) + ((g90) & (!g74) & (!g281) & (g513) & (!g635) & (!g1310)) + ((g90) & (!g74) & (!g281) & (g513) & (g635) & (!g1310)) + ((g90) & (!g74) & (g281) & (!g513) & (!g635) & (!g1310)) + ((g90) & (!g74) & (g281) & (!g513) & (g635) & (!g1310)) + ((g90) & (!g74) & (g281) & (g513) & (!g635) & (!g1310)) + ((g90) & (!g74) & (g281) & (g513) & (g635) & (!g1310)));
	assign g1312 = (((!sk[62]) & (!g673) & (!g926) & (g1045) & (!g1309) & (g1311)) + ((!sk[62]) & (!g673) & (!g926) & (g1045) & (g1309) & (!g1311)) + ((!sk[62]) & (!g673) & (!g926) & (g1045) & (g1309) & (g1311)) + ((!sk[62]) & (!g673) & (g926) & (!g1045) & (!g1309) & (!g1311)) + ((!sk[62]) & (!g673) & (g926) & (!g1045) & (!g1309) & (g1311)) + ((!sk[62]) & (!g673) & (g926) & (!g1045) & (g1309) & (!g1311)) + ((!sk[62]) & (!g673) & (g926) & (!g1045) & (g1309) & (g1311)) + ((!sk[62]) & (!g673) & (g926) & (g1045) & (!g1309) & (!g1311)) + ((!sk[62]) & (!g673) & (g926) & (g1045) & (!g1309) & (g1311)) + ((!sk[62]) & (!g673) & (g926) & (g1045) & (g1309) & (!g1311)) + ((!sk[62]) & (!g673) & (g926) & (g1045) & (g1309) & (g1311)) + ((!sk[62]) & (g673) & (!g926) & (g1045) & (!g1309) & (g1311)) + ((!sk[62]) & (g673) & (!g926) & (g1045) & (g1309) & (!g1311)) + ((!sk[62]) & (g673) & (!g926) & (g1045) & (g1309) & (g1311)) + ((!sk[62]) & (g673) & (g926) & (!g1045) & (!g1309) & (!g1311)) + ((!sk[62]) & (g673) & (g926) & (!g1045) & (!g1309) & (g1311)) + ((!sk[62]) & (g673) & (g926) & (!g1045) & (g1309) & (!g1311)) + ((!sk[62]) & (g673) & (g926) & (!g1045) & (g1309) & (g1311)) + ((!sk[62]) & (g673) & (g926) & (g1045) & (!g1309) & (!g1311)) + ((!sk[62]) & (g673) & (g926) & (g1045) & (!g1309) & (g1311)) + ((!sk[62]) & (g673) & (g926) & (g1045) & (g1309) & (!g1311)) + ((!sk[62]) & (g673) & (g926) & (g1045) & (g1309) & (g1311)) + ((sk[62]) & (!g673) & (g926) & (g1045) & (g1309) & (g1311)));
	assign g1313 = (((!i_12_) & (!i_13_) & (!i_14_) & (!g35) & (g36) & (g74)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g35) & (g36) & (g74)) + ((!i_12_) & (!i_13_) & (i_14_) & (g35) & (!g36) & (g74)) + ((!i_12_) & (!i_13_) & (i_14_) & (g35) & (g36) & (g74)) + ((!i_12_) & (i_13_) & (!i_14_) & (g35) & (!g36) & (g74)) + ((!i_12_) & (i_13_) & (!i_14_) & (g35) & (g36) & (g74)) + ((!i_12_) & (i_13_) & (i_14_) & (g35) & (!g36) & (g74)) + ((!i_12_) & (i_13_) & (i_14_) & (g35) & (g36) & (g74)) + ((i_12_) & (!i_13_) & (i_14_) & (!g35) & (g36) & (g74)) + ((i_12_) & (!i_13_) & (i_14_) & (g35) & (g36) & (g74)) + ((i_12_) & (i_13_) & (!i_14_) & (!g35) & (g36) & (g74)) + ((i_12_) & (i_13_) & (!i_14_) & (g35) & (g36) & (g74)) + ((i_12_) & (i_13_) & (i_14_) & (g35) & (!g36) & (g74)) + ((i_12_) & (i_13_) & (i_14_) & (g35) & (g36) & (g74)));
	assign g1314 = (((!g35) & (!g339) & (!g460) & (sk[64]) & (!g641)) + ((!g35) & (!g339) & (g460) & (!sk[64]) & (!g641)) + ((!g35) & (!g339) & (g460) & (!sk[64]) & (g641)) + ((!g35) & (!g339) & (g460) & (sk[64]) & (!g641)) + ((!g35) & (g339) & (g460) & (!sk[64]) & (!g641)) + ((!g35) & (g339) & (g460) & (!sk[64]) & (g641)) + ((g35) & (!g339) & (g460) & (!sk[64]) & (!g641)) + ((g35) & (!g339) & (g460) & (!sk[64]) & (g641)) + ((g35) & (!g339) & (g460) & (sk[64]) & (!g641)) + ((g35) & (g339) & (g460) & (!sk[64]) & (!g641)) + ((g35) & (g339) & (g460) & (!sk[64]) & (g641)));
	assign g1315 = (((!sk[65]) & (!i_8_) & (!i_7_) & (g924) & (!g394)) + ((!sk[65]) & (!i_8_) & (!i_7_) & (g924) & (g394)) + ((!sk[65]) & (!i_8_) & (i_7_) & (g924) & (!g394)) + ((!sk[65]) & (!i_8_) & (i_7_) & (g924) & (g394)) + ((!sk[65]) & (i_8_) & (!i_7_) & (g924) & (!g394)) + ((!sk[65]) & (i_8_) & (!i_7_) & (g924) & (g394)) + ((!sk[65]) & (i_8_) & (i_7_) & (g924) & (!g394)) + ((!sk[65]) & (i_8_) & (i_7_) & (g924) & (g394)) + ((sk[65]) & (!i_8_) & (i_7_) & (g924) & (g394)));
	assign g1316 = (((!g135) & (!g1314) & (!sk[66]) & (g1315) & (!g204)) + ((!g135) & (!g1314) & (!sk[66]) & (g1315) & (g204)) + ((!g135) & (g1314) & (!sk[66]) & (g1315) & (!g204)) + ((!g135) & (g1314) & (!sk[66]) & (g1315) & (g204)) + ((!g135) & (g1314) & (sk[66]) & (!g1315) & (g204)) + ((g135) & (!g1314) & (!sk[66]) & (g1315) & (!g204)) + ((g135) & (!g1314) & (!sk[66]) & (g1315) & (g204)) + ((g135) & (!g1314) & (sk[66]) & (!g1315) & (g204)) + ((g135) & (g1314) & (!sk[66]) & (g1315) & (!g204)) + ((g135) & (g1314) & (!sk[66]) & (g1315) & (g204)) + ((g135) & (g1314) & (sk[66]) & (!g1315) & (g204)));
	assign g1317 = (((!g313) & (!g348) & (!g514) & (sk[67]) & (g746)) + ((!g313) & (!g348) & (g514) & (!sk[67]) & (!g746)) + ((!g313) & (!g348) & (g514) & (!sk[67]) & (g746)) + ((!g313) & (g348) & (!g514) & (sk[67]) & (g746)) + ((!g313) & (g348) & (g514) & (!sk[67]) & (!g746)) + ((!g313) & (g348) & (g514) & (!sk[67]) & (g746)) + ((!g313) & (g348) & (g514) & (sk[67]) & (g746)) + ((g313) & (!g348) & (!g514) & (sk[67]) & (g746)) + ((g313) & (!g348) & (g514) & (!sk[67]) & (!g746)) + ((g313) & (!g348) & (g514) & (!sk[67]) & (g746)) + ((g313) & (g348) & (!g514) & (sk[67]) & (g746)) + ((g313) & (g348) & (g514) & (!sk[67]) & (!g746)) + ((g313) & (g348) & (g514) & (!sk[67]) & (g746)));
	assign g1318 = (((!g257) & (!g605) & (!sk[68]) & (g1313) & (!g1316) & (g1317)) + ((!g257) & (!g605) & (!sk[68]) & (g1313) & (g1316) & (!g1317)) + ((!g257) & (!g605) & (!sk[68]) & (g1313) & (g1316) & (g1317)) + ((!g257) & (!g605) & (sk[68]) & (!g1313) & (g1316) & (g1317)) + ((!g257) & (g605) & (!sk[68]) & (!g1313) & (!g1316) & (!g1317)) + ((!g257) & (g605) & (!sk[68]) & (!g1313) & (!g1316) & (g1317)) + ((!g257) & (g605) & (!sk[68]) & (!g1313) & (g1316) & (!g1317)) + ((!g257) & (g605) & (!sk[68]) & (!g1313) & (g1316) & (g1317)) + ((!g257) & (g605) & (!sk[68]) & (g1313) & (!g1316) & (!g1317)) + ((!g257) & (g605) & (!sk[68]) & (g1313) & (!g1316) & (g1317)) + ((!g257) & (g605) & (!sk[68]) & (g1313) & (g1316) & (!g1317)) + ((!g257) & (g605) & (!sk[68]) & (g1313) & (g1316) & (g1317)) + ((!g257) & (g605) & (sk[68]) & (!g1313) & (g1316) & (g1317)) + ((g257) & (!g605) & (!sk[68]) & (g1313) & (!g1316) & (g1317)) + ((g257) & (!g605) & (!sk[68]) & (g1313) & (g1316) & (!g1317)) + ((g257) & (!g605) & (!sk[68]) & (g1313) & (g1316) & (g1317)) + ((g257) & (!g605) & (sk[68]) & (!g1313) & (g1316) & (g1317)) + ((g257) & (g605) & (!sk[68]) & (!g1313) & (!g1316) & (!g1317)) + ((g257) & (g605) & (!sk[68]) & (!g1313) & (!g1316) & (g1317)) + ((g257) & (g605) & (!sk[68]) & (!g1313) & (g1316) & (!g1317)) + ((g257) & (g605) & (!sk[68]) & (!g1313) & (g1316) & (g1317)) + ((g257) & (g605) & (!sk[68]) & (g1313) & (!g1316) & (!g1317)) + ((g257) & (g605) & (!sk[68]) & (g1313) & (!g1316) & (g1317)) + ((g257) & (g605) & (!sk[68]) & (g1313) & (g1316) & (!g1317)) + ((g257) & (g605) & (!sk[68]) & (g1313) & (g1316) & (g1317)));
	assign g1319 = (((g1010) & (g506) & (g1297) & (g1304) & (g1312) & (g1318)));
	assign g1320 = (((!i_14_) & (!g27) & (!sk[70]) & (g102)) + ((!i_14_) & (g27) & (!sk[70]) & (!g102)) + ((!i_14_) & (g27) & (!sk[70]) & (g102)) + ((i_14_) & (!g27) & (!sk[70]) & (g102)) + ((i_14_) & (g27) & (!sk[70]) & (!g102)) + ((i_14_) & (g27) & (!sk[70]) & (g102)) + ((i_14_) & (g27) & (sk[70]) & (g102)));
	assign g1321 = (((!sk[71]) & (!g17) & (!g76) & (g135) & (!g460)) + ((!sk[71]) & (!g17) & (!g76) & (g135) & (g460)) + ((!sk[71]) & (!g17) & (g76) & (g135) & (!g460)) + ((!sk[71]) & (!g17) & (g76) & (g135) & (g460)) + ((!sk[71]) & (g17) & (!g76) & (g135) & (!g460)) + ((!sk[71]) & (g17) & (!g76) & (g135) & (g460)) + ((!sk[71]) & (g17) & (g76) & (g135) & (!g460)) + ((!sk[71]) & (g17) & (g76) & (g135) & (g460)) + ((sk[71]) & (g17) & (!g76) & (!g135) & (!g460)) + ((sk[71]) & (g17) & (!g76) & (!g135) & (g460)) + ((sk[71]) & (g17) & (g76) & (!g135) & (!g460)));
	assign g1322 = (((!g159) & (!sk[72]) & (!g253) & (g334) & (!g875)) + ((!g159) & (!sk[72]) & (!g253) & (g334) & (g875)) + ((!g159) & (!sk[72]) & (g253) & (g334) & (!g875)) + ((!g159) & (!sk[72]) & (g253) & (g334) & (g875)) + ((!g159) & (sk[72]) & (!g253) & (g334) & (!g875)) + ((!g159) & (sk[72]) & (g253) & (g334) & (!g875)) + ((g159) & (!sk[72]) & (!g253) & (g334) & (!g875)) + ((g159) & (!sk[72]) & (!g253) & (g334) & (g875)) + ((g159) & (!sk[72]) & (g253) & (g334) & (!g875)) + ((g159) & (!sk[72]) & (g253) & (g334) & (g875)) + ((g159) & (sk[72]) & (!g253) & (g334) & (!g875)) + ((g159) & (sk[72]) & (!g253) & (g334) & (g875)) + ((g159) & (sk[72]) & (g253) & (!g334) & (!g875)) + ((g159) & (sk[72]) & (g253) & (!g334) & (g875)) + ((g159) & (sk[72]) & (g253) & (g334) & (!g875)) + ((g159) & (sk[72]) & (g253) & (g334) & (g875)));
	assign g1323 = (((!sk[73]) & (!g135) & (!g185) & (g180) & (!g1321) & (g1322)) + ((!sk[73]) & (!g135) & (!g185) & (g180) & (g1321) & (!g1322)) + ((!sk[73]) & (!g135) & (!g185) & (g180) & (g1321) & (g1322)) + ((!sk[73]) & (!g135) & (g185) & (!g180) & (!g1321) & (!g1322)) + ((!sk[73]) & (!g135) & (g185) & (!g180) & (!g1321) & (g1322)) + ((!sk[73]) & (!g135) & (g185) & (!g180) & (g1321) & (!g1322)) + ((!sk[73]) & (!g135) & (g185) & (!g180) & (g1321) & (g1322)) + ((!sk[73]) & (!g135) & (g185) & (g180) & (!g1321) & (!g1322)) + ((!sk[73]) & (!g135) & (g185) & (g180) & (!g1321) & (g1322)) + ((!sk[73]) & (!g135) & (g185) & (g180) & (g1321) & (!g1322)) + ((!sk[73]) & (!g135) & (g185) & (g180) & (g1321) & (g1322)) + ((!sk[73]) & (g135) & (!g185) & (g180) & (!g1321) & (g1322)) + ((!sk[73]) & (g135) & (!g185) & (g180) & (g1321) & (!g1322)) + ((!sk[73]) & (g135) & (!g185) & (g180) & (g1321) & (g1322)) + ((!sk[73]) & (g135) & (g185) & (!g180) & (!g1321) & (!g1322)) + ((!sk[73]) & (g135) & (g185) & (!g180) & (!g1321) & (g1322)) + ((!sk[73]) & (g135) & (g185) & (!g180) & (g1321) & (!g1322)) + ((!sk[73]) & (g135) & (g185) & (!g180) & (g1321) & (g1322)) + ((!sk[73]) & (g135) & (g185) & (g180) & (!g1321) & (!g1322)) + ((!sk[73]) & (g135) & (g185) & (g180) & (!g1321) & (g1322)) + ((!sk[73]) & (g135) & (g185) & (g180) & (g1321) & (!g1322)) + ((!sk[73]) & (g135) & (g185) & (g180) & (g1321) & (g1322)) + ((sk[73]) & (!g135) & (!g185) & (!g180) & (!g1321) & (g1322)) + ((sk[73]) & (g135) & (!g185) & (!g180) & (!g1321) & (g1322)) + ((sk[73]) & (g135) & (!g185) & (g180) & (!g1321) & (g1322)) + ((sk[73]) & (g135) & (g185) & (!g180) & (!g1321) & (g1322)) + ((sk[73]) & (g135) & (g185) & (g180) & (!g1321) & (g1322)));
	assign g1324 = (((!sk[74]) & (!g74) & (!g180) & (g461) & (!g1320) & (g1323)) + ((!sk[74]) & (!g74) & (!g180) & (g461) & (g1320) & (!g1323)) + ((!sk[74]) & (!g74) & (!g180) & (g461) & (g1320) & (g1323)) + ((!sk[74]) & (!g74) & (g180) & (!g461) & (!g1320) & (!g1323)) + ((!sk[74]) & (!g74) & (g180) & (!g461) & (!g1320) & (g1323)) + ((!sk[74]) & (!g74) & (g180) & (!g461) & (g1320) & (!g1323)) + ((!sk[74]) & (!g74) & (g180) & (!g461) & (g1320) & (g1323)) + ((!sk[74]) & (!g74) & (g180) & (g461) & (!g1320) & (!g1323)) + ((!sk[74]) & (!g74) & (g180) & (g461) & (!g1320) & (g1323)) + ((!sk[74]) & (!g74) & (g180) & (g461) & (g1320) & (!g1323)) + ((!sk[74]) & (!g74) & (g180) & (g461) & (g1320) & (g1323)) + ((!sk[74]) & (g74) & (!g180) & (g461) & (!g1320) & (g1323)) + ((!sk[74]) & (g74) & (!g180) & (g461) & (g1320) & (!g1323)) + ((!sk[74]) & (g74) & (!g180) & (g461) & (g1320) & (g1323)) + ((!sk[74]) & (g74) & (g180) & (!g461) & (!g1320) & (!g1323)) + ((!sk[74]) & (g74) & (g180) & (!g461) & (!g1320) & (g1323)) + ((!sk[74]) & (g74) & (g180) & (!g461) & (g1320) & (!g1323)) + ((!sk[74]) & (g74) & (g180) & (!g461) & (g1320) & (g1323)) + ((!sk[74]) & (g74) & (g180) & (g461) & (!g1320) & (!g1323)) + ((!sk[74]) & (g74) & (g180) & (g461) & (!g1320) & (g1323)) + ((!sk[74]) & (g74) & (g180) & (g461) & (g1320) & (!g1323)) + ((!sk[74]) & (g74) & (g180) & (g461) & (g1320) & (g1323)) + ((sk[74]) & (!g74) & (!g180) & (!g461) & (!g1320) & (g1323)) + ((sk[74]) & (!g74) & (!g180) & (g461) & (!g1320) & (g1323)) + ((sk[74]) & (!g74) & (g180) & (!g461) & (!g1320) & (g1323)) + ((sk[74]) & (!g74) & (g180) & (g461) & (!g1320) & (g1323)) + ((sk[74]) & (g74) & (!g180) & (!g461) & (!g1320) & (g1323)));
	assign g1325 = (((!sk[75]) & (!g28) & (!g135) & (g275)) + ((!sk[75]) & (!g28) & (g135) & (!g275)) + ((!sk[75]) & (!g28) & (g135) & (g275)) + ((!sk[75]) & (g28) & (!g135) & (g275)) + ((!sk[75]) & (g28) & (g135) & (!g275)) + ((!sk[75]) & (g28) & (g135) & (g275)) + ((sk[75]) & (!g28) & (!g135) & (g275)) + ((sk[75]) & (g28) & (!g135) & (!g275)) + ((sk[75]) & (g28) & (!g135) & (g275)));
	assign g1326 = (((!sk[76]) & (!i_12_) & (!i_13_) & (i_14_) & (!g17) & (g102)) + ((!sk[76]) & (!i_12_) & (!i_13_) & (i_14_) & (g17) & (!g102)) + ((!sk[76]) & (!i_12_) & (!i_13_) & (i_14_) & (g17) & (g102)) + ((!sk[76]) & (!i_12_) & (i_13_) & (!i_14_) & (!g17) & (!g102)) + ((!sk[76]) & (!i_12_) & (i_13_) & (!i_14_) & (!g17) & (g102)) + ((!sk[76]) & (!i_12_) & (i_13_) & (!i_14_) & (g17) & (!g102)) + ((!sk[76]) & (!i_12_) & (i_13_) & (!i_14_) & (g17) & (g102)) + ((!sk[76]) & (!i_12_) & (i_13_) & (i_14_) & (!g17) & (!g102)) + ((!sk[76]) & (!i_12_) & (i_13_) & (i_14_) & (!g17) & (g102)) + ((!sk[76]) & (!i_12_) & (i_13_) & (i_14_) & (g17) & (!g102)) + ((!sk[76]) & (!i_12_) & (i_13_) & (i_14_) & (g17) & (g102)) + ((!sk[76]) & (i_12_) & (!i_13_) & (i_14_) & (!g17) & (g102)) + ((!sk[76]) & (i_12_) & (!i_13_) & (i_14_) & (g17) & (!g102)) + ((!sk[76]) & (i_12_) & (!i_13_) & (i_14_) & (g17) & (g102)) + ((!sk[76]) & (i_12_) & (i_13_) & (!i_14_) & (!g17) & (!g102)) + ((!sk[76]) & (i_12_) & (i_13_) & (!i_14_) & (!g17) & (g102)) + ((!sk[76]) & (i_12_) & (i_13_) & (!i_14_) & (g17) & (!g102)) + ((!sk[76]) & (i_12_) & (i_13_) & (!i_14_) & (g17) & (g102)) + ((!sk[76]) & (i_12_) & (i_13_) & (i_14_) & (!g17) & (!g102)) + ((!sk[76]) & (i_12_) & (i_13_) & (i_14_) & (!g17) & (g102)) + ((!sk[76]) & (i_12_) & (i_13_) & (i_14_) & (g17) & (!g102)) + ((!sk[76]) & (i_12_) & (i_13_) & (i_14_) & (g17) & (g102)) + ((sk[76]) & (!i_12_) & (!i_13_) & (i_14_) & (g17) & (g102)) + ((sk[76]) & (!i_12_) & (i_13_) & (!i_14_) & (g17) & (g102)) + ((sk[76]) & (!i_12_) & (i_13_) & (i_14_) & (g17) & (g102)) + ((sk[76]) & (i_12_) & (!i_13_) & (i_14_) & (g17) & (g102)) + ((sk[76]) & (i_12_) & (i_13_) & (i_14_) & (g17) & (g102)));
	assign g1327 = (((!i_8_) & (!g73) & (!sk[77]) & (g578) & (!g993)) + ((!i_8_) & (!g73) & (!sk[77]) & (g578) & (g993)) + ((!i_8_) & (g73) & (!sk[77]) & (g578) & (!g993)) + ((!i_8_) & (g73) & (!sk[77]) & (g578) & (g993)) + ((!i_8_) & (g73) & (sk[77]) & (!g578) & (g993)) + ((!i_8_) & (g73) & (sk[77]) & (g578) & (!g993)) + ((!i_8_) & (g73) & (sk[77]) & (g578) & (g993)) + ((i_8_) & (!g73) & (!sk[77]) & (g578) & (!g993)) + ((i_8_) & (!g73) & (!sk[77]) & (g578) & (g993)) + ((i_8_) & (g73) & (!sk[77]) & (g578) & (!g993)) + ((i_8_) & (g73) & (!sk[77]) & (g578) & (g993)));
	assign g1328 = (((!i_12_) & (!i_13_) & (!i_14_) & (g17) & (!g159) & (!g131)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g17) & (!g159) & (g131)) + ((!i_12_) & (!i_13_) & (!i_14_) & (g17) & (g159) & (!g131)) + ((!i_12_) & (!i_13_) & (i_14_) & (g17) & (!g159) & (!g131)) + ((!i_12_) & (!i_13_) & (i_14_) & (g17) & (!g159) & (g131)) + ((!i_12_) & (i_13_) & (i_14_) & (g17) & (!g159) & (!g131)) + ((!i_12_) & (i_13_) & (i_14_) & (g17) & (!g159) & (g131)) + ((!i_12_) & (i_13_) & (i_14_) & (g17) & (g159) & (!g131)) + ((i_12_) & (!i_13_) & (!i_14_) & (g17) & (!g159) & (!g131)) + ((i_12_) & (!i_13_) & (!i_14_) & (g17) & (!g159) & (g131)) + ((i_12_) & (!i_13_) & (!i_14_) & (g17) & (g159) & (!g131)) + ((i_12_) & (!i_13_) & (i_14_) & (g17) & (!g159) & (!g131)) + ((i_12_) & (!i_13_) & (i_14_) & (g17) & (!g159) & (g131)) + ((i_12_) & (!i_13_) & (i_14_) & (g17) & (g159) & (!g131)) + ((i_12_) & (i_13_) & (!i_14_) & (g17) & (!g159) & (!g131)) + ((i_12_) & (i_13_) & (!i_14_) & (g17) & (!g159) & (g131)) + ((i_12_) & (i_13_) & (!i_14_) & (g17) & (g159) & (!g131)));
	assign g1329 = (((!g1325) & (!g277) & (!sk[79]) & (g1326) & (!g1327) & (g1328)) + ((!g1325) & (!g277) & (!sk[79]) & (g1326) & (g1327) & (!g1328)) + ((!g1325) & (!g277) & (!sk[79]) & (g1326) & (g1327) & (g1328)) + ((!g1325) & (!g277) & (sk[79]) & (!g1326) & (!g1327) & (!g1328)) + ((!g1325) & (g277) & (!sk[79]) & (!g1326) & (!g1327) & (!g1328)) + ((!g1325) & (g277) & (!sk[79]) & (!g1326) & (!g1327) & (g1328)) + ((!g1325) & (g277) & (!sk[79]) & (!g1326) & (g1327) & (!g1328)) + ((!g1325) & (g277) & (!sk[79]) & (!g1326) & (g1327) & (g1328)) + ((!g1325) & (g277) & (!sk[79]) & (g1326) & (!g1327) & (!g1328)) + ((!g1325) & (g277) & (!sk[79]) & (g1326) & (!g1327) & (g1328)) + ((!g1325) & (g277) & (!sk[79]) & (g1326) & (g1327) & (!g1328)) + ((!g1325) & (g277) & (!sk[79]) & (g1326) & (g1327) & (g1328)) + ((g1325) & (!g277) & (!sk[79]) & (g1326) & (!g1327) & (g1328)) + ((g1325) & (!g277) & (!sk[79]) & (g1326) & (g1327) & (!g1328)) + ((g1325) & (!g277) & (!sk[79]) & (g1326) & (g1327) & (g1328)) + ((g1325) & (g277) & (!sk[79]) & (!g1326) & (!g1327) & (!g1328)) + ((g1325) & (g277) & (!sk[79]) & (!g1326) & (!g1327) & (g1328)) + ((g1325) & (g277) & (!sk[79]) & (!g1326) & (g1327) & (!g1328)) + ((g1325) & (g277) & (!sk[79]) & (!g1326) & (g1327) & (g1328)) + ((g1325) & (g277) & (!sk[79]) & (g1326) & (!g1327) & (!g1328)) + ((g1325) & (g277) & (!sk[79]) & (g1326) & (!g1327) & (g1328)) + ((g1325) & (g277) & (!sk[79]) & (g1326) & (g1327) & (!g1328)) + ((g1325) & (g277) & (!sk[79]) & (g1326) & (g1327) & (g1328)));
	assign g1330 = (((!g74) & (!g402) & (!g337) & (!g605) & (!g993) & (g1107)) + ((!g74) & (!g402) & (!g337) & (g605) & (!g993) & (g1107)) + ((!g74) & (!g402) & (g337) & (!g605) & (!g993) & (g1107)) + ((!g74) & (!g402) & (g337) & (g605) & (!g993) & (g1107)) + ((!g74) & (g402) & (!g337) & (!g605) & (!g993) & (!g1107)) + ((!g74) & (g402) & (!g337) & (!g605) & (!g993) & (g1107)) + ((!g74) & (g402) & (!g337) & (!g605) & (g993) & (!g1107)) + ((!g74) & (g402) & (!g337) & (!g605) & (g993) & (g1107)) + ((!g74) & (g402) & (!g337) & (g605) & (!g993) & (!g1107)) + ((!g74) & (g402) & (!g337) & (g605) & (!g993) & (g1107)) + ((!g74) & (g402) & (!g337) & (g605) & (g993) & (!g1107)) + ((!g74) & (g402) & (!g337) & (g605) & (g993) & (g1107)) + ((!g74) & (g402) & (g337) & (!g605) & (!g993) & (!g1107)) + ((!g74) & (g402) & (g337) & (!g605) & (!g993) & (g1107)) + ((!g74) & (g402) & (g337) & (!g605) & (g993) & (!g1107)) + ((!g74) & (g402) & (g337) & (!g605) & (g993) & (g1107)) + ((!g74) & (g402) & (g337) & (g605) & (!g993) & (!g1107)) + ((!g74) & (g402) & (g337) & (g605) & (!g993) & (g1107)) + ((!g74) & (g402) & (g337) & (g605) & (g993) & (!g1107)) + ((!g74) & (g402) & (g337) & (g605) & (g993) & (g1107)) + ((g74) & (!g402) & (!g337) & (!g605) & (!g993) & (g1107)) + ((g74) & (g402) & (!g337) & (!g605) & (!g993) & (g1107)) + ((g74) & (g402) & (!g337) & (!g605) & (g993) & (g1107)));
	assign g1331 = (((!g130) & (!g131) & (!sk[81]) & (g334) & (!g875)) + ((!g130) & (!g131) & (!sk[81]) & (g334) & (g875)) + ((!g130) & (!g131) & (sk[81]) & (g334) & (!g875)) + ((!g130) & (g131) & (!sk[81]) & (g334) & (!g875)) + ((!g130) & (g131) & (!sk[81]) & (g334) & (g875)) + ((!g130) & (g131) & (sk[81]) & (g334) & (!g875)) + ((g130) & (!g131) & (!sk[81]) & (g334) & (!g875)) + ((g130) & (!g131) & (!sk[81]) & (g334) & (g875)) + ((g130) & (!g131) & (sk[81]) & (g334) & (!g875)) + ((g130) & (g131) & (!sk[81]) & (g334) & (!g875)) + ((g130) & (g131) & (!sk[81]) & (g334) & (g875)) + ((g130) & (g131) & (sk[81]) & (!g334) & (!g875)) + ((g130) & (g131) & (sk[81]) & (!g334) & (g875)) + ((g130) & (g131) & (sk[81]) & (g334) & (!g875)) + ((g130) & (g131) & (sk[81]) & (g334) & (g875)));
	assign g1332 = (((!g18) & (!g33) & (!g74) & (sk[82]) & (g1331) & (!g937)) + ((!g18) & (!g33) & (g74) & (!sk[82]) & (!g1331) & (g937)) + ((!g18) & (!g33) & (g74) & (!sk[82]) & (g1331) & (!g937)) + ((!g18) & (!g33) & (g74) & (!sk[82]) & (g1331) & (g937)) + ((!g18) & (!g33) & (g74) & (sk[82]) & (g1331) & (!g937)) + ((!g18) & (g33) & (!g74) & (!sk[82]) & (!g1331) & (!g937)) + ((!g18) & (g33) & (!g74) & (!sk[82]) & (!g1331) & (g937)) + ((!g18) & (g33) & (!g74) & (!sk[82]) & (g1331) & (!g937)) + ((!g18) & (g33) & (!g74) & (!sk[82]) & (g1331) & (g937)) + ((!g18) & (g33) & (!g74) & (sk[82]) & (g1331) & (!g937)) + ((!g18) & (g33) & (g74) & (!sk[82]) & (!g1331) & (!g937)) + ((!g18) & (g33) & (g74) & (!sk[82]) & (!g1331) & (g937)) + ((!g18) & (g33) & (g74) & (!sk[82]) & (g1331) & (!g937)) + ((!g18) & (g33) & (g74) & (!sk[82]) & (g1331) & (g937)) + ((g18) & (!g33) & (!g74) & (sk[82]) & (g1331) & (!g937)) + ((g18) & (!g33) & (g74) & (!sk[82]) & (!g1331) & (g937)) + ((g18) & (!g33) & (g74) & (!sk[82]) & (g1331) & (!g937)) + ((g18) & (!g33) & (g74) & (!sk[82]) & (g1331) & (g937)) + ((g18) & (g33) & (!g74) & (!sk[82]) & (!g1331) & (!g937)) + ((g18) & (g33) & (!g74) & (!sk[82]) & (!g1331) & (g937)) + ((g18) & (g33) & (!g74) & (!sk[82]) & (g1331) & (!g937)) + ((g18) & (g33) & (!g74) & (!sk[82]) & (g1331) & (g937)) + ((g18) & (g33) & (!g74) & (sk[82]) & (g1331) & (!g937)) + ((g18) & (g33) & (g74) & (!sk[82]) & (!g1331) & (!g937)) + ((g18) & (g33) & (g74) & (!sk[82]) & (!g1331) & (g937)) + ((g18) & (g33) & (g74) & (!sk[82]) & (g1331) & (!g937)) + ((g18) & (g33) & (g74) & (!sk[82]) & (g1331) & (g937)));
	assign g1333 = (((!g1095) & (!sk[83]) & (!g1005) & (g1329) & (!g1330) & (g1332)) + ((!g1095) & (!sk[83]) & (!g1005) & (g1329) & (g1330) & (!g1332)) + ((!g1095) & (!sk[83]) & (!g1005) & (g1329) & (g1330) & (g1332)) + ((!g1095) & (!sk[83]) & (g1005) & (!g1329) & (!g1330) & (!g1332)) + ((!g1095) & (!sk[83]) & (g1005) & (!g1329) & (!g1330) & (g1332)) + ((!g1095) & (!sk[83]) & (g1005) & (!g1329) & (g1330) & (!g1332)) + ((!g1095) & (!sk[83]) & (g1005) & (!g1329) & (g1330) & (g1332)) + ((!g1095) & (!sk[83]) & (g1005) & (g1329) & (!g1330) & (!g1332)) + ((!g1095) & (!sk[83]) & (g1005) & (g1329) & (!g1330) & (g1332)) + ((!g1095) & (!sk[83]) & (g1005) & (g1329) & (g1330) & (!g1332)) + ((!g1095) & (!sk[83]) & (g1005) & (g1329) & (g1330) & (g1332)) + ((!g1095) & (sk[83]) & (!g1005) & (g1329) & (g1330) & (g1332)) + ((g1095) & (!sk[83]) & (!g1005) & (g1329) & (!g1330) & (g1332)) + ((g1095) & (!sk[83]) & (!g1005) & (g1329) & (g1330) & (!g1332)) + ((g1095) & (!sk[83]) & (!g1005) & (g1329) & (g1330) & (g1332)) + ((g1095) & (!sk[83]) & (g1005) & (!g1329) & (!g1330) & (!g1332)) + ((g1095) & (!sk[83]) & (g1005) & (!g1329) & (!g1330) & (g1332)) + ((g1095) & (!sk[83]) & (g1005) & (!g1329) & (g1330) & (!g1332)) + ((g1095) & (!sk[83]) & (g1005) & (!g1329) & (g1330) & (g1332)) + ((g1095) & (!sk[83]) & (g1005) & (g1329) & (!g1330) & (!g1332)) + ((g1095) & (!sk[83]) & (g1005) & (g1329) & (!g1330) & (g1332)) + ((g1095) & (!sk[83]) & (g1005) & (g1329) & (g1330) & (!g1332)) + ((g1095) & (!sk[83]) & (g1005) & (g1329) & (g1330) & (g1332)));
	assign g1334 = (((!sk[84]) & (!g97) & (!g98) & (g135)) + ((!sk[84]) & (!g97) & (g98) & (!g135)) + ((!sk[84]) & (!g97) & (g98) & (g135)) + ((!sk[84]) & (g97) & (!g98) & (g135)) + ((!sk[84]) & (g97) & (g98) & (!g135)) + ((!sk[84]) & (g97) & (g98) & (g135)) + ((sk[84]) & (!g97) & (!g98) & (!g135)) + ((sk[84]) & (!g97) & (g98) & (!g135)) + ((sk[84]) & (g97) & (g98) & (!g135)));
	assign g1335 = (((!g102) & (!g212) & (!sk[85]) & (g484)) + ((!g102) & (g212) & (!sk[85]) & (!g484)) + ((!g102) & (g212) & (!sk[85]) & (g484)) + ((g102) & (!g212) & (!sk[85]) & (g484)) + ((g102) & (!g212) & (sk[85]) & (g484)) + ((g102) & (g212) & (!sk[85]) & (!g484)) + ((g102) & (g212) & (!sk[85]) & (g484)) + ((g102) & (g212) & (sk[85]) & (!g484)) + ((g102) & (g212) & (sk[85]) & (g484)));
	assign g1336 = (((!i_4_) & (!i_3_) & (!i_5_) & (g71) & (sk[86]) & (g101)) + ((!i_4_) & (!i_3_) & (i_5_) & (!g71) & (!sk[86]) & (g101)) + ((!i_4_) & (!i_3_) & (i_5_) & (g71) & (!sk[86]) & (!g101)) + ((!i_4_) & (!i_3_) & (i_5_) & (g71) & (!sk[86]) & (g101)) + ((!i_4_) & (i_3_) & (!i_5_) & (!g71) & (!sk[86]) & (!g101)) + ((!i_4_) & (i_3_) & (!i_5_) & (!g71) & (!sk[86]) & (g101)) + ((!i_4_) & (i_3_) & (!i_5_) & (g71) & (!sk[86]) & (!g101)) + ((!i_4_) & (i_3_) & (!i_5_) & (g71) & (!sk[86]) & (g101)) + ((!i_4_) & (i_3_) & (i_5_) & (!g71) & (!sk[86]) & (!g101)) + ((!i_4_) & (i_3_) & (i_5_) & (!g71) & (!sk[86]) & (g101)) + ((!i_4_) & (i_3_) & (i_5_) & (g71) & (!sk[86]) & (!g101)) + ((!i_4_) & (i_3_) & (i_5_) & (g71) & (!sk[86]) & (g101)) + ((i_4_) & (!i_3_) & (i_5_) & (!g71) & (!sk[86]) & (g101)) + ((i_4_) & (!i_3_) & (i_5_) & (g71) & (!sk[86]) & (!g101)) + ((i_4_) & (!i_3_) & (i_5_) & (g71) & (!sk[86]) & (g101)) + ((i_4_) & (!i_3_) & (i_5_) & (g71) & (sk[86]) & (g101)) + ((i_4_) & (i_3_) & (!i_5_) & (!g71) & (!sk[86]) & (!g101)) + ((i_4_) & (i_3_) & (!i_5_) & (!g71) & (!sk[86]) & (g101)) + ((i_4_) & (i_3_) & (!i_5_) & (g71) & (!sk[86]) & (!g101)) + ((i_4_) & (i_3_) & (!i_5_) & (g71) & (!sk[86]) & (g101)) + ((i_4_) & (i_3_) & (i_5_) & (!g71) & (!sk[86]) & (!g101)) + ((i_4_) & (i_3_) & (i_5_) & (!g71) & (!sk[86]) & (g101)) + ((i_4_) & (i_3_) & (i_5_) & (g71) & (!sk[86]) & (!g101)) + ((i_4_) & (i_3_) & (i_5_) & (g71) & (!sk[86]) & (g101)));
	assign g1337 = (((!i_9_) & (!sk[87]) & (!i_10_) & (i_11_) & (!g1336)) + ((!i_9_) & (!sk[87]) & (!i_10_) & (i_11_) & (g1336)) + ((!i_9_) & (!sk[87]) & (i_10_) & (i_11_) & (!g1336)) + ((!i_9_) & (!sk[87]) & (i_10_) & (i_11_) & (g1336)) + ((i_9_) & (!sk[87]) & (!i_10_) & (i_11_) & (!g1336)) + ((i_9_) & (!sk[87]) & (!i_10_) & (i_11_) & (g1336)) + ((i_9_) & (!sk[87]) & (i_10_) & (i_11_) & (!g1336)) + ((i_9_) & (!sk[87]) & (i_10_) & (i_11_) & (g1336)) + ((i_9_) & (sk[87]) & (!i_10_) & (!i_11_) & (g1336)));
	assign g1338 = (((!g4) & (!sk[88]) & (!g27) & (g394) & (!g1337)) + ((!g4) & (!sk[88]) & (!g27) & (g394) & (g1337)) + ((!g4) & (!sk[88]) & (g27) & (g394) & (!g1337)) + ((!g4) & (!sk[88]) & (g27) & (g394) & (g1337)) + ((!g4) & (sk[88]) & (!g27) & (g394) & (g1337)) + ((!g4) & (sk[88]) & (g27) & (g394) & (g1337)) + ((g4) & (!sk[88]) & (!g27) & (g394) & (!g1337)) + ((g4) & (!sk[88]) & (!g27) & (g394) & (g1337)) + ((g4) & (!sk[88]) & (g27) & (g394) & (!g1337)) + ((g4) & (!sk[88]) & (g27) & (g394) & (g1337)) + ((g4) & (sk[88]) & (!g27) & (g394) & (g1337)) + ((g4) & (sk[88]) & (g27) & (!g394) & (g1337)) + ((g4) & (sk[88]) & (g27) & (g394) & (g1337)));
	assign g1339 = (((!g18) & (!g33) & (!sk[89]) & (g135) & (!g130) & (g624)) + ((!g18) & (!g33) & (!sk[89]) & (g135) & (g130) & (!g624)) + ((!g18) & (!g33) & (!sk[89]) & (g135) & (g130) & (g624)) + ((!g18) & (!g33) & (sk[89]) & (!g135) & (!g130) & (g624)) + ((!g18) & (!g33) & (sk[89]) & (!g135) & (g130) & (!g624)) + ((!g18) & (!g33) & (sk[89]) & (!g135) & (g130) & (g624)) + ((!g18) & (!g33) & (sk[89]) & (g135) & (!g130) & (g624)) + ((!g18) & (!g33) & (sk[89]) & (g135) & (g130) & (!g624)) + ((!g18) & (!g33) & (sk[89]) & (g135) & (g130) & (g624)) + ((!g18) & (g33) & (!sk[89]) & (!g135) & (!g130) & (!g624)) + ((!g18) & (g33) & (!sk[89]) & (!g135) & (!g130) & (g624)) + ((!g18) & (g33) & (!sk[89]) & (!g135) & (g130) & (!g624)) + ((!g18) & (g33) & (!sk[89]) & (!g135) & (g130) & (g624)) + ((!g18) & (g33) & (!sk[89]) & (g135) & (!g130) & (!g624)) + ((!g18) & (g33) & (!sk[89]) & (g135) & (!g130) & (g624)) + ((!g18) & (g33) & (!sk[89]) & (g135) & (g130) & (!g624)) + ((!g18) & (g33) & (!sk[89]) & (g135) & (g130) & (g624)) + ((!g18) & (g33) & (sk[89]) & (g135) & (!g130) & (g624)) + ((!g18) & (g33) & (sk[89]) & (g135) & (g130) & (!g624)) + ((!g18) & (g33) & (sk[89]) & (g135) & (g130) & (g624)) + ((g18) & (!g33) & (!sk[89]) & (g135) & (!g130) & (g624)) + ((g18) & (!g33) & (!sk[89]) & (g135) & (g130) & (!g624)) + ((g18) & (!g33) & (!sk[89]) & (g135) & (g130) & (g624)) + ((g18) & (!g33) & (sk[89]) & (g135) & (!g130) & (g624)) + ((g18) & (!g33) & (sk[89]) & (g135) & (g130) & (!g624)) + ((g18) & (!g33) & (sk[89]) & (g135) & (g130) & (g624)) + ((g18) & (g33) & (!sk[89]) & (!g135) & (!g130) & (!g624)) + ((g18) & (g33) & (!sk[89]) & (!g135) & (!g130) & (g624)) + ((g18) & (g33) & (!sk[89]) & (!g135) & (g130) & (!g624)) + ((g18) & (g33) & (!sk[89]) & (!g135) & (g130) & (g624)) + ((g18) & (g33) & (!sk[89]) & (g135) & (!g130) & (!g624)) + ((g18) & (g33) & (!sk[89]) & (g135) & (!g130) & (g624)) + ((g18) & (g33) & (!sk[89]) & (g135) & (g130) & (!g624)) + ((g18) & (g33) & (!sk[89]) & (g135) & (g130) & (g624)) + ((g18) & (g33) & (sk[89]) & (g135) & (!g130) & (g624)) + ((g18) & (g33) & (sk[89]) & (g135) & (g130) & (!g624)) + ((g18) & (g33) & (sk[89]) & (g135) & (g130) & (g624)));
	assign g1340 = (((!g1334) & (!g383) & (!g993) & (!g1335) & (!g1338) & (g1339)) + ((!g1334) & (g383) & (!g993) & (!g1335) & (!g1338) & (g1339)) + ((!g1334) & (g383) & (g993) & (!g1335) & (!g1338) & (g1339)));
	assign g1341 = (((!g179) & (!sk[91]) & (!g461) & (g605) & (!g487)) + ((!g179) & (!sk[91]) & (!g461) & (g605) & (g487)) + ((!g179) & (!sk[91]) & (g461) & (g605) & (!g487)) + ((!g179) & (!sk[91]) & (g461) & (g605) & (g487)) + ((!g179) & (sk[91]) & (!g461) & (!g605) & (!g487)) + ((g179) & (!sk[91]) & (!g461) & (g605) & (!g487)) + ((g179) & (!sk[91]) & (!g461) & (g605) & (g487)) + ((g179) & (!sk[91]) & (g461) & (g605) & (!g487)) + ((g179) & (!sk[91]) & (g461) & (g605) & (g487)));
	assign g1342 = (((!g135) & (!g313) & (!sk[92]) & (g477) & (!g1341) & (g990)) + ((!g135) & (!g313) & (!sk[92]) & (g477) & (g1341) & (!g990)) + ((!g135) & (!g313) & (!sk[92]) & (g477) & (g1341) & (g990)) + ((!g135) & (!g313) & (sk[92]) & (!g477) & (g1341) & (!g990)) + ((!g135) & (!g313) & (sk[92]) & (g477) & (g1341) & (!g990)) + ((!g135) & (g313) & (!sk[92]) & (!g477) & (!g1341) & (!g990)) + ((!g135) & (g313) & (!sk[92]) & (!g477) & (!g1341) & (g990)) + ((!g135) & (g313) & (!sk[92]) & (!g477) & (g1341) & (!g990)) + ((!g135) & (g313) & (!sk[92]) & (!g477) & (g1341) & (g990)) + ((!g135) & (g313) & (!sk[92]) & (g477) & (!g1341) & (!g990)) + ((!g135) & (g313) & (!sk[92]) & (g477) & (!g1341) & (g990)) + ((!g135) & (g313) & (!sk[92]) & (g477) & (g1341) & (!g990)) + ((!g135) & (g313) & (!sk[92]) & (g477) & (g1341) & (g990)) + ((!g135) & (g313) & (sk[92]) & (!g477) & (g1341) & (!g990)) + ((g135) & (!g313) & (!sk[92]) & (g477) & (!g1341) & (g990)) + ((g135) & (!g313) & (!sk[92]) & (g477) & (g1341) & (!g990)) + ((g135) & (!g313) & (!sk[92]) & (g477) & (g1341) & (g990)) + ((g135) & (!g313) & (sk[92]) & (!g477) & (!g1341) & (!g990)) + ((g135) & (!g313) & (sk[92]) & (!g477) & (g1341) & (!g990)) + ((g135) & (!g313) & (sk[92]) & (g477) & (!g1341) & (!g990)) + ((g135) & (!g313) & (sk[92]) & (g477) & (g1341) & (!g990)) + ((g135) & (g313) & (!sk[92]) & (!g477) & (!g1341) & (!g990)) + ((g135) & (g313) & (!sk[92]) & (!g477) & (!g1341) & (g990)) + ((g135) & (g313) & (!sk[92]) & (!g477) & (g1341) & (!g990)) + ((g135) & (g313) & (!sk[92]) & (!g477) & (g1341) & (g990)) + ((g135) & (g313) & (!sk[92]) & (g477) & (!g1341) & (!g990)) + ((g135) & (g313) & (!sk[92]) & (g477) & (!g1341) & (g990)) + ((g135) & (g313) & (!sk[92]) & (g477) & (g1341) & (!g990)) + ((g135) & (g313) & (!sk[92]) & (g477) & (g1341) & (g990)) + ((g135) & (g313) & (sk[92]) & (!g477) & (!g1341) & (!g990)) + ((g135) & (g313) & (sk[92]) & (!g477) & (g1341) & (!g990)));
	assign g1343 = (((!g97) & (!g98) & (!g74) & (!g257) & (sk[93]) & (!g489)) + ((!g97) & (!g98) & (!g74) & (!g257) & (sk[93]) & (g489)) + ((!g97) & (!g98) & (!g74) & (g257) & (sk[93]) & (!g489)) + ((!g97) & (!g98) & (g74) & (!g257) & (!sk[93]) & (g489)) + ((!g97) & (!g98) & (g74) & (g257) & (!sk[93]) & (!g489)) + ((!g97) & (!g98) & (g74) & (g257) & (!sk[93]) & (g489)) + ((!g97) & (g98) & (!g74) & (!g257) & (!sk[93]) & (!g489)) + ((!g97) & (g98) & (!g74) & (!g257) & (!sk[93]) & (g489)) + ((!g97) & (g98) & (!g74) & (!g257) & (sk[93]) & (!g489)) + ((!g97) & (g98) & (!g74) & (!g257) & (sk[93]) & (g489)) + ((!g97) & (g98) & (!g74) & (g257) & (!sk[93]) & (!g489)) + ((!g97) & (g98) & (!g74) & (g257) & (!sk[93]) & (g489)) + ((!g97) & (g98) & (!g74) & (g257) & (sk[93]) & (!g489)) + ((!g97) & (g98) & (g74) & (!g257) & (!sk[93]) & (!g489)) + ((!g97) & (g98) & (g74) & (!g257) & (!sk[93]) & (g489)) + ((!g97) & (g98) & (g74) & (g257) & (!sk[93]) & (!g489)) + ((!g97) & (g98) & (g74) & (g257) & (!sk[93]) & (g489)) + ((g97) & (!g98) & (!g74) & (!g257) & (sk[93]) & (!g489)) + ((g97) & (!g98) & (!g74) & (!g257) & (sk[93]) & (g489)) + ((g97) & (!g98) & (!g74) & (g257) & (sk[93]) & (!g489)) + ((g97) & (!g98) & (g74) & (!g257) & (!sk[93]) & (g489)) + ((g97) & (!g98) & (g74) & (!g257) & (sk[93]) & (!g489)) + ((g97) & (!g98) & (g74) & (g257) & (!sk[93]) & (!g489)) + ((g97) & (!g98) & (g74) & (g257) & (!sk[93]) & (g489)) + ((g97) & (!g98) & (g74) & (g257) & (sk[93]) & (!g489)) + ((g97) & (g98) & (!g74) & (!g257) & (!sk[93]) & (!g489)) + ((g97) & (g98) & (!g74) & (!g257) & (!sk[93]) & (g489)) + ((g97) & (g98) & (!g74) & (!g257) & (sk[93]) & (!g489)) + ((g97) & (g98) & (!g74) & (!g257) & (sk[93]) & (g489)) + ((g97) & (g98) & (!g74) & (g257) & (!sk[93]) & (!g489)) + ((g97) & (g98) & (!g74) & (g257) & (!sk[93]) & (g489)) + ((g97) & (g98) & (!g74) & (g257) & (sk[93]) & (!g489)) + ((g97) & (g98) & (g74) & (!g257) & (!sk[93]) & (!g489)) + ((g97) & (g98) & (g74) & (!g257) & (!sk[93]) & (g489)) + ((g97) & (g98) & (g74) & (g257) & (!sk[93]) & (!g489)) + ((g97) & (g98) & (g74) & (g257) & (!sk[93]) & (g489)));
	assign g1344 = (((!g1027) & (!sk[94]) & (!g995) & (g1340) & (!g1342) & (g1343)) + ((!g1027) & (!sk[94]) & (!g995) & (g1340) & (g1342) & (!g1343)) + ((!g1027) & (!sk[94]) & (!g995) & (g1340) & (g1342) & (g1343)) + ((!g1027) & (!sk[94]) & (g995) & (!g1340) & (!g1342) & (!g1343)) + ((!g1027) & (!sk[94]) & (g995) & (!g1340) & (!g1342) & (g1343)) + ((!g1027) & (!sk[94]) & (g995) & (!g1340) & (g1342) & (!g1343)) + ((!g1027) & (!sk[94]) & (g995) & (!g1340) & (g1342) & (g1343)) + ((!g1027) & (!sk[94]) & (g995) & (g1340) & (!g1342) & (!g1343)) + ((!g1027) & (!sk[94]) & (g995) & (g1340) & (!g1342) & (g1343)) + ((!g1027) & (!sk[94]) & (g995) & (g1340) & (g1342) & (!g1343)) + ((!g1027) & (!sk[94]) & (g995) & (g1340) & (g1342) & (g1343)) + ((!g1027) & (sk[94]) & (g995) & (g1340) & (g1342) & (g1343)) + ((g1027) & (!sk[94]) & (!g995) & (g1340) & (!g1342) & (g1343)) + ((g1027) & (!sk[94]) & (!g995) & (g1340) & (g1342) & (!g1343)) + ((g1027) & (!sk[94]) & (!g995) & (g1340) & (g1342) & (g1343)) + ((g1027) & (!sk[94]) & (g995) & (!g1340) & (!g1342) & (!g1343)) + ((g1027) & (!sk[94]) & (g995) & (!g1340) & (!g1342) & (g1343)) + ((g1027) & (!sk[94]) & (g995) & (!g1340) & (g1342) & (!g1343)) + ((g1027) & (!sk[94]) & (g995) & (!g1340) & (g1342) & (g1343)) + ((g1027) & (!sk[94]) & (g995) & (g1340) & (!g1342) & (!g1343)) + ((g1027) & (!sk[94]) & (g995) & (g1340) & (!g1342) & (g1343)) + ((g1027) & (!sk[94]) & (g995) & (g1340) & (g1342) & (!g1343)) + ((g1027) & (!sk[94]) & (g995) & (g1340) & (g1342) & (g1343)));
	assign g1345 = (((!g955) & (!sk[95]) & (!g982) & (g1324) & (!g1333) & (g1344)) + ((!g955) & (!sk[95]) & (!g982) & (g1324) & (g1333) & (!g1344)) + ((!g955) & (!sk[95]) & (!g982) & (g1324) & (g1333) & (g1344)) + ((!g955) & (!sk[95]) & (g982) & (!g1324) & (!g1333) & (!g1344)) + ((!g955) & (!sk[95]) & (g982) & (!g1324) & (!g1333) & (g1344)) + ((!g955) & (!sk[95]) & (g982) & (!g1324) & (g1333) & (!g1344)) + ((!g955) & (!sk[95]) & (g982) & (!g1324) & (g1333) & (g1344)) + ((!g955) & (!sk[95]) & (g982) & (g1324) & (!g1333) & (!g1344)) + ((!g955) & (!sk[95]) & (g982) & (g1324) & (!g1333) & (g1344)) + ((!g955) & (!sk[95]) & (g982) & (g1324) & (g1333) & (!g1344)) + ((!g955) & (!sk[95]) & (g982) & (g1324) & (g1333) & (g1344)) + ((g955) & (!sk[95]) & (!g982) & (g1324) & (!g1333) & (g1344)) + ((g955) & (!sk[95]) & (!g982) & (g1324) & (g1333) & (!g1344)) + ((g955) & (!sk[95]) & (!g982) & (g1324) & (g1333) & (g1344)) + ((g955) & (!sk[95]) & (g982) & (!g1324) & (!g1333) & (!g1344)) + ((g955) & (!sk[95]) & (g982) & (!g1324) & (!g1333) & (g1344)) + ((g955) & (!sk[95]) & (g982) & (!g1324) & (g1333) & (!g1344)) + ((g955) & (!sk[95]) & (g982) & (!g1324) & (g1333) & (g1344)) + ((g955) & (!sk[95]) & (g982) & (g1324) & (!g1333) & (!g1344)) + ((g955) & (!sk[95]) & (g982) & (g1324) & (!g1333) & (g1344)) + ((g955) & (!sk[95]) & (g982) & (g1324) & (g1333) & (!g1344)) + ((g955) & (!sk[95]) & (g982) & (g1324) & (g1333) & (g1344)) + ((g955) & (sk[95]) & (g982) & (g1324) & (g1333) & (g1344)));
	assign g1346 = (((g1172) & (g1183) & (g1207) & (g1295) & (g1319) & (g1345)));
	assign g1347 = (((!g123) & (!sk[97]) & (!g852) & (g853)) + ((!g123) & (!sk[97]) & (g852) & (!g853)) + ((!g123) & (!sk[97]) & (g852) & (g853)) + ((!g123) & (sk[97]) & (!g852) & (g853)) + ((!g123) & (sk[97]) & (g852) & (!g853)) + ((!g123) & (sk[97]) & (g852) & (g853)) + ((g123) & (!sk[97]) & (!g852) & (g853)) + ((g123) & (!sk[97]) & (g852) & (!g853)) + ((g123) & (!sk[97]) & (g852) & (g853)));
	assign g1348 = (((!g113) & (!g174) & (!g408) & (sk[98]) & (!g857)) + ((!g113) & (!g174) & (!g408) & (sk[98]) & (g857)) + ((!g113) & (!g174) & (g408) & (!sk[98]) & (!g857)) + ((!g113) & (!g174) & (g408) & (!sk[98]) & (g857)) + ((!g113) & (g174) & (!g408) & (sk[98]) & (g857)) + ((!g113) & (g174) & (g408) & (!sk[98]) & (!g857)) + ((!g113) & (g174) & (g408) & (!sk[98]) & (g857)) + ((g113) & (!g174) & (!g408) & (sk[98]) & (g857)) + ((g113) & (!g174) & (g408) & (!sk[98]) & (!g857)) + ((g113) & (!g174) & (g408) & (!sk[98]) & (g857)) + ((g113) & (g174) & (!g408) & (sk[98]) & (g857)) + ((g113) & (g174) & (g408) & (!sk[98]) & (!g857)) + ((g113) & (g174) & (g408) & (!sk[98]) & (g857)));
	assign g1349 = (((!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g112) & (!g123)) + ((i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g112) & (!g123)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g112) & (!g123)) + ((i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g112) & (!g123)));
	assign g1350 = (((!g130) & (!sk[100]) & (!g742) & (g1347) & (!g1348) & (g1349)) + ((!g130) & (!sk[100]) & (!g742) & (g1347) & (g1348) & (!g1349)) + ((!g130) & (!sk[100]) & (!g742) & (g1347) & (g1348) & (g1349)) + ((!g130) & (!sk[100]) & (g742) & (!g1347) & (!g1348) & (!g1349)) + ((!g130) & (!sk[100]) & (g742) & (!g1347) & (!g1348) & (g1349)) + ((!g130) & (!sk[100]) & (g742) & (!g1347) & (g1348) & (!g1349)) + ((!g130) & (!sk[100]) & (g742) & (!g1347) & (g1348) & (g1349)) + ((!g130) & (!sk[100]) & (g742) & (g1347) & (!g1348) & (!g1349)) + ((!g130) & (!sk[100]) & (g742) & (g1347) & (!g1348) & (g1349)) + ((!g130) & (!sk[100]) & (g742) & (g1347) & (g1348) & (!g1349)) + ((!g130) & (!sk[100]) & (g742) & (g1347) & (g1348) & (g1349)) + ((!g130) & (sk[100]) & (g742) & (!g1347) & (!g1348) & (!g1349)) + ((g130) & (!sk[100]) & (!g742) & (g1347) & (!g1348) & (g1349)) + ((g130) & (!sk[100]) & (!g742) & (g1347) & (g1348) & (!g1349)) + ((g130) & (!sk[100]) & (!g742) & (g1347) & (g1348) & (g1349)) + ((g130) & (!sk[100]) & (g742) & (!g1347) & (!g1348) & (!g1349)) + ((g130) & (!sk[100]) & (g742) & (!g1347) & (!g1348) & (g1349)) + ((g130) & (!sk[100]) & (g742) & (!g1347) & (g1348) & (!g1349)) + ((g130) & (!sk[100]) & (g742) & (!g1347) & (g1348) & (g1349)) + ((g130) & (!sk[100]) & (g742) & (g1347) & (!g1348) & (!g1349)) + ((g130) & (!sk[100]) & (g742) & (g1347) & (!g1348) & (g1349)) + ((g130) & (!sk[100]) & (g742) & (g1347) & (g1348) & (!g1349)) + ((g130) & (!sk[100]) & (g742) & (g1347) & (g1348) & (g1349)) + ((g130) & (sk[100]) & (!g742) & (!g1347) & (!g1348) & (!g1349)) + ((g130) & (sk[100]) & (g742) & (!g1347) & (!g1348) & (!g1349)));
	assign g1351 = (((!g123) & (!sk[101]) & (!g113) & (g130) & (!g507) & (g974)) + ((!g123) & (!sk[101]) & (!g113) & (g130) & (g507) & (!g974)) + ((!g123) & (!sk[101]) & (!g113) & (g130) & (g507) & (g974)) + ((!g123) & (!sk[101]) & (g113) & (!g130) & (!g507) & (!g974)) + ((!g123) & (!sk[101]) & (g113) & (!g130) & (!g507) & (g974)) + ((!g123) & (!sk[101]) & (g113) & (!g130) & (g507) & (!g974)) + ((!g123) & (!sk[101]) & (g113) & (!g130) & (g507) & (g974)) + ((!g123) & (!sk[101]) & (g113) & (g130) & (!g507) & (!g974)) + ((!g123) & (!sk[101]) & (g113) & (g130) & (!g507) & (g974)) + ((!g123) & (!sk[101]) & (g113) & (g130) & (g507) & (!g974)) + ((!g123) & (!sk[101]) & (g113) & (g130) & (g507) & (g974)) + ((!g123) & (sk[101]) & (!g113) & (!g130) & (!g507) & (g974)) + ((!g123) & (sk[101]) & (!g113) & (!g130) & (g507) & (!g974)) + ((!g123) & (sk[101]) & (!g113) & (!g130) & (g507) & (g974)) + ((!g123) & (sk[101]) & (!g113) & (g130) & (!g507) & (g974)) + ((!g123) & (sk[101]) & (!g113) & (g130) & (g507) & (g974)) + ((!g123) & (sk[101]) & (g113) & (!g130) & (!g507) & (g974)) + ((!g123) & (sk[101]) & (g113) & (!g130) & (g507) & (g974)) + ((!g123) & (sk[101]) & (g113) & (g130) & (!g507) & (g974)) + ((!g123) & (sk[101]) & (g113) & (g130) & (g507) & (g974)) + ((g123) & (!sk[101]) & (!g113) & (g130) & (!g507) & (g974)) + ((g123) & (!sk[101]) & (!g113) & (g130) & (g507) & (!g974)) + ((g123) & (!sk[101]) & (!g113) & (g130) & (g507) & (g974)) + ((g123) & (!sk[101]) & (g113) & (!g130) & (!g507) & (!g974)) + ((g123) & (!sk[101]) & (g113) & (!g130) & (!g507) & (g974)) + ((g123) & (!sk[101]) & (g113) & (!g130) & (g507) & (!g974)) + ((g123) & (!sk[101]) & (g113) & (!g130) & (g507) & (g974)) + ((g123) & (!sk[101]) & (g113) & (g130) & (!g507) & (!g974)) + ((g123) & (!sk[101]) & (g113) & (g130) & (!g507) & (g974)) + ((g123) & (!sk[101]) & (g113) & (g130) & (g507) & (!g974)) + ((g123) & (!sk[101]) & (g113) & (g130) & (g507) & (g974)) + ((g123) & (sk[101]) & (!g113) & (!g130) & (!g507) & (g974)) + ((g123) & (sk[101]) & (!g113) & (!g130) & (g507) & (!g974)) + ((g123) & (sk[101]) & (!g113) & (!g130) & (g507) & (g974)) + ((g123) & (sk[101]) & (g113) & (!g130) & (!g507) & (g974)) + ((g123) & (sk[101]) & (g113) & (!g130) & (g507) & (g974)));
	assign g1352 = (((!g24) & (!g113) & (!sk[102]) & (g408) & (!g1350) & (g1351)) + ((!g24) & (!g113) & (!sk[102]) & (g408) & (g1350) & (!g1351)) + ((!g24) & (!g113) & (!sk[102]) & (g408) & (g1350) & (g1351)) + ((!g24) & (!g113) & (sk[102]) & (g408) & (g1350) & (!g1351)) + ((!g24) & (g113) & (!sk[102]) & (!g408) & (!g1350) & (!g1351)) + ((!g24) & (g113) & (!sk[102]) & (!g408) & (!g1350) & (g1351)) + ((!g24) & (g113) & (!sk[102]) & (!g408) & (g1350) & (!g1351)) + ((!g24) & (g113) & (!sk[102]) & (!g408) & (g1350) & (g1351)) + ((!g24) & (g113) & (!sk[102]) & (g408) & (!g1350) & (!g1351)) + ((!g24) & (g113) & (!sk[102]) & (g408) & (!g1350) & (g1351)) + ((!g24) & (g113) & (!sk[102]) & (g408) & (g1350) & (!g1351)) + ((!g24) & (g113) & (!sk[102]) & (g408) & (g1350) & (g1351)) + ((!g24) & (g113) & (sk[102]) & (!g408) & (g1350) & (!g1351)) + ((!g24) & (g113) & (sk[102]) & (g408) & (g1350) & (!g1351)) + ((g24) & (!g113) & (!sk[102]) & (g408) & (!g1350) & (g1351)) + ((g24) & (!g113) & (!sk[102]) & (g408) & (g1350) & (!g1351)) + ((g24) & (!g113) & (!sk[102]) & (g408) & (g1350) & (g1351)) + ((g24) & (!g113) & (sk[102]) & (!g408) & (g1350) & (!g1351)) + ((g24) & (!g113) & (sk[102]) & (g408) & (g1350) & (!g1351)) + ((g24) & (g113) & (!sk[102]) & (!g408) & (!g1350) & (!g1351)) + ((g24) & (g113) & (!sk[102]) & (!g408) & (!g1350) & (g1351)) + ((g24) & (g113) & (!sk[102]) & (!g408) & (g1350) & (!g1351)) + ((g24) & (g113) & (!sk[102]) & (!g408) & (g1350) & (g1351)) + ((g24) & (g113) & (!sk[102]) & (g408) & (!g1350) & (!g1351)) + ((g24) & (g113) & (!sk[102]) & (g408) & (!g1350) & (g1351)) + ((g24) & (g113) & (!sk[102]) & (g408) & (g1350) & (!g1351)) + ((g24) & (g113) & (!sk[102]) & (g408) & (g1350) & (g1351)) + ((g24) & (g113) & (sk[102]) & (!g408) & (g1350) & (!g1351)) + ((g24) & (g113) & (sk[102]) & (g408) & (g1350) & (!g1351)));
	assign g1353 = (((!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (!g73) & (g112)) + ((!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g73) & (g112)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g73) & (g112)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g73) & (g112)) + ((!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g73) & (g112)) + ((!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g73) & (g112)) + ((i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (!g73) & (g112)) + ((i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g73) & (g112)) + ((i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g73) & (g112)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g73) & (g112)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g73) & (g112)) + ((i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g73) & (g112)) + ((i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g73) & (g112)) + ((i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g73) & (g112)) + ((i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g73) & (g112)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g73) & (g112)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g73) & (g112)) + ((i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g73) & (g112)) + ((i_15_) & (i_12_) & (i_13_) & (i_14_) & (g73) & (g112)));
	assign g1354 = (((!g10) & (!g72) & (g101) & (!sk[104]) & (!g1102)) + ((!g10) & (!g72) & (g101) & (!sk[104]) & (g1102)) + ((!g10) & (g72) & (g101) & (!sk[104]) & (!g1102)) + ((!g10) & (g72) & (g101) & (!sk[104]) & (g1102)) + ((!g10) & (g72) & (g101) & (sk[104]) & (!g1102)) + ((!g10) & (g72) & (g101) & (sk[104]) & (g1102)) + ((g10) & (!g72) & (g101) & (!sk[104]) & (!g1102)) + ((g10) & (!g72) & (g101) & (!sk[104]) & (g1102)) + ((g10) & (g72) & (!g101) & (sk[104]) & (g1102)) + ((g10) & (g72) & (g101) & (!sk[104]) & (!g1102)) + ((g10) & (g72) & (g101) & (!sk[104]) & (g1102)) + ((g10) & (g72) & (g101) & (sk[104]) & (!g1102)) + ((g10) & (g72) & (g101) & (sk[104]) & (g1102)));
	assign g1355 = (((!i_8_) & (!g73) & (g125) & (!sk[105]) & (!g857) & (g1029)) + ((!i_8_) & (!g73) & (g125) & (!sk[105]) & (g857) & (!g1029)) + ((!i_8_) & (!g73) & (g125) & (!sk[105]) & (g857) & (g1029)) + ((!i_8_) & (!g73) & (g125) & (sk[105]) & (g857) & (!g1029)) + ((!i_8_) & (!g73) & (g125) & (sk[105]) & (g857) & (g1029)) + ((!i_8_) & (g73) & (!g125) & (!sk[105]) & (!g857) & (!g1029)) + ((!i_8_) & (g73) & (!g125) & (!sk[105]) & (!g857) & (g1029)) + ((!i_8_) & (g73) & (!g125) & (!sk[105]) & (g857) & (!g1029)) + ((!i_8_) & (g73) & (!g125) & (!sk[105]) & (g857) & (g1029)) + ((!i_8_) & (g73) & (!g125) & (sk[105]) & (g857) & (!g1029)) + ((!i_8_) & (g73) & (!g125) & (sk[105]) & (g857) & (g1029)) + ((!i_8_) & (g73) & (g125) & (!sk[105]) & (!g857) & (!g1029)) + ((!i_8_) & (g73) & (g125) & (!sk[105]) & (!g857) & (g1029)) + ((!i_8_) & (g73) & (g125) & (!sk[105]) & (g857) & (!g1029)) + ((!i_8_) & (g73) & (g125) & (!sk[105]) & (g857) & (g1029)) + ((!i_8_) & (g73) & (g125) & (sk[105]) & (g857) & (!g1029)) + ((!i_8_) & (g73) & (g125) & (sk[105]) & (g857) & (g1029)) + ((i_8_) & (!g73) & (g125) & (!sk[105]) & (!g857) & (g1029)) + ((i_8_) & (!g73) & (g125) & (!sk[105]) & (g857) & (!g1029)) + ((i_8_) & (!g73) & (g125) & (!sk[105]) & (g857) & (g1029)) + ((i_8_) & (!g73) & (g125) & (sk[105]) & (g857) & (!g1029)) + ((i_8_) & (!g73) & (g125) & (sk[105]) & (g857) & (g1029)) + ((i_8_) & (g73) & (!g125) & (!sk[105]) & (!g857) & (!g1029)) + ((i_8_) & (g73) & (!g125) & (!sk[105]) & (!g857) & (g1029)) + ((i_8_) & (g73) & (!g125) & (!sk[105]) & (g857) & (!g1029)) + ((i_8_) & (g73) & (!g125) & (!sk[105]) & (g857) & (g1029)) + ((i_8_) & (g73) & (!g125) & (sk[105]) & (!g857) & (!g1029)) + ((i_8_) & (g73) & (!g125) & (sk[105]) & (g857) & (!g1029)) + ((i_8_) & (g73) & (g125) & (!sk[105]) & (!g857) & (!g1029)) + ((i_8_) & (g73) & (g125) & (!sk[105]) & (!g857) & (g1029)) + ((i_8_) & (g73) & (g125) & (!sk[105]) & (g857) & (!g1029)) + ((i_8_) & (g73) & (g125) & (!sk[105]) & (g857) & (g1029)) + ((i_8_) & (g73) & (g125) & (sk[105]) & (!g857) & (!g1029)) + ((i_8_) & (g73) & (g125) & (sk[105]) & (g857) & (!g1029)) + ((i_8_) & (g73) & (g125) & (sk[105]) & (g857) & (g1029)));
	assign g1356 = (((g102) & (!g200) & (!g212) & (!g484) & (!g684) & (!g881)) + ((g102) & (!g200) & (!g212) & (!g484) & (!g684) & (g881)) + ((g102) & (!g200) & (!g212) & (!g484) & (g684) & (g881)) + ((g102) & (!g200) & (!g212) & (g484) & (!g684) & (!g881)) + ((g102) & (!g200) & (!g212) & (g484) & (!g684) & (g881)) + ((g102) & (!g200) & (!g212) & (g484) & (g684) & (!g881)) + ((g102) & (!g200) & (!g212) & (g484) & (g684) & (g881)) + ((g102) & (!g200) & (g212) & (!g484) & (!g684) & (!g881)) + ((g102) & (!g200) & (g212) & (!g484) & (!g684) & (g881)) + ((g102) & (!g200) & (g212) & (!g484) & (g684) & (!g881)) + ((g102) & (!g200) & (g212) & (!g484) & (g684) & (g881)) + ((g102) & (!g200) & (g212) & (g484) & (!g684) & (!g881)) + ((g102) & (!g200) & (g212) & (g484) & (!g684) & (g881)) + ((g102) & (!g200) & (g212) & (g484) & (g684) & (!g881)) + ((g102) & (!g200) & (g212) & (g484) & (g684) & (g881)) + ((g102) & (g200) & (!g212) & (!g484) & (!g684) & (!g881)) + ((g102) & (g200) & (!g212) & (!g484) & (!g684) & (g881)) + ((g102) & (g200) & (!g212) & (!g484) & (g684) & (!g881)) + ((g102) & (g200) & (!g212) & (!g484) & (g684) & (g881)) + ((g102) & (g200) & (!g212) & (g484) & (!g684) & (!g881)) + ((g102) & (g200) & (!g212) & (g484) & (!g684) & (g881)) + ((g102) & (g200) & (!g212) & (g484) & (g684) & (!g881)) + ((g102) & (g200) & (!g212) & (g484) & (g684) & (g881)) + ((g102) & (g200) & (g212) & (!g484) & (!g684) & (!g881)) + ((g102) & (g200) & (g212) & (!g484) & (!g684) & (g881)) + ((g102) & (g200) & (g212) & (!g484) & (g684) & (!g881)) + ((g102) & (g200) & (g212) & (!g484) & (g684) & (g881)) + ((g102) & (g200) & (g212) & (g484) & (!g684) & (!g881)) + ((g102) & (g200) & (g212) & (g484) & (!g684) & (g881)) + ((g102) & (g200) & (g212) & (g484) & (g684) & (!g881)) + ((g102) & (g200) & (g212) & (g484) & (g684) & (g881)));
	assign g1357 = (((!sk[107]) & (!g105) & (!g984) & (g943) & (!g957) & (g1356)) + ((!sk[107]) & (!g105) & (!g984) & (g943) & (g957) & (!g1356)) + ((!sk[107]) & (!g105) & (!g984) & (g943) & (g957) & (g1356)) + ((!sk[107]) & (!g105) & (g984) & (!g943) & (!g957) & (!g1356)) + ((!sk[107]) & (!g105) & (g984) & (!g943) & (!g957) & (g1356)) + ((!sk[107]) & (!g105) & (g984) & (!g943) & (g957) & (!g1356)) + ((!sk[107]) & (!g105) & (g984) & (!g943) & (g957) & (g1356)) + ((!sk[107]) & (!g105) & (g984) & (g943) & (!g957) & (!g1356)) + ((!sk[107]) & (!g105) & (g984) & (g943) & (!g957) & (g1356)) + ((!sk[107]) & (!g105) & (g984) & (g943) & (g957) & (!g1356)) + ((!sk[107]) & (!g105) & (g984) & (g943) & (g957) & (g1356)) + ((!sk[107]) & (g105) & (!g984) & (g943) & (!g957) & (g1356)) + ((!sk[107]) & (g105) & (!g984) & (g943) & (g957) & (!g1356)) + ((!sk[107]) & (g105) & (!g984) & (g943) & (g957) & (g1356)) + ((!sk[107]) & (g105) & (g984) & (!g943) & (!g957) & (!g1356)) + ((!sk[107]) & (g105) & (g984) & (!g943) & (!g957) & (g1356)) + ((!sk[107]) & (g105) & (g984) & (!g943) & (g957) & (!g1356)) + ((!sk[107]) & (g105) & (g984) & (!g943) & (g957) & (g1356)) + ((!sk[107]) & (g105) & (g984) & (g943) & (!g957) & (!g1356)) + ((!sk[107]) & (g105) & (g984) & (g943) & (!g957) & (g1356)) + ((!sk[107]) & (g105) & (g984) & (g943) & (g957) & (!g1356)) + ((!sk[107]) & (g105) & (g984) & (g943) & (g957) & (g1356)) + ((sk[107]) & (!g105) & (!g984) & (!g943) & (!g957) & (!g1356)) + ((sk[107]) & (g105) & (!g984) & (!g943) & (!g957) & (!g1356)) + ((sk[107]) & (g105) & (g984) & (!g943) & (!g957) & (!g1356)));
	assign g1358 = (((!sk[108]) & (!g940) & (!g1353) & (g1354) & (!g1355) & (g1357)) + ((!sk[108]) & (!g940) & (!g1353) & (g1354) & (g1355) & (!g1357)) + ((!sk[108]) & (!g940) & (!g1353) & (g1354) & (g1355) & (g1357)) + ((!sk[108]) & (!g940) & (g1353) & (!g1354) & (!g1355) & (!g1357)) + ((!sk[108]) & (!g940) & (g1353) & (!g1354) & (!g1355) & (g1357)) + ((!sk[108]) & (!g940) & (g1353) & (!g1354) & (g1355) & (!g1357)) + ((!sk[108]) & (!g940) & (g1353) & (!g1354) & (g1355) & (g1357)) + ((!sk[108]) & (!g940) & (g1353) & (g1354) & (!g1355) & (!g1357)) + ((!sk[108]) & (!g940) & (g1353) & (g1354) & (!g1355) & (g1357)) + ((!sk[108]) & (!g940) & (g1353) & (g1354) & (g1355) & (!g1357)) + ((!sk[108]) & (!g940) & (g1353) & (g1354) & (g1355) & (g1357)) + ((!sk[108]) & (g940) & (!g1353) & (g1354) & (!g1355) & (g1357)) + ((!sk[108]) & (g940) & (!g1353) & (g1354) & (g1355) & (!g1357)) + ((!sk[108]) & (g940) & (!g1353) & (g1354) & (g1355) & (g1357)) + ((!sk[108]) & (g940) & (g1353) & (!g1354) & (!g1355) & (!g1357)) + ((!sk[108]) & (g940) & (g1353) & (!g1354) & (!g1355) & (g1357)) + ((!sk[108]) & (g940) & (g1353) & (!g1354) & (g1355) & (!g1357)) + ((!sk[108]) & (g940) & (g1353) & (!g1354) & (g1355) & (g1357)) + ((!sk[108]) & (g940) & (g1353) & (g1354) & (!g1355) & (!g1357)) + ((!sk[108]) & (g940) & (g1353) & (g1354) & (!g1355) & (g1357)) + ((!sk[108]) & (g940) & (g1353) & (g1354) & (g1355) & (!g1357)) + ((!sk[108]) & (g940) & (g1353) & (g1354) & (g1355) & (g1357)) + ((sk[108]) & (g940) & (!g1353) & (!g1354) & (!g1355) & (g1357)) + ((sk[108]) & (g940) & (!g1353) & (g1354) & (!g1355) & (g1357)) + ((sk[108]) & (g940) & (g1353) & (!g1354) & (!g1355) & (g1357)));
	assign g1359 = (((!sk[109]) & (!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[109]) & (!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[109]) & (!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g112)) + ((!sk[109]) & (!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g112)) + ((!sk[109]) & (!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((!sk[109]) & (!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g112)) + ((!sk[109]) & (!i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g112)) + ((!sk[109]) & (!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g112)) + ((!sk[109]) & (!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[109]) & (!i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[109]) & (!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g112)) + ((!sk[109]) & (i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[109]) & (i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[109]) & (i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g112)) + ((!sk[109]) & (i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (!g112)) + ((!sk[109]) & (i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((!sk[109]) & (i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g112)) + ((!sk[109]) & (i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g112)) + ((!sk[109]) & (i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g112)) + ((!sk[109]) & (i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!sk[109]) & (i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!sk[109]) & (i_15_) & (i_12_) & (i_13_) & (i_14_) & (g112)) + ((sk[109]) & (!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g112)) + ((sk[109]) & (!i_15_) & (!i_12_) & (i_13_) & (!i_14_) & (g112)) + ((sk[109]) & (!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g112)) + ((sk[109]) & (!i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((sk[109]) & (!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112)) + ((sk[109]) & (!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g112)) + ((sk[109]) & (i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((sk[109]) & (i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g112)) + ((sk[109]) & (i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g112)) + ((sk[109]) & (i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((sk[109]) & (i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g112)) + ((sk[109]) & (i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g112)));
	assign g1360 = (((!i_15_) & (!sk[110]) & (!i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!i_15_) & (!sk[110]) & (!i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!i_15_) & (!sk[110]) & (!i_12_) & (i_13_) & (i_14_) & (g112)) + ((!i_15_) & (!sk[110]) & (i_12_) & (!i_13_) & (!i_14_) & (!g112)) + ((!i_15_) & (!sk[110]) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((!i_15_) & (!sk[110]) & (i_12_) & (!i_13_) & (i_14_) & (!g112)) + ((!i_15_) & (!sk[110]) & (i_12_) & (!i_13_) & (i_14_) & (g112)) + ((!i_15_) & (!sk[110]) & (i_12_) & (i_13_) & (!i_14_) & (!g112)) + ((!i_15_) & (!sk[110]) & (i_12_) & (i_13_) & (!i_14_) & (g112)) + ((!i_15_) & (!sk[110]) & (i_12_) & (i_13_) & (i_14_) & (!g112)) + ((!i_15_) & (!sk[110]) & (i_12_) & (i_13_) & (i_14_) & (g112)) + ((!i_15_) & (sk[110]) & (!i_12_) & (!i_13_) & (i_14_) & (g112)) + ((!i_15_) & (sk[110]) & (!i_12_) & (i_13_) & (i_14_) & (g112)) + ((!i_15_) & (sk[110]) & (i_12_) & (i_13_) & (!i_14_) & (g112)) + ((i_15_) & (!sk[110]) & (!i_12_) & (i_13_) & (!i_14_) & (g112)) + ((i_15_) & (!sk[110]) & (!i_12_) & (i_13_) & (i_14_) & (!g112)) + ((i_15_) & (!sk[110]) & (!i_12_) & (i_13_) & (i_14_) & (g112)) + ((i_15_) & (!sk[110]) & (i_12_) & (!i_13_) & (!i_14_) & (!g112)) + ((i_15_) & (!sk[110]) & (i_12_) & (!i_13_) & (!i_14_) & (g112)) + ((i_15_) & (!sk[110]) & (i_12_) & (!i_13_) & (i_14_) & (!g112)) + ((i_15_) & (!sk[110]) & (i_12_) & (!i_13_) & (i_14_) & (g112)) + ((i_15_) & (!sk[110]) & (i_12_) & (i_13_) & (!i_14_) & (!g112)) + ((i_15_) & (!sk[110]) & (i_12_) & (i_13_) & (!i_14_) & (g112)) + ((i_15_) & (!sk[110]) & (i_12_) & (i_13_) & (i_14_) & (!g112)) + ((i_15_) & (!sk[110]) & (i_12_) & (i_13_) & (i_14_) & (g112)) + ((i_15_) & (sk[110]) & (!i_12_) & (!i_13_) & (i_14_) & (g112)) + ((i_15_) & (sk[110]) & (i_12_) & (i_13_) & (!i_14_) & (g112)));
	assign g1361 = (((!i_8_) & (!g107) & (g735) & (!sk[111]) & (!g1267) & (g1360)) + ((!i_8_) & (!g107) & (g735) & (!sk[111]) & (g1267) & (!g1360)) + ((!i_8_) & (!g107) & (g735) & (!sk[111]) & (g1267) & (g1360)) + ((!i_8_) & (g107) & (!g735) & (!sk[111]) & (!g1267) & (!g1360)) + ((!i_8_) & (g107) & (!g735) & (!sk[111]) & (!g1267) & (g1360)) + ((!i_8_) & (g107) & (!g735) & (!sk[111]) & (g1267) & (!g1360)) + ((!i_8_) & (g107) & (!g735) & (!sk[111]) & (g1267) & (g1360)) + ((!i_8_) & (g107) & (g735) & (!sk[111]) & (!g1267) & (!g1360)) + ((!i_8_) & (g107) & (g735) & (!sk[111]) & (!g1267) & (g1360)) + ((!i_8_) & (g107) & (g735) & (!sk[111]) & (g1267) & (!g1360)) + ((!i_8_) & (g107) & (g735) & (!sk[111]) & (g1267) & (g1360)) + ((i_8_) & (!g107) & (!g735) & (sk[111]) & (!g1267) & (!g1360)) + ((i_8_) & (!g107) & (g735) & (!sk[111]) & (!g1267) & (g1360)) + ((i_8_) & (!g107) & (g735) & (!sk[111]) & (g1267) & (!g1360)) + ((i_8_) & (!g107) & (g735) & (!sk[111]) & (g1267) & (g1360)) + ((i_8_) & (g107) & (!g735) & (!sk[111]) & (!g1267) & (!g1360)) + ((i_8_) & (g107) & (!g735) & (!sk[111]) & (!g1267) & (g1360)) + ((i_8_) & (g107) & (!g735) & (!sk[111]) & (g1267) & (!g1360)) + ((i_8_) & (g107) & (!g735) & (!sk[111]) & (g1267) & (g1360)) + ((i_8_) & (g107) & (!g735) & (sk[111]) & (!g1267) & (!g1360)) + ((i_8_) & (g107) & (g735) & (!sk[111]) & (!g1267) & (!g1360)) + ((i_8_) & (g107) & (g735) & (!sk[111]) & (!g1267) & (g1360)) + ((i_8_) & (g107) & (g735) & (!sk[111]) & (g1267) & (!g1360)) + ((i_8_) & (g107) & (g735) & (!sk[111]) & (g1267) & (g1360)) + ((i_8_) & (g107) & (g735) & (sk[111]) & (!g1267) & (!g1360)));
	assign g1362 = (((!sk[112]) & (!i_8_) & (!g165) & (g487) & (!g1359) & (g1361)) + ((!sk[112]) & (!i_8_) & (!g165) & (g487) & (g1359) & (!g1361)) + ((!sk[112]) & (!i_8_) & (!g165) & (g487) & (g1359) & (g1361)) + ((!sk[112]) & (!i_8_) & (g165) & (!g487) & (!g1359) & (!g1361)) + ((!sk[112]) & (!i_8_) & (g165) & (!g487) & (!g1359) & (g1361)) + ((!sk[112]) & (!i_8_) & (g165) & (!g487) & (g1359) & (!g1361)) + ((!sk[112]) & (!i_8_) & (g165) & (!g487) & (g1359) & (g1361)) + ((!sk[112]) & (!i_8_) & (g165) & (g487) & (!g1359) & (!g1361)) + ((!sk[112]) & (!i_8_) & (g165) & (g487) & (!g1359) & (g1361)) + ((!sk[112]) & (!i_8_) & (g165) & (g487) & (g1359) & (!g1361)) + ((!sk[112]) & (!i_8_) & (g165) & (g487) & (g1359) & (g1361)) + ((!sk[112]) & (i_8_) & (!g165) & (g487) & (!g1359) & (g1361)) + ((!sk[112]) & (i_8_) & (!g165) & (g487) & (g1359) & (!g1361)) + ((!sk[112]) & (i_8_) & (!g165) & (g487) & (g1359) & (g1361)) + ((!sk[112]) & (i_8_) & (g165) & (!g487) & (!g1359) & (!g1361)) + ((!sk[112]) & (i_8_) & (g165) & (!g487) & (!g1359) & (g1361)) + ((!sk[112]) & (i_8_) & (g165) & (!g487) & (g1359) & (!g1361)) + ((!sk[112]) & (i_8_) & (g165) & (!g487) & (g1359) & (g1361)) + ((!sk[112]) & (i_8_) & (g165) & (g487) & (!g1359) & (!g1361)) + ((!sk[112]) & (i_8_) & (g165) & (g487) & (!g1359) & (g1361)) + ((!sk[112]) & (i_8_) & (g165) & (g487) & (g1359) & (!g1361)) + ((!sk[112]) & (i_8_) & (g165) & (g487) & (g1359) & (g1361)) + ((sk[112]) & (!i_8_) & (g165) & (!g487) & (g1359) & (!g1361)) + ((sk[112]) & (!i_8_) & (g165) & (g487) & (!g1359) & (!g1361)) + ((sk[112]) & (!i_8_) & (g165) & (g487) & (g1359) & (!g1361)) + ((sk[112]) & (i_8_) & (g165) & (!g487) & (!g1359) & (!g1361)) + ((sk[112]) & (i_8_) & (g165) & (!g487) & (g1359) & (!g1361)) + ((sk[112]) & (i_8_) & (g165) & (g487) & (!g1359) & (!g1361)) + ((sk[112]) & (i_8_) & (g165) & (g487) & (g1359) & (!g1361)));
	assign g1363 = (((!sk[113]) & (!g135) & (!g122) & (g185) & (!g562)) + ((!sk[113]) & (!g135) & (!g122) & (g185) & (g562)) + ((!sk[113]) & (!g135) & (g122) & (g185) & (!g562)) + ((!sk[113]) & (!g135) & (g122) & (g185) & (g562)) + ((!sk[113]) & (g135) & (!g122) & (g185) & (!g562)) + ((!sk[113]) & (g135) & (!g122) & (g185) & (g562)) + ((!sk[113]) & (g135) & (g122) & (g185) & (!g562)) + ((!sk[113]) & (g135) & (g122) & (g185) & (g562)) + ((sk[113]) & (!g135) & (!g122) & (g185) & (!g562)) + ((sk[113]) & (!g135) & (!g122) & (g185) & (g562)) + ((sk[113]) & (!g135) & (g122) & (!g185) & (g562)) + ((sk[113]) & (!g135) & (g122) & (g185) & (!g562)) + ((sk[113]) & (!g135) & (g122) & (g185) & (g562)) + ((sk[113]) & (g135) & (g122) & (!g185) & (g562)) + ((sk[113]) & (g135) & (g122) & (g185) & (g562)));
	assign g1364 = (((!g165) & (!g122) & (!g114) & (!g286) & (!g557) & (!g983)) + ((!g165) & (!g122) & (!g114) & (!g286) & (!g557) & (g983)) + ((!g165) & (!g122) & (!g114) & (!g286) & (g557) & (!g983)) + ((!g165) & (!g122) & (!g114) & (!g286) & (g557) & (g983)) + ((!g165) & (!g122) & (!g114) & (g286) & (!g557) & (!g983)) + ((!g165) & (!g122) & (!g114) & (g286) & (!g557) & (g983)) + ((!g165) & (!g122) & (!g114) & (g286) & (g557) & (!g983)) + ((!g165) & (!g122) & (!g114) & (g286) & (g557) & (g983)) + ((!g165) & (!g122) & (g114) & (!g286) & (!g557) & (!g983)) + ((!g165) & (!g122) & (g114) & (!g286) & (!g557) & (g983)) + ((!g165) & (!g122) & (g114) & (!g286) & (g557) & (!g983)) + ((!g165) & (!g122) & (g114) & (!g286) & (g557) & (g983)) + ((!g165) & (!g122) & (g114) & (g286) & (!g557) & (!g983)) + ((!g165) & (!g122) & (g114) & (g286) & (!g557) & (g983)) + ((!g165) & (!g122) & (g114) & (g286) & (g557) & (!g983)) + ((!g165) & (!g122) & (g114) & (g286) & (g557) & (g983)) + ((!g165) & (g122) & (g114) & (!g286) & (!g557) & (!g983)) + ((!g165) & (g122) & (g114) & (!g286) & (!g557) & (g983)) + ((g165) & (!g122) & (!g114) & (!g286) & (!g557) & (!g983)) + ((g165) & (!g122) & (!g114) & (!g286) & (g557) & (!g983)) + ((g165) & (!g122) & (!g114) & (g286) & (!g557) & (!g983)) + ((g165) & (!g122) & (!g114) & (g286) & (g557) & (!g983)) + ((g165) & (!g122) & (g114) & (!g286) & (!g557) & (!g983)) + ((g165) & (!g122) & (g114) & (!g286) & (g557) & (!g983)) + ((g165) & (!g122) & (g114) & (g286) & (!g557) & (!g983)) + ((g165) & (!g122) & (g114) & (g286) & (g557) & (!g983)) + ((g165) & (g122) & (g114) & (!g286) & (!g557) & (!g983)));
	assign g1365 = (((!g122) & (!g197) & (!g200) & (!g715) & (!g1363) & (g1364)) + ((!g122) & (!g197) & (g200) & (!g715) & (!g1363) & (g1364)) + ((!g122) & (g197) & (!g200) & (!g715) & (!g1363) & (g1364)) + ((!g122) & (g197) & (g200) & (!g715) & (!g1363) & (g1364)) + ((g122) & (!g197) & (!g200) & (!g715) & (!g1363) & (g1364)));
	assign g1366 = (((!g1025) & (!sk[116]) & (!g1031) & (g1362) & (!g1365)) + ((!g1025) & (!sk[116]) & (!g1031) & (g1362) & (g1365)) + ((!g1025) & (!sk[116]) & (g1031) & (g1362) & (!g1365)) + ((!g1025) & (!sk[116]) & (g1031) & (g1362) & (g1365)) + ((g1025) & (!sk[116]) & (!g1031) & (g1362) & (!g1365)) + ((g1025) & (!sk[116]) & (!g1031) & (g1362) & (g1365)) + ((g1025) & (!sk[116]) & (g1031) & (g1362) & (!g1365)) + ((g1025) & (!sk[116]) & (g1031) & (g1362) & (g1365)) + ((g1025) & (sk[116]) & (g1031) & (!g1362) & (g1365)));
	assign g1367 = (((!g1184) & (!g527) & (g1009) & (!g1185) & (g1187) & (g1188)));
	assign g1368 = (((g987) & (g1099) & (g1352) & (g1358) & (g1366) & (g1367)));
	assign g1369 = (((!g165) & (!sk[119]) & (!g122) & (g343) & (!g626) & (g945)) + ((!g165) & (!sk[119]) & (!g122) & (g343) & (g626) & (!g945)) + ((!g165) & (!sk[119]) & (!g122) & (g343) & (g626) & (g945)) + ((!g165) & (!sk[119]) & (g122) & (!g343) & (!g626) & (!g945)) + ((!g165) & (!sk[119]) & (g122) & (!g343) & (!g626) & (g945)) + ((!g165) & (!sk[119]) & (g122) & (!g343) & (g626) & (!g945)) + ((!g165) & (!sk[119]) & (g122) & (!g343) & (g626) & (g945)) + ((!g165) & (!sk[119]) & (g122) & (g343) & (!g626) & (!g945)) + ((!g165) & (!sk[119]) & (g122) & (g343) & (!g626) & (g945)) + ((!g165) & (!sk[119]) & (g122) & (g343) & (g626) & (!g945)) + ((!g165) & (!sk[119]) & (g122) & (g343) & (g626) & (g945)) + ((!g165) & (sk[119]) & (!g122) & (!g343) & (!g626) & (!g945)) + ((!g165) & (sk[119]) & (!g122) & (!g343) & (!g626) & (g945)) + ((!g165) & (sk[119]) & (!g122) & (!g343) & (g626) & (!g945)) + ((!g165) & (sk[119]) & (!g122) & (!g343) & (g626) & (g945)) + ((!g165) & (sk[119]) & (!g122) & (g343) & (!g626) & (!g945)) + ((!g165) & (sk[119]) & (!g122) & (g343) & (!g626) & (g945)) + ((!g165) & (sk[119]) & (!g122) & (g343) & (g626) & (!g945)) + ((!g165) & (sk[119]) & (!g122) & (g343) & (g626) & (g945)) + ((!g165) & (sk[119]) & (g122) & (g343) & (!g626) & (!g945)) + ((!g165) & (sk[119]) & (g122) & (g343) & (!g626) & (g945)) + ((g165) & (!sk[119]) & (!g122) & (g343) & (!g626) & (g945)) + ((g165) & (!sk[119]) & (!g122) & (g343) & (g626) & (!g945)) + ((g165) & (!sk[119]) & (!g122) & (g343) & (g626) & (g945)) + ((g165) & (!sk[119]) & (g122) & (!g343) & (!g626) & (!g945)) + ((g165) & (!sk[119]) & (g122) & (!g343) & (!g626) & (g945)) + ((g165) & (!sk[119]) & (g122) & (!g343) & (g626) & (!g945)) + ((g165) & (!sk[119]) & (g122) & (!g343) & (g626) & (g945)) + ((g165) & (!sk[119]) & (g122) & (g343) & (!g626) & (!g945)) + ((g165) & (!sk[119]) & (g122) & (g343) & (!g626) & (g945)) + ((g165) & (!sk[119]) & (g122) & (g343) & (g626) & (!g945)) + ((g165) & (!sk[119]) & (g122) & (g343) & (g626) & (g945)) + ((g165) & (sk[119]) & (!g122) & (!g343) & (!g626) & (g945)) + ((g165) & (sk[119]) & (!g122) & (!g343) & (g626) & (g945)) + ((g165) & (sk[119]) & (!g122) & (g343) & (!g626) & (g945)) + ((g165) & (sk[119]) & (!g122) & (g343) & (g626) & (g945)) + ((g165) & (sk[119]) & (g122) & (g343) & (!g626) & (g945)));
	assign g1370 = (((!g135) & (!sk[120]) & (!g605) & (g761) & (!g1369)) + ((!g135) & (!sk[120]) & (!g605) & (g761) & (g1369)) + ((!g135) & (!sk[120]) & (g605) & (g761) & (!g1369)) + ((!g135) & (!sk[120]) & (g605) & (g761) & (g1369)) + ((!g135) & (sk[120]) & (!g605) & (g761) & (g1369)) + ((g135) & (!sk[120]) & (!g605) & (g761) & (!g1369)) + ((g135) & (!sk[120]) & (!g605) & (g761) & (g1369)) + ((g135) & (!sk[120]) & (g605) & (g761) & (!g1369)) + ((g135) & (!sk[120]) & (g605) & (g761) & (g1369)) + ((g135) & (sk[120]) & (!g605) & (!g761) & (g1369)) + ((g135) & (sk[120]) & (!g605) & (g761) & (g1369)) + ((g135) & (sk[120]) & (g605) & (!g761) & (g1369)) + ((g135) & (sk[120]) & (g605) & (g761) & (g1369)));
	assign g1371 = (((!g159) & (!g253) & (!sk[121]) & (g333) & (!g865)) + ((!g159) & (!g253) & (!sk[121]) & (g333) & (g865)) + ((!g159) & (!g253) & (sk[121]) & (!g333) & (!g865)) + ((!g159) & (g253) & (!sk[121]) & (g333) & (!g865)) + ((!g159) & (g253) & (!sk[121]) & (g333) & (g865)) + ((!g159) & (g253) & (sk[121]) & (!g333) & (!g865)) + ((g159) & (!g253) & (!sk[121]) & (g333) & (!g865)) + ((g159) & (!g253) & (!sk[121]) & (g333) & (g865)) + ((g159) & (!g253) & (sk[121]) & (!g333) & (!g865)) + ((g159) & (!g253) & (sk[121]) & (!g333) & (g865)) + ((g159) & (g253) & (!sk[121]) & (g333) & (!g865)) + ((g159) & (g253) & (!sk[121]) & (g333) & (g865)) + ((g159) & (g253) & (sk[121]) & (!g333) & (!g865)) + ((g159) & (g253) & (sk[121]) & (!g333) & (g865)) + ((g159) & (g253) & (sk[121]) & (g333) & (!g865)) + ((g159) & (g253) & (sk[121]) & (g333) & (g865)));
	assign g1372 = (((!g20) & (!g24) & (g74) & (!sk[122]) & (!g460)) + ((!g20) & (!g24) & (g74) & (!sk[122]) & (g460)) + ((!g20) & (g24) & (g74) & (!sk[122]) & (!g460)) + ((!g20) & (g24) & (g74) & (!sk[122]) & (g460)) + ((g20) & (!g24) & (g74) & (!sk[122]) & (!g460)) + ((g20) & (!g24) & (g74) & (!sk[122]) & (g460)) + ((g20) & (!g24) & (g74) & (sk[122]) & (!g460)) + ((g20) & (!g24) & (g74) & (sk[122]) & (g460)) + ((g20) & (g24) & (g74) & (!sk[122]) & (!g460)) + ((g20) & (g24) & (g74) & (!sk[122]) & (g460)) + ((g20) & (g24) & (g74) & (sk[122]) & (!g460)));
	assign g1373 = (((!i_12_) & (!i_13_) & (!i_14_) & (sk[123]) & (!g22) & (g102)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[123]) & (!g22) & (g102)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[123]) & (g22) & (!g102)) + ((!i_12_) & (!i_13_) & (i_14_) & (!sk[123]) & (g22) & (g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[123]) & (!g22) & (!g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[123]) & (!g22) & (g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[123]) & (g22) & (!g102)) + ((!i_12_) & (i_13_) & (!i_14_) & (!sk[123]) & (g22) & (g102)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[123]) & (!g22) & (!g102)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[123]) & (!g22) & (g102)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[123]) & (g22) & (!g102)) + ((!i_12_) & (i_13_) & (i_14_) & (!sk[123]) & (g22) & (g102)) + ((!i_12_) & (i_13_) & (i_14_) & (sk[123]) & (!g22) & (g102)) + ((i_12_) & (!i_13_) & (!i_14_) & (sk[123]) & (!g22) & (g102)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[123]) & (!g22) & (g102)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[123]) & (g22) & (!g102)) + ((i_12_) & (!i_13_) & (i_14_) & (!sk[123]) & (g22) & (g102)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[123]) & (!g22) & (!g102)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[123]) & (!g22) & (g102)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[123]) & (g22) & (!g102)) + ((i_12_) & (i_13_) & (!i_14_) & (!sk[123]) & (g22) & (g102)) + ((i_12_) & (i_13_) & (!i_14_) & (sk[123]) & (!g22) & (g102)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[123]) & (!g22) & (!g102)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[123]) & (!g22) & (g102)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[123]) & (g22) & (!g102)) + ((i_12_) & (i_13_) & (i_14_) & (!sk[123]) & (g22) & (g102)));
	assign g1374 = (((!sk[124]) & (!g257) & (!g313) & (g278) & (!g333)) + ((!sk[124]) & (!g257) & (!g313) & (g278) & (g333)) + ((!sk[124]) & (!g257) & (g313) & (g278) & (!g333)) + ((!sk[124]) & (!g257) & (g313) & (g278) & (g333)) + ((!sk[124]) & (g257) & (!g313) & (g278) & (!g333)) + ((!sk[124]) & (g257) & (!g313) & (g278) & (g333)) + ((!sk[124]) & (g257) & (g313) & (g278) & (!g333)) + ((!sk[124]) & (g257) & (g313) & (g278) & (g333)) + ((sk[124]) & (!g257) & (!g313) & (!g278) & (!g333)) + ((sk[124]) & (!g257) & (!g313) & (!g278) & (g333)) + ((sk[124]) & (!g257) & (!g313) & (g278) & (!g333)) + ((sk[124]) & (!g257) & (!g313) & (g278) & (g333)) + ((sk[124]) & (!g257) & (g313) & (!g278) & (!g333)) + ((sk[124]) & (g257) & (!g313) & (!g278) & (!g333)) + ((sk[124]) & (g257) & (!g313) & (!g278) & (g333)) + ((sk[124]) & (g257) & (g313) & (!g278) & (!g333)));
	assign g1375 = (((!g122) & (!g1314) & (g1371) & (!g1372) & (!g1373) & (g1374)) + ((!g122) & (g1314) & (g1371) & (!g1372) & (!g1373) & (g1374)) + ((g122) & (g1314) & (g1371) & (!g1372) & (!g1373) & (g1374)));
	assign g1376 = (((!g125) & (!g159) & (!sk[126]) & (g521) & (!g642)) + ((!g125) & (!g159) & (!sk[126]) & (g521) & (g642)) + ((!g125) & (!g159) & (sk[126]) & (g521) & (!g642)) + ((!g125) & (!g159) & (sk[126]) & (g521) & (g642)) + ((!g125) & (g159) & (!sk[126]) & (g521) & (!g642)) + ((!g125) & (g159) & (!sk[126]) & (g521) & (g642)) + ((g125) & (!g159) & (!sk[126]) & (g521) & (!g642)) + ((g125) & (!g159) & (!sk[126]) & (g521) & (g642)) + ((g125) & (!g159) & (sk[126]) & (!g521) & (g642)) + ((g125) & (!g159) & (sk[126]) & (g521) & (!g642)) + ((g125) & (!g159) & (sk[126]) & (g521) & (g642)) + ((g125) & (g159) & (!sk[126]) & (g521) & (!g642)) + ((g125) & (g159) & (!sk[126]) & (g521) & (g642)) + ((g125) & (g159) & (sk[126]) & (!g521) & (g642)) + ((g125) & (g159) & (sk[126]) & (g521) & (g642)));
	assign g1377 = (((!g23) & (!g157) & (g130) & (!g175) & (!g449) & (!g1376)) + ((!g23) & (!g157) & (g130) & (!g175) & (g449) & (!g1376)) + ((!g23) & (!g157) & (g130) & (g175) & (!g449) & (!g1376)) + ((!g23) & (!g157) & (g130) & (g175) & (g449) & (!g1376)) + ((!g23) & (g157) & (g130) & (!g175) & (g449) & (!g1376)) + ((!g23) & (g157) & (g130) & (g175) & (g449) & (!g1376)) + ((g23) & (!g157) & (!g130) & (!g175) & (!g449) & (!g1376)) + ((g23) & (!g157) & (!g130) & (!g175) & (g449) & (!g1376)) + ((g23) & (!g157) & (g130) & (!g175) & (!g449) & (!g1376)) + ((g23) & (!g157) & (g130) & (!g175) & (g449) & (!g1376)) + ((g23) & (!g157) & (g130) & (g175) & (!g449) & (!g1376)) + ((g23) & (!g157) & (g130) & (g175) & (g449) & (!g1376)) + ((g23) & (g157) & (!g130) & (!g175) & (g449) & (!g1376)) + ((g23) & (g157) & (g130) & (!g175) & (g449) & (!g1376)) + ((g23) & (g157) & (g130) & (g175) & (g449) & (!g1376)));
	assign g1378 = (((!g165) & (!g257) & (!g738) & (!g777) & (sk[0]) & (g1377)) + ((!g165) & (!g257) & (!g738) & (g777) & (sk[0]) & (g1377)) + ((!g165) & (!g257) & (g738) & (!g777) & (!sk[0]) & (g1377)) + ((!g165) & (!g257) & (g738) & (!g777) & (sk[0]) & (g1377)) + ((!g165) & (!g257) & (g738) & (g777) & (!sk[0]) & (!g1377)) + ((!g165) & (!g257) & (g738) & (g777) & (!sk[0]) & (g1377)) + ((!g165) & (!g257) & (g738) & (g777) & (sk[0]) & (g1377)) + ((!g165) & (g257) & (!g738) & (!g777) & (!sk[0]) & (!g1377)) + ((!g165) & (g257) & (!g738) & (!g777) & (!sk[0]) & (g1377)) + ((!g165) & (g257) & (!g738) & (!g777) & (sk[0]) & (g1377)) + ((!g165) & (g257) & (!g738) & (g777) & (!sk[0]) & (!g1377)) + ((!g165) & (g257) & (!g738) & (g777) & (!sk[0]) & (g1377)) + ((!g165) & (g257) & (!g738) & (g777) & (sk[0]) & (g1377)) + ((!g165) & (g257) & (g738) & (!g777) & (!sk[0]) & (!g1377)) + ((!g165) & (g257) & (g738) & (!g777) & (!sk[0]) & (g1377)) + ((!g165) & (g257) & (g738) & (g777) & (!sk[0]) & (!g1377)) + ((!g165) & (g257) & (g738) & (g777) & (!sk[0]) & (g1377)) + ((g165) & (!g257) & (!g738) & (!g777) & (sk[0]) & (g1377)) + ((g165) & (!g257) & (g738) & (!g777) & (!sk[0]) & (g1377)) + ((g165) & (!g257) & (g738) & (!g777) & (sk[0]) & (g1377)) + ((g165) & (!g257) & (g738) & (g777) & (!sk[0]) & (!g1377)) + ((g165) & (!g257) & (g738) & (g777) & (!sk[0]) & (g1377)) + ((g165) & (g257) & (!g738) & (!g777) & (!sk[0]) & (!g1377)) + ((g165) & (g257) & (!g738) & (!g777) & (!sk[0]) & (g1377)) + ((g165) & (g257) & (!g738) & (!g777) & (sk[0]) & (g1377)) + ((g165) & (g257) & (!g738) & (g777) & (!sk[0]) & (!g1377)) + ((g165) & (g257) & (!g738) & (g777) & (!sk[0]) & (g1377)) + ((g165) & (g257) & (g738) & (!g777) & (!sk[0]) & (!g1377)) + ((g165) & (g257) & (g738) & (!g777) & (!sk[0]) & (g1377)) + ((g165) & (g257) & (g738) & (g777) & (!sk[0]) & (!g1377)) + ((g165) & (g257) & (g738) & (g777) & (!sk[0]) & (g1377)));
	assign g1379 = (((!g425) & (!g408) & (g945) & (!sk[1]) & (!g1248) & (g1111)) + ((!g425) & (!g408) & (g945) & (!sk[1]) & (g1248) & (!g1111)) + ((!g425) & (!g408) & (g945) & (!sk[1]) & (g1248) & (g1111)) + ((!g425) & (!g408) & (g945) & (sk[1]) & (!g1248) & (!g1111)) + ((!g425) & (g408) & (!g945) & (!sk[1]) & (!g1248) & (!g1111)) + ((!g425) & (g408) & (!g945) & (!sk[1]) & (!g1248) & (g1111)) + ((!g425) & (g408) & (!g945) & (!sk[1]) & (g1248) & (!g1111)) + ((!g425) & (g408) & (!g945) & (!sk[1]) & (g1248) & (g1111)) + ((!g425) & (g408) & (g945) & (!sk[1]) & (!g1248) & (!g1111)) + ((!g425) & (g408) & (g945) & (!sk[1]) & (!g1248) & (g1111)) + ((!g425) & (g408) & (g945) & (!sk[1]) & (g1248) & (!g1111)) + ((!g425) & (g408) & (g945) & (!sk[1]) & (g1248) & (g1111)) + ((!g425) & (g408) & (g945) & (sk[1]) & (!g1248) & (!g1111)) + ((!g425) & (g408) & (g945) & (sk[1]) & (g1248) & (!g1111)) + ((g425) & (!g408) & (!g945) & (sk[1]) & (!g1248) & (!g1111)) + ((g425) & (!g408) & (g945) & (!sk[1]) & (!g1248) & (g1111)) + ((g425) & (!g408) & (g945) & (!sk[1]) & (g1248) & (!g1111)) + ((g425) & (!g408) & (g945) & (!sk[1]) & (g1248) & (g1111)) + ((g425) & (!g408) & (g945) & (sk[1]) & (!g1248) & (!g1111)) + ((g425) & (g408) & (!g945) & (!sk[1]) & (!g1248) & (!g1111)) + ((g425) & (g408) & (!g945) & (!sk[1]) & (!g1248) & (g1111)) + ((g425) & (g408) & (!g945) & (!sk[1]) & (g1248) & (!g1111)) + ((g425) & (g408) & (!g945) & (!sk[1]) & (g1248) & (g1111)) + ((g425) & (g408) & (!g945) & (sk[1]) & (!g1248) & (!g1111)) + ((g425) & (g408) & (!g945) & (sk[1]) & (g1248) & (!g1111)) + ((g425) & (g408) & (g945) & (!sk[1]) & (!g1248) & (!g1111)) + ((g425) & (g408) & (g945) & (!sk[1]) & (!g1248) & (g1111)) + ((g425) & (g408) & (g945) & (!sk[1]) & (g1248) & (!g1111)) + ((g425) & (g408) & (g945) & (!sk[1]) & (g1248) & (g1111)) + ((g425) & (g408) & (g945) & (sk[1]) & (!g1248) & (!g1111)) + ((g425) & (g408) & (g945) & (sk[1]) & (g1248) & (!g1111)));
	assign g1380 = (((!g74) & (!g521) & (!sk[2]) & (g1041) & (!g388)) + ((!g74) & (!g521) & (!sk[2]) & (g1041) & (g388)) + ((!g74) & (!g521) & (sk[2]) & (!g1041) & (!g388)) + ((!g74) & (!g521) & (sk[2]) & (g1041) & (!g388)) + ((!g74) & (g521) & (!sk[2]) & (g1041) & (!g388)) + ((!g74) & (g521) & (!sk[2]) & (g1041) & (g388)) + ((!g74) & (g521) & (sk[2]) & (!g1041) & (!g388)) + ((!g74) & (g521) & (sk[2]) & (g1041) & (!g388)) + ((g74) & (!g521) & (!sk[2]) & (g1041) & (!g388)) + ((g74) & (!g521) & (!sk[2]) & (g1041) & (g388)) + ((g74) & (!g521) & (sk[2]) & (g1041) & (!g388)) + ((g74) & (g521) & (!sk[2]) & (g1041) & (!g388)) + ((g74) & (g521) & (!sk[2]) & (g1041) & (g388)));
	assign g1381 = (((!sk[3]) & (!g1370) & (!g1375) & (g1378) & (!g1379) & (g1380)) + ((!sk[3]) & (!g1370) & (!g1375) & (g1378) & (g1379) & (!g1380)) + ((!sk[3]) & (!g1370) & (!g1375) & (g1378) & (g1379) & (g1380)) + ((!sk[3]) & (!g1370) & (g1375) & (!g1378) & (!g1379) & (!g1380)) + ((!sk[3]) & (!g1370) & (g1375) & (!g1378) & (!g1379) & (g1380)) + ((!sk[3]) & (!g1370) & (g1375) & (!g1378) & (g1379) & (!g1380)) + ((!sk[3]) & (!g1370) & (g1375) & (!g1378) & (g1379) & (g1380)) + ((!sk[3]) & (!g1370) & (g1375) & (g1378) & (!g1379) & (!g1380)) + ((!sk[3]) & (!g1370) & (g1375) & (g1378) & (!g1379) & (g1380)) + ((!sk[3]) & (!g1370) & (g1375) & (g1378) & (g1379) & (!g1380)) + ((!sk[3]) & (!g1370) & (g1375) & (g1378) & (g1379) & (g1380)) + ((!sk[3]) & (g1370) & (!g1375) & (g1378) & (!g1379) & (g1380)) + ((!sk[3]) & (g1370) & (!g1375) & (g1378) & (g1379) & (!g1380)) + ((!sk[3]) & (g1370) & (!g1375) & (g1378) & (g1379) & (g1380)) + ((!sk[3]) & (g1370) & (g1375) & (!g1378) & (!g1379) & (!g1380)) + ((!sk[3]) & (g1370) & (g1375) & (!g1378) & (!g1379) & (g1380)) + ((!sk[3]) & (g1370) & (g1375) & (!g1378) & (g1379) & (!g1380)) + ((!sk[3]) & (g1370) & (g1375) & (!g1378) & (g1379) & (g1380)) + ((!sk[3]) & (g1370) & (g1375) & (g1378) & (!g1379) & (!g1380)) + ((!sk[3]) & (g1370) & (g1375) & (g1378) & (!g1379) & (g1380)) + ((!sk[3]) & (g1370) & (g1375) & (g1378) & (g1379) & (!g1380)) + ((!sk[3]) & (g1370) & (g1375) & (g1378) & (g1379) & (g1380)) + ((sk[3]) & (g1370) & (g1375) & (g1378) & (g1379) & (g1380)));
	assign g1382 = (((!i_8_) & (!i_6_) & (g120) & (!sk[4]) & (!g761)) + ((!i_8_) & (!i_6_) & (g120) & (!sk[4]) & (g761)) + ((!i_8_) & (!i_6_) & (g120) & (sk[4]) & (!g761)) + ((!i_8_) & (i_6_) & (g120) & (!sk[4]) & (!g761)) + ((!i_8_) & (i_6_) & (g120) & (!sk[4]) & (g761)) + ((i_8_) & (!i_6_) & (g120) & (!sk[4]) & (!g761)) + ((i_8_) & (!i_6_) & (g120) & (!sk[4]) & (g761)) + ((i_8_) & (i_6_) & (g120) & (!sk[4]) & (!g761)) + ((i_8_) & (i_6_) & (g120) & (!sk[4]) & (g761)));
	assign g1383 = (((!g21) & (!g23) & (!sk[5]) & (g74) & (!g495) & (g1382)) + ((!g21) & (!g23) & (!sk[5]) & (g74) & (g495) & (!g1382)) + ((!g21) & (!g23) & (!sk[5]) & (g74) & (g495) & (g1382)) + ((!g21) & (!g23) & (sk[5]) & (!g74) & (!g495) & (!g1382)) + ((!g21) & (!g23) & (sk[5]) & (!g74) & (g495) & (!g1382)) + ((!g21) & (g23) & (!sk[5]) & (!g74) & (!g495) & (!g1382)) + ((!g21) & (g23) & (!sk[5]) & (!g74) & (!g495) & (g1382)) + ((!g21) & (g23) & (!sk[5]) & (!g74) & (g495) & (!g1382)) + ((!g21) & (g23) & (!sk[5]) & (!g74) & (g495) & (g1382)) + ((!g21) & (g23) & (!sk[5]) & (g74) & (!g495) & (!g1382)) + ((!g21) & (g23) & (!sk[5]) & (g74) & (!g495) & (g1382)) + ((!g21) & (g23) & (!sk[5]) & (g74) & (g495) & (!g1382)) + ((!g21) & (g23) & (!sk[5]) & (g74) & (g495) & (g1382)) + ((!g21) & (g23) & (sk[5]) & (!g74) & (!g495) & (!g1382)) + ((!g21) & (g23) & (sk[5]) & (!g74) & (g495) & (!g1382)) + ((!g21) & (g23) & (sk[5]) & (g74) & (!g495) & (!g1382)) + ((g21) & (!g23) & (!sk[5]) & (g74) & (!g495) & (g1382)) + ((g21) & (!g23) & (!sk[5]) & (g74) & (g495) & (!g1382)) + ((g21) & (!g23) & (!sk[5]) & (g74) & (g495) & (g1382)) + ((g21) & (!g23) & (sk[5]) & (!g74) & (!g495) & (!g1382)) + ((g21) & (!g23) & (sk[5]) & (!g74) & (g495) & (!g1382)) + ((g21) & (g23) & (!sk[5]) & (!g74) & (!g495) & (!g1382)) + ((g21) & (g23) & (!sk[5]) & (!g74) & (!g495) & (g1382)) + ((g21) & (g23) & (!sk[5]) & (!g74) & (g495) & (!g1382)) + ((g21) & (g23) & (!sk[5]) & (!g74) & (g495) & (g1382)) + ((g21) & (g23) & (!sk[5]) & (g74) & (!g495) & (!g1382)) + ((g21) & (g23) & (!sk[5]) & (g74) & (!g495) & (g1382)) + ((g21) & (g23) & (!sk[5]) & (g74) & (g495) & (!g1382)) + ((g21) & (g23) & (!sk[5]) & (g74) & (g495) & (g1382)) + ((g21) & (g23) & (sk[5]) & (!g74) & (!g495) & (!g1382)) + ((g21) & (g23) & (sk[5]) & (!g74) & (g495) & (!g1382)));
	assign g1384 = (((!g78) & (!g74) & (!sk[6]) & (g79)) + ((!g78) & (g74) & (!sk[6]) & (!g79)) + ((!g78) & (g74) & (!sk[6]) & (g79)) + ((!g78) & (g74) & (sk[6]) & (!g79)) + ((!g78) & (g74) & (sk[6]) & (g79)) + ((g78) & (!g74) & (!sk[6]) & (g79)) + ((g78) & (g74) & (!sk[6]) & (!g79)) + ((g78) & (g74) & (!sk[6]) & (g79)) + ((g78) & (g74) & (sk[6]) & (!g79)));
	assign g1385 = (((!sk[7]) & (!g74) & (!g175) & (g278)) + ((!sk[7]) & (!g74) & (g175) & (!g278)) + ((!sk[7]) & (!g74) & (g175) & (g278)) + ((!sk[7]) & (g74) & (!g175) & (g278)) + ((!sk[7]) & (g74) & (g175) & (!g278)) + ((!sk[7]) & (g74) & (g175) & (g278)) + ((sk[7]) & (g74) & (!g175) & (g278)) + ((sk[7]) & (g74) & (g175) & (!g278)) + ((sk[7]) & (g74) & (g175) & (g278)));
	assign g1386 = (((!g159) & (!sk[8]) & (!g131) & (g253) & (!g625)) + ((!g159) & (!sk[8]) & (!g131) & (g253) & (g625)) + ((!g159) & (!sk[8]) & (g131) & (g253) & (!g625)) + ((!g159) & (!sk[8]) & (g131) & (g253) & (g625)) + ((!g159) & (sk[8]) & (!g131) & (!g253) & (g625)) + ((!g159) & (sk[8]) & (!g131) & (g253) & (g625)) + ((!g159) & (sk[8]) & (g131) & (!g253) & (g625)) + ((!g159) & (sk[8]) & (g131) & (g253) & (g625)) + ((g159) & (!sk[8]) & (!g131) & (g253) & (!g625)) + ((g159) & (!sk[8]) & (!g131) & (g253) & (g625)) + ((g159) & (!sk[8]) & (g131) & (g253) & (!g625)) + ((g159) & (!sk[8]) & (g131) & (g253) & (g625)) + ((g159) & (sk[8]) & (!g131) & (!g253) & (g625)) + ((g159) & (sk[8]) & (!g131) & (g253) & (g625)) + ((g159) & (sk[8]) & (g131) & (!g253) & (g625)));
	assign g1387 = (((!i_8_) & (!i_6_) & (i_7_) & (!sk[9]) & (!g428) & (g394)) + ((!i_8_) & (!i_6_) & (i_7_) & (!sk[9]) & (g428) & (!g394)) + ((!i_8_) & (!i_6_) & (i_7_) & (!sk[9]) & (g428) & (g394)) + ((!i_8_) & (!i_6_) & (i_7_) & (sk[9]) & (!g428) & (g394)) + ((!i_8_) & (i_6_) & (!i_7_) & (!sk[9]) & (!g428) & (!g394)) + ((!i_8_) & (i_6_) & (!i_7_) & (!sk[9]) & (!g428) & (g394)) + ((!i_8_) & (i_6_) & (!i_7_) & (!sk[9]) & (g428) & (!g394)) + ((!i_8_) & (i_6_) & (!i_7_) & (!sk[9]) & (g428) & (g394)) + ((!i_8_) & (i_6_) & (!i_7_) & (sk[9]) & (!g428) & (g394)) + ((!i_8_) & (i_6_) & (i_7_) & (!sk[9]) & (!g428) & (!g394)) + ((!i_8_) & (i_6_) & (i_7_) & (!sk[9]) & (!g428) & (g394)) + ((!i_8_) & (i_6_) & (i_7_) & (!sk[9]) & (g428) & (!g394)) + ((!i_8_) & (i_6_) & (i_7_) & (!sk[9]) & (g428) & (g394)) + ((i_8_) & (!i_6_) & (i_7_) & (!sk[9]) & (!g428) & (g394)) + ((i_8_) & (!i_6_) & (i_7_) & (!sk[9]) & (g428) & (!g394)) + ((i_8_) & (!i_6_) & (i_7_) & (!sk[9]) & (g428) & (g394)) + ((i_8_) & (i_6_) & (!i_7_) & (!sk[9]) & (!g428) & (!g394)) + ((i_8_) & (i_6_) & (!i_7_) & (!sk[9]) & (!g428) & (g394)) + ((i_8_) & (i_6_) & (!i_7_) & (!sk[9]) & (g428) & (!g394)) + ((i_8_) & (i_6_) & (!i_7_) & (!sk[9]) & (g428) & (g394)) + ((i_8_) & (i_6_) & (i_7_) & (!sk[9]) & (!g428) & (!g394)) + ((i_8_) & (i_6_) & (i_7_) & (!sk[9]) & (!g428) & (g394)) + ((i_8_) & (i_6_) & (i_7_) & (!sk[9]) & (g428) & (!g394)) + ((i_8_) & (i_6_) & (i_7_) & (!sk[9]) & (g428) & (g394)));
	assign g1388 = (((!g25) & (!sk[10]) & (!g102) & (g79) & (!g278) & (g1387)) + ((!g25) & (!sk[10]) & (!g102) & (g79) & (g278) & (!g1387)) + ((!g25) & (!sk[10]) & (!g102) & (g79) & (g278) & (g1387)) + ((!g25) & (!sk[10]) & (g102) & (!g79) & (!g278) & (!g1387)) + ((!g25) & (!sk[10]) & (g102) & (!g79) & (!g278) & (g1387)) + ((!g25) & (!sk[10]) & (g102) & (!g79) & (g278) & (!g1387)) + ((!g25) & (!sk[10]) & (g102) & (!g79) & (g278) & (g1387)) + ((!g25) & (!sk[10]) & (g102) & (g79) & (!g278) & (!g1387)) + ((!g25) & (!sk[10]) & (g102) & (g79) & (!g278) & (g1387)) + ((!g25) & (!sk[10]) & (g102) & (g79) & (g278) & (!g1387)) + ((!g25) & (!sk[10]) & (g102) & (g79) & (g278) & (g1387)) + ((!g25) & (sk[10]) & (!g102) & (!g79) & (!g278) & (!g1387)) + ((!g25) & (sk[10]) & (!g102) & (!g79) & (g278) & (!g1387)) + ((!g25) & (sk[10]) & (!g102) & (g79) & (!g278) & (!g1387)) + ((!g25) & (sk[10]) & (!g102) & (g79) & (g278) & (!g1387)) + ((g25) & (!sk[10]) & (!g102) & (g79) & (!g278) & (g1387)) + ((g25) & (!sk[10]) & (!g102) & (g79) & (g278) & (!g1387)) + ((g25) & (!sk[10]) & (!g102) & (g79) & (g278) & (g1387)) + ((g25) & (!sk[10]) & (g102) & (!g79) & (!g278) & (!g1387)) + ((g25) & (!sk[10]) & (g102) & (!g79) & (!g278) & (g1387)) + ((g25) & (!sk[10]) & (g102) & (!g79) & (g278) & (!g1387)) + ((g25) & (!sk[10]) & (g102) & (!g79) & (g278) & (g1387)) + ((g25) & (!sk[10]) & (g102) & (g79) & (!g278) & (!g1387)) + ((g25) & (!sk[10]) & (g102) & (g79) & (!g278) & (g1387)) + ((g25) & (!sk[10]) & (g102) & (g79) & (g278) & (!g1387)) + ((g25) & (!sk[10]) & (g102) & (g79) & (g278) & (g1387)) + ((g25) & (sk[10]) & (!g102) & (!g79) & (!g278) & (!g1387)) + ((g25) & (sk[10]) & (!g102) & (!g79) & (g278) & (!g1387)) + ((g25) & (sk[10]) & (!g102) & (g79) & (!g278) & (!g1387)) + ((g25) & (sk[10]) & (!g102) & (g79) & (g278) & (!g1387)) + ((g25) & (sk[10]) & (g102) & (g79) & (!g278) & (!g1387)));
	assign g1389 = (((!g131) & (!g177) & (g551) & (!g1386) & (!sk[11]) & (g1388)) + ((!g131) & (!g177) & (g551) & (!g1386) & (sk[11]) & (g1388)) + ((!g131) & (!g177) & (g551) & (g1386) & (!sk[11]) & (!g1388)) + ((!g131) & (!g177) & (g551) & (g1386) & (!sk[11]) & (g1388)) + ((!g131) & (g177) & (!g551) & (!g1386) & (!sk[11]) & (!g1388)) + ((!g131) & (g177) & (!g551) & (!g1386) & (!sk[11]) & (g1388)) + ((!g131) & (g177) & (!g551) & (g1386) & (!sk[11]) & (!g1388)) + ((!g131) & (g177) & (!g551) & (g1386) & (!sk[11]) & (g1388)) + ((!g131) & (g177) & (g551) & (!g1386) & (!sk[11]) & (!g1388)) + ((!g131) & (g177) & (g551) & (!g1386) & (!sk[11]) & (g1388)) + ((!g131) & (g177) & (g551) & (g1386) & (!sk[11]) & (!g1388)) + ((!g131) & (g177) & (g551) & (g1386) & (!sk[11]) & (g1388)) + ((g131) & (!g177) & (!g551) & (!g1386) & (sk[11]) & (g1388)) + ((g131) & (!g177) & (g551) & (!g1386) & (!sk[11]) & (g1388)) + ((g131) & (!g177) & (g551) & (!g1386) & (sk[11]) & (g1388)) + ((g131) & (!g177) & (g551) & (g1386) & (!sk[11]) & (!g1388)) + ((g131) & (!g177) & (g551) & (g1386) & (!sk[11]) & (g1388)) + ((g131) & (g177) & (!g551) & (!g1386) & (!sk[11]) & (!g1388)) + ((g131) & (g177) & (!g551) & (!g1386) & (!sk[11]) & (g1388)) + ((g131) & (g177) & (!g551) & (!g1386) & (sk[11]) & (g1388)) + ((g131) & (g177) & (!g551) & (g1386) & (!sk[11]) & (!g1388)) + ((g131) & (g177) & (!g551) & (g1386) & (!sk[11]) & (g1388)) + ((g131) & (g177) & (g551) & (!g1386) & (!sk[11]) & (!g1388)) + ((g131) & (g177) & (g551) & (!g1386) & (!sk[11]) & (g1388)) + ((g131) & (g177) & (g551) & (!g1386) & (sk[11]) & (g1388)) + ((g131) & (g177) & (g551) & (g1386) & (!sk[11]) & (!g1388)) + ((g131) & (g177) & (g551) & (g1386) & (!sk[11]) & (g1388)));
	assign g1390 = (((!g21) & (!g122) & (!g413) & (sk[12]) & (!g931)) + ((!g21) & (!g122) & (g413) & (!sk[12]) & (!g931)) + ((!g21) & (!g122) & (g413) & (!sk[12]) & (g931)) + ((!g21) & (!g122) & (g413) & (sk[12]) & (!g931)) + ((!g21) & (!g122) & (g413) & (sk[12]) & (g931)) + ((!g21) & (g122) & (!g413) & (sk[12]) & (!g931)) + ((!g21) & (g122) & (g413) & (!sk[12]) & (!g931)) + ((!g21) & (g122) & (g413) & (!sk[12]) & (g931)) + ((!g21) & (g122) & (g413) & (sk[12]) & (!g931)) + ((g21) & (!g122) & (g413) & (!sk[12]) & (!g931)) + ((g21) & (!g122) & (g413) & (!sk[12]) & (g931)) + ((g21) & (!g122) & (g413) & (sk[12]) & (!g931)) + ((g21) & (!g122) & (g413) & (sk[12]) & (g931)) + ((g21) & (g122) & (g413) & (!sk[12]) & (!g931)) + ((g21) & (g122) & (g413) & (!sk[12]) & (g931)) + ((g21) & (g122) & (g413) & (sk[12]) & (!g931)));
	assign g1391 = (((!g1384) & (!g238) & (g1131) & (!g1385) & (g1389) & (g1390)));
	assign g1392 = (((!g1042) & (g1467) & (!g1006) & (g1270) & (g1383) & (g1391)));
	assign g1393 = (((g1172) & (g1224) & (g1319) & (g1368) & (g1381) & (g1392)));
	assign g1394 = (((!g74) & (!sk[16]) & (!g182) & (g183) & (!g699)) + ((!g74) & (!sk[16]) & (!g182) & (g183) & (g699)) + ((!g74) & (!sk[16]) & (g182) & (g183) & (!g699)) + ((!g74) & (!sk[16]) & (g182) & (g183) & (g699)) + ((g74) & (!sk[16]) & (!g182) & (g183) & (!g699)) + ((g74) & (!sk[16]) & (!g182) & (g183) & (g699)) + ((g74) & (!sk[16]) & (g182) & (g183) & (!g699)) + ((g74) & (!sk[16]) & (g182) & (g183) & (g699)) + ((g74) & (sk[16]) & (!g182) & (!g183) & (!g699)) + ((g74) & (sk[16]) & (!g182) & (g183) & (!g699)) + ((g74) & (sk[16]) & (!g182) & (g183) & (g699)) + ((g74) & (sk[16]) & (g182) & (!g183) & (!g699)) + ((g74) & (sk[16]) & (g182) & (!g183) & (g699)) + ((g74) & (sk[16]) & (g182) & (g183) & (!g699)) + ((g74) & (sk[16]) & (g182) & (g183) & (g699)));
	assign g1395 = (((!g355) & (!g83) & (!g356) & (!g629) & (sk[17]) & (!g1394)) + ((!g355) & (!g83) & (!g356) & (g629) & (sk[17]) & (!g1394)) + ((!g355) & (!g83) & (g356) & (!g629) & (!sk[17]) & (g1394)) + ((!g355) & (!g83) & (g356) & (!g629) & (sk[17]) & (!g1394)) + ((!g355) & (!g83) & (g356) & (g629) & (!sk[17]) & (!g1394)) + ((!g355) & (!g83) & (g356) & (g629) & (!sk[17]) & (g1394)) + ((!g355) & (g83) & (!g356) & (!g629) & (!sk[17]) & (!g1394)) + ((!g355) & (g83) & (!g356) & (!g629) & (!sk[17]) & (g1394)) + ((!g355) & (g83) & (!g356) & (!g629) & (sk[17]) & (!g1394)) + ((!g355) & (g83) & (!g356) & (g629) & (!sk[17]) & (!g1394)) + ((!g355) & (g83) & (!g356) & (g629) & (!sk[17]) & (g1394)) + ((!g355) & (g83) & (!g356) & (g629) & (sk[17]) & (!g1394)) + ((!g355) & (g83) & (g356) & (!g629) & (!sk[17]) & (!g1394)) + ((!g355) & (g83) & (g356) & (!g629) & (!sk[17]) & (g1394)) + ((!g355) & (g83) & (g356) & (!g629) & (sk[17]) & (!g1394)) + ((!g355) & (g83) & (g356) & (g629) & (!sk[17]) & (!g1394)) + ((!g355) & (g83) & (g356) & (g629) & (!sk[17]) & (g1394)) + ((g355) & (!g83) & (!g356) & (!g629) & (sk[17]) & (!g1394)) + ((g355) & (!g83) & (!g356) & (g629) & (sk[17]) & (!g1394)) + ((g355) & (!g83) & (g356) & (!g629) & (!sk[17]) & (g1394)) + ((g355) & (!g83) & (g356) & (!g629) & (sk[17]) & (!g1394)) + ((g355) & (!g83) & (g356) & (g629) & (!sk[17]) & (!g1394)) + ((g355) & (!g83) & (g356) & (g629) & (!sk[17]) & (g1394)) + ((g355) & (g83) & (!g356) & (!g629) & (!sk[17]) & (!g1394)) + ((g355) & (g83) & (!g356) & (!g629) & (!sk[17]) & (g1394)) + ((g355) & (g83) & (!g356) & (!g629) & (sk[17]) & (!g1394)) + ((g355) & (g83) & (!g356) & (g629) & (!sk[17]) & (!g1394)) + ((g355) & (g83) & (!g356) & (g629) & (!sk[17]) & (g1394)) + ((g355) & (g83) & (!g356) & (g629) & (sk[17]) & (!g1394)) + ((g355) & (g83) & (g356) & (!g629) & (!sk[17]) & (!g1394)) + ((g355) & (g83) & (g356) & (!g629) & (!sk[17]) & (g1394)) + ((g355) & (g83) & (g356) & (g629) & (!sk[17]) & (!g1394)) + ((g355) & (g83) & (g356) & (g629) & (!sk[17]) & (g1394)));
	assign g1396 = (((!g102) & (!g699) & (!sk[18]) & (g700)) + ((!g102) & (g699) & (!sk[18]) & (!g700)) + ((!g102) & (g699) & (!sk[18]) & (g700)) + ((g102) & (!g699) & (!sk[18]) & (g700)) + ((g102) & (!g699) & (sk[18]) & (!g700)) + ((g102) & (!g699) & (sk[18]) & (g700)) + ((g102) & (g699) & (!sk[18]) & (!g700)) + ((g102) & (g699) & (!sk[18]) & (g700)) + ((g102) & (g699) & (sk[18]) & (!g700)));
	assign g1397 = (((!g24) & (!g74) & (!sk[19]) & (g445)) + ((!g24) & (g74) & (!sk[19]) & (!g445)) + ((!g24) & (g74) & (!sk[19]) & (g445)) + ((!g24) & (g74) & (sk[19]) & (g445)) + ((g24) & (!g74) & (!sk[19]) & (g445)) + ((g24) & (g74) & (!sk[19]) & (!g445)) + ((g24) & (g74) & (!sk[19]) & (g445)));
	assign g1398 = (((!g24) & (!g68) & (!sk[20]) & (g102) & (!g83)) + ((!g24) & (!g68) & (!sk[20]) & (g102) & (g83)) + ((!g24) & (!g68) & (sk[20]) & (g102) & (g83)) + ((!g24) & (g68) & (!sk[20]) & (g102) & (!g83)) + ((!g24) & (g68) & (!sk[20]) & (g102) & (g83)) + ((!g24) & (g68) & (sk[20]) & (g102) & (g83)) + ((g24) & (!g68) & (!sk[20]) & (g102) & (!g83)) + ((g24) & (!g68) & (!sk[20]) & (g102) & (g83)) + ((g24) & (!g68) & (sk[20]) & (g102) & (g83)) + ((g24) & (g68) & (!sk[20]) & (g102) & (!g83)) + ((g24) & (g68) & (!sk[20]) & (g102) & (g83)));
	assign g1399 = (((!g102) & (!g501) & (!sk[21]) & (g543)) + ((!g102) & (g501) & (!sk[21]) & (!g543)) + ((!g102) & (g501) & (!sk[21]) & (g543)) + ((g102) & (!g501) & (!sk[21]) & (g543)) + ((g102) & (!g501) & (sk[21]) & (g543)) + ((g102) & (g501) & (!sk[21]) & (!g543)) + ((g102) & (g501) & (!sk[21]) & (g543)) + ((g102) & (g501) & (sk[21]) & (!g543)) + ((g102) & (g501) & (sk[21]) & (g543)));
	assign g1400 = (((!i_8_) & (!g19) & (!sk[22]) & (g73) & (!g76) & (g83)) + ((!i_8_) & (!g19) & (!sk[22]) & (g73) & (g76) & (!g83)) + ((!i_8_) & (!g19) & (!sk[22]) & (g73) & (g76) & (g83)) + ((!i_8_) & (!g19) & (sk[22]) & (g73) & (!g76) & (g83)) + ((!i_8_) & (g19) & (!sk[22]) & (!g73) & (!g76) & (!g83)) + ((!i_8_) & (g19) & (!sk[22]) & (!g73) & (!g76) & (g83)) + ((!i_8_) & (g19) & (!sk[22]) & (!g73) & (g76) & (!g83)) + ((!i_8_) & (g19) & (!sk[22]) & (!g73) & (g76) & (g83)) + ((!i_8_) & (g19) & (!sk[22]) & (g73) & (!g76) & (!g83)) + ((!i_8_) & (g19) & (!sk[22]) & (g73) & (!g76) & (g83)) + ((!i_8_) & (g19) & (!sk[22]) & (g73) & (g76) & (!g83)) + ((!i_8_) & (g19) & (!sk[22]) & (g73) & (g76) & (g83)) + ((!i_8_) & (g19) & (sk[22]) & (g73) & (!g76) & (g83)) + ((!i_8_) & (g19) & (sk[22]) & (g73) & (g76) & (g83)) + ((i_8_) & (!g19) & (!sk[22]) & (g73) & (!g76) & (g83)) + ((i_8_) & (!g19) & (!sk[22]) & (g73) & (g76) & (!g83)) + ((i_8_) & (!g19) & (!sk[22]) & (g73) & (g76) & (g83)) + ((i_8_) & (g19) & (!sk[22]) & (!g73) & (!g76) & (!g83)) + ((i_8_) & (g19) & (!sk[22]) & (!g73) & (!g76) & (g83)) + ((i_8_) & (g19) & (!sk[22]) & (!g73) & (g76) & (!g83)) + ((i_8_) & (g19) & (!sk[22]) & (!g73) & (g76) & (g83)) + ((i_8_) & (g19) & (!sk[22]) & (g73) & (!g76) & (!g83)) + ((i_8_) & (g19) & (!sk[22]) & (g73) & (!g76) & (g83)) + ((i_8_) & (g19) & (!sk[22]) & (g73) & (g76) & (!g83)) + ((i_8_) & (g19) & (!sk[22]) & (g73) & (g76) & (g83)));
	assign g1401 = (((!i_8_) & (!i_6_) & (!sk[23]) & (i_7_) & (!g445) & (g394)) + ((!i_8_) & (!i_6_) & (!sk[23]) & (i_7_) & (g445) & (!g394)) + ((!i_8_) & (!i_6_) & (!sk[23]) & (i_7_) & (g445) & (g394)) + ((!i_8_) & (!i_6_) & (sk[23]) & (i_7_) & (g445) & (g394)) + ((!i_8_) & (i_6_) & (!sk[23]) & (!i_7_) & (!g445) & (!g394)) + ((!i_8_) & (i_6_) & (!sk[23]) & (!i_7_) & (!g445) & (g394)) + ((!i_8_) & (i_6_) & (!sk[23]) & (!i_7_) & (g445) & (!g394)) + ((!i_8_) & (i_6_) & (!sk[23]) & (!i_7_) & (g445) & (g394)) + ((!i_8_) & (i_6_) & (!sk[23]) & (i_7_) & (!g445) & (!g394)) + ((!i_8_) & (i_6_) & (!sk[23]) & (i_7_) & (!g445) & (g394)) + ((!i_8_) & (i_6_) & (!sk[23]) & (i_7_) & (g445) & (!g394)) + ((!i_8_) & (i_6_) & (!sk[23]) & (i_7_) & (g445) & (g394)) + ((!i_8_) & (i_6_) & (sk[23]) & (!i_7_) & (g445) & (g394)) + ((i_8_) & (!i_6_) & (!sk[23]) & (i_7_) & (!g445) & (g394)) + ((i_8_) & (!i_6_) & (!sk[23]) & (i_7_) & (g445) & (!g394)) + ((i_8_) & (!i_6_) & (!sk[23]) & (i_7_) & (g445) & (g394)) + ((i_8_) & (i_6_) & (!sk[23]) & (!i_7_) & (!g445) & (!g394)) + ((i_8_) & (i_6_) & (!sk[23]) & (!i_7_) & (!g445) & (g394)) + ((i_8_) & (i_6_) & (!sk[23]) & (!i_7_) & (g445) & (!g394)) + ((i_8_) & (i_6_) & (!sk[23]) & (!i_7_) & (g445) & (g394)) + ((i_8_) & (i_6_) & (!sk[23]) & (i_7_) & (!g445) & (!g394)) + ((i_8_) & (i_6_) & (!sk[23]) & (i_7_) & (!g445) & (g394)) + ((i_8_) & (i_6_) & (!sk[23]) & (i_7_) & (g445) & (!g394)) + ((i_8_) & (i_6_) & (!sk[23]) & (i_7_) & (g445) & (g394)));
	assign g1402 = (((!i_8_) & (!sk[24]) & (!g73) & (g82) & (!g295) & (g1401)) + ((!i_8_) & (!sk[24]) & (!g73) & (g82) & (g295) & (!g1401)) + ((!i_8_) & (!sk[24]) & (!g73) & (g82) & (g295) & (g1401)) + ((!i_8_) & (!sk[24]) & (g73) & (!g82) & (!g295) & (!g1401)) + ((!i_8_) & (!sk[24]) & (g73) & (!g82) & (!g295) & (g1401)) + ((!i_8_) & (!sk[24]) & (g73) & (!g82) & (g295) & (!g1401)) + ((!i_8_) & (!sk[24]) & (g73) & (!g82) & (g295) & (g1401)) + ((!i_8_) & (!sk[24]) & (g73) & (g82) & (!g295) & (!g1401)) + ((!i_8_) & (!sk[24]) & (g73) & (g82) & (!g295) & (g1401)) + ((!i_8_) & (!sk[24]) & (g73) & (g82) & (g295) & (!g1401)) + ((!i_8_) & (!sk[24]) & (g73) & (g82) & (g295) & (g1401)) + ((!i_8_) & (sk[24]) & (!g73) & (!g82) & (!g295) & (!g1401)) + ((!i_8_) & (sk[24]) & (!g73) & (!g82) & (g295) & (!g1401)) + ((!i_8_) & (sk[24]) & (!g73) & (g82) & (!g295) & (!g1401)) + ((!i_8_) & (sk[24]) & (!g73) & (g82) & (g295) & (!g1401)) + ((!i_8_) & (sk[24]) & (g73) & (!g82) & (!g295) & (!g1401)) + ((i_8_) & (!sk[24]) & (!g73) & (g82) & (!g295) & (g1401)) + ((i_8_) & (!sk[24]) & (!g73) & (g82) & (g295) & (!g1401)) + ((i_8_) & (!sk[24]) & (!g73) & (g82) & (g295) & (g1401)) + ((i_8_) & (!sk[24]) & (g73) & (!g82) & (!g295) & (!g1401)) + ((i_8_) & (!sk[24]) & (g73) & (!g82) & (!g295) & (g1401)) + ((i_8_) & (!sk[24]) & (g73) & (!g82) & (g295) & (!g1401)) + ((i_8_) & (!sk[24]) & (g73) & (!g82) & (g295) & (g1401)) + ((i_8_) & (!sk[24]) & (g73) & (g82) & (!g295) & (!g1401)) + ((i_8_) & (!sk[24]) & (g73) & (g82) & (!g295) & (g1401)) + ((i_8_) & (!sk[24]) & (g73) & (g82) & (g295) & (!g1401)) + ((i_8_) & (!sk[24]) & (g73) & (g82) & (g295) & (g1401)) + ((i_8_) & (sk[24]) & (!g73) & (!g82) & (!g295) & (!g1401)) + ((i_8_) & (sk[24]) & (!g73) & (!g82) & (g295) & (!g1401)) + ((i_8_) & (sk[24]) & (!g73) & (g82) & (!g295) & (!g1401)) + ((i_8_) & (sk[24]) & (!g73) & (g82) & (g295) & (!g1401)) + ((i_8_) & (sk[24]) & (g73) & (!g82) & (!g295) & (!g1401)) + ((i_8_) & (sk[24]) & (g73) & (!g82) & (g295) & (!g1401)) + ((i_8_) & (sk[24]) & (g73) & (g82) & (!g295) & (!g1401)) + ((i_8_) & (sk[24]) & (g73) & (g82) & (g295) & (!g1401)));
	assign g1403 = (((!g1398) & (!g1399) & (!g583) & (!g1400) & (sk[25]) & (g1402)) + ((!g1398) & (!g1399) & (g583) & (!g1400) & (!sk[25]) & (g1402)) + ((!g1398) & (!g1399) & (g583) & (g1400) & (!sk[25]) & (!g1402)) + ((!g1398) & (!g1399) & (g583) & (g1400) & (!sk[25]) & (g1402)) + ((!g1398) & (g1399) & (!g583) & (!g1400) & (!sk[25]) & (!g1402)) + ((!g1398) & (g1399) & (!g583) & (!g1400) & (!sk[25]) & (g1402)) + ((!g1398) & (g1399) & (!g583) & (g1400) & (!sk[25]) & (!g1402)) + ((!g1398) & (g1399) & (!g583) & (g1400) & (!sk[25]) & (g1402)) + ((!g1398) & (g1399) & (g583) & (!g1400) & (!sk[25]) & (!g1402)) + ((!g1398) & (g1399) & (g583) & (!g1400) & (!sk[25]) & (g1402)) + ((!g1398) & (g1399) & (g583) & (g1400) & (!sk[25]) & (!g1402)) + ((!g1398) & (g1399) & (g583) & (g1400) & (!sk[25]) & (g1402)) + ((g1398) & (!g1399) & (g583) & (!g1400) & (!sk[25]) & (g1402)) + ((g1398) & (!g1399) & (g583) & (g1400) & (!sk[25]) & (!g1402)) + ((g1398) & (!g1399) & (g583) & (g1400) & (!sk[25]) & (g1402)) + ((g1398) & (g1399) & (!g583) & (!g1400) & (!sk[25]) & (!g1402)) + ((g1398) & (g1399) & (!g583) & (!g1400) & (!sk[25]) & (g1402)) + ((g1398) & (g1399) & (!g583) & (g1400) & (!sk[25]) & (!g1402)) + ((g1398) & (g1399) & (!g583) & (g1400) & (!sk[25]) & (g1402)) + ((g1398) & (g1399) & (g583) & (!g1400) & (!sk[25]) & (!g1402)) + ((g1398) & (g1399) & (g583) & (!g1400) & (!sk[25]) & (g1402)) + ((g1398) & (g1399) & (g583) & (g1400) & (!sk[25]) & (!g1402)) + ((g1398) & (g1399) & (g583) & (g1400) & (!sk[25]) & (g1402)));
	assign g1404 = (((!sk[26]) & (!g131) & (!g182) & (g183) & (!g295) & (g700)) + ((!sk[26]) & (!g131) & (!g182) & (g183) & (g295) & (!g700)) + ((!sk[26]) & (!g131) & (!g182) & (g183) & (g295) & (g700)) + ((!sk[26]) & (!g131) & (g182) & (!g183) & (!g295) & (!g700)) + ((!sk[26]) & (!g131) & (g182) & (!g183) & (!g295) & (g700)) + ((!sk[26]) & (!g131) & (g182) & (!g183) & (g295) & (!g700)) + ((!sk[26]) & (!g131) & (g182) & (!g183) & (g295) & (g700)) + ((!sk[26]) & (!g131) & (g182) & (g183) & (!g295) & (!g700)) + ((!sk[26]) & (!g131) & (g182) & (g183) & (!g295) & (g700)) + ((!sk[26]) & (!g131) & (g182) & (g183) & (g295) & (!g700)) + ((!sk[26]) & (!g131) & (g182) & (g183) & (g295) & (g700)) + ((!sk[26]) & (g131) & (!g182) & (g183) & (!g295) & (g700)) + ((!sk[26]) & (g131) & (!g182) & (g183) & (g295) & (!g700)) + ((!sk[26]) & (g131) & (!g182) & (g183) & (g295) & (g700)) + ((!sk[26]) & (g131) & (g182) & (!g183) & (!g295) & (!g700)) + ((!sk[26]) & (g131) & (g182) & (!g183) & (!g295) & (g700)) + ((!sk[26]) & (g131) & (g182) & (!g183) & (g295) & (!g700)) + ((!sk[26]) & (g131) & (g182) & (!g183) & (g295) & (g700)) + ((!sk[26]) & (g131) & (g182) & (g183) & (!g295) & (!g700)) + ((!sk[26]) & (g131) & (g182) & (g183) & (!g295) & (g700)) + ((!sk[26]) & (g131) & (g182) & (g183) & (g295) & (!g700)) + ((!sk[26]) & (g131) & (g182) & (g183) & (g295) & (g700)) + ((sk[26]) & (!g131) & (!g182) & (!g183) & (!g295) & (!g700)) + ((sk[26]) & (!g131) & (!g182) & (!g183) & (g295) & (!g700)) + ((sk[26]) & (!g131) & (!g182) & (!g183) & (g295) & (g700)) + ((sk[26]) & (!g131) & (!g182) & (g183) & (!g295) & (!g700)) + ((sk[26]) & (!g131) & (!g182) & (g183) & (!g295) & (g700)) + ((sk[26]) & (!g131) & (!g182) & (g183) & (g295) & (!g700)) + ((sk[26]) & (!g131) & (!g182) & (g183) & (g295) & (g700)) + ((sk[26]) & (!g131) & (g182) & (!g183) & (!g295) & (!g700)) + ((sk[26]) & (!g131) & (g182) & (!g183) & (!g295) & (g700)) + ((sk[26]) & (!g131) & (g182) & (!g183) & (g295) & (!g700)) + ((sk[26]) & (!g131) & (g182) & (!g183) & (g295) & (g700)) + ((sk[26]) & (!g131) & (g182) & (g183) & (!g295) & (!g700)) + ((sk[26]) & (!g131) & (g182) & (g183) & (!g295) & (g700)) + ((sk[26]) & (!g131) & (g182) & (g183) & (g295) & (!g700)) + ((sk[26]) & (!g131) & (g182) & (g183) & (g295) & (g700)));
	assign g1405 = (((!g157) & (!g74) & (!g183) & (!g892) & (!g608) & (!g1404)) + ((!g157) & (!g74) & (!g183) & (!g892) & (g608) & (!g1404)) + ((!g157) & (!g74) & (!g183) & (g892) & (!g608) & (!g1404)) + ((!g157) & (!g74) & (!g183) & (g892) & (g608) & (!g1404)) + ((!g157) & (!g74) & (g183) & (!g892) & (!g608) & (!g1404)) + ((!g157) & (!g74) & (g183) & (!g892) & (g608) & (!g1404)) + ((!g157) & (!g74) & (g183) & (g892) & (!g608) & (!g1404)) + ((!g157) & (!g74) & (g183) & (g892) & (g608) & (!g1404)) + ((!g157) & (g74) & (!g183) & (!g892) & (!g608) & (!g1404)) + ((!g157) & (g74) & (!g183) & (!g892) & (g608) & (!g1404)) + ((!g157) & (g74) & (g183) & (!g892) & (!g608) & (!g1404)) + ((!g157) & (g74) & (g183) & (!g892) & (g608) & (!g1404)) + ((g157) & (!g74) & (!g183) & (!g892) & (g608) & (!g1404)) + ((g157) & (g74) & (!g183) & (!g892) & (g608) & (!g1404)));
	assign g1406 = (((!g159) & (!g214) & (!g438) & (!g770) & (sk[28]) & (g930)) + ((!g159) & (!g214) & (g438) & (!g770) & (!sk[28]) & (g930)) + ((!g159) & (!g214) & (g438) & (!g770) & (sk[28]) & (!g930)) + ((!g159) & (!g214) & (g438) & (!g770) & (sk[28]) & (g930)) + ((!g159) & (!g214) & (g438) & (g770) & (!sk[28]) & (!g930)) + ((!g159) & (!g214) & (g438) & (g770) & (!sk[28]) & (g930)) + ((!g159) & (g214) & (!g438) & (!g770) & (!sk[28]) & (!g930)) + ((!g159) & (g214) & (!g438) & (!g770) & (!sk[28]) & (g930)) + ((!g159) & (g214) & (!g438) & (g770) & (!sk[28]) & (!g930)) + ((!g159) & (g214) & (!g438) & (g770) & (!sk[28]) & (g930)) + ((!g159) & (g214) & (g438) & (!g770) & (!sk[28]) & (!g930)) + ((!g159) & (g214) & (g438) & (!g770) & (!sk[28]) & (g930)) + ((!g159) & (g214) & (g438) & (g770) & (!sk[28]) & (!g930)) + ((!g159) & (g214) & (g438) & (g770) & (!sk[28]) & (g930)) + ((g159) & (!g214) & (!g438) & (!g770) & (sk[28]) & (g930)) + ((g159) & (!g214) & (g438) & (!g770) & (!sk[28]) & (g930)) + ((g159) & (!g214) & (g438) & (!g770) & (sk[28]) & (!g930)) + ((g159) & (!g214) & (g438) & (!g770) & (sk[28]) & (g930)) + ((g159) & (!g214) & (g438) & (g770) & (!sk[28]) & (!g930)) + ((g159) & (!g214) & (g438) & (g770) & (!sk[28]) & (g930)) + ((g159) & (!g214) & (g438) & (g770) & (sk[28]) & (!g930)) + ((g159) & (!g214) & (g438) & (g770) & (sk[28]) & (g930)) + ((g159) & (g214) & (!g438) & (!g770) & (!sk[28]) & (!g930)) + ((g159) & (g214) & (!g438) & (!g770) & (!sk[28]) & (g930)) + ((g159) & (g214) & (!g438) & (g770) & (!sk[28]) & (!g930)) + ((g159) & (g214) & (!g438) & (g770) & (!sk[28]) & (g930)) + ((g159) & (g214) & (g438) & (!g770) & (!sk[28]) & (!g930)) + ((g159) & (g214) & (g438) & (!g770) & (!sk[28]) & (g930)) + ((g159) & (g214) & (g438) & (g770) & (!sk[28]) & (!g930)) + ((g159) & (g214) & (g438) & (g770) & (!sk[28]) & (g930)));
	assign g1407 = (((!sk[29]) & (!g1396) & (!g1397) & (g1403) & (!g1405) & (g1406)) + ((!sk[29]) & (!g1396) & (!g1397) & (g1403) & (g1405) & (!g1406)) + ((!sk[29]) & (!g1396) & (!g1397) & (g1403) & (g1405) & (g1406)) + ((!sk[29]) & (!g1396) & (g1397) & (!g1403) & (!g1405) & (!g1406)) + ((!sk[29]) & (!g1396) & (g1397) & (!g1403) & (!g1405) & (g1406)) + ((!sk[29]) & (!g1396) & (g1397) & (!g1403) & (g1405) & (!g1406)) + ((!sk[29]) & (!g1396) & (g1397) & (!g1403) & (g1405) & (g1406)) + ((!sk[29]) & (!g1396) & (g1397) & (g1403) & (!g1405) & (!g1406)) + ((!sk[29]) & (!g1396) & (g1397) & (g1403) & (!g1405) & (g1406)) + ((!sk[29]) & (!g1396) & (g1397) & (g1403) & (g1405) & (!g1406)) + ((!sk[29]) & (!g1396) & (g1397) & (g1403) & (g1405) & (g1406)) + ((!sk[29]) & (g1396) & (!g1397) & (g1403) & (!g1405) & (g1406)) + ((!sk[29]) & (g1396) & (!g1397) & (g1403) & (g1405) & (!g1406)) + ((!sk[29]) & (g1396) & (!g1397) & (g1403) & (g1405) & (g1406)) + ((!sk[29]) & (g1396) & (g1397) & (!g1403) & (!g1405) & (!g1406)) + ((!sk[29]) & (g1396) & (g1397) & (!g1403) & (!g1405) & (g1406)) + ((!sk[29]) & (g1396) & (g1397) & (!g1403) & (g1405) & (!g1406)) + ((!sk[29]) & (g1396) & (g1397) & (!g1403) & (g1405) & (g1406)) + ((!sk[29]) & (g1396) & (g1397) & (g1403) & (!g1405) & (!g1406)) + ((!sk[29]) & (g1396) & (g1397) & (g1403) & (!g1405) & (g1406)) + ((!sk[29]) & (g1396) & (g1397) & (g1403) & (g1405) & (!g1406)) + ((!sk[29]) & (g1396) & (g1397) & (g1403) & (g1405) & (g1406)) + ((sk[29]) & (!g1396) & (!g1397) & (g1403) & (g1405) & (g1406)));
	assign g1408 = (((!i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g445) & (!g130)) + ((!i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g445) & (!g130)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g445) & (!g130)) + ((i_15_) & (!i_12_) & (!i_13_) & (!i_14_) & (g445) & (!g130)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g445) & (!g130)) + ((i_15_) & (i_12_) & (!i_13_) & (!i_14_) & (g445) & (!g130)) + ((i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g445) & (!g130)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g445) & (!g130)));
	assign g1409 = (((!g157) & (!g131) & (!g501) & (sk[31]) & (g543)) + ((!g157) & (!g131) & (g501) & (!sk[31]) & (!g543)) + ((!g157) & (!g131) & (g501) & (!sk[31]) & (g543)) + ((!g157) & (!g131) & (g501) & (sk[31]) & (g543)) + ((!g157) & (g131) & (g501) & (!sk[31]) & (!g543)) + ((!g157) & (g131) & (g501) & (!sk[31]) & (g543)) + ((g157) & (!g131) & (!g501) & (sk[31]) & (g543)) + ((g157) & (!g131) & (g501) & (!sk[31]) & (!g543)) + ((g157) & (!g131) & (g501) & (!sk[31]) & (g543)) + ((g157) & (!g131) & (g501) & (sk[31]) & (!g543)) + ((g157) & (!g131) & (g501) & (sk[31]) & (g543)) + ((g157) & (g131) & (g501) & (!sk[31]) & (!g543)) + ((g157) & (g131) & (g501) & (!sk[31]) & (g543)) + ((g157) & (g131) & (g501) & (sk[31]) & (!g543)) + ((g157) & (g131) & (g501) & (sk[31]) & (g543)));
	assign g1410 = (((!g157) & (!g159) & (!g253) & (!g335) & (!g597) & (!g850)) + ((!g157) & (!g159) & (g253) & (!g335) & (!g597) & (!g850)) + ((!g157) & (!g159) & (g253) & (g335) & (!g597) & (!g850)) + ((!g157) & (g159) & (!g253) & (!g335) & (!g597) & (!g850)) + ((!g157) & (g159) & (!g253) & (!g335) & (!g597) & (g850)) + ((!g157) & (g159) & (!g253) & (!g335) & (g597) & (!g850)) + ((!g157) & (g159) & (!g253) & (!g335) & (g597) & (g850)) + ((!g157) & (g159) & (g253) & (!g335) & (!g597) & (!g850)) + ((!g157) & (g159) & (g253) & (!g335) & (!g597) & (g850)) + ((!g157) & (g159) & (g253) & (!g335) & (g597) & (!g850)) + ((!g157) & (g159) & (g253) & (!g335) & (g597) & (g850)) + ((!g157) & (g159) & (g253) & (g335) & (!g597) & (!g850)) + ((!g157) & (g159) & (g253) & (g335) & (!g597) & (g850)) + ((!g157) & (g159) & (g253) & (g335) & (g597) & (!g850)) + ((!g157) & (g159) & (g253) & (g335) & (g597) & (g850)) + ((g157) & (!g159) & (!g253) & (!g335) & (!g597) & (!g850)) + ((g157) & (!g159) & (g253) & (!g335) & (!g597) & (!g850)) + ((g157) & (!g159) & (g253) & (g335) & (!g597) & (!g850)) + ((g157) & (g159) & (!g253) & (!g335) & (!g597) & (!g850)) + ((g157) & (g159) & (!g253) & (!g335) & (!g597) & (g850)) + ((g157) & (g159) & (g253) & (!g335) & (!g597) & (!g850)) + ((g157) & (g159) & (g253) & (!g335) & (!g597) & (g850)) + ((g157) & (g159) & (g253) & (g335) & (!g597) & (!g850)) + ((g157) & (g159) & (g253) & (g335) & (!g597) & (g850)));
	assign g1411 = (((!sk[33]) & (!g103) & (!g253) & (g237) & (!g629) & (g1410)) + ((!sk[33]) & (!g103) & (!g253) & (g237) & (g629) & (!g1410)) + ((!sk[33]) & (!g103) & (!g253) & (g237) & (g629) & (g1410)) + ((!sk[33]) & (!g103) & (g253) & (!g237) & (!g629) & (!g1410)) + ((!sk[33]) & (!g103) & (g253) & (!g237) & (!g629) & (g1410)) + ((!sk[33]) & (!g103) & (g253) & (!g237) & (g629) & (!g1410)) + ((!sk[33]) & (!g103) & (g253) & (!g237) & (g629) & (g1410)) + ((!sk[33]) & (!g103) & (g253) & (g237) & (!g629) & (!g1410)) + ((!sk[33]) & (!g103) & (g253) & (g237) & (!g629) & (g1410)) + ((!sk[33]) & (!g103) & (g253) & (g237) & (g629) & (!g1410)) + ((!sk[33]) & (!g103) & (g253) & (g237) & (g629) & (g1410)) + ((!sk[33]) & (g103) & (!g253) & (g237) & (!g629) & (g1410)) + ((!sk[33]) & (g103) & (!g253) & (g237) & (g629) & (!g1410)) + ((!sk[33]) & (g103) & (!g253) & (g237) & (g629) & (g1410)) + ((!sk[33]) & (g103) & (g253) & (!g237) & (!g629) & (!g1410)) + ((!sk[33]) & (g103) & (g253) & (!g237) & (!g629) & (g1410)) + ((!sk[33]) & (g103) & (g253) & (!g237) & (g629) & (!g1410)) + ((!sk[33]) & (g103) & (g253) & (!g237) & (g629) & (g1410)) + ((!sk[33]) & (g103) & (g253) & (g237) & (!g629) & (!g1410)) + ((!sk[33]) & (g103) & (g253) & (g237) & (!g629) & (g1410)) + ((!sk[33]) & (g103) & (g253) & (g237) & (g629) & (!g1410)) + ((!sk[33]) & (g103) & (g253) & (g237) & (g629) & (g1410)) + ((sk[33]) & (!g103) & (!g253) & (!g237) & (!g629) & (g1410)) + ((sk[33]) & (!g103) & (g253) & (!g237) & (!g629) & (g1410)) + ((sk[33]) & (!g103) & (g253) & (!g237) & (g629) & (g1410)));
	assign g1412 = (((!sk[34]) & (!i_4_) & (!i_3_) & (i_5_) & (!g83) & (g735)) + ((!sk[34]) & (!i_4_) & (!i_3_) & (i_5_) & (g83) & (!g735)) + ((!sk[34]) & (!i_4_) & (!i_3_) & (i_5_) & (g83) & (g735)) + ((!sk[34]) & (!i_4_) & (i_3_) & (!i_5_) & (!g83) & (!g735)) + ((!sk[34]) & (!i_4_) & (i_3_) & (!i_5_) & (!g83) & (g735)) + ((!sk[34]) & (!i_4_) & (i_3_) & (!i_5_) & (g83) & (!g735)) + ((!sk[34]) & (!i_4_) & (i_3_) & (!i_5_) & (g83) & (g735)) + ((!sk[34]) & (!i_4_) & (i_3_) & (i_5_) & (!g83) & (!g735)) + ((!sk[34]) & (!i_4_) & (i_3_) & (i_5_) & (!g83) & (g735)) + ((!sk[34]) & (!i_4_) & (i_3_) & (i_5_) & (g83) & (!g735)) + ((!sk[34]) & (!i_4_) & (i_3_) & (i_5_) & (g83) & (g735)) + ((!sk[34]) & (i_4_) & (!i_3_) & (i_5_) & (!g83) & (g735)) + ((!sk[34]) & (i_4_) & (!i_3_) & (i_5_) & (g83) & (!g735)) + ((!sk[34]) & (i_4_) & (!i_3_) & (i_5_) & (g83) & (g735)) + ((!sk[34]) & (i_4_) & (i_3_) & (!i_5_) & (!g83) & (!g735)) + ((!sk[34]) & (i_4_) & (i_3_) & (!i_5_) & (!g83) & (g735)) + ((!sk[34]) & (i_4_) & (i_3_) & (!i_5_) & (g83) & (!g735)) + ((!sk[34]) & (i_4_) & (i_3_) & (!i_5_) & (g83) & (g735)) + ((!sk[34]) & (i_4_) & (i_3_) & (i_5_) & (!g83) & (!g735)) + ((!sk[34]) & (i_4_) & (i_3_) & (i_5_) & (!g83) & (g735)) + ((!sk[34]) & (i_4_) & (i_3_) & (i_5_) & (g83) & (!g735)) + ((!sk[34]) & (i_4_) & (i_3_) & (i_5_) & (g83) & (g735)) + ((sk[34]) & (!i_4_) & (!i_3_) & (i_5_) & (g83) & (g735)) + ((sk[34]) & (i_4_) & (!i_3_) & (!i_5_) & (g83) & (g735)));
	assign g1413 = (((!g2) & (!g54) & (g71) & (!g723) & (!sk[35]) & (g1412)) + ((!g2) & (!g54) & (g71) & (g723) & (!sk[35]) & (!g1412)) + ((!g2) & (!g54) & (g71) & (g723) & (!sk[35]) & (g1412)) + ((!g2) & (g54) & (!g71) & (!g723) & (!sk[35]) & (!g1412)) + ((!g2) & (g54) & (!g71) & (!g723) & (!sk[35]) & (g1412)) + ((!g2) & (g54) & (!g71) & (g723) & (!sk[35]) & (!g1412)) + ((!g2) & (g54) & (!g71) & (g723) & (!sk[35]) & (g1412)) + ((!g2) & (g54) & (g71) & (!g723) & (!sk[35]) & (!g1412)) + ((!g2) & (g54) & (g71) & (!g723) & (!sk[35]) & (g1412)) + ((!g2) & (g54) & (g71) & (g723) & (!sk[35]) & (!g1412)) + ((!g2) & (g54) & (g71) & (g723) & (!sk[35]) & (g1412)) + ((g2) & (!g54) & (g71) & (!g723) & (!sk[35]) & (g1412)) + ((g2) & (!g54) & (g71) & (!g723) & (sk[35]) & (g1412)) + ((g2) & (!g54) & (g71) & (g723) & (!sk[35]) & (!g1412)) + ((g2) & (!g54) & (g71) & (g723) & (!sk[35]) & (g1412)) + ((g2) & (g54) & (!g71) & (!g723) & (!sk[35]) & (!g1412)) + ((g2) & (g54) & (!g71) & (!g723) & (!sk[35]) & (g1412)) + ((g2) & (g54) & (!g71) & (g723) & (!sk[35]) & (!g1412)) + ((g2) & (g54) & (!g71) & (g723) & (!sk[35]) & (g1412)) + ((g2) & (g54) & (g71) & (!g723) & (!sk[35]) & (!g1412)) + ((g2) & (g54) & (g71) & (!g723) & (!sk[35]) & (g1412)) + ((g2) & (g54) & (g71) & (!g723) & (sk[35]) & (g1412)) + ((g2) & (g54) & (g71) & (g723) & (!sk[35]) & (!g1412)) + ((g2) & (g54) & (g71) & (g723) & (!sk[35]) & (g1412)) + ((g2) & (g54) & (g71) & (g723) & (sk[35]) & (!g1412)) + ((g2) & (g54) & (g71) & (g723) & (sk[35]) & (g1412)));
	assign g1414 = (((!g102) & (!g350) & (!g608) & (!g898) & (sk[36]) & (!g1413)) + ((!g102) & (!g350) & (!g608) & (g898) & (sk[36]) & (!g1413)) + ((!g102) & (!g350) & (g608) & (!g898) & (!sk[36]) & (g1413)) + ((!g102) & (!g350) & (g608) & (!g898) & (sk[36]) & (!g1413)) + ((!g102) & (!g350) & (g608) & (g898) & (!sk[36]) & (!g1413)) + ((!g102) & (!g350) & (g608) & (g898) & (!sk[36]) & (g1413)) + ((!g102) & (!g350) & (g608) & (g898) & (sk[36]) & (!g1413)) + ((!g102) & (g350) & (!g608) & (!g898) & (!sk[36]) & (!g1413)) + ((!g102) & (g350) & (!g608) & (!g898) & (!sk[36]) & (g1413)) + ((!g102) & (g350) & (!g608) & (g898) & (!sk[36]) & (!g1413)) + ((!g102) & (g350) & (!g608) & (g898) & (!sk[36]) & (g1413)) + ((!g102) & (g350) & (g608) & (!g898) & (!sk[36]) & (!g1413)) + ((!g102) & (g350) & (g608) & (!g898) & (!sk[36]) & (g1413)) + ((!g102) & (g350) & (g608) & (g898) & (!sk[36]) & (!g1413)) + ((!g102) & (g350) & (g608) & (g898) & (!sk[36]) & (g1413)) + ((!g102) & (g350) & (g608) & (g898) & (sk[36]) & (!g1413)) + ((g102) & (!g350) & (g608) & (!g898) & (!sk[36]) & (g1413)) + ((g102) & (!g350) & (g608) & (g898) & (!sk[36]) & (!g1413)) + ((g102) & (!g350) & (g608) & (g898) & (!sk[36]) & (g1413)) + ((g102) & (!g350) & (g608) & (g898) & (sk[36]) & (!g1413)) + ((g102) & (g350) & (!g608) & (!g898) & (!sk[36]) & (!g1413)) + ((g102) & (g350) & (!g608) & (!g898) & (!sk[36]) & (g1413)) + ((g102) & (g350) & (!g608) & (g898) & (!sk[36]) & (!g1413)) + ((g102) & (g350) & (!g608) & (g898) & (!sk[36]) & (g1413)) + ((g102) & (g350) & (g608) & (!g898) & (!sk[36]) & (!g1413)) + ((g102) & (g350) & (g608) & (!g898) & (!sk[36]) & (g1413)) + ((g102) & (g350) & (g608) & (g898) & (!sk[36]) & (!g1413)) + ((g102) & (g350) & (g608) & (g898) & (!sk[36]) & (g1413)) + ((g102) & (g350) & (g608) & (g898) & (sk[36]) & (!g1413)));
	assign g1415 = (((!g774) & (!g1408) & (!g1409) & (sk[37]) & (g1411) & (g1414)) + ((!g774) & (!g1408) & (g1409) & (!sk[37]) & (!g1411) & (g1414)) + ((!g774) & (!g1408) & (g1409) & (!sk[37]) & (g1411) & (!g1414)) + ((!g774) & (!g1408) & (g1409) & (!sk[37]) & (g1411) & (g1414)) + ((!g774) & (g1408) & (!g1409) & (!sk[37]) & (!g1411) & (!g1414)) + ((!g774) & (g1408) & (!g1409) & (!sk[37]) & (!g1411) & (g1414)) + ((!g774) & (g1408) & (!g1409) & (!sk[37]) & (g1411) & (!g1414)) + ((!g774) & (g1408) & (!g1409) & (!sk[37]) & (g1411) & (g1414)) + ((!g774) & (g1408) & (g1409) & (!sk[37]) & (!g1411) & (!g1414)) + ((!g774) & (g1408) & (g1409) & (!sk[37]) & (!g1411) & (g1414)) + ((!g774) & (g1408) & (g1409) & (!sk[37]) & (g1411) & (!g1414)) + ((!g774) & (g1408) & (g1409) & (!sk[37]) & (g1411) & (g1414)) + ((g774) & (!g1408) & (g1409) & (!sk[37]) & (!g1411) & (g1414)) + ((g774) & (!g1408) & (g1409) & (!sk[37]) & (g1411) & (!g1414)) + ((g774) & (!g1408) & (g1409) & (!sk[37]) & (g1411) & (g1414)) + ((g774) & (g1408) & (!g1409) & (!sk[37]) & (!g1411) & (!g1414)) + ((g774) & (g1408) & (!g1409) & (!sk[37]) & (!g1411) & (g1414)) + ((g774) & (g1408) & (!g1409) & (!sk[37]) & (g1411) & (!g1414)) + ((g774) & (g1408) & (!g1409) & (!sk[37]) & (g1411) & (g1414)) + ((g774) & (g1408) & (g1409) & (!sk[37]) & (!g1411) & (!g1414)) + ((g774) & (g1408) & (g1409) & (!sk[37]) & (!g1411) & (g1414)) + ((g774) & (g1408) & (g1409) & (!sk[37]) & (g1411) & (!g1414)) + ((g774) & (g1408) & (g1409) & (!sk[37]) & (g1411) & (g1414)));
	assign g1416 = (((!sk[38]) & (!g1460) & (!g1004) & (g1395) & (!g1407) & (g1415)) + ((!sk[38]) & (!g1460) & (!g1004) & (g1395) & (g1407) & (!g1415)) + ((!sk[38]) & (!g1460) & (!g1004) & (g1395) & (g1407) & (g1415)) + ((!sk[38]) & (!g1460) & (g1004) & (!g1395) & (!g1407) & (!g1415)) + ((!sk[38]) & (!g1460) & (g1004) & (!g1395) & (!g1407) & (g1415)) + ((!sk[38]) & (!g1460) & (g1004) & (!g1395) & (g1407) & (!g1415)) + ((!sk[38]) & (!g1460) & (g1004) & (!g1395) & (g1407) & (g1415)) + ((!sk[38]) & (!g1460) & (g1004) & (g1395) & (!g1407) & (!g1415)) + ((!sk[38]) & (!g1460) & (g1004) & (g1395) & (!g1407) & (g1415)) + ((!sk[38]) & (!g1460) & (g1004) & (g1395) & (g1407) & (!g1415)) + ((!sk[38]) & (!g1460) & (g1004) & (g1395) & (g1407) & (g1415)) + ((!sk[38]) & (g1460) & (!g1004) & (g1395) & (!g1407) & (g1415)) + ((!sk[38]) & (g1460) & (!g1004) & (g1395) & (g1407) & (!g1415)) + ((!sk[38]) & (g1460) & (!g1004) & (g1395) & (g1407) & (g1415)) + ((!sk[38]) & (g1460) & (g1004) & (!g1395) & (!g1407) & (!g1415)) + ((!sk[38]) & (g1460) & (g1004) & (!g1395) & (!g1407) & (g1415)) + ((!sk[38]) & (g1460) & (g1004) & (!g1395) & (g1407) & (!g1415)) + ((!sk[38]) & (g1460) & (g1004) & (!g1395) & (g1407) & (g1415)) + ((!sk[38]) & (g1460) & (g1004) & (g1395) & (!g1407) & (!g1415)) + ((!sk[38]) & (g1460) & (g1004) & (g1395) & (!g1407) & (g1415)) + ((!sk[38]) & (g1460) & (g1004) & (g1395) & (g1407) & (!g1415)) + ((!sk[38]) & (g1460) & (g1004) & (g1395) & (g1407) & (g1415)) + ((sk[38]) & (g1460) & (!g1004) & (g1395) & (g1407) & (g1415)));
	assign g1417 = (((!g1152) & (!g1183) & (g1295) & (!g1368) & (!sk[39]) & (g1416)) + ((!g1152) & (!g1183) & (g1295) & (g1368) & (!sk[39]) & (!g1416)) + ((!g1152) & (!g1183) & (g1295) & (g1368) & (!sk[39]) & (g1416)) + ((!g1152) & (g1183) & (!g1295) & (!g1368) & (!sk[39]) & (!g1416)) + ((!g1152) & (g1183) & (!g1295) & (!g1368) & (!sk[39]) & (g1416)) + ((!g1152) & (g1183) & (!g1295) & (g1368) & (!sk[39]) & (!g1416)) + ((!g1152) & (g1183) & (!g1295) & (g1368) & (!sk[39]) & (g1416)) + ((!g1152) & (g1183) & (g1295) & (!g1368) & (!sk[39]) & (!g1416)) + ((!g1152) & (g1183) & (g1295) & (!g1368) & (!sk[39]) & (g1416)) + ((!g1152) & (g1183) & (g1295) & (g1368) & (!sk[39]) & (!g1416)) + ((!g1152) & (g1183) & (g1295) & (g1368) & (!sk[39]) & (g1416)) + ((g1152) & (!g1183) & (g1295) & (!g1368) & (!sk[39]) & (g1416)) + ((g1152) & (!g1183) & (g1295) & (g1368) & (!sk[39]) & (!g1416)) + ((g1152) & (!g1183) & (g1295) & (g1368) & (!sk[39]) & (g1416)) + ((g1152) & (g1183) & (!g1295) & (!g1368) & (!sk[39]) & (!g1416)) + ((g1152) & (g1183) & (!g1295) & (!g1368) & (!sk[39]) & (g1416)) + ((g1152) & (g1183) & (!g1295) & (g1368) & (!sk[39]) & (!g1416)) + ((g1152) & (g1183) & (!g1295) & (g1368) & (!sk[39]) & (g1416)) + ((g1152) & (g1183) & (g1295) & (!g1368) & (!sk[39]) & (!g1416)) + ((g1152) & (g1183) & (g1295) & (!g1368) & (!sk[39]) & (g1416)) + ((g1152) & (g1183) & (g1295) & (g1368) & (!sk[39]) & (!g1416)) + ((g1152) & (g1183) & (g1295) & (g1368) & (!sk[39]) & (g1416)) + ((g1152) & (g1183) & (g1295) & (g1368) & (sk[39]) & (g1416)));
	assign g1418 = (((!g109) & (!g161) & (!g392) & (!g569) & (!g1149) & (g374)) + ((!g109) & (!g161) & (!g392) & (!g569) & (g1149) & (g374)) + ((!g109) & (!g161) & (g392) & (!g569) & (g1149) & (g374)) + ((!g109) & (g161) & (!g392) & (!g569) & (!g1149) & (g374)) + ((!g109) & (g161) & (!g392) & (!g569) & (g1149) & (g374)) + ((!g109) & (g161) & (g392) & (!g569) & (g1149) & (g374)) + ((g109) & (!g161) & (!g392) & (!g569) & (!g1149) & (g374)) + ((g109) & (!g161) & (!g392) & (!g569) & (g1149) & (g374)) + ((g109) & (!g161) & (g392) & (!g569) & (g1149) & (g374)));
	assign g1419 = (((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g429) & (!g445)) + ((!i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g429) & (g445)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (!g429) & (g445)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g429) & (!g445)) + ((!i_15_) & (i_12_) & (i_13_) & (i_14_) & (g429) & (g445)) + ((i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (!g429) & (g445)) + ((i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g429) & (!g445)) + ((i_15_) & (!i_12_) & (!i_13_) & (i_14_) & (g429) & (g445)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (!g429) & (g445)) + ((i_15_) & (!i_12_) & (i_13_) & (i_14_) & (g429) & (g445)) + ((i_15_) & (i_12_) & (!i_13_) & (i_14_) & (!g429) & (g445)) + ((i_15_) & (i_12_) & (!i_13_) & (i_14_) & (g429) & (g445)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (!g429) & (g445)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g429) & (!g445)) + ((i_15_) & (i_12_) & (i_13_) & (!i_14_) & (g429) & (g445)) + ((i_15_) & (i_12_) & (i_13_) & (i_14_) & (g429) & (!g445)) + ((i_15_) & (i_12_) & (i_13_) & (i_14_) & (g429) & (g445)));
	assign g1420 = (((!g24) & (!g35) & (!g36) & (sk[42]) & (!g68)) + ((!g24) & (!g35) & (!g36) & (sk[42]) & (g68)) + ((!g24) & (!g35) & (g36) & (!sk[42]) & (!g68)) + ((!g24) & (!g35) & (g36) & (!sk[42]) & (g68)) + ((!g24) & (!g35) & (g36) & (sk[42]) & (g68)) + ((!g24) & (g35) & (g36) & (!sk[42]) & (!g68)) + ((!g24) & (g35) & (g36) & (!sk[42]) & (g68)) + ((g24) & (!g35) & (!g36) & (sk[42]) & (!g68)) + ((g24) & (!g35) & (!g36) & (sk[42]) & (g68)) + ((g24) & (!g35) & (g36) & (!sk[42]) & (!g68)) + ((g24) & (!g35) & (g36) & (!sk[42]) & (g68)) + ((g24) & (!g35) & (g36) & (sk[42]) & (g68)) + ((g24) & (g35) & (!g36) & (sk[42]) & (g68)) + ((g24) & (g35) & (g36) & (!sk[42]) & (!g68)) + ((g24) & (g35) & (g36) & (!sk[42]) & (g68)) + ((g24) & (g35) & (g36) & (sk[42]) & (g68)));
	assign g1421 = (((!g157) & (!g343) & (!sk[43]) & (g502) & (!g1419) & (g1420)) + ((!g157) & (!g343) & (!sk[43]) & (g502) & (g1419) & (!g1420)) + ((!g157) & (!g343) & (!sk[43]) & (g502) & (g1419) & (g1420)) + ((!g157) & (!g343) & (sk[43]) & (!g502) & (!g1419) & (!g1420)) + ((!g157) & (!g343) & (sk[43]) & (!g502) & (!g1419) & (g1420)) + ((!g157) & (!g343) & (sk[43]) & (!g502) & (g1419) & (!g1420)) + ((!g157) & (!g343) & (sk[43]) & (!g502) & (g1419) & (g1420)) + ((!g157) & (g343) & (!sk[43]) & (!g502) & (!g1419) & (!g1420)) + ((!g157) & (g343) & (!sk[43]) & (!g502) & (!g1419) & (g1420)) + ((!g157) & (g343) & (!sk[43]) & (!g502) & (g1419) & (!g1420)) + ((!g157) & (g343) & (!sk[43]) & (!g502) & (g1419) & (g1420)) + ((!g157) & (g343) & (!sk[43]) & (g502) & (!g1419) & (!g1420)) + ((!g157) & (g343) & (!sk[43]) & (g502) & (!g1419) & (g1420)) + ((!g157) & (g343) & (!sk[43]) & (g502) & (g1419) & (!g1420)) + ((!g157) & (g343) & (!sk[43]) & (g502) & (g1419) & (g1420)) + ((!g157) & (g343) & (sk[43]) & (!g502) & (!g1419) & (!g1420)) + ((!g157) & (g343) & (sk[43]) & (!g502) & (!g1419) & (g1420)) + ((!g157) & (g343) & (sk[43]) & (!g502) & (g1419) & (!g1420)) + ((!g157) & (g343) & (sk[43]) & (!g502) & (g1419) & (g1420)) + ((g157) & (!g343) & (!sk[43]) & (g502) & (!g1419) & (g1420)) + ((g157) & (!g343) & (!sk[43]) & (g502) & (g1419) & (!g1420)) + ((g157) & (!g343) & (!sk[43]) & (g502) & (g1419) & (g1420)) + ((g157) & (g343) & (!sk[43]) & (!g502) & (!g1419) & (!g1420)) + ((g157) & (g343) & (!sk[43]) & (!g502) & (!g1419) & (g1420)) + ((g157) & (g343) & (!sk[43]) & (!g502) & (g1419) & (!g1420)) + ((g157) & (g343) & (!sk[43]) & (!g502) & (g1419) & (g1420)) + ((g157) & (g343) & (!sk[43]) & (g502) & (!g1419) & (!g1420)) + ((g157) & (g343) & (!sk[43]) & (g502) & (!g1419) & (g1420)) + ((g157) & (g343) & (!sk[43]) & (g502) & (g1419) & (!g1420)) + ((g157) & (g343) & (!sk[43]) & (g502) & (g1419) & (g1420)) + ((g157) & (g343) & (sk[43]) & (!g502) & (!g1419) & (g1420)));
	assign g1422 = (((!g250) & (!g454) & (g1179) & (!sk[44]) & (!g1418) & (g1421)) + ((!g250) & (!g454) & (g1179) & (!sk[44]) & (g1418) & (!g1421)) + ((!g250) & (!g454) & (g1179) & (!sk[44]) & (g1418) & (g1421)) + ((!g250) & (g454) & (!g1179) & (!sk[44]) & (!g1418) & (!g1421)) + ((!g250) & (g454) & (!g1179) & (!sk[44]) & (!g1418) & (g1421)) + ((!g250) & (g454) & (!g1179) & (!sk[44]) & (g1418) & (!g1421)) + ((!g250) & (g454) & (!g1179) & (!sk[44]) & (g1418) & (g1421)) + ((!g250) & (g454) & (g1179) & (!sk[44]) & (!g1418) & (!g1421)) + ((!g250) & (g454) & (g1179) & (!sk[44]) & (!g1418) & (g1421)) + ((!g250) & (g454) & (g1179) & (!sk[44]) & (g1418) & (!g1421)) + ((!g250) & (g454) & (g1179) & (!sk[44]) & (g1418) & (g1421)) + ((g250) & (!g454) & (g1179) & (!sk[44]) & (!g1418) & (g1421)) + ((g250) & (!g454) & (g1179) & (!sk[44]) & (g1418) & (!g1421)) + ((g250) & (!g454) & (g1179) & (!sk[44]) & (g1418) & (g1421)) + ((g250) & (g454) & (!g1179) & (!sk[44]) & (!g1418) & (!g1421)) + ((g250) & (g454) & (!g1179) & (!sk[44]) & (!g1418) & (g1421)) + ((g250) & (g454) & (!g1179) & (!sk[44]) & (g1418) & (!g1421)) + ((g250) & (g454) & (!g1179) & (!sk[44]) & (g1418) & (g1421)) + ((g250) & (g454) & (!g1179) & (sk[44]) & (g1418) & (g1421)) + ((g250) & (g454) & (g1179) & (!sk[44]) & (!g1418) & (!g1421)) + ((g250) & (g454) & (g1179) & (!sk[44]) & (!g1418) & (g1421)) + ((g250) & (g454) & (g1179) & (!sk[44]) & (g1418) & (!g1421)) + ((g250) & (g454) & (g1179) & (!sk[44]) & (g1418) & (g1421)));
	assign g1423 = (((!g5) & (!sk[45]) & (!g16) & (g30) & (!g49)) + ((!g5) & (!sk[45]) & (!g16) & (g30) & (g49)) + ((!g5) & (!sk[45]) & (g16) & (g30) & (!g49)) + ((!g5) & (!sk[45]) & (g16) & (g30) & (g49)) + ((g5) & (!sk[45]) & (!g16) & (g30) & (!g49)) + ((g5) & (!sk[45]) & (!g16) & (g30) & (g49)) + ((g5) & (!sk[45]) & (g16) & (g30) & (!g49)) + ((g5) & (!sk[45]) & (g16) & (g30) & (g49)) + ((g5) & (sk[45]) & (g16) & (!g30) & (g49)) + ((g5) & (sk[45]) & (g16) & (g30) & (!g49)) + ((g5) & (sk[45]) & (g16) & (g30) & (g49)));
	assign g1424 = (((!sk[46]) & (!g2) & (!g14) & (g62) & (!g1126) & (g1423)) + ((!sk[46]) & (!g2) & (!g14) & (g62) & (g1126) & (!g1423)) + ((!sk[46]) & (!g2) & (!g14) & (g62) & (g1126) & (g1423)) + ((!sk[46]) & (!g2) & (g14) & (!g62) & (!g1126) & (!g1423)) + ((!sk[46]) & (!g2) & (g14) & (!g62) & (!g1126) & (g1423)) + ((!sk[46]) & (!g2) & (g14) & (!g62) & (g1126) & (!g1423)) + ((!sk[46]) & (!g2) & (g14) & (!g62) & (g1126) & (g1423)) + ((!sk[46]) & (!g2) & (g14) & (g62) & (!g1126) & (!g1423)) + ((!sk[46]) & (!g2) & (g14) & (g62) & (!g1126) & (g1423)) + ((!sk[46]) & (!g2) & (g14) & (g62) & (g1126) & (!g1423)) + ((!sk[46]) & (!g2) & (g14) & (g62) & (g1126) & (g1423)) + ((!sk[46]) & (g2) & (!g14) & (g62) & (!g1126) & (g1423)) + ((!sk[46]) & (g2) & (!g14) & (g62) & (g1126) & (!g1423)) + ((!sk[46]) & (g2) & (!g14) & (g62) & (g1126) & (g1423)) + ((!sk[46]) & (g2) & (g14) & (!g62) & (!g1126) & (!g1423)) + ((!sk[46]) & (g2) & (g14) & (!g62) & (!g1126) & (g1423)) + ((!sk[46]) & (g2) & (g14) & (!g62) & (g1126) & (!g1423)) + ((!sk[46]) & (g2) & (g14) & (!g62) & (g1126) & (g1423)) + ((!sk[46]) & (g2) & (g14) & (g62) & (!g1126) & (!g1423)) + ((!sk[46]) & (g2) & (g14) & (g62) & (!g1126) & (g1423)) + ((!sk[46]) & (g2) & (g14) & (g62) & (g1126) & (!g1423)) + ((!sk[46]) & (g2) & (g14) & (g62) & (g1126) & (g1423)) + ((sk[46]) & (!g2) & (!g14) & (!g62) & (!g1126) & (!g1423)) + ((sk[46]) & (!g2) & (!g14) & (!g62) & (g1126) & (!g1423)) + ((sk[46]) & (!g2) & (!g14) & (g62) & (!g1126) & (!g1423)) + ((sk[46]) & (!g2) & (!g14) & (g62) & (g1126) & (!g1423)) + ((sk[46]) & (!g2) & (g14) & (!g62) & (!g1126) & (!g1423)) + ((sk[46]) & (!g2) & (g14) & (!g62) & (g1126) & (!g1423)) + ((sk[46]) & (!g2) & (g14) & (g62) & (!g1126) & (!g1423)) + ((sk[46]) & (!g2) & (g14) & (g62) & (g1126) & (!g1423)) + ((sk[46]) & (g2) & (!g14) & (!g62) & (!g1126) & (!g1423)) + ((sk[46]) & (g2) & (!g14) & (!g62) & (g1126) & (!g1423)) + ((sk[46]) & (g2) & (!g14) & (g62) & (!g1126) & (!g1423)) + ((sk[46]) & (g2) & (!g14) & (g62) & (g1126) & (!g1423)) + ((sk[46]) & (g2) & (g14) & (!g62) & (!g1126) & (!g1423)) + ((sk[46]) & (g2) & (g14) & (!g62) & (g1126) & (!g1423)) + ((sk[46]) & (g2) & (g14) & (g62) & (g1126) & (!g1423)));
	assign o_41_ = (((!g80) & (!sk[47]) & (!i_11_) & (g7) & (!g101)) + ((!g80) & (!sk[47]) & (!i_11_) & (g7) & (g101)) + ((!g80) & (!sk[47]) & (i_11_) & (g7) & (!g101)) + ((!g80) & (!sk[47]) & (i_11_) & (g7) & (g101)) + ((g80) & (!sk[47]) & (!i_11_) & (g7) & (!g101)) + ((g80) & (!sk[47]) & (!i_11_) & (g7) & (g101)) + ((g80) & (!sk[47]) & (i_11_) & (g7) & (!g101)) + ((g80) & (!sk[47]) & (i_11_) & (g7) & (g101)) + ((g80) & (sk[47]) & (!i_11_) & (g7) & (g101)));
	assign g1426 = (((!g395) & (sk[48]) & (!g1459)) + ((g395) & (!sk[48]) & (!g1459)) + ((g395) & (!sk[48]) & (g1459)));
	assign g1427 = (((!sk[49]) & (g774) & (!g779)) + ((!sk[49]) & (g774) & (g779)) + ((sk[49]) & (!g774) & (g779)));
	assign g1428 = (((!g135) & (!g299) & (!g342) & (!g681) & (g301) & (g302)) + ((g135) & (!g299) & (!g342) & (!g681) & (g301) & (g302)) + ((g135) & (!g299) & (g342) & (!g681) & (g301) & (g302)));
	assign g1429 = (((!g122) & (!g948) & (!sk[51]) & (g1184) & (!g1268)) + ((!g122) & (!g948) & (!sk[51]) & (g1184) & (g1268)) + ((!g122) & (!g948) & (sk[51]) & (!g1184) & (!g1268)) + ((!g122) & (g948) & (!sk[51]) & (g1184) & (!g1268)) + ((!g122) & (g948) & (!sk[51]) & (g1184) & (g1268)) + ((!g122) & (g948) & (sk[51]) & (!g1184) & (!g1268)) + ((g122) & (!g948) & (!sk[51]) & (g1184) & (!g1268)) + ((g122) & (!g948) & (!sk[51]) & (g1184) & (g1268)) + ((g122) & (g948) & (!sk[51]) & (g1184) & (!g1268)) + ((g122) & (g948) & (!sk[51]) & (g1184) & (g1268)) + ((g122) & (g948) & (sk[51]) & (!g1184) & (!g1268)));
	assign g1430 = (((g122) & (!sk[52]) & (!g898)) + ((g122) & (!sk[52]) & (g898)) + ((g122) & (sk[52]) & (!g898)));
	assign g1431 = (((!g221) & (!g222) & (!g1430) & (g223) & (g224) & (!g1178)));
	assign g1432 = (((!g637) & (g138) & (g1554) & (g862) & (g1429) & (g1431)));
	assign g1433 = (((!i_8_) & (!g333) & (!sk[55]) & (g898) & (!g1015) & (g1032)) + ((!i_8_) & (!g333) & (!sk[55]) & (g898) & (g1015) & (!g1032)) + ((!i_8_) & (!g333) & (!sk[55]) & (g898) & (g1015) & (g1032)) + ((!i_8_) & (!g333) & (sk[55]) & (!g898) & (!g1015) & (!g1032)) + ((!i_8_) & (!g333) & (sk[55]) & (!g898) & (!g1015) & (g1032)) + ((!i_8_) & (!g333) & (sk[55]) & (!g898) & (g1015) & (!g1032)) + ((!i_8_) & (!g333) & (sk[55]) & (!g898) & (g1015) & (g1032)) + ((!i_8_) & (!g333) & (sk[55]) & (g898) & (!g1015) & (!g1032)) + ((!i_8_) & (!g333) & (sk[55]) & (g898) & (!g1015) & (g1032)) + ((!i_8_) & (!g333) & (sk[55]) & (g898) & (g1015) & (!g1032)) + ((!i_8_) & (g333) & (!sk[55]) & (!g898) & (!g1015) & (!g1032)) + ((!i_8_) & (g333) & (!sk[55]) & (!g898) & (!g1015) & (g1032)) + ((!i_8_) & (g333) & (!sk[55]) & (!g898) & (g1015) & (!g1032)) + ((!i_8_) & (g333) & (!sk[55]) & (!g898) & (g1015) & (g1032)) + ((!i_8_) & (g333) & (!sk[55]) & (g898) & (!g1015) & (!g1032)) + ((!i_8_) & (g333) & (!sk[55]) & (g898) & (!g1015) & (g1032)) + ((!i_8_) & (g333) & (!sk[55]) & (g898) & (g1015) & (!g1032)) + ((!i_8_) & (g333) & (!sk[55]) & (g898) & (g1015) & (g1032)) + ((!i_8_) & (g333) & (sk[55]) & (!g898) & (!g1015) & (!g1032)) + ((!i_8_) & (g333) & (sk[55]) & (!g898) & (!g1015) & (g1032)) + ((!i_8_) & (g333) & (sk[55]) & (!g898) & (g1015) & (!g1032)) + ((!i_8_) & (g333) & (sk[55]) & (!g898) & (g1015) & (g1032)) + ((!i_8_) & (g333) & (sk[55]) & (g898) & (!g1015) & (!g1032)) + ((!i_8_) & (g333) & (sk[55]) & (g898) & (!g1015) & (g1032)) + ((!i_8_) & (g333) & (sk[55]) & (g898) & (g1015) & (!g1032)) + ((!i_8_) & (g333) & (sk[55]) & (g898) & (g1015) & (g1032)) + ((i_8_) & (!g333) & (!sk[55]) & (g898) & (!g1015) & (g1032)) + ((i_8_) & (!g333) & (!sk[55]) & (g898) & (g1015) & (!g1032)) + ((i_8_) & (!g333) & (!sk[55]) & (g898) & (g1015) & (g1032)) + ((i_8_) & (g333) & (!sk[55]) & (!g898) & (!g1015) & (!g1032)) + ((i_8_) & (g333) & (!sk[55]) & (!g898) & (!g1015) & (g1032)) + ((i_8_) & (g333) & (!sk[55]) & (!g898) & (g1015) & (!g1032)) + ((i_8_) & (g333) & (!sk[55]) & (!g898) & (g1015) & (g1032)) + ((i_8_) & (g333) & (!sk[55]) & (g898) & (!g1015) & (!g1032)) + ((i_8_) & (g333) & (!sk[55]) & (g898) & (!g1015) & (g1032)) + ((i_8_) & (g333) & (!sk[55]) & (g898) & (g1015) & (!g1032)) + ((i_8_) & (g333) & (!sk[55]) & (g898) & (g1015) & (g1032)));
	assign g1434 = (((!sk[56]) & (!g514) & (!g725) & (g641) & (!g1203)) + ((!sk[56]) & (!g514) & (!g725) & (g641) & (g1203)) + ((!sk[56]) & (!g514) & (g725) & (g641) & (!g1203)) + ((!sk[56]) & (!g514) & (g725) & (g641) & (g1203)) + ((!sk[56]) & (g514) & (!g725) & (g641) & (!g1203)) + ((!sk[56]) & (g514) & (!g725) & (g641) & (g1203)) + ((!sk[56]) & (g514) & (g725) & (g641) & (!g1203)) + ((!sk[56]) & (g514) & (g725) & (g641) & (g1203)) + ((sk[56]) & (!g514) & (g725) & (!g641) & (g1203)));
	assign g1435 = (((!g165) & (!g933) & (!g1433) & (!g1434) & (!g1362) & (g1365)) + ((!g165) & (!g933) & (!g1433) & (g1434) & (!g1362) & (g1365)) + ((!g165) & (!g933) & (g1433) & (!g1434) & (!g1362) & (g1365)) + ((!g165) & (!g933) & (g1433) & (g1434) & (!g1362) & (g1365)) + ((!g165) & (g933) & (!g1433) & (!g1434) & (!g1362) & (g1365)) + ((!g165) & (g933) & (!g1433) & (g1434) & (!g1362) & (g1365)) + ((!g165) & (g933) & (g1433) & (!g1434) & (!g1362) & (g1365)) + ((!g165) & (g933) & (g1433) & (g1434) & (!g1362) & (g1365)) + ((g165) & (g933) & (!g1433) & (g1434) & (!g1362) & (g1365)));
	assign g1436 = (((g1427) & (g787) & (g1370) & (g1428) & (g1432) & (g1435)));
	assign g1437 = (((!g135) & (!sk[59]) & (!g337) & (g635) & (!g1001) & (g1436)) + ((!g135) & (!sk[59]) & (!g337) & (g635) & (g1001) & (!g1436)) + ((!g135) & (!sk[59]) & (!g337) & (g635) & (g1001) & (g1436)) + ((!g135) & (!sk[59]) & (g337) & (!g635) & (!g1001) & (!g1436)) + ((!g135) & (!sk[59]) & (g337) & (!g635) & (!g1001) & (g1436)) + ((!g135) & (!sk[59]) & (g337) & (!g635) & (g1001) & (!g1436)) + ((!g135) & (!sk[59]) & (g337) & (!g635) & (g1001) & (g1436)) + ((!g135) & (!sk[59]) & (g337) & (g635) & (!g1001) & (!g1436)) + ((!g135) & (!sk[59]) & (g337) & (g635) & (!g1001) & (g1436)) + ((!g135) & (!sk[59]) & (g337) & (g635) & (g1001) & (!g1436)) + ((!g135) & (!sk[59]) & (g337) & (g635) & (g1001) & (g1436)) + ((!g135) & (sk[59]) & (!g337) & (!g635) & (g1001) & (g1436)) + ((g135) & (!sk[59]) & (!g337) & (g635) & (!g1001) & (g1436)) + ((g135) & (!sk[59]) & (!g337) & (g635) & (g1001) & (!g1436)) + ((g135) & (!sk[59]) & (!g337) & (g635) & (g1001) & (g1436)) + ((g135) & (!sk[59]) & (g337) & (!g635) & (!g1001) & (!g1436)) + ((g135) & (!sk[59]) & (g337) & (!g635) & (!g1001) & (g1436)) + ((g135) & (!sk[59]) & (g337) & (!g635) & (g1001) & (!g1436)) + ((g135) & (!sk[59]) & (g337) & (!g635) & (g1001) & (g1436)) + ((g135) & (!sk[59]) & (g337) & (g635) & (!g1001) & (!g1436)) + ((g135) & (!sk[59]) & (g337) & (g635) & (!g1001) & (g1436)) + ((g135) & (!sk[59]) & (g337) & (g635) & (g1001) & (!g1436)) + ((g135) & (!sk[59]) & (g337) & (g635) & (g1001) & (g1436)) + ((g135) & (sk[59]) & (!g337) & (!g635) & (g1001) & (g1436)) + ((g135) & (sk[59]) & (!g337) & (g635) & (g1001) & (g1436)) + ((g135) & (sk[59]) & (g337) & (!g635) & (g1001) & (g1436)) + ((g135) & (sk[59]) & (g337) & (g635) & (g1001) & (g1436)));
	assign g1438 = (((!sk[60]) & (!g17) & (!g23) & (g507) & (!g624) & (g1036)) + ((!sk[60]) & (!g17) & (!g23) & (g507) & (g624) & (!g1036)) + ((!sk[60]) & (!g17) & (!g23) & (g507) & (g624) & (g1036)) + ((!sk[60]) & (!g17) & (g23) & (!g507) & (!g624) & (!g1036)) + ((!sk[60]) & (!g17) & (g23) & (!g507) & (!g624) & (g1036)) + ((!sk[60]) & (!g17) & (g23) & (!g507) & (g624) & (!g1036)) + ((!sk[60]) & (!g17) & (g23) & (!g507) & (g624) & (g1036)) + ((!sk[60]) & (!g17) & (g23) & (g507) & (!g624) & (!g1036)) + ((!sk[60]) & (!g17) & (g23) & (g507) & (!g624) & (g1036)) + ((!sk[60]) & (!g17) & (g23) & (g507) & (g624) & (!g1036)) + ((!sk[60]) & (!g17) & (g23) & (g507) & (g624) & (g1036)) + ((!sk[60]) & (g17) & (!g23) & (g507) & (!g624) & (g1036)) + ((!sk[60]) & (g17) & (!g23) & (g507) & (g624) & (!g1036)) + ((!sk[60]) & (g17) & (!g23) & (g507) & (g624) & (g1036)) + ((!sk[60]) & (g17) & (g23) & (!g507) & (!g624) & (!g1036)) + ((!sk[60]) & (g17) & (g23) & (!g507) & (!g624) & (g1036)) + ((!sk[60]) & (g17) & (g23) & (!g507) & (g624) & (!g1036)) + ((!sk[60]) & (g17) & (g23) & (!g507) & (g624) & (g1036)) + ((!sk[60]) & (g17) & (g23) & (g507) & (!g624) & (!g1036)) + ((!sk[60]) & (g17) & (g23) & (g507) & (!g624) & (g1036)) + ((!sk[60]) & (g17) & (g23) & (g507) & (g624) & (!g1036)) + ((!sk[60]) & (g17) & (g23) & (g507) & (g624) & (g1036)) + ((sk[60]) & (!g17) & (g23) & (!g507) & (g624) & (g1036)) + ((sk[60]) & (!g17) & (g23) & (g507) & (g624) & (g1036)) + ((sk[60]) & (g17) & (g23) & (!g507) & (g624) & (g1036)));
	assign g1439 = (((!g408) & (!g605) & (!sk[61]) & (g971) & (!g1248) & (g1181)) + ((!g408) & (!g605) & (!sk[61]) & (g971) & (g1248) & (!g1181)) + ((!g408) & (!g605) & (!sk[61]) & (g971) & (g1248) & (g1181)) + ((!g408) & (!g605) & (sk[61]) & (g971) & (!g1248) & (!g1181)) + ((!g408) & (g605) & (!sk[61]) & (!g971) & (!g1248) & (!g1181)) + ((!g408) & (g605) & (!sk[61]) & (!g971) & (!g1248) & (g1181)) + ((!g408) & (g605) & (!sk[61]) & (!g971) & (g1248) & (!g1181)) + ((!g408) & (g605) & (!sk[61]) & (!g971) & (g1248) & (g1181)) + ((!g408) & (g605) & (!sk[61]) & (g971) & (!g1248) & (!g1181)) + ((!g408) & (g605) & (!sk[61]) & (g971) & (!g1248) & (g1181)) + ((!g408) & (g605) & (!sk[61]) & (g971) & (g1248) & (!g1181)) + ((!g408) & (g605) & (!sk[61]) & (g971) & (g1248) & (g1181)) + ((g408) & (!g605) & (!sk[61]) & (g971) & (!g1248) & (g1181)) + ((g408) & (!g605) & (!sk[61]) & (g971) & (g1248) & (!g1181)) + ((g408) & (!g605) & (!sk[61]) & (g971) & (g1248) & (g1181)) + ((g408) & (!g605) & (sk[61]) & (!g971) & (!g1248) & (!g1181)) + ((g408) & (!g605) & (sk[61]) & (!g971) & (g1248) & (!g1181)) + ((g408) & (!g605) & (sk[61]) & (g971) & (!g1248) & (!g1181)) + ((g408) & (!g605) & (sk[61]) & (g971) & (g1248) & (!g1181)) + ((g408) & (g605) & (!sk[61]) & (!g971) & (!g1248) & (!g1181)) + ((g408) & (g605) & (!sk[61]) & (!g971) & (!g1248) & (g1181)) + ((g408) & (g605) & (!sk[61]) & (!g971) & (g1248) & (!g1181)) + ((g408) & (g605) & (!sk[61]) & (!g971) & (g1248) & (g1181)) + ((g408) & (g605) & (!sk[61]) & (g971) & (!g1248) & (!g1181)) + ((g408) & (g605) & (!sk[61]) & (g971) & (!g1248) & (g1181)) + ((g408) & (g605) & (!sk[61]) & (g971) & (g1248) & (!g1181)) + ((g408) & (g605) & (!sk[61]) & (g971) & (g1248) & (g1181)) + ((g408) & (g605) & (sk[61]) & (!g971) & (!g1248) & (!g1181)) + ((g408) & (g605) & (sk[61]) & (!g971) & (g1248) & (!g1181)) + ((g408) & (g605) & (sk[61]) & (g971) & (!g1248) & (!g1181)) + ((g408) & (g605) & (sk[61]) & (g971) & (g1248) & (!g1181)));
	assign g1440 = (((!g130) & (!g965) & (!sk[62]) & (g1438) & (!g1185) & (g1439)) + ((!g130) & (!g965) & (!sk[62]) & (g1438) & (g1185) & (!g1439)) + ((!g130) & (!g965) & (!sk[62]) & (g1438) & (g1185) & (g1439)) + ((!g130) & (g965) & (!sk[62]) & (!g1438) & (!g1185) & (!g1439)) + ((!g130) & (g965) & (!sk[62]) & (!g1438) & (!g1185) & (g1439)) + ((!g130) & (g965) & (!sk[62]) & (!g1438) & (g1185) & (!g1439)) + ((!g130) & (g965) & (!sk[62]) & (!g1438) & (g1185) & (g1439)) + ((!g130) & (g965) & (!sk[62]) & (g1438) & (!g1185) & (!g1439)) + ((!g130) & (g965) & (!sk[62]) & (g1438) & (!g1185) & (g1439)) + ((!g130) & (g965) & (!sk[62]) & (g1438) & (g1185) & (!g1439)) + ((!g130) & (g965) & (!sk[62]) & (g1438) & (g1185) & (g1439)) + ((!g130) & (g965) & (sk[62]) & (g1438) & (!g1185) & (g1439)) + ((g130) & (!g965) & (!sk[62]) & (g1438) & (!g1185) & (g1439)) + ((g130) & (!g965) & (!sk[62]) & (g1438) & (g1185) & (!g1439)) + ((g130) & (!g965) & (!sk[62]) & (g1438) & (g1185) & (g1439)) + ((g130) & (!g965) & (sk[62]) & (!g1438) & (!g1185) & (g1439)) + ((g130) & (!g965) & (sk[62]) & (g1438) & (!g1185) & (g1439)) + ((g130) & (g965) & (!sk[62]) & (!g1438) & (!g1185) & (!g1439)) + ((g130) & (g965) & (!sk[62]) & (!g1438) & (!g1185) & (g1439)) + ((g130) & (g965) & (!sk[62]) & (!g1438) & (g1185) & (!g1439)) + ((g130) & (g965) & (!sk[62]) & (!g1438) & (g1185) & (g1439)) + ((g130) & (g965) & (!sk[62]) & (g1438) & (!g1185) & (!g1439)) + ((g130) & (g965) & (!sk[62]) & (g1438) & (!g1185) & (g1439)) + ((g130) & (g965) & (!sk[62]) & (g1438) & (g1185) & (!g1439)) + ((g130) & (g965) & (!sk[62]) & (g1438) & (g1185) & (g1439)) + ((g130) & (g965) & (sk[62]) & (!g1438) & (!g1185) & (g1439)) + ((g130) & (g965) & (sk[62]) & (g1438) & (!g1185) & (g1439)));
	assign g1441 = (((!g123) & (!g850) & (!sk[63]) & (g1154)) + ((!g123) & (!g850) & (sk[63]) & (!g1154)) + ((!g123) & (g850) & (!sk[63]) & (!g1154)) + ((!g123) & (g850) & (!sk[63]) & (g1154)) + ((g123) & (!g850) & (!sk[63]) & (g1154)) + ((g123) & (!g850) & (sk[63]) & (!g1154)) + ((g123) & (g850) & (!sk[63]) & (!g1154)) + ((g123) & (g850) & (!sk[63]) & (g1154)) + ((g123) & (g850) & (sk[63]) & (!g1154)));
	assign g1442 = (((!sk[64]) & (!g597) & (!g489) & (g624) & (!g629)) + ((!sk[64]) & (!g597) & (!g489) & (g624) & (g629)) + ((!sk[64]) & (!g597) & (g489) & (g624) & (!g629)) + ((!sk[64]) & (!g597) & (g489) & (g624) & (g629)) + ((!sk[64]) & (g597) & (!g489) & (g624) & (!g629)) + ((!sk[64]) & (g597) & (!g489) & (g624) & (g629)) + ((!sk[64]) & (g597) & (g489) & (g624) & (!g629)) + ((!sk[64]) & (g597) & (g489) & (g624) & (g629)) + ((sk[64]) & (!g597) & (!g489) & (g624) & (!g629)));
	assign g1443 = (((!g70) & (!g335) & (!g468) & (!g770) & (sk[65]) & (!g877)) + ((!g70) & (!g335) & (g468) & (!g770) & (!sk[65]) & (g877)) + ((!g70) & (!g335) & (g468) & (g770) & (!sk[65]) & (!g877)) + ((!g70) & (!g335) & (g468) & (g770) & (!sk[65]) & (g877)) + ((!g70) & (g335) & (!g468) & (!g770) & (!sk[65]) & (!g877)) + ((!g70) & (g335) & (!g468) & (!g770) & (!sk[65]) & (g877)) + ((!g70) & (g335) & (!g468) & (g770) & (!sk[65]) & (!g877)) + ((!g70) & (g335) & (!g468) & (g770) & (!sk[65]) & (g877)) + ((!g70) & (g335) & (g468) & (!g770) & (!sk[65]) & (!g877)) + ((!g70) & (g335) & (g468) & (!g770) & (!sk[65]) & (g877)) + ((!g70) & (g335) & (g468) & (g770) & (!sk[65]) & (!g877)) + ((!g70) & (g335) & (g468) & (g770) & (!sk[65]) & (g877)) + ((g70) & (!g335) & (g468) & (!g770) & (!sk[65]) & (g877)) + ((g70) & (!g335) & (g468) & (g770) & (!sk[65]) & (!g877)) + ((g70) & (!g335) & (g468) & (g770) & (!sk[65]) & (g877)) + ((g70) & (g335) & (!g468) & (!g770) & (!sk[65]) & (!g877)) + ((g70) & (g335) & (!g468) & (!g770) & (!sk[65]) & (g877)) + ((g70) & (g335) & (!g468) & (g770) & (!sk[65]) & (!g877)) + ((g70) & (g335) & (!g468) & (g770) & (!sk[65]) & (g877)) + ((g70) & (g335) & (g468) & (!g770) & (!sk[65]) & (!g877)) + ((g70) & (g335) & (g468) & (!g770) & (!sk[65]) & (g877)) + ((g70) & (g335) & (g468) & (g770) & (!sk[65]) & (!g877)) + ((g70) & (g335) & (g468) & (g770) & (!sk[65]) & (g877)));
	assign g1444 = (((!g334) & (!g875) & (g928) & (!sk[66]) & (!g1442) & (g1443)) + ((!g334) & (!g875) & (g928) & (!sk[66]) & (g1442) & (!g1443)) + ((!g334) & (!g875) & (g928) & (!sk[66]) & (g1442) & (g1443)) + ((!g334) & (g875) & (!g928) & (!sk[66]) & (!g1442) & (!g1443)) + ((!g334) & (g875) & (!g928) & (!sk[66]) & (!g1442) & (g1443)) + ((!g334) & (g875) & (!g928) & (!sk[66]) & (g1442) & (!g1443)) + ((!g334) & (g875) & (!g928) & (!sk[66]) & (g1442) & (g1443)) + ((!g334) & (g875) & (g928) & (!sk[66]) & (!g1442) & (!g1443)) + ((!g334) & (g875) & (g928) & (!sk[66]) & (!g1442) & (g1443)) + ((!g334) & (g875) & (g928) & (!sk[66]) & (g1442) & (!g1443)) + ((!g334) & (g875) & (g928) & (!sk[66]) & (g1442) & (g1443)) + ((g334) & (!g875) & (g928) & (!sk[66]) & (!g1442) & (g1443)) + ((g334) & (!g875) & (g928) & (!sk[66]) & (g1442) & (!g1443)) + ((g334) & (!g875) & (g928) & (!sk[66]) & (g1442) & (g1443)) + ((g334) & (!g875) & (g928) & (sk[66]) & (g1442) & (g1443)) + ((g334) & (g875) & (!g928) & (!sk[66]) & (!g1442) & (!g1443)) + ((g334) & (g875) & (!g928) & (!sk[66]) & (!g1442) & (g1443)) + ((g334) & (g875) & (!g928) & (!sk[66]) & (g1442) & (!g1443)) + ((g334) & (g875) & (!g928) & (!sk[66]) & (g1442) & (g1443)) + ((g334) & (g875) & (g928) & (!sk[66]) & (!g1442) & (!g1443)) + ((g334) & (g875) & (g928) & (!sk[66]) & (!g1442) & (g1443)) + ((g334) & (g875) & (g928) & (!sk[66]) & (g1442) & (!g1443)) + ((g334) & (g875) & (g928) & (!sk[66]) & (g1442) & (g1443)));
	assign g1445 = (((!sk[67]) & (!g123) & (!g552) & (g511) & (!g654)) + ((!sk[67]) & (!g123) & (!g552) & (g511) & (g654)) + ((!sk[67]) & (!g123) & (g552) & (g511) & (!g654)) + ((!sk[67]) & (!g123) & (g552) & (g511) & (g654)) + ((!sk[67]) & (g123) & (!g552) & (g511) & (!g654)) + ((!sk[67]) & (g123) & (!g552) & (g511) & (g654)) + ((!sk[67]) & (g123) & (g552) & (g511) & (!g654)) + ((!sk[67]) & (g123) & (g552) & (g511) & (g654)) + ((sk[67]) & (!g123) & (!g552) & (!g511) & (!g654)) + ((sk[67]) & (!g123) & (!g552) & (!g511) & (g654)) + ((sk[67]) & (!g123) & (!g552) & (g511) & (!g654)) + ((sk[67]) & (!g123) & (!g552) & (g511) & (g654)) + ((sk[67]) & (!g123) & (g552) & (!g511) & (g654)) + ((sk[67]) & (!g123) & (g552) & (g511) & (!g654)) + ((sk[67]) & (!g123) & (g552) & (g511) & (g654)));
	assign g1446 = (((!g77) & (!g123) & (!g270) & (sk[68]) & (!g1287) & (!g1445)) + ((!g77) & (!g123) & (g270) & (!sk[68]) & (!g1287) & (g1445)) + ((!g77) & (!g123) & (g270) & (!sk[68]) & (g1287) & (!g1445)) + ((!g77) & (!g123) & (g270) & (!sk[68]) & (g1287) & (g1445)) + ((!g77) & (g123) & (!g270) & (!sk[68]) & (!g1287) & (!g1445)) + ((!g77) & (g123) & (!g270) & (!sk[68]) & (!g1287) & (g1445)) + ((!g77) & (g123) & (!g270) & (!sk[68]) & (g1287) & (!g1445)) + ((!g77) & (g123) & (!g270) & (!sk[68]) & (g1287) & (g1445)) + ((!g77) & (g123) & (!g270) & (sk[68]) & (!g1287) & (!g1445)) + ((!g77) & (g123) & (g270) & (!sk[68]) & (!g1287) & (!g1445)) + ((!g77) & (g123) & (g270) & (!sk[68]) & (!g1287) & (g1445)) + ((!g77) & (g123) & (g270) & (!sk[68]) & (g1287) & (!g1445)) + ((!g77) & (g123) & (g270) & (!sk[68]) & (g1287) & (g1445)) + ((!g77) & (g123) & (g270) & (sk[68]) & (!g1287) & (!g1445)) + ((g77) & (!g123) & (g270) & (!sk[68]) & (!g1287) & (g1445)) + ((g77) & (!g123) & (g270) & (!sk[68]) & (g1287) & (!g1445)) + ((g77) & (!g123) & (g270) & (!sk[68]) & (g1287) & (g1445)) + ((g77) & (g123) & (!g270) & (!sk[68]) & (!g1287) & (!g1445)) + ((g77) & (g123) & (!g270) & (!sk[68]) & (!g1287) & (g1445)) + ((g77) & (g123) & (!g270) & (!sk[68]) & (g1287) & (!g1445)) + ((g77) & (g123) & (!g270) & (!sk[68]) & (g1287) & (g1445)) + ((g77) & (g123) & (!g270) & (sk[68]) & (!g1287) & (!g1445)) + ((g77) & (g123) & (g270) & (!sk[68]) & (!g1287) & (!g1445)) + ((g77) & (g123) & (g270) & (!sk[68]) & (!g1287) & (g1445)) + ((g77) & (g123) & (g270) & (!sk[68]) & (g1287) & (!g1445)) + ((g77) & (g123) & (g270) & (!sk[68]) & (g1287) & (g1445)) + ((g77) & (g123) & (g270) & (sk[68]) & (!g1287) & (!g1445)));
	assign g1447 = (((!g123) & (!g198) & (g1107) & (g1444) & (!g1222) & (g1446)) + ((g123) & (!g198) & (!g1107) & (!g1444) & (!g1222) & (g1446)) + ((g123) & (!g198) & (!g1107) & (g1444) & (!g1222) & (g1446)) + ((g123) & (!g198) & (g1107) & (!g1444) & (!g1222) & (g1446)) + ((g123) & (!g198) & (g1107) & (g1444) & (!g1222) & (g1446)));
	assign g1448 = (((!g1254) & (!g1352) & (g1408) & (!sk[70]) & (!g1441) & (g1447)) + ((!g1254) & (!g1352) & (g1408) & (!sk[70]) & (g1441) & (!g1447)) + ((!g1254) & (!g1352) & (g1408) & (!sk[70]) & (g1441) & (g1447)) + ((!g1254) & (g1352) & (!g1408) & (!sk[70]) & (!g1441) & (!g1447)) + ((!g1254) & (g1352) & (!g1408) & (!sk[70]) & (!g1441) & (g1447)) + ((!g1254) & (g1352) & (!g1408) & (!sk[70]) & (g1441) & (!g1447)) + ((!g1254) & (g1352) & (!g1408) & (!sk[70]) & (g1441) & (g1447)) + ((!g1254) & (g1352) & (!g1408) & (sk[70]) & (g1441) & (g1447)) + ((!g1254) & (g1352) & (g1408) & (!sk[70]) & (!g1441) & (!g1447)) + ((!g1254) & (g1352) & (g1408) & (!sk[70]) & (!g1441) & (g1447)) + ((!g1254) & (g1352) & (g1408) & (!sk[70]) & (g1441) & (!g1447)) + ((!g1254) & (g1352) & (g1408) & (!sk[70]) & (g1441) & (g1447)) + ((g1254) & (!g1352) & (g1408) & (!sk[70]) & (!g1441) & (g1447)) + ((g1254) & (!g1352) & (g1408) & (!sk[70]) & (g1441) & (!g1447)) + ((g1254) & (!g1352) & (g1408) & (!sk[70]) & (g1441) & (g1447)) + ((g1254) & (g1352) & (!g1408) & (!sk[70]) & (!g1441) & (!g1447)) + ((g1254) & (g1352) & (!g1408) & (!sk[70]) & (!g1441) & (g1447)) + ((g1254) & (g1352) & (!g1408) & (!sk[70]) & (g1441) & (!g1447)) + ((g1254) & (g1352) & (!g1408) & (!sk[70]) & (g1441) & (g1447)) + ((g1254) & (g1352) & (g1408) & (!sk[70]) & (!g1441) & (!g1447)) + ((g1254) & (g1352) & (g1408) & (!sk[70]) & (!g1441) & (g1447)) + ((g1254) & (g1352) & (g1408) & (!sk[70]) & (g1441) & (!g1447)) + ((g1254) & (g1352) & (g1408) & (!sk[70]) & (g1441) & (g1447)));
	assign g1449 = (((!g1456) & (!g1297) & (!sk[71]) & (g1436) & (!g1440) & (g1448)) + ((!g1456) & (!g1297) & (!sk[71]) & (g1436) & (g1440) & (!g1448)) + ((!g1456) & (!g1297) & (!sk[71]) & (g1436) & (g1440) & (g1448)) + ((!g1456) & (g1297) & (!sk[71]) & (!g1436) & (!g1440) & (!g1448)) + ((!g1456) & (g1297) & (!sk[71]) & (!g1436) & (!g1440) & (g1448)) + ((!g1456) & (g1297) & (!sk[71]) & (!g1436) & (g1440) & (!g1448)) + ((!g1456) & (g1297) & (!sk[71]) & (!g1436) & (g1440) & (g1448)) + ((!g1456) & (g1297) & (!sk[71]) & (g1436) & (!g1440) & (!g1448)) + ((!g1456) & (g1297) & (!sk[71]) & (g1436) & (!g1440) & (g1448)) + ((!g1456) & (g1297) & (!sk[71]) & (g1436) & (g1440) & (!g1448)) + ((!g1456) & (g1297) & (!sk[71]) & (g1436) & (g1440) & (g1448)) + ((g1456) & (!g1297) & (!sk[71]) & (g1436) & (!g1440) & (g1448)) + ((g1456) & (!g1297) & (!sk[71]) & (g1436) & (g1440) & (!g1448)) + ((g1456) & (!g1297) & (!sk[71]) & (g1436) & (g1440) & (g1448)) + ((g1456) & (g1297) & (!sk[71]) & (!g1436) & (!g1440) & (!g1448)) + ((g1456) & (g1297) & (!sk[71]) & (!g1436) & (!g1440) & (g1448)) + ((g1456) & (g1297) & (!sk[71]) & (!g1436) & (g1440) & (!g1448)) + ((g1456) & (g1297) & (!sk[71]) & (!g1436) & (g1440) & (g1448)) + ((g1456) & (g1297) & (!sk[71]) & (g1436) & (!g1440) & (!g1448)) + ((g1456) & (g1297) & (!sk[71]) & (g1436) & (!g1440) & (g1448)) + ((g1456) & (g1297) & (!sk[71]) & (g1436) & (g1440) & (!g1448)) + ((g1456) & (g1297) & (!sk[71]) & (g1436) & (g1440) & (g1448)) + ((g1456) & (g1297) & (sk[71]) & (g1436) & (g1440) & (g1448)));
	assign g1450 = (((!g2) & (!sk[72]) & (!g16) & (g43) & (!g38) & (g1070)) + ((!g2) & (!sk[72]) & (!g16) & (g43) & (g38) & (!g1070)) + ((!g2) & (!sk[72]) & (!g16) & (g43) & (g38) & (g1070)) + ((!g2) & (!sk[72]) & (g16) & (!g43) & (!g38) & (!g1070)) + ((!g2) & (!sk[72]) & (g16) & (!g43) & (!g38) & (g1070)) + ((!g2) & (!sk[72]) & (g16) & (!g43) & (g38) & (!g1070)) + ((!g2) & (!sk[72]) & (g16) & (!g43) & (g38) & (g1070)) + ((!g2) & (!sk[72]) & (g16) & (g43) & (!g38) & (!g1070)) + ((!g2) & (!sk[72]) & (g16) & (g43) & (!g38) & (g1070)) + ((!g2) & (!sk[72]) & (g16) & (g43) & (g38) & (!g1070)) + ((!g2) & (!sk[72]) & (g16) & (g43) & (g38) & (g1070)) + ((!g2) & (sk[72]) & (!g16) & (!g43) & (!g38) & (!g1070)) + ((!g2) & (sk[72]) & (!g16) & (g43) & (!g38) & (!g1070)) + ((!g2) & (sk[72]) & (g16) & (!g43) & (!g38) & (!g1070)) + ((!g2) & (sk[72]) & (g16) & (g43) & (!g38) & (!g1070)) + ((!g2) & (sk[72]) & (g16) & (g43) & (!g38) & (g1070)) + ((g2) & (!sk[72]) & (!g16) & (g43) & (!g38) & (g1070)) + ((g2) & (!sk[72]) & (!g16) & (g43) & (g38) & (!g1070)) + ((g2) & (!sk[72]) & (!g16) & (g43) & (g38) & (g1070)) + ((g2) & (!sk[72]) & (g16) & (!g43) & (!g38) & (!g1070)) + ((g2) & (!sk[72]) & (g16) & (!g43) & (!g38) & (g1070)) + ((g2) & (!sk[72]) & (g16) & (!g43) & (g38) & (!g1070)) + ((g2) & (!sk[72]) & (g16) & (!g43) & (g38) & (g1070)) + ((g2) & (!sk[72]) & (g16) & (g43) & (!g38) & (!g1070)) + ((g2) & (!sk[72]) & (g16) & (g43) & (!g38) & (g1070)) + ((g2) & (!sk[72]) & (g16) & (g43) & (g38) & (!g1070)) + ((g2) & (!sk[72]) & (g16) & (g43) & (g38) & (g1070)) + ((g2) & (sk[72]) & (!g16) & (!g43) & (!g38) & (!g1070)) + ((g2) & (sk[72]) & (!g16) & (g43) & (!g38) & (!g1070)) + ((g2) & (sk[72]) & (g16) & (!g43) & (!g38) & (!g1070)) + ((g2) & (sk[72]) & (g16) & (!g43) & (!g38) & (g1070)) + ((g2) & (sk[72]) & (g16) & (g43) & (!g38) & (!g1070)) + ((g2) & (sk[72]) & (g16) & (g43) & (!g38) & (g1070)));
	assign g1451 = (((g100) & (g711) & (g961) & (g1117) & (g1123) & (!g1450)));
	assign g1452 = (((!g91) & (!g107) & (!sk[74]) & (i_14_) & (!g164)) + ((!g91) & (!g107) & (!sk[74]) & (i_14_) & (g164)) + ((!g91) & (!g107) & (sk[74]) & (!i_14_) & (g164)) + ((!g91) & (!g107) & (sk[74]) & (i_14_) & (g164)) + ((!g91) & (g107) & (!sk[74]) & (i_14_) & (!g164)) + ((!g91) & (g107) & (!sk[74]) & (i_14_) & (g164)) + ((!g91) & (g107) & (sk[74]) & (!i_14_) & (g164)) + ((!g91) & (g107) & (sk[74]) & (i_14_) & (g164)) + ((g91) & (!g107) & (!sk[74]) & (i_14_) & (!g164)) + ((g91) & (!g107) & (!sk[74]) & (i_14_) & (g164)) + ((g91) & (!g107) & (sk[74]) & (i_14_) & (g164)) + ((g91) & (g107) & (!sk[74]) & (i_14_) & (!g164)) + ((g91) & (g107) & (!sk[74]) & (i_14_) & (g164)));
	assign g1453 = (((!g88) & (!g154) & (!g86) & (g1180) & (!g1179) & (!g1178)) + ((!g88) & (g154) & (!g86) & (g1180) & (!g1179) & (!g1178)) + ((!g88) & (g154) & (g86) & (g1180) & (!g1179) & (!g1178)) + ((g88) & (g154) & (!g86) & (g1180) & (!g1179) & (!g1178)) + ((g88) & (g154) & (g86) & (g1180) & (!g1179) & (!g1178)));
	assign g1454 = (((!g48) & (!i_7_) & (!i_8_) & (!g1068) & (!g1067) & (!g16)) + ((!g48) & (!i_7_) & (!i_8_) & (!g1068) & (!g1067) & (g16)) + ((!g48) & (!i_7_) & (!i_8_) & (!g1068) & (g1067) & (!g16)) + ((!g48) & (!i_7_) & (!i_8_) & (!g1068) & (g1067) & (g16)) + ((!g48) & (!i_7_) & (!i_8_) & (g1068) & (g1067) & (!g16)) + ((!g48) & (!i_7_) & (!i_8_) & (g1068) & (g1067) & (g16)) + ((!g48) & (!i_7_) & (i_8_) & (!g1068) & (!g1067) & (!g16)) + ((!g48) & (!i_7_) & (i_8_) & (!g1068) & (!g1067) & (g16)) + ((!g48) & (!i_7_) & (i_8_) & (!g1068) & (g1067) & (!g16)) + ((!g48) & (!i_7_) & (i_8_) & (!g1068) & (g1067) & (g16)) + ((!g48) & (!i_7_) & (i_8_) & (g1068) & (g1067) & (!g16)) + ((!g48) & (!i_7_) & (i_8_) & (g1068) & (g1067) & (g16)) + ((!g48) & (i_7_) & (!i_8_) & (!g1068) & (!g1067) & (!g16)) + ((!g48) & (i_7_) & (!i_8_) & (!g1068) & (!g1067) & (g16)) + ((!g48) & (i_7_) & (!i_8_) & (!g1068) & (g1067) & (!g16)) + ((!g48) & (i_7_) & (!i_8_) & (!g1068) & (g1067) & (g16)) + ((!g48) & (i_7_) & (!i_8_) & (g1068) & (g1067) & (!g16)) + ((!g48) & (i_7_) & (!i_8_) & (g1068) & (g1067) & (g16)) + ((!g48) & (i_7_) & (i_8_) & (!g1068) & (!g1067) & (!g16)) + ((!g48) & (i_7_) & (i_8_) & (!g1068) & (!g1067) & (g16)) + ((!g48) & (i_7_) & (i_8_) & (!g1068) & (g1067) & (!g16)) + ((!g48) & (i_7_) & (i_8_) & (!g1068) & (g1067) & (g16)) + ((!g48) & (i_7_) & (i_8_) & (g1068) & (g1067) & (!g16)) + ((!g48) & (i_7_) & (i_8_) & (g1068) & (g1067) & (g16)) + ((g48) & (!i_7_) & (!i_8_) & (!g1068) & (!g1067) & (!g16)) + ((g48) & (!i_7_) & (!i_8_) & (!g1068) & (!g1067) & (g16)) + ((g48) & (!i_7_) & (!i_8_) & (!g1068) & (g1067) & (!g16)) + ((g48) & (!i_7_) & (!i_8_) & (!g1068) & (g1067) & (g16)) + ((g48) & (!i_7_) & (!i_8_) & (g1068) & (g1067) & (!g16)) + ((g48) & (!i_7_) & (!i_8_) & (g1068) & (g1067) & (g16)) + ((g48) & (!i_7_) & (i_8_) & (!g1068) & (!g1067) & (!g16)) + ((g48) & (!i_7_) & (i_8_) & (!g1068) & (g1067) & (!g16)) + ((g48) & (!i_7_) & (i_8_) & (g1068) & (g1067) & (!g16)) + ((g48) & (i_7_) & (!i_8_) & (!g1068) & (!g1067) & (!g16)) + ((g48) & (i_7_) & (!i_8_) & (!g1068) & (!g1067) & (g16)) + ((g48) & (i_7_) & (!i_8_) & (!g1068) & (g1067) & (!g16)) + ((g48) & (i_7_) & (!i_8_) & (!g1068) & (g1067) & (g16)) + ((g48) & (i_7_) & (!i_8_) & (g1068) & (g1067) & (!g16)) + ((g48) & (i_7_) & (!i_8_) & (g1068) & (g1067) & (g16)) + ((g48) & (i_7_) & (i_8_) & (!g1068) & (!g1067) & (!g16)) + ((g48) & (i_7_) & (i_8_) & (!g1068) & (!g1067) & (g16)) + ((g48) & (i_7_) & (i_8_) & (!g1068) & (g1067) & (!g16)) + ((g48) & (i_7_) & (i_8_) & (!g1068) & (g1067) & (g16)) + ((g48) & (i_7_) & (i_8_) & (g1068) & (g1067) & (!g16)) + ((g48) & (i_7_) & (i_8_) & (g1068) & (g1067) & (g16)));
	assign g1455 = (((!g36) & (!sk[77]) & (!g35) & (i_14_) & (!g154)) + ((!g36) & (!sk[77]) & (!g35) & (i_14_) & (g154)) + ((!g36) & (!sk[77]) & (g35) & (i_14_) & (!g154)) + ((!g36) & (!sk[77]) & (g35) & (i_14_) & (g154)) + ((!g36) & (sk[77]) & (g35) & (i_14_) & (!g154)) + ((g36) & (!sk[77]) & (!g35) & (i_14_) & (!g154)) + ((g36) & (!sk[77]) & (!g35) & (i_14_) & (g154)) + ((g36) & (!sk[77]) & (g35) & (i_14_) & (!g154)) + ((g36) & (!sk[77]) & (g35) & (i_14_) & (g154)) + ((g36) & (sk[77]) & (!g35) & (!i_14_) & (!g154)) + ((g36) & (sk[77]) & (!g35) & (i_14_) & (!g154)) + ((g36) & (sk[77]) & (g35) & (!i_14_) & (!g154)) + ((g36) & (sk[77]) & (g35) & (i_14_) & (!g154)));
	assign g1456 = (((!i_10_) & (!i_9_) & (!g118) & (!g10) & (!i_8_) & (!i_11_)) + ((!i_10_) & (!i_9_) & (!g118) & (!g10) & (!i_8_) & (i_11_)) + ((!i_10_) & (!i_9_) & (!g118) & (!g10) & (i_8_) & (!i_11_)) + ((!i_10_) & (!i_9_) & (!g118) & (!g10) & (i_8_) & (i_11_)) + ((!i_10_) & (!i_9_) & (!g118) & (g10) & (!i_8_) & (!i_11_)) + ((!i_10_) & (!i_9_) & (!g118) & (g10) & (!i_8_) & (i_11_)) + ((!i_10_) & (!i_9_) & (!g118) & (g10) & (i_8_) & (!i_11_)) + ((!i_10_) & (!i_9_) & (!g118) & (g10) & (i_8_) & (i_11_)) + ((!i_10_) & (!i_9_) & (g118) & (!g10) & (!i_8_) & (!i_11_)) + ((!i_10_) & (!i_9_) & (g118) & (!g10) & (!i_8_) & (i_11_)) + ((!i_10_) & (!i_9_) & (g118) & (!g10) & (i_8_) & (!i_11_)) + ((!i_10_) & (!i_9_) & (g118) & (!g10) & (i_8_) & (i_11_)) + ((!i_10_) & (!i_9_) & (g118) & (g10) & (!i_8_) & (!i_11_)) + ((!i_10_) & (!i_9_) & (g118) & (g10) & (i_8_) & (i_11_)) + ((!i_10_) & (i_9_) & (!g118) & (!g10) & (!i_8_) & (!i_11_)) + ((!i_10_) & (i_9_) & (!g118) & (!g10) & (!i_8_) & (i_11_)) + ((!i_10_) & (i_9_) & (!g118) & (!g10) & (i_8_) & (!i_11_)) + ((!i_10_) & (i_9_) & (!g118) & (!g10) & (i_8_) & (i_11_)) + ((!i_10_) & (i_9_) & (!g118) & (g10) & (!i_8_) & (!i_11_)) + ((!i_10_) & (i_9_) & (!g118) & (g10) & (!i_8_) & (i_11_)) + ((!i_10_) & (i_9_) & (!g118) & (g10) & (i_8_) & (!i_11_)) + ((!i_10_) & (i_9_) & (!g118) & (g10) & (i_8_) & (i_11_)) + ((!i_10_) & (i_9_) & (g118) & (!g10) & (!i_8_) & (!i_11_)) + ((!i_10_) & (i_9_) & (g118) & (!g10) & (!i_8_) & (i_11_)) + ((!i_10_) & (i_9_) & (g118) & (!g10) & (i_8_) & (!i_11_)) + ((!i_10_) & (i_9_) & (g118) & (!g10) & (i_8_) & (i_11_)) + ((!i_10_) & (i_9_) & (g118) & (g10) & (!i_8_) & (i_11_)) + ((!i_10_) & (i_9_) & (g118) & (g10) & (i_8_) & (!i_11_)) + ((!i_10_) & (i_9_) & (g118) & (g10) & (i_8_) & (i_11_)) + ((i_10_) & (!i_9_) & (!g118) & (!g10) & (!i_8_) & (!i_11_)) + ((i_10_) & (!i_9_) & (!g118) & (!g10) & (!i_8_) & (i_11_)) + ((i_10_) & (!i_9_) & (!g118) & (!g10) & (i_8_) & (!i_11_)) + ((i_10_) & (!i_9_) & (!g118) & (!g10) & (i_8_) & (i_11_)) + ((i_10_) & (!i_9_) & (!g118) & (g10) & (!i_8_) & (!i_11_)) + ((i_10_) & (!i_9_) & (!g118) & (g10) & (!i_8_) & (i_11_)) + ((i_10_) & (!i_9_) & (!g118) & (g10) & (i_8_) & (!i_11_)) + ((i_10_) & (!i_9_) & (!g118) & (g10) & (i_8_) & (i_11_)) + ((i_10_) & (!i_9_) & (g118) & (!g10) & (!i_8_) & (!i_11_)) + ((i_10_) & (!i_9_) & (g118) & (!g10) & (!i_8_) & (i_11_)) + ((i_10_) & (!i_9_) & (g118) & (!g10) & (i_8_) & (!i_11_)) + ((i_10_) & (!i_9_) & (g118) & (!g10) & (i_8_) & (i_11_)) + ((i_10_) & (!i_9_) & (g118) & (g10) & (!i_8_) & (i_11_)) + ((i_10_) & (!i_9_) & (g118) & (g10) & (i_8_) & (!i_11_)) + ((i_10_) & (!i_9_) & (g118) & (g10) & (i_8_) & (i_11_)) + ((i_10_) & (i_9_) & (!g118) & (!g10) & (!i_8_) & (!i_11_)) + ((i_10_) & (i_9_) & (!g118) & (!g10) & (!i_8_) & (i_11_)) + ((i_10_) & (i_9_) & (!g118) & (!g10) & (i_8_) & (!i_11_)) + ((i_10_) & (i_9_) & (!g118) & (!g10) & (i_8_) & (i_11_)) + ((i_10_) & (i_9_) & (!g118) & (g10) & (!i_8_) & (!i_11_)) + ((i_10_) & (i_9_) & (!g118) & (g10) & (!i_8_) & (i_11_)) + ((i_10_) & (i_9_) & (!g118) & (g10) & (i_8_) & (!i_11_)) + ((i_10_) & (i_9_) & (!g118) & (g10) & (i_8_) & (i_11_)) + ((i_10_) & (i_9_) & (g118) & (!g10) & (!i_8_) & (!i_11_)) + ((i_10_) & (i_9_) & (g118) & (!g10) & (!i_8_) & (i_11_)) + ((i_10_) & (i_9_) & (g118) & (!g10) & (i_8_) & (!i_11_)) + ((i_10_) & (i_9_) & (g118) & (!g10) & (i_8_) & (i_11_)) + ((i_10_) & (i_9_) & (g118) & (g10) & (!i_8_) & (!i_11_)) + ((i_10_) & (i_9_) & (g118) & (g10) & (!i_8_) & (i_11_)) + ((i_10_) & (i_9_) & (g118) & (g10) & (i_8_) & (!i_11_)) + ((i_10_) & (i_9_) & (g118) & (g10) & (i_8_) & (i_11_)));
	assign g1457 = (((!i_14_) & (!g682) & (!sk[79]) & (g681) & (!g226) & (g69)) + ((!i_14_) & (!g682) & (!sk[79]) & (g681) & (g226) & (!g69)) + ((!i_14_) & (!g682) & (!sk[79]) & (g681) & (g226) & (g69)) + ((!i_14_) & (g682) & (!sk[79]) & (!g681) & (!g226) & (!g69)) + ((!i_14_) & (g682) & (!sk[79]) & (!g681) & (!g226) & (g69)) + ((!i_14_) & (g682) & (!sk[79]) & (!g681) & (g226) & (!g69)) + ((!i_14_) & (g682) & (!sk[79]) & (!g681) & (g226) & (g69)) + ((!i_14_) & (g682) & (!sk[79]) & (g681) & (!g226) & (!g69)) + ((!i_14_) & (g682) & (!sk[79]) & (g681) & (!g226) & (g69)) + ((!i_14_) & (g682) & (!sk[79]) & (g681) & (g226) & (!g69)) + ((!i_14_) & (g682) & (!sk[79]) & (g681) & (g226) & (g69)) + ((!i_14_) & (g682) & (sk[79]) & (!g681) & (!g226) & (!g69)) + ((!i_14_) & (g682) & (sk[79]) & (!g681) & (g226) & (!g69)) + ((!i_14_) & (g682) & (sk[79]) & (!g681) & (g226) & (g69)) + ((i_14_) & (!g682) & (!sk[79]) & (g681) & (!g226) & (g69)) + ((i_14_) & (!g682) & (!sk[79]) & (g681) & (g226) & (!g69)) + ((i_14_) & (!g682) & (!sk[79]) & (g681) & (g226) & (g69)) + ((i_14_) & (g682) & (!sk[79]) & (!g681) & (!g226) & (!g69)) + ((i_14_) & (g682) & (!sk[79]) & (!g681) & (!g226) & (g69)) + ((i_14_) & (g682) & (!sk[79]) & (!g681) & (g226) & (!g69)) + ((i_14_) & (g682) & (!sk[79]) & (!g681) & (g226) & (g69)) + ((i_14_) & (g682) & (!sk[79]) & (g681) & (!g226) & (!g69)) + ((i_14_) & (g682) & (!sk[79]) & (g681) & (!g226) & (g69)) + ((i_14_) & (g682) & (!sk[79]) & (g681) & (g226) & (!g69)) + ((i_14_) & (g682) & (!sk[79]) & (g681) & (g226) & (g69)) + ((i_14_) & (g682) & (sk[79]) & (!g681) & (!g226) & (!g69)) + ((i_14_) & (g682) & (sk[79]) & (!g681) & (!g226) & (g69)) + ((i_14_) & (g682) & (sk[79]) & (!g681) & (g226) & (!g69)) + ((i_14_) & (g682) & (sk[79]) & (!g681) & (g226) & (g69)));
	assign g1458 = (((!g605) & (!g73) & (!g606) & (!g604) & (!g603) & (!g602)) + ((!g605) & (g73) & (!g606) & (!g604) & (!g603) & (!g602)) + ((g605) & (!g73) & (!g606) & (!g604) & (!g603) & (!g602)));
	assign g1459 = (((g71) & (g15) & (!i_7_) & (i_6_) & (i_11_) & (!i_10_)) + ((g71) & (g15) & (i_7_) & (!i_6_) & (i_11_) & (!i_10_)));
	assign g1460 = (((!sk[82]) & (g73) & (!g1461)) + ((!sk[82]) & (g73) & (g1461)) + ((sk[82]) & (g73) & (!g1461)));
	assign g1461 = (((!sk[83]) & (g73) & (!g1462)) + ((!sk[83]) & (g73) & (g1462)) + ((sk[83]) & (g73) & (g1462)));
	assign g1462 = (((!g1463) & (sk[84]) & (!g1464)) + ((g1463) & (!sk[84]) & (!g1464)) + ((g1463) & (!sk[84]) & (g1464)));
	assign g1463 = (((!i_8_) & (sk[85]) & (g1465)) + ((i_8_) & (!sk[85]) & (!g1465)) + ((i_8_) & (!sk[85]) & (g1465)));
	assign g1464 = (((i_8_) & (!sk[86]) & (!g1466)) + ((i_8_) & (!sk[86]) & (g1466)) + ((i_8_) & (sk[86]) & (g1466)));
	assign g1465 = (((!g628) & (!g608) & (g898) & (!sk[87]) & (!g340)) + ((!g628) & (!g608) & (g898) & (!sk[87]) & (g340)) + ((!g628) & (g608) & (g898) & (!sk[87]) & (!g340)) + ((!g628) & (g608) & (g898) & (!sk[87]) & (g340)) + ((g628) & (!g608) & (g898) & (!sk[87]) & (!g340)) + ((g628) & (!g608) & (g898) & (!sk[87]) & (g340)) + ((g628) & (g608) & (g898) & (!sk[87]) & (!g340)) + ((g628) & (g608) & (g898) & (!sk[87]) & (g340)) + ((g628) & (g608) & (g898) & (sk[87]) & (g340)));
	assign g1466 = (((!sk[88]) & (g608) & (!g847)) + ((!sk[88]) & (g608) & (g847)) + ((sk[88]) & (g608) & (g847)));
	assign g1467 = (((!sk[89]) & (g1468) & (!g1469)) + ((!sk[89]) & (g1468) & (g1469)) + ((sk[89]) & (!g1468) & (!g1469)));
	assign g1468 = (((!sk[90]) & (g168) & (!g1470)) + ((!sk[90]) & (g168) & (g1470)) + ((sk[90]) & (!g168) & (g1470)));
	assign g1469 = (((!sk[91]) & (g168) & (!g1472)) + ((!sk[91]) & (g168) & (g1472)) + ((sk[91]) & (g168) & (g1472)));
	assign g1470 = (((!g105) & (sk[92]) & (!g1471)) + ((g105) & (!sk[92]) & (!g1471)) + ((g105) & (!sk[92]) & (g1471)));
	assign g1471 = (((!g105) & (sk[93]) & (g1475)) + ((g105) & (!sk[93]) & (!g1475)) + ((g105) & (!sk[93]) & (g1475)));
	assign g1472 = (((!g1473) & (sk[94]) & (!g1474)) + ((g1473) & (!sk[94]) & (!g1474)) + ((g1473) & (!sk[94]) & (g1474)));
	assign g1473 = (((!g105) & (sk[95]) & (g1476)) + ((g105) & (!sk[95]) & (!g1476)) + ((g105) & (!sk[95]) & (g1476)));
	assign g1474 = (((g105) & (!sk[96]) & (!g1477)) + ((g105) & (!sk[96]) & (g1477)) + ((g105) & (sk[96]) & (g1477)));
	assign g1475 = (((!sk[97]) & (!g626) & (!g343) & (g851)) + ((!sk[97]) & (!g626) & (g343) & (!g851)) + ((!sk[97]) & (!g626) & (g343) & (g851)) + ((!sk[97]) & (g626) & (!g343) & (g851)) + ((!sk[97]) & (g626) & (g343) & (!g851)) + ((!sk[97]) & (g626) & (g343) & (g851)) + ((sk[97]) & (!g626) & (g343) & (g851)));
	assign g1476 = (((!g626) & (!g343) & (!sk[98]) & (g851) & (!g945)) + ((!g626) & (!g343) & (!sk[98]) & (g851) & (g945)) + ((!g626) & (g343) & (!sk[98]) & (g851) & (!g945)) + ((!g626) & (g343) & (!sk[98]) & (g851) & (g945)) + ((!g626) & (g343) & (sk[98]) & (g851) & (g945)) + ((g626) & (!g343) & (!sk[98]) & (g851) & (!g945)) + ((g626) & (!g343) & (!sk[98]) & (g851) & (g945)) + ((g626) & (g343) & (!sk[98]) & (g851) & (!g945)) + ((g626) & (g343) & (!sk[98]) & (g851) & (g945)));
	assign g1477 = (((!g626) & (!g343) & (!g102) & (sk[99]) & (g945)) + ((!g626) & (!g343) & (g102) & (!sk[99]) & (!g945)) + ((!g626) & (!g343) & (g102) & (!sk[99]) & (g945)) + ((!g626) & (g343) & (!g102) & (sk[99]) & (g945)) + ((!g626) & (g343) & (g102) & (!sk[99]) & (!g945)) + ((!g626) & (g343) & (g102) & (!sk[99]) & (g945)) + ((!g626) & (g343) & (g102) & (sk[99]) & (g945)) + ((g626) & (!g343) & (!g102) & (sk[99]) & (g945)) + ((g626) & (!g343) & (g102) & (!sk[99]) & (!g945)) + ((g626) & (!g343) & (g102) & (!sk[99]) & (g945)) + ((g626) & (g343) & (!g102) & (sk[99]) & (g945)) + ((g626) & (g343) & (g102) & (!sk[99]) & (!g945)) + ((g626) & (g343) & (g102) & (!sk[99]) & (g945)));
	assign g1478 = (((!g1479) & (sk[100]) & (!g1480)) + ((g1479) & (!sk[100]) & (!g1480)) + ((g1479) & (!sk[100]) & (g1480)));
	assign g1479 = (((!g23) & (sk[101]) & (g1481)) + ((g23) & (!sk[101]) & (!g1481)) + ((g23) & (!sk[101]) & (g1481)));
	assign g1480 = (((g23) & (!sk[102]) & (!g1482)) + ((g23) & (!sk[102]) & (g1482)) + ((g23) & (sk[102]) & (g1482)));
	assign g1481 = (((g142) & (!sk[103]) & (!g1485)) + ((g142) & (!sk[103]) & (g1485)) + ((g142) & (sk[103]) & (g1485)));
	assign g1482 = (((!g1483) & (sk[104]) & (!g1484)) + ((g1483) & (!sk[104]) & (!g1484)) + ((g1483) & (!sk[104]) & (g1484)));
	assign g1483 = (((!g142) & (sk[105]) & (g1486)) + ((g142) & (!sk[105]) & (!g1486)) + ((g142) & (!sk[105]) & (g1486)));
	assign g1484 = (((g142) & (!sk[106]) & (!g1487)) + ((g142) & (!sk[106]) & (g1487)) + ((g142) & (sk[106]) & (g1487)));
	assign g1485 = (((!g703) & (!sk[107]) & (!g518) & (g154) & (!g896)) + ((!g703) & (!sk[107]) & (!g518) & (g154) & (g896)) + ((!g703) & (!sk[107]) & (g518) & (g154) & (!g896)) + ((!g703) & (!sk[107]) & (g518) & (g154) & (g896)) + ((!g703) & (sk[107]) & (!g518) & (g154) & (g896)) + ((g703) & (!sk[107]) & (!g518) & (g154) & (!g896)) + ((g703) & (!sk[107]) & (!g518) & (g154) & (g896)) + ((g703) & (!sk[107]) & (g518) & (g154) & (!g896)) + ((g703) & (!sk[107]) & (g518) & (g154) & (g896)) + ((g703) & (sk[107]) & (!g518) & (g154) & (g896)) + ((g703) & (sk[107]) & (g518) & (g154) & (g896)));
	assign g1486 = (((!g703) & (!g518) & (!sk[108]) & (g25) & (!g896)) + ((!g703) & (!g518) & (!sk[108]) & (g25) & (g896)) + ((!g703) & (!g518) & (sk[108]) & (g25) & (g896)) + ((!g703) & (g518) & (!sk[108]) & (g25) & (!g896)) + ((!g703) & (g518) & (!sk[108]) & (g25) & (g896)) + ((g703) & (!g518) & (!sk[108]) & (g25) & (!g896)) + ((g703) & (!g518) & (!sk[108]) & (g25) & (g896)) + ((g703) & (!g518) & (sk[108]) & (g25) & (g896)) + ((g703) & (g518) & (!sk[108]) & (g25) & (!g896)) + ((g703) & (g518) & (!sk[108]) & (g25) & (g896)) + ((g703) & (g518) & (sk[108]) & (g25) & (g896)));
	assign g1487 = (((!sk[109]) & (!g703) & (!g518) & (g896)) + ((!sk[109]) & (!g703) & (g518) & (!g896)) + ((!sk[109]) & (!g703) & (g518) & (g896)) + ((!sk[109]) & (g703) & (!g518) & (g896)) + ((!sk[109]) & (g703) & (g518) & (!g896)) + ((!sk[109]) & (g703) & (g518) & (g896)) + ((sk[109]) & (!g703) & (!g518) & (g896)) + ((sk[109]) & (g703) & (!g518) & (g896)) + ((sk[109]) & (g703) & (g518) & (g896)));
	assign g1488 = (((!g1489) & (sk[110]) & (!g1490)) + ((g1489) & (!sk[110]) & (!g1490)) + ((g1489) & (!sk[110]) & (g1490)));
	assign g1489 = (((!sk[111]) & (g130) & (!g1491)) + ((!sk[111]) & (g130) & (g1491)) + ((sk[111]) & (!g130) & (g1491)));
	assign g1490 = (((!sk[112]) & (g130) & (!g1494)) + ((!sk[112]) & (g130) & (g1494)) + ((sk[112]) & (g130) & (g1494)));
	assign g1491 = (((!sk[113]) & (g1492) & (!g1493)) + ((!sk[113]) & (g1492) & (g1493)) + ((sk[113]) & (!g1492) & (!g1493)));
	assign g1492 = (((!g123) & (sk[114]) & (g1497)) + ((g123) & (!sk[114]) & (!g1497)) + ((g123) & (!sk[114]) & (g1497)));
	assign g1493 = (((g123) & (!sk[115]) & (!g1498)) + ((g123) & (!sk[115]) & (g1498)) + ((g123) & (sk[115]) & (g1498)));
	assign g1494 = (((!g1495) & (sk[116]) & (!g1496)) + ((g1495) & (!sk[116]) & (!g1496)) + ((g1495) & (!sk[116]) & (g1496)));
	assign g1495 = (((!sk[117]) & (g123) & (!g1499)) + ((!sk[117]) & (g123) & (g1499)) + ((sk[117]) & (!g123) & (g1499)));
	assign g1496 = (((!sk[118]) & (g123) & (!g1500)) + ((!sk[118]) & (g123) & (g1500)) + ((sk[118]) & (g123) & (g1500)));
	assign g1497 = (((!g872) & (!g868) & (!sk[119]) & (g847) & (!g848)) + ((!g872) & (!g868) & (!sk[119]) & (g847) & (g848)) + ((!g872) & (g868) & (!sk[119]) & (g847) & (!g848)) + ((!g872) & (g868) & (!sk[119]) & (g847) & (g848)) + ((g872) & (!g868) & (!sk[119]) & (g847) & (!g848)) + ((g872) & (!g868) & (!sk[119]) & (g847) & (g848)) + ((g872) & (g868) & (!sk[119]) & (g847) & (!g848)) + ((g872) & (g868) & (!sk[119]) & (g847) & (g848)) + ((g872) & (g868) & (sk[119]) & (g847) & (g848)));
	assign g1498 = (((!sk[120]) & (!g872) & (!g868) & (g848)) + ((!sk[120]) & (!g872) & (g868) & (!g848)) + ((!sk[120]) & (!g872) & (g868) & (g848)) + ((!sk[120]) & (g872) & (!g868) & (g848)) + ((!sk[120]) & (g872) & (g868) & (!g848)) + ((!sk[120]) & (g872) & (g868) & (g848)) + ((sk[120]) & (g872) & (g868) & (g848)));
	assign g1499 = (((!g872) & (!sk[121]) & (!g868) & (g847) & (!g848)) + ((!g872) & (!sk[121]) & (!g868) & (g847) & (g848)) + ((!g872) & (!sk[121]) & (g868) & (g847) & (!g848)) + ((!g872) & (!sk[121]) & (g868) & (g847) & (g848)) + ((g872) & (!sk[121]) & (!g868) & (g847) & (!g848)) + ((g872) & (!sk[121]) & (!g868) & (g847) & (g848)) + ((g872) & (!sk[121]) & (g868) & (g847) & (!g848)) + ((g872) & (!sk[121]) & (g868) & (g847) & (g848)) + ((g872) & (sk[121]) & (g868) & (g847) & (g848)));
	assign g1500 = (((!g872) & (!g868) & (!sk[122]) & (g159) & (!g848)) + ((!g872) & (!g868) & (!sk[122]) & (g159) & (g848)) + ((!g872) & (g868) & (!sk[122]) & (g159) & (!g848)) + ((!g872) & (g868) & (!sk[122]) & (g159) & (g848)) + ((g872) & (!g868) & (!sk[122]) & (g159) & (!g848)) + ((g872) & (!g868) & (!sk[122]) & (g159) & (g848)) + ((g872) & (g868) & (!sk[122]) & (g159) & (!g848)) + ((g872) & (g868) & (!sk[122]) & (g159) & (g848)) + ((g872) & (g868) & (sk[122]) & (!g159) & (g848)) + ((g872) & (g868) & (sk[122]) & (g159) & (!g848)) + ((g872) & (g868) & (sk[122]) & (g159) & (g848)));
	assign g1501 = (((!sk[123]) & (g1502) & (!g1503)) + ((!sk[123]) & (g1502) & (g1503)) + ((sk[123]) & (!g1502) & (!g1503)));
	assign g1502 = (((!sk[124]) & (g253) & (!g1504)) + ((!sk[124]) & (g253) & (g1504)) + ((sk[124]) & (!g253) & (g1504)));
	assign g1503 = (((g253) & (!sk[125]) & (!g1505)) + ((g253) & (!sk[125]) & (g1505)) + ((g253) & (sk[125]) & (g1505)));
	assign g1504 = (((g851) & (!sk[126]) & (!g1508)) + ((g851) & (!sk[126]) & (g1508)) + ((g851) & (sk[126]) & (g1508)));
	assign g1505 = (((!sk[127]) & (g1506) & (!g1507)) + ((!sk[127]) & (g1506) & (g1507)) + ((sk[127]) & (!g1506) & (!g1507)));
	assign g1506 = (((!g851) & (sk[0]) & (g1509)) + ((g851) & (!sk[0]) & (!g1509)) + ((g851) & (!sk[0]) & (g1509)));
	assign g1507 = (((g851) & (!sk[1]) & (!g1510)) + ((g851) & (!sk[1]) & (g1510)) + ((g851) & (sk[1]) & (g1510)));
	assign g1508 = (((!sk[2]) & (g862) & (!g684)) + ((!sk[2]) & (g862) & (g684)) + ((sk[2]) & (g862) & (g684)));
	assign g1509 = (((!g75) & (!g862) & (!sk[3]) & (g408) & (!g356)) + ((!g75) & (!g862) & (!sk[3]) & (g408) & (g356)) + ((!g75) & (g862) & (!sk[3]) & (g408) & (!g356)) + ((!g75) & (g862) & (!sk[3]) & (g408) & (g356)) + ((g75) & (!g862) & (!sk[3]) & (g408) & (!g356)) + ((g75) & (!g862) & (!sk[3]) & (g408) & (g356)) + ((g75) & (g862) & (!sk[3]) & (g408) & (!g356)) + ((g75) & (g862) & (!sk[3]) & (g408) & (g356)) + ((g75) & (g862) & (sk[3]) & (g408) & (!g356)));
	assign g1510 = (((!g862) & (!g684) & (!sk[4]) & (g356)) + ((!g862) & (g684) & (!sk[4]) & (!g356)) + ((!g862) & (g684) & (!sk[4]) & (g356)) + ((g862) & (!g684) & (!sk[4]) & (g356)) + ((g862) & (!g684) & (sk[4]) & (!g356)) + ((g862) & (g684) & (!sk[4]) & (!g356)) + ((g862) & (g684) & (!sk[4]) & (g356)) + ((g862) & (g684) & (sk[4]) & (!g356)) + ((g862) & (g684) & (sk[4]) & (g356)));
	assign g1511 = (((!sk[5]) & (g76) & (!g1512)) + ((!sk[5]) & (g76) & (g1512)) + ((sk[5]) & (!g76) & (!g1512)));
	assign g1512 = (((!sk[6]) & (g76) & (!g1513)) + ((!sk[6]) & (g76) & (g1513)) + ((sk[6]) & (!g76) & (g1513)));
	assign g1513 = (((!g1514) & (sk[7]) & (!g1515)) + ((g1514) & (!sk[7]) & (!g1515)) + ((g1514) & (!sk[7]) & (g1515)));
	assign g1514 = (((!i_11_) & (sk[8]) & (g1516)) + ((i_11_) & (!sk[8]) & (!g1516)) + ((i_11_) & (!sk[8]) & (g1516)));
	assign g1515 = (((i_11_) & (!sk[9]) & (!g1517)) + ((i_11_) & (!sk[9]) & (g1517)) + ((i_11_) & (sk[9]) & (g1517)));
	assign g1516 = (((!i_15_) & (!i_10_) & (!sk[10]) & (g436) & (!i_9_)) + ((!i_15_) & (!i_10_) & (!sk[10]) & (g436) & (i_9_)) + ((!i_15_) & (!i_10_) & (sk[10]) & (!g436) & (!i_9_)) + ((!i_15_) & (!i_10_) & (sk[10]) & (!g436) & (i_9_)) + ((!i_15_) & (!i_10_) & (sk[10]) & (g436) & (i_9_)) + ((!i_15_) & (i_10_) & (!sk[10]) & (g436) & (!i_9_)) + ((!i_15_) & (i_10_) & (!sk[10]) & (g436) & (i_9_)) + ((!i_15_) & (i_10_) & (sk[10]) & (!g436) & (!i_9_)) + ((!i_15_) & (i_10_) & (sk[10]) & (!g436) & (i_9_)) + ((!i_15_) & (i_10_) & (sk[10]) & (g436) & (!i_9_)) + ((!i_15_) & (i_10_) & (sk[10]) & (g436) & (i_9_)) + ((i_15_) & (!i_10_) & (!sk[10]) & (g436) & (!i_9_)) + ((i_15_) & (!i_10_) & (!sk[10]) & (g436) & (i_9_)) + ((i_15_) & (!i_10_) & (sk[10]) & (!g436) & (!i_9_)) + ((i_15_) & (!i_10_) & (sk[10]) & (!g436) & (i_9_)) + ((i_15_) & (!i_10_) & (sk[10]) & (g436) & (!i_9_)) + ((i_15_) & (!i_10_) & (sk[10]) & (g436) & (i_9_)) + ((i_15_) & (i_10_) & (!sk[10]) & (g436) & (!i_9_)) + ((i_15_) & (i_10_) & (!sk[10]) & (g436) & (i_9_)) + ((i_15_) & (i_10_) & (sk[10]) & (!g436) & (!i_9_)) + ((i_15_) & (i_10_) & (sk[10]) & (!g436) & (i_9_)) + ((i_15_) & (i_10_) & (sk[10]) & (g436) & (!i_9_)) + ((i_15_) & (i_10_) & (sk[10]) & (g436) & (i_9_)));
	assign g1517 = (((!sk[11]) & (!i_15_) & (!i_10_) & (g422) & (!i_9_)) + ((!sk[11]) & (!i_15_) & (!i_10_) & (g422) & (i_9_)) + ((!sk[11]) & (!i_15_) & (i_10_) & (g422) & (!i_9_)) + ((!sk[11]) & (!i_15_) & (i_10_) & (g422) & (i_9_)) + ((!sk[11]) & (i_15_) & (!i_10_) & (g422) & (!i_9_)) + ((!sk[11]) & (i_15_) & (!i_10_) & (g422) & (i_9_)) + ((!sk[11]) & (i_15_) & (i_10_) & (g422) & (!i_9_)) + ((!sk[11]) & (i_15_) & (i_10_) & (g422) & (i_9_)) + ((sk[11]) & (!i_15_) & (!i_10_) & (!g422) & (!i_9_)) + ((sk[11]) & (!i_15_) & (!i_10_) & (!g422) & (i_9_)) + ((sk[11]) & (!i_15_) & (!i_10_) & (g422) & (!i_9_)) + ((sk[11]) & (!i_15_) & (!i_10_) & (g422) & (i_9_)) + ((sk[11]) & (!i_15_) & (i_10_) & (!g422) & (!i_9_)) + ((sk[11]) & (!i_15_) & (i_10_) & (!g422) & (i_9_)) + ((sk[11]) & (!i_15_) & (i_10_) & (g422) & (!i_9_)) + ((sk[11]) & (i_15_) & (!i_10_) & (!g422) & (!i_9_)) + ((sk[11]) & (i_15_) & (!i_10_) & (!g422) & (i_9_)) + ((sk[11]) & (i_15_) & (!i_10_) & (g422) & (!i_9_)) + ((sk[11]) & (i_15_) & (!i_10_) & (g422) & (i_9_)) + ((sk[11]) & (i_15_) & (i_10_) & (!g422) & (!i_9_)) + ((sk[11]) & (i_15_) & (i_10_) & (!g422) & (i_9_)) + ((sk[11]) & (i_15_) & (i_10_) & (g422) & (!i_9_)) + ((sk[11]) & (i_15_) & (i_10_) & (g422) & (i_9_)));
	assign g1518 = (((!sk[12]) & (g1519) & (!g1520)) + ((!sk[12]) & (g1519) & (g1520)) + ((sk[12]) & (!g1519) & (!g1520)));
	assign g1519 = (((!g125) & (sk[13]) & (g1521)) + ((g125) & (!sk[13]) & (!g1521)) + ((g125) & (!sk[13]) & (g1521)));
	assign g1520 = (((!sk[14]) & (g125) & (!g1524)) + ((!sk[14]) & (g125) & (g1524)) + ((sk[14]) & (g125) & (g1524)));
	assign g1521 = (((!sk[15]) & (g1522) & (!g1523)) + ((!sk[15]) & (g1522) & (g1523)) + ((sk[15]) & (!g1522) & (!g1523)));
	assign g1522 = (((!sk[16]) & (g154) & (!g1527)) + ((!sk[16]) & (g154) & (g1527)) + ((sk[16]) & (!g154) & (g1527)));
	assign g1523 = (((!sk[17]) & (g154) & (!g1528)) + ((!sk[17]) & (g154) & (g1528)) + ((sk[17]) & (g154) & (g1528)));
	assign g1524 = (((!sk[18]) & (g1525) & (!g1526)) + ((!sk[18]) & (g1525) & (g1526)) + ((sk[18]) & (!g1525) & (!g1526)));
	assign g1525 = (((!sk[19]) & (g154) & (!g1529)) + ((!sk[19]) & (g154) & (g1529)) + ((sk[19]) & (!g154) & (g1529)));
	assign g1526 = (((g154) & (!sk[20]) & (!g1530)) + ((g154) & (!sk[20]) & (g1530)) + ((g154) & (sk[20]) & (g1530)));
	assign g1527 = (((!sk[21]) & (!g731) & (!g641) & (g339) & (!g640)) + ((!sk[21]) & (!g731) & (!g641) & (g339) & (g640)) + ((!sk[21]) & (!g731) & (g641) & (g339) & (!g640)) + ((!sk[21]) & (!g731) & (g641) & (g339) & (g640)) + ((!sk[21]) & (g731) & (!g641) & (g339) & (!g640)) + ((!sk[21]) & (g731) & (!g641) & (g339) & (g640)) + ((!sk[21]) & (g731) & (g641) & (g339) & (!g640)) + ((!sk[21]) & (g731) & (g641) & (g339) & (g640)) + ((sk[21]) & (g731) & (!g641) & (!g339) & (!g640)));
	assign g1528 = (((!g731) & (!g641) & (!sk[22]) & (g122) & (!g640)) + ((!g731) & (!g641) & (!sk[22]) & (g122) & (g640)) + ((!g731) & (g641) & (!sk[22]) & (g122) & (!g640)) + ((!g731) & (g641) & (!sk[22]) & (g122) & (g640)) + ((g731) & (!g641) & (!sk[22]) & (g122) & (!g640)) + ((g731) & (!g641) & (!sk[22]) & (g122) & (g640)) + ((g731) & (!g641) & (sk[22]) & (!g122) & (!g640)) + ((g731) & (!g641) & (sk[22]) & (!g122) & (g640)) + ((g731) & (!g641) & (sk[22]) & (g122) & (!g640)) + ((g731) & (g641) & (!sk[22]) & (g122) & (!g640)) + ((g731) & (g641) & (!sk[22]) & (g122) & (g640)) + ((g731) & (g641) & (sk[22]) & (!g122) & (!g640)) + ((g731) & (g641) & (sk[22]) & (!g122) & (g640)));
	assign g1529 = (((!g731) & (!sk[23]) & (!g641) & (g339) & (!g640)) + ((!g731) & (!sk[23]) & (!g641) & (g339) & (g640)) + ((!g731) & (!sk[23]) & (g641) & (g339) & (!g640)) + ((!g731) & (!sk[23]) & (g641) & (g339) & (g640)) + ((g731) & (!sk[23]) & (!g641) & (g339) & (!g640)) + ((g731) & (!sk[23]) & (!g641) & (g339) & (g640)) + ((g731) & (!sk[23]) & (g641) & (g339) & (!g640)) + ((g731) & (!sk[23]) & (g641) & (g339) & (g640)) + ((g731) & (sk[23]) & (!g641) & (!g339) & (!g640)));
	assign g1530 = (((!sk[24]) & (!g731) & (!g641) & (g122) & (!g640)) + ((!sk[24]) & (!g731) & (!g641) & (g122) & (g640)) + ((!sk[24]) & (!g731) & (g641) & (g122) & (!g640)) + ((!sk[24]) & (!g731) & (g641) & (g122) & (g640)) + ((!sk[24]) & (g731) & (!g641) & (g122) & (!g640)) + ((!sk[24]) & (g731) & (!g641) & (g122) & (g640)) + ((!sk[24]) & (g731) & (g641) & (g122) & (!g640)) + ((!sk[24]) & (g731) & (g641) & (g122) & (g640)) + ((sk[24]) & (g731) & (!g641) & (!g122) & (!g640)) + ((sk[24]) & (g731) & (!g641) & (g122) & (!g640)) + ((sk[24]) & (g731) & (g641) & (!g122) & (!g640)));
	assign g1531 = (((!sk[25]) & (g1532) & (!g1533)) + ((!sk[25]) & (g1532) & (g1533)) + ((sk[25]) & (!g1532) & (!g1533)));
	assign g1532 = (((!g634) & (sk[26]) & (g1534)) + ((g634) & (!sk[26]) & (!g1534)) + ((g634) & (!sk[26]) & (g1534)));
	assign g1533 = (((!sk[27]) & (g634) & (!g1537)) + ((!sk[27]) & (g634) & (g1537)) + ((sk[27]) & (g634) & (g1537)));
	assign g1534 = (((!sk[28]) & (g1535) & (!g1536)) + ((!sk[28]) & (g1535) & (g1536)) + ((sk[28]) & (!g1535) & (!g1536)));
	assign g1535 = (((!i_8_) & (sk[29]) & (!g73)) + ((i_8_) & (!sk[29]) & (!g73)) + ((i_8_) & (!sk[29]) & (g73)));
	assign g1536 = (((!sk[30]) & (i_8_) & (!g1540)) + ((!sk[30]) & (i_8_) & (g1540)) + ((sk[30]) & (i_8_) & (g1540)));
	assign g1537 = (((!sk[31]) & (g1538) & (!g1539)) + ((!sk[31]) & (g1538) & (g1539)) + ((sk[31]) & (!g1538) & (!g1539)));
	assign g1538 = (((!i_8_) & (sk[32]) & (g1541)) + ((i_8_) & (!sk[32]) & (!g1541)) + ((i_8_) & (!sk[32]) & (g1541)));
	assign g1539 = (((!sk[33]) & (i_8_) & (!g1542)) + ((!sk[33]) & (i_8_) & (g1542)) + ((sk[33]) & (i_8_) & (g1542)));
	assign g1540 = (((!g700) & (!sk[34]) & (!g699) & (g73)) + ((!g700) & (!sk[34]) & (g699) & (!g73)) + ((!g700) & (!sk[34]) & (g699) & (g73)) + ((!g700) & (sk[34]) & (!g699) & (!g73)) + ((!g700) & (sk[34]) & (g699) & (!g73)) + ((g700) & (!sk[34]) & (!g699) & (g73)) + ((g700) & (!sk[34]) & (g699) & (!g73)) + ((g700) & (!sk[34]) & (g699) & (g73)) + ((g700) & (sk[34]) & (!g699) & (!g73)) + ((g700) & (sk[34]) & (g699) & (!g73)) + ((g700) & (sk[34]) & (g699) & (g73)));
	assign g1541 = (((!sk[35]) & (!g701) & (!g700) & (g37) & (!g73)) + ((!sk[35]) & (!g701) & (!g700) & (g37) & (g73)) + ((!sk[35]) & (!g701) & (g700) & (g37) & (!g73)) + ((!sk[35]) & (!g701) & (g700) & (g37) & (g73)) + ((!sk[35]) & (g701) & (!g700) & (g37) & (!g73)) + ((!sk[35]) & (g701) & (!g700) & (g37) & (g73)) + ((!sk[35]) & (g701) & (g700) & (g37) & (!g73)) + ((!sk[35]) & (g701) & (g700) & (g37) & (g73)) + ((sk[35]) & (!g701) & (!g700) & (!g37) & (!g73)) + ((sk[35]) & (!g701) & (!g700) & (g37) & (!g73)) + ((sk[35]) & (!g701) & (g700) & (!g37) & (!g73)) + ((sk[35]) & (!g701) & (g700) & (g37) & (!g73)) + ((sk[35]) & (g701) & (!g700) & (!g37) & (!g73)) + ((sk[35]) & (g701) & (!g700) & (g37) & (!g73)) + ((sk[35]) & (g701) & (g700) & (!g37) & (!g73)) + ((sk[35]) & (g701) & (g700) & (g37) & (!g73)) + ((sk[35]) & (g701) & (g700) & (g37) & (g73)));
	assign g1542 = (((!g700) & (!g699) & (!sk[36]) & (g73)) + ((!g700) & (!g699) & (sk[36]) & (!g73)) + ((!g700) & (g699) & (!sk[36]) & (!g73)) + ((!g700) & (g699) & (!sk[36]) & (g73)) + ((!g700) & (g699) & (sk[36]) & (!g73)) + ((g700) & (!g699) & (!sk[36]) & (g73)) + ((g700) & (!g699) & (sk[36]) & (!g73)) + ((g700) & (g699) & (!sk[36]) & (!g73)) + ((g700) & (g699) & (!sk[36]) & (g73)) + ((g700) & (g699) & (sk[36]) & (!g73)) + ((g700) & (g699) & (sk[36]) & (g73)));
	assign g1543 = (((!sk[37]) & (g1544) & (!g1545)) + ((!sk[37]) & (g1544) & (g1545)) + ((sk[37]) & (!g1544) & (!g1545)));
	assign g1544 = (((!sk[38]) & (g102) & (!g1546)) + ((!sk[38]) & (g102) & (g1546)) + ((sk[38]) & (!g102) & (g1546)));
	assign g1545 = (((g102) & (!sk[39]) & (!g1549)) + ((g102) & (!sk[39]) & (g1549)) + ((g102) & (sk[39]) & (g1549)));
	assign g1546 = (((!sk[40]) & (g1547) & (!g1548)) + ((!sk[40]) & (g1547) & (g1548)) + ((sk[40]) & (!g1547) & (!g1548)));
	assign g1547 = (((!sk[41]) & (g22) & (!g556)) + ((!sk[41]) & (g22) & (g556)) + ((sk[41]) & (!g22) & (g556)));
	assign g1548 = (((!sk[42]) & (g22) & (!g556)) + ((!sk[42]) & (g22) & (g556)) + ((sk[42]) & (g22) & (g556)));
	assign g1549 = (((!sk[43]) & (g1550) & (!g1551)) + ((!sk[43]) & (g1550) & (g1551)) + ((sk[43]) & (!g1550) & (!g1551)));
	assign g1550 = (((!g22) & (sk[44]) & (g1552)) + ((g22) & (!sk[44]) & (!g1552)) + ((g22) & (!sk[44]) & (g1552)));
	assign g1551 = (((g22) & (!sk[45]) & (!g1553)) + ((g22) & (!sk[45]) & (g1553)) + ((g22) & (sk[45]) & (g1553)));
	assign g1552 = (((!g460) & (!sk[46]) & (!g76) & (g556)) + ((!g460) & (!sk[46]) & (g76) & (!g556)) + ((!g460) & (!sk[46]) & (g76) & (g556)) + ((g460) & (!sk[46]) & (!g76) & (g556)) + ((g460) & (!sk[46]) & (g76) & (!g556)) + ((g460) & (!sk[46]) & (g76) & (g556)) + ((g460) & (sk[46]) & (g76) & (g556)));
	assign g1553 = (((!g460) & (!sk[47]) & (!g91) & (g113) & (!g556)) + ((!g460) & (!sk[47]) & (!g91) & (g113) & (g556)) + ((!g460) & (!sk[47]) & (g91) & (g113) & (!g556)) + ((!g460) & (!sk[47]) & (g91) & (g113) & (g556)) + ((!g460) & (sk[47]) & (g91) & (g113) & (g556)) + ((g460) & (!sk[47]) & (!g91) & (g113) & (!g556)) + ((g460) & (!sk[47]) & (!g91) & (g113) & (g556)) + ((g460) & (!sk[47]) & (g91) & (g113) & (!g556)) + ((g460) & (!sk[47]) & (g91) & (g113) & (g556)) + ((g460) & (sk[47]) & (!g91) & (!g113) & (g556)) + ((g460) & (sk[47]) & (!g91) & (g113) & (g556)) + ((g460) & (sk[47]) & (g91) & (!g113) & (g556)) + ((g460) & (sk[47]) & (g91) & (g113) & (g556)));
	assign g1554 = (((!sk[48]) & (g1555) & (!g1556)) + ((!sk[48]) & (g1555) & (g1556)) + ((sk[48]) & (!g1555) & (!g1556)));
	assign g1555 = (((!sk[49]) & (g513) & (!g1557)) + ((!sk[49]) & (g513) & (g1557)) + ((sk[49]) & (!g513) & (g1557)));
	assign g1556 = (((g513) & (!sk[50]) & (!g1558)) + ((g513) & (!sk[50]) & (g1558)) + ((g513) & (sk[50]) & (g1558)));
	assign g1557 = (((!sk[51]) & (g122) & (!g1561)) + ((!sk[51]) & (g122) & (g1561)) + ((sk[51]) & (!g122) & (g1561)));
	assign g1558 = (((!sk[52]) & (g1559) & (!g1560)) + ((!sk[52]) & (g1559) & (g1560)) + ((sk[52]) & (!g1559) & (!g1560)));
	assign g1559 = (((!g122) & (sk[53]) & (g1562)) + ((g122) & (!sk[53]) & (!g1562)) + ((g122) & (!sk[53]) & (g1562)));
	assign g1560 = (((g122) & (!sk[54]) & (!g1563)) + ((g122) & (!sk[54]) & (g1563)) + ((g122) & (sk[54]) & (g1563)));
	assign g1561 = (((!g554) & (!g135) & (!sk[55]) & (g553)) + ((!g554) & (g135) & (!sk[55]) & (!g553)) + ((!g554) & (g135) & (!sk[55]) & (g553)) + ((g554) & (!g135) & (!sk[55]) & (g553)) + ((g554) & (g135) & (!sk[55]) & (!g553)) + ((g554) & (g135) & (!sk[55]) & (g553)) + ((g554) & (g135) & (sk[55]) & (g553)));
	assign g1562 = (((!sk[56]) & (g554) & (!g553)) + ((!sk[56]) & (g554) & (g553)) + ((sk[56]) & (g554) & (g553)));
	assign g1563 = (((!g552) & (!g554) & (g551) & (!sk[57]) & (!g553)) + ((!g552) & (!g554) & (g551) & (!sk[57]) & (g553)) + ((!g552) & (g554) & (g551) & (!sk[57]) & (!g553)) + ((!g552) & (g554) & (g551) & (!sk[57]) & (g553)) + ((g552) & (!g554) & (g551) & (!sk[57]) & (!g553)) + ((g552) & (!g554) & (g551) & (!sk[57]) & (g553)) + ((g552) & (g554) & (g551) & (!sk[57]) & (!g553)) + ((g552) & (g554) & (g551) & (!sk[57]) & (g553)) + ((g552) & (g554) & (g551) & (sk[57]) & (g553)));
	assign g1564 = (((!sk[58]) & (g1565) & (!g1566)) + ((!sk[58]) & (g1565) & (g1566)) + ((sk[58]) & (!g1565) & (!g1566)));
	assign g1565 = (((!g392) & (sk[59]) & (g1567)) + ((g392) & (!sk[59]) & (!g1567)) + ((g392) & (!sk[59]) & (g1567)));
	assign g1566 = (((g392) & (!sk[60]) & (!g1570)) + ((g392) & (!sk[60]) & (g1570)) + ((g392) & (sk[60]) & (g1570)));
	assign g1567 = (((!g1568) & (sk[61]) & (!g1569)) + ((g1568) & (!sk[61]) & (!g1569)) + ((g1568) & (!sk[61]) & (g1569)));
	assign g1568 = (((!i_15_) & (sk[62]) & (g1573)) + ((i_15_) & (!sk[62]) & (!g1573)) + ((i_15_) & (!sk[62]) & (g1573)));
	assign g1569 = (((!sk[63]) & (i_15_) & (!g1574)) + ((!sk[63]) & (i_15_) & (g1574)) + ((sk[63]) & (i_15_) & (g1574)));
	assign g1570 = (((!sk[64]) & (g1571) & (!g1572)) + ((!sk[64]) & (g1571) & (g1572)) + ((sk[64]) & (!g1571) & (!g1572)));
	assign g1571 = (((!sk[65]) & (i_15_) & (!g1575)) + ((!sk[65]) & (i_15_) & (g1575)) + ((sk[65]) & (!i_15_) & (g1575)));
	assign g1572 = (((!sk[66]) & (i_15_) & (!g1576)) + ((!sk[66]) & (i_15_) & (g1576)) + ((sk[66]) & (i_15_) & (g1576)));
	assign g1573 = (((!g174) & (!g428) & (g142) & (!sk[67]) & (!g524)) + ((!g174) & (!g428) & (g142) & (!sk[67]) & (g524)) + ((!g174) & (!g428) & (g142) & (sk[67]) & (g524)) + ((!g174) & (g428) & (!g142) & (sk[67]) & (g524)) + ((!g174) & (g428) & (g142) & (!sk[67]) & (!g524)) + ((!g174) & (g428) & (g142) & (!sk[67]) & (g524)) + ((!g174) & (g428) & (g142) & (sk[67]) & (g524)) + ((g174) & (!g428) & (!g142) & (sk[67]) & (g524)) + ((g174) & (!g428) & (g142) & (!sk[67]) & (!g524)) + ((g174) & (!g428) & (g142) & (!sk[67]) & (g524)) + ((g174) & (!g428) & (g142) & (sk[67]) & (g524)) + ((g174) & (g428) & (!g142) & (sk[67]) & (g524)) + ((g174) & (g428) & (g142) & (!sk[67]) & (!g524)) + ((g174) & (g428) & (g142) & (!sk[67]) & (g524)) + ((g174) & (g428) & (g142) & (sk[67]) & (g524)));
	assign g1574 = (((!sk[68]) & (!g174) & (!g520) & (g524)) + ((!sk[68]) & (!g174) & (g520) & (!g524)) + ((!sk[68]) & (!g174) & (g520) & (g524)) + ((!sk[68]) & (g174) & (!g520) & (g524)) + ((!sk[68]) & (g174) & (g520) & (!g524)) + ((!sk[68]) & (g174) & (g520) & (g524)) + ((sk[68]) & (!g174) & (g520) & (g524)) + ((sk[68]) & (g174) & (!g520) & (g524)) + ((sk[68]) & (g174) & (g520) & (g524)));
	assign g1575 = (((!sk[69]) & (!g174) & (!g428) & (g524)) + ((!sk[69]) & (!g174) & (g428) & (!g524)) + ((!sk[69]) & (!g174) & (g428) & (g524)) + ((!sk[69]) & (g174) & (!g428) & (g524)) + ((!sk[69]) & (g174) & (g428) & (!g524)) + ((!sk[69]) & (g174) & (g428) & (g524)) + ((sk[69]) & (!g174) & (g428) & (g524)) + ((sk[69]) & (g174) & (!g428) & (g524)) + ((sk[69]) & (g174) & (g428) & (g524)));
	assign g1576 = (((!g174) & (!sk[70]) & (!g520) & (g524)) + ((!g174) & (!sk[70]) & (g520) & (!g524)) + ((!g174) & (!sk[70]) & (g520) & (g524)) + ((!g174) & (sk[70]) & (g520) & (g524)) + ((g174) & (!sk[70]) & (!g520) & (g524)) + ((g174) & (!sk[70]) & (g520) & (!g524)) + ((g174) & (!sk[70]) & (g520) & (g524)) + ((g174) & (sk[70]) & (!g520) & (g524)) + ((g174) & (sk[70]) & (g520) & (g524)));
	assign g1577 = (((!sk[71]) & (g174) & (!g1578)) + ((!sk[71]) & (g174) & (g1578)) + ((sk[71]) & (!g174) & (!g1578)));
	assign g1578 = (((!g174) & (sk[72]) & (g1579)) + ((g174) & (!sk[72]) & (!g1579)) + ((g174) & (!sk[72]) & (g1579)));
	assign g1579 = (((!g1580) & (sk[73]) & (!g1581)) + ((g1580) & (!sk[73]) & (!g1581)) + ((g1580) & (!sk[73]) & (g1581)));
	assign g1580 = (((!i_9_) & (sk[74]) & (g1582)) + ((i_9_) & (!sk[74]) & (!g1582)) + ((i_9_) & (!sk[74]) & (g1582)));
	assign g1581 = (((i_9_) & (!sk[75]) & (!g1583)) + ((i_9_) & (!sk[75]) & (g1583)) + ((i_9_) & (sk[75]) & (g1583)));
	assign g1582 = (((!i_15_) & (!i_11_) & (!g262) & (sk[76]) & (!i_10_)) + ((!i_15_) & (!i_11_) & (!g262) & (sk[76]) & (i_10_)) + ((!i_15_) & (!i_11_) & (g262) & (!sk[76]) & (!i_10_)) + ((!i_15_) & (!i_11_) & (g262) & (!sk[76]) & (i_10_)) + ((!i_15_) & (!i_11_) & (g262) & (sk[76]) & (!i_10_)) + ((!i_15_) & (!i_11_) & (g262) & (sk[76]) & (i_10_)) + ((!i_15_) & (i_11_) & (!g262) & (sk[76]) & (!i_10_)) + ((!i_15_) & (i_11_) & (!g262) & (sk[76]) & (i_10_)) + ((!i_15_) & (i_11_) & (g262) & (!sk[76]) & (!i_10_)) + ((!i_15_) & (i_11_) & (g262) & (!sk[76]) & (i_10_)) + ((!i_15_) & (i_11_) & (g262) & (sk[76]) & (i_10_)) + ((i_15_) & (!i_11_) & (!g262) & (sk[76]) & (!i_10_)) + ((i_15_) & (!i_11_) & (!g262) & (sk[76]) & (i_10_)) + ((i_15_) & (!i_11_) & (g262) & (!sk[76]) & (!i_10_)) + ((i_15_) & (!i_11_) & (g262) & (!sk[76]) & (i_10_)) + ((i_15_) & (!i_11_) & (g262) & (sk[76]) & (!i_10_)) + ((i_15_) & (!i_11_) & (g262) & (sk[76]) & (i_10_)) + ((i_15_) & (i_11_) & (!g262) & (sk[76]) & (!i_10_)) + ((i_15_) & (i_11_) & (!g262) & (sk[76]) & (i_10_)) + ((i_15_) & (i_11_) & (g262) & (!sk[76]) & (!i_10_)) + ((i_15_) & (i_11_) & (g262) & (!sk[76]) & (i_10_)) + ((i_15_) & (i_11_) & (g262) & (sk[76]) & (!i_10_)) + ((i_15_) & (i_11_) & (g262) & (sk[76]) & (i_10_)));
	assign g1583 = (((!sk[77]) & (!i_15_) & (!i_11_) & (g518) & (!i_10_)) + ((!sk[77]) & (!i_15_) & (!i_11_) & (g518) & (i_10_)) + ((!sk[77]) & (!i_15_) & (i_11_) & (g518) & (!i_10_)) + ((!sk[77]) & (!i_15_) & (i_11_) & (g518) & (i_10_)) + ((!sk[77]) & (i_15_) & (!i_11_) & (g518) & (!i_10_)) + ((!sk[77]) & (i_15_) & (!i_11_) & (g518) & (i_10_)) + ((!sk[77]) & (i_15_) & (i_11_) & (g518) & (!i_10_)) + ((!sk[77]) & (i_15_) & (i_11_) & (g518) & (i_10_)) + ((sk[77]) & (!i_15_) & (!i_11_) & (!g518) & (!i_10_)) + ((sk[77]) & (!i_15_) & (!i_11_) & (!g518) & (i_10_)) + ((sk[77]) & (!i_15_) & (!i_11_) & (g518) & (!i_10_)) + ((sk[77]) & (!i_15_) & (!i_11_) & (g518) & (i_10_)) + ((sk[77]) & (!i_15_) & (i_11_) & (!g518) & (!i_10_)) + ((sk[77]) & (!i_15_) & (i_11_) & (!g518) & (i_10_)) + ((sk[77]) & (!i_15_) & (i_11_) & (g518) & (i_10_)) + ((sk[77]) & (i_15_) & (!i_11_) & (!g518) & (!i_10_)) + ((sk[77]) & (i_15_) & (!i_11_) & (!g518) & (i_10_)) + ((sk[77]) & (i_15_) & (!i_11_) & (g518) & (!i_10_)) + ((sk[77]) & (i_15_) & (!i_11_) & (g518) & (i_10_)) + ((sk[77]) & (i_15_) & (i_11_) & (!g518) & (!i_10_)) + ((sk[77]) & (i_15_) & (i_11_) & (!g518) & (i_10_)) + ((sk[77]) & (i_15_) & (i_11_) & (g518) & (!i_10_)) + ((sk[77]) & (i_15_) & (i_11_) & (g518) & (i_10_)));
	assign g1584 = (((!g1585) & (sk[78]) & (!g1586)) + ((g1585) & (!sk[78]) & (!g1586)) + ((g1585) & (!sk[78]) & (g1586)));
	assign g1585 = (((!sk[79]) & (i_15_) & (!g1587)) + ((!sk[79]) & (i_15_) & (g1587)) + ((sk[79]) & (!i_15_) & (g1587)));
	assign g1586 = (((!sk[80]) & (i_15_) & (!g1589)) + ((!sk[80]) & (i_15_) & (g1589)) + ((sk[80]) & (i_15_) & (g1589)));
	assign g1587 = (((!sk[81]) & (i_11_) & (!g1588)) + ((!sk[81]) & (i_11_) & (g1588)) + ((sk[81]) & (i_11_) & (!g1588)));
	assign g1588 = (((!sk[82]) & (i_11_) & (!g1591)) + ((!sk[82]) & (i_11_) & (g1591)) + ((sk[82]) & (i_11_) & (g1591)));
	assign g1589 = (((!i_11_) & (sk[83]) & (!g1590)) + ((i_11_) & (!sk[83]) & (!g1590)) + ((i_11_) & (!sk[83]) & (g1590)));
	assign g1590 = (((!i_11_) & (sk[84]) & (g1592)) + ((i_11_) & (!sk[84]) & (!g1592)) + ((i_11_) & (!sk[84]) & (g1592)));
	assign g1591 = (((!g176) & (!sk[85]) & (!i_10_) & (g443) & (!i_9_)) + ((!g176) & (!sk[85]) & (!i_10_) & (g443) & (i_9_)) + ((!g176) & (!sk[85]) & (i_10_) & (g443) & (!i_9_)) + ((!g176) & (!sk[85]) & (i_10_) & (g443) & (i_9_)) + ((!g176) & (sk[85]) & (!i_10_) & (!g443) & (!i_9_)) + ((!g176) & (sk[85]) & (!i_10_) & (!g443) & (i_9_)) + ((!g176) & (sk[85]) & (!i_10_) & (g443) & (!i_9_)) + ((!g176) & (sk[85]) & (!i_10_) & (g443) & (i_9_)) + ((!g176) & (sk[85]) & (i_10_) & (!g443) & (i_9_)) + ((!g176) & (sk[85]) & (i_10_) & (g443) & (!i_9_)) + ((!g176) & (sk[85]) & (i_10_) & (g443) & (i_9_)) + ((g176) & (!sk[85]) & (!i_10_) & (g443) & (!i_9_)) + ((g176) & (!sk[85]) & (!i_10_) & (g443) & (i_9_)) + ((g176) & (!sk[85]) & (i_10_) & (g443) & (!i_9_)) + ((g176) & (!sk[85]) & (i_10_) & (g443) & (i_9_)) + ((g176) & (sk[85]) & (!i_10_) & (!g443) & (!i_9_)) + ((g176) & (sk[85]) & (!i_10_) & (!g443) & (i_9_)) + ((g176) & (sk[85]) & (!i_10_) & (g443) & (!i_9_)) + ((g176) & (sk[85]) & (!i_10_) & (g443) & (i_9_)) + ((g176) & (sk[85]) & (i_10_) & (!g443) & (!i_9_)) + ((g176) & (sk[85]) & (i_10_) & (!g443) & (i_9_)) + ((g176) & (sk[85]) & (i_10_) & (g443) & (!i_9_)) + ((g176) & (sk[85]) & (i_10_) & (g443) & (i_9_)));
	assign g1592 = (((!g176) & (!sk[86]) & (!i_10_) & (g444) & (!i_9_)) + ((!g176) & (!sk[86]) & (!i_10_) & (g444) & (i_9_)) + ((!g176) & (!sk[86]) & (i_10_) & (g444) & (!i_9_)) + ((!g176) & (!sk[86]) & (i_10_) & (g444) & (i_9_)) + ((!g176) & (sk[86]) & (!i_10_) & (!g444) & (!i_9_)) + ((!g176) & (sk[86]) & (!i_10_) & (!g444) & (i_9_)) + ((!g176) & (sk[86]) & (!i_10_) & (g444) & (!i_9_)) + ((!g176) & (sk[86]) & (!i_10_) & (g444) & (i_9_)) + ((!g176) & (sk[86]) & (i_10_) & (!g444) & (i_9_)) + ((!g176) & (sk[86]) & (i_10_) & (g444) & (!i_9_)) + ((!g176) & (sk[86]) & (i_10_) & (g444) & (i_9_)) + ((g176) & (!sk[86]) & (!i_10_) & (g444) & (!i_9_)) + ((g176) & (!sk[86]) & (!i_10_) & (g444) & (i_9_)) + ((g176) & (!sk[86]) & (i_10_) & (g444) & (!i_9_)) + ((g176) & (!sk[86]) & (i_10_) & (g444) & (i_9_)) + ((g176) & (sk[86]) & (!i_10_) & (!g444) & (!i_9_)) + ((g176) & (sk[86]) & (!i_10_) & (!g444) & (i_9_)) + ((g176) & (sk[86]) & (!i_10_) & (g444) & (!i_9_)) + ((g176) & (sk[86]) & (!i_10_) & (g444) & (i_9_)) + ((g176) & (sk[86]) & (i_10_) & (!g444) & (!i_9_)) + ((g176) & (sk[86]) & (i_10_) & (!g444) & (i_9_)) + ((g176) & (sk[86]) & (i_10_) & (g444) & (!i_9_)) + ((g176) & (sk[86]) & (i_10_) & (g444) & (i_9_)));
	assign g1593 = (((!sk[87]) & (g1594) & (!g1595)) + ((!sk[87]) & (g1594) & (g1595)) + ((sk[87]) & (!g1594) & (!g1595)));
	assign g1594 = (((!sk[88]) & (g78) & (!g1596)) + ((!sk[88]) & (g78) & (g1596)) + ((sk[88]) & (!g78) & (g1596)));
	assign g1595 = (((g78) & (!sk[89]) & (!g1599)) + ((g78) & (!sk[89]) & (g1599)) + ((g78) & (sk[89]) & (g1599)));
	assign g1596 = (((!sk[90]) & (g1597) & (!g1598)) + ((!sk[90]) & (g1597) & (g1598)) + ((sk[90]) & (!g1597) & (!g1598)));
	assign g1597 = (((!sk[91]) & (g97) & (!g1602)) + ((!sk[91]) & (g97) & (g1602)) + ((sk[91]) & (!g97) & (g1602)));
	assign g1598 = (((g97) & (!sk[92]) & (!g1603)) + ((g97) & (!sk[92]) & (g1603)) + ((g97) & (sk[92]) & (g1603)));
	assign g1599 = (((!g1600) & (sk[93]) & (!g1601)) + ((g1600) & (!sk[93]) & (!g1601)) + ((g1600) & (!sk[93]) & (g1601)));
	assign g1600 = (((!g97) & (sk[94]) & (g1604)) + ((g97) & (!sk[94]) & (!g1604)) + ((g97) & (!sk[94]) & (g1604)));
	assign g1601 = (((g97) & (!sk[95]) & (!g1605)) + ((g97) & (!sk[95]) & (g1605)) + ((g97) & (sk[95]) & (g1605)));
	assign g1602 = (((!g144) & (!sk[96]) & (!g425) & (g226) & (!g142)) + ((!g144) & (!sk[96]) & (!g425) & (g226) & (g142)) + ((!g144) & (!sk[96]) & (g425) & (g226) & (!g142)) + ((!g144) & (!sk[96]) & (g425) & (g226) & (g142)) + ((!g144) & (sk[96]) & (g425) & (g226) & (g142)) + ((g144) & (!sk[96]) & (!g425) & (g226) & (!g142)) + ((g144) & (!sk[96]) & (!g425) & (g226) & (g142)) + ((g144) & (!sk[96]) & (g425) & (g226) & (!g142)) + ((g144) & (!sk[96]) & (g425) & (g226) & (g142)));
	assign g1603 = (((!g144) & (!g425) & (g114) & (!sk[97]) & (!g142)) + ((!g144) & (!g425) & (g114) & (!sk[97]) & (g142)) + ((!g144) & (g425) & (!g114) & (sk[97]) & (g142)) + ((!g144) & (g425) & (g114) & (!sk[97]) & (!g142)) + ((!g144) & (g425) & (g114) & (!sk[97]) & (g142)) + ((!g144) & (g425) & (g114) & (sk[97]) & (g142)) + ((g144) & (!g425) & (g114) & (!sk[97]) & (!g142)) + ((g144) & (!g425) & (g114) & (!sk[97]) & (g142)) + ((g144) & (g425) & (g114) & (!sk[97]) & (!g142)) + ((g144) & (g425) & (g114) & (!sk[97]) & (g142)) + ((g144) & (g425) & (g114) & (sk[97]) & (g142)));
	assign g1604 = (((!g144) & (!sk[98]) & (!g425) & (g226)) + ((!g144) & (!sk[98]) & (g425) & (!g226)) + ((!g144) & (!sk[98]) & (g425) & (g226)) + ((!g144) & (sk[98]) & (g425) & (g226)) + ((g144) & (!sk[98]) & (!g425) & (g226)) + ((g144) & (!sk[98]) & (g425) & (!g226)) + ((g144) & (!sk[98]) & (g425) & (g226)));
	assign g1605 = (((!g144) & (!sk[99]) & (!g425) & (g114)) + ((!g144) & (!sk[99]) & (g425) & (!g114)) + ((!g144) & (!sk[99]) & (g425) & (g114)) + ((!g144) & (sk[99]) & (!g425) & (g114)) + ((!g144) & (sk[99]) & (g425) & (!g114)) + ((!g144) & (sk[99]) & (g425) & (g114)) + ((g144) & (!sk[99]) & (!g425) & (g114)) + ((g144) & (!sk[99]) & (g425) & (!g114)) + ((g144) & (!sk[99]) & (g425) & (g114)) + ((g144) & (sk[99]) & (!g425) & (g114)) + ((g144) & (sk[99]) & (g425) & (g114)));
	assign g1606 = (((!g24) & (sk[100]) & (!g1607)) + ((g24) & (!sk[100]) & (!g1607)) + ((g24) & (!sk[100]) & (g1607)));
	assign g1607 = (((!g24) & (sk[101]) & (g1608)) + ((g24) & (!sk[101]) & (!g1608)) + ((g24) & (!sk[101]) & (g1608)));
	assign g1608 = (((!sk[102]) & (g1609) & (!g1610)) + ((!sk[102]) & (g1609) & (g1610)) + ((sk[102]) & (!g1609) & (!g1610)));
	assign g1609 = (((!sk[103]) & (i_11_) & (!g1611)) + ((!sk[103]) & (i_11_) & (g1611)) + ((sk[103]) & (!i_11_) & (g1611)));
	assign g1610 = (((!sk[104]) & (i_11_) & (!g1612)) + ((!sk[104]) & (i_11_) & (g1612)) + ((sk[104]) & (i_11_) & (g1612)));
	assign g1611 = (((!i_15_) & (!sk[105]) & (!i_10_) & (g144) & (!i_9_)) + ((!i_15_) & (!sk[105]) & (!i_10_) & (g144) & (i_9_)) + ((!i_15_) & (!sk[105]) & (i_10_) & (g144) & (!i_9_)) + ((!i_15_) & (!sk[105]) & (i_10_) & (g144) & (i_9_)) + ((!i_15_) & (sk[105]) & (!i_10_) & (!g144) & (!i_9_)) + ((!i_15_) & (sk[105]) & (!i_10_) & (!g144) & (i_9_)) + ((!i_15_) & (sk[105]) & (!i_10_) & (g144) & (!i_9_)) + ((!i_15_) & (sk[105]) & (i_10_) & (!g144) & (!i_9_)) + ((!i_15_) & (sk[105]) & (i_10_) & (!g144) & (i_9_)) + ((!i_15_) & (sk[105]) & (i_10_) & (g144) & (!i_9_)) + ((!i_15_) & (sk[105]) & (i_10_) & (g144) & (i_9_)) + ((i_15_) & (!sk[105]) & (!i_10_) & (g144) & (!i_9_)) + ((i_15_) & (!sk[105]) & (!i_10_) & (g144) & (i_9_)) + ((i_15_) & (!sk[105]) & (i_10_) & (g144) & (!i_9_)) + ((i_15_) & (!sk[105]) & (i_10_) & (g144) & (i_9_)) + ((i_15_) & (sk[105]) & (!i_10_) & (!g144) & (!i_9_)) + ((i_15_) & (sk[105]) & (!i_10_) & (!g144) & (i_9_)) + ((i_15_) & (sk[105]) & (!i_10_) & (g144) & (!i_9_)) + ((i_15_) & (sk[105]) & (!i_10_) & (g144) & (i_9_)) + ((i_15_) & (sk[105]) & (i_10_) & (!g144) & (!i_9_)) + ((i_15_) & (sk[105]) & (i_10_) & (!g144) & (i_9_)) + ((i_15_) & (sk[105]) & (i_10_) & (g144) & (!i_9_)) + ((i_15_) & (sk[105]) & (i_10_) & (g144) & (i_9_)));
	assign g1612 = (((!i_15_) & (!sk[106]) & (!i_10_) & (g165) & (!i_9_)) + ((!i_15_) & (!sk[106]) & (!i_10_) & (g165) & (i_9_)) + ((!i_15_) & (!sk[106]) & (i_10_) & (g165) & (!i_9_)) + ((!i_15_) & (!sk[106]) & (i_10_) & (g165) & (i_9_)) + ((!i_15_) & (sk[106]) & (!i_10_) & (!g165) & (!i_9_)) + ((!i_15_) & (sk[106]) & (!i_10_) & (!g165) & (i_9_)) + ((!i_15_) & (sk[106]) & (!i_10_) & (g165) & (!i_9_)) + ((!i_15_) & (sk[106]) & (i_10_) & (!g165) & (!i_9_)) + ((!i_15_) & (sk[106]) & (i_10_) & (!g165) & (i_9_)) + ((!i_15_) & (sk[106]) & (i_10_) & (g165) & (!i_9_)) + ((!i_15_) & (sk[106]) & (i_10_) & (g165) & (i_9_)) + ((i_15_) & (!sk[106]) & (!i_10_) & (g165) & (!i_9_)) + ((i_15_) & (!sk[106]) & (!i_10_) & (g165) & (i_9_)) + ((i_15_) & (!sk[106]) & (i_10_) & (g165) & (!i_9_)) + ((i_15_) & (!sk[106]) & (i_10_) & (g165) & (i_9_)) + ((i_15_) & (sk[106]) & (!i_10_) & (!g165) & (!i_9_)) + ((i_15_) & (sk[106]) & (!i_10_) & (!g165) & (i_9_)) + ((i_15_) & (sk[106]) & (!i_10_) & (g165) & (!i_9_)) + ((i_15_) & (sk[106]) & (!i_10_) & (g165) & (i_9_)) + ((i_15_) & (sk[106]) & (i_10_) & (!g165) & (!i_9_)) + ((i_15_) & (sk[106]) & (i_10_) & (!g165) & (i_9_)) + ((i_15_) & (sk[106]) & (i_10_) & (g165) & (!i_9_)) + ((i_15_) & (sk[106]) & (i_10_) & (g165) & (i_9_)));
	assign g1613 = (((!sk[107]) & (g1614) & (!g1615)) + ((!sk[107]) & (g1614) & (g1615)) + ((sk[107]) & (!g1614) & (!g1615)));
	assign g1614 = (((!g102) & (sk[108]) & (g1616)) + ((g102) & (!sk[108]) & (!g1616)) + ((g102) & (!sk[108]) & (g1616)));
	assign g1615 = (((!sk[109]) & (g102) & (!g1619)) + ((!sk[109]) & (g102) & (g1619)) + ((sk[109]) & (g102) & (g1619)));
	assign g1616 = (((!g1617) & (sk[110]) & (!g1618)) + ((g1617) & (!sk[110]) & (!g1618)) + ((g1617) & (!sk[110]) & (g1618)));
	assign g1617 = (((!g155) & (sk[111]) & (g1622)) + ((g155) & (!sk[111]) & (!g1622)) + ((g155) & (!sk[111]) & (g1622)));
	assign g1618 = (((!sk[112]) & (g155) & (!g1623)) + ((!sk[112]) & (g155) & (g1623)) + ((sk[112]) & (g155) & (g1623)));
	assign g1619 = (((!sk[113]) & (g1620) & (!g1621)) + ((!sk[113]) & (g1620) & (g1621)) + ((sk[113]) & (!g1620) & (!g1621)));
	assign g1620 = (((!sk[114]) & (g155) & (!g323)) + ((!sk[114]) & (g155) & (g323)) + ((sk[114]) & (!g155) & (g323)));
	assign g1621 = (((g155) & (!sk[115]) & (!g1624)) + ((g155) & (!sk[115]) & (g1624)) + ((g155) & (sk[115]) & (g1624)));
	assign g1622 = (((!g24) & (!sk[116]) & (!g323) & (g107) & (!g254)) + ((!g24) & (!sk[116]) & (!g323) & (g107) & (g254)) + ((!g24) & (!sk[116]) & (g323) & (g107) & (!g254)) + ((!g24) & (!sk[116]) & (g323) & (g107) & (g254)) + ((!g24) & (sk[116]) & (!g323) & (g107) & (g254)) + ((!g24) & (sk[116]) & (g323) & (!g107) & (!g254)) + ((!g24) & (sk[116]) & (g323) & (!g107) & (g254)) + ((!g24) & (sk[116]) & (g323) & (g107) & (!g254)) + ((!g24) & (sk[116]) & (g323) & (g107) & (g254)) + ((g24) & (!sk[116]) & (!g323) & (g107) & (!g254)) + ((g24) & (!sk[116]) & (!g323) & (g107) & (g254)) + ((g24) & (!sk[116]) & (g323) & (g107) & (!g254)) + ((g24) & (!sk[116]) & (g323) & (g107) & (g254)) + ((g24) & (sk[116]) & (!g323) & (!g107) & (g254)) + ((g24) & (sk[116]) & (!g323) & (g107) & (g254)) + ((g24) & (sk[116]) & (g323) & (!g107) & (!g254)) + ((g24) & (sk[116]) & (g323) & (!g107) & (g254)) + ((g24) & (sk[116]) & (g323) & (g107) & (!g254)) + ((g24) & (sk[116]) & (g323) & (g107) & (g254)));
	assign g1623 = (((!sk[117]) & (!g24) & (!g323) & (g126) & (!g254)) + ((!sk[117]) & (!g24) & (!g323) & (g126) & (g254)) + ((!sk[117]) & (!g24) & (g323) & (g126) & (!g254)) + ((!sk[117]) & (!g24) & (g323) & (g126) & (g254)) + ((!sk[117]) & (g24) & (!g323) & (g126) & (!g254)) + ((!sk[117]) & (g24) & (!g323) & (g126) & (g254)) + ((!sk[117]) & (g24) & (g323) & (g126) & (!g254)) + ((!sk[117]) & (g24) & (g323) & (g126) & (g254)) + ((sk[117]) & (!g24) & (!g323) & (!g126) & (g254)) + ((sk[117]) & (!g24) & (!g323) & (g126) & (!g254)) + ((sk[117]) & (!g24) & (!g323) & (g126) & (g254)) + ((sk[117]) & (!g24) & (g323) & (!g126) & (!g254)) + ((sk[117]) & (!g24) & (g323) & (!g126) & (g254)) + ((sk[117]) & (!g24) & (g323) & (g126) & (!g254)) + ((sk[117]) & (!g24) & (g323) & (g126) & (g254)) + ((sk[117]) & (g24) & (!g323) & (!g126) & (!g254)) + ((sk[117]) & (g24) & (!g323) & (!g126) & (g254)) + ((sk[117]) & (g24) & (!g323) & (g126) & (!g254)) + ((sk[117]) & (g24) & (!g323) & (g126) & (g254)) + ((sk[117]) & (g24) & (g323) & (!g126) & (!g254)) + ((sk[117]) & (g24) & (g323) & (!g126) & (g254)) + ((sk[117]) & (g24) & (g323) & (g126) & (!g254)) + ((sk[117]) & (g24) & (g323) & (g126) & (g254)));
	assign g1624 = (((!g24) & (!sk[118]) & (!g323) & (g126)) + ((!g24) & (!sk[118]) & (g323) & (!g126)) + ((!g24) & (!sk[118]) & (g323) & (g126)) + ((!g24) & (sk[118]) & (!g323) & (g126)) + ((!g24) & (sk[118]) & (g323) & (!g126)) + ((!g24) & (sk[118]) & (g323) & (g126)) + ((g24) & (!sk[118]) & (!g323) & (g126)) + ((g24) & (!sk[118]) & (g323) & (!g126)) + ((g24) & (!sk[118]) & (g323) & (g126)) + ((g24) & (sk[118]) & (!g323) & (!g126)) + ((g24) & (sk[118]) & (!g323) & (g126)) + ((g24) & (sk[118]) & (g323) & (!g126)) + ((g24) & (sk[118]) & (g323) & (g126)));
	assign g1625 = (((!g68) & (sk[119]) & (!g1626)) + ((g68) & (!sk[119]) & (!g1626)) + ((g68) & (!sk[119]) & (g1626)));
	assign g1626 = (((!g68) & (sk[120]) & (g1627)) + ((g68) & (!sk[120]) & (!g1627)) + ((g68) & (!sk[120]) & (g1627)));
	assign g1627 = (((!g1628) & (sk[121]) & (!g1629)) + ((g1628) & (!sk[121]) & (!g1629)) + ((g1628) & (!sk[121]) & (g1629)));
	assign g1628 = (((!sk[122]) & (i_11_) & (!g1630)) + ((!sk[122]) & (i_11_) & (g1630)) + ((sk[122]) & (!i_11_) & (g1630)));
	assign g1629 = (((!sk[123]) & (i_11_) & (!g1631)) + ((!sk[123]) & (i_11_) & (g1631)) + ((sk[123]) & (i_11_) & (g1631)));
	assign g1630 = (((!sk[124]) & (!i_15_) & (!i_10_) & (g157) & (!i_9_)) + ((!sk[124]) & (!i_15_) & (!i_10_) & (g157) & (i_9_)) + ((!sk[124]) & (!i_15_) & (i_10_) & (g157) & (!i_9_)) + ((!sk[124]) & (!i_15_) & (i_10_) & (g157) & (i_9_)) + ((!sk[124]) & (i_15_) & (!i_10_) & (g157) & (!i_9_)) + ((!sk[124]) & (i_15_) & (!i_10_) & (g157) & (i_9_)) + ((!sk[124]) & (i_15_) & (i_10_) & (g157) & (!i_9_)) + ((!sk[124]) & (i_15_) & (i_10_) & (g157) & (i_9_)) + ((sk[124]) & (!i_15_) & (!i_10_) & (!g157) & (!i_9_)) + ((sk[124]) & (!i_15_) & (!i_10_) & (!g157) & (i_9_)) + ((sk[124]) & (!i_15_) & (!i_10_) & (g157) & (!i_9_)) + ((sk[124]) & (!i_15_) & (!i_10_) & (g157) & (i_9_)) + ((sk[124]) & (!i_15_) & (i_10_) & (!g157) & (!i_9_)) + ((sk[124]) & (!i_15_) & (i_10_) & (!g157) & (i_9_)) + ((sk[124]) & (!i_15_) & (i_10_) & (g157) & (!i_9_)) + ((sk[124]) & (i_15_) & (!i_10_) & (!g157) & (!i_9_)) + ((sk[124]) & (i_15_) & (!i_10_) & (!g157) & (i_9_)) + ((sk[124]) & (i_15_) & (!i_10_) & (g157) & (!i_9_)) + ((sk[124]) & (i_15_) & (!i_10_) & (g157) & (i_9_)) + ((sk[124]) & (i_15_) & (i_10_) & (!g157) & (!i_9_)) + ((sk[124]) & (i_15_) & (i_10_) & (!g157) & (i_9_)) + ((sk[124]) & (i_15_) & (i_10_) & (g157) & (!i_9_)) + ((sk[124]) & (i_15_) & (i_10_) & (g157) & (i_9_)));
	assign g1631 = (((!i_15_) & (!sk[125]) & (!i_10_) & (g254) & (!i_9_)) + ((!i_15_) & (!sk[125]) & (!i_10_) & (g254) & (i_9_)) + ((!i_15_) & (!sk[125]) & (i_10_) & (g254) & (!i_9_)) + ((!i_15_) & (!sk[125]) & (i_10_) & (g254) & (i_9_)) + ((!i_15_) & (sk[125]) & (!i_10_) & (!g254) & (!i_9_)) + ((!i_15_) & (sk[125]) & (!i_10_) & (!g254) & (i_9_)) + ((!i_15_) & (sk[125]) & (!i_10_) & (g254) & (!i_9_)) + ((!i_15_) & (sk[125]) & (!i_10_) & (g254) & (i_9_)) + ((!i_15_) & (sk[125]) & (i_10_) & (!g254) & (i_9_)) + ((!i_15_) & (sk[125]) & (i_10_) & (g254) & (!i_9_)) + ((!i_15_) & (sk[125]) & (i_10_) & (g254) & (i_9_)) + ((i_15_) & (!sk[125]) & (!i_10_) & (g254) & (!i_9_)) + ((i_15_) & (!sk[125]) & (!i_10_) & (g254) & (i_9_)) + ((i_15_) & (!sk[125]) & (i_10_) & (g254) & (!i_9_)) + ((i_15_) & (!sk[125]) & (i_10_) & (g254) & (i_9_)) + ((i_15_) & (sk[125]) & (!i_10_) & (!g254) & (!i_9_)) + ((i_15_) & (sk[125]) & (!i_10_) & (!g254) & (i_9_)) + ((i_15_) & (sk[125]) & (!i_10_) & (g254) & (!i_9_)) + ((i_15_) & (sk[125]) & (!i_10_) & (g254) & (i_9_)) + ((i_15_) & (sk[125]) & (i_10_) & (!g254) & (!i_9_)) + ((i_15_) & (sk[125]) & (i_10_) & (!g254) & (i_9_)) + ((i_15_) & (sk[125]) & (i_10_) & (g254) & (!i_9_)) + ((i_15_) & (sk[125]) & (i_10_) & (g254) & (i_9_)));
	assign g1632 = (((!sk[126]) & (g68) & (!g1633)) + ((!sk[126]) & (g68) & (g1633)) + ((sk[126]) & (!g68) & (!g1633)));
	assign g1633 = (((!g68) & (sk[127]) & (g1634)) + ((g68) & (!sk[127]) & (!g1634)) + ((g68) & (!sk[127]) & (g1634)));
	assign g1634 = (((!g1635) & (sk[0]) & (!g1636)) + ((g1635) & (!sk[0]) & (!g1636)) + ((g1635) & (!sk[0]) & (g1636)));
	assign g1635 = (((!sk[1]) & (i_11_) & (!g1637)) + ((!sk[1]) & (i_11_) & (g1637)) + ((sk[1]) & (!i_11_) & (g1637)));
	assign g1636 = (((!sk[2]) & (i_11_) & (!g1638)) + ((!sk[2]) & (i_11_) & (g1638)) + ((sk[2]) & (i_11_) & (g1638)));
	assign g1637 = (((!sk[3]) & (!i_15_) & (!i_10_) & (g131) & (!i_9_)) + ((!sk[3]) & (!i_15_) & (!i_10_) & (g131) & (i_9_)) + ((!sk[3]) & (!i_15_) & (i_10_) & (g131) & (!i_9_)) + ((!sk[3]) & (!i_15_) & (i_10_) & (g131) & (i_9_)) + ((!sk[3]) & (i_15_) & (!i_10_) & (g131) & (!i_9_)) + ((!sk[3]) & (i_15_) & (!i_10_) & (g131) & (i_9_)) + ((!sk[3]) & (i_15_) & (i_10_) & (g131) & (!i_9_)) + ((!sk[3]) & (i_15_) & (i_10_) & (g131) & (i_9_)) + ((sk[3]) & (!i_15_) & (!i_10_) & (!g131) & (!i_9_)) + ((sk[3]) & (!i_15_) & (!i_10_) & (g131) & (!i_9_)) + ((sk[3]) & (!i_15_) & (!i_10_) & (g131) & (i_9_)) + ((sk[3]) & (!i_15_) & (i_10_) & (!g131) & (!i_9_)) + ((sk[3]) & (!i_15_) & (i_10_) & (!g131) & (i_9_)) + ((sk[3]) & (!i_15_) & (i_10_) & (g131) & (!i_9_)) + ((sk[3]) & (!i_15_) & (i_10_) & (g131) & (i_9_)) + ((sk[3]) & (i_15_) & (!i_10_) & (!g131) & (!i_9_)) + ((sk[3]) & (i_15_) & (!i_10_) & (!g131) & (i_9_)) + ((sk[3]) & (i_15_) & (!i_10_) & (g131) & (!i_9_)) + ((sk[3]) & (i_15_) & (!i_10_) & (g131) & (i_9_)) + ((sk[3]) & (i_15_) & (i_10_) & (!g131) & (!i_9_)) + ((sk[3]) & (i_15_) & (i_10_) & (!g131) & (i_9_)) + ((sk[3]) & (i_15_) & (i_10_) & (g131) & (!i_9_)) + ((sk[3]) & (i_15_) & (i_10_) & (g131) & (i_9_)));
	assign g1638 = (((!i_15_) & (!i_10_) & (!g122) & (sk[4]) & (!i_9_)) + ((!i_15_) & (!i_10_) & (!g122) & (sk[4]) & (i_9_)) + ((!i_15_) & (!i_10_) & (g122) & (!sk[4]) & (!i_9_)) + ((!i_15_) & (!i_10_) & (g122) & (!sk[4]) & (i_9_)) + ((!i_15_) & (!i_10_) & (g122) & (sk[4]) & (!i_9_)) + ((!i_15_) & (!i_10_) & (g122) & (sk[4]) & (i_9_)) + ((!i_15_) & (i_10_) & (!g122) & (sk[4]) & (!i_9_)) + ((!i_15_) & (i_10_) & (!g122) & (sk[4]) & (i_9_)) + ((!i_15_) & (i_10_) & (g122) & (!sk[4]) & (!i_9_)) + ((!i_15_) & (i_10_) & (g122) & (!sk[4]) & (i_9_)) + ((!i_15_) & (i_10_) & (g122) & (sk[4]) & (!i_9_)) + ((i_15_) & (!i_10_) & (!g122) & (sk[4]) & (!i_9_)) + ((i_15_) & (!i_10_) & (!g122) & (sk[4]) & (i_9_)) + ((i_15_) & (!i_10_) & (g122) & (!sk[4]) & (!i_9_)) + ((i_15_) & (!i_10_) & (g122) & (!sk[4]) & (i_9_)) + ((i_15_) & (!i_10_) & (g122) & (sk[4]) & (!i_9_)) + ((i_15_) & (!i_10_) & (g122) & (sk[4]) & (i_9_)) + ((i_15_) & (i_10_) & (!g122) & (sk[4]) & (!i_9_)) + ((i_15_) & (i_10_) & (!g122) & (sk[4]) & (i_9_)) + ((i_15_) & (i_10_) & (g122) & (!sk[4]) & (!i_9_)) + ((i_15_) & (i_10_) & (g122) & (!sk[4]) & (i_9_)) + ((i_15_) & (i_10_) & (g122) & (sk[4]) & (!i_9_)) + ((i_15_) & (i_10_) & (g122) & (sk[4]) & (i_9_)));
	assign g1639 = (((!g1640) & (sk[5]) & (!g1641)) + ((g1640) & (!sk[5]) & (!g1641)) + ((g1640) & (!sk[5]) & (g1641)));
	assign g1640 = (((!sk[6]) & (g75) & (!g1642)) + ((!sk[6]) & (g75) & (g1642)) + ((sk[6]) & (!g75) & (g1642)));
	assign g1641 = (((g75) & (!sk[7]) & (!g1643)) + ((g75) & (!sk[7]) & (g1643)) + ((g75) & (sk[7]) & (g1643)));
	assign g1642 = (((g87) & (!sk[8]) & (!g1646)) + ((g87) & (!sk[8]) & (g1646)) + ((g87) & (sk[8]) & (g1646)));
	assign g1643 = (((!sk[9]) & (g1644) & (!g1645)) + ((!sk[9]) & (g1644) & (g1645)) + ((sk[9]) & (!g1644) & (!g1645)));
	assign g1644 = (((!sk[10]) & (g87) & (!g1647)) + ((!sk[10]) & (g87) & (g1647)) + ((sk[10]) & (!g87) & (g1647)));
	assign g1645 = (((!sk[11]) & (g87) & (!g1648)) + ((!sk[11]) & (g87) & (g1648)) + ((sk[11]) & (g87) & (g1648)));
	assign g1646 = (((!sk[12]) & (!g79) & (!g89) & (g125)) + ((!sk[12]) & (!g79) & (g89) & (!g125)) + ((!sk[12]) & (!g79) & (g89) & (g125)) + ((!sk[12]) & (g79) & (!g89) & (g125)) + ((!sk[12]) & (g79) & (g89) & (!g125)) + ((!sk[12]) & (g79) & (g89) & (g125)) + ((sk[12]) & (!g79) & (g89) & (!g125)) + ((sk[12]) & (g79) & (g89) & (!g125)) + ((sk[12]) & (g79) & (g89) & (g125)));
	assign g1647 = (((!g131) & (!g79) & (g130) & (!sk[13]) & (!g125)) + ((!g131) & (!g79) & (g130) & (!sk[13]) & (g125)) + ((!g131) & (g79) & (g130) & (!sk[13]) & (!g125)) + ((!g131) & (g79) & (g130) & (!sk[13]) & (g125)) + ((g131) & (!g79) & (g130) & (!sk[13]) & (!g125)) + ((g131) & (!g79) & (g130) & (!sk[13]) & (g125)) + ((g131) & (!g79) & (g130) & (sk[13]) & (!g125)) + ((g131) & (g79) & (g130) & (!sk[13]) & (!g125)) + ((g131) & (g79) & (g130) & (!sk[13]) & (g125)) + ((g131) & (g79) & (g130) & (sk[13]) & (!g125)) + ((g131) & (g79) & (g130) & (sk[13]) & (g125)));
	assign g1648 = (((!g79) & (sk[14]) & (!g125)) + ((g79) & (!sk[14]) & (!g125)) + ((g79) & (!sk[14]) & (g125)) + ((g79) & (sk[14]) & (!g125)) + ((g79) & (sk[14]) & (g125)));

endmodule