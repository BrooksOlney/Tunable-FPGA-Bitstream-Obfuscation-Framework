module seq_qmap_map (sk, i_37_, i_7_, i_5_, i_36_, i_34_, i_35_, i_33_, i_32_, i_31_, i_16_, i_9_, i_40_, i_38_, i_39_, i_11_, i_12_, i_15_, i_24_, i_17_, i_22_, i_2_, i_1_, i_3_, i_4_, i_13_, i_0_, i_10_, i_27_, i_25_, i_26_, i_18_, i_19_, i_30_, i_28_, i_29_, i_21_, i_23_, i_14_, i_20_, i_8_, i_6_, o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_, o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_, o_31_, o_32_, o_33_, o_34_);

	input i_37_;
	input i_7_;
	input i_5_;
	input i_36_;
	input i_34_;
	input i_35_;
	input i_33_;
	input i_32_;
	input i_31_;
	input i_16_;
	input i_9_;
	input i_40_;
	input i_38_;
	input i_39_;
	input i_11_;
	input i_12_;
	input i_15_;
	input i_24_;
	input i_17_;
	input i_22_;
	input i_2_;
	input i_1_;
	input i_3_;
	input i_4_;
	input i_13_;
	input i_0_;
	input i_10_;
	input i_27_;
	input i_25_;
	input i_26_;
	input i_18_;
	input i_19_;
	input i_30_;
	input i_28_;
	input i_29_;
	input i_21_;
	input i_23_;
	input i_14_;
	input i_20_;
	input i_8_;
	input i_6_;
	output o_0_;
	output o_1_;
	output o_2_;
	output o_3_;
	output o_4_;
	output o_5_;
	output o_6_;
	output o_7_;
	output o_8_;
	output o_9_;
	output o_10_;
	output o_11_;
	output o_12_;
	output o_13_;
	output o_14_;
	output o_15_;
	output o_16_;
	output o_17_;
	output o_18_;
	output o_19_;
	output o_20_;
	output o_21_;
	output o_22_;
	output o_23_;
	output o_24_;
	output o_25_;
	output o_26_;
	output o_27_;
	output o_28_;
	output o_29_;
	output o_30_;
	output o_31_;
	output o_32_;
	output o_33_;
	output o_34_;



	wire g159, g207, g230, g287, g328, g421, g439, g440, g441, g453, g458, g459, g184, g469, g519, g526, g554, g565, g597, g613, g616;
	wire g617, g607, g615, g619, g610, g660, g689, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14;
	wire g15, g16, g17, g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29, g30, g31, g32, g33, g34, g35;
	wire g36, g37, g38, g39, g40, g41, g42, g43, g44, g45, g46, g47, g48, g49, g50, g51, g52, g53, g54, g55, g56;
	wire g57, g58, g59, g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g70, g71, g72, g73, g74, g75, g76, g77;
	wire g78, g79, g80, g81, g82, g83, g84, g85, g86, g87, g88, g89, g90, g91, g92, g93, g94, g95, g96, g97, g98;
	wire g99, g100, g101, g102, g103, g104, g105, g106, g107, g108, g109, g110, g692, g111, g112, g113, g114, g115, g116, g117, g118;
	wire g119, g120, g121, g122, g123, g124, g125, g126, g127, g128, g129, g130, g131, g132, g133, g134, g135, g136, g137, g138, g139;
	wire g140, g141, g142, g143, g144, g145, g146, g147, g148, g149, g150, g151, g152, g153, g154, g155, g156, g157, g747, g158, g160;
	wire g161, g162, g163, g164, g165, g166, g167, g168, g169, g170, g171, g172, g173, g174, g175, g176, g177, g178, g691, g179, g180;
	wire g181, g182, g183, g185, g186, g187, g188, g189, g190, g191, g192, g193, g194, g195, g196, g197, g198, g199, g200, g201, g202;
	wire g203, g204, g205, g206, g208, g209, g210, g211, g212, g213, g214, g215, g216, g217, g218, g219, g220, g221, g222, g223, g224;
	wire g225, g226, g227, g228, g229, g231, g232, g233, g234, g235, g236, g237, g238, g239, g240, g241, g242, g243, g244, g245, g246;
	wire g247, g248, g249, g250, g251, g252, g253, g254, g255, g256, g257, g258, g259, g260, g261, g262, g740, g263, g264, g265, g266;
	wire g267, g268, g269, g270, g729, g271, g272, g273, g274, g275, g276, g277, g278, g279, g280, g281, g282, g283, g284, g285, g286;
	wire g288, g289, g290, g291, g292, g293, g294, g295, g296, g297, g298, g299, g300, g301, g302, g303, g304, g305, g306, g307, g308;
	wire g309, g310, g311, g312, g313, g314, g315, g316, g317, g318, g319, g320, g321, g322, g323, g324, g325, g326, g327, g329, g330;
	wire g331, g332, g333, g334, g335, g336, g337, g338, g339, g340, g341, g342, g343, g344, g345, g346, g347, g348, g349, g350, g351;
	wire g352, g353, g354, g355, g356, g357, g723, g358, g359, g360, g361, g362, g363, g364, g365, g366, g367, g368, g369, g370, g371;
	wire g372, g373, g374, g375, g376, g377, g378, g379, g381, g382, g383, g384, g385, g386, g387, g388, g389, g390, g391, g392, g393;
	wire g394, g395, g396, g397, g398, g399, g400, g401, g402, g403, g404, g405, g406, g407, g408, g409, g410, g411, g412, g413, g414;
	wire g415, g416, g417, g418, g419, g420, g422, g423, g424, g425, g426, g427, g428, g429, g430, g431, g432, g433, g434, g435, g436;
	wire g437, g438, g442, g443, g444, g445, g446, g447, g449, g450, g451, g452, g454, g455, g457, g460, g461, g462, g463, g464, g465;
	wire g466, g467, g468, g470, g471, g472, g473, g474, g475, g476, g477, g478, g479, g480, g481, g482, g483, g484, g485, g486, g487;
	wire g488, g489, g491, g492, g493, g494, g495, g496, g497, g498, g499, g500, g501, g502, g503, g504, g505, g506, g507, g508, g509;
	wire g510, g511, g512, g513, g514, g515, g516, g517, g518, g520, g521, g522, g523, g524, g525, g712, g527, g528, g529, g530, g531;
	wire g532, g533, g534, g535, g536, g537, g538, g539, g540, g541, g542, g543, g544, g545, g546, g547, g548, g549, g550, g551, g552;
	wire g553, g555, g556, g557, g558, g559, g560, g561, g562, g563, g564, g566, g567, g568, g569, g570, g571, g572, g573, g574, g576;
	wire g577, g578, g704, g579, g580, g581, g582, g583, g584, g585, g586, g587, g588, g589, g590, g591, g592, g593, g594, g595, g693;
	wire g596, g598, g599, g600, g601, g602, g603, g604, g605, g606, g608, g609, g611, g612, g614, g618, g620, g621, g622, g623, g624;
	wire g626, g627, g629, g630, g631, g632, g633, g634, g635, g636, g637, g638, g639, g640, g641, g642, g643, g644, g645, g646, g647;
	wire g648, g649, g650, g651, g652, g653, g654, g655, g656, g657, g658, g659, g661, g662, g663, g664, g665, g666, g667, g668, g669;
	wire g670, g671, g672, g673, g674, g675, g676, g677, g678, g679, g680, g681, g682, g683, g684, g685, g686, g687, g688, g690, g694;
	wire g695, g696, g699, g697, g698, g702, g703, g700, g701, g705, g706, g707, g709, g708, g711, g710, g713, g714, g715, g717, g716;
	wire g720, g718, g719, g721, g722, g724, g725, g726, g727, g728, g730, g731, g732, g735, g733, g734, g737, g738, g736, g739, g741;
	wire g742, g743, g744, g745, g746, g748, g749, g750, g753, g751, g752, g756, g757, g754, g755, g758, g759;

	lut_sub lut_5 ({g159}, o_0_);
	defparam lut_5.LUT_SIZE = 1;
	defparam lut_5.mask = 2'b10;

	lut_sub lut_9 ({g207}, o_1_);
	defparam lut_9.LUT_SIZE = 1;
	defparam lut_9.mask = 2'b10;

	lut_sub lut_13 ({g230}, o_2_);
	defparam lut_13.LUT_SIZE = 1;
	defparam lut_13.mask = 2'b10;

	lut_sub lut_17 ({g287}, o_3_);
	defparam lut_17.LUT_SIZE = 1;
	defparam lut_17.mask = 2'b10;

	lut_sub lut_21 ({g328}, o_4_);
	defparam lut_21.LUT_SIZE = 1;
	defparam lut_21.mask = 2'b10;

	lut_sub lut_25 ({g421}, o_6_);
	defparam lut_25.LUT_SIZE = 1;
	defparam lut_25.mask = 2'b10;

	lut_sub lut_29 ({g439}, o_7_);
	defparam lut_29.LUT_SIZE = 1;
	defparam lut_29.mask = 2'b10;

	lut_sub lut_33 ({g440}, o_8_);
	defparam lut_33.LUT_SIZE = 1;
	defparam lut_33.mask = 2'b10;

	lut_sub lut_37 ({g441}, o_9_);
	defparam lut_37.LUT_SIZE = 1;
	defparam lut_37.mask = 2'b10;

	lut_sub lut_41 ({g453}, o_11_);
	defparam lut_41.LUT_SIZE = 1;
	defparam lut_41.mask = 2'b10;

	lut_sub lut_45 ({g458}, o_13_);
	defparam lut_45.LUT_SIZE = 1;
	defparam lut_45.mask = 2'b10;

	lut_sub lut_49 ({g459}, o_14_);
	defparam lut_49.LUT_SIZE = 1;
	defparam lut_49.mask = 2'b10;

	lut_sub lut_53 ({g184}, o_15_);
	defparam lut_53.LUT_SIZE = 1;
	defparam lut_53.mask = 2'b10;

	lut_sub lut_57 ({g469}, o_16_);
	defparam lut_57.LUT_SIZE = 1;
	defparam lut_57.mask = 2'b10;

	lut_sub lut_61 ({g519}, o_18_);
	defparam lut_61.LUT_SIZE = 1;
	defparam lut_61.mask = 2'b10;

	lut_sub lut_65 ({g526}, o_19_);
	defparam lut_65.LUT_SIZE = 1;
	defparam lut_65.mask = 2'b10;

	lut_sub lut_69 ({g554}, o_20_);
	defparam lut_69.LUT_SIZE = 1;
	defparam lut_69.mask = 2'b10;

	lut_sub lut_73 ({g565}, o_21_);
	defparam lut_73.LUT_SIZE = 1;
	defparam lut_73.mask = 2'b10;

	lut_sub lut_77 ({g597}, o_23_);
	defparam lut_77.LUT_SIZE = 1;
	defparam lut_77.mask = 2'b10;

	lut_sub lut_81 ({g613}, o_24_);
	defparam lut_81.LUT_SIZE = 1;
	defparam lut_81.mask = 2'b10;

	lut_sub lut_85 ({g616}, o_25_);
	defparam lut_85.LUT_SIZE = 1;
	defparam lut_85.mask = 2'b10;

	lut_sub lut_89 ({g617}, o_26_);
	defparam lut_89.LUT_SIZE = 1;
	defparam lut_89.mask = 2'b10;

	lut_sub lut_93 ({g607}, o_27_);
	defparam lut_93.LUT_SIZE = 1;
	defparam lut_93.mask = 2'b10;

	lut_sub lut_97 ({g615}, o_28_);
	defparam lut_97.LUT_SIZE = 1;
	defparam lut_97.mask = 2'b10;

	lut_sub lut_101 ({g619}, o_29_);
	defparam lut_101.LUT_SIZE = 1;
	defparam lut_101.mask = 2'b10;

	lut_sub lut_105 ({g610}, o_32_);
	defparam lut_105.LUT_SIZE = 1;
	defparam lut_105.mask = 2'b10;

	lut_sub lut_109 ({g660}, o_33_);
	defparam lut_109.LUT_SIZE = 1;
	defparam lut_109.mask = 2'b10;

	lut_sub lut_113 ({g689}, o_34_);
	defparam lut_113.LUT_SIZE = 1;
	defparam lut_113.mask = 2'b10;

	lut_sub lut_117 ({i_7_, i_5_}, g1);
	defparam lut_117.LUT_SIZE = 2;
	defparam lut_117.mask = 4'b0111;

	lut_sub lut_123 ({i_36_, i_34_, i_35_}, g2);
	defparam lut_123.LUT_SIZE = 3;
	defparam lut_123.mask = 8'h80;

	lut_sub lut_127 ({i_33_, i_32_, i_31_}, g3);
	defparam lut_127.LUT_SIZE = 3;
	defparam lut_127.mask = 8'h08;

	lut_sub lut_134 ({g1, g2, g3, i_16_, i_9_}, g4);
	defparam lut_134.LUT_SIZE = 5;
	defparam lut_134.mask = 32'h00080000;

	lut_sub lut_138 ({i_34_, i_35_}, g5);
	defparam lut_138.LUT_SIZE = 2;
	defparam lut_138.mask = 4'b0100;

	lut_sub lut_142 ({i_7_, i_33_, i_32_}, g6);
	defparam lut_142.LUT_SIZE = 3;
	defparam lut_142.mask = 8'h20;

	lut_sub lut_148 ({i_36_, g5, g6}, g7);
	defparam lut_148.LUT_SIZE = 3;
	defparam lut_148.mask = 8'h01;

	lut_sub lut_152 ({i_37_, i_38_, i_39_}, g8);
	defparam lut_152.LUT_SIZE = 3;
	defparam lut_152.mask = 8'h04;

	lut_sub lut_158 ({i_40_, g7, g8}, g9);
	defparam lut_158.LUT_SIZE = 3;
	defparam lut_158.mask = 8'h10;

	lut_sub lut_162 ({i_33_, i_34_, i_35_}, g10);
	defparam lut_162.LUT_SIZE = 3;
	defparam lut_162.mask = 8'hfb;

	lut_sub lut_172 ({i_32_, i_15_}, g11);
	defparam lut_172.LUT_SIZE = 2;
	defparam lut_172.mask = 4'b0100;

	lut_sub lut_178 ({g10, g11, i_24_}, g12);
	defparam lut_178.LUT_SIZE = 3;
	defparam lut_178.mask = 8'h20;

	lut_sub lut_182 ({i_36_, i_37_, i_38_, i_39_, i_40_}, g13);
	defparam lut_182.LUT_SIZE = 5;
	defparam lut_182.mask = 32'hc0400000;

	lut_sub lut_188 ({i_38_, i_39_}, g14);
	defparam lut_188.LUT_SIZE = 2;
	defparam lut_188.mask = 4'b1000;

	lut_sub lut_192 ({i_36_, i_37_, i_38_, i_39_}, g15);
	defparam lut_192.LUT_SIZE = 4;
	defparam lut_192.mask = 16'h9000;

	lut_sub lut_199 ({i_36_, i_40_, g14, g15}, g16);
	defparam lut_199.LUT_SIZE = 4;
	defparam lut_199.mask = 16'ha8aa;

	lut_sub lut_213 ({i_11_, g1, i_12_, g12, g13, g16}, g17);
	defparam lut_213.LUT_SIZE = 6;
	defparam lut_213.mask = 64'h000300000a0b0000;

	lut_sub lut_223 ({i_11_, i_12_, i_15_}, g18);
	defparam lut_223.LUT_SIZE = 3;
	defparam lut_223.mask = 8'h15;

	lut_sub lut_230 ({i_38_, i_40_, g18}, g19);
	defparam lut_230.LUT_SIZE = 3;
	defparam lut_230.mask = 8'h04;

	lut_sub lut_238 ({i_37_, g4, g9, g17, g19}, g20);
	defparam lut_238.LUT_SIZE = 5;
	defparam lut_238.mask = 32'hc080c0c0;

	lut_sub lut_248 ({i_37_, i_38_, i_39_}, g21);
	defparam lut_248.LUT_SIZE = 3;
	defparam lut_248.mask = 8'h08;

	lut_sub lut_252 ({i_11_, i_12_}, g22);
	defparam lut_252.LUT_SIZE = 2;
	defparam lut_252.mask = 4'b1000;

	lut_sub lut_258 ({g1, g22, i_15_}, g23);
	defparam lut_258.LUT_SIZE = 3;
	defparam lut_258.mask = 8'h40;

	lut_sub lut_262 ({i_16_, i_17_}, g24);
	defparam lut_262.LUT_SIZE = 2;
	defparam lut_262.mask = 4'b1000;

	lut_sub lut_269 ({g3, g23, g24}, g25);
	defparam lut_269.LUT_SIZE = 3;
	defparam lut_269.mask = 8'h01;

	lut_sub lut_273 ({i_11_, i_15_}, g26);
	defparam lut_273.LUT_SIZE = 2;
	defparam lut_273.mask = 4'b0001;

	lut_sub lut_277 ({i_36_, i_37_, i_38_}, g27);
	defparam lut_277.LUT_SIZE = 3;
	defparam lut_277.mask = 8'h40;

	lut_sub lut_282 ({i_39_, g27}, g28);
	defparam lut_282.LUT_SIZE = 2;
	defparam lut_282.mask = 4'b0001;

	lut_sub lut_289 ({g1, i_12_, g28, g12}, g29);
	defparam lut_289.LUT_SIZE = 4;
	defparam lut_289.mask = 16'h0100;

	lut_sub lut_293 ({i_38_, i_40_}, g30);
	defparam lut_293.LUT_SIZE = 2;
	defparam lut_293.mask = 4'b1011;

	lut_sub lut_302 ({g1, g2, g3}, g31);
	defparam lut_302.LUT_SIZE = 3;
	defparam lut_302.mask = 8'h10;

	lut_sub lut_306 ({i_38_, i_39_, i_17_}, g32);
	defparam lut_306.LUT_SIZE = 3;
	defparam lut_306.mask = 8'h02;

	lut_sub lut_314 ({g30, g31, i_9_, g4, g32}, g33);
	defparam lut_314.LUT_SIZE = 5;
	defparam lut_314.mask = 32'h33730050;

	lut_sub lut_329 ({g1, i_9_}, g34);
	defparam lut_329.LUT_SIZE = 2;
	defparam lut_329.mask = 4'b1000;

	lut_sub lut_336 ({g2, g21, g18}, g35);
	defparam lut_336.LUT_SIZE = 3;
	defparam lut_336.mask = 8'h01;

	lut_sub lut_343 ({g3, i_16_, i_17_, g34, g35}, g36);
	defparam lut_343.LUT_SIZE = 5;
	defparam lut_343.mask = 32'h00001110;

	lut_sub lut_349 ({i_12_, i_15_}, g37);
	defparam lut_349.LUT_SIZE = 2;
	defparam lut_349.mask = 4'b0001;

	lut_sub lut_357 ({i_37_, i_39_, g30, g26, g4, g37}, g38);
	defparam lut_357.LUT_SIZE = 6;
	defparam lut_357.mask = 64'h1100131311001100;

	lut_sub lut_372 ({i_37_, i_38_, i_39_, i_40_}, g39);
	defparam lut_372.LUT_SIZE = 4;
	defparam lut_372.mask = 16'h0203;

	lut_sub lut_382 ({g31, i_9_, g32, g37, g39}, g40);
	defparam lut_382.LUT_SIZE = 5;
	defparam lut_382.mask = 32'h00005700;

	lut_sub lut_396 ({g26, g29, g33, g36, g38, g40}, g41);
	defparam lut_396.LUT_SIZE = 6;
	defparam lut_396.mask = 64'h8080000080000000;

	lut_sub lut_404 ({i_22_, g10, g11}, g42);
	defparam lut_404.LUT_SIZE = 3;
	defparam lut_404.mask = 8'h40;

	lut_sub lut_410 ({g1, g22}, g43);
	defparam lut_410.LUT_SIZE = 2;
	defparam lut_410.mask = 4'b1000;

	lut_sub lut_416 ({g42, g43}, g44);
	defparam lut_416.LUT_SIZE = 2;
	defparam lut_416.mask = 4'b0001;

	lut_sub lut_420 ({i_36_, i_37_, i_38_}, g45);
	defparam lut_420.LUT_SIZE = 3;
	defparam lut_420.mask = 8'h20;

	lut_sub lut_425 ({i_39_, g45}, g46);
	defparam lut_425.LUT_SIZE = 2;
	defparam lut_425.mask = 4'b0100;

	lut_sub lut_429 ({i_2_, i_1_, i_3_, i_4_}, g47);
	defparam lut_429.LUT_SIZE = 4;
	defparam lut_429.mask = 16'h8000;

	lut_sub lut_433 ({i_7_, i_32_}, g48);
	defparam lut_433.LUT_SIZE = 2;
	defparam lut_433.mask = 4'b1000;

	lut_sub lut_437 ({i_33_, i_34_, i_35_}, g49);
	defparam lut_437.LUT_SIZE = 3;
	defparam lut_437.mask = 8'hfd;

	lut_sub lut_452 ({g28, g46, g47, g48, g49}, g50);
	defparam lut_452.LUT_SIZE = 5;
	defparam lut_452.mask = 32'h00202020;

	lut_sub lut_458 ({i_36_, i_35_}, g51);
	defparam lut_458.LUT_SIZE = 2;
	defparam lut_458.mask = 4'b1000;

	lut_sub lut_463 ({i_37_, i_38_, i_39_, i_40_, g51}, g52);
	defparam lut_463.LUT_SIZE = 5;
	defparam lut_463.mask = 32'h15055100;

	lut_sub lut_474 ({i_33_, i_34_, i_32_, i_31_}, g53);
	defparam lut_474.LUT_SIZE = 4;
	defparam lut_474.mask = 16'h0080;

	lut_sub lut_478 ({i_7_, i_11_, i_5_, i_12_}, g54);
	defparam lut_478.LUT_SIZE = 4;
	defparam lut_478.mask = 16'h8000;

	lut_sub lut_484 ({g53, g54, i_13_}, g55);
	defparam lut_484.LUT_SIZE = 3;
	defparam lut_484.mask = 8'h01;

	lut_sub lut_488 ({i_33_, i_34_, i_35_}, g56);
	defparam lut_488.LUT_SIZE = 3;
	defparam lut_488.mask = 8'h08;

	lut_sub lut_492 ({i_7_, i_5_, i_13_, i_15_}, g57);
	defparam lut_492.LUT_SIZE = 4;
	defparam lut_492.mask = 16'h2000;

	lut_sub lut_498 ({g56, i_32_, i_31_, g57}, g58);
	defparam lut_498.LUT_SIZE = 4;
	defparam lut_498.mask = 16'h0040;

	lut_sub lut_502 ({i_36_, i_37_, i_38_, i_39_, i_40_}, g59);
	defparam lut_502.LUT_SIZE = 5;
	defparam lut_502.mask = 32'h73d00000;

	lut_sub lut_517 ({g52, g55, g58, g59}, g60);
	defparam lut_517.LUT_SIZE = 4;
	defparam lut_517.mask = 16'h111f;

	lut_sub lut_527 ({i_37_, i_38_, i_39_, i_40_}, g61);
	defparam lut_527.LUT_SIZE = 4;
	defparam lut_527.mask = 16'h0200;

	lut_sub lut_534 ({i_11_, g1, i_12_, i_15_, g31, g61}, g62);
	defparam lut_534.LUT_SIZE = 6;
	defparam lut_534.mask = 64'h1111111111101100;

	lut_sub lut_555 ({g28, g44, g50, g60, g62}, g63);
	defparam lut_555.LUT_SIZE = 5;
	defparam lut_555.mask = 32'h80808000;

	lut_sub lut_566 ({g2, g21, g25, g41, g63}, g64);
	defparam lut_566.LUT_SIZE = 5;
	defparam lut_566.mask = 32'h11111110;

	lut_sub lut_576 ({i_33_, i_34_, i_32_}, g65);
	defparam lut_576.LUT_SIZE = 3;
	defparam lut_576.mask = 8'h08;

	lut_sub lut_581 ({i_36_, i_37_, i_35_, g65}, g66);
	defparam lut_581.LUT_SIZE = 4;
	defparam lut_581.mask = 16'h0001;

	lut_sub lut_585 ({i_3_, i_4_}, g67);
	defparam lut_585.LUT_SIZE = 2;
	defparam lut_585.mask = 4'b0100;

	lut_sub lut_590 ({i_7_, i_2_, i_1_, i_0_, g67}, g68);
	defparam lut_590.LUT_SIZE = 5;
	defparam lut_590.mask = 32'h32330000;

	lut_sub lut_600 ({i_38_, i_40_}, g69);
	defparam lut_600.LUT_SIZE = 2;
	defparam lut_600.mask = 4'b1000;

	lut_sub lut_605 ({i_7_, g65}, g70);
	defparam lut_605.LUT_SIZE = 2;
	defparam lut_605.mask = 4'b0100;

	lut_sub lut_609 ({i_36_, i_37_, i_35_}, g71);
	defparam lut_609.LUT_SIZE = 3;
	defparam lut_609.mask = 8'h08;

	lut_sub lut_615 ({g70, i_10_, i_27_, g71}, g72);
	defparam lut_615.LUT_SIZE = 4;
	defparam lut_615.mask = 16'h0001;

	lut_sub lut_619 ({i_39_, i_40_}, g73);
	defparam lut_619.LUT_SIZE = 2;
	defparam lut_619.mask = 4'b1000;

	lut_sub lut_625 ({i_38_, g72, g73}, g74);
	defparam lut_625.LUT_SIZE = 3;
	defparam lut_625.mask = 8'h01;

	lut_sub lut_629 ({i_1_, i_3_, i_4_}, g75);
	defparam lut_629.LUT_SIZE = 3;
	defparam lut_629.mask = 8'h80;

	lut_sub lut_633 ({i_39_, i_40_}, g76);
	defparam lut_633.LUT_SIZE = 2;
	defparam lut_633.mask = 4'b0100;

	lut_sub lut_638 ({i_38_, g76}, g77);
	defparam lut_638.LUT_SIZE = 2;
	defparam lut_638.mask = 4'b0001;

	lut_sub lut_642 ({i_36_, i_35_}, g78);
	defparam lut_642.LUT_SIZE = 2;
	defparam lut_642.mask = 4'b0010;

	lut_sub lut_646 ({i_38_, i_39_, i_40_}, g79);
	defparam lut_646.LUT_SIZE = 3;
	defparam lut_646.mask = 8'h01;

	lut_sub lut_653 ({i_37_, g77, g78, g79}, g80);
	defparam lut_653.LUT_SIZE = 4;
	defparam lut_653.mask = 16'h1103;

	lut_sub lut_663 ({i_2_, g75, g70, i_0_, g80}, g81);
	defparam lut_663.LUT_SIZE = 5;
	defparam lut_663.mask = 32'h01000101;

	lut_sub lut_674 ({g66, g68, g69, g74, g81}, g82);
	defparam lut_674.LUT_SIZE = 5;
	defparam lut_674.mask = 32'h88888880;

	lut_sub lut_684 ({i_36_, i_37_, i_35_}, g83);
	defparam lut_684.LUT_SIZE = 3;
	defparam lut_684.mask = 8'h10;

	lut_sub lut_691 ({i_38_, g65, g76, g83}, g84);
	defparam lut_691.LUT_SIZE = 4;
	defparam lut_691.mask = 16'h0100;

	lut_sub lut_697 ({i_22_, g23, i_24_, g84}, g85);
	defparam lut_697.LUT_SIZE = 4;
	defparam lut_697.mask = 16'h0100;

	lut_sub lut_703 ({i_36_, i_37_, i_38_, g10, g49}, g86);
	defparam lut_703.LUT_SIZE = 5;
	defparam lut_703.mask = 32'ha000000c;

	lut_sub lut_710 ({i_2_, i_1_, i_3_, i_0_}, g87);
	defparam lut_710.LUT_SIZE = 4;
	defparam lut_710.mask = 16'h0040;

	lut_sub lut_714 ({i_36_, i_37_, i_35_}, g88);
	defparam lut_714.LUT_SIZE = 3;
	defparam lut_714.mask = 8'h04;

	lut_sub lut_721 ({g14, g70, g88, i_25_, i_26_}, g89);
	defparam lut_721.LUT_SIZE = 5;
	defparam lut_721.mask = 32'h00000008;

	lut_sub lut_729 ({g48, g86, g87, g89}, g90);
	defparam lut_729.LUT_SIZE = 4;
	defparam lut_729.mask = 16'haaa8;

	lut_sub lut_742 ({g23, g34, g18, i_18_, i_19_}, g91);
	defparam lut_742.LUT_SIZE = 5;
	defparam lut_742.mask = 32'h000a888a;

	lut_sub lut_752 ({i_1_, i_4_, i_0_}, g92);
	defparam lut_752.LUT_SIZE = 3;
	defparam lut_752.mask = 8'h40;

	lut_sub lut_758 ({g92, g7}, g93);
	defparam lut_758.LUT_SIZE = 2;
	defparam lut_758.mask = 4'b0001;

	lut_sub lut_762 ({i_36_, i_34_, i_35_}, g94);
	defparam lut_762.LUT_SIZE = 3;
	defparam lut_762.mask = 8'hdf;

	lut_sub lut_774 ({g6, g94}, g95);
	defparam lut_774.LUT_SIZE = 2;
	defparam lut_774.mask = 4'b0010;

	lut_sub lut_780 ({g92, g95}, g96);
	defparam lut_780.LUT_SIZE = 2;
	defparam lut_780.mask = 4'b0001;

	lut_sub lut_786 ({i_37_, i_38_, g93, g96}, g97);
	defparam lut_786.LUT_SIZE = 4;
	defparam lut_786.mask = 16'h5003;

	lut_sub lut_793 ({i_37_, i_38_, i_39_}, g98);
	defparam lut_793.LUT_SIZE = 3;
	defparam lut_793.mask = 8'h40;

	lut_sub lut_800 ({i_40_, g95, g77, g98}, g99);
	defparam lut_800.LUT_SIZE = 4;
	defparam lut_800.mask = 16'h0307;

	lut_sub lut_808 ({i_37_, i_38_}, g100);
	defparam lut_808.LUT_SIZE = 2;
	defparam lut_808.mask = 4'b1000;

	lut_sub lut_812 ({i_39_, i_40_}, g101);
	defparam lut_812.LUT_SIZE = 2;
	defparam lut_812.mask = 4'b0001;

	lut_sub lut_817 ({g56, i_32_}, g102);
	defparam lut_817.LUT_SIZE = 2;
	defparam lut_817.mask = 4'b0010;

	lut_sub lut_824 ({i_36_, g100, g101, g102}, g103);
	defparam lut_824.LUT_SIZE = 4;
	defparam lut_824.mask = 16'h0001;

	lut_sub lut_828 ({i_38_, i_39_}, g104);
	defparam lut_828.LUT_SIZE = 2;
	defparam lut_828.mask = 4'b0010;

	lut_sub lut_833 ({i_36_, i_40_, g104}, g105);
	defparam lut_833.LUT_SIZE = 3;
	defparam lut_833.mask = 8'h10;

	lut_sub lut_837 ({i_33_, i_35_, i_32_}, g106);
	defparam lut_837.LUT_SIZE = 3;
	defparam lut_837.mask = 8'h08;

	lut_sub lut_842 ({g1, i_30_, i_28_, i_29_}, g107);
	defparam lut_842.LUT_SIZE = 4;
	defparam lut_842.mask = 16'h0400;

	lut_sub lut_847 ({g1, i_30_, i_28_, i_29_}, g108);
	defparam lut_847.LUT_SIZE = 4;
	defparam lut_847.mask = 16'h2000;

	lut_sub lut_855 ({i_31_, g105, g106, g107, g108}, g109);
	defparam lut_855.LUT_SIZE = 5;
	defparam lut_855.mask = 32'h00070000;

	lut_sub lut_864 ({i_7_, i_11_, g99, g103, g109}, g110);
	defparam lut_864.LUT_SIZE = 5;
	defparam lut_864.mask = 32'ha080a0a0;

	lut_sub lut_879 ({g85, g90, g692, g97, g110}, g111);
	defparam lut_879.LUT_SIZE = 5;
	defparam lut_879.mask = 32'h00400000;

	lut_sub lut_883 ({i_37_, i_38_, i_39_}, g112);
	defparam lut_883.LUT_SIZE = 3;
	defparam lut_883.mask = 8'h10;

	lut_sub lut_888 ({i_40_, g112}, g113);
	defparam lut_888.LUT_SIZE = 2;
	defparam lut_888.mask = 4'b0001;

	lut_sub lut_896 ({g24, g31, g37, g113}, g114);
	defparam lut_896.LUT_SIZE = 4;
	defparam lut_896.mask = 16'h0001;

	lut_sub lut_900 ({i_39_, i_40_}, g115);
	defparam lut_900.LUT_SIZE = 2;
	defparam lut_900.mask = 4'b0010;

	lut_sub lut_904 ({i_37_, i_38_}, g116);
	defparam lut_904.LUT_SIZE = 2;
	defparam lut_904.mask = 4'b0001;

	lut_sub lut_911 ({i_36_, g10, g48, g116, i_0_}, g117);
	defparam lut_911.LUT_SIZE = 5;
	defparam lut_911.mask = 32'h01000000;

	lut_sub lut_916 ({i_38_, g115}, g118);
	defparam lut_916.LUT_SIZE = 2;
	defparam lut_916.mask = 4'b0100;

	lut_sub lut_922 ({i_37_, g51, g118}, g119);
	defparam lut_922.LUT_SIZE = 3;
	defparam lut_922.mask = 8'h01;

	lut_sub lut_932 ({g53, g115, g117, g107, g108, g119}, g120);
	defparam lut_932.LUT_SIZE = 6;
	defparam lut_932.mask = 64'h000000ff151515ff;

	lut_sub lut_960 ({i_36_, i_34_, i_35_}, g121);
	defparam lut_960.LUT_SIZE = 3;
	defparam lut_960.mask = 8'h40;

	lut_sub lut_964 ({i_33_, i_32_}, g122);
	defparam lut_964.LUT_SIZE = 2;
	defparam lut_964.mask = 4'b1101;

	lut_sub lut_972 ({g122, i_22_, g23, i_24_, i_21_}, g123);
	defparam lut_972.LUT_SIZE = 5;
	defparam lut_972.mask = 32'h00010000;

	lut_sub lut_977 ({i_40_, g21}, g124);
	defparam lut_977.LUT_SIZE = 2;
	defparam lut_977.mask = 4'b0001;

	lut_sub lut_983 ({g122, g121}, g125);
	defparam lut_983.LUT_SIZE = 2;
	defparam lut_983.mask = 4'b0100;

	lut_sub lut_988 ({i_37_, i_38_, i_39_, i_40_, g125}, g126);
	defparam lut_988.LUT_SIZE = 5;
	defparam lut_988.mask = 32'h40040000;

	lut_sub lut_998 ({g23, g121, g123, g124, g126}, g127);
	defparam lut_998.LUT_SIZE = 5;
	defparam lut_998.mask = 32'h00035557;

	lut_sub lut_1014 ({i_32_, g54, i_13_, g10}, g128);
	defparam lut_1014.LUT_SIZE = 4;
	defparam lut_1014.mask = 16'h0200;

	lut_sub lut_1019 ({i_36_, i_40_, g14}, g129);
	defparam lut_1019.LUT_SIZE = 3;
	defparam lut_1019.mask = 8'h10;

	lut_sub lut_1025 ({g122, g94}, g130);
	defparam lut_1025.LUT_SIZE = 2;
	defparam lut_1025.mask = 4'b1000;

	lut_sub lut_1029 ({i_38_, i_39_, i_40_}, g131);
	defparam lut_1029.LUT_SIZE = 3;
	defparam lut_1029.mask = 8'h10;

	lut_sub lut_1035 ({g130, g131}, g132);
	defparam lut_1035.LUT_SIZE = 2;
	defparam lut_1035.mask = 4'b0001;

	lut_sub lut_1043 ({g23, g128, g129, g132}, g133);
	defparam lut_1043.LUT_SIZE = 4;
	defparam lut_1043.mask = 16'h0357;

	lut_sub lut_1055 ({i_34_, g51, g122}, g134);
	defparam lut_1055.LUT_SIZE = 3;
	defparam lut_1055.mask = 8'h02;

	lut_sub lut_1061 ({i_38_, g101, g134}, g135);
	defparam lut_1061.LUT_SIZE = 3;
	defparam lut_1061.mask = 8'h10;

	lut_sub lut_1065 ({i_36_, i_37_, i_35_}, g136);
	defparam lut_1065.LUT_SIZE = 3;
	defparam lut_1065.mask = 8'h80;

	lut_sub lut_1071 ({i_38_, i_40_, g55, g136}, g137);
	defparam lut_1071.LUT_SIZE = 4;
	defparam lut_1071.mask = 16'h0010;

	lut_sub lut_1076 ({g56, i_32_, i_31_}, g138);
	defparam lut_1076.LUT_SIZE = 3;
	defparam lut_1076.mask = 8'h08;

	lut_sub lut_1081 ({i_38_, g76}, g139);
	defparam lut_1081.LUT_SIZE = 2;
	defparam lut_1081.mask = 4'b0100;

	lut_sub lut_1090 ({i_40_, g27, g138, g57, g139, g125}, g140);
	defparam lut_1090.LUT_SIZE = 6;
	defparam lut_1090.mask = 64'h0101010f01010101;

	lut_sub lut_1108 ({g1, i_13_, g135, g137, g140}, g141);
	defparam lut_1108.LUT_SIZE = 5;
	defparam lut_1108.mask = 32'h88808888;

	lut_sub lut_1123 ({g114, g120, g127, g133, g141}, g142);
	defparam lut_1123.LUT_SIZE = 5;
	defparam lut_1123.mask = 32'h40000000;

	lut_sub lut_1129 ({g10, g11}, g143);
	defparam lut_1129.LUT_SIZE = 2;
	defparam lut_1129.mask = 4'b0100;

	lut_sub lut_1135 ({g143, g43}, g144);
	defparam lut_1135.LUT_SIZE = 2;
	defparam lut_1135.mask = 4'b0001;

	lut_sub lut_1141 ({i_11_, g1, i_12_, g24}, g145);
	defparam lut_1141.LUT_SIZE = 4;
	defparam lut_1141.mask = 16'h0040;

	lut_sub lut_1148 ({g56, i_31_, g11, g145}, g146);
	defparam lut_1148.LUT_SIZE = 4;
	defparam lut_1148.mask = 16'h0010;

	lut_sub lut_1154 ({i_37_, i_38_, i_39_, g57, g125}, g147);
	defparam lut_1154.LUT_SIZE = 5;
	defparam lut_1154.mask = 32'h10010000;

	lut_sub lut_1161 ({i_34_, g6, g78}, g148);
	defparam lut_1161.LUT_SIZE = 3;
	defparam lut_1161.mask = 8'h10;

	lut_sub lut_1166 ({i_37_, i_38_, i_39_, i_40_, g148}, g149);
	defparam lut_1166.LUT_SIZE = 5;
	defparam lut_1166.mask = 32'h00000004;

	lut_sub lut_1174 ({g128, g147, g15, g149}, g150);
	defparam lut_1174.LUT_SIZE = 4;
	defparam lut_1174.mask = 16'ha080;

	lut_sub lut_1180 ({i_36_, i_37_, i_35_}, g151);
	defparam lut_1180.LUT_SIZE = 3;
	defparam lut_1180.mask = 8'h40;

	lut_sub lut_1186 ({i_38_, i_39_, g65, g151}, g152);
	defparam lut_1186.LUT_SIZE = 4;
	defparam lut_1186.mask = 16'hfffe;

	lut_sub lut_1204 ({i_22_, i_24_, i_21_}, g153);
	defparam lut_1204.LUT_SIZE = 3;
	defparam lut_1204.mask = 8'h02;

	lut_sub lut_1210 ({g18, i_23_, g153}, g154);
	defparam lut_1210.LUT_SIZE = 3;
	defparam lut_1210.mask = 8'h04;

	lut_sub lut_1215 ({g1, i_9_}, g155);
	defparam lut_1215.LUT_SIZE = 2;
	defparam lut_1215.mask = 4'b0100;

	lut_sub lut_1222 ({g125, i_18_, g124, g155, i_19_}, g156);
	defparam lut_1222.LUT_SIZE = 5;
	defparam lut_1222.mask = 32'h00000103;

	lut_sub lut_1231 ({i_32_, g10, g45, g76}, g157);
	defparam lut_1231.LUT_SIZE = 4;
	defparam lut_1231.mask = 16'h1000;

	lut_sub lut_1240 ({g28, i_21_, g144, g146, g150, g747}, g158);
	defparam lut_1240.LUT_SIZE = 6;
	defparam lut_1240.mask = 64'h1111111110101000;

	lut_sub lut_1260 ({g20, g64, g82, g111, g142, g158}, g159);
	defparam lut_1260.LUT_SIZE = 6;
	defparam lut_1260.mask = 64'h0000000000000001;

	lut_sub lut_1265 ({i_36_, g5}, g160);
	defparam lut_1265.LUT_SIZE = 2;
	defparam lut_1265.mask = 4'b0001;

	lut_sub lut_1272 ({g100, g122, i_25_, i_26_, g160}, g161);
	defparam lut_1272.LUT_SIZE = 5;
	defparam lut_1272.mask = 32'h00001500;

	lut_sub lut_1278 ({i_33_, i_34_}, g162);
	defparam lut_1278.LUT_SIZE = 2;
	defparam lut_1278.mask = 4'b1101;

	lut_sub lut_1284 ({i_11_, i_36_, i_12_}, g163);
	defparam lut_1284.LUT_SIZE = 3;
	defparam lut_1284.mask = 8'h10;

	lut_sub lut_1291 ({i_40_, g162, i_32_, g98, g163}, g164);
	defparam lut_1291.LUT_SIZE = 5;
	defparam lut_1291.mask = 32'h00001000;

	lut_sub lut_1297 ({g101, g27}, g165);
	defparam lut_1297.LUT_SIZE = 2;
	defparam lut_1297.mask = 4'b0001;

	lut_sub lut_1302 ({i_5_, i_16_, i_17_, i_9_, g18}, g166);
	defparam lut_1302.LUT_SIZE = 5;
	defparam lut_1302.mask = 32'h01150000;

	lut_sub lut_1312 ({g102, g165, g166}, g167);
	defparam lut_1312.LUT_SIZE = 3;
	defparam lut_1312.mask = 8'h01;

	lut_sub lut_1318 ({i_37_, g51, g14}, g168);
	defparam lut_1318.LUT_SIZE = 3;
	defparam lut_1318.mask = 8'h01;

	lut_sub lut_1322 ({i_5_, i_15_, i_16_, i_17_, i_9_}, g169);
	defparam lut_1322.LUT_SIZE = 5;
	defparam lut_1322.mask = 32'h00170000;

	lut_sub lut_1330 ({i_12_, i_14_, g169}, g170);
	defparam lut_1330.LUT_SIZE = 3;
	defparam lut_1330.mask = 8'h04;

	lut_sub lut_1334 ({i_16_, i_17_}, g171);
	defparam lut_1334.LUT_SIZE = 2;
	defparam lut_1334.mask = 4'b0001;

	lut_sub lut_1338 ({i_5_, i_13_, i_15_}, g172);
	defparam lut_1338.LUT_SIZE = 3;
	defparam lut_1338.mask = 8'h80;

	lut_sub lut_1342 ({i_36_, i_37_, i_38_, i_39_, i_40_, i_35_}, g173);
	defparam lut_1342.LUT_SIZE = 6;
	defparam lut_1342.mask = 64'h7a02a00000000000;

	lut_sub lut_1355 ({g51, i_31_, i_5_, g37}, g174);
	defparam lut_1355.LUT_SIZE = 4;
	defparam lut_1355.mask = 16'h0008;

	lut_sub lut_1361 ({i_38_, i_39_, g83, g174}, g175);
	defparam lut_1361.LUT_SIZE = 4;
	defparam lut_1361.mask = 16'ha8aa;

	lut_sub lut_1371 ({i_36_, i_37_, i_38_, i_39_, i_40_, i_35_}, g176);
	defparam lut_1371.LUT_SIZE = 6;
	defparam lut_1371.mask = 64'h0010014105140002;

	lut_sub lut_1387 ({g172, g173, g175, g176}, g177);
	defparam lut_1387.LUT_SIZE = 4;
	defparam lut_1387.mask = 16'h2220;

	lut_sub lut_1397 ({i_34_, g51, g122, g47, g113}, g178);
	defparam lut_1397.LUT_SIZE = 5;
	defparam lut_1397.mask = 32'hf0f00010;

	lut_sub lut_1414 ({i_34_, g168, g170, g691, g177, g178}, g179);
	defparam lut_1414.LUT_SIZE = 6;
	defparam lut_1414.mask = 64'h4444455555555555;

	lut_sub lut_1447 ({g27, g106, g73}, g180);
	defparam lut_1447.LUT_SIZE = 3;
	defparam lut_1447.mask = 8'h01;

	lut_sub lut_1455 ({g101, g45, g152, g106}, g181);
	defparam lut_1455.LUT_SIZE = 4;
	defparam lut_1455.mask = 16'h3332;

	lut_sub lut_1468 ({g30, g65, g83}, g182);
	defparam lut_1468.LUT_SIZE = 3;
	defparam lut_1468.mask = 8'h10;

	lut_sub lut_1473 ({i_36_, i_32_, i_31_, i_5_, g21}, g183);
	defparam lut_1473.LUT_SIZE = 5;
	defparam lut_1473.mask = 32'h08000000;

	lut_sub lut_1477 ({i_7_, i_33_}, g184);
	defparam lut_1477.LUT_SIZE = 2;
	defparam lut_1477.mask = 4'b1110;

	lut_sub lut_1485 ({g122, i_5_, g22, i_13_}, g185);
	defparam lut_1485.LUT_SIZE = 4;
	defparam lut_1485.mask = 16'h2000;

	lut_sub lut_1492 ({i_37_, g51, g131, g185}, g186);
	defparam lut_1492.LUT_SIZE = 4;
	defparam lut_1492.mask = 16'h0001;

	lut_sub lut_1496 ({i_38_, i_39_, i_40_}, g187);
	defparam lut_1496.LUT_SIZE = 3;
	defparam lut_1496.mask = 8'h80;

	lut_sub lut_1503 ({i_34_, g122, g71, g187}, g188);
	defparam lut_1503.LUT_SIZE = 4;
	defparam lut_1503.mask = 16'h0010;

	lut_sub lut_1509 ({i_38_, g136, g73}, g189);
	defparam lut_1509.LUT_SIZE = 3;
	defparam lut_1509.mask = 8'h01;

	lut_sub lut_1513 ({i_37_, i_38_, i_39_, i_40_}, g190);
	defparam lut_1513.LUT_SIZE = 4;
	defparam lut_1513.mask = 16'h71c0;

	lut_sub lut_1527 ({g2, g188, g185, g189, g190}, g191);
	defparam lut_1527.LUT_SIZE = 5;
	defparam lut_1527.mask = 32'hfc00f800;

	lut_sub lut_1546 ({g56, g183, g184, g186, g191}, g192);
	defparam lut_1546.LUT_SIZE = 5;
	defparam lut_1546.mask = 32'h04040400;

	lut_sub lut_1557 ({g180, g172, g181, g182, g192}, g193);
	defparam lut_1557.LUT_SIZE = 5;
	defparam lut_1557.mask = 32'h55045500;

	lut_sub lut_1571 ({i_31_, g122, g2}, g194);
	defparam lut_1571.LUT_SIZE = 3;
	defparam lut_1571.mask = 8'h04;

	lut_sub lut_1575 ({i_16_, i_17_, i_9_}, g195);
	defparam lut_1575.LUT_SIZE = 3;
	defparam lut_1575.mask = 8'he8;

	lut_sub lut_1584 ({g194, g195}, g196);
	defparam lut_1584.LUT_SIZE = 2;
	defparam lut_1584.mask = 4'b0001;

	lut_sub lut_1589 ({i_34_, g122}, g197);
	defparam lut_1589.LUT_SIZE = 2;
	defparam lut_1589.mask = 4'b0010;

	lut_sub lut_1594 ({i_5_, g18}, g198);
	defparam lut_1594.LUT_SIZE = 2;
	defparam lut_1594.mask = 4'b0100;

	lut_sub lut_1599 ({i_37_, g76}, g199);
	defparam lut_1599.LUT_SIZE = 2;
	defparam lut_1599.mask = 4'b0100;

	lut_sub lut_1608 ({i_24_, g125, g197, g189, g198, g199}, g200);
	defparam lut_1608.LUT_SIZE = 6;
	defparam lut_1608.mask = 64'h000f000f000f111f;

	lut_sub lut_1630 ({i_11_, i_12_, i_14_}, g201);
	defparam lut_1630.LUT_SIZE = 3;
	defparam lut_1630.mask = 8'h01;

	lut_sub lut_1635 ({i_15_, i_16_, i_17_, i_9_, g201}, g202);
	defparam lut_1635.LUT_SIZE = 5;
	defparam lut_1635.mask = 32'h00000115;

	lut_sub lut_1646 ({g65, g136, g79, g202}, g203);
	defparam lut_1646.LUT_SIZE = 4;
	defparam lut_1646.mask = 16'h0001;

	lut_sub lut_1652 ({i_5_, g22, i_13_, g125}, g204);
	defparam lut_1652.LUT_SIZE = 4;
	defparam lut_1652.mask = 16'h0400;

	lut_sub lut_1657 ({i_37_, i_38_, i_39_, i_40_, g204}, g205);
	defparam lut_1657.LUT_SIZE = 5;
	defparam lut_1657.mask = 32'h50051100;

	lut_sub lut_1670 ({i_5_, g196, g200, g203, g205}, g206);
	defparam lut_1670.LUT_SIZE = 5;
	defparam lut_1670.mask = 32'h80008080;

	lut_sub lut_1682 ({g161, g164, g167, g179, g193, g206}, g207);
	defparam lut_1682.LUT_SIZE = 6;
	defparam lut_1682.mask = 64'h1000000000000000;

	lut_sub lut_1692 ({g2, g21, g3, g113, g184, g691}, g208);
	defparam lut_1692.LUT_SIZE = 6;
	defparam lut_1692.mask = 64'h3333333333323322;

	lut_sub lut_1725 ({i_5_, g3, i_30_, i_28_, i_29_}, g209);
	defparam lut_1725.LUT_SIZE = 5;
	defparam lut_1725.mask = 32'h00db0000;

	lut_sub lut_1738 ({g2, g77, g119, g209}, g210);
	defparam lut_1738.LUT_SIZE = 4;
	defparam lut_1738.mask = 16'h1115;

	lut_sub lut_1749 ({g14, g65, g83}, g211);
	defparam lut_1749.LUT_SIZE = 3;
	defparam lut_1749.mask = 8'h01;

	lut_sub lut_1754 ({i_5_, i_9_, g18, i_18_, i_19_}, g212);
	defparam lut_1754.LUT_SIZE = 5;
	defparam lut_1754.mask = 32'h01070000;

	lut_sub lut_1763 ({i_23_, g153, g212}, g213);
	defparam lut_1763.LUT_SIZE = 3;
	defparam lut_1763.mask = 8'h01;

	lut_sub lut_1769 ({i_34_, g122, g78}, g214);
	defparam lut_1769.LUT_SIZE = 3;
	defparam lut_1769.mask = 8'h40;

	lut_sub lut_1774 ({i_37_, g104}, g215);
	defparam lut_1774.LUT_SIZE = 2;
	defparam lut_1774.mask = 4'b0100;

	lut_sub lut_1778 ({i_36_, i_37_, i_38_}, g216);
	defparam lut_1778.LUT_SIZE = 3;
	defparam lut_1778.mask = 8'h04;

	lut_sub lut_1785 ({g65, g76, g216}, g217);
	defparam lut_1785.LUT_SIZE = 3;
	defparam lut_1785.mask = 8'h01;

	lut_sub lut_1792 ({i_10_, i_27_, g214, g215, g217}, g218);
	defparam lut_1792.LUT_SIZE = 5;
	defparam lut_1792.mask = 32'ha8a8a8aa;

	lut_sub lut_1810 ({i_37_, g51, g197}, g219);
	defparam lut_1810.LUT_SIZE = 3;
	defparam lut_1810.mask = 8'h01;

	lut_sub lut_1816 ({g112, g124}, g220);
	defparam lut_1816.LUT_SIZE = 2;
	defparam lut_1816.mask = 4'b1000;

	lut_sub lut_1825 ({g47, g130, g118, g219, g220}, g221);
	defparam lut_1825.LUT_SIZE = 5;
	defparam lut_1825.mask = 32'h030303ab;

	lut_sub lut_1840 ({i_5_, i_9_, g18, i_18_}, g222);
	defparam lut_1840.LUT_SIZE = 4;
	defparam lut_1840.mask = 16'h1300;

	lut_sub lut_1852 ({g125, g153, g79, g204, g199, g222}, g223);
	defparam lut_1852.LUT_SIZE = 6;
	defparam lut_1852.mask = 64'h0303030303030357;

	lut_sub lut_1879 ({g211, g213, g218, g221, g223}, g224);
	defparam lut_1879.LUT_SIZE = 5;
	defparam lut_1879.mask = 32'h08080800;

	lut_sub lut_1886 ({i_37_, g14}, g225);
	defparam lut_1886.LUT_SIZE = 2;
	defparam lut_1886.mask = 4'b0100;

	lut_sub lut_1893 ({g122, g160, g225}, g226);
	defparam lut_1893.LUT_SIZE = 3;
	defparam lut_1893.mask = 8'h10;

	lut_sub lut_1897 ({i_36_, i_37_, i_38_, i_39_, i_40_, i_35_}, g227);
	defparam lut_1897.LUT_SIZE = 6;
	defparam lut_1897.mask = 64'h0010400100142a00;

	lut_sub lut_1912 ({g76, g151, g172, g227}, g228);
	defparam lut_1912.LUT_SIZE = 4;
	defparam lut_1912.mask = 16'haaa8;

	lut_sub lut_1925 ({g65, i_25_, i_26_, g226, g228}, g229);
	defparam lut_1925.LUT_SIZE = 5;
	defparam lut_1925.mask = 32'hfccc5444;

	lut_sub lut_1948 ({g200, g208, g210, g224, g229}, g230);
	defparam lut_1948.LUT_SIZE = 5;
	defparam lut_1948.mask = 32'h00100000;

	lut_sub lut_1955 ({i_22_, g112, g125, g198}, g231);
	defparam lut_1955.LUT_SIZE = 4;
	defparam lut_1955.mask = 16'h0100;

	lut_sub lut_1959 ({i_5_, i_9_}, g232);
	defparam lut_1959.LUT_SIZE = 2;
	defparam lut_1959.mask = 4'b1000;

	lut_sub lut_1964 ({i_11_, i_38_, i_39_, g232}, g233);
	defparam lut_1964.LUT_SIZE = 4;
	defparam lut_1964.mask = 16'h0010;

	lut_sub lut_1968 ({i_36_, i_37_, i_38_, i_39_}, g234);
	defparam lut_1968.LUT_SIZE = 4;
	defparam lut_1968.mask = 16'h001f;

	lut_sub lut_1978 ({i_40_, i_32_, g47, i_0_, g234}, g235);
	defparam lut_1978.LUT_SIZE = 5;
	defparam lut_1978.mask = 32'h00001000;

	lut_sub lut_1985 ({i_36_, g11, i_16_, g233, g235}, g236);
	defparam lut_1985.LUT_SIZE = 5;
	defparam lut_1985.mask = 32'haa8aaaaa;

	lut_sub lut_2005 ({i_11_, i_36_, g30, i_12_, g232}, g237);
	defparam lut_2005.LUT_SIZE = 5;
	defparam lut_2005.mask = 32'h11115111;

	lut_sub lut_2021 ({i_39_, g30, g22, g45, g232}, g238);
	defparam lut_2021.LUT_SIZE = 5;
	defparam lut_2021.mask = 32'h8ccc0000;

	lut_sub lut_2034 ({i_36_, g11, i_16_, g237, g238}, g239);
	defparam lut_2034.LUT_SIZE = 5;
	defparam lut_2034.mask = 32'h00200000;

	lut_sub lut_2043 ({g56, g183, g231, g236, g239}, g240);
	defparam lut_2043.LUT_SIZE = 5;
	defparam lut_2043.mask = 32'hf0f02000;

	lut_sub lut_2057 ({g10, i_2_, i_1_, i_0_, g67}, g241);
	defparam lut_2057.LUT_SIZE = 5;
	defparam lut_2057.mask = 32'h32330000;

	lut_sub lut_2070 ({i_37_, i_32_, i_25_, g69, g226, g241}, g242);
	defparam lut_2070.LUT_SIZE = 6;
	defparam lut_2070.mask = 64'h3300330037053300;

	lut_sub lut_2094 ({i_22_, g125, i_21_, g198}, g243);
	defparam lut_2094.LUT_SIZE = 4;
	defparam lut_2094.mask = 16'h0504;

	lut_sub lut_2102 ({i_37_, i_38_, g187, g243}, g244);
	defparam lut_2102.LUT_SIZE = 4;
	defparam lut_2102.mask = 16'h1151;

	lut_sub lut_2111 ({i_37_, i_38_, i_39_, i_40_, g92}, g245);
	defparam lut_2111.LUT_SIZE = 5;
	defparam lut_2111.mask = 32'h40cf3000;

	lut_sub lut_2125 ({g27, g115}, g246);
	defparam lut_2125.LUT_SIZE = 2;
	defparam lut_2125.mask = 4'b0001;

	lut_sub lut_2132 ({i_13_, g45, g76, g246}, g247);
	defparam lut_2132.LUT_SIZE = 4;
	defparam lut_2132.mask = 16'ha8aa;

	lut_sub lut_2142 ({i_5_, i_12_, i_13_, i_15_}, g248);
	defparam lut_2142.LUT_SIZE = 4;
	defparam lut_2142.mask = 16'hd800;

	lut_sub lut_2154 ({g106, g202, g165, g247, g248}, g249);
	defparam lut_2154.LUT_SIZE = 5;
	defparam lut_2154.mask = 32'h0000444f;

	lut_sub lut_2165 ({i_37_, i_38_, i_39_, i_34_, g51}, g250);
	defparam lut_2165.LUT_SIZE = 5;
	defparam lut_2165.mask = 32'h00054000;

	lut_sub lut_2172 ({i_2_, i_1_, g49, i_0_}, g251);
	defparam lut_2172.LUT_SIZE = 4;
	defparam lut_2172.mask = 16'h0040;

	lut_sub lut_2177 ({i_11_, g122, i_5_, i_12_, i_15_}, g252);
	defparam lut_2177.LUT_SIZE = 5;
	defparam lut_2177.mask = 32'h10004000;

	lut_sub lut_2183 ({i_36_, i_37_, i_40_, i_32_, g67}, g253);
	defparam lut_2183.LUT_SIZE = 5;
	defparam lut_2183.mask = 32'h40000000;

	lut_sub lut_2191 ({g250, g251, g252, g253}, g254);
	defparam lut_2191.LUT_SIZE = 4;
	defparam lut_2191.mask = 16'h0537;

	lut_sub lut_2202 ({i_33_, g51}, g255);
	defparam lut_2202.LUT_SIZE = 2;
	defparam lut_2202.mask = 4'b1110;

	lut_sub lut_2210 ({i_12_, g11, i_17_, g232}, g256);
	defparam lut_2210.LUT_SIZE = 4;
	defparam lut_2210.mask = 16'h0004;

	lut_sub lut_2216 ({i_32_, i_5_, g24, g37}, g257);
	defparam lut_2216.LUT_SIZE = 4;
	defparam lut_2216.mask = 16'h1000;

	lut_sub lut_2226 ({g56, g46, g113, g255, g256, g257}, g258);
	defparam lut_2226.LUT_SIZE = 6;
	defparam lut_2226.mask = 64'h0050005000507777;

	lut_sub lut_2253 ({g134, g244, g245, g249, g254, g258}, g259);
	defparam lut_2253.LUT_SIZE = 6;
	defparam lut_2253.mask = 64'h8080000080000000;

	lut_sub lut_2259 ({i_38_, i_39_, i_40_}, g260);
	defparam lut_2259.LUT_SIZE = 3;
	defparam lut_2259.mask = 8'h02;

	lut_sub lut_2265 ({g51, i_31_, i_5_, i_9_, g260, i_14_}, g261);
	defparam lut_2265.LUT_SIZE = 6;
	defparam lut_2265.mask = 64'h000000003000ba00;

	lut_sub lut_2275 ({i_36_, i_37_, i_38_, i_39_, i_40_, i_35_}, g262);
	defparam lut_2275.LUT_SIZE = 6;
	defparam lut_2275.mask = 64'h0000440000142e0a;

	lut_sub lut_2293 ({g65, g175, g740, g261, g262}, g263);
	defparam lut_2293.LUT_SIZE = 5;
	defparam lut_2293.mask = 32'h0000fff7;

	lut_sub lut_2312 ({i_37_, i_38_, g65, i_5_}, g264);
	defparam lut_2312.LUT_SIZE = 4;
	defparam lut_2312.mask = 16'h0020;

	lut_sub lut_2319 ({i_37_, g115, g125, i_0_, g264}, g265);
	defparam lut_2319.LUT_SIZE = 5;
	defparam lut_2319.mask = 32'h00550057;

	lut_sub lut_2332 ({g260, i_21_, i_23_}, g266);
	defparam lut_2332.LUT_SIZE = 3;
	defparam lut_2332.mask = 8'h0e;

	lut_sub lut_2339 ({g122, i_22_, i_21_}, g267);
	defparam lut_2339.LUT_SIZE = 3;
	defparam lut_2339.mask = 8'he0;

	lut_sub lut_2347 ({i_40_, i_32_, i_16_, g215, g255}, g268);
	defparam lut_2347.LUT_SIZE = 5;
	defparam lut_2347.mask = 32'h20000000;

	lut_sub lut_2353 ({g22, i_15_, g232}, g269);
	defparam lut_2353.LUT_SIZE = 3;
	defparam lut_2353.mask = 8'h10;

	lut_sub lut_2360 ({i_18_, g152, i_21_, g268, g269}, g270);
	defparam lut_2360.LUT_SIZE = 5;
	defparam lut_2360.mask = 32'h51111111;

	lut_sub lut_2377 ({g198, g263, g265, g729, g270}, g271);
	defparam lut_2377.LUT_SIZE = 5;
	defparam lut_2377.mask = 32'ha0002000;

	lut_sub lut_2385 ({i_24_, g125, g198}, g272);
	defparam lut_2385.LUT_SIZE = 3;
	defparam lut_2385.mask = 8'h10;

	lut_sub lut_2389 ({i_30_, i_28_, i_29_}, g273);
	defparam lut_2389.LUT_SIZE = 3;
	defparam lut_2389.mask = 8'h80;

	lut_sub lut_2394 ({i_37_, i_38_, i_39_, g232}, g274);
	defparam lut_2394.LUT_SIZE = 4;
	defparam lut_2394.mask = 16'h0001;

	lut_sub lut_2398 ({i_36_, i_38_, i_39_}, g275);
	defparam lut_2398.LUT_SIZE = 3;
	defparam lut_2398.mask = 8'h10;

	lut_sub lut_2404 ({i_12_, i_15_, i_17_, g232, g275}, g276);
	defparam lut_2404.LUT_SIZE = 5;
	defparam lut_2404.mask = 32'h00000010;

	lut_sub lut_2412 ({g131, g163, g274, g276}, g277);
	defparam lut_2412.LUT_SIZE = 4;
	defparam lut_2412.mask = 16'h8880;

	lut_sub lut_2421 ({i_5_, g105, g273, g277}, g278);
	defparam lut_2421.LUT_SIZE = 4;
	defparam lut_2421.mask = 16'h5155;

	lut_sub lut_2434 ({g102, i_10_, i_27_, g73, g216}, g279);
	defparam lut_2434.LUT_SIZE = 5;
	defparam lut_2434.mask = 32'h00000001;

	lut_sub lut_2440 ({i_36_, g10, g116}, g280);
	defparam lut_2440.LUT_SIZE = 3;
	defparam lut_2440.mask = 8'h04;

	lut_sub lut_2445 ({i_36_, g14}, g281);
	defparam lut_2445.LUT_SIZE = 2;
	defparam lut_2445.mask = 4'b0100;

	lut_sub lut_2450 ({i_32_, i_2_, i_1_, i_0_, g67}, g282);
	defparam lut_2450.LUT_SIZE = 5;
	defparam lut_2450.mask = 32'h00100000;

	lut_sub lut_2458 ({g49, g280, g281, g282}, g283);
	defparam lut_2458.LUT_SIZE = 4;
	defparam lut_2458.mask = 16'h1505;

	lut_sub lut_2470 ({g21, g47, g130, g184}, g284);
	defparam lut_2470.LUT_SIZE = 4;
	defparam lut_2470.mask = 16'h5545;

	lut_sub lut_2485 ({g112, g272, g279, g283, g284}, g285);
	defparam lut_2485.LUT_SIZE = 5;
	defparam lut_2485.mask = 32'h40404000;

	lut_sub lut_2496 ({g102, g14, g272, g278, g285}, g286);
	defparam lut_2496.LUT_SIZE = 5;
	defparam lut_2496.mask = 32'h55501110;

	lut_sub lut_2513 ({g240, g242, g259, g271, g286}, g287);
	defparam lut_2513.LUT_SIZE = 5;
	defparam lut_2513.mask = 32'h00000100;

	lut_sub lut_2517 ({i_7_, i_5_, i_30_, i_28_, i_29_}, g288);
	defparam lut_2517.LUT_SIZE = 5;
	defparam lut_2517.mask = 32'h9b000000;

	lut_sub lut_2527 ({g1, i_30_, i_29_, g288}, g289);
	defparam lut_2527.LUT_SIZE = 4;
	defparam lut_2527.mask = 16'h8aaa;

	lut_sub lut_2540 ({g65, g1, i_15_, i_24_, g151}, g290);
	defparam lut_2540.LUT_SIZE = 5;
	defparam lut_2540.mask = 32'h00005100;

	lut_sub lut_2551 ({g122, g139, g119, g289, g290}, g291);
	defparam lut_2551.LUT_SIZE = 5;
	defparam lut_2551.mask = 32'h0c5d0055;

	lut_sub lut_2568 ({i_9_, i_18_, g153, g144, g165}, g292);
	defparam lut_2568.LUT_SIZE = 5;
	defparam lut_2568.mask = 32'h00010101;

	lut_sub lut_2576 ({i_36_, g56, g48}, g293);
	defparam lut_2576.LUT_SIZE = 3;
	defparam lut_2576.mask = 8'h10;

	lut_sub lut_2584 ({g102, g1, g105, g273}, g294);
	defparam lut_2584.LUT_SIZE = 4;
	defparam lut_2584.mask = 16'h0010;

	lut_sub lut_2591 ({i_31_, i_5_, g24, g293, g294}, g295);
	defparam lut_2591.LUT_SIZE = 5;
	defparam lut_2591.mask = 32'haaaaa8aa;

	lut_sub lut_2613 ({i_40_, g117, g95, g8, g215}, g296);
	defparam lut_2613.LUT_SIZE = 5;
	defparam lut_2613.mask = 32'h07ff0000;

	lut_sub lut_2629 ({g1, i_12_, i_15_, g194}, g297);
	defparam lut_2629.LUT_SIZE = 4;
	defparam lut_2629.mask = 16'h5400;

	lut_sub lut_2639 ({g57, g130, g8, g297}, g298);
	defparam lut_2639.LUT_SIZE = 4;
	defparam lut_2639.mask = 16'haaa8;

	lut_sub lut_2651 ({i_37_, i_38_, i_39_, i_40_, g93, g96}, g299);
	defparam lut_2651.LUT_SIZE = 6;
	defparam lut_2651.mask = 64'h0550030000500300;

	lut_sub lut_2669 ({g292, g295, g296, g298, g299}, g300);
	defparam lut_2669.LUT_SIZE = 5;
	defparam lut_2669.mask = 32'h00200000;

	lut_sub lut_2675 ({g122, g1, i_13_, i_15_}, g301);
	defparam lut_2675.LUT_SIZE = 4;
	defparam lut_2675.mask = 16'h8000;

	lut_sub lut_2684 ({g2, g45, g128, g98, g301}, g302);
	defparam lut_2684.LUT_SIZE = 5;
	defparam lut_2684.mask = 32'h000f111f;

	lut_sub lut_2701 ({i_36_, g100, g10, g48, i_25_, i_26_}, g303);
	defparam lut_2701.LUT_SIZE = 6;
	defparam lut_2701.mask = 64'h0000000000000b00;

	lut_sub lut_2709 ({i_7_, g102, i_10_, i_27_, g216}, g304);
	defparam lut_2709.LUT_SIZE = 5;
	defparam lut_2709.mask = 32'h00540000;

	lut_sub lut_2718 ({i_40_, i_34_, g6, g78, g225}, g305);
	defparam lut_2718.LUT_SIZE = 5;
	defparam lut_2718.mask = 32'h00010000;

	lut_sub lut_2725 ({i_38_, g101, i_35_, g70, g163}, g306);
	defparam lut_2725.LUT_SIZE = 5;
	defparam lut_2725.mask = 32'h00100000;

	lut_sub lut_2730 ({i_7_, i_33_, g11}, g307);
	defparam lut_2730.LUT_SIZE = 3;
	defparam lut_2730.mask = 8'h10;

	lut_sub lut_2735 ({i_5_, g22, i_16_, i_17_, i_9_}, g308);
	defparam lut_2735.LUT_SIZE = 5;
	defparam lut_2735.mask = 32'h17000000;

	lut_sub lut_2747 ({g2, g21, g113, g307, g308}, g309);
	defparam lut_2747.LUT_SIZE = 5;
	defparam lut_2747.mask = 32'h00000111;

	lut_sub lut_2756 ({i_37_, i_35_, g65, g21, g79}, g310);
	defparam lut_2756.LUT_SIZE = 5;
	defparam lut_2756.mask = 32'h08000c00;

	lut_sub lut_2763 ({i_36_, i_31_, g1}, g311);
	defparam lut_2763.LUT_SIZE = 3;
	defparam lut_2763.mask = 8'h20;

	lut_sub lut_2771 ({g102, i_9_, g171, g310, g311}, g312);
	defparam lut_2771.LUT_SIZE = 5;
	defparam lut_2771.mask = 32'h11115111;

	lut_sub lut_2788 ({g201, g305, g306, g309, g312}, g313);
	defparam lut_2788.LUT_SIZE = 5;
	defparam lut_2788.mask = 32'h8000a000;

	lut_sub lut_2798 ({i_39_, i_40_, g302, g303, g304, g313}, g314);
	defparam lut_2798.LUT_SIZE = 6;
	defparam lut_2798.mask = 64'h4040400055555500;

	lut_sub lut_2817 ({i_40_, g8}, g315);
	defparam lut_2817.LUT_SIZE = 2;
	defparam lut_2817.mask = 4'b0001;

	lut_sub lut_2822 ({i_37_, i_38_, i_39_, i_40_, g121}, g316);
	defparam lut_2822.LUT_SIZE = 5;
	defparam lut_2822.mask = 32'h00004140;

	lut_sub lut_2830 ({i_36_, i_37_, i_34_, g77, g316}, g317);
	defparam lut_2830.LUT_SIZE = 5;
	defparam lut_2830.mask = 32'haaaa8aaa;

	lut_sub lut_2850 ({i_37_, g260, g5}, g318);
	defparam lut_2850.LUT_SIZE = 3;
	defparam lut_2850.mask = 8'h01;

	lut_sub lut_2858 ({g61, g92, g160, g318}, g319);
	defparam lut_2858.LUT_SIZE = 4;
	defparam lut_2858.mask = 16'h0537;

	lut_sub lut_2872 ({i_34_, g78, g315, g317, g319}, g320);
	defparam lut_2872.LUT_SIZE = 5;
	defparam lut_2872.mask = 32'h22202222;

	lut_sub lut_2884 ({i_7_, i_33_, i_32_, g150, g320}, g321);
	defparam lut_2884.LUT_SIZE = 5;
	defparam lut_2884.mask = 32'h33133333;

	lut_sub lut_2905 ({i_36_, g100, g101, g102, i_13_}, g322);
	defparam lut_2905.LUT_SIZE = 5;
	defparam lut_2905.mask = 32'h00020000;

	lut_sub lut_2911 ({i_39_, i_32_, i_13_, g45, g49}, g323);
	defparam lut_2911.LUT_SIZE = 5;
	defparam lut_2911.mask = 32'h00000200;

	lut_sub lut_2919 ({i_40_, g125, g225, g322, g323}, g324);
	defparam lut_2919.LUT_SIZE = 5;
	defparam lut_2919.mask = 32'h88888880;

	lut_sub lut_2932 ({g23, g18, i_18_, g155, i_19_}, g325);
	defparam lut_2932.LUT_SIZE = 5;
	defparam lut_2932.mask = 32'h00130517;

	lut_sub lut_2948 ({g57, g125, i_23_, g153, g325}, g326);
	defparam lut_2948.LUT_SIZE = 5;
	defparam lut_2948.mask = 32'h000100ff;

	lut_sub lut_2964 ({i_37_, g30, g54, g324, g326}, g327);
	defparam lut_2964.LUT_SIZE = 5;
	defparam lut_2964.mask = 32'h0c0c5d0c;

	lut_sub lut_2983 ({g291, g300, g314, g321, g327}, g328);
	defparam lut_2983.LUT_SIZE = 5;
	defparam lut_2983.mask = 32'h00020000;

	lut_sub lut_2990 ({g25, g136, g79}, g329);
	defparam lut_2990.LUT_SIZE = 3;
	defparam lut_2990.mask = 8'h01;

	lut_sub lut_2995 ({i_7_, i_2_, i_1_, i_0_, g67}, g330);
	defparam lut_2995.LUT_SIZE = 5;
	defparam lut_2995.mask = 32'h00100000;

	lut_sub lut_3001 ({i_38_, g66, g330}, g331);
	defparam lut_3001.LUT_SIZE = 3;
	defparam lut_3001.mask = 8'h01;

	lut_sub lut_3008 ({g124, g148, g331}, g332);
	defparam lut_3008.LUT_SIZE = 3;
	defparam lut_3008.mask = 8'ha8;

	lut_sub lut_3016 ({i_32_, g54, i_13_, g10}, g333);
	defparam lut_3016.LUT_SIZE = 4;
	defparam lut_3016.mask = 16'h0800;

	lut_sub lut_3023 ({i_36_, g100, g76, g333}, g334);
	defparam lut_3023.LUT_SIZE = 4;
	defparam lut_3023.mask = 16'h0100;

	lut_sub lut_3030 ({i_31_, g54, i_13_, g180, g334}, g335);
	defparam lut_3030.LUT_SIZE = 5;
	defparam lut_3030.mask = 32'haaa8aaaa;

	lut_sub lut_3049 ({g138, i_30_, i_29_}, g336);
	defparam lut_3049.LUT_SIZE = 3;
	defparam lut_3049.mask = 8'h08;

	lut_sub lut_3058 ({g1, g44, g46, g105, g336}, g337);
	defparam lut_3058.LUT_SIZE = 5;
	defparam lut_3058.mask = 32'h111f000f;

	lut_sub lut_3074 ({i_38_, g51, g76}, g338);
	defparam lut_3074.LUT_SIZE = 3;
	defparam lut_3074.mask = 8'h01;

	lut_sub lut_3081 ({g53, g107, g338}, g339);
	defparam lut_3081.LUT_SIZE = 3;
	defparam lut_3081.mask = 8'h01;

	lut_sub lut_3086 ({i_36_, i_38_, i_39_, g92}, g340);
	defparam lut_3086.LUT_SIZE = 4;
	defparam lut_3086.mask = 16'h0ece;

	lut_sub lut_3097 ({i_36_, i_37_, i_38_, i_35_}, g341);
	defparam lut_3097.LUT_SIZE = 4;
	defparam lut_3097.mask = 16'h054d;

	lut_sub lut_3108 ({i_37_, i_40_, i_34_, g6, g341}, g342);
	defparam lut_3108.LUT_SIZE = 5;
	defparam lut_3108.mask = 32'h10101000;

	lut_sub lut_3116 ({i_37_, i_39_, i_40_, g7, g95}, g343);
	defparam lut_3116.LUT_SIZE = 5;
	defparam lut_3116.mask = 32'h00350000;

	lut_sub lut_3128 ({g303, g339, g340, g342, g343}, g344);
	defparam lut_3128.LUT_SIZE = 5;
	defparam lut_3128.mask = 32'h8a000000;

	lut_sub lut_3139 ({g329, g332, g335, g337, g344}, g345);
	defparam lut_3139.LUT_SIZE = 5;
	defparam lut_3139.mask = 32'h00040000;

	lut_sub lut_3144 ({i_37_, g104}, g346);
	defparam lut_3144.LUT_SIZE = 2;
	defparam lut_3144.mask = 4'b0001;

	lut_sub lut_3150 ({i_38_, g70, g78}, g347);
	defparam lut_3150.LUT_SIZE = 3;
	defparam lut_3150.mask = 8'h01;

	lut_sub lut_3158 ({g47, i_0_, g93, g346, g347}, g348);
	defparam lut_3158.LUT_SIZE = 5;
	defparam lut_3158.mask = 32'h03570303;

	lut_sub lut_3175 ({i_37_, i_38_, i_39_, g121, g148, g301}, g349);
	defparam lut_3175.LUT_SIZE = 6;
	defparam lut_3175.mask = 64'hfaffccffffffffcc;

	lut_sub lut_3233 ({i_33_, i_32_, g51, i_31_}, g350);
	defparam lut_3233.LUT_SIZE = 4;
	defparam lut_3233.mask = 16'h0020;

	lut_sub lut_3240 ({i_36_, g162, g48, g98}, g351);
	defparam lut_3240.LUT_SIZE = 4;
	defparam lut_3240.mask = 16'h0010;

	lut_sub lut_3248 ({i_40_, g44, g281, g95, g215}, g352);
	defparam lut_3248.LUT_SIZE = 5;
	defparam lut_3248.mask = 32'heee00000;

	lut_sub lut_3261 ({i_37_, i_38_, i_35_, g65}, g353);
	defparam lut_3261.LUT_SIZE = 4;
	defparam lut_3261.mask = 16'h0010;

	lut_sub lut_3270 ({g57, g68, g215, g350, g353}, g354);
	defparam lut_3270.LUT_SIZE = 5;
	defparam lut_3270.mask = 32'h00550357;

	lut_sub lut_3286 ({g10, g11, i_21_}, g355);
	defparam lut_3286.LUT_SIZE = 3;
	defparam lut_3286.mask = 8'h20;

	lut_sub lut_3292 ({i_11_, g1, i_12_, g355}, g356);
	defparam lut_3292.LUT_SIZE = 4;
	defparam lut_3292.mask = 16'h1050;

	lut_sub lut_3302 ({i_11_, g1, g28, g12, g356}, g357);
	defparam lut_3302.LUT_SIZE = 5;
	defparam lut_3302.mask = 32'h05050705;

	lut_sub lut_3319 ({g348, g723, g352, g354, g357}, g358);
	defparam lut_3319.LUT_SIZE = 5;
	defparam lut_3319.mask = 32'h08aa0808;

	lut_sub lut_3331 ({i_11_, g1, g37, i_14_}, g359);
	defparam lut_3331.LUT_SIZE = 4;
	defparam lut_3331.mask = 16'h0020;

	lut_sub lut_3340 ({g2, g21, g136, g79, g359}, g360);
	defparam lut_3340.LUT_SIZE = 5;
	defparam lut_3340.mask = 32'h01010155;

	lut_sub lut_3351 ({g1, i_30_, i_28_, i_29_}, g361);
	defparam lut_3351.LUT_SIZE = 4;
	defparam lut_3351.mask = 16'h80a0;

	lut_sub lut_3359 ({i_37_, i_38_, i_34_, g1, g361}, g362);
	defparam lut_3359.LUT_SIZE = 5;
	defparam lut_3359.mask = 32'h00008000;

	lut_sub lut_3368 ({g100, g104, g72, g73, g96}, g363);
	defparam lut_3368.LUT_SIZE = 5;
	defparam lut_3368.mask = 32'h000f444f;

	lut_sub lut_3387 ({g3, g115, g360, g362, g363}, g364);
	defparam lut_3387.LUT_SIZE = 5;
	defparam lut_3387.mask = 32'haaaaa080;

	lut_sub lut_3403 ({g122, g1, i_9_, i_18_, i_21_}, g365);
	defparam lut_3403.LUT_SIZE = 5;
	defparam lut_3403.mask = 32'h80000000;

	lut_sub lut_3410 ({g26, g37, g365}, g366);
	defparam lut_3410.LUT_SIZE = 3;
	defparam lut_3410.mask = 8'h15;

	lut_sub lut_3420 ({g122, g121, i_21_, g91, g366}, g367);
	defparam lut_3420.LUT_SIZE = 5;
	defparam lut_3420.mask = 32'h00750055;

	lut_sub lut_3435 ({i_37_, g10, g48, g115, i_0_}, g368);
	defparam lut_3435.LUT_SIZE = 5;
	defparam lut_3435.mask = 32'h00000100;

	lut_sub lut_3441 ({i_11_, g1, i_12_, g12}, g369);
	defparam lut_3441.LUT_SIZE = 4;
	defparam lut_3441.mask = 16'h1050;

	lut_sub lut_3451 ({i_40_, g14, g356, g368, g369}, g370);
	defparam lut_3451.LUT_SIZE = 5;
	defparam lut_3451.mask = 32'hcc80cc88;

	lut_sub lut_3469 ({i_38_, g3, i_16_, g34, g18, g73}, g371);
	defparam lut_3469.LUT_SIZE = 6;
	defparam lut_3469.mask = 64'h0000000000000100;

	lut_sub lut_3476 ({g1, i_15_, g3, g131}, g372);
	defparam lut_3476.LUT_SIZE = 4;
	defparam lut_3476.mask = 16'h1000;

	lut_sub lut_3483 ({i_38_, g197, g330, g372}, g373);
	defparam lut_3483.LUT_SIZE = 4;
	defparam lut_3483.mask = 16'ha8aa;

	lut_sub lut_3494 ({i_15_, i_21_, i_23_, g211}, g374);
	defparam lut_3494.LUT_SIZE = 4;
	defparam lut_3494.mask = 16'h0040;

	lut_sub lut_3499 ({i_22_, g11, i_21_}, g375);
	defparam lut_3499.LUT_SIZE = 3;
	defparam lut_3499.mask = 8'h32;

	lut_sub lut_3507 ({i_36_, g49, g131}, g376);
	defparam lut_3507.LUT_SIZE = 3;
	defparam lut_3507.mask = 8'h40;

	lut_sub lut_3515 ({g143, g61, i_23_, g375, g376}, g377);
	defparam lut_3515.LUT_SIZE = 5;
	defparam lut_3515.mask = 32'h111111f1;

	lut_sub lut_3535 ({g43, g136, g371, g373, g374, g377}, g378);
	defparam lut_3535.LUT_SIZE = 6;
	defparam lut_3535.mask = 64'hffff0f0088880800;

	lut_sub lut_3567 ({i_36_, g21, g367, g370, g378}, g379);
	defparam lut_3567.LUT_SIZE = 5;
	defparam lut_3567.mask = 32'h11105550;

	lut_sub lut_3584 ({g64, g345, g358, g364, g379}, o_5_);
	defparam lut_3584.LUT_SIZE = 5;
	defparam lut_3584.mask = 32'hfffffffe;

	lut_sub lut_3620 ({i_15_, g31, g98}, g381);
	defparam lut_3620.LUT_SIZE = 3;
	defparam lut_3620.mask = 8'h10;

	lut_sub lut_3627 ({i_11_, g95, g346, g351}, g382);
	defparam lut_3627.LUT_SIZE = 4;
	defparam lut_3627.mask = 16'h0357;

	lut_sub lut_3641 ({i_40_, g45, g333, g381, g382}, g383);
	defparam lut_3641.LUT_SIZE = 5;
	defparam lut_3641.mask = 32'h0000777f;

	lut_sub lut_3659 ({i_40_, g105, g8}, g384);
	defparam lut_3659.LUT_SIZE = 3;
	defparam lut_3659.mask = 8'h8c;

	lut_sub lut_3665 ({i_11_, i_12_}, g385);
	defparam lut_3665.LUT_SIZE = 2;
	defparam lut_3665.mask = 4'b0001;

	lut_sub lut_3669 ({i_36_, i_37_, i_38_, i_39_, i_40_}, g386);
	defparam lut_3669.LUT_SIZE = 5;
	defparam lut_3669.mask = 32'h10400000;

	lut_sub lut_3679 ({g54, g155, g385, g246, g386}, g387);
	defparam lut_3679.LUT_SIZE = 5;
	defparam lut_3679.mask = 32'h00305575;

	lut_sub lut_3697 ({g102, i_31_, g288, g384, g387}, g388);
	defparam lut_3697.LUT_SIZE = 5;
	defparam lut_3697.mask = 32'h00005d00;

	lut_sub lut_3707 ({i_22_, i_24_, i_23_, g182, g325}, g389);
	defparam lut_3707.LUT_SIZE = 5;
	defparam lut_3707.mask = 32'h00000001;

	lut_sub lut_3712 ({i_22_, g23, i_21_}, g390);
	defparam lut_3712.LUT_SIZE = 3;
	defparam lut_3712.mask = 8'h01;

	lut_sub lut_3719 ({i_37_, g5, g6, g77}, g391);
	defparam lut_3719.LUT_SIZE = 4;
	defparam lut_3719.mask = 16'h0100;

	lut_sub lut_3725 ({i_32_, g28, g10, i_24_, i_23_}, g392);
	defparam lut_3725.LUT_SIZE = 5;
	defparam lut_3725.mask = 32'h00100000;

	lut_sub lut_3731 ({i_38_, g5, g6}, g393);
	defparam lut_3731.LUT_SIZE = 3;
	defparam lut_3731.mask = 8'h10;

	lut_sub lut_3737 ({i_36_, i_37_, i_39_, i_40_, g7, g393}, g394);
	defparam lut_3737.LUT_SIZE = 6;
	defparam lut_3737.mask = 64'h0030005555750000;

	lut_sub lut_3757 ({i_37_, g14, g5}, g395);
	defparam lut_3757.LUT_SIZE = 3;
	defparam lut_3757.mask = 8'h10;

	lut_sub lut_3765 ({i_24_, g123, g144, g199, g395}, g396);
	defparam lut_3765.LUT_SIZE = 5;
	defparam lut_3765.mask = 32'h00550357;

	lut_sub lut_3784 ({g390, g391, g392, g394, g396}, g397);
	defparam lut_3784.LUT_SIZE = 5;
	defparam lut_3784.mask = 32'h88008000;

	lut_sub lut_3790 ({i_37_, i_38_, i_39_, i_40_}, g398);
	defparam lut_3790.LUT_SIZE = 4;
	defparam lut_3790.mask = 16'h060e;

	lut_sub lut_3801 ({g101, g45, g49}, g399);
	defparam lut_3801.LUT_SIZE = 3;
	defparam lut_3801.mask = 8'h02;

	lut_sub lut_3807 ({i_32_, g54, i_13_, g399}, g400);
	defparam lut_3807.LUT_SIZE = 4;
	defparam lut_3807.mask = 16'h0400;

	lut_sub lut_3812 ({i_37_, i_38_, i_39_, i_40_, g51}, g401);
	defparam lut_3812.LUT_SIZE = 5;
	defparam lut_3812.mask = 32'h15015100;

	lut_sub lut_3827 ({i_40_, g55, g148, g8, g189, g401}, g402);
	defparam lut_3827.LUT_SIZE = 6;
	defparam lut_3827.mask = 64'h000f777f00007777;

	lut_sub lut_3862 ({i_15_, g138, g155, g246}, g403);
	defparam lut_3862.LUT_SIZE = 4;
	defparam lut_3862.mask = 16'h0100;

	lut_sub lut_3870 ({i_37_, g122, g57, g76, g5}, g404);
	defparam lut_3870.LUT_SIZE = 5;
	defparam lut_3870.mask = 32'h01000000;

	lut_sub lut_3876 ({g1, g22, i_9_, i_18_, i_21_}, g405);
	defparam lut_3876.LUT_SIZE = 5;
	defparam lut_3876.mask = 32'h7f000000;

	lut_sub lut_3886 ({i_37_, i_38_, i_40_, i_15_}, g406);
	defparam lut_3886.LUT_SIZE = 4;
	defparam lut_3886.mask = 16'h0100;

	lut_sub lut_3893 ({i_22_, i_24_, g125, g405, g406}, g407);
	defparam lut_3893.LUT_SIZE = 5;
	defparam lut_3893.mask = 32'h00000001;

	lut_sub lut_3900 ({g47, g48, g49}, g408);
	defparam lut_3900.LUT_SIZE = 3;
	defparam lut_3900.mask = 8'h02;

	lut_sub lut_3904 ({i_36_, i_37_, i_38_, i_39_, i_40_}, g409);
	defparam lut_3904.LUT_SIZE = 5;
	defparam lut_3904.mask = 32'h79d00000;

	lut_sub lut_3919 ({g58, g165, g408, g409}, g410);
	defparam lut_3919.LUT_SIZE = 4;
	defparam lut_3919.mask = 16'h0357;

	lut_sub lut_3934 ({i_40_, g28, g128, g199, g225, g333}, g411);
	defparam lut_3934.LUT_SIZE = 6;
	defparam lut_3934.mask = 64'h111f555f000f555f;

	lut_sub lut_3973 ({g403, g404, g407, g410, g411}, g412);
	defparam lut_3973.LUT_SIZE = 5;
	defparam lut_3973.mask = 32'h80000000;

	lut_sub lut_3982 ({g93, g398, g400, g402, g412}, g413);
	defparam lut_3982.LUT_SIZE = 5;
	defparam lut_3982.mask = 32'h40404000;

	lut_sub lut_3990 ({i_15_, g31, g124}, g414);
	defparam lut_3990.LUT_SIZE = 3;
	defparam lut_3990.mask = 8'h10;

	lut_sub lut_3997 ({g131, g219, g390}, g415);
	defparam lut_3997.LUT_SIZE = 3;
	defparam lut_3997.mask = 8'h01;

	lut_sub lut_4004 ({g1, g138, i_30_, i_29_, g384}, g416);
	defparam lut_4004.LUT_SIZE = 5;
	defparam lut_4004.mask = 32'h00200000;

	lut_sub lut_4009 ({i_36_, i_37_, i_38_, i_39_, i_40_, g5}, g417);
	defparam lut_4009.LUT_SIZE = 6;
	defparam lut_4009.mask = 64'h4005110040000000;

	lut_sub lut_4022 ({g94, g315, g301, g417}, g418);
	defparam lut_4022.LUT_SIZE = 4;
	defparam lut_4022.mask = 16'h1311;

	lut_sub lut_4034 ({i_37_, g30, g121, g123, g418}, g419);
	defparam lut_4034.LUT_SIZE = 5;
	defparam lut_4034.mask = 32'haaaaa8aa;

	lut_sub lut_4058 ({g73, g304, g414, g415, g416, g419}, g420);
	defparam lut_4058.LUT_SIZE = 6;
	defparam lut_4058.mask = 64'h4000400040000000;

	lut_sub lut_4070 ({g383, g388, g389, g397, g413, g420}, g421);
	defparam lut_4070.LUT_SIZE = 6;
	defparam lut_4070.mask = 64'h0100000000000000;

	lut_sub lut_4075 ({i_11_, i_12_, g103}, g422);
	defparam lut_4075.LUT_SIZE = 3;
	defparam lut_4075.mask = 8'h10;

	lut_sub lut_4081 ({g65, i_22_, i_24_, i_21_, g198}, g423);
	defparam lut_4081.LUT_SIZE = 5;
	defparam lut_4081.mask = 32'h00000001;

	lut_sub lut_4089 ({g151, g79, g187, g423}, g424);
	defparam lut_4089.LUT_SIZE = 4;
	defparam lut_4089.mask = 16'h0015;

	lut_sub lut_4096 ({i_5_, i_9_, g18, i_18_, i_19_}, g425);
	defparam lut_4096.LUT_SIZE = 5;
	defparam lut_4096.mask = 32'h010f0000;

	lut_sub lut_4104 ({i_24_, i_18_, i_23_, i_19_}, g426);
	defparam lut_4104.LUT_SIZE = 4;
	defparam lut_4104.mask = 16'h0013;

	lut_sub lut_4113 ({g112, i_24_, g125, i_21_, i_23_, g198}, g427);
	defparam lut_4113.LUT_SIZE = 6;
	defparam lut_4113.mask = 64'h0000000000000001;

	lut_sub lut_4119 ({i_32_, i_21_, g198, g376}, g428);
	defparam lut_4119.LUT_SIZE = 4;
	defparam lut_4119.mask = 16'h0100;

	lut_sub lut_4128 ({g157, g425, g426, g427, g428}, g429);
	defparam lut_4128.LUT_SIZE = 5;
	defparam lut_4128.mask = 32'h88888880;

	lut_sub lut_4141 ({i_5_, g45, g115, i_28_, g336}, g430);
	defparam lut_4141.LUT_SIZE = 5;
	defparam lut_4141.mask = 32'h00040000;

	lut_sub lut_4148 ({i_5_, g77, g273, g350}, g431);
	defparam lut_4148.LUT_SIZE = 4;
	defparam lut_4148.mask = 16'h0100;

	lut_sub lut_4154 ({g139, g83}, g432);
	defparam lut_4154.LUT_SIZE = 2;
	defparam lut_4154.mask = 4'b0001;

	lut_sub lut_4162 ({g136, g131, g104, g338}, g433);
	defparam lut_4162.LUT_SIZE = 4;
	defparam lut_4162.mask = 16'haa80;

	lut_sub lut_4174 ({g197, g423, g432, g433}, g434);
	defparam lut_4174.LUT_SIZE = 4;
	defparam lut_4174.mask = 16'h03ab;

	lut_sub lut_4188 ({i_22_, g429, g430, g431, g434}, g435);
	defparam lut_4188.LUT_SIZE = 5;
	defparam lut_4188.mask = 32'h80800080;

	lut_sub lut_4195 ({i_22_, i_24_, g222}, g436);
	defparam lut_4195.LUT_SIZE = 3;
	defparam lut_4195.mask = 8'h01;

	lut_sub lut_4201 ({i_38_, i_39_, i_40_, g65, g88}, g437);
	defparam lut_4201.LUT_SIZE = 5;
	defparam lut_4201.mask = 32'h00000110;

	lut_sub lut_4211 ({g65, g151, g79, g436, g437}, g438);
	defparam lut_4211.LUT_SIZE = 5;
	defparam lut_4211.mask = 32'haaaaaaa8;

	lut_sub lut_4234 ({g422, g424, g208, g435, g438}, g439);
	defparam lut_4234.LUT_SIZE = 5;
	defparam lut_4234.mask = 32'h01000000;

	lut_sub lut_4242 ({g77, g184, g219, g422}, g440);
	defparam lut_4242.LUT_SIZE = 4;
	defparam lut_4242.mask = 16'h0a08;

	lut_sub lut_4252 ({g84, g213, g208, g430}, g441);
	defparam lut_4252.LUT_SIZE = 4;
	defparam lut_4252.mask = 16'h2220;

	lut_sub lut_4260 ({i_36_, g100, g73}, g442);
	defparam lut_4260.LUT_SIZE = 3;
	defparam lut_4260.mask = 8'h10;

	lut_sub lut_4269 ({g10, g45, g76, g165, g442}, g443);
	defparam lut_4269.LUT_SIZE = 5;
	defparam lut_4269.mask = 32'h777f0000;

	lut_sub lut_4288 ({g11, g43, i_25_, i_20_, g443}, g444);
	defparam lut_4288.LUT_SIZE = 5;
	defparam lut_4288.mask = 32'h00000015;

	lut_sub lut_4296 ({i_24_, g152, g132, i_23_}, g445);
	defparam lut_4296.LUT_SIZE = 4;
	defparam lut_4296.mask = 16'hcc8c;

	lut_sub lut_4309 ({i_40_, g95, g98, g215}, g446);
	defparam lut_4309.LUT_SIZE = 4;
	defparam lut_4309.mask = 16'h0507;

	lut_sub lut_4320 ({i_25_, g390, i_20_, g445, g446}, g447);
	defparam lut_4320.LUT_SIZE = 5;
	defparam lut_4320.mask = 32'haaa2aa22;

	lut_sub lut_4338 ({i_22_, i_24_, i_21_, g444, g447}, o_10_);
	defparam lut_4338.LUT_SIZE = 5;
	defparam lut_4338.mask = 32'haaaaaaab;

	lut_sub lut_4362 ({i_31_, g1, g105, g106, g273}, g449);
	defparam lut_4362.LUT_SIZE = 5;
	defparam lut_4362.mask = 32'h01000000;

	lut_sub lut_4369 ({g56, g46, g165}, g450);
	defparam lut_4369.LUT_SIZE = 3;
	defparam lut_4369.mask = 8'h07;

	lut_sub lut_4377 ({i_11_, i_31_, i_12_, g11, g450}, g451);
	defparam lut_4377.LUT_SIZE = 5;
	defparam lut_4377.mask = 32'h01001000;

	lut_sub lut_4384 ({g1, i_16_, i_17_, i_9_, g451}, g452);
	defparam lut_4384.LUT_SIZE = 5;
	defparam lut_4384.mask = 32'h01150000;

	lut_sub lut_4397 ({g95, g99, g215, g292, g449, g452}, g453);
	defparam lut_4397.LUT_SIZE = 6;
	defparam lut_4397.mask = 64'h8080000080000000;

	lut_sub lut_4403 ({i_7_, i_5_, i_0_}, g454);
	defparam lut_4403.LUT_SIZE = 3;
	defparam lut_4403.mask = 8'h20;

	lut_sub lut_4409 ({i_37_, i_38_, i_40_, g160, g94}, g455);
	defparam lut_4409.LUT_SIZE = 5;
	defparam lut_4409.mask = 32'ha0000030;

	lut_sub lut_4419 ({g122, g454, i_8_, g455}, o_12_);
	defparam lut_4419.LUT_SIZE = 4;
	defparam lut_4419.mask = 16'h0100;

	lut_sub lut_4426 ({i_38_, i_39_, i_40_, g65, g151, g184}, g457);
	defparam lut_4426.LUT_SIZE = 6;
	defparam lut_4426.mask = 64'h5555555454555555;

	lut_sub lut_4463 ({g14, g65, g88, g457}, g458);
	defparam lut_4463.LUT_SIZE = 4;
	defparam lut_4463.mask = 16'h5554;

	lut_sub lut_4475 ({i_13_, g226, g457}, g459);
	defparam lut_4475.LUT_SIZE = 3;
	defparam lut_4475.mask = 8'h54;

	lut_sub lut_4482 ({i_37_, i_38_, i_39_, i_40_, g95}, g460);
	defparam lut_4482.LUT_SIZE = 5;
	defparam lut_4482.mask = 32'h00000004;

	lut_sub lut_4486 ({i_2_, i_1_, i_0_}, g461);
	defparam lut_4486.LUT_SIZE = 3;
	defparam lut_4486.mask = 8'h40;

	lut_sub lut_4491 ({i_3_, i_4_, g461}, g462);
	defparam lut_4491.LUT_SIZE = 3;
	defparam lut_4491.mask = 8'h40;

	lut_sub lut_4499 ({i_37_, g104, g78, g79, g462}, g463);
	defparam lut_4499.LUT_SIZE = 5;
	defparam lut_4499.mask = 32'h01010005;

	lut_sub lut_4511 ({g30, g22, g70, g71, g463}, g464);
	defparam lut_4511.LUT_SIZE = 5;
	defparam lut_4511.mask = 32'h05070505;

	lut_sub lut_4523 ({i_2_, i_1_, i_0_}, g465);
	defparam lut_4523.LUT_SIZE = 3;
	defparam lut_4523.mask = 8'h10;

	lut_sub lut_4529 ({i_7_, g67, g465}, g466);
	defparam lut_4529.LUT_SIZE = 3;
	defparam lut_4529.mask = 8'h10;

	lut_sub lut_4534 ({i_36_, i_40_, i_34_, i_35_, g6}, g467);
	defparam lut_4534.LUT_SIZE = 5;
	defparam lut_4534.mask = 32'h00104000;

	lut_sub lut_4544 ({g66, g187, g346, g466, g467}, g468);
	defparam lut_4544.LUT_SIZE = 5;
	defparam lut_4544.mask = 32'h05050537;

	lut_sub lut_4563 ({g148, g225, g460, g464, g468}, g469);
	defparam lut_4563.LUT_SIZE = 5;
	defparam lut_4563.mask = 32'h80808000;

	lut_sub lut_4570 ({i_37_, i_38_, i_39_, g51}, g470);
	defparam lut_4570.LUT_SIZE = 4;
	defparam lut_4570.mask = 16'h0001;

	lut_sub lut_4578 ({i_38_, g51, g115, g232, g470}, g471);
	defparam lut_4578.LUT_SIZE = 5;
	defparam lut_4578.mask = 32'h11111113;

	lut_sub lut_4591 ({i_37_, i_38_, i_39_, g51, i_17_}, g472);
	defparam lut_4591.LUT_SIZE = 5;
	defparam lut_4591.mask = 32'h00022002;

	lut_sub lut_4598 ({i_37_, i_38_, i_39_, i_40_, g51}, g473);
	defparam lut_4598.LUT_SIZE = 5;
	defparam lut_4598.mask = 32'h15455105;

	lut_sub lut_4616 ({i_16_, g269, g471, g472, g473}, g474);
	defparam lut_4616.LUT_SIZE = 5;
	defparam lut_4616.mask = 32'hf080f0c0;

	lut_sub lut_4633 ({i_36_, i_37_, i_38_, g67, g241, g251}, g475);
	defparam lut_4633.LUT_SIZE = 6;
	defparam lut_4633.mask = 64'h0500000000003300;

	lut_sub lut_4643 ({i_40_, i_32_, g475}, g476);
	defparam lut_4643.LUT_SIZE = 3;
	defparam lut_4643.mask = 8'h40;

	lut_sub lut_4650 ({g94, g267, g315}, g477);
	defparam lut_4650.LUT_SIZE = 3;
	defparam lut_4650.mask = 8'h10;

	lut_sub lut_4657 ({g168, g136, g79}, g478);
	defparam lut_4657.LUT_SIZE = 3;
	defparam lut_4657.mask = 8'he0;

	lut_sub lut_4668 ({g53, g24, g198, g477, g478}, g479);
	defparam lut_4668.LUT_SIZE = 5;
	defparam lut_4668.mask = 32'h0303030b;

	lut_sub lut_4683 ({g139, g225, g272}, g480);
	defparam lut_4683.LUT_SIZE = 3;
	defparam lut_4683.mask = 8'h15;

	lut_sub lut_4691 ({i_40_, g121, i_23_, g198}, g481);
	defparam lut_4691.LUT_SIZE = 4;
	defparam lut_4691.mask = 16'h0400;

	lut_sub lut_4700 ({g122, g112, g47, g94, g481}, g482);
	defparam lut_4700.LUT_SIZE = 5;
	defparam lut_4700.mask = 32'h00d50000;

	lut_sub lut_4709 ({g56, i_32_, i_31_, i_30_, i_28_, i_29_}, g483);
	defparam lut_4709.LUT_SIZE = 6;
	defparam lut_4709.mask = 64'h0000000024000000;

	lut_sub lut_4718 ({i_5_, g45, g115, g105, g483}, g484);
	defparam lut_4718.LUT_SIZE = 5;
	defparam lut_4718.mask = 32'h11150000;

	lut_sub lut_4727 ({i_32_, g47, i_0_}, g485);
	defparam lut_4727.LUT_SIZE = 3;
	defparam lut_4727.mask = 8'h40;

	lut_sub lut_4731 ({i_36_, i_37_, i_38_, i_39_, i_40_}, g486);
	defparam lut_4731.LUT_SIZE = 5;
	defparam lut_4731.mask = 32'h00000104;

	lut_sub lut_4741 ({g56, g118, g66, g485, g486}, g487);
	defparam lut_4741.LUT_SIZE = 5;
	defparam lut_4741.mask = 32'h000f111f;

	lut_sub lut_4759 ({i_40_, g220, g225, g243, g487}, g488);
	defparam lut_4759.LUT_SIZE = 5;
	defparam lut_4759.mask = 32'h88a888aa;

	lut_sub lut_4778 ({g479, g480, g482, g484, g488}, g489);
	defparam lut_4778.LUT_SIZE = 5;
	defparam lut_4778.mask = 32'h40000000;

	lut_sub lut_4787 ({g53, g474, g476, g285, g489}, o_17_);
	defparam lut_4787.LUT_SIZE = 5;
	defparam lut_4787.mask = 32'hefefffef;

	lut_sub lut_4820 ({i_37_, i_38_, i_31_, g1}, g491);
	defparam lut_4820.LUT_SIZE = 4;
	defparam lut_4820.mask = 16'h8008;

	lut_sub lut_4829 ({i_36_, g56, g353, g466, g491}, g492);
	defparam lut_4829.LUT_SIZE = 5;
	defparam lut_4829.mask = 32'h03570303;

	lut_sub lut_4844 ({g24, i_9_}, g493);
	defparam lut_4844.LUT_SIZE = 2;
	defparam lut_4844.mask = 4'b0100;

	lut_sub lut_4850 ({i_11_, i_12_, i_15_, g171, g493}, g494);
	defparam lut_4850.LUT_SIZE = 5;
	defparam lut_4850.mask = 32'h00000007;

	lut_sub lut_4859 ({i_7_, g162, i_14_, g478, g494}, g495);
	defparam lut_4859.LUT_SIZE = 5;
	defparam lut_4859.mask = 32'h04000000;

	lut_sub lut_4863 ({i_36_, i_37_, i_38_, i_39_, i_40_}, g496);
	defparam lut_4863.LUT_SIZE = 5;
	defparam lut_4863.mask = 32'hf8180000;

	lut_sub lut_4874 ({i_31_, g1, i_16_, i_9_}, g497);
	defparam lut_4874.LUT_SIZE = 4;
	defparam lut_4874.mask = 16'h7000;

	lut_sub lut_4884 ({g56, g18, g496, g497}, g498);
	defparam lut_4884.LUT_SIZE = 4;
	defparam lut_4884.mask = 16'h0001;

	lut_sub lut_4892 ({i_40_, g95, g104, g347, g462}, g499);
	defparam lut_4892.LUT_SIZE = 5;
	defparam lut_4892.mask = 32'h000f111f;

	lut_sub lut_4911 ({g5, g116, g92, g71, g187}, g500);
	defparam lut_4911.LUT_SIZE = 5;
	defparam lut_4911.mask = 32'h1111111f;

	lut_sub lut_4929 ({g116, g6, g467, g500}, g501);
	defparam lut_4929.LUT_SIZE = 4;
	defparam lut_4929.mask = 16'h0537;

	lut_sub lut_4940 ({i_37_, i_38_, i_39_, i_40_, g148}, g502);
	defparam lut_4940.LUT_SIZE = 5;
	defparam lut_4940.mask = 32'h10141505;

	lut_sub lut_4952 ({i_7_, i_33_, i_32_, g2}, g503);
	defparam lut_4952.LUT_SIZE = 4;
	defparam lut_4952.mask = 16'h0100;

	lut_sub lut_4960 ({i_37_, g76, g5, g301, g503}, g504);
	defparam lut_4960.LUT_SIZE = 5;
	defparam lut_4960.mask = 32'haaa8aaaa;

	lut_sub lut_4980 ({i_37_, i_38_, i_39_, i_40_, g95, g333}, g505);
	defparam lut_4980.LUT_SIZE = 6;
	defparam lut_4980.mask = 64'h0503050000300030;

	lut_sub lut_4994 ({i_33_, i_31_, g2}, g506);
	defparam lut_4994.LUT_SIZE = 3;
	defparam lut_4994.mask = 8'h04;

	lut_sub lut_5002 ({i_40_, g77, g8, g289, g506}, g507);
	defparam lut_5002.LUT_SIZE = 5;
	defparam lut_5002.mask = 32'h04440044;

	lut_sub lut_5015 ({g117, g502, g504, g505, g507}, g508);
	defparam lut_5015.LUT_SIZE = 5;
	defparam lut_5015.mask = 32'h08000000;

	lut_sub lut_5024 ({g495, g498, g499, g501, g508}, g509);
	defparam lut_5024.LUT_SIZE = 5;
	defparam lut_5024.mask = 32'h40000000;

	lut_sub lut_5030 ({i_37_, i_39_, g118, g96}, g510);
	defparam lut_5030.LUT_SIZE = 4;
	defparam lut_5030.mask = 16'h5111;

	lut_sub lut_5040 ({i_37_, i_38_, i_39_, i_40_, g123, g6}, g511);
	defparam lut_5040.LUT_SIZE = 6;
	defparam lut_5040.mask = 64'h0000030373735703;

	lut_sub lut_5064 ({i_7_, i_11_, i_38_, i_40_, i_10_, i_27_}, g512);
	defparam lut_5064.LUT_SIZE = 6;
	defparam lut_5064.mask = 64'h0fe000e000000000;

	lut_sub lut_5077 ({i_37_, i_38_, i_39_, i_40_}, g513);
	defparam lut_5077.LUT_SIZE = 4;
	defparam lut_5077.mask = 16'he4b1;

	lut_sub lut_5092 ({i_36_, g102, g408, g512, g513}, g514);
	defparam lut_5092.LUT_SIZE = 5;
	defparam lut_5092.mask = 32'h0a0a0033;

	lut_sub lut_5105 ({i_38_, i_40_, g51, i_15_, g385}, g515);
	defparam lut_5105.LUT_SIZE = 5;
	defparam lut_5105.mask = 32'h00000100;

	lut_sub lut_5111 ({g162, i_31_, g155}, g516);
	defparam lut_5111.LUT_SIZE = 3;
	defparam lut_5111.mask = 8'h40;

	lut_sub lut_5120 ({g135, g390, g470, g515, g516}, g517);
	defparam lut_5120.LUT_SIZE = 5;
	defparam lut_5120.mask = 32'heaeaea00;

	lut_sub lut_5143 ({g121, g510, g511, g514, g517}, g518);
	defparam lut_5143.LUT_SIZE = 5;
	defparam lut_5143.mask = 32'h44004000;

	lut_sub lut_5154 ({g73, g492, g397, g509, g518}, g519);
	defparam lut_5154.LUT_SIZE = 5;
	defparam lut_5154.mask = 32'h01010100;

	lut_sub lut_5162 ({i_7_, g67, g461}, g520);
	defparam lut_5162.LUT_SIZE = 3;
	defparam lut_5162.mask = 8'h10;

	lut_sub lut_5171 ({i_38_, g101, g197, g136, g66, g520}, g521);
	defparam lut_5171.LUT_SIZE = 6;
	defparam lut_5171.mask = 64'h0005000011111111;

	lut_sub lut_5187 ({g45, g73, g408}, g522);
	defparam lut_5187.LUT_SIZE = 3;
	defparam lut_5187.mask = 8'h01;

	lut_sub lut_5192 ({i_38_, i_39_, i_40_, g121}, g523);
	defparam lut_5192.LUT_SIZE = 4;
	defparam lut_5192.mask = 16'h0140;

	lut_sub lut_5201 ({i_40_, g21, g7, g148, g8}, g524);
	defparam lut_5201.LUT_SIZE = 5;
	defparam lut_5201.mask = 32'h00330505;

	lut_sub lut_5216 ({i_37_, g6, g522, g523, g524}, g525);
	defparam lut_5216.LUT_SIZE = 5;
	defparam lut_5216.mask = 32'ha080a0a0;

	lut_sub lut_5230 ({g48, i_6_, g712, g521, g525}, g526);
	defparam lut_5230.LUT_SIZE = 5;
	defparam lut_5230.mask = 32'h44444404;

	lut_sub lut_5245 ({g122, g2, g21, g24, g112}, g527);
	defparam lut_5245.LUT_SIZE = 5;
	defparam lut_5245.mask = 32'h004c0000;

	lut_sub lut_5255 ({g65, i_9_, g260, g136, g527}, g528);
	defparam lut_5255.LUT_SIZE = 5;
	defparam lut_5255.mask = 32'h00550057;

	lut_sub lut_5267 ({i_36_, i_37_, i_38_, i_39_, i_40_}, g529);
	defparam lut_5267.LUT_SIZE = 5;
	defparam lut_5267.mask = 32'h02020004;

	lut_sub lut_5273 ({i_37_, i_35_, i_13_}, g530);
	defparam lut_5273.LUT_SIZE = 3;
	defparam lut_5273.mask = 8'h20;

	lut_sub lut_5279 ({i_36_, i_38_, i_39_, i_40_, g136, g530}, g531);
	defparam lut_5279.LUT_SIZE = 6;
	defparam lut_5279.mask = 64'h0a22000000000000;

	lut_sub lut_5292 ({g168, g151, g187, g189, g165, g531}, g532);
	defparam lut_5292.LUT_SIZE = 6;
	defparam lut_5292.mask = 64'h8080800000000000;

	lut_sub lut_5303 ({g65, g22, g454, g529, g532}, g533);
	defparam lut_5303.LUT_SIZE = 5;
	defparam lut_5303.mask = 32'h000003ab;

	lut_sub lut_5317 ({g122, g2, g21, g113}, g534);
	defparam lut_5317.LUT_SIZE = 4;
	defparam lut_5317.mask = 16'h0700;

	lut_sub lut_5327 ({g171, g493, i_14_, g385, g534}, g535);
	defparam lut_5327.LUT_SIZE = 5;
	defparam lut_5327.mask = 32'h00505454;

	lut_sub lut_5342 ({i_12_, g196, g528, g533, g535}, g536);
	defparam lut_5342.LUT_SIZE = 5;
	defparam lut_5342.mask = 32'h80008800;

	lut_sub lut_5352 ({g28, g10, g255, g315}, g537);
	defparam lut_5352.LUT_SIZE = 4;
	defparam lut_5352.mask = 16'h44f4;

	lut_sub lut_5362 ({i_36_, i_37_, i_38_, i_39_, i_40_}, g538);
	defparam lut_5362.LUT_SIZE = 5;
	defparam lut_5362.mask = 32'h78400000;

	lut_sub lut_5374 ({g162, i_35_, g46, g442, g538}, g539);
	defparam lut_5374.LUT_SIZE = 5;
	defparam lut_5374.mask = 32'h5f330000;

	lut_sub lut_5387 ({i_37_, i_38_, i_39_, i_40_}, g540);
	defparam lut_5387.LUT_SIZE = 4;
	defparam lut_5387.mask = 16'h0140;

	lut_sub lut_5394 ({i_13_, g28, i_9_, g129}, g541);
	defparam lut_5394.LUT_SIZE = 4;
	defparam lut_5394.mask = 16'h0357;

	lut_sub lut_5408 ({i_36_, g162, g70, g540, g541}, g542);
	defparam lut_5408.LUT_SIZE = 5;
	defparam lut_5408.mask = 32'h37050505;

	lut_sub lut_5426 ({i_15_, g48, g537, g539, g542}, g543);
	defparam lut_5426.LUT_SIZE = 5;
	defparam lut_5426.mask = 32'h007f0000;

	lut_sub lut_5438 ({i_37_, i_40_, g162, i_35_, g281}, g544);
	defparam lut_5438.LUT_SIZE = 5;
	defparam lut_5438.mask = 32'h50500010;

	lut_sub lut_5449 ({i_36_, i_37_, i_38_, g101, g106, g66}, g545);
	defparam lut_5449.LUT_SIZE = 6;
	defparam lut_5449.mask = 64'h3055005500550055;

	lut_sub lut_5475 ({g65, g71, g79, g454, g545}, g546);
	defparam lut_5475.LUT_SIZE = 5;
	defparam lut_5475.mask = 32'h11111113;

	lut_sub lut_5491 ({i_5_, g48, g537, g544, g546}, g547);
	defparam lut_5491.LUT_SIZE = 5;
	defparam lut_5491.mask = 32'haaaaaa80;

	lut_sub lut_5510 ({i_7_, g122, i_5_, g2, g195}, g548);
	defparam lut_5510.LUT_SIZE = 5;
	defparam lut_5510.mask = 32'h01000000;

	lut_sub lut_5517 ({i_36_, g162, i_5_, g61, g48}, g549);
	defparam lut_5517.LUT_SIZE = 5;
	defparam lut_5517.mask = 32'h01000000;

	lut_sub lut_5521 ({i_37_, i_38_, i_39_, i_40_, i_31_}, g550);
	defparam lut_5521.LUT_SIZE = 5;
	defparam lut_5521.mask = 32'h000bf000;

	lut_sub lut_5534 ({i_31_, i_5_, g293, g549, g550}, g551);
	defparam lut_5534.LUT_SIZE = 5;
	defparam lut_5534.mask = 32'hccc4c4c4;

	lut_sub lut_5554 ({i_7_, g22, g181, g548, g551}, g552);
	defparam lut_5554.LUT_SIZE = 5;
	defparam lut_5554.mask = 32'h44044444;

	lut_sub lut_5567 ({i_7_, i_11_, g103, g528, g552}, g553);
	defparam lut_5567.LUT_SIZE = 5;
	defparam lut_5567.mask = 32'h44505555;

	lut_sub lut_5586 ({i_7_, g536, g543, g547, g553}, g554);
	defparam lut_5586.LUT_SIZE = 5;
	defparam lut_5586.mask = 32'h00101010;

	lut_sub lut_5593 ({i_36_, i_38_, i_39_, i_40_, g88, i_6_}, g555);
	defparam lut_5593.LUT_SIZE = 6;
	defparam lut_5593.mask = 64'h000000000a000002;

	lut_sub lut_5601 ({i_36_, i_37_, i_0_, g187, g555}, g556);
	defparam lut_5601.LUT_SIZE = 5;
	defparam lut_5601.mask = 32'haaaaaa8a;

	lut_sub lut_5621 ({i_36_, i_37_, g5, g79}, g557);
	defparam lut_5621.LUT_SIZE = 4;
	defparam lut_5621.mask = 16'h1113;

	lut_sub lut_5631 ({i_36_, g100, i_35_, g73}, g558);
	defparam lut_5631.LUT_SIZE = 4;
	defparam lut_5631.mask = 16'h0004;

	lut_sub lut_5637 ({i_37_, i_34_, g51, g79, i_6_}, g559);
	defparam lut_5637.LUT_SIZE = 5;
	defparam lut_5637.mask = 32'h00000002;

	lut_sub lut_5644 ({i_34_, i_32_, g51, g558, g559}, g560);
	defparam lut_5644.LUT_SIZE = 5;
	defparam lut_5644.mask = 32'haa08aa80;

	lut_sub lut_5659 ({i_34_, g113, g78}, g561);
	defparam lut_5659.LUT_SIZE = 3;
	defparam lut_5659.mask = 8'h10;

	lut_sub lut_5667 ({i_37_, i_38_, g101, g160, g94, g318}, g562);
	defparam lut_5667.LUT_SIZE = 6;
	defparam lut_5667.mask = 64'h22aaaaaaaaaaa0a0;

	lut_sub lut_5698 ({i_36_, i_37_, i_34_, g77, g562}, g563);
	defparam lut_5698.LUT_SIZE = 5;
	defparam lut_5698.mask = 32'h55555545;

	lut_sub lut_5719 ({i_33_, g1, i_0_, g561, g563}, g564);
	defparam lut_5719.LUT_SIZE = 5;
	defparam lut_5719.mask = 32'h00004fff;

	lut_sub lut_5739 ({i_7_, g556, g557, g560, g564}, g565);
	defparam lut_5739.LUT_SIZE = 5;
	defparam lut_5739.mask = 32'h10115555;

	lut_sub lut_5753 ({i_37_, i_40_, i_31_, i_9_}, g566);
	defparam lut_5753.LUT_SIZE = 4;
	defparam lut_5753.mask = 16'h4000;

	lut_sub lut_5758 ({i_11_, i_5_, i_12_, i_15_, i_14_, g566}, g567);
	defparam lut_5758.LUT_SIZE = 6;
	defparam lut_5758.mask = 64'hffff0000fffa0002;

	lut_sub lut_5792 ({i_37_, i_38_, i_39_, i_40_}, g568);
	defparam lut_5792.LUT_SIZE = 4;
	defparam lut_5792.mask = 16'hc1c0;

	lut_sub lut_5801 ({i_16_, i_17_, i_9_, g568}, g569);
	defparam lut_5801.LUT_SIZE = 4;
	defparam lut_5801.mask = 16'h0115;

	lut_sub lut_5810 ({i_33_, i_5_, g2, g569}, g570);
	defparam lut_5810.LUT_SIZE = 4;
	defparam lut_5810.mask = 16'h0002;

	lut_sub lut_5815 ({i_16_, i_9_, g18}, g571);
	defparam lut_5815.LUT_SIZE = 3;
	defparam lut_5815.mask = 8'h15;

	lut_sub lut_5823 ({i_37_, i_38_, i_39_, i_40_, g506, g571}, g572);
	defparam lut_5823.LUT_SIZE = 6;
	defparam lut_5823.mask = 64'h3111100000013000;

	lut_sub lut_5839 ({i_36_, g56, g567, g570, g572}, g573);
	defparam lut_5839.LUT_SIZE = 5;
	defparam lut_5839.mask = 32'h88088888;

	lut_sub lut_5852 ({i_39_, i_40_, i_35_, g65, g116, g454}, g574);
	defparam lut_5852.LUT_SIZE = 6;
	defparam lut_5852.mask = 64'h0000010000010000;

	lut_sub lut_5861 ({i_7_, g573, g503, g547, g574}, o_22_);
	defparam lut_5861.LUT_SIZE = 5;
	defparam lut_5861.mask = 32'hffdfdfdf;

	lut_sub lut_5896 ({i_36_, g100, g106, g73}, g576);
	defparam lut_5896.LUT_SIZE = 4;
	defparam lut_5896.mask = 16'h0001;

	lut_sub lut_5903 ({i_38_, i_39_, g122, g136, g385}, g577);
	defparam lut_5903.LUT_SIZE = 5;
	defparam lut_5903.mask = 32'h00000020;

	lut_sub lut_5910 ({i_37_, g122, g5, i_0_, g69}, g578);
	defparam lut_5910.LUT_SIZE = 5;
	defparam lut_5910.mask = 32'h00000100;

	lut_sub lut_5917 ({i_38_, g73, g219, g704}, g579);
	defparam lut_5917.LUT_SIZE = 4;
	defparam lut_5917.mask = 16'h4555;

	lut_sub lut_5930 ({i_37_, i_38_, g47, g87, g130}, g580);
	defparam lut_5930.LUT_SIZE = 5;
	defparam lut_5930.mask = 32'h11005100;

	lut_sub lut_5941 ({i_31_, g122, i_5_, g2, g580}, g581);
	defparam lut_5941.LUT_SIZE = 5;
	defparam lut_5941.mask = 32'ha8aa88aa;

	lut_sub lut_5959 ({i_34_, g30, i_15_, g106}, g582);
	defparam lut_5959.LUT_SIZE = 4;
	defparam lut_5959.mask = 16'h4000;

	lut_sub lut_5967 ({i_40_, g27, g105, g106, g582}, g583);
	defparam lut_5967.LUT_SIZE = 5;
	defparam lut_5967.mask = 32'ha8a8a888;

	lut_sub lut_5984 ({i_38_, g101, g134, g152}, g584);
	defparam lut_5984.LUT_SIZE = 4;
	defparam lut_5984.mask = 16'h5445;

	lut_sub lut_5995 ({i_38_, i_39_, g122, i_15_, g2}, g585);
	defparam lut_5995.LUT_SIZE = 5;
	defparam lut_5995.mask = 32'h00400050;

	lut_sub lut_6004 ({i_37_, i_38_, g134, g92, g585}, g586);
	defparam lut_6004.LUT_SIZE = 5;
	defparam lut_6004.mask = 32'h57035500;

	lut_sub lut_6023 ({g184, g581, g583, g584, g586}, g587);
	defparam lut_6023.LUT_SIZE = 5;
	defparam lut_6023.mask = 32'h00000002;

	lut_sub lut_6029 ({g22, i_16_, i_9_, g255}, g588);
	defparam lut_6029.LUT_SIZE = 4;
	defparam lut_6029.mask = 16'h7f55;

	lut_sub lut_6047 ({i_37_, g51, g122, i_15_, g5, g87}, g589);
	defparam lut_6047.LUT_SIZE = 6;
	defparam lut_6047.mask = 64'h0000f00011001100;

	lut_sub lut_6061 ({i_34_, i_5_, i_0_, g106, g214, g589}, g590);
	defparam lut_6061.LUT_SIZE = 6;
	defparam lut_6061.mask = 64'haa88a080aa88aa88;

	lut_sub lut_6086 ({i_37_, i_38_, i_39_, i_40_, g92}, g591);
	defparam lut_6086.LUT_SIZE = 5;
	defparam lut_6086.mask = 32'hf03c0c55;

	lut_sub lut_6103 ({i_36_, i_37_, i_38_, i_39_, i_40_, i_35_}, g592);
	defparam lut_6103.LUT_SIZE = 6;
	defparam lut_6103.mask = 64'h0000fd5177a82a8a;

	lut_sub lut_6132 ({i_38_, i_39_, i_40_, g22, i_16_, i_9_}, g593);
	defparam lut_6132.LUT_SIZE = 6;
	defparam lut_6132.mask = 64'h888f8f8f88888888;

	lut_sub lut_6163 ({i_36_, i_39_, g102, g30, g593}, g594);
	defparam lut_6163.LUT_SIZE = 5;
	defparam lut_6163.mask = 32'h04050404;

	lut_sub lut_6175 ({i_35_, g65, g591, g592, g594}, g595);
	defparam lut_6175.LUT_SIZE = 5;
	defparam lut_6175.mask = 32'haa88aa80;

	lut_sub lut_6192 ({i_38_, i_9_, g585, g693, g595}, g596);
	defparam lut_6192.LUT_SIZE = 5;
	defparam lut_6192.mask = 32'h50551011;

	lut_sub lut_6210 ({g576, g577, g578, g579, g587, g596}, g597);
	defparam lut_6210.LUT_SIZE = 6;
	defparam lut_6210.mask = 64'h0100000000000000;

	lut_sub lut_6218 ({g112, g18, g121, g365}, g598);
	defparam lut_6218.LUT_SIZE = 4;
	defparam lut_6218.mask = 16'h0001;

	lut_sub lut_6224 ({g23, g84, i_21_, i_23_}, g599);
	defparam lut_6224.LUT_SIZE = 4;
	defparam lut_6224.mask = 16'h0008;

	lut_sub lut_6231 ({g43, g375, g399}, g600);
	defparam lut_6231.LUT_SIZE = 3;
	defparam lut_6231.mask = 8'h01;

	lut_sub lut_6238 ({g143, g43, i_23_, g246}, g601);
	defparam lut_6238.LUT_SIZE = 4;
	defparam lut_6238.mask = 16'h0004;

	lut_sub lut_6242 ({i_36_, i_37_, i_38_, i_39_, i_40_}, g602);
	defparam lut_6242.LUT_SIZE = 5;
	defparam lut_6242.mask = 32'h80400000;

	lut_sub lut_6251 ({i_11_, g1, i_12_, g28, g42, g602}, g603);
	defparam lut_6251.LUT_SIZE = 6;
	defparam lut_6251.mask = 64'h0013000013130000;

	lut_sub lut_6267 ({i_11_, g1, i_12_, g246, g355, g442}, g604);
	defparam lut_6267.LUT_SIZE = 6;
	defparam lut_6267.mask = 64'h0013000013130000;

	lut_sub lut_6285 ({g2, g21, g3, g23, g24, g113}, g605);
	defparam lut_6285.LUT_SIZE = 6;
	defparam lut_6285.mask = 64'h0000000000010003;

	lut_sub lut_6297 ({g599, g600, g601, g603, g604, g605}, g606);
	defparam lut_6297.LUT_SIZE = 6;
	defparam lut_6297.mask = 64'h8000000000000000;

	lut_sub lut_6307 ({g124, g367, g41, g20, g598, g606}, g607);
	defparam lut_6307.LUT_SIZE = 6;
	defparam lut_6307.mask = 64'h0004000400040000;

	lut_sub lut_6318 ({g53, g107, g108, g119, g338}, g608);
	defparam lut_6318.LUT_SIZE = 5;
	defparam lut_6318.mask = 32'h00000777;

	lut_sub lut_6334 ({g197, g136, g69, g330}, g609);
	defparam lut_6334.LUT_SIZE = 4;
	defparam lut_6334.mask = 16'h0001;

	lut_sub lut_6341 ({i_40_, g121, g6, g346}, g610);
	defparam lut_6341.LUT_SIZE = 4;
	defparam lut_6341.mask = 16'hfeff;

	lut_sub lut_6363 ({g331, g609, g50, g610}, g611);
	defparam lut_6363.LUT_SIZE = 4;
	defparam lut_6363.mask = 16'h4000;

	lut_sub lut_6371 ({g14, g134, g330, g611}, g612);
	defparam lut_6371.LUT_SIZE = 4;
	defparam lut_6371.mask = 16'h5554;

	lut_sub lut_6386 ({g607, g305, g608, g82, g612}, g613);
	defparam lut_6386.LUT_SIZE = 5;
	defparam lut_6386.mask = 32'h00001000;

	lut_sub lut_6394 ({g14, g197, g136, g330}, g614);
	defparam lut_6394.LUT_SIZE = 4;
	defparam lut_6394.mask = 16'h0001;

	lut_sub lut_6402 ({g74, g331, g609, g614}, g615);
	defparam lut_6402.LUT_SIZE = 4;
	defparam lut_6402.mask = 16'h8000;

	lut_sub lut_6410 ({g607, g305, g608, g615}, g616);
	defparam lut_6410.LUT_SIZE = 4;
	defparam lut_6410.mask = 16'h0040;

	lut_sub lut_6420 ({g66, g68, g81, g187, g305, g50}, g617);
	defparam lut_6420.LUT_SIZE = 6;
	defparam lut_6420.mask = 64'h8800880088008000;

	lut_sub lut_6434 ({g23, i_24_, g131, g126, g219}, g618);
	defparam lut_6434.LUT_SIZE = 5;
	defparam lut_6434.mask = 32'h00000537;

	lut_sub lut_6447 ({i_22_, i_21_, g9, g608, g618}, g619);
	defparam lut_6447.LUT_SIZE = 5;
	defparam lut_6447.mask = 32'hc0c080c0;

	lut_sub lut_6457 ({i_38_, i_39_, i_40_}, g620);
	defparam lut_6457.LUT_SIZE = 3;
	defparam lut_6457.mask = 8'h83;

	lut_sub lut_6467 ({i_22_, g151, g266, g432, g620}, g621);
	defparam lut_6467.LUT_SIZE = 5;
	defparam lut_6467.mask = 32'h337f000f;

	lut_sub lut_6488 ({g151, i_21_, g187, g621}, g622);
	defparam lut_6488.LUT_SIZE = 4;
	defparam lut_6488.mask = 16'haa8a;

	lut_sub lut_6499 ({i_24_, g84, i_21_, i_23_}, g623);
	defparam lut_6499.LUT_SIZE = 4;
	defparam lut_6499.mask = 16'h0008;

	lut_sub lut_6507 ({g74, g325, g600, g623}, g624);
	defparam lut_6507.LUT_SIZE = 4;
	defparam lut_6507.mask = 16'hc800;

	lut_sub lut_6517 ({g65, g23, i_24_, g622, g624}, o_30_);
	defparam lut_6517.LUT_SIZE = 5;
	defparam lut_6517.mask = 32'haaaaaaae;

	lut_sub lut_6539 ({i_22_, g84, i_21_, g325}, g626);
	defparam lut_6539.LUT_SIZE = 4;
	defparam lut_6539.mask = 16'h0004;

	lut_sub lut_6547 ({g61, g125, g390, g626}, g627);
	defparam lut_6547.LUT_SIZE = 4;
	defparam lut_6547.mask = 16'haaa8;

	lut_sub lut_6561 ({g29, i_23_, g17, g615, g627}, o_31_);
	defparam lut_6561.LUT_SIZE = 5;
	defparam lut_6561.mask = 32'hefcfffff;

	lut_sub lut_6594 ({i_31_, i_5_, i_15_, g401}, g629);
	defparam lut_6594.LUT_SIZE = 4;
	defparam lut_6594.mask = 16'h4000;

	lut_sub lut_6601 ({g100, i_35_, g73, g172}, g630);
	defparam lut_6601.LUT_SIZE = 4;
	defparam lut_6601.mask = 16'h0001;

	lut_sub lut_6605 ({i_36_, i_37_, i_38_, i_39_, i_40_, i_35_}, g631);
	defparam lut_6605.LUT_SIZE = 6;
	defparam lut_6605.mask = 64'h00000000000c8100;

	lut_sub lut_6617 ({g101, g151, g204, g220, g436}, g632);
	defparam lut_6617.LUT_SIZE = 5;
	defparam lut_6617.mask = 32'h0c0c0c5d;

	lut_sub lut_6636 ({g65, g629, g630, g631, g632}, g633);
	defparam lut_6636.LUT_SIZE = 5;
	defparam lut_6636.mask = 32'h00007fff;

	lut_sub lut_6656 ({i_37_, i_34_, i_35_, g3, g260}, g634);
	defparam lut_6656.LUT_SIZE = 5;
	defparam lut_6656.mask = 32'h10000000;

	lut_sub lut_6663 ({g56, i_32_, i_31_, g24, g46}, g635);
	defparam lut_6663.LUT_SIZE = 5;
	defparam lut_6663.mask = 32'h00004000;

	lut_sub lut_6672 ({g24, g138, g275, g634, g635}, g636);
	defparam lut_6672.LUT_SIZE = 5;
	defparam lut_6672.mask = 32'h88808888;

	lut_sub lut_6683 ({i_31_, i_5_, i_15_, g180}, g637);
	defparam lut_6683.LUT_SIZE = 4;
	defparam lut_6683.mask = 16'h4000;

	lut_sub lut_6688 ({i_5_, i_9_, g637}, g638);
	defparam lut_6688.LUT_SIZE = 3;
	defparam lut_6688.mask = 8'h8a;

	lut_sub lut_6697 ({i_40_, g56, g46, g275}, g639);
	defparam lut_6697.LUT_SIZE = 4;
	defparam lut_6697.mask = 16'h0357;

	lut_sub lut_6709 ({g24, g138, i_14_}, g640);
	defparam lut_6709.LUT_SIZE = 3;
	defparam lut_6709.mask = 8'h20;

	lut_sub lut_6718 ({g53, g470, g637, g639, g640}, g641);
	defparam lut_6718.LUT_SIZE = 5;
	defparam lut_6718.mask = 32'he0e0e000;

	lut_sub lut_6734 ({i_12_, i_15_, g634, g636, g638, g641}, g642);
	defparam lut_6734.LUT_SIZE = 6;
	defparam lut_6734.mask = 64'hc8ccc8c888cc8888;

	lut_sub lut_6762 ({g100, i_40_, g122, i_6_}, g643);
	defparam lut_6762.LUT_SIZE = 4;
	defparam lut_6762.mask = 16'h0400;

	lut_sub lut_6770 ({g116, g160, g94, g643}, g644);
	defparam lut_6770.LUT_SIZE = 4;
	defparam lut_6770.mask = 16'h0544;

	lut_sub lut_6777 ({i_37_, i_38_, i_39_, i_40_}, g645);
	defparam lut_6777.LUT_SIZE = 4;
	defparam lut_6777.mask = 16'h71d0;

	lut_sub lut_6790 ({i_37_, g122, i_13_, g5, g187}, g646);
	defparam lut_6790.LUT_SIZE = 5;
	defparam lut_6790.mask = 32'h10000000;

	lut_sub lut_6799 ({g2, g3, g189, g645, g646}, g647);
	defparam lut_6799.LUT_SIZE = 5;
	defparam lut_6799.mask = 32'haaa0aa80;

	lut_sub lut_6817 ({i_5_, g22, i_13_, g132, g644, g647}, g648);
	defparam lut_6817.LUT_SIZE = 6;
	defparam lut_6817.mask = 64'hcccc4044cccccccc;

	lut_sub lut_6849 ({i_32_, i_31_, i_5_, g171, g201}, g649);
	defparam lut_6849.LUT_SIZE = 5;
	defparam lut_6849.mask = 32'h20000000;

	lut_sub lut_6855 ({g100, i_39_, i_40_, i_35_, g151}, g650);
	defparam lut_6855.LUT_SIZE = 5;
	defparam lut_6855.mask = 32'h00053005;

	lut_sub lut_6867 ({i_36_, i_32_, g10, g67, g187}, g651);
	defparam lut_6867.LUT_SIZE = 5;
	defparam lut_6867.mask = 32'h00001000;

	lut_sub lut_6875 ({g423, g465, g650, g651}, g652);
	defparam lut_6875.LUT_SIZE = 4;
	defparam lut_6875.mask = 16'h0537;

	lut_sub lut_6887 ({i_40_, g98, g214}, g653);
	defparam lut_6887.LUT_SIZE = 3;
	defparam lut_6887.mask = 8'h01;

	lut_sub lut_6895 ({i_40_, g122, g21, g47, g94}, g654);
	defparam lut_6895.LUT_SIZE = 5;
	defparam lut_6895.mask = 32'h02000000;

	lut_sub lut_6903 ({i_33_, i_32_, g86, g67, g461, g654}, g655);
	defparam lut_6903.LUT_SIZE = 6;
	defparam lut_6903.mask = 64'haaa80000aaa8aaaa;

	lut_sub lut_6932 ({g22, g218, g653, g655}, g656);
	defparam lut_6932.LUT_SIZE = 4;
	defparam lut_6932.mask = 16'h0405;

	lut_sub lut_6943 ({g450, g458, g649, g652, g656}, g657);
	defparam lut_6943.LUT_SIZE = 5;
	defparam lut_6943.mask = 32'h00440040;

	lut_sub lut_6953 ({g135, g84, g152, g172}, g658);
	defparam lut_6953.LUT_SIZE = 4;
	defparam lut_6953.mask = 16'h4555;

	lut_sub lut_6965 ({i_11_, i_5_, i_9_, g636, g658}, g659);
	defparam lut_6965.LUT_SIZE = 5;
	defparam lut_6965.mask = 32'ha2aaaaaa;

	lut_sub lut_6989 ({g633, g642, g648, g435, g657, g659}, g660);
	defparam lut_6989.LUT_SIZE = 6;
	defparam lut_6989.mask = 64'h0001000000000000;

	lut_sub lut_6994 ({i_36_, i_37_, i_38_, i_39_, i_40_, g462}, g661);
	defparam lut_6994.LUT_SIZE = 6;
	defparam lut_6994.mask = 64'h0000000000050010;

	lut_sub lut_7002 ({i_36_, i_5_, i_15_, g201, g661}, g662);
	defparam lut_7002.LUT_SIZE = 5;
	defparam lut_7002.mask = 32'haa02aaaa;

	lut_sub lut_7021 ({i_36_, g162, i_35_, g112, g260}, g663);
	defparam lut_7021.LUT_SIZE = 5;
	defparam lut_7021.mask = 32'h75003000;

	lut_sub lut_7036 ({g100, g101, g280, g255, g663}, g664);
	defparam lut_7036.LUT_SIZE = 5;
	defparam lut_7036.mask = 32'ha0a020a0;

	lut_sub lut_7049 ({i_36_, i_40_, g162, g346, g664}, g665);
	defparam lut_7049.LUT_SIZE = 5;
	defparam lut_7049.mask = 32'h55555545;

	lut_sub lut_7070 ({i_36_, i_40_, g162, g21, g465}, g666);
	defparam lut_7070.LUT_SIZE = 5;
	defparam lut_7070.mask = 32'h00001000;

	lut_sub lut_7077 ({i_36_, g100, g101, g49}, g667);
	defparam lut_7077.LUT_SIZE = 4;
	defparam lut_7077.mask = 16'h0800;

	lut_sub lut_7086 ({g280, g67, g461, g666, g667}, g668);
	defparam lut_7086.LUT_SIZE = 5;
	defparam lut_7086.mask = 32'h0037003f;

	lut_sub lut_7102 ({i_32_, i_5_, i_0_, g665, g668}, g669);
	defparam lut_7102.LUT_SIZE = 5;
	defparam lut_7102.mask = 32'h55d50000;

	lut_sub lut_7116 ({i_37_, i_35_, g53, i_9_, g260}, g670);
	defparam lut_7116.LUT_SIZE = 5;
	defparam lut_7116.mask = 32'h01000000;

	lut_sub lut_7123 ({i_11_, i_38_, g73, g219, g653}, g671);
	defparam lut_7123.LUT_SIZE = 5;
	defparam lut_7123.mask = 32'h00035557;

	lut_sub lut_7141 ({g2, g21, g3, g201}, g672);
	defparam lut_7141.LUT_SIZE = 4;
	defparam lut_7141.mask = 16'h0002;

	lut_sub lut_7149 ({g53, g136, g79, g672}, g673);
	defparam lut_7149.LUT_SIZE = 4;
	defparam lut_7149.mask = 16'haaa8;

	lut_sub lut_7161 ({i_39_, g53, i_15_, i_9_, g136}, g674);
	defparam lut_7161.LUT_SIZE = 5;
	defparam lut_7161.mask = 32'h00000010;

	lut_sub lut_7170 ({g171, g493, g673, g203, g674}, g675);
	defparam lut_7170.LUT_SIZE = 5;
	defparam lut_7170.mask = 32'h88080808;

	lut_sub lut_7183 ({g385, g457, g670, g671, g675}, g676);
	defparam lut_7183.LUT_SIZE = 5;
	defparam lut_7183.mask = 32'h00400044;

	lut_sub lut_7191 ({i_37_, i_38_, i_39_, i_40_, g160, g94}, g677);
	defparam lut_7191.LUT_SIZE = 6;
	defparam lut_7191.mask = 64'h000000030300000a;

	lut_sub lut_7202 ({i_36_, i_37_, i_40_, g162, g104}, g678);
	defparam lut_7202.LUT_SIZE = 5;
	defparam lut_7202.mask = 32'h40000000;

	lut_sub lut_7207 ({i_36_, i_37_, i_38_, i_39_, i_40_, g56}, g679);
	defparam lut_7207.LUT_SIZE = 6;
	defparam lut_7207.mask = 64'h1501510000000000;

	lut_sub lut_7219 ({i_32_, i_31_, i_15_, g678, g679}, g680);
	defparam lut_7219.LUT_SIZE = 5;
	defparam lut_7219.mask = 32'h70000000;

	lut_sub lut_7229 ({i_31_, g22, g27, g73, g401}, g681);
	defparam lut_7229.LUT_SIZE = 5;
	defparam lut_7229.mask = 32'h00570000;

	lut_sub lut_7240 ({i_37_, g260, g78, g187}, g682);
	defparam lut_7240.LUT_SIZE = 4;
	defparam lut_7240.mask = 16'h0311;

	lut_sub lut_7250 ({g51, i_5_, g195, g682}, g683);
	defparam lut_7250.LUT_SIZE = 4;
	defparam lut_7250.mask = 16'haaa8;

	lut_sub lut_7260 ({i_36_, i_37_, i_38_, i_39_, i_34_, i_35_}, g684);
	defparam lut_7260.LUT_SIZE = 6;
	defparam lut_7260.mask = 64'hc88c088800000000;

	lut_sub lut_7275 ({i_37_, g51, g131, g684}, g685);
	defparam lut_7275.LUT_SIZE = 4;
	defparam lut_7275.mask = 16'haaa8;

	lut_sub lut_7289 ({g122, i_5_, g139, g121, g685}, g686);
	defparam lut_7289.LUT_SIZE = 5;
	defparam lut_7289.mask = 32'h00ab0000;

	lut_sub lut_7301 ({g65, g681, g683, g686}, g687);
	defparam lut_7301.LUT_SIZE = 4;
	defparam lut_7301.mask = 16'haa20;

	lut_sub lut_7313 ({g122, i_6_, g677, g680, g687}, g688);
	defparam lut_7313.LUT_SIZE = 5;
	defparam lut_7313.mask = 32'h44404444;

	lut_sub lut_7328 ({g102, g662, g669, g676, g688}, g689);
	defparam lut_7328.LUT_SIZE = 5;
	defparam lut_7328.mask = 32'h10100010;

	lut_sub lut_7334 ({i_17_, i_16_, i_15_, i_12_, i_11_, i_9_}, g690);
	defparam lut_7334.LUT_SIZE = 6;
	defparam lut_7334.mask = 64'h000000140014003c;

	lut_sub lut_7346 ({g690, i_5_}, g691);
	defparam lut_7346.LUT_SIZE = 2;
	defparam lut_7346.mask = 4'b0010;

	lut_sub lut_7354 ({i_19_, g23, i_18_, g18, g34, g84}, g692);
	defparam lut_7354.LUT_SIZE = 6;
	defparam lut_7354.mask = 64'h0101550101000100;

	lut_sub lut_7368 ({g694, g695}, g693);
	defparam lut_7368.LUT_SIZE = 2;
	defparam lut_7368.mask = 4'b1000;

	lut_sub lut_7373 ({i_32_, g696}, g694);
	defparam lut_7373.LUT_SIZE = 2;
	defparam lut_7373.mask = 4'b0100;

	lut_sub lut_7378 ({i_32_, g699}, g695);
	defparam lut_7378.LUT_SIZE = 2;
	defparam lut_7378.mask = 4'b0001;

	lut_sub lut_7384 ({g697, g698}, g696);
	defparam lut_7384.LUT_SIZE = 2;
	defparam lut_7384.mask = 4'b1000;

	lut_sub lut_7389 ({i_37_, g702}, g697);
	defparam lut_7389.LUT_SIZE = 2;
	defparam lut_7389.mask = 4'b0100;

	lut_sub lut_7394 ({i_37_, g703}, g698);
	defparam lut_7394.LUT_SIZE = 2;
	defparam lut_7394.mask = 4'b0001;

	lut_sub lut_7400 ({g700, g701}, g699);
	defparam lut_7400.LUT_SIZE = 2;
	defparam lut_7400.mask = 4'b1000;

	lut_sub lut_7405 ({i_37_, g590}, g700);
	defparam lut_7405.LUT_SIZE = 2;
	defparam lut_7405.mask = 4'b0100;

	lut_sub lut_7410 ({i_37_, g590}, g701);
	defparam lut_7410.LUT_SIZE = 2;
	defparam lut_7410.mask = 4'b0001;

	lut_sub lut_7416 ({g588, g590}, g702);
	defparam lut_7416.LUT_SIZE = 2;
	defparam lut_7416.mask = 4'b0001;

	lut_sub lut_7422 ({i_5_, g162, i_0_, g590}, g703);
	defparam lut_7422.LUT_SIZE = 4;
	defparam lut_7422.mask = 16'h5515;

	lut_sub lut_7434 ({g705, g706}, g704);
	defparam lut_7434.LUT_SIZE = 2;
	defparam lut_7434.mask = 4'b1000;

	lut_sub lut_7439 ({i_37_, g707}, g705);
	defparam lut_7439.LUT_SIZE = 2;
	defparam lut_7439.mask = 4'b0100;

	lut_sub lut_7444 ({i_37_, g709}, g706);
	defparam lut_7444.LUT_SIZE = 2;
	defparam lut_7444.mask = 4'b0001;

	lut_sub lut_7449 ({i_0_, g708}, g707);
	defparam lut_7449.LUT_SIZE = 2;
	defparam lut_7449.mask = 4'b1000;

	lut_sub lut_7454 ({i_0_, g711}, g708);
	defparam lut_7454.LUT_SIZE = 2;
	defparam lut_7454.mask = 4'b0100;

	lut_sub lut_7459 ({i_0_, g710}, g709);
	defparam lut_7459.LUT_SIZE = 2;
	defparam lut_7459.mask = 4'b0010;

	lut_sub lut_7464 ({i_0_, g125}, g710);
	defparam lut_7464.LUT_SIZE = 2;
	defparam lut_7464.mask = 4'b0010;

	lut_sub lut_7469 ({i_38_, g255, i_32_, i_5_}, g711);
	defparam lut_7469.LUT_SIZE = 4;
	defparam lut_7469.mask = 16'hbfff;

	lut_sub lut_7489 ({g713, g714}, g712);
	defparam lut_7489.LUT_SIZE = 2;
	defparam lut_7489.mask = 4'b1000;

	lut_sub lut_7494 ({i_37_, g715}, g713);
	defparam lut_7494.LUT_SIZE = 2;
	defparam lut_7494.mask = 4'b0100;

	lut_sub lut_7499 ({i_37_, g717}, g714);
	defparam lut_7499.LUT_SIZE = 2;
	defparam lut_7499.mask = 4'b0001;

	lut_sub lut_7504 ({i_36_, g716}, g715);
	defparam lut_7504.LUT_SIZE = 2;
	defparam lut_7504.mask = 4'b0010;

	lut_sub lut_7509 ({i_36_, g720}, g716);
	defparam lut_7509.LUT_SIZE = 2;
	defparam lut_7509.mask = 4'b0001;

	lut_sub lut_7515 ({g718, g719}, g717);
	defparam lut_7515.LUT_SIZE = 2;
	defparam lut_7515.mask = 4'b1000;

	lut_sub lut_7520 ({i_36_, g721}, g718);
	defparam lut_7520.LUT_SIZE = 2;
	defparam lut_7520.mask = 4'b0100;

	lut_sub lut_7525 ({i_36_, g722}, g719);
	defparam lut_7525.LUT_SIZE = 2;
	defparam lut_7525.mask = 4'b0001;

	lut_sub lut_7530 ({i_40_, i_39_, g10, i_38_}, g720);
	defparam lut_7530.LUT_SIZE = 4;
	defparam lut_7530.mask = 16'hfffb;

	lut_sub lut_7549 ({i_40_, i_39_, g49, i_38_}, g721);
	defparam lut_7549.LUT_SIZE = 4;
	defparam lut_7549.mask = 16'hfffb;

	lut_sub lut_7568 ({i_40_, g10, i_38_}, g722);
	defparam lut_7568.LUT_SIZE = 3;
	defparam lut_7568.mask = 8'hf7;

	lut_sub lut_7579 ({i_40_, g724}, g723);
	defparam lut_7579.LUT_SIZE = 2;
	defparam lut_7579.mask = 4'b0001;

	lut_sub lut_7585 ({g725, g726}, g724);
	defparam lut_7585.LUT_SIZE = 2;
	defparam lut_7585.mask = 4'b1000;

	lut_sub lut_7591 ({g22, g727}, g725);
	defparam lut_7591.LUT_SIZE = 2;
	defparam lut_7591.mask = 4'b0100;

	lut_sub lut_7597 ({g22, g728}, g726);
	defparam lut_7597.LUT_SIZE = 2;
	defparam lut_7597.mask = 4'b0001;

	lut_sub lut_7603 ({g351, g349}, g727);
	defparam lut_7603.LUT_SIZE = 2;
	defparam lut_7603.mask = 4'b0100;

	lut_sub lut_7611 ({g350, g98, g1, g349}, g728);
	defparam lut_7611.LUT_SIZE = 4;
	defparam lut_7611.mask = 16'h5551;

	lut_sub lut_7623 ({g730, g731}, g729);
	defparam lut_7623.LUT_SIZE = 2;
	defparam lut_7623.mask = 4'b1000;

	lut_sub lut_7629 ({g30, g732}, g730);
	defparam lut_7629.LUT_SIZE = 2;
	defparam lut_7629.mask = 4'b0100;

	lut_sub lut_7635 ({g30, g735}, g731);
	defparam lut_7635.LUT_SIZE = 2;
	defparam lut_7635.mask = 4'b0001;

	lut_sub lut_7641 ({g733, g734}, g732);
	defparam lut_7641.LUT_SIZE = 2;
	defparam lut_7641.mask = 4'b1000;

	lut_sub lut_7646 ({i_37_, g737}, g733);
	defparam lut_7646.LUT_SIZE = 2;
	defparam lut_7646.mask = 4'b0100;

	lut_sub lut_7651 ({i_37_, g738}, g734);
	defparam lut_7651.LUT_SIZE = 2;
	defparam lut_7651.mask = 4'b0001;

	lut_sub lut_7656 ({i_37_, g736}, g735);
	defparam lut_7656.LUT_SIZE = 2;
	defparam lut_7656.mask = 4'b1000;

	lut_sub lut_7661 ({i_37_, g739}, g736);
	defparam lut_7661.LUT_SIZE = 2;
	defparam lut_7661.mask = 4'b0100;

	lut_sub lut_7668 ({g5, g122, g266}, g737);
	defparam lut_7668.LUT_SIZE = 3;
	defparam lut_7668.mask = 8'hfb;

	lut_sub lut_7680 ({g267, g94}, g738);
	defparam lut_7680.LUT_SIZE = 2;
	defparam lut_7680.mask = 4'b1101;

	lut_sub lut_7689 ({g5, g122, g266}, g739);
	defparam lut_7689.LUT_SIZE = 3;
	defparam lut_7689.mask = 8'hfb;

	lut_sub lut_7700 ({i_36_, g741}, g740);
	defparam lut_7700.LUT_SIZE = 2;
	defparam lut_7700.mask = 4'b0010;

	lut_sub lut_7705 ({i_36_, g742}, g741);
	defparam lut_7705.LUT_SIZE = 2;
	defparam lut_7705.mask = 4'b0001;

	lut_sub lut_7711 ({g743, g744}, g742);
	defparam lut_7711.LUT_SIZE = 2;
	defparam lut_7711.mask = 4'b1000;

	lut_sub lut_7716 ({i_40_, g745}, g743);
	defparam lut_7716.LUT_SIZE = 2;
	defparam lut_7716.mask = 4'b0100;

	lut_sub lut_7721 ({i_40_, g746}, g744);
	defparam lut_7721.LUT_SIZE = 2;
	defparam lut_7721.mask = 4'b0001;

	lut_sub lut_7726 ({i_37_, i_39_, i_35_, g92}, g745);
	defparam lut_7726.LUT_SIZE = 4;
	defparam lut_7726.mask = 16'hffef;

	lut_sub lut_7745 ({i_37_, i_39_, i_38_, g92}, g746);
	defparam lut_7745.LUT_SIZE = 4;
	defparam lut_7745.mask = 16'hfffe;

	lut_sub lut_7765 ({g748, g749}, g747);
	defparam lut_7765.LUT_SIZE = 2;
	defparam lut_7765.mask = 4'b1000;

	lut_sub lut_7771 ({g152, g750}, g748);
	defparam lut_7771.LUT_SIZE = 2;
	defparam lut_7771.mask = 4'b0100;

	lut_sub lut_7777 ({g152, g753}, g749);
	defparam lut_7777.LUT_SIZE = 2;
	defparam lut_7777.mask = 4'b0001;

	lut_sub lut_7783 ({g751, g752}, g750);
	defparam lut_7783.LUT_SIZE = 2;
	defparam lut_7783.mask = 4'b1000;

	lut_sub lut_7788 ({i_18_, g756}, g751);
	defparam lut_7788.LUT_SIZE = 2;
	defparam lut_7788.mask = 4'b0100;

	lut_sub lut_7793 ({i_18_, g757}, g752);
	defparam lut_7793.LUT_SIZE = 2;
	defparam lut_7793.mask = 4'b0001;

	lut_sub lut_7799 ({g754, g755}, g753);
	defparam lut_7799.LUT_SIZE = 2;
	defparam lut_7799.mask = 4'b1000;

	lut_sub lut_7804 ({i_18_, g758}, g754);
	defparam lut_7804.LUT_SIZE = 2;
	defparam lut_7804.mask = 4'b0100;

	lut_sub lut_7809 ({i_18_, g759}, g755);
	defparam lut_7809.LUT_SIZE = 2;
	defparam lut_7809.mask = 4'b0001;

	lut_sub lut_7817 ({g34, g156, g18, g154}, g756);
	defparam lut_7817.LUT_SIZE = 4;
	defparam lut_7817.mask = 16'hfac8;

	lut_sub lut_7833 ({g34, g156, g157, g154}, g757);
	defparam lut_7833.LUT_SIZE = 4;
	defparam lut_7833.mask = 16'hfaea;

	lut_sub lut_7849 ({g156, g154}, g758);
	defparam lut_7849.LUT_SIZE = 2;
	defparam lut_7849.mask = 4'b1110;

	lut_sub lut_7859 ({g34, g156, g157, g154}, g759);
	defparam lut_7859.LUT_SIZE = 4;
	defparam lut_7859.mask = 16'hfaea;


endmodule