module ks_alu4_qmap_map (clk, sk, in, outreg);

input [13:0] in;
reg [13:0] inreg;
input clk;
output reg [7:0] outreg;
wire [7:0] out;

  wire a, b, c, d, e, f, g, h, i, j, k, l, m, n;
  wire o, p, q, r, s, t, u, v;

	input [127 : 0] sk /* synthesis noprune */;

always@(posedge clk)
begin
	inreg <= in;
	outreg <= out;
end

assign {a, b, c, d, e, f, g, h, i, j, k, l, m, n}=inreg;
assign out={o, p, q, r, s, t, u, v};

	wire g163, g121, g179, g1, g2, g3, g4, g182, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16, g17;
	wire g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29, g30, g31, g32, g33, g34, g35, g36, g37, g38;
	wire g39, g40, g41, g42, g43, g44, g45, g46, g47, g48, g49, g50, g51, g52, g53, g54, g55, g56, g57, g206, g58;
	wire g59, g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g70, g71, g72, g73, g74, g75, g76, g77, g78, g80;
	wire g81, g82, g83, g84, g85, g86, g87, g88, g89, g90, g91, g92, g93, g94, g95, g96, g97, g98, g99, g100, g101;
	wire g102, g103, g104, g105, g106, g107, g108, g109, g110, g111, g112, g113, g114, g115, g116, g117, g118, g119, g120, g122, g123;
	wire g124, g125, g126, g127, g128, g129, g130, g131, g132, g133, g134, g135, g136, g137, g138, g139, g140, g141, g142, g143, g144;
	wire g145, g146, g147, g148, g149, g150, g151, g152, g153, g154, g155, g156, g157, g158, g159, g160, g161, g164, g165, g166, g167;
	wire g168, g169, g170, g171, g183, g172, g173, g174, g175, g176, g178, g180, g181, g184, g185, g186, g189, g187, g188, g190, g191;
	wire g192, g194, g195, g196, g199, g197, g198, g202, g203, g200, g201, g204, g205, g207, g208, g209, g212, g210, g211, g215, g216;
	wire g213, g214, g217, g218, g220, g221, g222, g225, g223, g224, g228, g229, g226, g227, g230, g231;

	assign s = (((sk[0]) & (!g163)));
	assign t = (((sk[1]) & (g121)));
	assign v = (((sk[2]) & (!g179)));
	assign g1 = (((k) & (!sk[3]) & (!l)) + ((k) & (!sk[3]) & (!l)));
	assign g2 = (((k) & (!l) & (!n) & (!sk[4]) & (!i) & (!j)) + ((!k) & (!l) & (n) & (!sk[4]) & (!i) & (!j)) + ((!k) & (!l) & (!n) & (!sk[4]) & (i) & (!j)) + ((k) & (!l) & (!n) & (!sk[4]) & (i) & (j)) + ((!k) & (!l) & (n) & (!sk[4]) & (!i) & (j)) + ((!k) & (l) & (n) & (!sk[4]) & (!i) & (j)) + ((k) & (l) & (!n) & (!sk[4]) & (i) & (!j)));
	assign g3 = (((k) & (!l) & (!n) & (!i) & (!sk[5]) & (!j)) + ((!k) & (!l) & (n) & (!i) & (!sk[5]) & (!j)) + ((!k) & (!l) & (!n) & (i) & (!sk[5]) & (!j)) + ((!k) & (!l) & (!n) & (!i) & (sk[5]) & (!j)) + ((!k) & (!l) & (!n) & (!i) & (sk[5]) & (!j)));
	assign g4 = (((k) & (!l) & (!n) & (!i) & (!sk[6]) & (!j)) + ((!k) & (!l) & (n) & (!i) & (!sk[6]) & (!j)) + ((!k) & (!l) & (!n) & (i) & (!sk[6]) & (!j)) + ((k) & (!l) & (n) & (i) & (!sk[6]) & (!j)) + ((!k) & (!l) & (!n) & (i) & (!sk[6]) & (!j)));
	assign g5 = (((!k) & (l) & (!i) & (a) & (!e) & (!g182)) + ((k) & (l) & (!i) & (!a) & (!e) & (g182)) + ((!k) & (!l) & (!i) & (!a) & (!e) & (g182)) + ((k) & (!l) & (!i) & (!a) & (!e) & (!g182)) + ((!k) & (!l) & (i) & (!a) & (!e) & (!g182)) + ((k) & (!l) & (i) & (!a) & (!e) & (!g182)) + ((!k) & (l) & (i) & (!a) & (e) & (!g182)));
	assign g6 = (((!k) & (l) & (!i) & (!a) & (e) & (!g182)) + ((k) & (!l) & (i) & (a) & (!e) & (g182)) + ((k) & (!l) & (!i) & (!a) & (!e) & (!g182)));
	assign g7 = (((!n) & (!i) & (!sk[9]) & (j) & (!g1)) + ((!n) & (!i) & (!sk[9]) & (!j) & (g1)) + ((n) & (i) & (!sk[9]) & (!j) & (!g1)) + ((n) & (i) & (!sk[9]) & (!j) & (g1)));
	assign g8 = (((!sk[10]) & (i) & (!j)) + ((!sk[10]) & (i) & (j)));
	assign g9 = (((!n) & (!sk[11]) & (!g8) & (g1)) + ((n) & (!sk[11]) & (g8) & (!g1)) + ((n) & (!sk[11]) & (g8) & (g1)));
	assign g10 = (((!n) & (!sk[12]) & (!i) & (j) & (!g1)) + ((!n) & (!sk[12]) & (!i) & (!j) & (g1)) + ((n) & (!sk[12]) & (i) & (!j) & (!g1)) + ((n) & (!sk[12]) & (!i) & (!j) & (g1)));
	assign g11 = (((!n) & (!sk[13]) & (!i) & (j)) + ((n) & (!sk[13]) & (i) & (!j)) + ((n) & (!sk[13]) & (!i) & (j)));
	assign g12 = (((!sk[14]) & (l) & (!g11)) + ((!sk[14]) & (l) & (g11)));
	assign g13 = (((!sk[15]) & (a) & (!g182) & (!g9) & (!g10) & (!g12)) + ((!sk[15]) & (!a) & (!g182) & (g9) & (!g10) & (!g12)) + ((!sk[15]) & (!a) & (!g182) & (!g9) & (g10) & (!g12)) + ((sk[15]) & (!a) & (!g182) & (!g9) & (!g10) & (!g12)) + ((sk[15]) & (!a) & (g182) & (!g9) & (!g10) & (!g12)) + ((sk[15]) & (!a) & (g182) & (!g9) & (!g10) & (!g12)) + ((!sk[15]) & (a) & (!g182) & (!g9) & (!g10) & (!g12)));
	assign g14 = (((!a) & (!e) & (g7) & (!sk[16]) & (!g13)) + ((!a) & (!e) & (!g7) & (!sk[16]) & (g13)) + ((!a) & (!e) & (!g7) & (!sk[16]) & (g13)) + ((!a) & (!e) & (!g7) & (!sk[16]) & (g13)) + ((a) & (e) & (!g7) & (!sk[16]) & (!g13)));
	assign g15 = (((k) & (!sk[17]) & (!g12)) + ((!k) & (sk[17]) & (g12)));
	assign g16 = (((a) & (!e) & (!g7) & (!sk[18]) & (!g13) & (!g15)) + ((!a) & (!e) & (g7) & (!sk[18]) & (!g13) & (!g15)) + ((!a) & (!e) & (!g7) & (!sk[18]) & (g13) & (!g15)) + ((!a) & (!e) & (g7) & (!sk[18]) & (g13) & (!g15)) + ((!a) & (!e) & (g7) & (!sk[18]) & (g13) & (!g15)) + ((a) & (e) & (!g7) & (!sk[18]) & (!g13) & (g15)));
	assign g17 = (((!sk[19]) & (!k) & (!i) & (j)) + ((!sk[19]) & (k) & (i) & (!j)) + ((!sk[19]) & (!k) & (!i) & (j)));
	assign g18 = (((!sk[20]) & (l) & (!g17)) + ((!sk[20]) & (l) & (g17)));
	assign g19 = (((!l) & (!i) & (!j) & (a) & (!e) & (!g182)) + ((!l) & (i) & (!j) & (!a) & (e) & (!g182)) + ((!l) & (i) & (!j) & (a) & (!e) & (!g182)) + ((!l) & (!i) & (j) & (!a) & (!e) & (g182)) + ((!l) & (!i) & (!j) & (a) & (!e) & (!g182)));
	assign g20 = (((k) & (l) & (!i) & (!j) & (!a) & (g182)) + ((!k) & (l) & (!i) & (!j) & (!a) & (g182)) + ((k) & (l) & (!i) & (!j) & (a) & (!g182)) + ((k) & (l) & (!i) & (!j) & (a) & (!g182)));
	assign g21 = (((k) & (!g14) & (!g16) & (!g18) & (!g19) & (!g20)) + ((!k) & (!g14) & (!g16) & (!g18) & (!g19) & (!g20)) + ((k) & (!g14) & (g16) & (!g18) & (!g19) & (!g20)) + ((k) & (g14) & (!g16) & (!g18) & (!g19) & (!g20)) + ((!k) & (!g14) & (g16) & (!g18) & (!g19) & (!g20)) + ((!k) & (g14) & (!g16) & (!g18) & (!g19) & (!g20)));
	assign g22 = (((!sk[24]) & (!l) & (!n) & (j)) + ((!sk[24]) & (l) & (n) & (!j)) + ((sk[24]) & (!l) & (n) & (!j)));
	assign g23 = (((!k) & (!i) & (!sk[25]) & (g22)) + ((k) & (i) & (!sk[25]) & (!g22)) + ((k) & (i) & (!sk[25]) & (g22)));
	assign g24 = (((!g182) & (!sk[26]) & (!g16) & (g23)) + ((g182) & (!sk[26]) & (g16) & (!g23)) + ((!g182) & (!sk[26]) & (g16) & (g23)) + ((g182) & (!sk[26]) & (!g16) & (g23)));
	assign g25 = (((k) & (l) & (n) & (g8) & (!a) & (!g14)) + ((k) & (!l) & (n) & (g8) & (!a) & (g14)));
	assign g26 = (((i) & (!sk[28]) & (!g22)) + ((!i) & (sk[28]) & (g22)));
	assign g27 = (((!sk[29]) & (k) & (!l) & (!n) & (!i) & (!j)) + ((!sk[29]) & (!k) & (!l) & (n) & (!i) & (!j)) + ((!sk[29]) & (!k) & (!l) & (!n) & (i) & (!j)) + ((!sk[29]) & (!k) & (l) & (n) & (i) & (j)) + ((!sk[29]) & (k) & (!l) & (n) & (!i) & (j)));
	assign g28 = (((i) & (!sk[30]) & (!g22)) + ((i) & (!sk[30]) & (g22)));
	assign g29 = (((!sk[31]) & (k) & (!e) & (!g182) & (!g27) & (!g28)) + ((!sk[31]) & (!k) & (!e) & (g182) & (!g27) & (!g28)) + ((!sk[31]) & (!k) & (!e) & (!g182) & (g27) & (!g28)) + ((sk[31]) & (!k) & (e) & (!g182) & (!g27) & (g28)));
	assign g30 = (((k) & (!a) & (!sk[32]) & (!g14) & (!g26) & (!g29)) + ((!k) & (!a) & (!sk[32]) & (g14) & (!g26) & (!g29)) + ((!k) & (!a) & (!sk[32]) & (!g14) & (g26) & (!g29)) + ((!k) & (!a) & (!sk[32]) & (g14) & (!g26) & (!g29)) + ((!k) & (!a) & (sk[32]) & (!g14) & (!g26) & (!g29)) + ((!k) & (!a) & (sk[32]) & (!g14) & (!g26) & (!g29)) + ((!k) & (a) & (sk[32]) & (!g14) & (!g26) & (!g29)));
	assign g31 = (((!n) & (!g21) & (!sk[33]) & (g24) & (!g25) & (!g30)) + ((!n) & (!g21) & (!sk[33]) & (!g24) & (g25) & (!g30)) + ((n) & (!g21) & (!sk[33]) & (!g24) & (!g25) & (!g30)) + ((n) & (!g21) & (!sk[33]) & (!g24) & (!g25) & (!g30)) + ((!n) & (!g21) & (sk[33]) & (!g24) & (!g25) & (!g30)));
	assign g32 = (((!k) & (!n) & (!sk[34]) & (i)) + ((k) & (n) & (!sk[34]) & (!i)) + ((!k) & (!n) & (sk[34]) & (!i)));
	assign g33 = (((k) & (!l) & (!n) & (!sk[35]) & (!i) & (!j)) + ((!k) & (!l) & (n) & (!sk[35]) & (!i) & (!j)) + ((!k) & (!l) & (!n) & (!sk[35]) & (i) & (!j)) + ((!k) & (!l) & (n) & (!sk[35]) & (i) & (j)) + ((k) & (l) & (!n) & (!sk[35]) & (!i) & (!j)));
	assign g34 = (((k) & (!sk[36]) & (!l) & (!n) & (!i) & (!j)) + ((!k) & (!sk[36]) & (!l) & (n) & (!i) & (!j)) + ((!k) & (!sk[36]) & (!l) & (!n) & (i) & (!j)) + ((!k) & (sk[36]) & (l) & (!n) & (!i) & (j)) + ((k) & (!sk[36]) & (!l) & (!n) & (!i) & (j)));
	assign g35 = (((k) & (!sk[37]) & (!l) & (!n) & (!i) & (!j)) + ((!k) & (!sk[37]) & (!l) & (n) & (!i) & (!j)) + ((!k) & (!sk[37]) & (!l) & (!n) & (i) & (!j)) + ((k) & (!sk[37]) & (l) & (!n) & (!i) & (!j)) + ((!k) & (sk[37]) & (l) & (!n) & (!i) & (!j)));
	assign g36 = (((g33) & (!a) & (!e) & (!sk[38]) & (!g34) & (!g35)) + ((!g33) & (!a) & (e) & (!sk[38]) & (!g34) & (!g35)) + ((!g33) & (!a) & (!e) & (!sk[38]) & (g34) & (!g35)) + ((!g33) & (!a) & (!e) & (sk[38]) & (!g34) & (!g35)) + ((!g33) & (!a) & (!e) & (sk[38]) & (!g34) & (!g35)) + ((!g33) & (!a) & (!e) & (sk[38]) & (!g34) & (!g35)));
	assign g37 = (((!e) & (!g32) & (!g182) & (!sk[39]) & (g36)) + ((!e) & (!g32) & (!g182) & (sk[39]) & (!g36)) + ((e) & (g32) & (g182) & (!sk[39]) & (!g36)) + ((!e) & (!g32) & (g182) & (!sk[39]) & (!g36)) + ((e) & (g32) & (!g182) & (!sk[39]) & (!g36)));
	assign g38 = (((k) & (!sk[40]) & (!l) & (!n) & (!i) & (!j)) + ((!k) & (!sk[40]) & (!l) & (n) & (!i) & (!j)) + ((!k) & (!sk[40]) & (!l) & (!n) & (i) & (!j)) + ((k) & (!sk[40]) & (l) & (n) & (!i) & (!j)));
	assign g39 = (((a) & (!e) & (!g1) & (!sk[41]) & (!f) & (!b)) + ((!a) & (!e) & (g1) & (!sk[41]) & (!f) & (!b)) + ((!a) & (!e) & (!g1) & (!sk[41]) & (f) & (!b)) + ((a) & (!e) & (!g1) & (!sk[41]) & (!f) & (b)) + ((!a) & (!e) & (!g1) & (sk[41]) & (!f) & (b)) + ((a) & (!e) & (g1) & (!sk[41]) & (f) & (!b)) + ((!a) & (!e) & (g1) & (!sk[41]) & (f) & (!b)) + ((!a) & (e) & (!g1) & (sk[41]) & (!f) & (!b)));
	assign g40 = (((!g2) & (!sk[42]) & (!g3) & (f) & (!b)) + ((!g2) & (!sk[42]) & (!g3) & (!f) & (b)) + ((g2) & (sk[42]) & (!g3) & (!f) & (!b)) + ((!g2) & (sk[42]) & (g3) & (!f) & (!b)) + ((g2) & (!sk[42]) & (g3) & (!f) & (!b)));
	assign g41 = (((!sk[43]) & (k) & (!l) & (!n) & (!i) & (!j)) + ((!sk[43]) & (!k) & (!l) & (n) & (!i) & (!j)) + ((!sk[43]) & (!k) & (!l) & (!n) & (i) & (!j)) + ((!sk[43]) & (k) & (!l) & (n) & (!i) & (!j)) + ((!sk[43]) & (k) & (!l) & (!n) & (!i) & (!j)) + ((!sk[43]) & (!k) & (l) & (n) & (i) & (j)) + ((!sk[43]) & (!k) & (l) & (n) & (!i) & (!j)));
	assign g42 = (((n) & (!i) & (!sk[44]) & (!a) & (!e) & (!g1)) + ((!n) & (!i) & (!sk[44]) & (a) & (!e) & (!g1)) + ((!n) & (!i) & (!sk[44]) & (!a) & (e) & (!g1)) + ((n) & (!i) & (!sk[44]) & (!a) & (e) & (g1)));
	assign g43 = (((!sk[45]) & (g4) & (!f) & (!b) & (!g41) & (!g42)) + ((!sk[45]) & (g4) & (f) & (!b) & (!g41) & (!g42)) + ((!sk[45]) & (!g4) & (!f) & (b) & (!g41) & (!g42)) + ((!sk[45]) & (g4) & (!f) & (b) & (!g41) & (!g42)) + ((!sk[45]) & (!g4) & (!f) & (!b) & (g41) & (!g42)) + ((!sk[45]) & (!g4) & (f) & (b) & (g41) & (!g42)) + ((!sk[45]) & (!g4) & (f) & (b) & (!g41) & (g42)));
	assign g44 = (((!a) & (!g11) & (!g38) & (!g39) & (g40) & (!g43)) + ((!a) & (!g11) & (!g38) & (!g39) & (!g40) & (g43)) + ((a) & (!g11) & (g38) & (!g39) & (!g40) & (!g43)) + ((!a) & (g11) & (!g38) & (g39) & (!g40) & (!g43)));
	assign g45 = (((g7) & (!sk[47]) & (!f)) + ((g7) & (!sk[47]) & (f)));
	assign g46 = (((!g9) & (!g10) & (!g12) & (!b) & (g44) & (!g45)) + ((!g9) & (!g10) & (!g12) & (!b) & (!g44) & (!g45)) + ((!g9) & (!g10) & (!g12) & (!b) & (g44) & (!g45)) + ((!g9) & (!g10) & (!g12) & (!b) & (!g44) & (!g45)));
	assign g47 = (((!g15) & (!sk[49]) & (!f) & (b)) + ((g15) & (!sk[49]) & (f) & (!b)) + ((g15) & (!sk[49]) & (f) & (b)));
	assign g48 = (((!g7) & (!sk[50]) & (!g46) & (g47)) + ((g7) & (!sk[50]) & (g46) & (!g47)) + ((!g7) & (sk[50]) & (!g46) & (!g47)) + ((!g7) & (sk[50]) & (!g46) & (!g47)));
	assign g49 = (((!k) & (l) & (!i) & (j) & (a) & (e)));
	assign g50 = (((!sk[52]) & (a) & (!g182)) + ((!sk[52]) & (a) & (g182)));
	assign g51 = (((!k) & (!l) & (i) & (!sk[53]) & (!j)) + ((!k) & (!l) & (!i) & (!sk[53]) & (j)) + ((k) & (l) & (!i) & (!sk[53]) & (!j)) + ((k) & (l) & (!i) & (!sk[53]) & (!j)) + ((!k) & (l) & (!i) & (sk[53]) & (!j)));
	assign g52 = (((!g50) & (!sk[54]) & (!b) & (g44) & (!g51)) + ((!g50) & (!sk[54]) & (!b) & (!g44) & (g51)) + ((g50) & (!sk[54]) & (b) & (!g44) & (!g51)) + ((g50) & (!sk[54]) & (!b) & (!g44) & (g51)));
	assign g53 = (((!k) & (!sk[55]) & (!l) & (i) & (!j)) + ((!k) & (!sk[55]) & (!l) & (!i) & (j)) + ((k) & (!sk[55]) & (l) & (!i) & (!j)) + ((k) & (!sk[55]) & (l) & (!i) & (!j)) + ((!k) & (sk[55]) & (!l) & (!i) & (!j)));
	assign g54 = (((!sk[56]) & (l) & (!g17)) + ((sk[56]) & (!l) & (g17)));
	assign g55 = (((!k) & (!l) & (i) & (!sk[57]) & (!j)) + ((!k) & (!l) & (!i) & (!sk[57]) & (j)) + ((k) & (l) & (!i) & (!sk[57]) & (!j)) + ((!k) & (!l) & (!i) & (!sk[57]) & (j)) + ((!k) & (l) & (i) & (!sk[57]) & (j)));
	assign g56 = (((g182) & (g54) & (!sk[58]) & (!g55)) + ((!g182) & (g54) & (sk[58]) & (!g55)) + ((g182) & (!g54) & (!sk[58]) & (g55)) + ((!g182) & (!g54) & (!sk[58]) & (g55)));
	assign g57 = (((!k) & (!l) & (!sk[59]) & (g8)) + ((k) & (l) & (!sk[59]) & (!g8)) + ((!k) & (!l) & (sk[59]) & (!g8)));
	assign g58 = (((n) & (!g46) & (!g48) & (!g49) & (g52) & (!g206)) + ((n) & (!g46) & (!g48) & (!g49) & (!g52) & (g206)) + ((n) & (g46) & (g48) & (g49) & (!g52) & (!g206)));
	assign g59 = (((!sk[61]) & (g182) & (!g16) & (!g23) & (!g44) & (!g48)) + ((!sk[61]) & (!g182) & (!g16) & (g23) & (!g44) & (!g48)) + ((!sk[61]) & (!g182) & (!g16) & (!g23) & (g44) & (!g48)) + ((!sk[61]) & (!g182) & (!g16) & (g23) & (g44) & (g48)) + ((!sk[61]) & (!g182) & (!g16) & (g23) & (g44) & (g48)) + ((!sk[61]) & (!g182) & (!g16) & (g23) & (!g44) & (!g48)) + ((!sk[61]) & (!g182) & (!g16) & (g23) & (!g44) & (!g48)) + ((!sk[61]) & (g182) & (g16) & (g23) & (!g44) & (g48)) + ((!sk[61]) & (g182) & (g16) & (g23) & (g44) & (!g48)));
	assign g60 = (((!sk[62]) & (!k) & (!n) & (g8)) + ((!sk[62]) & (k) & (n) & (!g8)) + ((!sk[62]) & (k) & (n) & (g8)));
	assign g61 = (((l) & (!a) & (!g14) & (!b) & (!sk[63]) & (!g46)) + ((!l) & (!a) & (g14) & (!b) & (!sk[63]) & (!g46)) + ((!l) & (!a) & (!g14) & (b) & (!sk[63]) & (!g46)) + ((l) & (a) & (!g14) & (b) & (!sk[63]) & (!g46)) + ((l) & (!a) & (!g14) & (!b) & (!sk[63]) & (!g46)) + ((!l) & (!a) & (g14) & (!b) & (!sk[63]) & (g46)) + ((!l) & (!a) & (!g14) & (!b) & (sk[63]) & (!g46)));
	assign g62 = (((!sk[64]) & (g182) & (!g44)) + ((sk[64]) & (!g182) & (!g44)));
	assign g63 = (((!k) & (!sk[65]) & (!i) & (g22) & (!f)) + ((!k) & (!sk[65]) & (!i) & (!g22) & (f)) + ((k) & (!sk[65]) & (i) & (!g22) & (!f)) + ((!k) & (!sk[65]) & (i) & (g22) & (f)));
	assign g64 = (((l) & (!a) & (!e) & (!sk[66]) & (!f) & (!b)) + ((!l) & (!a) & (e) & (!sk[66]) & (!f) & (!b)) + ((!l) & (!a) & (!e) & (!sk[66]) & (f) & (!b)) + ((!l) & (!a) & (!e) & (!sk[66]) & (f) & (!b)) + ((!l) & (!a) & (!e) & (!sk[66]) & (f) & (!b)) + ((!l) & (a) & (e) & (!sk[66]) & (f) & (b)) + ((!l) & (!a) & (!e) & (sk[66]) & (!f) & (b)) + ((l) & (a) & (e) & (!sk[66]) & (!f) & (!b)) + ((!l) & (!a) & (!e) & (sk[66]) & (!f) & (b)));
	assign g65 = (((!k) & (!n) & (i) & (!sk[67]) & (!j)) + ((!k) & (!n) & (!i) & (!sk[67]) & (j)) + ((k) & (n) & (!i) & (!sk[67]) & (!j)) + ((!k) & (n) & (i) & (!sk[67]) & (!j)));
	assign g66 = (((g27) & (!g62) & (!g63) & (!g64) & (!sk[68]) & (!g65)) + ((!g27) & (!g62) & (g63) & (!g64) & (!sk[68]) & (!g65)) + ((!g27) & (!g62) & (!g63) & (g64) & (!sk[68]) & (!g65)) + ((!g27) & (!g62) & (!g63) & (!g64) & (sk[68]) & (!g65)) + ((!g27) & (!g62) & (!g63) & (!g64) & (sk[68]) & (!g65)) + ((!g27) & (!g62) & (!g63) & (!g64) & (sk[68]) & (!g65)) + ((!g27) & (!g62) & (!g63) & (!g64) & (sk[68]) & (!g65)));
	assign g67 = (((!a) & (!sk[69]) & (!e) & (g15)) + ((a) & (!sk[69]) & (e) & (!g15)) + ((a) & (!sk[69]) & (e) & (g15)));
	assign g68 = (((!sk[70]) & (!k) & (!l) & (g11)) + ((!sk[70]) & (k) & (l) & (!g11)) + ((!sk[70]) & (!k) & (l) & (g11)));
	assign g69 = (((!l) & (!sk[71]) & (!i) & (a) & (!e)) + ((!l) & (!sk[71]) & (!i) & (!a) & (e)) + ((l) & (!sk[71]) & (i) & (!a) & (!e)) + ((l) & (!sk[71]) & (!i) & (a) & (e)));
	assign g70 = (((!g7) & (!g67) & (!g46) & (g47) & (!g68) & (g69)) + ((!g7) & (!g67) & (g46) & (g47) & (g68) & (!g69)) + ((!g7) & (!g67) & (!g46) & (!g47) & (g68) & (!g69)) + ((g7) & (!g67) & (!g46) & (!g47) & (g68) & (!g69)));
	assign g71 = (((!k) & (!a) & (!g14) & (g26) & (b) & (g46)) + ((!k) & (!a) & (g14) & (g26) & (b) & (g46)) + ((!k) & (a) & (!g14) & (g26) & (b) & (!g46)) + ((k) & (!a) & (!g14) & (g26) & (!b) & (!g46)) + ((k) & (!a) & (g14) & (g26) & (!b) & (!g46)) + ((k) & (a) & (!g14) & (g26) & (!b) & (g46)));
	assign g72 = (((g60) & (!g61) & (!g66) & (!sk[74]) & (!g70) & (!g71)) + ((!g60) & (!g61) & (g66) & (!sk[74]) & (!g70) & (!g71)) + ((!g60) & (!g61) & (!g66) & (!sk[74]) & (g70) & (!g71)) + ((!g60) & (!g61) & (g66) & (!sk[74]) & (!g70) & (!g71)) + ((!g60) & (!g61) & (g66) & (!sk[74]) & (!g70) & (!g71)));
	assign g73 = (((!g58) & (!g59) & (!sk[75]) & (g72)) + ((g58) & (g59) & (!sk[75]) & (!g72)) + ((!g58) & (!g59) & (!sk[75]) & (g72)));
	assign g74 = (((!k) & (!l) & (i) & (!f) & (!b) & (g44)) + ((k) & (!l) & (!i) & (!f) & (!b) & (g44)) + ((!k) & (!l) & (!i) & (!f) & (!b) & (!g44)) + ((k) & (!l) & (i) & (f) & (!b) & (!g44)) + ((k) & (!l) & (i) & (f) & (!b) & (!g44)) + ((!k) & (!l) & (!i) & (f) & (!b) & (!g44)) + ((!k) & (!l) & (!i) & (!f) & (!b) & (!g44)) + ((!k) & (l) & (i) & (f) & (b) & (!g44)) + ((!k) & (l) & (i) & (!f) & (!b) & (!g44)) + ((k) & (l) & (i) & (!f) & (!b) & (!g44)));
	assign g75 = (((!k) & (l) & (!i) & (f) & (!b) & (!g44)) + ((k) & (!l) & (i) & (!f) & (b) & (g44)) + ((k) & (!l) & (!i) & (!f) & (!b) & (!g44)));
	assign g76 = (((!sk[78]) & (!g34) & (!g35) & (f) & (!b)) + ((!sk[78]) & (!g34) & (!g35) & (!f) & (b)) + ((!sk[78]) & (!g34) & (g35) & (!f) & (b)) + ((!sk[78]) & (g34) & (g35) & (!f) & (!b)) + ((!sk[78]) & (g34) & (!g35) & (f) & (b)));
	assign g77 = (((g33) & (!g32) & (!f) & (!g44) & (!sk[79]) & (!g76)) + ((!g33) & (!g32) & (f) & (!g44) & (!sk[79]) & (!g76)) + ((!g33) & (!g32) & (!f) & (g44) & (!sk[79]) & (!g76)) + ((!g33) & (!g32) & (!f) & (!g44) & (sk[79]) & (!g76)) + ((!g33) & (!g32) & (!f) & (!g44) & (sk[79]) & (!g76)) + ((!g33) & (!g32) & (!f) & (!g44) & (sk[79]) & (!g76)));
	assign g78 = (((n) & (!j) & (!g74) & (!g75) & (!sk[80]) & (!g77)) + ((!n) & (!j) & (g74) & (!g75) & (!sk[80]) & (!g77)) + ((!n) & (!j) & (!g74) & (g75) & (!sk[80]) & (!g77)) + ((n) & (!j) & (!g74) & (!g75) & (!sk[80]) & (g77)) + ((!n) & (!j) & (g74) & (!g75) & (!sk[80]) & (g77)) + ((!n) & (j) & (!g74) & (!g75) & (sk[80]) & (g77)));
	assign p = (((!sk[81]) & (!n) & (!m) & (g31) & (!g73) & (!g78)) + ((!sk[81]) & (!n) & (!m) & (!g31) & (g73) & (!g78)) + ((sk[81]) & (!n) & (!m) & (!g31) & (!g73) & (!g78)) + ((!sk[81]) & (n) & (m) & (!g31) & (!g73) & (!g78)) + ((!sk[81]) & (n) & (!m) & (!g31) & (!g73) & (!g78)) + ((!sk[81]) & (n) & (!m) & (g31) & (g73) & (!g78)));
	assign g80 = (((m) & (!g31) & (!g58) & (!g59) & (!sk[82]) & (!g72)) + ((!m) & (!g31) & (!g58) & (!g59) & (sk[82]) & (!g72)) + ((!m) & (!g31) & (g58) & (!g59) & (!sk[82]) & (!g72)) + ((!m) & (!g31) & (!g58) & (g59) & (!sk[82]) & (!g72)) + ((!m) & (!g31) & (!g58) & (!g59) & (sk[82]) & (g72)));
	assign g81 = (((!a) & (!sk[83]) & (!e) & (!f) & (b)) + ((!a) & (!sk[83]) & (!e) & (f) & (!b)) + ((a) & (!sk[83]) & (e) & (!f) & (!b)) + ((!a) & (!sk[83]) & (e) & (f) & (!b)) + ((!a) & (sk[83]) & (e) & (!f) & (!b)));
	assign g82 = (((g1) & (!sk[84]) & (!g11) & (!c) & (!g) & (!g81)) + ((!g1) & (!sk[84]) & (!g11) & (c) & (!g) & (!g81)) + ((!g1) & (!sk[84]) & (!g11) & (!c) & (g) & (!g81)) + ((!g1) & (!sk[84]) & (g11) & (c) & (!g) & (!g81)) + ((g1) & (!sk[84]) & (g11) & (!c) & (g) & (!g81)));
	assign g83 = (((!j) & (!g1) & (!sk[85]) & (c) & (!g)) + ((!j) & (!g1) & (!sk[85]) & (!c) & (g)) + ((!j) & (g1) & (!sk[85]) & (c) & (g)) + ((j) & (!g1) & (sk[85]) & (!c) & (!g)) + ((j) & (g1) & (!sk[85]) & (!c) & (!g)));
	assign g84 = (((!n) & (!i) & (g81) & (!sk[86]) & (!g83)) + ((!n) & (!i) & (!g81) & (!sk[86]) & (g83)) + ((n) & (i) & (!g81) & (!sk[86]) & (!g83)) + ((n) & (!i) & (g81) & (!sk[86]) & (g83)));
	assign g85 = (((!g2) & (!sk[87]) & (!g3) & (c) & (!g)) + ((!g2) & (!sk[87]) & (!g3) & (!c) & (g)) + ((!g2) & (sk[87]) & (g3) & (!c) & (!g)) + ((g2) & (sk[87]) & (!g3) & (!c) & (!g)) + ((g2) & (!sk[87]) & (g3) & (!c) & (!g)));
	assign g86 = (((g4) & (!sk[88]) & (!g41) & (c) & (!g)) + ((!g4) & (!sk[88]) & (!g41) & (c) & (!g)) + ((g4) & (!sk[88]) & (!g41) & (!c) & (g)) + ((!g4) & (!sk[88]) & (!g41) & (!c) & (g)) + ((g4) & (!sk[88]) & (g41) & (!c) & (!g)) + ((!g4) & (!sk[88]) & (g41) & (c) & (g)));
	assign g87 = (((b) & (!sk[89]) & (!g38) & (!g84) & (!g85) & (!g86)) + ((!b) & (!sk[89]) & (!g38) & (g84) & (!g85) & (!g86)) + ((!b) & (!sk[89]) & (!g38) & (!g84) & (g85) & (!g86)) + ((!b) & (sk[89]) & (!g38) & (!g84) & (!g85) & (!g86)) + ((!b) & (sk[89]) & (!g38) & (!g84) & (!g85) & (!g86)));
	assign g88 = (((!g9) & (!g12) & (!sk[90]) & (c)) + ((g9) & (g12) & (!sk[90]) & (!c)) + ((!g9) & (!g12) & (sk[90]) & (!c)) + ((!g9) & (!g12) & (!sk[90]) & (c)));
	assign g89 = (((!g7) & (!sk[91]) & (!g12) & (c) & (!g)) + ((!g7) & (!sk[91]) & (g12) & (c) & (!g)) + ((!g7) & (!sk[91]) & (!g12) & (!c) & (g)) + ((g7) & (!sk[91]) & (g12) & (!c) & (!g)) + ((g7) & (!sk[91]) & (!g12) & (c) & (g)));
	assign g90 = (((g10) & (!sk[92]) & (!g82) & (!g87) & (!g88) & (!g89)) + ((!g10) & (!sk[92]) & (!g82) & (g87) & (!g88) & (!g89)) + ((!g10) & (!sk[92]) & (!g82) & (!g87) & (g88) & (!g89)) + ((!g10) & (!sk[92]) & (g82) & (!g87) & (g88) & (!g89)) + ((!g10) & (!sk[92]) & (!g82) & (!g87) & (g88) & (!g89)) + ((!g10) & (!sk[92]) & (!g82) & (g87) & (!g88) & (!g89)));
	assign g91 = (((a) & (!sk[93]) & (!g14) & (!b) & (!g46) & (!g90)) + ((!a) & (!sk[93]) & (!g14) & (b) & (!g46) & (!g90)) + ((!a) & (!sk[93]) & (!g14) & (!b) & (g46) & (!g90)) + ((!a) & (!sk[93]) & (!g14) & (b) & (!g46) & (g90)) + ((!a) & (!sk[93]) & (!g14) & (!b) & (g46) & (!g90)) + ((!a) & (!sk[93]) & (g14) & (!b) & (g46) & (!g90)) + ((!a) & (!sk[93]) & (!g14) & (!b) & (g46) & (!g90)) + ((a) & (!sk[93]) & (!g14) & (b) & (!g46) & (g90)) + ((a) & (!sk[93]) & (!g14) & (!b) & (!g46) & (g90)) + ((!a) & (sk[93]) & (!g14) & (!b) & (!g46) & (!g90)) + ((!a) & (sk[93]) & (g14) & (!b) & (!g46) & (!g90)));
	assign g92 = (((g50) & (b) & (!sk[94]) & (!g44)) + ((g50) & (!b) & (!sk[94]) & (g44)) + ((!g50) & (b) & (!sk[94]) & (g44)) + ((!g50) & (!b) & (!sk[94]) & (g44)));
	assign g93 = (((g82) & (!sk[95]) & (!g87)) + ((!g82) & (sk[95]) & (g87)));
	assign g94 = (((n) & (!g53) & (g57) & (!sk[96]) & (!g92) & (!g93)) + ((n) & (!g53) & (!g57) & (!sk[96]) & (!g92) & (!g93)) + ((!n) & (!g53) & (g57) & (!sk[96]) & (!g92) & (!g93)) + ((!n) & (!g53) & (!g57) & (!sk[96]) & (g92) & (!g93)) + ((n) & (g53) & (!g57) & (!sk[96]) & (!g92) & (g93)));
	assign g95 = (((!sk[97]) & (!l) & (!a) & (b) & (!g60)) + ((!sk[97]) & (!l) & (!a) & (!b) & (g60)) + ((!sk[97]) & (l) & (a) & (!b) & (!g60)) + ((!sk[97]) & (l) & (a) & (!b) & (g60)) + ((!sk[97]) & (l) & (!a) & (b) & (g60)));
	assign g96 = (((!a) & (!e) & (f) & (!sk[98]) & (!b)) + ((!a) & (!e) & (f) & (!sk[98]) & (b)) + ((!a) & (!e) & (!f) & (!sk[98]) & (b)) + ((a) & (e) & (f) & (!sk[98]) & (!b)) + ((a) & (e) & (!f) & (!sk[98]) & (!b)) + ((a) & (e) & (!f) & (!sk[98]) & (b)));
	assign g97 = (((!g65) & (!sk[99]) & (!g) & (g95) & (!g96)) + ((!g65) & (sk[99]) & (!g) & (!g95) & (!g96)) + ((!g65) & (!sk[99]) & (!g) & (!g95) & (g96)) + ((!g65) & (!sk[99]) & (!g) & (!g95) & (g96)) + ((g65) & (!sk[99]) & (g) & (!g95) & (!g96)));
	assign g98 = (((g26) & (!sk[100]) & (!c) & (!g91) & (!g94) & (!g97)) + ((!g26) & (!sk[100]) & (!c) & (g91) & (!g94) & (!g97)) + ((!g26) & (!sk[100]) & (!c) & (!g91) & (g94) & (!g97)) + ((!g26) & (!sk[100]) & (c) & (!g91) & (g94) & (!g97)) + ((g26) & (!sk[100]) & (c) & (!g91) & (!g94) & (!g97)) + ((!g26) & (sk[100]) & (c) & (!g91) & (!g94) & (!g97)));
	assign g99 = (((!l) & (!g65) & (!sk[101]) & (g) & (!g96)) + ((!l) & (!g65) & (!sk[101]) & (!g) & (g96)) + ((l) & (g65) & (!sk[101]) & (!g) & (!g96)) + ((!l) & (g65) & (!sk[101]) & (g) & (!g96)) + ((l) & (g65) & (!sk[101]) & (!g) & (g96)));
	assign g100 = (((n) & (!g51) & (!sk[102]) & (!g92) & (!g93) & (!g99)) + ((!n) & (!g51) & (!sk[102]) & (g92) & (!g93) & (!g99)) + ((!n) & (!g51) & (!sk[102]) & (!g92) & (g93) & (!g99)) + ((!n) & (!g51) & (sk[102]) & (!g92) & (!g93) & (!g99)) + ((!n) & (!g51) & (sk[102]) & (!g92) & (!g93) & (!g99)) + ((!n) & (!g51) & (sk[102]) & (!g92) & (!g93) & (!g99)) + ((!n) & (!g51) & (sk[102]) & (!g92) & (!g93) & (!g99)));
	assign g101 = (((k) & (!g26) & (!c) & (!g91) & (!sk[103]) & (!g100)) + ((!k) & (!g26) & (c) & (!g91) & (!sk[103]) & (!g100)) + ((!k) & (!g26) & (!c) & (g91) & (!sk[103]) & (!g100)) + ((!k) & (!g26) & (!c) & (!g91) & (sk[103]) & (!g100)) + ((k) & (g26) & (!c) & (g91) & (!sk[103]) & (!g100)));
	assign g102 = (((!g15) & (!c) & (!sk[104]) & (g)) + ((g15) & (c) & (!sk[104]) & (!g)) + ((g15) & (c) & (!sk[104]) & (g)));
	assign g103 = (((!g7) & (!sk[105]) & (!g90) & (g102)) + ((g7) & (!sk[105]) & (g90) & (!g102)) + ((!g7) & (sk[105]) & (!g90) & (!g102)) + ((!g7) & (sk[105]) & (!g90) & (!g102)));
	assign g104 = (((!g182) & (!g7) & (!g16) & (g44) & (!g46) & (g47)) + ((g182) & (!g7) & (g16) & (g44) & (!g46) & (!g47)) + ((!g182) & (g7) & (!g16) & (g44) & (g46) & (!g47)) + ((g182) & (!g7) & (g16) & (!g44) & (!g46) & (g47)) + ((g182) & (g7) & (g16) & (!g44) & (g46) & (!g47)));
	assign g105 = (((!k) & (g28) & (g) & (!g93) & (!g103) & (!g104)) + ((k) & (g28) & (!g) & (g93) & (g103) & (g104)) + ((k) & (g28) & (!g) & (!g93) & (!g103) & (g104)) + ((k) & (g28) & (!g) & (!g93) & (g103) & (!g104)) + ((k) & (g28) & (!g) & (g93) & (!g103) & (!g104)));
	assign g106 = (((!sk[108]) & (!g7) & (!g67) & (g46) & (!g47)) + ((!sk[108]) & (!g7) & (!g67) & (!g46) & (g47)) + ((!sk[108]) & (g7) & (g67) & (!g46) & (!g47)) + ((sk[108]) & (!g7) & (!g67) & (!g46) & (!g47)) + ((!sk[108]) & (!g7) & (!g67) & (g46) & (!g47)));
	assign g107 = (((!g68) & (!g90) & (g103) & (!sk[109]) & (!g106)) + ((!g68) & (!g90) & (!g103) & (!sk[109]) & (g106)) + ((g68) & (g90) & (!g103) & (!sk[109]) & (!g106)) + ((g68) & (g90) & (!g103) & (!sk[109]) & (g106)) + ((g68) & (!g90) & (!g103) & (sk[109]) & (!g106)));
	assign g108 = (((l) & (!a) & (!b) & (!sk[110]) & (!g60) & (!c)) + ((!l) & (!a) & (b) & (!sk[110]) & (!g60) & (!c)) + ((!l) & (!a) & (!b) & (!sk[110]) & (g60) & (!c)) + ((l) & (!a) & (!b) & (!sk[110]) & (g60) & (!c)));
	assign g109 = (((!g27) & (!sk[111]) & (!g62) & (g93)) + ((g27) & (!sk[111]) & (g62) & (!g93)) + ((g27) & (!sk[111]) & (g62) & (g93)));
	assign g110 = (((l) & (!g14) & (!g46) & (!sk[112]) & (!g60) & (!g90)) + ((!l) & (!g14) & (g46) & (!sk[112]) & (!g60) & (!g90)) + ((!l) & (!g14) & (!g46) & (!sk[112]) & (g60) & (!g90)) + ((!l) & (!g14) & (!g46) & (!sk[112]) & (g60) & (!g90)) + ((!l) & (!g14) & (!g46) & (!sk[112]) & (g60) & (!g90)) + ((!l) & (g14) & (g46) & (!sk[112]) & (g60) & (g90)));
	assign g111 = (((!g182) & (!g44) & (g54) & (!sk[113]) & (!g55)) + ((!g182) & (!g44) & (!g54) & (!sk[113]) & (g55)) + ((!g182) & (!g44) & (!g54) & (sk[113]) & (!g55)) + ((!g182) & (!g44) & (!g54) & (!sk[113]) & (g55)) + ((g182) & (g44) & (!g54) & (!sk[113]) & (!g55)));
	assign g112 = (((!sk[114]) & (g51) & (!g53) & (!c) & (!g92) & (!g111)) + ((!sk[114]) & (!g51) & (!g53) & (c) & (!g92) & (!g111)) + ((!sk[114]) & (!g51) & (!g53) & (!c) & (g92) & (!g111)) + ((!sk[114]) & (!g51) & (!g53) & (!c) & (g92) & (g111)) + ((!sk[114]) & (!g51) & (!g53) & (c) & (!g92) & (g111)) + ((!sk[114]) & (!g51) & (!g53) & (!c) & (g92) & (g111)) + ((sk[114]) & (!g51) & (!g53) & (!c) & (!g92) & (g111)));
	assign g113 = (((!n) & (!g93) & (!g108) & (!g109) & (!g110) & (!g112)) + ((!n) & (g93) & (!g108) & (!g109) & (!g110) & (!g112)) + ((!n) & (!g93) & (!g108) & (!g109) & (!g110) & (g112)));
	assign g114 = (((!g68) & (!g90) & (g103) & (!sk[116]) & (!g106)) + ((!g68) & (!g90) & (!g103) & (!sk[116]) & (g106)) + ((g68) & (g90) & (!g103) & (!sk[116]) & (!g106)) + ((g68) & (!g90) & (g103) & (!sk[116]) & (g106)) + ((g68) & (g90) & (g103) & (!sk[116]) & (!g106)));
	assign g115 = (((g98) & (!g101) & (!g105) & (!g107) & (!g113) & (!g114)) + ((!g98) & (g101) & (!g105) & (!g107) & (!g113) & (!g114)) + ((!g98) & (!g101) & (g105) & (!g107) & (!g113) & (!g114)) + ((!g98) & (!g101) & (!g105) & (g107) & (!g113) & (!g114)) + ((!g98) & (!g101) & (!g105) & (!g107) & (!g113) & (!g114)) + ((!g98) & (!g101) & (!g105) & (!g107) & (!g113) & (g114)));
	assign g116 = (((!k) & (l) & (!i) & (c) & (!g) & (!g93)) + ((k) & (!l) & (!i) & (!c) & (!g) & (g93)) + ((k) & (l) & (!i) & (!c) & (!g) & (!g93)) + ((!k) & (!l) & (!i) & (!c) & (!g) & (!g93)) + ((!k) & (!l) & (i) & (!c) & (!g) & (g93)) + ((k) & (!l) & (i) & (!c) & (!g) & (!g93)) + ((!k) & (l) & (i) & (!c) & (g) & (!g93)));
	assign g117 = (((!k) & (l) & (!i) & (!c) & (g) & (!g93)) + ((k) & (!l) & (i) & (c) & (!g) & (!g93)) + ((k) & (!l) & (!i) & (!c) & (!g) & (!g93)));
	assign g118 = (((g34) & (!g32) & (!sk[120]) & (c) & (!g93)) + ((!g34) & (!g32) & (!sk[120]) & (c) & (!g93)) + ((!g34) & (!g32) & (!sk[120]) & (!c) & (g93)) + ((!g34) & (g32) & (sk[120]) & (!c) & (!g93)) + ((g34) & (g32) & (!sk[120]) & (!c) & (!g93)));
	assign g119 = (((!sk[121]) & (g33) & (!g35) & (!c) & (!g) & (!g118)) + ((!sk[121]) & (!g33) & (!g35) & (c) & (!g) & (!g118)) + ((!sk[121]) & (!g33) & (g35) & (c) & (!g) & (!g118)) + ((!sk[121]) & (!g33) & (!g35) & (!c) & (g) & (!g118)) + ((!sk[121]) & (!g33) & (!g35) & (!c) & (g) & (g118)));
	assign g120 = (((!sk[122]) & (!g14) & (!g46) & (g90)) + ((!sk[122]) & (g14) & (g46) & (!g90)) + ((!sk[122]) & (g14) & (g46) & (g90)));
	assign g121 = (((!sk[123]) & (d) & (!h)) + ((!sk[123]) & (d) & (h)));
	assign g122 = (((!c) & (!sk[124]) & (!g) & (g81)) + ((!c) & (!sk[124]) & (!g) & (g81)) + ((!c) & (!sk[124]) & (g) & (g81)) + ((!c) & (sk[124]) & (g) & (!g81)) + ((c) & (!sk[124]) & (g) & (!g81)));
	assign g123 = (((!sk[125]) & (k) & (!l) & (!i) & (!j) & (!g122)) + ((!sk[125]) & (!k) & (!l) & (i) & (!j) & (!g122)) + ((!sk[125]) & (!k) & (!l) & (!i) & (j) & (!g122)) + ((!sk[125]) & (k) & (!l) & (!i) & (!j) & (!g122)) + ((!sk[125]) & (!k) & (l) & (i) & (j) & (!g122)) + ((!sk[125]) & (k) & (!l) & (!i) & (!j) & (g122)) + ((sk[125]) & (!k) & (l) & (!i) & (!j) & (!g122)));
	assign g124 = (((!sk[126]) & (!n) & (!g121) & (g123)) + ((!sk[126]) & (n) & (g121) & (!g123)) + ((!sk[126]) & (n) & (g121) & (g123)));
	assign g125 = (((!n) & (!j) & (!sk[127]) & (h)) + ((n) & (j) & (!sk[127]) & (!h)));
	assign g126 = (((!k) & (!l) & (!sk[0]) & (n) & (!j)) + ((!k) & (!l) & (!sk[0]) & (!n) & (j)) + ((k) & (l) & (!sk[0]) & (!n) & (!j)) + ((!k) & (!l) & (sk[0]) & (!n) & (!j)) + ((!k) & (!l) & (!sk[0]) & (!n) & (j)));
	assign g127 = (((i) & (!d) & (!g122) & (!g125) & (!sk[1]) & (!g126)) + ((!i) & (!d) & (g122) & (!g125) & (!sk[1]) & (!g126)) + ((!i) & (!d) & (!g122) & (g125) & (!sk[1]) & (!g126)) + ((!i) & (!d) & (g122) & (g125) & (!sk[1]) & (!g126)) + ((!i) & (!d) & (!g122) & (!g125) & (sk[1]) & (g126)));
	assign g128 = (((!sk[2]) & (!g1) & (!d) & (h)) + ((!sk[2]) & (g1) & (!d) & (h)) + ((sk[2]) & (!g1) & (d) & (!h)) + ((!sk[2]) & (g1) & (d) & (!h)));
	assign g129 = (((k) & (!sk[3]) & (!l) & (!n) & (!c) & (!g121)) + ((!k) & (!sk[3]) & (!l) & (n) & (!c) & (!g121)) + ((!k) & (!sk[3]) & (!l) & (!n) & (c) & (!g121)) + ((k) & (!sk[3]) & (!l) & (!n) & (!c) & (g121)) + ((k) & (!sk[3]) & (l) & (n) & (c) & (!g121)));
	assign g130 = (((!g2) & (!g4) & (!sk[4]) & (d) & (!h)) + ((!g2) & (!g4) & (!sk[4]) & (!d) & (h)) + ((!g2) & (!g4) & (!sk[4]) & (!d) & (h)) + ((g2) & (g4) & (!sk[4]) & (!d) & (!h)) + ((!g2) & (!g4) & (sk[4]) & (!d) & (!h)) + ((!g2) & (!g4) & (!sk[4]) & (d) & (!h)));
	assign g131 = (((!i) & (!j) & (!sk[5]) & (g129) & (!g130)) + ((i) & (!j) & (!sk[5]) & (!g129) & (g130)) + ((!i) & (j) & (!sk[5]) & (!g129) & (g130)) + ((!i) & (!j) & (!sk[5]) & (!g129) & (g130)) + ((i) & (j) & (!sk[5]) & (!g129) & (!g130)));
	assign g132 = (((g11) & (!g122) & (!g127) & (!g128) & (!sk[6]) & (!g131)) + ((!g11) & (!g122) & (g127) & (!g128) & (!sk[6]) & (!g131)) + ((!g11) & (!g122) & (!g127) & (g128) & (!sk[6]) & (!g131)) + ((!g11) & (!g122) & (!g127) & (!g128) & (sk[6]) & (g131)) + ((!g11) & (g122) & (!g127) & (!g128) & (sk[6]) & (g131)) + ((!g11) & (!g122) & (!g127) & (!g128) & (sk[6]) & (g131)));
	assign g133 = (((!g9) & (!g12) & (!sk[7]) & (d)) + ((g9) & (g12) & (!sk[7]) & (!d)) + ((!g9) & (!g12) & (sk[7]) & (!d)) + ((!g9) & (!g12) & (!sk[7]) & (d)));
	assign g134 = (((!g7) & (g12) & (!sk[8]) & (d) & (!h)) + ((!g7) & (!g12) & (!sk[8]) & (d) & (!h)) + ((!g7) & (!g12) & (!sk[8]) & (!d) & (h)) + ((g7) & (g12) & (!sk[8]) & (!d) & (!h)) + ((g7) & (!g12) & (!sk[8]) & (d) & (h)));
	assign g135 = (((g10) & (!g124) & (!sk[9]) & (!g132) & (!g133) & (!g134)) + ((!g10) & (!g124) & (!sk[9]) & (g132) & (!g133) & (!g134)) + ((!g10) & (!g124) & (!sk[9]) & (!g132) & (g133) & (!g134)) + ((!g10) & (g124) & (!sk[9]) & (!g132) & (g133) & (!g134)) + ((!g10) & (!g124) & (!sk[9]) & (!g132) & (g133) & (!g134)) + ((!g10) & (!g124) & (!sk[9]) & (g132) & (!g133) & (!g134)));
	assign g136 = (((!a) & (!b) & (c) & (!sk[10]) & (!d)) + ((a) & (!b) & (!c) & (!sk[10]) & (d)) + ((!a) & (b) & (!c) & (!sk[10]) & (d)) + ((!a) & (!b) & (c) & (!sk[10]) & (d)) + ((!a) & (!b) & (!c) & (!sk[10]) & (d)) + ((a) & (b) & (!c) & (!sk[10]) & (!d)) + ((!a) & (!b) & (!c) & (sk[10]) & (!d)));
	assign g137 = (((l) & (!g60) & (!g120) & (!g135) & (!sk[11]) & (!g136)) + ((!l) & (!g60) & (g120) & (!g135) & (!sk[11]) & (!g136)) + ((!l) & (!g60) & (!g120) & (g135) & (!sk[11]) & (!g136)) + ((l) & (g60) & (!g120) & (!g135) & (!sk[11]) & (g136)) + ((!l) & (g60) & (g120) & (g135) & (!sk[11]) & (!g136)) + ((!l) & (g60) & (!g120) & (!g135) & (sk[11]) & (!g136)));
	assign g138 = (((!g7) & (g15) & (!sk[12]) & (g121) & (!g135)) + ((!g7) & (!g15) & (!sk[12]) & (g121) & (!g135)) + ((g7) & (!g15) & (!sk[12]) & (!g121) & (g135)) + ((!g7) & (!g15) & (!sk[12]) & (!g121) & (g135)) + ((g7) & (g15) & (!sk[12]) & (!g121) & (!g135)));
	assign g139 = (((!g7) & (!g67) & (g46) & (!g47) & (g90) & (!g102)) + ((!g7) & (!g67) & (!g46) & (!g47) & (g90) & (!g102)) + ((!g7) & (!g67) & (g46) & (!g47) & (!g90) & (!g102)) + ((!g7) & (!g67) & (!g46) & (!g47) & (!g90) & (!g102)) + ((!g7) & (!g67) & (!g46) & (!g47) & (g90) & (!g102)) + ((!g7) & (!g67) & (g46) & (!g47) & (g90) & (!g102)) + ((!g7) & (!g67) & (g46) & (!g47) & (!g90) & (!g102)));
	assign g140 = (((n) & (!sk[14]) & (!g18) & (!g135) & (!g138) & (!g139)) + ((!n) & (!sk[14]) & (!g18) & (g135) & (!g138) & (!g139)) + ((!n) & (!sk[14]) & (!g18) & (!g135) & (g138) & (!g139)) + ((n) & (!sk[14]) & (g18) & (g135) & (g138) & (g139)) + ((n) & (!sk[14]) & (g18) & (!g135) & (!g138) & (g139)) + ((n) & (!sk[14]) & (g18) & (!g135) & (g138) & (!g139)) + ((n) & (!sk[14]) & (g18) & (g135) & (!g138) & (!g139)));
	assign g141 = (((g124) & (!sk[15]) & (!g132)) + ((!g124) & (sk[15]) & (g132)));
	assign g142 = (((g7) & (g93) & (g103) & (!g104) & (g141) & (g138)) + ((g7) & (g93) & (!g103) & (!g104) & (g141) & (g138)) + ((g7) & (!g93) & (g103) & (!g104) & (g141) & (g138)) + ((g7) & (g93) & (g103) & (!g104) & (!g141) & (!g138)) + ((g7) & (g93) & (!g103) & (!g104) & (!g141) & (!g138)) + ((g7) & (!g93) & (g103) & (!g104) & (!g141) & (!g138)));
	assign g143 = (((g7) & (!g93) & (!g103) & (!g104) & (!g141) & (g138)) + ((g7) & (!g93) & (!g103) & (g104) & (!g141) & (g138)) + ((g7) & (!g93) & (!g103) & (g104) & (!g141) & (g138)) + ((g7) & (!g93) & (!g103) & (!g104) & (g141) & (!g138)) + ((g7) & (!g93) & (!g103) & (g104) & (g141) & (!g138)) + ((g7) & (!g93) & (!g103) & (g104) & (g141) & (!g138)));
	assign g144 = (((!g53) & (!g57) & (!c) & (!g92) & (!g93) & (!g141)) + ((!g53) & (!g57) & (c) & (g92) & (!g93) & (g141)) + ((!g53) & (!g57) & (c) & (!g92) & (!g93) & (g141)) + ((!g53) & (!g57) & (!c) & (g92) & (!g93) & (g141)) + ((!g53) & (!g57) & (!c) & (!g92) & (!g93) & (!g141)) + ((!g53) & (!g57) & (!c) & (!g92) & (g93) & (!g141)) + ((!g53) & (!g57) & (!c) & (!g92) & (g93) & (!g141)));
	assign g145 = (((n) & (!sk[19]) & (!d)) + ((n) & (!sk[19]) & (d)));
	assign g146 = (((n) & (!g62) & (g54) & (!g55) & (!g93) & (!g141)) + ((n) & (!g62) & (!g54) & (g55) & (!g93) & (!g141)) + ((n) & (!g62) & (!g54) & (g55) & (!g93) & (!g141)));
	assign g147 = (((!sk[21]) & (c) & (g) & (!g96)) + ((!sk[21]) & (!c) & (!g) & (g96)) + ((!sk[21]) & (c) & (!g) & (g96)) + ((!sk[21]) & (!c) & (g) & (g96)));
	assign g148 = (((l) & (!g65) & (!d) & (!h) & (!sk[22]) & (!g147)) + ((!l) & (!g65) & (d) & (!h) & (!sk[22]) & (!g147)) + ((!l) & (!g65) & (!d) & (h) & (!sk[22]) & (!g147)) + ((!l) & (g65) & (!d) & (h) & (!sk[22]) & (!g147)) + ((!l) & (g65) & (d) & (h) & (!sk[22]) & (g147)) + ((!l) & (g65) & (!d) & (h) & (!sk[22]) & (!g147)) + ((!l) & (g65) & (d) & (!h) & (!sk[22]) & (!g147)) + ((l) & (g65) & (!d) & (!h) & (!sk[22]) & (g147)));
	assign g149 = (((!sk[23]) & (!n) & (!g51) & (d)) + ((!sk[23]) & (n) & (g51) & (!d)));
	assign g150 = (((!c) & (!g92) & (!g93) & (!g141) & (!g148) & (!g149)) + ((!c) & (!g92) & (!g93) & (g141) & (!g148) & (!g149)) + ((!c) & (!g92) & (g93) & (g141) & (!g148) & (!g149)) + ((!c) & (!g92) & (g93) & (g141) & (!g148) & (!g149)) + ((c) & (g92) & (!g93) & (!g141) & (!g148) & (!g149)) + ((c) & (!g92) & (!g93) & (!g141) & (!g148) & (!g149)) + ((!c) & (g92) & (!g93) & (!g141) & (!g148) & (!g149)));
	assign g151 = (((!g109) & (!g141) & (g144) & (!g145) & (!g146) & (g150)) + ((!g109) & (!g141) & (g144) & (!g145) & (!g146) & (g150)) + ((!g109) & (!g141) & (!g144) & (!g145) & (!g146) & (g150)) + ((!g109) & (!g141) & (!g144) & (!g145) & (!g146) & (g150)));
	assign g152 = (((!a) & (!g14) & (!b) & (!g46) & (c) & (!g90)) + ((!a) & (!g14) & (b) & (!g46) & (c) & (!g90)) + ((!a) & (!g14) & (b) & (!g46) & (!c) & (!g90)) + ((a) & (!g14) & (b) & (!g46) & (c) & (!g90)) + ((a) & (!g14) & (!b) & (!g46) & (c) & (!g90)) + ((a) & (!g14) & (b) & (!g46) & (!c) & (!g90)) + ((a) & (!g14) & (!b) & (!g46) & (!c) & (!g90)));
	assign g153 = (((!sk[27]) & (!l) & (!i) & (j) & (!d)) + ((!sk[27]) & (!l) & (!i) & (!j) & (d)) + ((!sk[27]) & (l) & (i) & (!j) & (!d)) + ((!sk[27]) & (!l) & (!i) & (!j) & (d)));
	assign g154 = (((!i) & (!j) & (!sk[28]) & (g1) & (!d)) + ((!i) & (!j) & (!sk[28]) & (!g1) & (d)) + ((i) & (j) & (!sk[28]) & (!g1) & (!d)) + ((!i) & (!j) & (!sk[28]) & (g1) & (!d)));
	assign g155 = (((!sk[29]) & (n) & (!g135) & (!g152) & (!g153) & (!g154)) + ((!sk[29]) & (!n) & (!g135) & (g152) & (!g153) & (!g154)) + ((!sk[29]) & (!n) & (!g135) & (!g152) & (g153) & (!g154)) + ((!sk[29]) & (n) & (!g135) & (g152) & (g153) & (!g154)) + ((!sk[29]) & (n) & (g135) & (!g152) & (g153) & (!g154)) + ((!sk[29]) & (n) & (g135) & (g152) & (!g153) & (g154)) + ((!sk[29]) & (n) & (!g135) & (!g152) & (!g153) & (g154)));
	assign g156 = (((!g137) & (!g140) & (!g142) & (!g143) & (g151) & (!g155)));
	assign g157 = (((!k) & (!l) & (!i) & (!d) & (!h) & (g141)) + ((!k) & (!l) & (i) & (!d) & (!h) & (!g141)) + ((k) & (!l) & (!i) & (!d) & (!h) & (!g141)) + ((k) & (!l) & (i) & (!d) & (h) & (!g141)) + ((!k) & (!l) & (!i) & (!d) & (!h) & (g141)) + ((k) & (!l) & (i) & (!d) & (h) & (g141)) + ((!k) & (!l) & (!i) & (!d) & (h) & (g141)) + ((!k) & (l) & (i) & (d) & (h) & (!g141)) + ((!k) & (l) & (i) & (!d) & (!h) & (!g141)) + ((k) & (l) & (i) & (!d) & (!h) & (g141)));
	assign g158 = (((!k) & (l) & (!i) & (!d) & (h) & (!g141)) + ((k) & (!l) & (i) & (d) & (!h) & (!g141)) + ((k) & (!l) & (!i) & (!d) & (!h) & (!g141)));
	assign g159 = (((g33) & (!g34) & (!g35) & (!sk[33]) & (!d) & (!h)) + ((!g33) & (!g34) & (!g35) & (!sk[33]) & (d) & (!h)) + ((!g33) & (!g34) & (!g35) & (sk[33]) & (!d) & (!h)) + ((!g33) & (!g34) & (g35) & (!sk[33]) & (!d) & (!h)) + ((!g33) & (!g34) & (!g35) & (!sk[33]) & (d) & (!h)) + ((!g33) & (!g34) & (!g35) & (!sk[33]) & (d) & (!h)));
	assign g160 = (((!sk[34]) & (!g32) & (!h) & (g141) & (!g159)) + ((!sk[34]) & (!g32) & (!h) & (!g141) & (g159)) + ((!sk[34]) & (!g32) & (!h) & (!g141) & (g159)) + ((!sk[34]) & (!g32) & (!h) & (g141) & (g159)) + ((!sk[34]) & (g32) & (h) & (!g141) & (!g159)));
	assign g161 = (((n) & (!sk[35]) & (!j) & (!g157) & (!g158) & (!g160)) + ((!n) & (!sk[35]) & (!j) & (g157) & (!g158) & (!g160)) + ((!n) & (!sk[35]) & (!j) & (!g157) & (g158) & (!g160)) + ((n) & (!sk[35]) & (!j) & (!g157) & (!g158) & (g160)) + ((!n) & (!sk[35]) & (!j) & (g157) & (!g158) & (g160)) + ((!n) & (sk[35]) & (j) & (!g157) & (!g158) & (g160)));
	assign r = (((!n) & (!sk[36]) & (!g80) & (g115) & (!g156) & (!g161)) + ((!n) & (!sk[36]) & (!g80) & (!g115) & (g156) & (!g161)) + ((!n) & (sk[36]) & (!g80) & (!g115) & (!g156) & (!g161)) + ((n) & (!sk[36]) & (g80) & (!g115) & (!g156) & (!g161)) + ((n) & (!sk[36]) & (!g80) & (!g115) & (!g156) & (!g161)) + ((n) & (!sk[36]) & (!g80) & (g115) & (g156) & (!g161)));
	assign g163 = (((d) & (!sk[37]) & (!h)) + ((d) & (!sk[37]) & (!h)) + ((!d) & (sk[37]) & (h)));
	assign g164 = (((k) & (!l) & (!sk[38]) & (!g8) & (!g120) & (!g135)) + ((!k) & (!l) & (!sk[38]) & (g8) & (!g120) & (!g135)) + ((!k) & (!l) & (!sk[38]) & (!g8) & (g120) & (!g135)) + ((!k) & (!l) & (!sk[38]) & (g8) & (!g120) & (!g135)) + ((!k) & (!l) & (!sk[38]) & (g8) & (g120) & (g135)));
	assign g165 = (((!i) & (!sk[39]) & (!d) & (g135) & (!g152)) + ((!i) & (!sk[39]) & (!d) & (!g135) & (g152)) + ((i) & (!sk[39]) & (d) & (!g135) & (!g152)) + ((!i) & (!sk[39]) & (d) & (!g135) & (g152)) + ((!i) & (sk[39]) & (d) & (!g135) & (!g152)));
	assign g166 = (((i) & (!g93) & (!g103) & (!g104) & (!g141) & (!g138)) + ((i) & (!g93) & (!g103) & (g104) & (!g141) & (!g138)) + ((i) & (!g93) & (!g103) & (g104) & (!g141) & (!g138)) + ((i) & (!g93) & (!g103) & (!g104) & (!g141) & (g138)) + ((i) & (!g93) & (!g103) & (g104) & (!g141) & (g138)) + ((i) & (!g93) & (!g103) & (g104) & (!g141) & (g138)));
	assign g167 = (((i) & (!sk[41]) & (!g141) & (!g135) & (!g138) & (!g152)) + ((!i) & (!sk[41]) & (!g141) & (g135) & (!g138) & (!g152)) + ((!i) & (!sk[41]) & (!g141) & (!g135) & (g138) & (!g152)) + ((i) & (!sk[41]) & (!g141) & (!g135) & (g138) & (!g152)) + ((!i) & (sk[41]) & (!g141) & (!g135) & (!g138) & (g152)));
	assign g168 = (((!k) & (!sk[42]) & (!i) & (j)) + ((!k) & (sk[42]) & (!i) & (!j)) + ((k) & (!sk[42]) & (!i) & (j)) + ((k) & (!sk[42]) & (i) & (!j)));
	assign g169 = (((!c) & (!g92) & (!g93) & (d) & (!g141) & (g168)) + ((c) & (g92) & (!g93) & (d) & (!g141) & (g168)) + ((c) & (!g92) & (!g93) & (d) & (!g141) & (g168)) + ((!c) & (g92) & (!g93) & (d) & (!g141) & (g168)) + ((c) & (g92) & (!g93) & (!d) & (!g141) & (g168)) + ((c) & (!g92) & (!g93) & (!d) & (!g141) & (g168)) + ((!c) & (g92) & (!g93) & (!d) & (!g141) & (g168)));
	assign g170 = (((g7) & (!g15) & (g17) & (!sk[44]) & (!g121) & (!g135)) + ((g7) & (!g15) & (!g17) & (!sk[44]) & (!g121) & (!g135)) + ((!g7) & (!g15) & (g17) & (!sk[44]) & (!g121) & (!g135)) + ((!g7) & (!g15) & (!g17) & (!sk[44]) & (g121) & (!g135)) + ((!g7) & (!g15) & (g17) & (!sk[44]) & (!g121) & (!g135)) + ((!g7) & (g15) & (g17) & (!sk[44]) & (g121) & (!g135)));
	assign g171 = (((!sk[45]) & (!a) & (!b) & (c) & (!d)) + ((!sk[45]) & (!a) & (!b) & (!c) & (d)) + ((!sk[45]) & (a) & (b) & (!c) & (!d)) + ((sk[45]) & (!a) & (!b) & (!c) & (!d)));
	assign g172 = (((!k) & (!g8) & (!sk[46]) & (g171) & (!g183)) + ((!k) & (!g8) & (!sk[46]) & (!g171) & (g183)) + ((!k) & (!g8) & (!sk[46]) & (!g171) & (g183)) + ((k) & (g8) & (!sk[46]) & (!g171) & (!g183)) + ((k) & (g8) & (!sk[46]) & (g171) & (!g183)));
	assign g173 = (((!sk[47]) & (!k) & (!l) & (i) & (!j)) + ((!sk[47]) & (!k) & (!l) & (!i) & (j)) + ((!sk[47]) & (k) & (l) & (!i) & (!j)) + ((!sk[47]) & (!k) & (!l) & (i) & (j)) + ((!sk[47]) & (k) & (!l) & (!i) & (j)));
	assign g174 = (((!g62) & (!g93) & (!sk[48]) & (g141) & (!g173)) + ((!g62) & (!g93) & (!sk[48]) & (!g141) & (g173)) + ((g62) & (g93) & (!sk[48]) & (!g141) & (!g173)) + ((g62) & (g93) & (!sk[48]) & (g141) & (g173)));
	assign g175 = (((!l) & (!g139) & (!g169) & (!g170) & (!g172) & (!g174)) + ((!l) & (g139) & (!g169) & (!g170) & (!g172) & (!g174)) + ((!l) & (!g139) & (!g169) & (!g170) & (!g172) & (!g174)));
	assign g176 = (((j) & (!g1) & (!g165) & (!g166) & (!g167) & (g175)) + ((!j) & (!g1) & (!g165) & (!g166) & (!g167) & (g175)) + ((!j) & (!g1) & (!g165) & (!g166) & (!g167) & (g175)));
	assign u = (((n) & (!g80) & (!g115) & (!g156) & (g164) & (!g176)) + ((n) & (!g80) & (!g115) & (!g156) & (!g164) & (!g176)) + ((n) & (!g80) & (g115) & (!g156) & (!g164) & (!g176)));
	assign g178 = (((!a) & (!e) & (!sk[52]) & (g163)) + ((a) & (e) & (!sk[52]) & (!g163)) + ((!a) & (!e) & (sk[52]) & (!g163)));
	assign g179 = (((f) & (!b) & (!c) & (!sk[53]) & (!g) & (!g178)) + ((f) & (!b) & (!c) & (!sk[53]) & (!g) & (!g178)) + ((!f) & (!b) & (!c) & (!sk[53]) & (g) & (!g178)) + ((!f) & (!b) & (c) & (!sk[53]) & (!g) & (!g178)) + ((!f) & (!b) & (!c) & (sk[53]) & (!g) & (!g178)) + ((!f) & (b) & (!c) & (sk[53]) & (!g) & (!g178)) + ((!f) & (!b) & (!c) & (!sk[53]) & (g) & (!g178)));
	assign g180 = (((l) & (!k) & (!e) & (!a) & (j) & (n)) + ((!l) & (!k) & (!e) & (a) & (j) & (n)) + ((!l) & (!k) & (!e) & (!a) & (!j) & (!n)) + ((!l) & (!k) & (!e) & (!a) & (!j) & (!n)) + ((!l) & (k) & (e) & (a) & (!j) & (!n)) + ((!l) & (k) & (e) & (!a) & (j) & (n)) + ((l) & (!k) & (e) & (a) & (!j) & (n)) + ((!l) & (!k) & (!e) & (!a) & (j) & (!n)));
	assign g181 = (((!l) & (k) & (!e) & (!a) & (j) & (!n)) + ((!l) & (k) & (e) & (!a) & (!j) & (n)) + ((!l) & (!k) & (e) & (!a) & (!j) & (!n)) + ((l) & (k) & (!e) & (!a) & (!j) & (!n)) + ((!l) & (!k) & (!e) & (a) & (!j) & (!n)) + ((l) & (!k) & (e) & (a) & (j) & (n)) + ((!l) & (k) & (!e) & (a) & (!j) & (n)));
	assign g182 = (((g180) & (g181) & (!sk[56]) & (!i)) + ((!g180) & (g181) & (!sk[56]) & (i)) + ((!g180) & (!g181) & (!sk[56]) & (i)) + ((g180) & (!g181) & (sk[56]) & (!i)));
	assign g183 = (((g184) & (!sk[57]) & (!g185)) + ((!g184) & (sk[57]) & (!g185)));
	assign g184 = (((k) & (!sk[58]) & (!g186)) + ((!k) & (sk[58]) & (g186)));
	assign g185 = (((k) & (!sk[59]) & (!g189)) + ((k) & (!sk[59]) & (g189)));
	assign g186 = (((g187) & (!sk[60]) & (!g188)) + ((!g187) & (sk[60]) & (!g188)));
	assign g187 = (((!sk[61]) & (j) & (!g190)) + ((sk[61]) & (!j) & (g190)));
	assign g188 = (((j) & (!sk[62]) & (!g191)) + ((j) & (!sk[62]) & (g191)));
	assign g189 = (((!sk[63]) & (j) & (!g192)) + ((sk[63]) & (!j) & (g192)));
	assign g190 = (((!sk[64]) & (!h) & (!d) & (g147) & (!i)) + ((!sk[64]) & (!h) & (!d) & (!g147) & (i)) + ((!sk[64]) & (h) & (d) & (!g147) & (!i)) + ((!sk[64]) & (h) & (d) & (!g147) & (i)) + ((!sk[64]) & (h) & (!d) & (g147) & (i)) + ((!sk[64]) & (!h) & (d) & (g147) & (i)));
	assign g191 = (((!h) & (!sk[65]) & (!d) & (g12) & (!i)) + ((!h) & (!sk[65]) & (!d) & (!g12) & (i)) + ((h) & (!sk[65]) & (d) & (!g12) & (!i)) + ((h) & (!sk[65]) & (d) & (g12) & (!i)));
	assign g192 = (((!h) & (!d) & (!sk[66]) & (g147) & (!i)) + ((!h) & (!d) & (!sk[66]) & (!g147) & (i)) + ((h) & (d) & (!sk[66]) & (!g147) & (!i)) + ((h) & (d) & (!sk[66]) & (!g147) & (i)) + ((h) & (!d) & (!sk[66]) & (g147) & (i)) + ((!h) & (d) & (!sk[66]) & (g147) & (i)));
	assign q = (((!sk[67]) & (g194) & (!g195)) + ((sk[67]) & (!g194) & (!g195)));
	assign g194 = (((!sk[68]) & (n) & (!g196)) + ((sk[68]) & (!n) & (g196)));
	assign g195 = (((n) & (!sk[69]) & (!g199)) + ((n) & (!sk[69]) & (g199)));
	assign g196 = (((g197) & (!sk[70]) & (!g198)) + ((!g197) & (sk[70]) & (!g198)));
	assign g197 = (((!sk[71]) & (j) & (!g202)) + ((sk[71]) & (!j) & (g202)));
	assign g198 = (((!sk[72]) & (j) & (!g203)) + ((!sk[72]) & (j) & (g203)));
	assign g199 = (((!sk[73]) & (g200) & (!g201)) + ((sk[73]) & (!g200) & (!g201)));
	assign g200 = (((!sk[74]) & (j) & (!g204)) + ((sk[74]) & (!j) & (g204)));
	assign g201 = (((!sk[75]) & (j) & (!g205)) + ((!sk[75]) & (j) & (g205)));
	assign g202 = (((!sk[76]) & (g119) & (!g116)) + ((sk[76]) & (!g119) & (g116)));
	assign g203 = (((!sk[77]) & (g119) & (!g117)) + ((sk[77]) & (!g119) & (g117)));
	assign g204 = (((g119) & (g115) & (!sk[78]) & (!g80)) + ((!g119) & (g115) & (!sk[78]) & (g80)) + ((!g119) & (!g115) & (!sk[78]) & (g80)) + ((!g119) & (!g115) & (sk[78]) & (!g80)) + ((g119) & (!g115) & (!sk[78]) & (g80)));
	assign g205 = (((g119) & (!sk[79]) & (g115) & (!g80)) + ((!g119) & (!sk[79]) & (!g115) & (g80)) + ((!g119) & (!sk[79]) & (g115) & (g80)) + ((!g119) & (sk[79]) & (!g115) & (!g80)) + ((g119) & (!sk[79]) & (!g115) & (g80)));
	assign g206 = (((g207) & (!sk[80]) & (!g208)) + ((!g207) & (sk[80]) & (!g208)));
	assign g207 = (((!sk[81]) & (g50) & (!g209)) + ((sk[81]) & (!g50) & (g209)));
	assign g208 = (((!sk[82]) & (g50) & (!g212)) + ((!sk[82]) & (g50) & (g212)));
	assign g209 = (((!sk[83]) & (g210) & (!g211)) + ((sk[83]) & (!g210) & (!g211)));
	assign g210 = (((b) & (!sk[84]) & (!g215)) + ((!b) & (sk[84]) & (g215)));
	assign g211 = (((!sk[85]) & (b) & (!g216)) + ((!sk[85]) & (b) & (g216)));
	assign g212 = (((!sk[86]) & (g213) & (!g214)) + ((sk[86]) & (!g213) & (!g214)));
	assign g213 = (((!sk[87]) & (b) & (!g217)) + ((sk[87]) & (!b) & (g217)));
	assign g214 = (((!sk[88]) & (b) & (!g218)) + ((!sk[88]) & (b) & (g218)));
	assign g215 = (((g56) & (!sk[89]) & (!g51) & (g44)) + ((!g56) & (!sk[89]) & (!g51) & (g44)) + ((!g56) & (!sk[89]) & (g51) & (g44)) + ((g56) & (!sk[89]) & (g51) & (!g44)));
	assign g216 = (((sk[90]) & (!g56) & (g57) & (!g53) & (!g44)) + ((!sk[90]) & (g56) & (g57) & (!g53) & (!g44)) + ((!sk[90]) & (!g56) & (!g57) & (!g53) & (g44)) + ((!sk[90]) & (g56) & (!g57) & (!g53) & (g44)) + ((!sk[90]) & (!g56) & (!g57) & (g53) & (!g44)));
	assign g217 = (((g56) & (!sk[91]) & (!g44)) + ((g56) & (!sk[91]) & (g44)));
	assign g218 = (((sk[92]) & (!g56) & (g57) & (!g53) & (!g44)) + ((!sk[92]) & (g56) & (g57) & (!g53) & (!g44)) + ((!sk[92]) & (!g56) & (!g57) & (g53) & (!g44)) + ((!sk[92]) & (!g56) & (!g57) & (!g53) & (g44)) + ((!sk[92]) & (g56) & (!g57) & (!g53) & (g44)) + ((!sk[92]) & (!g56) & (!g57) & (g53) & (g44)));
	assign o = (((g220) & (!sk[93]) & (!g221)) + ((!g220) & (sk[93]) & (!g221)));
	assign g220 = (((!sk[94]) & (n) & (!g222)) + ((sk[94]) & (!n) & (g222)));
	assign g221 = (((!sk[95]) & (n) & (!g225)) + ((!sk[95]) & (n) & (g225)));
	assign g222 = (((!sk[96]) & (g223) & (!g224)) + ((sk[96]) & (!g223) & (!g224)));
	assign g223 = (((!sk[97]) & (j) & (!g228)) + ((sk[97]) & (!j) & (g228)));
	assign g224 = (((!sk[98]) & (j) & (!g229)) + ((!sk[98]) & (j) & (g229)));
	assign g225 = (((g226) & (!sk[99]) & (!g227)) + ((!g226) & (sk[99]) & (!g227)));
	assign g226 = (((!sk[100]) & (j) & (!g230)) + ((sk[100]) & (!j) & (g230)));
	assign g227 = (((j) & (!sk[101]) & (!g231)) + ((j) & (!sk[101]) & (g231)));
	assign g228 = (((!sk[102]) & (g37) & (!g5)) + ((sk[102]) & (!g37) & (g5)));
	assign g229 = (((g37) & (!sk[103]) & (!g6)) + ((!g37) & (sk[103]) & (g6)));
	assign g230 = (((g37) & (g31) & (!sk[104]) & (!m)) + ((!g37) & (g31) & (!sk[104]) & (m)) + ((!g37) & (!g31) & (!sk[104]) & (m)) + ((!g37) & (!g31) & (sk[104]) & (!m)) + ((g37) & (!g31) & (!sk[104]) & (m)));
	assign g231 = (((!sk[105]) & (g37) & (g31) & (!m)) + ((!sk[105]) & (!g37) & (!g31) & (m)) + ((!sk[105]) & (!g37) & (g31) & (m)) + ((sk[105]) & (!g37) & (!g31) & (!m)) + ((!sk[105]) & (g37) & (!g31) & (m)));

endmodule