module ex5px6xv (i_7_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_, o_1_, o_19_, o_2_, o_0_, o_29_, o_60_, o_39_, o_38_, o_25_, o_12_, o_37_, o_26_, o_11_, o_50_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_, o_34_, o_21_, o_16_, o_40_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_, o_31_, o_24_, o_17_, o_56_, o_43_, o_30_, o_55_, o_44_, o_58_, o_41_, o_57_, o_42_, o_20_, o_52_, o_47_, o_51_, o_48_, o_54_, o_45_, o_10_, o_53_, o_46_, o_61_, o_9_, o_62_, o_49_, o_7_, o_8_, o_5_, o_59_, o_6_, o_3_, o_4_);

	input i_7_;
	input i_5_;
	input i_6_;
	input i_3_;
	input i_4_;
	input i_1_;
	input i_2_;
	input i_0_;
	output o_1_;
	output o_19_;
	output o_2_;
	output o_0_;
	output o_29_;
	output o_60_;
	output o_39_;
	output o_38_;
	output o_25_;
	output o_12_;
	output o_37_;
	output o_26_;
	output o_11_;
	output o_50_;
	output o_36_;
	output o_27_;
	output o_14_;
	output o_35_;
	output o_28_;
	output o_13_;
	output o_34_;
	output o_21_;
	output o_16_;
	output o_40_;
	output o_33_;
	output o_22_;
	output o_15_;
	output o_32_;
	output o_23_;
	output o_18_;
	output o_31_;
	output o_24_;
	output o_17_;
	output o_56_;
	output o_43_;
	output o_30_;
	output o_55_;
	output o_44_;
	output o_58_;
	output o_41_;
	output o_57_;
	output o_42_;
	output o_20_;
	output o_52_;
	output o_47_;
	output o_51_;
	output o_48_;
	output o_54_;
	output o_45_;
	output o_10_;
	output o_53_;
	output o_46_;
	output o_61_;
	output o_9_;
	output o_62_;
	output o_49_;
	output o_7_;
	output o_8_;
	output o_5_;
	output o_59_;
	output o_6_;
	output o_3_;
	output o_4_;

	wire [127 : 0] sk /* synthesis noprune */;

	lut_sub lut_3 ({sk[0], i_7_, i_5_, i_6_}, o_1_);
	defparam lut_3.LUT_SIZE = 4;
	defparam lut_3.mask = 16'h5580;

	lut_sub lut_5 ({sk[1], i_7_, i_5_, i_6_, i_3_, i_4_, n_n0}, o_19_);
	defparam lut_5.LUT_SIZE = 7;
	defparam lut_5.mask = 128'h555f55ff5f5f5fff1010101010101010;

	lut_sub lut_14 ({sk[2], i_7_, i_6_, i_1_, i_2_, i_0_, n_n8}, o_2_);
	defparam lut_14.LUT_SIZE = 7;
	defparam lut_14.mask = 128'h555f55ff5f5f5fff5555000000000000;

	lut_sub lut_23 ({sk[3], i_5_, i_6_, i_3_, i_4_}, o_0_);
	defparam lut_23.LUT_SIZE = 5;
	defparam lut_23.mask = 32'h5757a000;

	lut_sub lut_26 ({sk[4], i_7_, i_5_, i_6_, i_3_, i_4_, n_n0}, o_29_);
	defparam lut_26.LUT_SIZE = 7;
	defparam lut_26.mask = 128'h555f55ff5f5f5fff0000000040000000;

	lut_sub lut_28 ({sk[5], i_3_, i_4_, x5121x, x5122x}, o_60_);
	defparam lut_28.LUT_SIZE = 5;
	defparam lut_28.mask = 32'h5757e7df;

	lut_sub lut_36 ({sk[6], i_7_, i_5_, i_6_, i_3_, i_4_, x5119x}, o_39_);
	defparam lut_36.LUT_SIZE = 7;
	defparam lut_36.mask = 128'h555f55ff5f5f5fffbbbbb3bbbbbbbbbb;

	lut_sub lut_43 ({sk[7], i_7_, i_6_, x5117x, x5118x}, o_38_);
	defparam lut_43.LUT_SIZE = 5;
	defparam lut_43.mask = 32'h57579a9b;

	lut_sub lut_48 ({sk[8], i_7_, i_6_, i_1_, i_2_, i_0_, n_n7}, o_25_);
	defparam lut_48.LUT_SIZE = 7;
	defparam lut_48.mask = 128'h555f55ff5f5f5fff0000004000000000;

	lut_sub lut_50 ({sk[9], i_1_, i_2_, i_0_, x82x}, o_12_);
	defparam lut_50.LUT_SIZE = 5;
	defparam lut_50.mask = 32'h57570100;

	lut_sub lut_52 ({sk[10], i_7_, i_5_, i_6_, i_3_, i_4_, x5115x}, o_37_);
	defparam lut_52.LUT_SIZE = 7;
	defparam lut_52.mask = 128'h555f55ff5f5f5fffaaa2aaaaaaaaaaaa;

	lut_sub lut_58 ({sk[11], i_1_, i_2_, i_0_, x121x}, o_26_);
	defparam lut_58.LUT_SIZE = 5;
	defparam lut_58.mask = 32'h57570101;

	lut_sub lut_61 ({sk[12], i_1_, i_2_, i_0_, x82x}, o_11_);
	defparam lut_61.LUT_SIZE = 5;
	defparam lut_61.mask = 32'h57570010;

	lut_sub lut_63 ({sk[13], i_7_, i_6_, x5114x}, o_50_);
	defparam lut_63.LUT_SIZE = 4;
	defparam lut_63.mask = 16'h55fe;

	lut_sub lut_67 ({sk[14], i_5_, i_4_, i_1_, i_2_, i_0_, x5112x}, o_36_);
	defparam lut_67.LUT_SIZE = 7;
	defparam lut_67.mask = 128'h555f55ff5f5f5ffffbfbdbfbfbfbfbfb;

	lut_sub lut_75 ({sk[15], i_7_, i_6_, i_1_, i_2_, i_0_, n_n7}, o_27_);
	defparam lut_75.LUT_SIZE = 7;
	defparam lut_75.mask = 128'h555f55ff5f5f5fff0000000400000000;

	lut_sub lut_77 ({sk[16], i_1_, i_2_, i_0_, x102x}, o_14_);
	defparam lut_77.LUT_SIZE = 5;
	defparam lut_77.mask = 32'h57571000;

	lut_sub lut_79 ({sk[17], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, o_35_);
	defparam lut_79.LUT_SIZE = 7;
	defparam lut_79.mask = 128'h555f55ff5f5f5fffff7fffffff3fff9f;

	lut_sub lut_88 ({sk[18], i_1_, i_2_, i_0_, x124x}, o_28_);
	defparam lut_88.LUT_SIZE = 5;
	defparam lut_88.mask = 32'h57570100;

	lut_sub lut_90 ({sk[19], i_1_, i_2_, i_0_, x102x}, o_13_);
	defparam lut_90.LUT_SIZE = 5;
	defparam lut_90.mask = 32'h57570040;

	lut_sub lut_92 ({sk[20], i_7_, i_6_, x5107x, x5108x, x5109x}, o_34_);
	defparam lut_92.LUT_SIZE = 6;
	defparam lut_92.mask = 64'h000fffffafcfefe0;

	lut_sub lut_100 ({sk[21], i_7_, i_6_, x3194x}, o_21_);
	defparam lut_100.LUT_SIZE = 4;
	defparam lut_100.mask = 16'h3f44;

	lut_sub lut_103 ({sk[22], i_1_, i_2_, i_0_, x102x}, o_16_);
	defparam lut_103.LUT_SIZE = 5;
	defparam lut_103.mask = 32'h33ff0010;

	lut_sub lut_105 ({sk[23], i_7_, i_6_, x5104x, x5105x, x5106x}, o_40_);
	defparam lut_105.LUT_SIZE = 6;
	defparam lut_105.mask = 64'h00ffffffcfd0cf9f;

	lut_sub lut_112 ({sk[24], i_2_, i_0_, x5103x}, o_33_);
	defparam lut_112.LUT_SIZE = 4;
	defparam lut_112.mask = 16'h3ffe;

	lut_sub lut_116 ({sk[25], i_1_, i_2_, i_0_, x124x, x121x}, o_22_);
	defparam lut_116.LUT_SIZE = 6;
	defparam lut_116.mask = 64'h00ffffff07000000;

	lut_sub lut_119 ({sk[26], i_1_, i_2_, i_0_, x102x}, o_15_);
	defparam lut_119.LUT_SIZE = 5;
	defparam lut_119.mask = 32'h33ff0004;

	lut_sub lut_121 ({sk[27], i_3_, i_4_, x5100x, x5101x, x5102x}, o_32_);
	defparam lut_121.LUT_SIZE = 6;
	defparam lut_121.mask = 64'h00fffffff0dfef9f;

	lut_sub lut_130 ({sk[28], i_7_, i_5_, i_6_, i_3_, i_4_, n_n0}, o_23_);
	defparam lut_130.LUT_SIZE = 7;
	defparam lut_130.mask = 128'h5f5f5f5f7f7f7f7f0000050500000505;

	lut_sub lut_136 ({sk[29], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, o_18_);
	defparam lut_136.LUT_SIZE = 7;
	defparam lut_136.mask = 128'h5f5f5f5f7f7f7f7f0000002000000000;

	lut_sub lut_138 ({sk[30], i_6_, x5098x, x5099x}, o_31_);
	defparam lut_138.LUT_SIZE = 4;
	defparam lut_138.mask = 16'h558b;

	lut_sub lut_141 ({sk[31], i_7_, i_6_, i_1_, i_2_, i_0_, n_n7}, o_24_);
	defparam lut_141.LUT_SIZE = 7;
	defparam lut_141.mask = 128'h7fff7fff7fff7fff0000400000000000;

	lut_sub lut_143 ({sk[32], i_7_, i_5_, i_6_, i_3_, i_4_, x5127x}, o_17_);
	defparam lut_143.LUT_SIZE = 7;
	defparam lut_143.mask = 128'h7fff7fff7fff7fffbabaaaaababaaaaa;

	lut_sub lut_152 ({sk[33], i_7_, i_6_, x5096x, x5097x}, o_56_);
	defparam lut_152.LUT_SIZE = 5;
	defparam lut_152.mask = 32'h5f5faba8;

	lut_sub lut_157 ({sk[34], i_7_, i_6_, x5093x, x5094x, x5095x}, o_43_);
	defparam lut_157.LUT_SIZE = 6;
	defparam lut_157.mask = 64'h33ffffff95bab5a5;

	lut_sub lut_166 ({sk[35], i_1_, i_2_, i_0_, x121x}, o_30_);
	defparam lut_166.LUT_SIZE = 5;
	defparam lut_166.mask = 32'h5f5f0001;

	lut_sub lut_168 ({sk[36], i_2_, i_0_, x5091x, x5092x}, o_55_);
	defparam lut_168.LUT_SIZE = 5;
	defparam lut_168.mask = 32'h5f5f676d;

	lut_sub lut_174 ({sk[37], i_3_, i_4_, i_1_, i_2_, i_0_, x5089x}, o_44_);
	defparam lut_174.LUT_SIZE = 7;
	defparam lut_174.mask = 128'h7fff7fff7fff7fffefef6fefefefefef;

	lut_sub lut_182 ({sk[38], i_3_, i_4_, i_1_, i_2_, i_0_, x5088x}, o_58_);
	defparam lut_182.LUT_SIZE = 7;
	defparam lut_182.mask = 128'h7fff7fff7fff7fffffffffff5559fff3;

	lut_sub lut_195 ({sk[39], i_5_, i_3_, i_1_, i_2_, i_0_}, o_41_);
	defparam lut_195.LUT_SIZE = 6;
	defparam lut_195.mask = 64'h33fffffffbfffbbf;

	lut_sub lut_206 ({sk[40], i_2_, i_0_, x5084x, x5085x}, o_57_);
	defparam lut_206.LUT_SIZE = 5;
	defparam lut_206.mask = 32'h5f5fe7df;

	lut_sub lut_214 ({sk[41], i_7_, i_5_, i_6_, i_4_, x5082x}, o_42_);
	defparam lut_214.LUT_SIZE = 6;
	defparam lut_214.mask = 64'h33ffffffff7ffafa;

	lut_sub lut_221 ({sk[42], i_7_, i_6_, i_1_, i_2_, i_0_, n_n7}, o_20_);
	defparam lut_221.LUT_SIZE = 7;
	defparam lut_221.mask = 128'h7fff7fff7fff7fff1000000010000000;

	lut_sub lut_224 ({sk[43], i_3_, i_4_, x5079x, x5080x, x5081x}, o_52_);
	defparam lut_224.LUT_SIZE = 6;
	defparam lut_224.mask = 64'h33ffffffaf2feaf0;

	lut_sub lut_233 ({sk[44], i_2_, i_0_, x5077x, x5078x}, o_47_);
	defparam lut_233.LUT_SIZE = 5;
	defparam lut_233.mask = 32'h5f5fef7d;

	lut_sub lut_241 ({sk[45], i_7_, i_6_, x5075x, x5076x}, o_51_);
	defparam lut_241.LUT_SIZE = 5;
	defparam lut_241.mask = 32'h5f5f5756;

	lut_sub lut_246 ({sk[46], i_2_, i_0_, x5074x}, o_48_);
	defparam lut_246.LUT_SIZE = 4;
	defparam lut_246.mask = 16'h55bf;

	lut_sub lut_250 ({sk[47], i_7_, i_6_, x5072x, x5073x}, o_54_);
	defparam lut_250.LUT_SIZE = 5;
	defparam lut_250.mask = 32'h5f5fcdc9;

	lut_sub lut_255 ({sk[48], i_2_, i_0_, x5070x, x5071x}, o_45_);
	defparam lut_255.LUT_SIZE = 5;
	defparam lut_255.mask = 32'h5f5fcf7f;

	lut_sub lut_261 ({sk[49], i_1_, i_2_, i_0_, x82x, x102x}, o_10_);
	defparam lut_261.LUT_SIZE = 6;
	defparam lut_261.mask = 64'h33ffffff00000070;

	lut_sub lut_264 ({sk[50], i_2_, i_0_, x5067x, x5068x, x5069x}, o_53_);
	defparam lut_264.LUT_SIZE = 6;
	defparam lut_264.mask = 64'h33ffffff707aef5f;

	lut_sub lut_274 ({sk[51], i_2_, i_0_, x5066x}, o_46_);
	defparam lut_274.LUT_SIZE = 4;
	defparam lut_274.mask = 16'h55bf;

	lut_sub lut_278 ({sk[52], i_2_, i_0_, x5065x}, o_61_);
	defparam lut_278.LUT_SIZE = 4;
	defparam lut_278.mask = 16'h55fe;

	lut_sub lut_282 ({sk[53], i_1_, i_2_, i_0_, x121x}, o_9_);
	defparam lut_282.LUT_SIZE = 5;
	defparam lut_282.mask = 32'h5f5f0400;

	lut_sub lut_284 ({sk[54], i_5_, i_6_, i_3_, i_4_, i_1_, i_0_}, o_62_);
	defparam lut_284.LUT_SIZE = 7;
	defparam lut_284.mask = 128'h7fff7fff7fff7fffeefffefffefffeff;

	lut_sub lut_292 ({sk[55], i_2_, i_0_, x5063x}, o_49_);
	defparam lut_292.LUT_SIZE = 4;
	defparam lut_292.mask = 16'h55fb;

	lut_sub lut_296 ({sk[56], i_1_, i_2_, i_0_, x82x}, o_7_);
	defparam lut_296.LUT_SIZE = 5;
	defparam lut_296.mask = 32'h5f5f0040;

	lut_sub lut_298 ({sk[57], i_1_, i_2_, i_0_, x82x}, o_8_);
	defparam lut_298.LUT_SIZE = 5;
	defparam lut_298.mask = 32'h5f5f0001;

	lut_sub lut_300 ({sk[58], i_1_, i_2_, i_0_, n_n8, n_n12, n_n16}, o_5_);
	defparam lut_300.LUT_SIZE = 7;
	defparam lut_300.mask = 128'h7fff7fff7fff7fff1515151515151515;

	lut_sub lut_317 ({sk[59], i_7_, i_6_, x5061x, x5062x}, o_59_);
	defparam lut_317.LUT_SIZE = 5;
	defparam lut_317.mask = 32'h5f5faba9;

	lut_sub lut_322 ({sk[60], i_7_, i_5_, i_6_, i_3_, i_4_, n_n1}, o_6_);
	defparam lut_322.LUT_SIZE = 7;
	defparam lut_322.mask = 128'h7fff7fff7fff7fff0400000004000000;

	lut_sub lut_325 ({sk[61], i_7_, i_5_, i_6_, i_3_, i_4_}, o_3_);
	defparam lut_325.LUT_SIZE = 6;
	defparam lut_325.mask = 64'h33ffffff00200000;

	lut_sub lut_327 ({sk[62], i_7_, i_6_, i_1_, i_2_, i_0_, n_n11}, o_4_);
	defparam lut_327.LUT_SIZE = 7;
	defparam lut_327.mask = 128'h7fff7fff7fff7fff0000555500000000;

	lut_sub lut_336 ({sk[63], i_1_, i_2_, i_0_}, n_n0);
	defparam lut_336.LUT_SIZE = 4;
	defparam lut_336.mask = 16'h5580;

	lut_sub lut_338 ({sk[64], i_5_, i_3_, i_4_}, n_n8);
	defparam lut_338.LUT_SIZE = 4;
	defparam lut_338.mask = 16'h5508;

	lut_sub lut_340 ({sk[65], i_7_, i_5_, i_6_, i_1_, i_0_}, x5121x);
	defparam lut_340.LUT_SIZE = 6;
	defparam lut_340.mask = 64'h33ffffff00000008;

	lut_sub lut_342 ({sk[66], i_7_, i_5_, i_6_, i_1_, i_2_, i_0_}, x5122x);
	defparam lut_342.LUT_SIZE = 7;
	defparam lut_342.mask = 128'h7fff7fff7fff7ffffafafafafafafada;

	lut_sub lut_349 ({sk[67], i_7_, i_5_, i_6_, i_1_, i_2_, i_0_}, x5119x);
	defparam lut_349.LUT_SIZE = 7;
	defparam lut_349.mask = 128'h7fff7fff7fff7fff0000000000400000;

	lut_sub lut_351 ({sk[68], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5117x);
	defparam lut_351.LUT_SIZE = 7;
	defparam lut_351.mask = 128'h7fff7fff7fff7fff8000400000000000;

	lut_sub lut_354 ({sk[69], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5118x);
	defparam lut_354.LUT_SIZE = 7;
	defparam lut_354.mask = 128'h7fff7fff7fff7fff8040006000400060;

	lut_sub lut_358 ({sk[70], i_5_, i_3_, i_4_}, n_n7);
	defparam lut_358.LUT_SIZE = 4;
	defparam lut_358.mask = 16'h5580;

	lut_sub lut_360 ({sk[71], i_7_, i_5_, i_6_, i_3_, i_4_}, x82x);
	defparam lut_360.LUT_SIZE = 6;
	defparam lut_360.mask = 64'h33ffffff00000008;

	lut_sub lut_362 ({sk[72], i_5_, i_3_, i_1_, i_2_, i_0_}, x5115x);
	defparam lut_362.LUT_SIZE = 6;
	defparam lut_362.mask = 64'h33ffffff04000440;

	lut_sub lut_365 ({sk[73], i_7_, i_5_, i_6_, i_3_, i_4_}, x121x);
	defparam lut_365.LUT_SIZE = 6;
	defparam lut_365.mask = 64'h33ffffff00000800;

	lut_sub lut_367 ({sk[74], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5114x);
	defparam lut_367.LUT_SIZE = 7;
	defparam lut_367.mask = 128'h7fff7fff7fff7fff88008c0000000000;

	lut_sub lut_371 ({sk[75], i_7_, i_5_, i_6_, i_3_, i_4_, i_1_}, x5112x);
	defparam lut_371.LUT_SIZE = 7;
	defparam lut_371.mask = 128'h7fff7fff7fff7fff0080000000000000;

	lut_sub lut_373 ({sk[76], i_7_, i_5_, i_6_, i_3_, i_4_}, x102x);
	defparam lut_373.LUT_SIZE = 6;
	defparam lut_373.mask = 64'h33ffffff00000002;

	lut_sub lut_375 ({sk[77], i_7_, i_5_, i_6_, i_3_, i_4_}, x124x);
	defparam lut_375.LUT_SIZE = 6;
	defparam lut_375.mask = 64'h33ffffff00000200;

	lut_sub lut_377 ({sk[78], i_5_, i_4_, i_1_, i_2_, i_0_}, x5107x);
	defparam lut_377.LUT_SIZE = 6;
	defparam lut_377.mask = 64'h33ffffff40000000;

	lut_sub lut_379 ({sk[79], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5108x);
	defparam lut_379.LUT_SIZE = 7;
	defparam lut_379.mask = 128'h7fff7fff7fff7fff2040004000000000;

	lut_sub lut_382 ({sk[80], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5109x);
	defparam lut_382.LUT_SIZE = 7;
	defparam lut_382.mask = 128'h7fff7fff7fff7fff004000400000ff00;

	lut_sub lut_388 ({sk[81], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x3194x);
	defparam lut_388.LUT_SIZE = 7;
	defparam lut_388.mask = 128'h7fff7fff7fff7fff0000400000000000;

	lut_sub lut_390 ({sk[82], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5104x);
	defparam lut_390.LUT_SIZE = 7;
	defparam lut_390.mask = 128'h7fff7fff7fff7fff8000000000000000;

	lut_sub lut_392 ({sk[83], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5105x);
	defparam lut_392.LUT_SIZE = 7;
	defparam lut_392.mask = 128'h7fff7fff7fff7fff4080402000c00060;

	lut_sub lut_397 ({sk[84], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5106x);
	defparam lut_397.LUT_SIZE = 7;
	defparam lut_397.mask = 128'h7fff7fff7fff7fff5100400000000000;

	lut_sub lut_401 ({sk[85], i_7_, i_5_, i_6_, i_3_, i_4_, i_1_}, x5103x);
	defparam lut_401.LUT_SIZE = 7;
	defparam lut_401.mask = 128'h7fff7fff7fff7fff0000000000c80044;

	lut_sub lut_405 ({sk[86], i_7_, i_5_, i_6_, i_1_, i_2_, i_0_}, x5100x);
	defparam lut_405.LUT_SIZE = 7;
	defparam lut_405.mask = 128'h7fff7fff7fff7fff0080000000000000;

	lut_sub lut_407 ({sk[87], i_5_, i_6_, i_1_, i_2_, i_0_}, x5101x);
	defparam lut_407.LUT_SIZE = 6;
	defparam lut_407.mask = 64'h33ffffff40004040;

	lut_sub lut_410 ({sk[88], i_5_, i_6_, i_1_, i_2_, i_0_}, x5102x);
	defparam lut_410.LUT_SIZE = 6;
	defparam lut_410.mask = 64'h33ffffff60202020;

	lut_sub lut_413 ({sk[89], i_5_, i_4_, i_1_, i_2_, i_0_}, x5098x);
	defparam lut_413.LUT_SIZE = 6;
	defparam lut_413.mask = 64'h33ffffff40000000;

	lut_sub lut_415 ({sk[90], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5099x);
	defparam lut_415.LUT_SIZE = 7;
	defparam lut_415.mask = 128'h7fff7fff7fff7fff0000000000c00060;

	lut_sub lut_419 ({sk[91], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5127x);
	defparam lut_419.LUT_SIZE = 7;
	defparam lut_419.mask = 128'h7fff7fff7fff7fffffffffbfffffffff;

	lut_sub lut_435 ({sk[92], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5096x);
	defparam lut_435.LUT_SIZE = 7;
	defparam lut_435.mask = 128'h7fff7fff7fff7fff0000080022000200;

	lut_sub lut_439 ({sk[93], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5097x);
	defparam lut_439.LUT_SIZE = 7;
	defparam lut_439.mask = 128'h7fff7fff7fff7fff0000080800000008;

	lut_sub lut_442 ({sk[94], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5093x);
	defparam lut_442.LUT_SIZE = 7;
	defparam lut_442.mask = 128'h7fff7fff7fff7fffc000400000000000;

	lut_sub lut_445 ({sk[95], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5094x);
	defparam lut_445.LUT_SIZE = 7;
	defparam lut_445.mask = 128'h7fff7fff7fff7fff11001000ff00ff00;

	lut_sub lut_449 ({sk[96], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5095x);
	defparam lut_449.LUT_SIZE = 7;
	defparam lut_449.mask = 128'h7fff7fff7fff7fff91c0106000c00060;

	lut_sub lut_460 ({sk[97], i_7_, i_5_, i_6_, i_3_, i_4_, i_1_}, x5091x);
	defparam lut_460.LUT_SIZE = 7;
	defparam lut_460.mask = 128'h7fff7fff7fff7fff5010101050101054;

	lut_sub lut_466 ({sk[98], i_7_, i_5_, i_6_, i_3_, i_4_, i_1_}, x5092x);
	defparam lut_466.LUT_SIZE = 7;
	defparam lut_466.mask = 128'h7fff7fff7fff7ffffafefefefafefeba;

	lut_sub lut_479 ({sk[99], i_5_, i_6_, i_3_, i_4_, i_1_}, x5089x);
	defparam lut_479.LUT_SIZE = 6;
	defparam lut_479.mask = 64'h33ffffff80000000;

	lut_sub lut_481 ({sk[100], i_7_, i_5_, i_6_, i_1_, i_2_, i_0_}, x5088x);
	defparam lut_481.LUT_SIZE = 7;
	defparam lut_481.mask = 128'h7fff7fff7fff7ffffffdfdfdff7dfdfc;

	lut_sub lut_492 ({sk[101], i_7_, i_5_, i_6_, i_3_, i_4_, i_1_}, x5084x);
	defparam lut_492.LUT_SIZE = 7;
	defparam lut_492.mask = 128'h7fff7fff7fff7fff501010105050105c;

	lut_sub lut_499 ({sk[102], i_7_, i_5_, i_6_, i_3_, i_4_, i_1_}, x5085x);
	defparam lut_499.LUT_SIZE = 7;
	defparam lut_499.mask = 128'h7fff7fff7fff7ffffafefefefafafeb2;

	lut_sub lut_512 ({sk[103], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5082x);
	defparam lut_512.LUT_SIZE = 7;
	defparam lut_512.mask = 128'h7fff7fff7fff7fff4000500000000000;

	lut_sub lut_515 ({sk[104], i_1_, i_2_, i_0_}, x5079x);
	defparam lut_515.LUT_SIZE = 4;
	defparam lut_515.mask = 16'h5580;

	lut_sub lut_517 ({sk[105], i_5_, i_6_, i_1_, i_2_, i_0_}, x5080x);
	defparam lut_517.LUT_SIZE = 6;
	defparam lut_517.mask = 64'h33ffffff6a4a4a4a;

	lut_sub lut_521 ({sk[106], i_5_, i_6_, i_1_, i_2_, i_0_}, x5081x);
	defparam lut_521.LUT_SIZE = 6;
	defparam lut_521.mask = 64'h33ffffffb5000000;

	lut_sub lut_525 ({sk[107], i_7_, i_5_, i_6_, i_3_, i_4_, i_1_}, x5077x);
	defparam lut_525.LUT_SIZE = 7;
	defparam lut_525.mask = 128'h7fff7fff7fff7fff0000000000880004;

	lut_sub lut_528 ({sk[108], i_7_, i_5_, i_6_, i_3_, i_4_, i_1_}, x5078x);
	defparam lut_528.LUT_SIZE = 7;
	defparam lut_528.mask = 128'h7fff7fff7fff7fffaaeeeeeeaaeeeeea;

	lut_sub lut_542 ({sk[109], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5075x);
	defparam lut_542.LUT_SIZE = 7;
	defparam lut_542.mask = 128'h7fff7fff7fff7fff0500a10004000000;

	lut_sub lut_546 ({sk[110], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5076x);
	defparam lut_546.LUT_SIZE = 7;
	defparam lut_546.mask = 128'h7fff7fff7fff7ffffafa5e7efffaff7e;

	lut_sub lut_561 ({sk[111], i_7_, i_5_, i_6_, i_3_, i_4_, i_1_}, x5074x);
	defparam lut_561.LUT_SIZE = 7;
	defparam lut_561.mask = 128'h7fff7fff7fff7fff0a0202020a02020a;

	lut_sub lut_569 ({sk[112], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5072x);
	defparam lut_569.LUT_SIZE = 7;
	defparam lut_569.mask = 128'h7fff7fff7fff7fff0808020200080002;

	lut_sub lut_574 ({sk[113], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5073x);
	defparam lut_574.LUT_SIZE = 7;
	defparam lut_574.mask = 128'h7fff7fff7fff7fff0800020027008a00;

	lut_sub lut_583 ({sk[114], i_7_, i_5_, i_6_, i_4_, i_1_}, x5070x);
	defparam lut_583.LUT_SIZE = 6;
	defparam lut_583.mask = 64'h33ffffff00000800;

	lut_sub lut_585 ({sk[115], i_7_, i_5_, i_6_, i_4_, i_1_}, x5071x);
	defparam lut_585.LUT_SIZE = 6;
	defparam lut_585.mask = 64'h33ffffffaeeea6ee;

	lut_sub lut_598 ({sk[116], i_7_, i_5_, i_6_, i_3_, i_4_}, x5067x);
	defparam lut_598.LUT_SIZE = 6;
	defparam lut_598.mask = 64'h33ffffff00000008;

	lut_sub lut_600 ({sk[117], i_7_, i_5_, i_6_, i_3_, i_4_, i_1_}, x5068x);
	defparam lut_600.LUT_SIZE = 7;
	defparam lut_600.mask = 128'h7fff7fff7fff7fff501010105010101c;

	lut_sub lut_605 ({sk[118], i_7_, i_5_, i_6_, i_3_, i_4_, i_1_}, x5069x);
	defparam lut_605.LUT_SIZE = 7;
	defparam lut_605.mask = 128'h7fff7fff7fff7ffffafefefefafefeba;

	lut_sub lut_618 ({sk[119], i_7_, i_5_, i_6_, i_3_, i_4_, i_1_}, x5066x);
	defparam lut_618.LUT_SIZE = 7;
	defparam lut_618.mask = 128'h7fff7fff7fff7fff5010101050501010;

	lut_sub lut_624 ({sk[120], i_5_, i_6_, i_3_, i_4_, i_1_}, x5065x);
	defparam lut_624.LUT_SIZE = 6;
	defparam lut_624.mask = 64'h33ffffff0a020202;

	lut_sub lut_628 ({sk[121], i_5_, i_6_, i_3_, i_4_, i_1_}, x5063x);
	defparam lut_628.LUT_SIZE = 6;
	defparam lut_628.mask = 64'h33ffffffa8202020;

	lut_sub lut_633 ({sk[122], i_5_, i_3_, i_4_}, n_n12);
	defparam lut_633.LUT_SIZE = 4;
	defparam lut_633.mask = 16'h5502;

	lut_sub lut_635 ({sk[123], i_7_, i_6_}, n_n16);
	defparam lut_635.LUT_SIZE = 3;
	defparam lut_635.mask = 8'h54;

	lut_sub lut_637 ({sk[124], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5061x);
	defparam lut_637.LUT_SIZE = 7;
	defparam lut_637.mask = 128'h7fff7fff7fff7fffa9009c0000000000;

	lut_sub lut_644 ({sk[125], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x5062x);
	defparam lut_644.LUT_SIZE = 7;
	defparam lut_644.mask = 128'h7fff7fff7fff7fff0101101000010010;

	lut_sub lut_649 ({sk[126], i_1_, i_2_, i_0_}, n_n1);
	defparam lut_649.LUT_SIZE = 4;
	defparam lut_649.mask = 16'h5520;

	lut_sub lut_651 ({sk[127], i_5_, i_3_, i_4_}, n_n11);
	defparam lut_651.LUT_SIZE = 4;
	defparam lut_651.mask = 16'h5520;


endmodule