module ex1010 (
	i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, 
	i_8_, i_9_, o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, 
	o_8_, o_9_);

input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_;

output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_;

wire n1, n2, n6, n4, n5, n3, n10, n8, n9, n7, n12, n13, n14, n15, n11, n17, n18, n19, n20, n21, n16, n25, n26, n23, n24, n22, n28, n29, n30, n31, n32, n33, n34, n35, n27, n37, n38, n39, n40, n41, n42, n36, n44, n45, n46, n47, n48, n43, n50, n51, n52, n53, n54, n49, n58, n59, n56, n57, n55, n63, n64, n61, n62, n60, n67, n68, n66, n65, n72, n70, n71, n69, n75, n74, n73, n77, n78, n79, n80, n76, n82, n83, n84, n85, n86, n87, n81, n89, n90, n91, n92, n93, n94, n88, n96, n97, n98, n99, n100, n101, n102, n103, n95, n105, n106, n107, n108, n109, n110, n104, n113, n114, n112, n111, n116, n117, n118, n115, n121, n122, n120, n119, n125, n126, n124, n123, n129, n128, n127, n132, n131, n130, n134, n135, n136, n137, n138, n139, n140, n141, n133, n143, n144, n145, n146, n142, n148, n149, n150, n151, n152, n153, n147, n155, n156, n157, n158, n159, n160, n154, n162, n163, n164, n165, n166, n167, n161, n170, n171, n169, n168, n174, n175, n173, n172, n177, n178, n176, n180, n181, n182, n183, n184, n185, n186, n187, n179, n190, n191, n189, n188, n195, n193, n194, n192, n197, n198, n199, n200, n201, n202, n203, n196, n205, n206, n207, n208, n209, n210, n211, n212, n204, n214, n215, n216, n217, n218, n219, n213, n222, n223, n221, n220, n226, n227, n225, n224, n231, n229, n230, n228, n234, n233, n232, n236, n237, n238, n239, n240, n241, n235, n244, n243, n242, n246, n247, n248, n249, n250, n251, n252, n253, n245, n255, n256, n257, n258, n254, n261, n262, n260, n259, n265, n266, n264, n263, n268, n269, n270, n271, n267, n272, n273, n274, n275, n276, n277, n281, n282, n279, n280, n278, n284, n285, n286, n287, n288, n289, n283, n291, n292, n293, n294, n295, n296, n297, n298, n290, n300, n301, n302, n303, n304, n305, n306, n307, n299, n310, n311, n309, n308, n313, n314, n315, n316, n317, n318, n319, n320, n312, n322, n323, n324, n325, n326, n327, n328, n321, n330, n331, n332, n333, n334, n335, n329, n337, n338, n339, n340, n341, n342, n336, n344, n345, n346, n347, n348, n349, n343, n351, n352, n353, n354, n355, n356, n350, n358, n359, n360, n361, n362, n363, n364, n365, n357, n367, n368, n369, n370, n371, n372, n373, n374, n366, n375, n376, n377, n378, n379, n380, n382, n383, n384, n385, n386, n387, n388, n389, n381, n391, n396, n398, n400, n402, n403, n404, n406, n407, n408, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n540, n541, n539, n542, n543, n544, n545, n546, n547, n548, n549, n551, n550, n552, n553, n555, n556, n554, n558, n557, n559, n560, n561, n563, n564, n562, n565, n566, n567, n569, n568, n570, n572, n573, n571, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n589, n588, n590, n591, n592, n594, n593, n596, n597, n595, n599, n598, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n614, n613, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n634, n633, n636, n635, n637, n638, n640, n639, n642, n641, n643, n644, n645, n647, n646, n648, n649, n651, n650, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n669, n668, n671, n670, n673, n672, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n696, n695, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n716, n715, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n742, n741, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n758, n757, n759, n760, n761, n763, n762, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n805, n804, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850;

assign o_0_ = ( (~ n381) ) ;
 assign o_1_ = ( (~ n2) ) ;
 assign o_2_ = ( (~ n366) ) ;
 assign o_3_ = ( (~ n343) ) ;
 assign o_4_ = ( (~ n312) ) ;
 assign o_5_ = ( (~ n1) ) ;
 assign o_6_ = ( (~ n235) ) ;
 assign o_7_ = ( (~ n179) ) ;
 assign o_8_ = ( (~ n133) ) ;
 assign o_9_ = ( (~ n76) ) ;
 assign n1 = ( n123  &  n16  &  n272  &  n273  &  n274  &  n275  &  n276  &  n277 ) ;
 assign n2 = ( n65  &  n375  &  n119  &  n376  &  n377  &  n378  &  n379  &  n380 ) ;
 assign n6 = ( n189  &  n417 ) | ( n460  &  n417 ) | ( n189  &  n439 ) | ( n460  &  n439 ) ;
 assign n4 = ( (~ i_9_) ) | ( n410 ) ;
 assign n5 = ( n402 ) | ( n427 ) ;
 assign n3 = ( n6  &  n4 ) | ( n6  &  n5 ) ;
 assign n10 = ( n15  &  n193 ) | ( n461  &  n193 ) | ( n15  &  n462 ) | ( n461  &  n462 ) ;
 assign n8 = ( (~ i_9_) ) | ( n391 ) ;
 assign n9 = ( n402 ) | ( n438 ) ;
 assign n7 = ( n10  &  n8 ) | ( n10  &  n9 ) ;
 assign n12 = ( i_9_ ) | ( n421 ) ;
 assign n13 = ( n396 ) | ( n422 ) ;
 assign n14 = ( n391 ) | ( n431 ) ;
 assign n15 = ( i_9_ ) | ( n398 ) ;
 assign n11 = ( n12  &  n14 ) | ( n13  &  n14 ) | ( n12  &  n15 ) | ( n13  &  n15 ) ;
 assign n17 = ( n189 ) | ( n74 ) ;
 assign n18 = ( n420 ) | ( n260 ) ;
 assign n19 = ( n546  &  n292  &  n547 ) ;
 assign n20 = ( n544  &  n545  &  n243 ) | ( n544  &  n545  &  n457 ) ;
 assign n21 = ( n542  &  n543  &  n97  &  n537  &  n539  &  n538 ) ;
 assign n16 = ( n17  &  n18  &  n11  &  n3  &  n7  &  n19  &  n20  &  n21 ) ;
 assign n25 = ( n12 ) | ( n437 ) ;
 assign n26 = ( n417 ) | ( n173 ) ;
 assign n23 = ( (~ i_9_) ) | ( n407 ) ;
 assign n24 = ( n406 ) | ( n427 ) ;
 assign n22 = ( n25  &  n26  &  n23 ) | ( n25  &  n26  &  n24 ) ;
 assign n28 = ( n8 ) | ( n233 ) ;
 assign n29 = ( n243 ) | ( n468 ) ;
 assign n30 = ( n291  &  n189 ) | ( n291  &  n469 ) ;
 assign n31 = ( n536  &  n22  &  n61 ) | ( n536  &  n22  &  n470 ) ;
 assign n32 = ( n23 ) | ( n62 ) ;
 assign n33 = ( n189 ) | ( n466 ) ;
 assign n34 = ( n4 ) | ( n467 ) ;
 assign n35 = ( n360  &  n535  &  n23 ) | ( n360  &  n535  &  n464 ) ;
 assign n27 = ( n28  &  n29  &  n30  &  n31  &  n32  &  n33  &  n34  &  n35 ) ;
 assign n37 = ( n533  &  n8 ) | ( n533  &  n471 ) ;
 assign n38 = ( n417 ) | ( n472 ) ;
 assign n39 = ( n66  &  n4 ) | ( n15  &  n4 ) | ( n66  &  n450 ) | ( n15  &  n450 ) ;
 assign n40 = ( n189 ) | ( n309 ) ;
 assign n41 = ( n420  &  n8 ) | ( n475  &  n8 ) | ( n420  &  n459 ) | ( n475  &  n459 ) ;
 assign n42 = ( n534  &  n300  &  n279 ) | ( n534  &  n300  &  n462 ) ;
 assign n36 = ( n37  &  n38  &  n39  &  n40  &  n41  &  n42 ) ;
 assign n44 = ( n61 ) | ( n477 ) ;
 assign n45 = ( n71 ) | ( n13 ) ;
 assign n46 = ( n193  &  n279 ) | ( n476  &  n279 ) | ( n193  &  n444 ) | ( n476  &  n444 ) ;
 assign n47 = ( n15  &  n193 ) | ( n225  &  n193 ) | ( n15  &  n444 ) | ( n225  &  n444 ) ;
 assign n48 = ( n15  &  n400 ) | ( n194  &  n400 ) | ( n15  &  n443 ) | ( n194  &  n443 ) ;
 assign n43 = ( n44  &  n45  &  n46  &  n47  &  n48 ) ;
 assign n50 = ( n189 ) | ( n479 ) ;
 assign n51 = ( n417 ) | ( n461 ) ;
 assign n52 = ( n193  &  n417 ) | ( n478  &  n417 ) | ( n193  &  n428 ) | ( n478  &  n428 ) ;
 assign n53 = ( n229  &  n56 ) | ( n480  &  n56 ) | ( n229  &  n456 ) | ( n480  &  n456 ) ;
 assign n54 = ( n12  &  n279 ) | ( n474  &  n279 ) | ( n12  &  n461 ) | ( n474  &  n461 ) ;
 assign n49 = ( n50  &  n51  &  n52  &  n53  &  n54 ) ;
 assign n58 = ( n443  &  n424 ) | ( n483  &  n424 ) | ( n443  &  n56 ) | ( n483  &  n56 ) ;
 assign n59 = ( n197  &  n532  &  n229 ) | ( n197  &  n532  &  n481 ) ;
 assign n56 = ( i_9_ ) | ( n441 ) ;
 assign n57 = ( n414 ) | ( n447 ) ;
 assign n55 = ( n58  &  n59  &  n56 ) | ( n58  &  n59  &  n57 ) ;
 assign n63 = ( n4  &  n193 ) | ( n120  &  n193 ) | ( n4  &  n173 ) | ( n120  &  n173 ) ;
 assign n64 = ( n530  &  n531  &  n189 ) | ( n530  &  n531  &  n169 ) ;
 assign n61 = ( (~ i_9_) ) | ( n447 ) ;
 assign n62 = ( n416 ) | ( n423 ) ;
 assign n60 = ( n63  &  n64  &  n61 ) | ( n63  &  n64  &  n62 ) ;
 assign n67 = ( n443 ) | ( n488 ) ;
 assign n68 = ( n529  &  n96  &  n71 ) | ( n529  &  n96  &  n487 ) ;
 assign n66 = ( n422 ) | ( n423 ) ;
 assign n65 = ( n67  &  n68  &  n66 ) | ( n67  &  n68  &  n56 ) ;
 assign n72 = ( n23  &  n189 ) | ( n450  &  n189 ) | ( n23  &  n62 ) | ( n450  &  n62 ) ;
 assign n70 = ( n412 ) | ( n413 ) ;
 assign n71 = ( i_9_ ) | ( n438 ) ;
 assign n69 = ( n72  &  n70 ) | ( n72  &  n71 ) ;
 assign n75 = ( n4  &  n71 ) | ( n470  &  n71 ) | ( n4  &  n489 ) | ( n470  &  n489 ) ;
 assign n74 = ( n402 ) | ( n441 ) ;
 assign n73 = ( n75  &  n8 ) | ( n75  &  n74 ) ;
 assign n77 = ( n445  &  n56 ) | ( n189  &  n56 ) | ( n445  &  n446 ) | ( n189  &  n446 ) ;
 assign n78 = ( n27  &  n36  &  n16  &  n49  &  n55  &  n43 ) ;
 assign n79 = ( n570  &  n574  &  n571  &  n567  &  n566  &  n568 ) ;
 assign n80 = ( n561  &  n565  &  n562  &  n560  &  n557  &  n554 ) ;
 assign n76 = ( n65  &  n69  &  n60  &  n77  &  n73  &  n78  &  n79  &  n80 ) ;
 assign n82 = ( n604  &  n71 ) | ( n604  &  n495 ) ;
 assign n83 = ( n8 ) | ( n488 ) ;
 assign n84 = ( n56 ) | ( n449  &  n473 ) ;
 assign n85 = ( n603  &  n443 ) | ( n603  &  n479 ) ;
 assign n86 = ( n601  &  n602  &  n15 ) | ( n601  &  n602  &  n280 ) ;
 assign n87 = ( n600  &  n257  &  n542  &  n181  &  n28  &  n598  &  n271  &  n595 ) ;
 assign n81 = ( n82  &  n83  &  n84  &  n85  &  n86  &  n87 ) ;
 assign n89 = ( n4  &  n8 ) | ( n501  &  n8 ) | ( n4  &  n452 ) | ( n501  &  n452 ) ;
 assign n90 = ( n23 ) | ( n5 ) ;
 assign n91 = ( n443  &  n61 ) | ( n469  &  n61 ) | ( n443  &  n504 ) | ( n469  &  n504 ) ;
 assign n92 = ( n590  &  n588  &  n71 ) | ( n590  &  n588  &  n456 ) ;
 assign n93 = ( n284  &  n593  &  n279 ) | ( n284  &  n593  &  n439 ) ;
 assign n94 = ( n592  &  n591  &  n428 ) | ( n592  &  n591  &  n15 ) ;
 assign n88 = ( n89  &  n90  &  n91  &  n92  &  n93  &  n94 ) ;
 assign n96 = ( n443 ) | ( n486 ) ;
 assign n97 = ( n15 ) | ( n449 ) ;
 assign n98 = ( n45  &  n193 ) | ( n45  &  n499 ) ;
 assign n99 = ( n243  &  n56 ) | ( n446  &  n56 ) | ( n243  &  n506 ) | ( n446  &  n506 ) ;
 assign n100 = ( n587  &  n279 ) | ( n587  &  n505 ) ;
 assign n101 = ( n584  &  n443 ) | ( n584  &  n507 ) ;
 assign n102 = ( n582  &  n583  &  n420 ) | ( n582  &  n583  &  n479 ) ;
 assign n103 = ( n586  &  n585  &  n8 ) | ( n586  &  n585  &  n442 ) ;
 assign n95 = ( n96  &  n97  &  n98  &  n99  &  n100  &  n101  &  n102  &  n103 ) ;
 assign n105 = ( n61  &  n243 ) | ( n74  &  n243 ) | ( n61  &  n476 ) | ( n74  &  n476 ) ;
 assign n106 = ( n435 ) | ( n71 ) ;
 assign n107 = ( n581  &  n279 ) | ( n581  &  n465 ) ;
 assign n108 = ( n443 ) | ( n458 ) ;
 assign n109 = ( n579  &  n580  &  n189 ) | ( n579  &  n580  &  n481 ) ;
 assign n110 = ( n577  &  n578  &  n193 ) | ( n577  &  n578  &  n14 ) ;
 assign n104 = ( n105  &  n106  &  n107  &  n108  &  n109  &  n110 ) ;
 assign n113 = ( n243  &  n61 ) | ( n509  &  n61 ) | ( n243  &  n492 ) | ( n509  &  n492 ) ;
 assign n114 = ( n575  &  n576  &  n61 ) | ( n575  &  n576  &  n5 ) ;
 assign n112 = ( n396 ) | ( n413 ) ;
 assign n111 = ( n113  &  n114  &  n56 ) | ( n113  &  n114  &  n112 ) ;
 assign n116 = ( n229  &  n243 ) | ( n484  &  n243 ) | ( n229  &  n510 ) | ( n484  &  n510 ) ;
 assign n117 = ( n56 ) | ( n511 ) ;
 assign n118 = ( n403  &  n23 ) | ( n443  &  n23 ) | ( n403  &  n74 ) | ( n443  &  n74 ) ;
 assign n115 = ( n116  &  n117  &  n118  &  n33 ) ;
 assign n121 = ( n417  &  n279 ) | ( n437  &  n279 ) | ( n417  &  n512 ) | ( n437  &  n512 ) ;
 assign n122 = ( n71  &  n56 ) | ( n453  &  n56 ) | ( n71  &  n513 ) | ( n453  &  n513 ) ;
 assign n120 = ( n398 ) | ( n423 ) ;
 assign n119 = ( n121  &  n122  &  n61 ) | ( n121  &  n122  &  n120 ) ;
 assign n125 = ( n514 ) | ( n12  &  n417 ) ;
 assign n126 = ( n352  &  n23 ) | ( n352  &  n477 ) ;
 assign n124 = ( n402 ) | ( n416 ) ;
 assign n123 = ( n125  &  n126  &  n61 ) | ( n125  &  n126  &  n124 ) ;
 assign n129 = ( n61  &  n71 ) | ( n515  &  n71 ) | ( n61  &  n512 ) | ( n515  &  n512 ) ;
 assign n128 = ( n406 ) | ( n447 ) ;
 assign n127 = ( n129  &  n56 ) | ( n129  &  n128 ) ;
 assign n132 = ( n61  &  n4 ) | ( n9  &  n4 ) | ( n61  &  n486 ) | ( n9  &  n486 ) ;
 assign n131 = ( n414 ) | ( n441 ) ;
 assign n130 = ( n132  &  n4 ) | ( n132  &  n131 ) ;
 assign n134 = ( n4  &  n417 ) | ( n62  &  n417 ) | ( n4  &  n494 ) | ( n62  &  n494 ) ;
 assign n135 = ( n193  &  n23 ) | ( n493  &  n23 ) | ( n193  &  n490 ) | ( n493  &  n490 ) ;
 assign n136 = ( n8  &  n193 ) | ( n448  &  n193 ) | ( n8  &  n494 ) | ( n448  &  n494 ) ;
 assign n137 = ( n15  &  n229 ) | ( n482  &  n229 ) | ( n15  &  n448 ) | ( n482  &  n448 ) ;
 assign n138 = ( n607  &  n606  &  n279 ) | ( n607  &  n606  &  n14 ) ;
 assign n139 = ( n613  &  n615  &  n612  &  n611  &  n610  &  n359  &  n609  &  n608 ) ;
 assign n140 = ( n104  &  n111  &  n115  &  n119  &  n88  &  n95  &  n81  &  n625 ) ;
 assign n141 = ( n621  &  n622  &  n620  &  n619  &  n618  &  n623  &  n617  &  n616 ) ;
 assign n133 = ( n134  &  n135  &  n136  &  n137  &  n138  &  n139  &  n140  &  n141 ) ;
 assign n143 = ( n15  &  n8 ) | ( n465  &  n8 ) | ( n15  &  n62 ) | ( n465  &  n62 ) ;
 assign n144 = ( n629  &  n630  &  n439 ) | ( n629  &  n630  &  n56 ) ;
 assign n145 = ( n628  &  n71 ) | ( n628  &  n264 ) ;
 assign n146 = ( n626  &  n627  &  n189 ) | ( n626  &  n627  &  n521 ) ;
 assign n142 = ( n143  &  n144  &  n145  &  n146 ) ;
 assign n148 = ( n4 ) | ( n458 ) ;
 assign n149 = ( n243 ) | ( n225 ) ;
 assign n150 = ( n433  &  n61 ) | ( n15  &  n61 ) | ( n433  &  n519 ) | ( n15  &  n519 ) ;
 assign n151 = ( n61 ) | ( n485 ) ;
 assign n152 = ( n229  &  n71 ) | ( n485  &  n71 ) | ( n229  &  n473 ) | ( n485  &  n473 ) ;
 assign n153 = ( n541  &  n23 ) | ( n541  &  n260 ) ;
 assign n147 = ( n148  &  n149  &  n150  &  n151  &  n152  &  n153 ) ;
 assign n155 = ( n408 ) | ( n71 ) ;
 assign n156 = ( n189 ) | ( n5 ) ;
 assign n157 = ( n15  &  n417 ) | ( n455  &  n417 ) | ( n15  &  n453 ) | ( n455  &  n453 ) ;
 assign n158 = ( n12 ) | ( n523 ) ;
 assign n159 = ( n426  &  n61 ) | ( n189  &  n61 ) | ( n426  &  n309 ) | ( n189  &  n309 ) ;
 assign n160 = ( n189  &  n12 ) | ( n486  &  n12 ) | ( n189  &  n506 ) | ( n486  &  n506 ) ;
 assign n154 = ( n155  &  n156  &  n157  &  n158  &  n159  &  n160 ) ;
 assign n162 = ( n417 ) | ( n506 ) ;
 assign n163 = ( n56 ) | ( n493 ) ;
 assign n164 = ( n417  &  n56 ) | ( n525  &  n56 ) | ( n417  &  n461 ) | ( n525  &  n461 ) ;
 assign n165 = ( n23 ) | ( n467 ) ;
 assign n166 = ( n279 ) | ( n524 ) ;
 assign n167 = ( n193  &  n229 ) | ( n264  &  n229 ) | ( n193  &  n221 ) | ( n264  &  n221 ) ;
 assign n161 = ( n162  &  n163  &  n164  &  n165  &  n166  &  n167 ) ;
 assign n170 = ( n243  &  n66 ) | ( n513  &  n66 ) | ( n243  &  n71 ) | ( n513  &  n71 ) ;
 assign n171 = ( n322  &  n323  &  n12 ) | ( n322  &  n323  &  n494 ) ;
 assign n169 = ( n431 ) | ( n438 ) ;
 assign n168 = ( n170  &  n171  &  n23 ) | ( n170  &  n171  &  n169 ) ;
 assign n174 = ( n8  &  n443 ) | ( n503  &  n443 ) | ( n8  &  n477 ) | ( n503  &  n477 ) ;
 assign n175 = ( n420  &  n279 ) | ( n520  &  n279 ) | ( n420  &  n498 ) | ( n520  &  n498 ) ;
 assign n173 = ( n402 ) | ( n413 ) ;
 assign n172 = ( n174  &  n175  &  n56 ) | ( n174  &  n175  &  n173 ) ;
 assign n177 = ( n243  &  n193 ) | ( n502  &  n193 ) | ( n243  &  n112 ) | ( n502  &  n112 ) ;
 assign n178 = ( n4  &  n420 ) | ( n451  &  n420 ) | ( n4  &  n477 ) | ( n451  &  n477 ) ;
 assign n176 = ( n177  &  n178 ) ;
 assign n180 = ( n71  &  n56 ) | ( n518  &  n56 ) | ( n71  &  n500 ) | ( n518  &  n500 ) ;
 assign n181 = ( n23 ) | ( n120 ) ;
 assign n182 = ( n655  &  n654  &  n243 ) | ( n655  &  n654  &  n495 ) ;
 assign n183 = ( n547  &  n544  &  n206  &  n586  &  n653  &  n652 ) ;
 assign n184 = ( n27  &  n104  &  n442 ) | ( n27  &  n104  &  n61 ) ;
 assign n185 = ( n657  &  n656  &  n23 ) | ( n657  &  n656  &  n520 ) ;
 assign n186 = ( n161  &  n168  &  n172  &  n176  &  n147  &  n154  &  n142 ) ;
 assign n187 = ( n650  &  n199  &  n649  &  n648  &  n644  &  n643  &  n646  &  n641 ) ;
 assign n179 = ( n180  &  n181  &  n182  &  n183  &  n184  &  n185  &  n186  &  n187 ) ;
 assign n190 = ( n229 ) | ( n62 ) ;
 assign n191 = ( n12  &  n279 ) | ( n499  &  n279 ) | ( n12  &  n523 ) | ( n499  &  n523 ) ;
 assign n189 = ( (~ i_9_) ) | ( n432 ) ;
 assign n188 = ( n190  &  n191  &  n189 ) | ( n190  &  n191  &  n9 ) ;
 assign n195 = ( n443  &  n56 ) | ( n526  &  n56 ) | ( n443  &  n494 ) | ( n526  &  n494 ) ;
 assign n193 = ( i_9_ ) | ( n404 ) ;
 assign n194 = ( n423 ) | ( n447 ) ;
 assign n192 = ( n195  &  n193 ) | ( n195  &  n194 ) ;
 assign n197 = ( n243 ) | ( n482 ) ;
 assign n198 = ( n419 ) | ( n420 ) ;
 assign n199 = ( n437 ) | ( n71 ) ;
 assign n200 = ( n17  &  n44  &  n15 ) | ( n17  &  n44  &  n506 ) ;
 assign n201 = ( n667  &  n666  &  n279 ) | ( n667  &  n666  &  n264 ) ;
 assign n202 = ( n248  &  n634  &  n665  &  n249 ) ;
 assign n203 = ( n192  &  n127  &  n188  &  n11  &  n375  &  n674  &  n672  &  n670 ) ;
 assign n196 = ( n197  &  n198  &  n199  &  n148  &  n200  &  n201  &  n202  &  n203 ) ;
 assign n205 = ( n415 ) | ( n4 ) ;
 assign n206 = ( n443 ) | ( n459 ) ;
 assign n207 = ( n655  &  n12 ) | ( n655  &  n517 ) ;
 assign n208 = ( n193  &  n229 ) | ( n491  &  n229 ) | ( n193  &  n508 ) | ( n491  &  n508 ) ;
 assign n209 = ( n4 ) | ( n504 ) ;
 assign n210 = ( n8  &  n12 ) | ( n230  &  n12 ) | ( n8  &  n500 ) | ( n230  &  n500 ) ;
 assign n211 = ( n420 ) | ( n309  &  n497 ) ;
 assign n212 = ( n663  &  n664  &  n71 ) | ( n663  &  n664  &  n522 ) ;
 assign n204 = ( n205  &  n206  &  n207  &  n208  &  n209  &  n210  &  n211  &  n212 ) ;
 assign n214 = ( n443  &  n23 ) | ( n24  &  n23 ) | ( n443  &  n515 ) | ( n24  &  n515 ) ;
 assign n215 = ( n66 ) | ( n243 ) ;
 assign n216 = ( n662  &  n56 ) | ( n662  &  n482 ) ;
 assign n217 = ( n15 ) | ( n472 ) ;
 assign n218 = ( n18  &  n597  &  n61 ) | ( n18  &  n597  &  n460 ) ;
 assign n219 = ( n660  &  n661  &  n417 ) | ( n660  &  n661  &  n489 ) ;
 assign n213 = ( n214  &  n215  &  n216  &  n217  &  n218  &  n219 ) ;
 assign n222 = ( n364  &  n12 ) | ( n364  &  n473 ) ;
 assign n223 = ( n659  &  n658  &  n4 ) | ( n659  &  n658  &  n527 ) ;
 assign n221 = ( n423 ) | ( n427 ) ;
 assign n220 = ( n222  &  n223  &  n23 ) | ( n222  &  n223  &  n221 ) ;
 assign n226 = ( n243 ) | ( n517 ) ;
 assign n227 = ( n56  &  n229 ) | ( n496  &  n229 ) | ( n56  &  n521 ) | ( n496  &  n521 ) ;
 assign n225 = ( n412 ) | ( n422 ) ;
 assign n224 = ( n226  &  n227  &  n12 ) | ( n226  &  n227  &  n225 ) ;
 assign n231 = ( n437  &  n61 ) | ( n15  &  n61 ) | ( n437  &  n501 ) | ( n15  &  n501 ) ;
 assign n229 = ( (~ i_9_) ) | ( n422 ) ;
 assign n230 = ( n396 ) | ( n421 ) ;
 assign n228 = ( n231  &  n229 ) | ( n231  &  n230 ) ;
 assign n234 = ( n229  &  n193 ) | ( n309  &  n193 ) | ( n229  &  n449 ) | ( n309  &  n449 ) ;
 assign n233 = ( n396 ) | ( n430 ) ;
 assign n232 = ( n234  &  n23 ) | ( n234  &  n233 ) ;
 assign n236 = ( n435  &  n8 ) | ( n56  &  n8 ) | ( n435  &  n260 ) | ( n56  &  n260 ) ;
 assign n237 = ( n4  &  n189 ) | ( n475  &  n189 ) | ( n4  &  n492 ) | ( n475  &  n492 ) ;
 assign n238 = ( n691  &  n690  &  n279 ) | ( n691  &  n690  &  n487 ) ;
 assign n239 = ( n694  &  n693  &  n4 ) | ( n694  &  n693  &  n460 ) ;
 assign n240 = ( n220  &  n224  &  n228  &  n232  &  n204  &  n213  &  n196  &  n698 ) ;
 assign n241 = ( n681  &  n149  &  n680  &  n679  &  n676  &  n675  &  n678  &  n689 ) ;
 assign n235 = ( n236  &  n237  &  n238  &  n239  &  n240  &  n241 ) ;
 assign n244 = ( n420  &  n71 ) | ( n221  &  n71 ) | ( n420  &  n516 ) | ( n221  &  n516 ) ;
 assign n243 = ( i_9_ ) | ( n430 ) ;
 assign n242 = ( n244  &  n243 ) | ( n244  &  n14 ) ;
 assign n246 = ( n61 ) | ( n527 ) ;
 assign n247 = ( n420 ) | ( n527 ) ;
 assign n248 = ( n417 ) | ( n457 ) ;
 assign n249 = ( n189 ) | ( n120 ) ;
 assign n250 = ( n226  &  n700  &  n279 ) | ( n226  &  n700  &  n509 ) ;
 assign n251 = ( n696  &  n61 ) | ( n696  &  n507 ) ;
 assign n252 = ( n293  &  n8 ) | ( n293  &  n419 ) ;
 assign n253 = ( n702  &  n701  &  n56 ) | ( n702  &  n701  &  n13 ) ;
 assign n245 = ( n246  &  n247  &  n248  &  n249  &  n250  &  n251  &  n252  &  n253 ) ;
 assign n255 = ( n189 ) | ( n459 ) ;
 assign n256 = ( n408 ) | ( n417 ) ;
 assign n257 = ( n71 ) | ( n502 ) ;
 assign n258 = ( n647  &  n436 ) | ( n647  &  n189 ) ;
 assign n254 = ( n130  &  n255  &  n232  &  n256  &  n257  &  n258 ) ;
 assign n261 = ( n8  &  n12 ) | ( n520  &  n12 ) | ( n8  &  n478 ) | ( n520  &  n478 ) ;
 assign n262 = ( n699  &  n189 ) | ( n699  &  n467 ) ;
 assign n260 = ( n434 ) | ( n441 ) ;
 assign n259 = ( n261  &  n262  &  n260 ) | ( n261  &  n262  &  n61 ) ;
 assign n265 = ( n15 ) | ( n457  &  n487 ) ;
 assign n266 = ( n667  &  n23 ) | ( n667  &  n454 ) ;
 assign n264 = ( n402 ) | ( n447 ) ;
 assign n263 = ( n265  &  n266  &  n243 ) | ( n265  &  n266  &  n264 ) ;
 assign n268 = ( n189 ) | ( n450 ) ;
 assign n269 = ( n71 ) | ( n514 ) ;
 assign n270 = ( n443  &  n243 ) | ( n467  &  n243 ) | ( n443  &  n524 ) | ( n467  &  n524 ) ;
 assign n271 = ( n436 ) | ( n23 ) ;
 assign n267 = ( n268  &  n269  &  n270  &  n271 ) ;
 assign n272 = ( n189  &  n417 ) | ( n528  &  n417 ) | ( n189  &  n510 ) | ( n528  &  n510 ) ;
 assign n273 = ( n730  &  n729  &  n61 ) | ( n730  &  n729  &  n497 ) ;
 assign n274 = ( n245  &  n254  &  n259  &  n263  &  n267  &  n220  &  n192  &  n161 ) ;
 assign n275 = ( n728  &  n727  &  n726  &  n725  &  n724  &  n723  &  n722  &  n721 ) ;
 assign n276 = ( n719  &  n720  &  n711  &  n713  &  n712  &  n718  &  n717  &  n715 ) ;
 assign n277 = ( n710  &  n709  &  n708  &  n707  &  n706  &  n705  &  n704  &  n703 ) ;
 assign n281 = ( n659  &  n189 ) | ( n659  &  n471 ) ;
 assign n282 = ( n440  &  n189 ) | ( n443  &  n189 ) | ( n440  &  n488 ) | ( n443  &  n488 ) ;
 assign n279 = ( i_9_ ) | ( n427 ) ;
 assign n280 = ( n391 ) | ( n414 ) ;
 assign n278 = ( n281  &  n282  &  n279 ) | ( n281  &  n282  &  n280 ) ;
 assign n284 = ( n23 ) | ( n484 ) ;
 assign n285 = ( n691  &  n614  &  n279 ) | ( n691  &  n614  &  n482 ) ;
 assign n286 = ( n734  &  n572  &  n162  &  n50  &  n51  &  n25 ) ;
 assign n287 = ( n450 ) | ( n61 ) ;
 assign n288 = ( n651  &  n630  &  n8 ) | ( n651  &  n630  &  n458 ) ;
 assign n289 = ( n732  &  n733  &  n420 ) | ( n732  &  n733  &  n62 ) ;
 assign n283 = ( n278  &  n284  &  n285  &  n286  &  n287  &  n206  &  n288  &  n289 ) ;
 assign n291 = ( n428 ) | ( n71 ) ;
 assign n292 = ( n189 ) | ( n458 ) ;
 assign n293 = ( n189 ) | ( n124 ) ;
 assign n294 = ( n71  &  n420 ) | ( n511  &  n420 ) | ( n71  &  n442 ) | ( n511  &  n442 ) ;
 assign n295 = ( n193 ) | ( n453 ) ;
 assign n296 = ( n636  &  n61 ) | ( n636  &  n230 ) ;
 assign n297 = ( n8  &  n193 ) | ( n463  &  n193 ) | ( n8  &  n518 ) | ( n463  &  n518 ) ;
 assign n298 = ( n731  &  n719  &  n243 ) | ( n731  &  n719  &  n465 ) ;
 assign n290 = ( n291  &  n292  &  n293  &  n294  &  n295  &  n296  &  n297  &  n298 ) ;
 assign n300 = ( n417 ) | ( n473 ) ;
 assign n301 = ( n23 ) | ( n470 ) ;
 assign n302 = ( n433 ) | ( n71 ) ;
 assign n303 = ( n243  &  n446 ) | ( n493  &  n446 ) | ( n243  &  n15 ) | ( n493  &  n15 ) ;
 assign n304 = ( n8  &  n420 ) | ( n508  &  n420 ) | ( n8  &  n519 ) | ( n508  &  n519 ) ;
 assign n305 = ( n443 ) | ( n519 ) ;
 assign n306 = ( n403  &  n443 ) | ( n189  &  n443 ) | ( n403  &  n501 ) | ( n189  &  n501 ) ;
 assign n307 = ( n229 ) | ( n471 ) ;
 assign n299 = ( n300  &  n301  &  n302  &  n303  &  n304  &  n305  &  n306  &  n307 ) ;
 assign n310 = ( n23 ) | ( n501 ) ;
 assign n311 = ( n15 ) | ( n173 ) ;
 assign n309 = ( n396 ) | ( n404 ) ;
 assign n308 = ( n310  &  n311  &  n23 ) | ( n310  &  n311  &  n309 ) ;
 assign n313 = ( n740  &  n739  &  n443 ) | ( n740  &  n739  &  n508 ) ;
 assign n314 = ( n583  &  n738  &  n229 ) | ( n583  &  n738  &  n460 ) ;
 assign n315 = ( n596  &  n737  &  n15 ) | ( n596  &  n737  &  n478 ) ;
 assign n316 = ( n736  &  n735  &  n15 ) | ( n736  &  n735  &  n264 ) ;
 assign n317 = ( n580  &  n246  &  n741  &  n744  &  n743  &  n746  &  n745  &  n747 ) ;
 assign n318 = ( n754  &  n602  &  n753  &  n752 ) ;
 assign n319 = ( n750  &  n751  &  n533  &  n543  &  n749  &  n748 ) ;
 assign n320 = ( n308  &  n267  &  n213  &  n188  &  n290  &  n299  &  n283  &  n757 ) ;
 assign n312 = ( n313  &  n314  &  n315  &  n316  &  n317  &  n318  &  n319  &  n320 ) ;
 assign n322 = ( n70 ) | ( n243 ) ;
 assign n323 = ( n443 ) | ( n74 ) ;
 assign n324 = ( n308  &  n440 ) | ( n308  &  n189 ) ;
 assign n325 = ( n4  &  n417 ) | ( n448  &  n417 ) | ( n4  &  n449 ) | ( n448  &  n449 ) ;
 assign n326 = ( n67  &  n564  &  n15 ) | ( n67  &  n564  &  n522 ) ;
 assign n327 = ( n287  &  n762  &  n229 ) | ( n287  &  n762  &  n492 ) ;
 assign n328 = ( n720  &  n761  &  n193 ) | ( n720  &  n761  &  n472 ) ;
 assign n321 = ( n269  &  n322  &  n323  &  n324  &  n325  &  n326  &  n327  &  n328 ) ;
 assign n330 = ( n61  &  n417 ) | ( n451  &  n417 ) | ( n61  &  n513 ) | ( n451  &  n513 ) ;
 assign n331 = ( n12 ) | ( n509 ) ;
 assign n332 = ( n403  &  n15 ) | ( n23  &  n15 ) | ( n403  &  n496 ) | ( n23  &  n496 ) ;
 assign n333 = ( n193 ) | ( n517 ) ;
 assign n334 = ( n760  &  n657  &  n71 ) | ( n760  &  n657  &  n112 ) ;
 assign n335 = ( n759  &  n742  &  n61 ) | ( n759  &  n742  &  n458 ) ;
 assign n329 = ( n330  &  n331  &  n332  &  n333  &  n334  &  n335 ) ;
 assign n337 = ( n417  &  n193 ) | ( n518  &  n193 ) | ( n417  &  n505 ) | ( n518  &  n505 ) ;
 assign n338 = ( n71 ) | ( n513 ) ;
 assign n339 = ( n12  &  n61 ) | ( n522  &  n61 ) | ( n12  &  n479 ) | ( n522  &  n479 ) ;
 assign n340 = ( n193  &  n4 ) | ( n522  &  n4 ) | ( n193  &  n124 ) | ( n522  &  n124 ) ;
 assign n341 = ( n23 ) | ( n483 ) ;
 assign n342 = ( n551  &  n417 ) | ( n551  &  n128 ) ;
 assign n336 = ( n337  &  n338  &  n339  &  n340  &  n341  &  n342 ) ;
 assign n344 = ( n782  &  n781  &  n436 ) | ( n782  &  n781  &  n443 ) ;
 assign n345 = ( n779  &  n778  &  n243 ) | ( n779  &  n778  &  n511 ) ;
 assign n346 = ( n329  &  n336  &  n321  &  n785  &  n55  &  n22  &  n81  &  n784 ) ;
 assign n347 = ( n776  &  n775  &  n260 ) | ( n776  &  n775  &  n189 ) ;
 assign n348 = ( n773  &  n772  &  n71 ) | ( n773  &  n772  &  n474 ) ;
 assign n349 = ( n769  &  n770  &  n768  &  n767  &  n766  &  n190  &  n765  &  n764 ) ;
 assign n343 = ( n344  &  n345  &  n346  &  n347  &  n348  &  n349 ) ;
 assign n351 = ( n443 ) | ( n425  &  n515 ) ;
 assign n352 = ( n229 ) | ( n488 ) ;
 assign n353 = ( n789  &  n23 ) | ( n789  &  n452 ) ;
 assign n354 = ( n790  &  n791  &  n71 ) | ( n790  &  n791  &  n482 ) ;
 assign n355 = ( n787  &  n788  &  n23 ) | ( n787  &  n788  &  n442 ) ;
 assign n356 = ( n740  &  n786  &  n12 ) | ( n740  &  n786  &  n465 ) ;
 assign n350 = ( n351  &  n352  &  n353  &  n354  &  n355  &  n356 ) ;
 assign n358 = ( n56 ) | ( n495 ) ;
 assign n359 = ( n189 ) | ( n477 ) ;
 assign n360 = ( n61 ) | ( n463 ) ;
 assign n361 = ( n69  &  n243 ) | ( n69  &  n500 ) ;
 assign n362 = ( n12 ) | ( n495 ) ;
 assign n363 = ( n8 ) | ( n124 ) ;
 assign n364 = ( n411 ) | ( n71 ) ;
 assign n365 = ( n577  &  n578  &  n420 ) | ( n577  &  n578  &  n501 ) ;
 assign n357 = ( n358  &  n359  &  n360  &  n361  &  n362  &  n363  &  n364  &  n365 ) ;
 assign n367 = ( n8  &  n193 ) | ( n309  &  n193 ) | ( n8  &  n428 ) | ( n309  &  n428 ) ;
 assign n368 = ( n15 ) | ( n435  &  n491 ) ;
 assign n369 = ( n792  &  n8 ) | ( n792  &  n415 ) ;
 assign n370 = ( n794  &  n443 ) | ( n794  &  n527 ) ;
 assign n371 = ( n793  &  n23 ) | ( n793  &  n479 ) ;
 assign n372 = ( n798  &  n799  &  n420 ) | ( n798  &  n799  &  n74 ) ;
 assign n373 = ( n797  &  n796  &  n243 ) | ( n797  &  n796  &  n489 ) ;
 assign n374 = ( n147  &  n111  &  n228  &  n808  &  n60  &  n809  &  n807  &  n803 ) ;
 assign n366 = ( n367  &  n368  &  n369  &  n370  &  n371  &  n372  &  n373  &  n374 ) ;
 assign n375 = ( n4 ) | ( n515 ) ;
 assign n376 = ( n56  &  n8 ) | ( n505  &  n8 ) | ( n56  &  n483 ) | ( n505  &  n483 ) ;
 assign n377 = ( n193  &  n71 ) | ( n435  &  n71 ) | ( n193  &  n499 ) | ( n435  &  n499 ) ;
 assign n378 = ( n283  &  n254  &  n224  &  n168  &  n357  &  n329  &  n242 ) ;
 assign n379 = ( n83  &  n587  &  n789  &  n830  &  n829  &  n828  &  n827  &  n826 ) ;
 assign n380 = ( n824  &  n545  &  n823  &  n821  &  n813  &  n812  &  n811  &  n817 ) ;
 assign n382 = ( n420  &  n56 ) | ( n169  &  n56 ) | ( n420  &  n514 ) | ( n169  &  n514 ) ;
 assign n383 = ( n419 ) | ( n61 ) ;
 assign n384 = ( n839  &  n536  &  n15 ) | ( n839  &  n536  &  n514 ) ;
 assign n385 = ( n702  &  n838  &  n71 ) | ( n702  &  n838  &  n498 ) ;
 assign n386 = ( n763  &  n837  &  n443 ) | ( n763  &  n837  &  n480 ) ;
 assign n387 = ( n836  &  n835  &  n279 ) | ( n836  &  n835  &  n449 ) ;
 assign n388 = ( n833  &  n832  &  n4 ) | ( n833  &  n832  &  n425 ) ;
 assign n389 = ( n95  &  n49  &  n142  &  n849  &  n848  &  n850  &  n847  &  n843 ) ;
 assign n381 = ( n382  &  n383  &  n384  &  n385  &  n386  &  n387  &  n388  &  n389 ) ;
 assign n391 = ( i_6_ ) | ( (~ i_7_) ) | ( i_8_ ) ;
 assign n396 = ( (~ i_3_) ) | ( i_4_ ) | ( (~ i_5_) ) ;
 assign n398 = ( (~ i_0_) ) | ( (~ i_1_) ) | ( (~ i_2_) ) ;
 assign n400 = ( n396 ) | ( n398 ) ;
 assign n402 = ( i_3_ ) | ( (~ i_4_) ) | ( i_5_ ) ;
 assign n403 = ( n398 ) | ( n402 ) ;
 assign n404 = ( (~ i_0_) ) | ( (~ i_1_) ) | ( i_2_ ) ;
 assign n406 = ( (~ i_3_) ) | ( (~ i_4_) ) | ( i_5_ ) ;
 assign n407 = ( (~ i_6_) ) | ( (~ i_7_) ) | ( i_8_ ) ;
 assign n408 = ( n406 ) | ( n407 ) ;
 assign n410 = ( (~ i_6_) ) | ( (~ i_7_) ) | ( (~ i_8_) ) ;
 assign n411 = ( n396 ) | ( n410 ) ;
 assign n412 = ( i_3_ ) | ( i_4_ ) | ( (~ i_5_) ) ;
 assign n413 = ( i_6_ ) | ( i_7_ ) | ( i_8_ ) ;
 assign n414 = ( i_3_ ) | ( i_4_ ) | ( i_5_ ) ;
 assign n415 = ( n404 ) | ( n414 ) ;
 assign n416 = ( (~ i_0_) ) | ( i_1_ ) | ( (~ i_2_) ) ;
 assign n417 = ( i_9_ ) | ( n416 ) ;
 assign n418 = ( (~ i_6_) ) | ( i_7_ ) | ( i_8_ ) ;
 assign n419 = ( n414 ) | ( n416 ) ;
 assign n420 = ( (~ i_9_) ) | ( n418 ) ;
 assign n421 = ( (~ i_0_) ) | ( i_1_ ) | ( i_2_ ) ;
 assign n422 = ( (~ i_6_) ) | ( i_7_ ) | ( (~ i_8_) ) ;
 assign n423 = ( (~ i_3_) ) | ( (~ i_4_) ) | ( (~ i_5_) ) ;
 assign n424 = ( n391 ) | ( n423 ) ;
 assign n425 = ( n412 ) | ( n421 ) ;
 assign n426 = ( n414 ) | ( n421 ) ;
 assign n427 = ( i_0_ ) | ( (~ i_1_) ) | ( (~ i_2_) ) ;
 assign n428 = ( n391 ) | ( n396 ) ;
 assign n429 = ( n412 ) | ( n418 ) ;
 assign n430 = ( i_0_ ) | ( (~ i_1_) ) | ( i_2_ ) ;
 assign n431 = ( (~ i_3_) ) | ( i_4_ ) | ( i_5_ ) ;
 assign n432 = ( i_6_ ) | ( (~ i_7_) ) | ( (~ i_8_) ) ;
 assign n433 = ( n431 ) | ( n432 ) ;
 assign n434 = ( i_3_ ) | ( (~ i_4_) ) | ( (~ i_5_) ) ;
 assign n435 = ( n410 ) | ( n434 ) ;
 assign n436 = ( n402 ) | ( n430 ) ;
 assign n437 = ( n402 ) | ( n422 ) ;
 assign n438 = ( i_0_ ) | ( i_1_ ) | ( (~ i_2_) ) ;
 assign n439 = ( n410 ) | ( n412 ) ;
 assign n440 = ( n414 ) | ( n438 ) ;
 assign n441 = ( i_0_ ) | ( i_1_ ) | ( i_2_ ) ;
 assign n442 = ( n431 ) | ( n441 ) ;
 assign n443 = ( (~ i_9_) ) | ( n413 ) ;
 assign n444 = ( n402 ) | ( n410 ) ;
 assign n445 = ( n412 ) | ( n441 ) ;
 assign n446 = ( n407 ) | ( n414 ) ;
 assign n447 = ( i_6_ ) | ( i_7_ ) | ( (~ i_8_) ) ;
 assign n448 = ( n398 ) | ( n431 ) ;
 assign n449 = ( n402 ) | ( n418 ) ;
 assign n450 = ( n398 ) | ( n412 ) ;
 assign n451 = ( n404 ) | ( n406 ) ;
 assign n452 = ( n404 ) | ( n434 ) ;
 assign n453 = ( n414 ) | ( n422 ) ;
 assign n454 = ( n406 ) | ( n421 ) ;
 assign n455 = ( n434 ) | ( n447 ) ;
 assign n456 = ( n402 ) | ( n432 ) ;
 assign n457 = ( n413 ) | ( n431 ) ;
 assign n458 = ( n406 ) | ( n438 ) ;
 assign n459 = ( n396 ) | ( n441 ) ;
 assign n460 = ( n396 ) | ( n416 ) ;
 assign n461 = ( n413 ) | ( n434 ) ;
 assign n462 = ( n406 ) | ( n410 ) ;
 assign n463 = ( n398 ) | ( n406 ) ;
 assign n464 = ( n398 ) | ( n434 ) ;
 assign n465 = ( n407 ) | ( n434 ) ;
 assign n466 = ( n404 ) | ( n412 ) ;
 assign n467 = ( n412 ) | ( n427 ) ;
 assign n468 = ( n396 ) | ( n407 ) ;
 assign n469 = ( n412 ) | ( n430 ) ;
 assign n470 = ( n434 ) | ( n438 ) ;
 assign n471 = ( n404 ) | ( n431 ) ;
 assign n472 = ( n396 ) | ( n447 ) ;
 assign n473 = ( n410 ) | ( n431 ) ;
 assign n474 = ( n422 ) | ( n434 ) ;
 assign n475 = ( n423 ) | ( n430 ) ;
 assign n476 = ( n410 ) | ( n414 ) ;
 assign n477 = ( n406 ) | ( n441 ) ;
 assign n478 = ( n412 ) | ( n447 ) ;
 assign n479 = ( n412 ) | ( n416 ) ;
 assign n480 = ( n430 ) | ( n434 ) ;
 assign n481 = ( n421 ) | ( n431 ) ;
 assign n482 = ( n423 ) | ( n432 ) ;
 assign n483 = ( n412 ) | ( n438 ) ;
 assign n484 = ( n402 ) | ( n421 ) ;
 assign n485 = ( n406 ) | ( n430 ) ;
 assign n486 = ( n416 ) | ( n434 ) ;
 assign n487 = ( n396 ) | ( n418 ) ;
 assign n488 = ( n423 ) | ( n441 ) ;
 assign n489 = ( n391 ) | ( n402 ) ;
 assign n490 = ( n402 ) | ( n404 ) ;
 assign n491 = ( n418 ) | ( n434 ) ;
 assign n492 = ( n396 ) | ( n438 ) ;
 assign n493 = ( n422 ) | ( n431 ) ;
 assign n494 = ( n391 ) | ( n406 ) ;
 assign n495 = ( n413 ) | ( n414 ) ;
 assign n496 = ( n414 ) | ( n432 ) ;
 assign n497 = ( n416 ) | ( n431 ) ;
 assign n498 = ( n406 ) | ( n432 ) ;
 assign n499 = ( n414 ) | ( n418 ) ;
 assign n500 = ( n432 ) | ( n434 ) ;
 assign n501 = ( n398 ) | ( n414 ) ;
 assign n502 = ( n418 ) | ( n423 ) ;
 assign n503 = ( n406 ) | ( n416 ) ;
 assign n504 = ( n423 ) | ( n438 ) ;
 assign n505 = ( n410 ) | ( n423 ) ;
 assign n506 = ( n407 ) | ( n423 ) ;
 assign n507 = ( n396 ) | ( n427 ) ;
 assign n508 = ( n421 ) | ( n423 ) ;
 assign n509 = ( n412 ) | ( n432 ) ;
 assign n510 = ( n406 ) | ( n422 ) ;
 assign n511 = ( n396 ) | ( n432 ) ;
 assign n512 = ( n418 ) | ( n431 ) ;
 assign n513 = ( n407 ) | ( n412 ) ;
 assign n514 = ( n407 ) | ( n431 ) ;
 assign n515 = ( n414 ) | ( n427 ) ;
 assign n516 = ( n391 ) | ( n434 ) ;
 assign n517 = ( n413 ) | ( n423 ) ;
 assign n518 = ( n402 ) | ( n407 ) ;
 assign n519 = ( n427 ) | ( n434 ) ;
 assign n520 = ( n430 ) | ( n431 ) ;
 assign n521 = ( n414 ) | ( n430 ) ;
 assign n522 = ( n406 ) | ( n413 ) ;
 assign n523 = ( n391 ) | ( n412 ) ;
 assign n524 = ( n406 ) | ( n418 ) ;
 assign n525 = ( n431 ) | ( n447 ) ;
 assign n526 = ( n427 ) | ( n431 ) ;
 assign n527 = ( n421 ) | ( n434 ) ;
 assign n528 = ( n404 ) | ( n423 ) ;
 assign n529 = ( n443 ) | ( n230 ) ;
 assign n530 = ( n420 ) | ( n485 ) ;
 assign n531 = ( n61 ) | ( n484 ) ;
 assign n532 = ( n403  &  n193 ) | ( n4  &  n193 ) | ( n403  &  n474 ) | ( n4  &  n474 ) ;
 assign n533 = ( n23 ) | ( n460 ) ;
 assign n534 = ( n417 ) | ( n474 ) ;
 assign n535 = ( n4  &  n193 ) | ( n309  &  n193 ) | ( n4  &  n465 ) | ( n309  &  n465 ) ;
 assign n536 = ( n437 ) | ( n56 ) ;
 assign n537 = ( n287  &  n311  &  n443 ) | ( n287  &  n311  &  n451 ) ;
 assign n538 = ( n295  &  n383  &  n4 ) | ( n295  &  n383  &  n452 ) ;
 assign n540 = ( n12 ) | ( n128 ) ;
 assign n541 = ( n61 ) | ( n454 ) ;
 assign n539 = ( n540  &  n541  &  n279 ) | ( n540  &  n541  &  n455 ) ;
 assign n542 = ( n23 ) | ( n448 ) ;
 assign n543 = ( n128 ) | ( n15 ) ;
 assign n544 = ( n279 ) | ( n456 ) ;
 assign n545 = ( n243 ) | ( n173 ) ;
 assign n546 = ( n408 ) | ( n56 ) ;
 assign n547 = ( n4 ) | ( n459 ) ;
 assign n548 = ( n400  &  n189 ) | ( n8  &  n189 ) | ( n400  &  n448 ) | ( n8  &  n448 ) ;
 assign n549 = ( n61  &  n8 ) | ( n464  &  n8 ) | ( n61  &  n403 ) | ( n464  &  n403 ) ;
 assign n551 = ( n193 ) | ( n411 ) ;
 assign n550 = ( n551  &  n408 ) | ( n551  &  n193 ) ;
 assign n552 = ( n229  &  n193 ) | ( n466  &  n193 ) | ( n229  &  n70 ) | ( n466  &  n70 ) ;
 assign n553 = ( n415  &  n417 ) | ( n420  &  n417 ) | ( n415  &  n491 ) | ( n420  &  n491 ) ;
 assign n555 = ( n70 ) | ( n417 ) ;
 assign n556 = ( n4 ) | ( n490 ) ;
 assign n554 = ( n553  &  n555  &  n552  &  n205  &  n550  &  n556  &  n549  &  n548 ) ;
 assign n558 = ( n66 ) | ( n12 ) ;
 assign n557 = ( n558  &  n198  &  n12 ) | ( n558  &  n198  &  n424 ) ;
 assign n559 = ( n8  &  n4 ) | ( n425  &  n4 ) | ( n8  &  n426 ) | ( n425  &  n426 ) ;
 assign n560 = ( n559  &  n420 ) | ( n559  &  n24 ) ;
 assign n561 = ( n279 ) | ( n428  &  n429 ) ;
 assign n563 = ( n243 ) | ( n435 ) ;
 assign n564 = ( n243 ) | ( n433 ) ;
 assign n562 = ( n563  &  n564  &  n243 ) | ( n563  &  n564  &  n474 ) ;
 assign n565 = ( n424 ) | ( n243 ) ;
 assign n566 = ( n436 ) | ( n4  &  n229 ) ;
 assign n567 = ( n243  &  n4 ) | ( n437  &  n4 ) | ( n243  &  n492 ) | ( n437  &  n492 ) ;
 assign n569 = ( n71 ) | ( n14 ) ;
 assign n568 = ( n569  &  n302  &  n71 ) | ( n569  &  n302  &  n173 ) ;
 assign n570 = ( n71  &  n440 ) | ( n439  &  n440 ) | ( n71  &  n23 ) | ( n439  &  n23 ) ;
 assign n572 = ( n444 ) | ( n56 ) ;
 assign n573 = ( n260 ) | ( n443 ) ;
 assign n571 = ( n572  &  n573  &  n429 ) | ( n572  &  n573  &  n56 ) ;
 assign n574 = ( n229 ) | ( n442 ) ;
 assign n575 = ( n12 ) | ( n457 ) ;
 assign n576 = ( n61 ) | ( n508 ) ;
 assign n577 = ( n439 ) | ( n15 ) ;
 assign n578 = ( n420 ) | ( n486 ) ;
 assign n579 = ( n12 ) | ( n505 ) ;
 assign n580 = ( n12 ) | ( n446 ) ;
 assign n581 = ( n61 ) | ( n233 ) ;
 assign n582 = ( n229 ) | ( n479 ) ;
 assign n583 = ( n417 ) | ( n194 ) ;
 assign n584 = ( n12 ) | ( n502 ) ;
 assign n585 = ( n279  &  n229 ) | ( n491  &  n229 ) | ( n279  &  n458 ) | ( n491  &  n458 ) ;
 assign n586 = ( n420 ) | ( n9 ) ;
 assign n587 = ( n411 ) | ( n417 ) ;
 assign n589 = ( n71 ) | ( n462 ) ;
 assign n588 = ( n589  &  n71 ) | ( n589  &  n465 ) ;
 assign n590 = ( n71 ) | ( n444 ) ;
 assign n591 = ( n530  &  n565  &  n15 ) | ( n530  &  n565  &  n502 ) ;
 assign n592 = ( n400 ) | ( n229 ) ;
 assign n594 = ( n193 ) | ( n437 ) ;
 assign n593 = ( n594  &  n420 ) | ( n594  &  n466 ) ;
 assign n596 = ( n189 ) | ( n501 ) ;
 assign n597 = ( n417 ) | ( n499 ) ;
 assign n595 = ( n596  &  n597  &  n189 ) | ( n596  &  n597  &  n451 ) ;
 assign n599 = ( n12 ) | ( n489 ) ;
 assign n598 = ( n599  &  n189 ) | ( n599  &  n484 ) ;
 assign n600 = ( n56 ) | ( n453 ) ;
 assign n601 = ( n193 ) | ( n424 ) ;
 assign n602 = ( n443 ) | ( n309 ) ;
 assign n603 = ( n420  &  n417 ) | ( n503  &  n417 ) | ( n420  &  n14 ) | ( n503  &  n14 ) ;
 assign n604 = ( n189 ) | ( n230 ) ;
 assign n605 = ( n12 ) | ( n472  &  n510 ) ;
 assign n606 = ( n363  &  n605  &  n417 ) | ( n363  &  n605  &  n495 ) ;
 assign n607 = ( n4  &  n12 ) | ( n481  &  n12 ) | ( n4  &  n439 ) | ( n481  &  n439 ) ;
 assign n608 = ( n229  &  n243 ) | ( n233  &  n243 ) | ( n229  &  n478 ) | ( n233  &  n478 ) ;
 assign n609 = ( n243  &  n4 ) | ( n57  &  n4 ) | ( n243  &  n9 ) | ( n57  &  n9 ) ;
 assign n610 = ( n71  &  n4 ) | ( n449  &  n4 ) | ( n71  &  n483 ) | ( n449  &  n483 ) ;
 assign n611 = ( n61  &  n4 ) | ( n459  &  n4 ) | ( n61  &  n442 ) | ( n459  &  n442 ) ;
 assign n612 = ( n56  &  n189 ) | ( n264  &  n189 ) | ( n56  &  n463 ) | ( n264  &  n463 ) ;
 assign n614 = ( n443 ) | ( n448 ) ;
 assign n613 = ( n614  &  n15 ) | ( n614  &  n476 ) ;
 assign n615 = ( n193 ) | ( n482 ) ;
 assign n616 = ( n193  &  n417 ) | ( n496  &  n417 ) | ( n193  &  n424 ) | ( n496  &  n424 ) ;
 assign n617 = ( n443  &  n8 ) | ( n62  &  n8 ) | ( n443  &  n460 ) | ( n62  &  n460 ) ;
 assign n618 = ( n8  &  n12 ) | ( n497  &  n12 ) | ( n8  &  n498 ) | ( n497  &  n498 ) ;
 assign n619 = ( n279 ) | ( n472  &  n478 ) ;
 assign n620 = ( n8  &  n243 ) | ( n480  &  n243 ) | ( n8  &  n499 ) | ( n480  &  n499 ) ;
 assign n621 = ( n189  &  n71 ) | ( n470  &  n71 ) | ( n189  &  n500 ) | ( n470  &  n500 ) ;
 assign n622 = ( n71 ) | ( n57 ) ;
 assign n623 = ( n61 ) | ( n221 ) ;
 assign n624 = ( n56  &  n229 ) | ( n516  &  n229 ) | ( n56  &  n445 ) | ( n516  &  n445 ) ;
 assign n625 = ( n127  &  n130  &  n123  &  n36  &  n3  &  n624 ) ;
 assign n626 = ( n417 ) | ( n435 ) ;
 assign n627 = ( n15 ) | ( n57 ) ;
 assign n628 = ( n243 ) | ( n280 ) ;
 assign n629 = ( n56 ) | ( n522 ) ;
 assign n630 = ( n420 ) | ( n483 ) ;
 assign n631 = ( n15 ) | ( n474  &  n494 ) ;
 assign n632 = ( n15  &  n229 ) | ( n456  &  n229 ) | ( n15  &  n501 ) | ( n456  &  n501 ) ;
 assign n634 = ( n23 ) | ( n451 ) ;
 assign n633 = ( n634  &  n420 ) | ( n634  &  n451 ) ;
 assign n636 = ( n193 ) | ( n513 ) ;
 assign n635 = ( n636  &  n61 ) | ( n636  &  n490 ) ;
 assign n637 = ( n193  &  n415 ) | ( n509  &  n415 ) | ( n193  &  n61 ) | ( n509  &  n61 ) ;
 assign n638 = ( n193  &  n417 ) | ( n57  &  n417 ) | ( n193  &  n517 ) | ( n57  &  n517 ) ;
 assign n640 = ( n417 ) | ( n465 ) ;
 assign n639 = ( n640  &  n443 ) | ( n640  &  n497 ) ;
 assign n642 = ( n443 ) | ( n124 ) ;
 assign n641 = ( n639  &  n642  &  n638  &  n637  &  n635  &  n633  &  n632  &  n631 ) ;
 assign n643 = ( n417  &  n12 ) | ( n446  &  n12 ) | ( n417  &  n14 ) | ( n446  &  n14 ) ;
 assign n644 = ( n12 ) | ( n491  &  n518 ) ;
 assign n645 = ( n12  &  n8 ) | ( n429  &  n8 ) | ( n12  &  n426 ) | ( n429  &  n426 ) ;
 assign n647 = ( n229 ) | ( n24 ) ;
 assign n646 = ( n647  &  n645  &  n279 ) | ( n647  &  n645  &  n517 ) ;
 assign n648 = ( n8  &  n243 ) | ( n5  &  n243 ) | ( n8  &  n498 ) | ( n5  &  n498 ) ;
 assign n649 = ( n23  &  n71 ) | ( n504  &  n71 ) | ( n23  &  n510 ) | ( n504  &  n510 ) ;
 assign n651 = ( n443 ) | ( n169 ) ;
 assign n650 = ( n651  &  n71 ) | ( n651  &  n494 ) ;
 assign n652 = ( n4  &  n8 ) | ( n508  &  n8 ) | ( n4  &  n484 ) | ( n508  &  n484 ) ;
 assign n653 = ( n425  &  n189 ) | ( n61  &  n189 ) | ( n425  &  n519 ) | ( n61  &  n519 ) ;
 assign n654 = ( n229  &  n243 ) | ( n5  &  n243 ) | ( n229  &  n505 ) | ( n5  &  n505 ) ;
 assign n655 = ( n243 ) | ( n444 ) ;
 assign n656 = ( n279  &  n189 ) | ( n128  &  n189 ) | ( n279  &  n507 ) | ( n128  &  n507 ) ;
 assign n657 = ( n420 ) | ( n488 ) ;
 assign n658 = ( n229  &  n420 ) | ( n120  &  n420 ) | ( n229  &  n460 ) | ( n120  &  n460 ) ;
 assign n659 = ( n279 ) | ( n518 ) ;
 assign n660 = ( n417 ) | ( n512 ) ;
 assign n661 = ( n411 ) | ( n15 ) ;
 assign n662 = ( n279 ) | ( n511 ) ;
 assign n663 = ( n243 ) | ( n473 ) ;
 assign n664 = ( n279 ) | ( n489 ) ;
 assign n665 = ( n189 ) | ( n464 ) ;
 assign n666 = ( n420  &  n4 ) | ( n454  &  n4 ) | ( n420  &  n526 ) | ( n454  &  n526 ) ;
 assign n667 = ( n4 ) | ( n469 ) ;
 assign n669 = ( n15 ) | ( n509 ) ;
 assign n668 = ( n669  &  n4 ) | ( n669  &  n471 ) ;
 assign n671 = ( n23 ) | ( n475 ) ;
 assign n670 = ( n671  &  n668  &  n23 ) | ( n671  &  n668  &  n508 ) ;
 assign n673 = ( n443 ) | ( n521 ) ;
 assign n672 = ( n673  &  n604  &  n243 ) | ( n673  &  n604  &  n516 ) ;
 assign n674 = ( n8  &  n189 ) | ( n504  &  n189 ) | ( n8  &  n490 ) | ( n504  &  n490 ) ;
 assign n675 = ( n15  &  n443 ) | ( n499  &  n443 ) | ( n15  &  n490 ) | ( n499  &  n490 ) ;
 assign n676 = ( n23  &  n12 ) | ( n486  &  n12 ) | ( n23  &  n468 ) | ( n486  &  n468 ) ;
 assign n677 = ( n12  &  n425 ) | ( n525  &  n425 ) | ( n12  &  n23 ) | ( n525  &  n23 ) ;
 assign n678 = ( n362  &  n677  &  n408 ) | ( n362  &  n677  &  n279 ) ;
 assign n679 = ( n229  &  n8 ) | ( n526  &  n8 ) | ( n229  &  n519 ) | ( n526  &  n519 ) ;
 assign n680 = ( n151  &  n61 ) | ( n151  &  n475 ) ;
 assign n681 = ( n243  &  n420 ) | ( n13  &  n420 ) | ( n243  &  n233 ) | ( n13  &  n233 ) ;
 assign n682 = ( n229  &  n61 ) | ( n504  &  n61 ) | ( n229  &  n169 ) | ( n504  &  n169 ) ;
 assign n683 = ( n71  &  n229 ) | ( n457  &  n229 ) | ( n71  &  n9 ) | ( n457  &  n9 ) ;
 assign n684 = ( n600  &  n56 ) | ( n600  &  n499 ) ;
 assign n685 = ( n15  &  n193 ) | ( n112  &  n193 ) | ( n15  &  n429 ) | ( n112  &  n429 ) ;
 assign n686 = ( n443  &  n417 ) | ( n503  &  n417 ) | ( n443  &  n511 ) | ( n503  &  n511 ) ;
 assign n687 = ( n189  &  n417 ) | ( n497  &  n417 ) | ( n189  &  n496 ) | ( n497  &  n496 ) ;
 assign n688 = ( n687  &  n417 ) | ( n687  &  n280 ) ;
 assign n689 = ( n531  &  n32  &  n684  &  n683  &  n682  &  n686  &  n685  &  n688 ) ;
 assign n690 = ( n23  &  n279 ) | ( n526  &  n279 ) | ( n23  &  n493 ) | ( n526  &  n493 ) ;
 assign n691 = ( n12 ) | ( n496 ) ;
 assign n692 = ( n323  &  n70 ) | ( n323  &  n56 ) ;
 assign n693 = ( n601  &  n692  &  n15 ) | ( n601  &  n692  &  n524 ) ;
 assign n694 = ( n61  &  n243 ) | ( n24  &  n243 ) | ( n61  &  n453 ) | ( n24  &  n453 ) ;
 assign n696 = ( n279 ) | ( n516 ) ;
 assign n695 = ( n696  &  n411 ) | ( n696  &  n12 ) ;
 assign n697 = ( n4  &  n189 ) | ( n521  &  n189 ) | ( n4  &  n475 ) | ( n521  &  n475 ) ;
 assign n698 = ( n176  &  n88  &  n73  &  n7  &  n697  &  n695 ) ;
 assign n699 = ( n229  &  n12 ) | ( n451  &  n12 ) | ( n229  &  n487 ) | ( n451  &  n487 ) ;
 assign n700 = ( n23  &  n243 ) | ( n480  &  n243 ) | ( n23  &  n523 ) | ( n480  &  n523 ) ;
 assign n701 = ( n15  &  n417 ) | ( n525  &  n417 ) | ( n15  &  n498 ) | ( n525  &  n498 ) ;
 assign n702 = ( n23 ) | ( n458 ) ;
 assign n703 = ( n420  &  n23 ) | ( n120  &  n23 ) | ( n420  &  n463 ) | ( n120  &  n463 ) ;
 assign n704 = ( n400  &  n420 ) | ( n189  &  n420 ) | ( n400  &  n464 ) | ( n189  &  n464 ) ;
 assign n705 = ( n403  &  n15 ) | ( n229  &  n15 ) | ( n403  &  n489 ) | ( n229  &  n489 ) ;
 assign n706 = ( n528 ) | ( n4  &  n229 ) ;
 assign n707 = ( n193 ) | ( n468  &  n524 ) ;
 assign n708 = ( n420  &  n4 ) | ( n471  &  n4 ) | ( n420  &  n497 ) | ( n471  &  n497 ) ;
 assign n709 = ( n579  &  n417 ) | ( n579  &  n509 ) ;
 assign n710 = ( n576  &  n443 ) | ( n576  &  n481 ) ;
 assign n711 = ( n8  &  n12 ) | ( n527  &  n12 ) | ( n8  &  n516 ) | ( n527  &  n516 ) ;
 assign n712 = ( n158  &  n279 ) | ( n158  &  n112 ) ;
 assign n713 = ( n279 ) | ( n225  &  n500 ) ;
 assign n714 = ( n279  &  n411 ) | ( n495  &  n411 ) | ( n279  &  n243 ) | ( n495  &  n243 ) ;
 assign n716 = ( n71 ) | ( n505 ) ;
 assign n715 = ( n716  &  n714  &  n243 ) | ( n716  &  n714  &  n456 ) ;
 assign n717 = ( n71  &  n229 ) | ( n517  &  n229 ) | ( n71  &  n470 ) | ( n517  &  n470 ) ;
 assign n718 = ( n443  &  n229 ) | ( n9  &  n229 ) | ( n443  &  n74 ) | ( n9  &  n74 ) ;
 assign n719 = ( n425 ) | ( n189 ) ;
 assign n720 = ( n443 ) | ( n484 ) ;
 assign n721 = ( n358  &  n229 ) | ( n358  &  n131 ) ;
 assign n722 = ( n15  &  n400 ) | ( n505  &  n400 ) | ( n15  &  n4 ) | ( n505  &  n4 ) ;
 assign n723 = ( n429  &  n193 ) | ( n15  &  n193 ) | ( n429  &  n502 ) | ( n15  &  n502 ) ;
 assign n724 = ( n417 ) | ( n476  &  n493 ) ;
 assign n725 = ( n662  &  n8 ) | ( n662  &  n475 ) ;
 assign n726 = ( n243  &  n189 ) | ( n522  &  n189 ) | ( n243  &  n504 ) | ( n522  &  n504 ) ;
 assign n727 = ( n229  &  n8 ) | ( n169  &  n8 ) | ( n229  &  n477 ) | ( n169  &  n477 ) ;
 assign n728 = ( n594  &  n415 ) | ( n594  &  n229 ) ;
 assign n729 = ( n243  &  n189 ) | ( n518  &  n189 ) | ( n243  &  n483 ) | ( n518  &  n483 ) ;
 assign n730 = ( n189 ) | ( n503 ) ;
 assign n731 = ( n189 ) | ( n233 ) ;
 assign n732 = ( n15  &  n193 ) | ( n453  &  n193 ) | ( n15  &  n487 ) | ( n453  &  n487 ) ;
 assign n733 = ( n576  &  n166  &  n417 ) | ( n576  &  n166  &  n429 ) ;
 assign n734 = ( n443 ) | ( n452 ) ;
 assign n735 = ( n15  &  n229 ) | ( n512  &  n229 ) | ( n15  &  n464 ) | ( n512  &  n464 ) ;
 assign n736 = ( n403 ) | ( n61 ) ;
 assign n737 = ( n193 ) | ( n510  &  n511 ) ;
 assign n738 = ( n193  &  n415 ) | ( n523  &  n415 ) | ( n193  &  n189 ) | ( n523  &  n189 ) ;
 assign n739 = ( n417  &  n8 ) | ( n264  &  n8 ) | ( n417  &  n479 ) | ( n264  &  n479 ) ;
 assign n740 = ( n229 ) | ( n527 ) ;
 assign n742 = ( n12 ) | ( n453 ) ;
 assign n741 = ( n742  &  n426 ) | ( n742  &  n229 ) ;
 assign n743 = ( n420  &  n279 ) | ( n426  &  n279 ) | ( n420  &  n506 ) | ( n426  &  n506 ) ;
 assign n744 = ( n443  &  n279 ) | ( n221  &  n279 ) | ( n443  &  n474 ) | ( n221  &  n474 ) ;
 assign n745 = ( n90  &  n189 ) | ( n90  &  n515 ) ;
 assign n746 = ( n243 ) | ( n128  &  n487 ) ;
 assign n747 = ( n581  &  n589  &  n4 ) | ( n581  &  n589  &  n520 ) ;
 assign n748 = ( n8  &  n56 ) | ( n492  &  n56 ) | ( n8  &  n517 ) | ( n492  &  n517 ) ;
 assign n749 = ( n56  &  n189 ) | ( n498  &  n189 ) | ( n56  &  n131 ) | ( n498  &  n131 ) ;
 assign n750 = ( n193 ) | ( n500 ) ;
 assign n751 = ( n193 ) | ( n506 ) ;
 assign n752 = ( n12 ) | ( n449  &  n524 ) ;
 assign n753 = ( n4  &  n61 ) | ( n507  &  n61 ) | ( n4  &  n467 ) | ( n507  &  n467 ) ;
 assign n754 = ( n71 ) | ( n476  &  n525 ) ;
 assign n755 = ( n193  &  n417 ) | ( n498  &  n417 ) | ( n193  &  n523 ) | ( n498  &  n523 ) ;
 assign n756 = ( n12  &  n420 ) | ( n444  &  n420 ) | ( n12  &  n5 ) | ( n444  &  n5 ) ;
 assign n758 = ( n229 ) | ( n515 ) ;
 assign n757 = ( n154  &  n115  &  n43  &  n758  &  n756  &  n755 ) ;
 assign n759 = ( n279 ) | ( n457 ) ;
 assign n760 = ( n417 ) | ( n500 ) ;
 assign n761 = ( n661  &  n634  &  n4 ) | ( n661  &  n634  &  n464 ) ;
 assign n763 = ( n420 ) | ( n480 ) ;
 assign n762 = ( n763  &  n716  &  n8 ) | ( n763  &  n716  &  n467 ) ;
 assign n764 = ( n15  &  n400 ) | ( n498  &  n400 ) | ( n15  &  n23 ) | ( n498  &  n23 ) ;
 assign n765 = ( n229  &  n193 ) | ( n450  &  n193 ) | ( n229  &  n433 ) | ( n450  &  n433 ) ;
 assign n766 = ( n443  &  n193 ) | ( n471  &  n193 ) | ( n443  &  n516 ) | ( n471  &  n516 ) ;
 assign n767 = ( n61  &  n417 ) | ( n503  &  n417 ) | ( n61  &  n456 ) | ( n503  &  n456 ) ;
 assign n768 = ( n4  &  n419 ) | ( n479  &  n419 ) | ( n4  &  n189 ) | ( n479  &  n189 ) ;
 assign n769 = ( n8  &  n189 ) | ( n481  &  n189 ) | ( n8  &  n527 ) | ( n481  &  n527 ) ;
 assign n770 = ( n426 ) | ( n61 ) ;
 assign n771 = ( n8  &  n428 ) | ( n485  &  n428 ) | ( n8  &  n243 ) | ( n485  &  n243 ) ;
 assign n772 = ( n156  &  n771  &  n12 ) | ( n156  &  n771  &  n57 ) ;
 assign n773 = ( n469 ) | ( n23  &  n229 ) ;
 assign n774 = ( n61  &  n71 ) | ( n483  &  n71 ) | ( n61  &  n280 ) | ( n483  &  n280 ) ;
 assign n775 = ( n774  &  n56 ) | ( n774  &  n194 ) ;
 assign n776 = ( n56 ) | ( n472  &  n510 ) ;
 assign n777 = ( n540  &  n56 ) | ( n540  &  n518 ) ;
 assign n778 = ( n750  &  n777  &  n15 ) | ( n750  &  n777  &  n523 ) ;
 assign n779 = ( n734  &  n229 ) | ( n734  &  n497 ) ;
 assign n780 = ( n71  &  n229 ) | ( n493  &  n229 ) | ( n71  &  n507 ) | ( n493  &  n507 ) ;
 assign n781 = ( n673  &  n780  &  n243 ) | ( n673  &  n780  &  n512 ) ;
 assign n782 = ( n4  &  n243 ) | ( n485  &  n243 ) | ( n4  &  n472 ) | ( n485  &  n472 ) ;
 assign n783 = ( n8  &  n56 ) | ( n169  &  n56 ) | ( n8  &  n280 ) | ( n169  &  n280 ) ;
 assign n784 = ( n11  &  n783  &  n420 ) | ( n11  &  n783  &  n458 ) ;
 assign n785 = ( n204  &  n172  &  n245 ) ;
 assign n786 = ( n640  &  n736  &  n61 ) | ( n640  &  n736  &  n481 ) ;
 assign n787 = ( n23  &  n440 ) | ( n485  &  n440 ) | ( n23  &  n61 ) | ( n485  &  n61 ) ;
 assign n788 = ( n29  &  n189 ) | ( n29  &  n452 ) ;
 assign n789 = ( n400 ) | ( n420 ) ;
 assign n790 = ( n730  &  n193 ) | ( n730  &  n446 ) ;
 assign n791 = ( n443  &  n408 ) | ( n120  &  n408 ) | ( n443  &  n15 ) | ( n120  &  n15 ) ;
 assign n792 = ( n193  &  n8 ) | ( n514  &  n8 ) | ( n193  &  n466 ) | ( n514  &  n466 ) ;
 assign n793 = ( n417 ) | ( n444  &  n505 ) ;
 assign n794 = ( n12 ) | ( n112  &  n511 ) ;
 assign n795 = ( n425  &  n426 ) | ( n229  &  n426 ) | ( n425  &  n443 ) | ( n229  &  n443 ) ;
 assign n796 = ( n795  &  n424 ) | ( n795  &  n279 ) ;
 assign n797 = ( n279  &  n243 ) | ( n510  &  n243 ) | ( n279  &  n462 ) | ( n510  &  n462 ) ;
 assign n798 = ( n23  &  n229 ) | ( n492  &  n229 ) | ( n23  &  n459 ) | ( n492  &  n459 ) ;
 assign n799 = ( n40  &  n34  &  n420 ) | ( n40  &  n34  &  n131 ) ;
 assign n800 = ( n443  &  n448 ) | ( n463  &  n448 ) | ( n443  &  n61 ) | ( n463  &  n61 ) ;
 assign n801 = ( n669  &  n800  &  n420 ) | ( n669  &  n800  &  n490 ) ;
 assign n802 = ( n23  &  n4 ) | ( n497  &  n4 ) | ( n23  &  n454 ) | ( n497  &  n454 ) ;
 assign n803 = ( n802  &  n801  &  n12 ) | ( n802  &  n801  &  n512 ) ;
 assign n805 = ( n61 ) | ( n480 ) ;
 assign n804 = ( n805  &  n671  &  n23 ) | ( n805  &  n671  &  n521 ) ;
 assign n806 = ( n56  &  n417 ) | ( n476  &  n417 ) | ( n56  &  n524 ) | ( n476  &  n524 ) ;
 assign n807 = ( n806  &  n804  &  n229 ) | ( n806  &  n804  &  n486 ) ;
 assign n808 = ( n408  &  n14 ) | ( n243  &  n14 ) | ( n408  &  n56 ) | ( n243  &  n56 ) ;
 assign n809 = ( n357  &  n321  &  n350  &  n278  &  n263  &  n299 ) ;
 assign n810 = ( n443  &  n15 ) | ( n464  &  n15 ) | ( n443  &  n495 ) | ( n464  &  n495 ) ;
 assign n811 = ( n665  &  n810  &  n424 ) | ( n665  &  n810  &  n15 ) ;
 assign n812 = ( n193  &  n61 ) | ( n13  &  n61 ) | ( n193  &  n471 ) | ( n13  &  n471 ) ;
 assign n813 = ( n443  &  n417 ) | ( n466  &  n417 ) | ( n443  &  n482 ) | ( n466  &  n482 ) ;
 assign n814 = ( n4  &  n417 ) | ( n503  &  n417 ) | ( n4  &  n13 ) | ( n503  &  n13 ) ;
 assign n815 = ( n626  &  n814  &  n419 ) | ( n626  &  n814  &  n229 ) ;
 assign n816 = ( n584  &  n12 ) | ( n584  &  n455 ) ;
 assign n817 = ( n816  &  n815  &  n279 ) | ( n816  &  n815  &  n502 ) ;
 assign n818 = ( n243  &  n189 ) | ( n112  &  n189 ) | ( n243  &  n480 ) | ( n112  &  n480 ) ;
 assign n819 = ( n664  &  n818  &  n443 ) | ( n664  &  n818  &  n233 ) ;
 assign n820 = ( n436  &  n243 ) | ( n61  &  n243 ) | ( n436  &  n439 ) | ( n61  &  n439 ) ;
 assign n821 = ( n820  &  n819  &  n420 ) | ( n820  &  n819  &  n469 ) ;
 assign n822 = ( n628  &  n71 ) | ( n628  &  n194 ) ;
 assign n823 = ( n590  &  n822  &  n420 ) | ( n590  &  n822  &  n492 ) ;
 assign n824 = ( n4 ) | ( n440  &  n445 ) ;
 assign n825 = ( n23  &  n417 ) | ( n471  &  n417 ) | ( n23  &  n487 ) | ( n471  &  n487 ) ;
 assign n826 = ( n546  &  n825  &  n15 ) | ( n546  &  n825  &  n13 ) ;
 assign n827 = ( n61  &  n189 ) | ( n486  &  n189 ) | ( n61  &  n221 ) | ( n486  &  n221 ) ;
 assign n828 = ( n8 ) | ( n24  &  n221 ) ;
 assign n829 = ( n411  &  n420 ) | ( n279  &  n420 ) | ( n411  &  n521 ) | ( n279  &  n521 ) ;
 assign n830 = ( n592  &  n443 ) | ( n592  &  n445 ) ;
 assign n831 = ( n15  &  n417 ) | ( n468  &  n417 ) | ( n15  &  n516 ) | ( n468  &  n516 ) ;
 assign n832 = ( n247  &  n831  &  n12 ) | ( n247  &  n831  &  n433 ) ;
 assign n833 = ( n599  &  n12 ) | ( n599  &  n456 ) ;
 assign n834 = ( n12  &  n66 ) | ( n280  &  n66 ) | ( n12  &  n279 ) | ( n280  &  n279 ) ;
 assign n835 = ( n834  &  n279 ) | ( n834  &  n473 ) ;
 assign n836 = ( n279  &  n229 ) | ( n525  &  n229 ) | ( n279  &  n519 ) | ( n525  &  n519 ) ;
 assign n837 = ( n443  &  n189 ) | ( n475  &  n189 ) | ( n443  &  n485 ) | ( n475  &  n485 ) ;
 assign n838 = ( n8 ) | ( n436 ) ;
 assign n839 = ( n15 ) | ( n517 ) ;
 assign n840 = ( n528 ) | ( n8  &  n23 ) ;
 assign n841 = ( n760  &  n840  &  n193 ) | ( n760  &  n840  &  n489 ) ;
 assign n842 = ( n23 ) | ( n124  &  n230 ) ;
 assign n843 = ( n842  &  n841  &  n12 ) | ( n842  &  n841  &  n493 ) ;
 assign n844 = ( n420  &  n23 ) | ( n481  &  n23 ) | ( n420  &  n519 ) | ( n481  &  n519 ) ;
 assign n845 = ( n844  &  n71 ) | ( n844  &  n524 ) ;
 assign n846 = ( n71  &  n443 ) | ( n491  &  n443 ) | ( n71  &  n470 ) | ( n491  &  n470 ) ;
 assign n847 = ( n846  &  n845  &  n429 ) | ( n846  &  n845  &  n71 ) ;
 assign n848 = ( n443  &  n417 ) | ( n5  &  n417 ) | ( n443  &  n462 ) | ( n5  &  n462 ) ;
 assign n849 = ( n229  &  n417 ) | ( n475  &  n417 ) | ( n229  &  n455 ) | ( n475  &  n455 ) ;
 assign n850 = ( n350  &  n336  &  n242  &  n259  &  n196  &  n290 ) ;


endmodule

