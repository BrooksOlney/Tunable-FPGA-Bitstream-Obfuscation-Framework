`timescale 10ns/1ns
module TOP (/* input clk, */ input i_0_, input i_1_, input i_2_, input i_3_, input i_4_, input i_5_, input i_6_, input i_7_, input i_8_, input i_9_, input i_10_, input i_11_, input i_12_, input i_13_output wire o_0_, output wire o_1_, output wire o_2_, output wire o_3_, output wire o_4_, output wire o_5_, output wire o_6_, output wire o_7_);

//reg [13:0] inputs;
//reg [7:0] outputs;
//always @(posedge clk) inputs = {i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_};
//always @(posedge clk) outputs = {o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_};

	wire n19, n636, n627, n611, n18, n10, n11, n12, n14, n16, n817;
	wire n819, n820, n9, n1, n2, n3, n5, n8, n717, n791, n792;
	wire n177, n180, n182, n50, n522, n264, n296, n776, n47, n771, n773;
	wire n267, n270, n275, n279, n283, n288, n782, n783, n328, n332, n333;
	wire n317, n445, n807, n448, n326, n61, n666, n701, n806, n42, n334;
	wire n804, n574, n577, n585, n596, n597, n599, n600, n601, n23, n641;
	wire n640, n21, n24, n542, n53, n39, n125, n655, n35, n557, n118;
	wire n33, n31, n32, n247, n36, n233, n38, n40, n43, n45, n46;
	wire n471, n763, n653, n174, n497, n765, n223, n57, n421, n63, n73;
	wire n364, n65, n99, n74, n216, n77, n78, n69, n72, n778, n58;
	wire n197, n196, n406, n650, n656, n62, n79, n83, n84, n85, n87;
	wire n88, n144, n98, n173, n91, n90, n101, n654, n652, n93, n94;
	wire n102, n108, n96, n95, n453, n104, n757, n185, n106, n107, n114;
	wire n110, n111, n113, n376, n116, n181, n684, n685, n749, n649, n124;
	wire n268, n748, n692, n693, n690, n691, n220, n287, n565, n383, n658;
	wire n123, n681, n683, n127, n132, n133, n134, n135, n136, n138, n139;
	wire n499, n164, n688, n188, n165, n746, n747, n682, n687, n146, n147;
	wire n145, n149, n151, n241, n686, n179, n217, n680, n157, n158, n159;
	wire n160, n161, n162, n744, n745, n222, n315, n166, n167, n189, n742;
	wire n743, n677, n170, n171, n178, n172, n175, n186, n675, n559, n673;
	wire n548, n190, n191, n193, n194, n195, n578, n582, n738, n740, n667;
	wire n201, n202, n199, n481, n409, n669, n668, n206, n204, n205, n402;
	wire n670, n671, n672, n602, n210, n211, n209, n214, n236, n219, n226;
	wire n945, n651, n229, n230, n225, n228, n234, n238, n239, n242, n237;
	wire n240, n248, n249, n246, n252, n255, n604, n257, n696, n259, n260;
	wire n775, n261, n256, n506, n89, n271, n720, n148, n152, n276, n659;
	wire n479, n212, n280, n723, n662, n726, n730, n732, n734, n198, n203;
	wire n207, n759, n761, n762, n302, n303, n306, n307, n384, n304, n308;
	wire n698, n301, n311, n915, n313, n314, n318, n323, n324, n322, n339;
	wire n316, n695, n794, n327, n312, n330, n331, n946, n802, n803, n309;
	wire n335, n398, n657, n920, n337, n338, n341, n340, n344, n346, n342;
	wire n345, n349, n348, n704, n705, n352, n351, n353, n951, n354, n719;
	wire n357, n362, n365, n674, n367, n718, n347, n350, n360, n363, n366;
	wire n816, n370, n336, n371, n372, n373, n664, n380, n381, n377, n702;
	wire n382, n387, n388, n389, n390, n391, n626, n697, n379, n385, n393;
	wire n394, n648, n396, n397, n403, n809, n399, n401, n921, n500, n433;
	wire n700, n395, n404, n408, n411, n412, n415, n417, n488, n813, n814;
	wire n416, n419, n424, n426, n713, n647, n451, n455, n454, n712, n109;
	wire n449, n452, n457, n458, n460, n461, n462, n927, n703, n923, n463;
	wire n852, n467, n468, n105, n470, n552, n851, n478, n480, n485, n483;
	wire n490, n492, n493, n489, n429, n476, n901, n835, n502, n504, n508;
	wire n529, n834, n833, n513, n514, n517, n518, n521, n524, n520, n507;
	wire n511, n515, n76, n519, n832, n523, n830, n525, n528, n532, n533;
	wire n534, n535, n537, n538, n56, n235, n541, n708, n551, n553, n556;
	wire n848, n849, n568, n570, n572, n573, n575, n823, n709, n824, n584;
	wire n825, n710, n826, n711, n827, n547, n543, n550, n564, n581, n874;
	wire n872, n567, n871, n869, n571, n876, n878, n879, n882, n884, n885;
	wire n932, n933, n736, n603, n896, n607, n608, n437, n942, n606, n714;
	wire n232, n898, n899, n894, n891, n539, n540, n612, n613, n614, n615;
	wire n616, n617, n620, n619, n943, n944, n622, n624, n618, n621, n41;
	wire n905, n909, n900, n904, n908, n906, n250, n628, n629, n630, n631;
	wire n633, n632, n635, n910, n911, n637, n638, n639, n487, n660, n112;
	wire n82, n912, n722, n725, n251, n661, n727, n231, n243, n728, n20;
	wire n224, n227, n733, n663, n218, n215, n221, n428, n168, n140, n665;
	wire n751, n115, n750, n752, n119, n754, n92, n97, n100, n758, n44;
	wire n764, n766, n37, n768, n26, n767, n30, n34, n716, n772, n51;
	wire n769, n770, n777, n258, n779, n253, n781, n780, n192, n292, n785;
	wire n187, n169, n788, n163, n156, n143, n790, n789, n131, n297, n753;
	wire n755, n320, n914, n796, n799, n795, n797, n916, n805, n425, n808;
	wire n810, n812, n699, n818, n434, n410, n422, n369, n392, n430, n821;
	wire n822, n934, n838, n496, n495, n841, n494, n844, n486, n843, n845;
	wire n491, n482, n857, n469, n472, n856, n922, n863, n862, n456, n466;
	wire n867, n930, n870, n707, n873, n569, n588, n828, n829, n554, n591;
	wire n592, n531, n886, n940, n609, n890, n895, n893, n610, n903, n902;
	wire n625, n623, n798, n854, n558, n561, n858, n861, n865, n840, n837;
	wire n498, n646, n846, n847, n935, n937, n941;


	lut_sub lut_0 ({n19}, o_0_);
	defparam lut_0.LUT_SIZE = 1;
	defparam lut_0.mask = 2'b01;

	lut_sub lut_1 ({n636}, o_1_);
	defparam lut_1.LUT_SIZE = 1;
	defparam lut_1.mask = 2'b01;

	lut_sub lut_2 ({n627}, o_2_);
	defparam lut_2.LUT_SIZE = 1;
	defparam lut_2.mask = 2'b01;

	lut_sub lut_3 ({n611}, o_3_);
	defparam lut_3.LUT_SIZE = 1;
	defparam lut_3.mask = 2'b01;

	lut_sub lut_4 ({n18}, o_4_);
	defparam lut_4.LUT_SIZE = 1;
	defparam lut_4.mask = 2'b01;

	lut_sub lut_5 ({n10, n11, n12, n14, n16, n817, n819, n820}, o_5_);
	defparam lut_5.LUT_SIZE = 8;
	defparam lut_5.mask = 256'HFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F;

	lut_sub lut_6 ({n9}, o_6_);
	defparam lut_6.LUT_SIZE = 1;
	defparam lut_6.mask = 2'b01;

	lut_sub lut_7 ({n1, n2, n3, n5, n8, n717, n791, n792}, o_7_);
	defparam lut_7.LUT_SIZE = 8;
	defparam lut_7.mask = 256'HFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F;

	lut_sub lut_8 ({i_9_, n177, n180, n182}, n1);
	defparam lut_8.LUT_SIZE = 4;
	defparam lut_8.mask = 16'H00EF;

	lut_sub lut_9 ({n50, n522, i_9_}, n2);
	defparam lut_9.LUT_SIZE = 3;
	defparam lut_9.mask = 8'H80;

	lut_sub lut_10 ({i_5_, n264, n296, n776}, n3);
	defparam lut_10.LUT_SIZE = 4;
	defparam lut_10.mask = 16'H005D;

	lut_sub lut_11 ({i_9_, n47, n771, n773}, n5);
	defparam lut_11.LUT_SIZE = 4;
	defparam lut_11.mask = 16'HF700;

	lut_sub lut_12 ({n267, n270, n275, n279, n283, n288, n782, n783}, n8);
	defparam lut_12.LUT_SIZE = 8;
	defparam lut_12.mask = 256'HFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7;

	lut_sub lut_13 ({i_2_, n328, n332, n333}, n9);
	defparam lut_13.LUT_SIZE = 4;
	defparam lut_13.mask = 16'H8088;

	lut_sub lut_14 ({i_11_, n317, n445, n807}, n10);
	defparam lut_14.LUT_SIZE = 4;
	defparam lut_14.mask = 16'H5D00;

	lut_sub lut_15 ({n448, n326, i_2_}, n11);
	defparam lut_15.LUT_SIZE = 3;
	defparam lut_15.mask = 8'H80;

	lut_sub lut_16 ({n61, n666}, n12);
	defparam lut_16.LUT_SIZE = 2;
	defparam lut_16.mask = 4'b0001;

	lut_sub lut_17 ({i_13_, n666, n701, n806}, n14);
	defparam lut_17.LUT_SIZE = 4;
	defparam lut_17.mask = 16'H1113;

	lut_sub lut_18 ({i_4_, n42, n334, n804}, n16);
	defparam lut_18.LUT_SIZE = 4;
	defparam lut_18.mask = 16'H0057;

	lut_sub lut_19 ({n574, n577, n585, n596, n597, n599, n600, n601}, n18);
	defparam lut_19.LUT_SIZE = 8;
	defparam lut_19.mask = 256'H0000000000000000000000000000000000000000000000000000000080000000;

	lut_sub lut_20 ({i_0_, n23, n641, n640}, n19);
	defparam lut_20.LUT_SIZE = 4;
	defparam lut_20.mask = 16'H080C;

	lut_sub lut_21 ({i_1_, i_3_}, n21);
	defparam lut_21.LUT_SIZE = 2;
	defparam lut_21.mask = 4'b0111;

	lut_sub lut_22 ({i_5_, n21}, n20);
	defparam lut_22.LUT_SIZE = 2;
	defparam lut_22.mask = 4'b1011;

	lut_sub lut_23 ({i_8_, i_10_}, n24);
	defparam lut_23.LUT_SIZE = 2;
	defparam lut_23.mask = 4'b0010;

	lut_sub lut_24 ({i_3_, n24, n542}, n23);
	defparam lut_24.LUT_SIZE = 3;
	defparam lut_24.mask = 8'HD0;

	lut_sub lut_25 ({i_6_, i_10_, n53}, n26);
	defparam lut_25.LUT_SIZE = 3;
	defparam lut_25.mask = 8'H15;

	lut_sub lut_26 ({n39, n125, n655, n35}, n33);
	defparam lut_26.LUT_SIZE = 4;
	defparam lut_26.mask = 16'HEEE0;

	lut_sub lut_27 ({i_1_, n557}, n31);
	defparam lut_27.LUT_SIZE = 2;
	defparam lut_27.mask = 4'b1110;

	lut_sub lut_28 ({i_11_, n118}, n32);
	defparam lut_28.LUT_SIZE = 2;
	defparam lut_28.mask = 4'b1110;

	lut_sub lut_29 ({n33, n31, n32}, n30);
	defparam lut_29.LUT_SIZE = 3;
	defparam lut_29.mask = 8'HE0;

	lut_sub lut_30 ({i_12_, n118}, n35);
	defparam lut_30.LUT_SIZE = 2;
	defparam lut_30.mask = 4'b1110;

	lut_sub lut_31 ({i_0_, n247}, n36);
	defparam lut_31.LUT_SIZE = 2;
	defparam lut_31.mask = 4'b1110;

	lut_sub lut_32 ({n31, n35, i_11_, n36}, n34);
	defparam lut_32.LUT_SIZE = 4;
	defparam lut_32.mask = 16'HEEE0;

	lut_sub lut_33 ({i_6_, i_7_}, n38);
	defparam lut_33.LUT_SIZE = 2;
	defparam lut_33.mask = 4'b1011;

	lut_sub lut_34 ({i_0_, n233}, n39);
	defparam lut_34.LUT_SIZE = 2;
	defparam lut_34.mask = 4'b1110;

	lut_sub lut_35 ({i_0_, i_1_, i_2_}, n40);
	defparam lut_35.LUT_SIZE = 3;
	defparam lut_35.mask = 8'HFD;

	lut_sub lut_36 ({n38, n39, i_6_, n40}, n37);
	defparam lut_36.LUT_SIZE = 4;
	defparam lut_36.mask = 16'HEEE0;

	lut_sub lut_37 ({i_3_, n247}, n42);
	defparam lut_37.LUT_SIZE = 2;
	defparam lut_37.mask = 4'b1011;

	lut_sub lut_38 ({i_3_, n557}, n43);
	defparam lut_38.LUT_SIZE = 2;
	defparam lut_38.mask = 4'b1011;

	lut_sub lut_39 ({i_5_, i_6_, n42, n43}, n41);
	defparam lut_39.LUT_SIZE = 4;
	defparam lut_39.mask = 16'H8CAF;

	lut_sub lut_40 ({i_0_, n45}, n46);
	defparam lut_40.LUT_SIZE = 2;
	defparam lut_40.mask = 4'b1110;

	lut_sub lut_41 ({i_3_, i_2_}, n45);
	defparam lut_41.LUT_SIZE = 2;
	defparam lut_41.mask = 4'b1110;

	lut_sub lut_42 ({i_5_, n46, n45}, n44);
	defparam lut_42.LUT_SIZE = 3;
	defparam lut_42.mask = 8'H8C;

	lut_sub lut_43 ({i_12_, i_13_}, n50);
	defparam lut_43.LUT_SIZE = 2;
	defparam lut_43.mask = 4'b0010;

	lut_sub lut_44 ({i_8_, n50, n471, n763}, n47);
	defparam lut_44.LUT_SIZE = 4;
	defparam lut_44.mask = 16'H7050;

	lut_sub lut_45 ({i_6_, n653}, n53);
	defparam lut_45.LUT_SIZE = 2;
	defparam lut_45.mask = 4'b1000;

	lut_sub lut_46 ({n53, n174, n497, n765}, n51);
	defparam lut_46.LUT_SIZE = 4;
	defparam lut_46.mask = 16'H0705;

	lut_sub lut_47 ({i_6_, n46, i_7_, n223}, n57);
	defparam lut_47.LUT_SIZE = 4;
	defparam lut_47.mask = 16'HEEE0;

	lut_sub lut_48 ({n57, i_8_, n39}, n56);
	defparam lut_48.LUT_SIZE = 3;
	defparam lut_48.mask = 8'HE0;

	lut_sub lut_49 ({i_12_, n118}, n61);
	defparam lut_49.LUT_SIZE = 2;
	defparam lut_49.mask = 4'b1011;

	lut_sub lut_50 ({i_1_, i_6_, n61, n421}, n58);
	defparam lut_50.LUT_SIZE = 4;
	defparam lut_50.mask = 16'H4C5F;

	lut_sub lut_51 ({i_1_, i_6_}, n63);
	defparam lut_51.LUT_SIZE = 2;
	defparam lut_51.mask = 4'b0010;

	lut_sub lut_52 ({i_0_, i_1_, i_5_, n63}, n62);
	defparam lut_52.LUT_SIZE = 4;
	defparam lut_52.mask = 16'H8ACF;

	lut_sub lut_53 ({i_9_, n73, n364}, n65);
	defparam lut_53.LUT_SIZE = 3;
	defparam lut_53.mask = 8'H01;

	lut_sub lut_54 ({i_3_, n61, n65, n99}, n69);
	defparam lut_54.LUT_SIZE = 4;
	defparam lut_54.mask = 16'HCD00;

	lut_sub lut_55 ({i_11_, n118}, n73);
	defparam lut_55.LUT_SIZE = 2;
	defparam lut_55.mask = 4'b1011;

	lut_sub lut_56 ({i_8_, i_6_}, n74);
	defparam lut_56.LUT_SIZE = 2;
	defparam lut_56.mask = 4'b1110;

	lut_sub lut_57 ({i_2_, i_9_, n73, n74}, n72);
	defparam lut_57.LUT_SIZE = 4;
	defparam lut_57.mask = 16'HFEFF;

	lut_sub lut_58 ({i_0_, n45}, n77);
	defparam lut_58.LUT_SIZE = 2;
	defparam lut_58.mask = 4'b1011;

	lut_sub lut_59 ({i_0_, n216}, n78);
	defparam lut_59.LUT_SIZE = 2;
	defparam lut_59.mask = 4'b1011;

	lut_sub lut_60 ({i_6_, n77, i_7_, n78}, n76);
	defparam lut_60.LUT_SIZE = 4;
	defparam lut_60.mask = 16'HEEE0;

	lut_sub lut_61 ({i_0_, n69, n72, n778}, n79);
	defparam lut_61.LUT_SIZE = 4;
	defparam lut_61.mask = 16'HF700;

	lut_sub lut_62 ({i_3_, i_11_, n39, n421}, n83);
	defparam lut_62.LUT_SIZE = 4;
	defparam lut_62.mask = 16'HFFDF;

	lut_sub lut_63 ({i_3_, i_9_, n118, n497}, n84);
	defparam lut_63.LUT_SIZE = 4;
	defparam lut_63.mask = 16'HFEFF;

	lut_sub lut_64 ({i_5_, n58, n197}, n85);
	defparam lut_64.LUT_SIZE = 3;
	defparam lut_64.mask = 8'HEF;

	lut_sub lut_65 ({n196, n406, n650}, n87);
	defparam lut_65.LUT_SIZE = 3;
	defparam lut_65.mask = 8'HFB;

	lut_sub lut_66 ({n656, n73, i_9_, n62}, n88);
	defparam lut_66.LUT_SIZE = 4;
	defparam lut_66.mask = 16'HFFFE;

	lut_sub lut_67 ({n79, n83, n84, n85, n87, n88}, n82);
	defparam lut_67.LUT_SIZE = 6;
	defparam lut_67.mask = 64'H0000000080000000;

	lut_sub lut_68 ({n144, n655, n98, n173}, n91);
	defparam lut_68.LUT_SIZE = 4;
	defparam lut_68.mask = 16'HEEE0;

	lut_sub lut_69 ({i_6_, n656}, n90);
	defparam lut_69.LUT_SIZE = 2;
	defparam lut_69.mask = 4'b1011;

	lut_sub lut_70 ({n91, n90, n31}, n89);
	defparam lut_70.LUT_SIZE = 3;
	defparam lut_70.mask = 8'HE0;

	lut_sub lut_71 ({n53, n101, n173, n655}, n93);
	defparam lut_71.LUT_SIZE = 4;
	defparam lut_71.mask = 16'H8CAF;

	lut_sub lut_72 ({n654, n497, n652, n31}, n94);
	defparam lut_72.LUT_SIZE = 4;
	defparam lut_72.mask = 16'HEEE0;

	lut_sub lut_73 ({n93, n94}, n92);
	defparam lut_73.LUT_SIZE = 2;
	defparam lut_73.mask = 4'b1000;

	lut_sub lut_74 ({n36, n102, n108, n144}, n96);
	defparam lut_74.LUT_SIZE = 4;
	defparam lut_74.mask = 16'HAF8C;

	lut_sub lut_75 ({n96, n40, n90}, n95);
	defparam lut_75.LUT_SIZE = 3;
	defparam lut_75.mask = 8'HE0;

	lut_sub lut_76 ({i_6_, n326}, n99);
	defparam lut_76.LUT_SIZE = 2;
	defparam lut_76.mask = 4'b1011;

	lut_sub lut_77 ({i_6_, i_7_, i_8_}, n98);
	defparam lut_77.LUT_SIZE = 3;
	defparam lut_77.mask = 8'HBF;

	lut_sub lut_78 ({n99, n95, n98, n39}, n97);
	defparam lut_78.LUT_SIZE = 4;
	defparam lut_78.mask = 16'HE000;

	lut_sub lut_79 ({i_5_, n453}, n104);
	defparam lut_79.LUT_SIZE = 2;
	defparam lut_79.mask = 4'b1000;

	lut_sub lut_80 ({i_6_, n653}, n101);
	defparam lut_80.LUT_SIZE = 2;
	defparam lut_80.mask = 4'b0010;

	lut_sub lut_81 ({i_0_, i_1_, i_2_}, n102);
	defparam lut_81.LUT_SIZE = 3;
	defparam lut_81.mask = 8'H04;

	lut_sub lut_82 ({n104, n101, n102, n757}, n100);
	defparam lut_82.LUT_SIZE = 4;
	defparam lut_82.mask = 16'HD500;

	lut_sub lut_83 ({i_11_, n185}, n106);
	defparam lut_83.LUT_SIZE = 2;
	defparam lut_83.mask = 4'b1101;

	lut_sub lut_84 ({i_10_, n364}, n107);
	defparam lut_84.LUT_SIZE = 2;
	defparam lut_84.mask = 4'b1110;

	lut_sub lut_85 ({i_6_, n656}, n108);
	defparam lut_85.LUT_SIZE = 2;
	defparam lut_85.mask = 4'b1110;

	lut_sub lut_86 ({n106, n107, n108, n32}, n105);
	defparam lut_86.LUT_SIZE = 4;
	defparam lut_86.mask = 16'HEEE0;

	lut_sub lut_87 ({i_12_, n114}, n110);
	defparam lut_87.LUT_SIZE = 2;
	defparam lut_87.mask = 4'b1110;

	lut_sub lut_88 ({i_11_, n114}, n111);
	defparam lut_88.LUT_SIZE = 2;
	defparam lut_88.mask = 4'b1110;

	lut_sub lut_89 ({n53, n98, n110, n111}, n109);
	defparam lut_89.LUT_SIZE = 4;
	defparam lut_89.mask = 16'HC8FA;

	lut_sub lut_90 ({i_11_, i_12_}, n113);
	defparam lut_90.LUT_SIZE = 2;
	defparam lut_90.mask = 4'b1110;

	lut_sub lut_91 ({i_9_, i_13_}, n114);
	defparam lut_91.LUT_SIZE = 2;
	defparam lut_91.mask = 4'b1110;

	lut_sub lut_92 ({n113, n114, i_3_, i_10_}, n112);
	defparam lut_92.LUT_SIZE = 4;
	defparam lut_92.mask = 16'HFFFE;

	lut_sub lut_93 ({i_5_, n376}, n116);
	defparam lut_93.LUT_SIZE = 2;
	defparam lut_93.mask = 4'b1110;

	lut_sub lut_94 ({i_10_, i_13_}, n118);
	defparam lut_94.LUT_SIZE = 2;
	defparam lut_94.mask = 4'b1110;

	lut_sub lut_95 ({i_10_, n116, n118, n181}, n115);
	defparam lut_95.LUT_SIZE = 4;
	defparam lut_95.mask = 16'HD0DD;

	lut_sub lut_96 ({i_13_, n684, n685, n749}, n119);
	defparam lut_96.LUT_SIZE = 4;
	defparam lut_96.mask = 16'H5700;

	lut_sub lut_97 ({i_5_, n649}, n124);
	defparam lut_97.LUT_SIZE = 2;
	defparam lut_97.mask = 4'b1110;

	lut_sub lut_98 ({i_12_, n406}, n125);
	defparam lut_98.LUT_SIZE = 2;
	defparam lut_98.mask = 4'b1101;

	lut_sub lut_99 ({n124, n125, n181, n268}, n123);
	defparam lut_99.LUT_SIZE = 4;
	defparam lut_99.mask = 16'H7770;

	lut_sub lut_100 ({i_3_, i_11_, n50, n748}, n127);
	defparam lut_100.LUT_SIZE = 4;
	defparam lut_100.mask = 16'H444C;

	lut_sub lut_101 ({n652, n692, n693}, n132);
	defparam lut_101.LUT_SIZE = 3;
	defparam lut_101.mask = 8'HFE;

	lut_sub lut_102 ({n144, n690, n691}, n133);
	defparam lut_102.LUT_SIZE = 3;
	defparam lut_102.mask = 8'HFE;

	lut_sub lut_103 ({n220, n287, n656}, n134);
	defparam lut_103.LUT_SIZE = 3;
	defparam lut_103.mask = 8'HFB;

	lut_sub lut_104 ({n53, n104, n421}, n135);
	defparam lut_104.LUT_SIZE = 3;
	defparam lut_104.mask = 8'H7F;

	lut_sub lut_105 ({n108, n406, n565}, n136);
	defparam lut_105.LUT_SIZE = 3;
	defparam lut_105.mask = 8'HFB;

	lut_sub lut_106 ({n98, n383, n658}, n138);
	defparam lut_106.LUT_SIZE = 3;
	defparam lut_106.mask = 8'HFB;

	lut_sub lut_107 ({n123, n654, n681, n683}, n139);
	defparam lut_107.LUT_SIZE = 4;
	defparam lut_107.mask = 16'HEEE0;

	lut_sub lut_108 ({n127, n132, n133, n134, n135, n136, n138, n139}, n131);
	defparam lut_108.LUT_SIZE = 8;
	defparam lut_108.mask = 256'H0000000000000000000000000000000080000000000000000000000000000000;

	lut_sub lut_109 ({n90, n108, n499, n522}, n140);
	defparam lut_109.LUT_SIZE = 4;
	defparam lut_109.mask = 16'HF531;

	lut_sub lut_110 ({n164, n688, n188, n165}, n146);
	defparam lut_110.LUT_SIZE = 4;
	defparam lut_110.mask = 16'HEEE0;

	lut_sub lut_111 ({n746, n747, n682, n687}, n147);
	defparam lut_111.LUT_SIZE = 4;
	defparam lut_111.mask = 16'HE000;

	lut_sub lut_112 ({i_7_, n74}, n144);
	defparam lut_112.LUT_SIZE = 2;
	defparam lut_112.mask = 4'b1011;

	lut_sub lut_113 ({n104, n268}, n145);
	defparam lut_113.LUT_SIZE = 2;
	defparam lut_113.mask = 4'b0111;

	lut_sub lut_114 ({n146, n147, n144, n145}, n143);
	defparam lut_114.LUT_SIZE = 4;
	defparam lut_114.mask = 16'HE000;

	lut_sub lut_115 ({i_0_, i_1_, i_4_}, n149);
	defparam lut_115.LUT_SIZE = 3;
	defparam lut_115.mask = 8'HBF;

	lut_sub lut_116 ({i_4_, n557}, n151);
	defparam lut_116.LUT_SIZE = 2;
	defparam lut_116.mask = 4'b1110;

	lut_sub lut_117 ({i_6_, i_7_, n149, n151}, n148);
	defparam lut_117.LUT_SIZE = 4;
	defparam lut_117.mask = 16'H8ACF;

	lut_sub lut_118 ({i_2_, i_8_, n241, n658}, n152);
	defparam lut_118.LUT_SIZE = 4;
	defparam lut_118.mask = 16'H0100;

	lut_sub lut_119 ({n683, n686}, n157);
	defparam lut_119.LUT_SIZE = 2;
	defparam lut_119.mask = 4'b1110;

	lut_sub lut_120 ({n108, n174, n179}, n158);
	defparam lut_120.LUT_SIZE = 3;
	defparam lut_120.mask = 8'HFE;

	lut_sub lut_121 ({n101, n692, n693}, n159);
	defparam lut_121.LUT_SIZE = 3;
	defparam lut_121.mask = 8'HEF;

	lut_sub lut_122 ({n90, n690, n691}, n160);
	defparam lut_122.LUT_SIZE = 3;
	defparam lut_122.mask = 8'HFE;

	lut_sub lut_123 ({n220, n688, n217, n165}, n161);
	defparam lut_123.LUT_SIZE = 4;
	defparam lut_123.mask = 16'HEEE0;

	lut_sub lut_124 ({n684, n687, n144, n680}, n162);
	defparam lut_124.LUT_SIZE = 4;
	defparam lut_124.mask = 16'HEEE0;

	lut_sub lut_125 ({n157, n158, n159, n160, n161, n162}, n156);
	defparam lut_125.LUT_SIZE = 6;
	defparam lut_125.mask = 64'H8000000000000000;

	lut_sub lut_126 ({n98, n680, n188, n688}, n166);
	defparam lut_126.LUT_SIZE = 4;
	defparam lut_126.mask = 16'HEEE0;

	lut_sub lut_127 ({n744, n745, n682, n686}, n167);
	defparam lut_127.LUT_SIZE = 4;
	defparam lut_127.mask = 16'HE000;

	lut_sub lut_128 ({i_5_, n222}, n164);
	defparam lut_128.LUT_SIZE = 2;
	defparam lut_128.mask = 4'b1011;

	lut_sub lut_129 ({n50, n315}, n165);
	defparam lut_129.LUT_SIZE = 2;
	defparam lut_129.mask = 4'b0111;

	lut_sub lut_130 ({n166, n167, n164, n165}, n163);
	defparam lut_130.LUT_SIZE = 4;
	defparam lut_130.mask = 16'HE000;

	lut_sub lut_131 ({n90, n98, n499, n522}, n168);
	defparam lut_131.LUT_SIZE = 4;
	defparam lut_131.mask = 16'HF351;

	lut_sub lut_132 ({n189, n220, n681, n684}, n170);
	defparam lut_132.LUT_SIZE = 4;
	defparam lut_132.mask = 16'HEEE0;

	lut_sub lut_133 ({n742, n743, n677, n683}, n171);
	defparam lut_133.LUT_SIZE = 4;
	defparam lut_133.mask = 16'HE000;

	lut_sub lut_134 ({n170, n171, n90, n145}, n169);
	defparam lut_134.LUT_SIZE = 4;
	defparam lut_134.mask = 16'HE000;

	lut_sub lut_135 ({i_0_, n233}, n173);
	defparam lut_135.LUT_SIZE = 2;
	defparam lut_135.mask = 4'b1011;

	lut_sub lut_136 ({i_5_, n376}, n174);
	defparam lut_136.LUT_SIZE = 2;
	defparam lut_136.mask = 4'b1011;

	lut_sub lut_137 ({n173, n144, n174}, n172);
	defparam lut_137.LUT_SIZE = 3;
	defparam lut_137.mask = 8'HFE;

	lut_sub lut_138 ({n98, n102, n116}, n175);
	defparam lut_138.LUT_SIZE = 3;
	defparam lut_138.mask = 8'HFB;

	lut_sub lut_139 ({i_2_, n376}, n178);
	defparam lut_139.LUT_SIZE = 2;
	defparam lut_139.mask = 4'b1110;

	lut_sub lut_140 ({i_10_, n383}, n179);
	defparam lut_140.LUT_SIZE = 2;
	defparam lut_140.mask = 4'b0111;

	lut_sub lut_141 ({i_5_, n90, n178, n179}, n177);
	defparam lut_141.LUT_SIZE = 4;
	defparam lut_141.mask = 16'HFEFF;

	lut_sub lut_142 ({i_3_, i_4_, i_5_}, n181);
	defparam lut_142.LUT_SIZE = 3;
	defparam lut_142.mask = 8'H40;

	lut_sub lut_143 ({i_1_, i_7_, n73, n181}, n180);
	defparam lut_143.LUT_SIZE = 4;
	defparam lut_143.mask = 16'H0200;

	lut_sub lut_144 ({i_12_, i_13_}, n185);
	defparam lut_144.LUT_SIZE = 2;
	defparam lut_144.mask = 4'b0001;

	lut_sub lut_145 ({i_10_, i_11_}, n186);
	defparam lut_145.LUT_SIZE = 2;
	defparam lut_145.mask = 4'b1000;

	lut_sub lut_146 ({n172, n175, n185, n186}, n182);
	defparam lut_146.LUT_SIZE = 4;
	defparam lut_146.mask = 16'H0888;

	lut_sub lut_147 ({n675, n164, n677, n682}, n190);
	defparam lut_147.LUT_SIZE = 4;
	defparam lut_147.mask = 16'HEEE0;

	lut_sub lut_148 ({n108, n145, n559, n681}, n191);
	defparam lut_148.LUT_SIZE = 4;
	defparam lut_148.mask = 16'HBBB0;

	lut_sub lut_149 ({i_3_, n673}, n188);
	defparam lut_149.LUT_SIZE = 2;
	defparam lut_149.mask = 4'b1110;

	lut_sub lut_150 ({n50, n548}, n189);
	defparam lut_150.LUT_SIZE = 2;
	defparam lut_150.mask = 4'b0111;

	lut_sub lut_151 ({n190, n191, n188, n189}, n187);
	defparam lut_151.LUT_SIZE = 4;
	defparam lut_151.mask = 16'HE000;

	lut_sub lut_152 ({n188, n559, n675, n677}, n193);
	defparam lut_152.LUT_SIZE = 4;
	defparam lut_152.mask = 16'HAF8C;

	lut_sub lut_153 ({n90, n680, n681, n682}, n194);
	defparam lut_153.LUT_SIZE = 4;
	defparam lut_153.mask = 16'HEEE0;

	lut_sub lut_154 ({n193, n194, n189, n164}, n192);
	defparam lut_154.LUT_SIZE = 4;
	defparam lut_154.mask = 16'HE000;

	lut_sub lut_155 ({i_10_, n656}, n196);
	defparam lut_155.LUT_SIZE = 2;
	defparam lut_155.mask = 4'b1110;

	lut_sub lut_156 ({i_8_, n326}, n197);
	defparam lut_156.LUT_SIZE = 2;
	defparam lut_156.mask = 4'b1011;

	lut_sub lut_157 ({n196, n197}, n195);
	defparam lut_157.LUT_SIZE = 2;
	defparam lut_157.mask = 4'b1000;

	lut_sub lut_158 ({n195, n578, n582, n738}, n201);
	defparam lut_158.LUT_SIZE = 4;
	defparam lut_158.mask = 16'HAF23;

	lut_sub lut_159 ({n740, n667, n39}, n202);
	defparam lut_159.LUT_SIZE = 3;
	defparam lut_159.mask = 8'HE0;

	lut_sub lut_160 ({n107, n99}, n199);
	defparam lut_160.LUT_SIZE = 2;
	defparam lut_160.mask = 4'b1000;

	lut_sub lut_161 ({n201, n202, n199, n481}, n198);
	defparam lut_161.LUT_SIZE = 4;
	defparam lut_161.mask = 16'HD000;

	lut_sub lut_162 ({n107, n409, n565, n669}, n206);
	defparam lut_162.LUT_SIZE = 4;
	defparam lut_162.mask = 16'HAF8C;

	lut_sub lut_163 ({i_8_, n668}, n204);
	defparam lut_163.LUT_SIZE = 2;
	defparam lut_163.mask = 4'b1110;

	lut_sub lut_164 ({i_4_, n233}, n205);
	defparam lut_164.LUT_SIZE = 2;
	defparam lut_164.mask = 4'b1011;

	lut_sub lut_165 ({n206, n204, n205}, n203);
	defparam lut_165.LUT_SIZE = 3;
	defparam lut_165.mask = 8'HE0;

	lut_sub lut_166 ({n402, n670, n671, n672}, n210);
	defparam lut_166.LUT_SIZE = 4;
	defparam lut_166.mask = 16'HCF8A;

	lut_sub lut_167 ({n99, n104, n205, n602}, n211);
	defparam lut_167.LUT_SIZE = 4;
	defparam lut_167.mask = 16'HEE0E;

	lut_sub lut_168 ({i_5_, n326}, n209);
	defparam lut_168.LUT_SIZE = 2;
	defparam lut_168.mask = 4'b1011;

	lut_sub lut_169 ({n210, n211, n209, n409}, n207);
	defparam lut_169.LUT_SIZE = 4;
	defparam lut_169.mask = 16'HD000;

	lut_sub lut_170 ({n654, n173, n652, n655}, n214);
	defparam lut_170.LUT_SIZE = 4;
	defparam lut_170.mask = 16'HEEE0;

	lut_sub lut_171 ({n31, n101, n214}, n212);
	defparam lut_171.LUT_SIZE = 3;
	defparam lut_171.mask = 8'HA2;

	lut_sub lut_172 ({i_3_, n236}, n217);
	defparam lut_172.LUT_SIZE = 2;
	defparam lut_172.mask = 4'b1110;

	lut_sub lut_173 ({i_1_, i_3_}, n216);
	defparam lut_173.LUT_SIZE = 2;
	defparam lut_173.mask = 4'b1110;

	lut_sub lut_174 ({i_5_, n217, n216}, n215);
	defparam lut_174.LUT_SIZE = 3;
	defparam lut_174.mask = 8'H8C;

	lut_sub lut_175 ({i_0_, i_3_, i_6_}, n218);
	defparam lut_175.LUT_SIZE = 3;
	defparam lut_175.mask = 8'HFD;

	lut_sub lut_176 ({i_3_, n650}, n220);
	defparam lut_176.LUT_SIZE = 2;
	defparam lut_176.mask = 4'b1110;

	lut_sub lut_177 ({n220, i_5_, n216}, n219);
	defparam lut_177.LUT_SIZE = 3;
	defparam lut_177.mask = 8'HE0;

	lut_sub lut_178 ({i_0_, n216}, n223);
	defparam lut_178.LUT_SIZE = 2;
	defparam lut_178.mask = 4'b1110;

	lut_sub lut_179 ({i_3_, i_6_}, n222);
	defparam lut_179.LUT_SIZE = 2;
	defparam lut_179.mask = 4'b1110;

	lut_sub lut_180 ({n223, n219, i_0_, n222}, n221);
	defparam lut_180.LUT_SIZE = 4;
	defparam lut_180.mask = 16'HE000;

	lut_sub lut_181 ({i_0_, i_3_, i_6_}, n224);
	defparam lut_181.LUT_SIZE = 3;
	defparam lut_181.mask = 8'H7F;

	lut_sub lut_182 ({i_1_, i_6_}, n226);
	defparam lut_182.LUT_SIZE = 2;
	defparam lut_182.mask = 4'b0100;

	lut_sub lut_183 ({i_2_, i_6_, i_7_, n226}, n225);
	defparam lut_183.LUT_SIZE = 4;
	defparam lut_183.mask = 16'HBB0B;

	lut_sub lut_184 ({i_6_, n945, n651}, n229);
	defparam lut_184.LUT_SIZE = 3;
	defparam lut_184.mask = 8'HFE;

	lut_sub lut_185 ({i_1_, i_7_, n651}, n230);
	defparam lut_185.LUT_SIZE = 3;
	defparam lut_185.mask = 8'HFE;

	lut_sub lut_186 ({i_11_, n542}, n228);
	defparam lut_186.LUT_SIZE = 2;
	defparam lut_186.mask = 4'b1110;

	lut_sub lut_187 ({n229, n230, n225, n228}, n227);
	defparam lut_187.LUT_SIZE = 4;
	defparam lut_187.mask = 16'HE000;

	lut_sub lut_188 ({i_5_, n45}, n231);
	defparam lut_188.LUT_SIZE = 2;
	defparam lut_188.mask = 4'b1110;

	lut_sub lut_189 ({i_2_, n650}, n234);
	defparam lut_189.LUT_SIZE = 2;
	defparam lut_189.mask = 4'b1110;

	lut_sub lut_190 ({i_1_, i_2_}, n233);
	defparam lut_190.LUT_SIZE = 2;
	defparam lut_190.mask = 4'b1110;

	lut_sub lut_191 ({n234, i_5_, n233}, n232);
	defparam lut_191.LUT_SIZE = 3;
	defparam lut_191.mask = 8'HE0;

	lut_sub lut_192 ({i_5_, i_6_}, n236);
	defparam lut_192.LUT_SIZE = 2;
	defparam lut_192.mask = 4'b0111;

	lut_sub lut_193 ({i_2_, i_5_, n233, n236}, n235);
	defparam lut_193.LUT_SIZE = 4;
	defparam lut_193.mask = 16'HCF8A;

	lut_sub lut_194 ({i_2_, i_5_, n236, n247}, n238);
	defparam lut_194.LUT_SIZE = 4;
	defparam lut_194.mask = 16'H8CAF;

	lut_sub lut_195 ({i_6_, n557}, n239);
	defparam lut_195.LUT_SIZE = 2;
	defparam lut_195.mask = 4'b1011;

	lut_sub lut_196 ({n238, n239}, n237);
	defparam lut_196.LUT_SIZE = 2;
	defparam lut_196.mask = 4'b1000;

	lut_sub lut_197 ({i_1_, i_5_, i_7_}, n242);
	defparam lut_197.LUT_SIZE = 3;
	defparam lut_197.mask = 8'H7F;

	lut_sub lut_198 ({i_1_, i_6_}, n241);
	defparam lut_198.LUT_SIZE = 2;
	defparam lut_198.mask = 4'b0001;

	lut_sub lut_199 ({i_0_, i_7_, n242, n241}, n240);
	defparam lut_199.LUT_SIZE = 4;
	defparam lut_199.mask = 16'H8CCC;

	lut_sub lut_200 ({i_10_, n237, n240, n542}, n243);
	defparam lut_200.LUT_SIZE = 4;
	defparam lut_200.mask = 16'H1500;

	lut_sub lut_201 ({i_2_, n650}, n248);
	defparam lut_201.LUT_SIZE = 2;
	defparam lut_201.mask = 4'b1011;

	lut_sub lut_202 ({i_6_, n557}, n249);
	defparam lut_202.LUT_SIZE = 2;
	defparam lut_202.mask = 4'b1110;

	lut_sub lut_203 ({i_1_, i_2_}, n247);
	defparam lut_203.LUT_SIZE = 2;
	defparam lut_203.mask = 4'b0111;

	lut_sub lut_204 ({n248, n249, i_5_, n247}, n246);
	defparam lut_204.LUT_SIZE = 4;
	defparam lut_204.mask = 16'HE000;

	lut_sub lut_205 ({n246, i_7_, n62}, n250);
	defparam lut_205.LUT_SIZE = 3;
	defparam lut_205.mask = 8'HE0;

	lut_sub lut_206 ({i_0_, i_1_, i_5_, i_6_}, n251);
	defparam lut_206.LUT_SIZE = 4;
	defparam lut_206.mask = 16'H8ACF;

	lut_sub lut_207 ({i_7_, n149, i_6_, n151}, n252);
	defparam lut_207.LUT_SIZE = 4;
	defparam lut_207.mask = 16'HEEE0;

	lut_sub lut_208 ({i_2_, i_8_, n63, n124}, n255);
	defparam lut_208.LUT_SIZE = 4;
	defparam lut_208.mask = 16'HEFFF;

	lut_sub lut_209 ({n252, n255, n604}, n253);
	defparam lut_209.LUT_SIZE = 3;
	defparam lut_209.mask = 8'HC4;

	lut_sub lut_210 ({n36, n53, n102, n652}, n257);
	defparam lut_210.LUT_SIZE = 4;
	defparam lut_210.mask = 16'HBB0B;

	lut_sub lut_211 ({n40, n101, n257}, n256);
	defparam lut_211.LUT_SIZE = 3;
	defparam lut_211.mask = 8'HA2;

	lut_sub lut_212 ({i_4_, n247}, n259);
	defparam lut_212.LUT_SIZE = 2;
	defparam lut_212.mask = 4'b1011;

	lut_sub lut_213 ({i_4_, n696}, n260);
	defparam lut_213.LUT_SIZE = 2;
	defparam lut_213.mask = 4'b1011;

	lut_sub lut_214 ({i_8_, n259, i_6_, n260}, n258);
	defparam lut_214.LUT_SIZE = 4;
	defparam lut_214.mask = 16'HEEE0;

	lut_sub lut_215 ({i_1_, i_4_, n196, n775}, n261);
	defparam lut_215.LUT_SIZE = 4;
	defparam lut_215.mask = 16'H5070;

	lut_sub lut_216 ({i_6_, i_10_, n261, n670}, n264);
	defparam lut_216.LUT_SIZE = 4;
	defparam lut_216.mask = 16'H3331;

	lut_sub lut_217 ({i_9_, n406}, n268);
	defparam lut_217.LUT_SIZE = 2;
	defparam lut_217.mask = 4'b0010;

	lut_sub lut_218 ({n181, n256, n268}, n267);
	defparam lut_218.LUT_SIZE = 3;
	defparam lut_218.mask = 8'H20;

	lut_sub lut_219 ({i_10_, i_13_, n506}, n271);
	defparam lut_219.LUT_SIZE = 3;
	defparam lut_219.mask = 8'H02;

	lut_sub lut_220 ({n89, n124, n271, n720}, n270);
	defparam lut_220.LUT_SIZE = 4;
	defparam lut_220.mask = 16'H050D;

	lut_sub lut_221 ({i_3_, i_8_}, n276);
	defparam lut_221.LUT_SIZE = 2;
	defparam lut_221.mask = 4'b0001;

	lut_sub lut_222 ({n148, n152, n276, n659}, n275);
	defparam lut_222.LUT_SIZE = 4;
	defparam lut_222.mask = 16'H5054;

	lut_sub lut_223 ({i_9_, i_13_, n479}, n280);
	defparam lut_223.LUT_SIZE = 3;
	defparam lut_223.mask = 8'H02;

	lut_sub lut_224 ({n212, n280, n658, n723}, n279);
	defparam lut_224.LUT_SIZE = 4;
	defparam lut_224.mask = 16'H1131;

	lut_sub lut_225 ({i_11_, i_13_}, n287);
	defparam lut_225.LUT_SIZE = 2;
	defparam lut_225.mask = 4'b0010;

	lut_sub lut_226 ({n248, n287, n662, n726}, n283);
	defparam lut_226.LUT_SIZE = 4;
	defparam lut_226.mask = 16'H5070;

	lut_sub lut_227 ({n50, n730, n732, n734}, n288);
	defparam lut_227.LUT_SIZE = 4;
	defparam lut_227.mask = 16'H7F00;

	lut_sub lut_228 ({n406, i_12_}, n296);
	defparam lut_228.LUT_SIZE = 2;
	defparam lut_228.mask = 4'b1000;

	lut_sub lut_229 ({n198, n203, n207, n296}, n292);
	defparam lut_229.LUT_SIZE = 4;
	defparam lut_229.mask = 16'H2AAA;

	lut_sub lut_230 ({n61, n759, n761, n762}, n297);
	defparam lut_230.LUT_SIZE = 4;
	defparam lut_230.mask = 16'H007F;

	lut_sub lut_231 ({i_4_, i_8_, n287, n506}, n302);
	defparam lut_231.LUT_SIZE = 4;
	defparam lut_231.mask = 16'H3313;

	lut_sub lut_232 ({i_3_, n228, n406, n667}, n303);
	defparam lut_232.LUT_SIZE = 4;
	defparam lut_232.mask = 16'HB0BB;

	lut_sub lut_233 ({n125, n302, n303, n604}, n301);
	defparam lut_233.LUT_SIZE = 4;
	defparam lut_233.mask = 16'HC040;

	lut_sub lut_234 ({i_7_, i_10_}, n306);
	defparam lut_234.LUT_SIZE = 2;
	defparam lut_234.mask = 4'b1011;

	lut_sub lut_235 ({i_4_, n479}, n307);
	defparam lut_235.LUT_SIZE = 2;
	defparam lut_235.mask = 4'b1101;

	lut_sub lut_236 ({i_7_, n306, n307, n384}, n304);
	defparam lut_236.LUT_SIZE = 4;
	defparam lut_236.mask = 16'HC4F5;

	lut_sub lut_237 ({i_7_, n24}, n308);
	defparam lut_237.LUT_SIZE = 2;
	defparam lut_237.mask = 4'b1000;

	lut_sub lut_238 ({i_8_, n304, n308, n698}, n311);
	defparam lut_238.LUT_SIZE = 4;
	defparam lut_238.mask = 16'HBBB0;

	lut_sub lut_239 ({i_7_, n301, n311, n915}, n309);
	defparam lut_239.LUT_SIZE = 4;
	defparam lut_239.mask = 16'H4440;

	lut_sub lut_240 ({i_7_, i_9_}, n313);
	defparam lut_240.LUT_SIZE = 2;
	defparam lut_240.mask = 4'b0111;

	lut_sub lut_241 ({i_7_, i_10_, n313}, n312);
	defparam lut_241.LUT_SIZE = 3;
	defparam lut_241.mask = 8'HA2;

	lut_sub lut_242 ({i_7_, i_8_, i_10_}, n315);
	defparam lut_242.LUT_SIZE = 3;
	defparam lut_242.mask = 8'H08;

	lut_sub lut_243 ({i_12_, n315, n685}, n314);
	defparam lut_243.LUT_SIZE = 3;
	defparam lut_243.mask = 8'HD0;

	lut_sub lut_244 ({i_10_, n656}, n317);
	defparam lut_244.LUT_SIZE = 2;
	defparam lut_244.mask = 4'b1011;

	lut_sub lut_245 ({i_8_, n313}, n318);
	defparam lut_245.LUT_SIZE = 2;
	defparam lut_245.mask = 4'b1110;

	lut_sub lut_246 ({i_11_, n314, n317, n318}, n316);
	defparam lut_246.LUT_SIZE = 4;
	defparam lut_246.mask = 16'H080F;

	lut_sub lut_247 ({n110, n111, n276, n604}, n320);
	defparam lut_247.LUT_SIZE = 4;
	defparam lut_247.mask = 16'HF351;

	lut_sub lut_248 ({i_4_, n118}, n323);
	defparam lut_248.LUT_SIZE = 2;
	defparam lut_248.mask = 4'b1011;

	lut_sub lut_249 ({i_8_, n35, n323}, n322);
	defparam lut_249.LUT_SIZE = 3;
	defparam lut_249.mask = 8'H8A;

	lut_sub lut_250 ({i_7_, i_9_}, n326);
	defparam lut_250.LUT_SIZE = 2;
	defparam lut_250.mask = 4'b1011;

	lut_sub lut_251 ({i_4_, n326}, n324);
	defparam lut_251.LUT_SIZE = 2;
	defparam lut_251.mask = 4'b1011;

	lut_sub lut_252 ({i_13_, n324, i_7_, n322}, n327);
	defparam lut_252.LUT_SIZE = 4;
	defparam lut_252.mask = 16'HEEE0;

	lut_sub lut_253 ({n339, i_4_, n316}, n330);
	defparam lut_253.LUT_SIZE = 3;
	defparam lut_253.mask = 8'HE0;

	lut_sub lut_254 ({n695, n794, i_3_, n327}, n331);
	defparam lut_254.LUT_SIZE = 4;
	defparam lut_254.mask = 16'HE000;

	lut_sub lut_255 ({i_13_, n312, n330, n331}, n328);
	defparam lut_255.LUT_SIZE = 4;
	defparam lut_255.mask = 16'H8088;

	lut_sub lut_256 ({n685, n698, n946}, n332);
	defparam lut_256.LUT_SIZE = 3;
	defparam lut_256.mask = 8'H54;

	lut_sub lut_257 ({n802, n803, i_2_, n309}, n333);
	defparam lut_257.LUT_SIZE = 4;
	defparam lut_257.mask = 16'HE000;

	lut_sub lut_258 ({i_6_, i_9_}, n335);
	defparam lut_258.LUT_SIZE = 2;
	defparam lut_258.mask = 4'b0111;

	lut_sub lut_259 ({i_6_, i_10_, n335}, n334);
	defparam lut_259.LUT_SIZE = 3;
	defparam lut_259.mask = 8'HA2;

	lut_sub lut_260 ({n398, n118}, n339);
	defparam lut_260.LUT_SIZE = 2;
	defparam lut_260.mask = 4'b1110;

	lut_sub lut_261 ({i_7_, n657, n920}, n337);
	defparam lut_261.LUT_SIZE = 3;
	defparam lut_261.mask = 8'HAC;

	lut_sub lut_262 ({i_2_, i_13_}, n338);
	defparam lut_262.LUT_SIZE = 2;
	defparam lut_262.mask = 4'b1110;

	lut_sub lut_263 ({n339, n337, n338}, n336);
	defparam lut_263.LUT_SIZE = 3;
	defparam lut_263.mask = 8'HE0;

	lut_sub lut_264 ({i_10_, i_7_}, n341);
	defparam lut_264.LUT_SIZE = 2;
	defparam lut_264.mask = 4'b1110;

	lut_sub lut_265 ({i_11_, n341}, n340);
	defparam lut_265.LUT_SIZE = 2;
	defparam lut_265.mask = 4'b1110;

	lut_sub lut_266 ({i_11_, i_13_}, n344);
	defparam lut_266.LUT_SIZE = 2;
	defparam lut_266.mask = 4'b1110;

	lut_sub lut_267 ({n185, n196, n340, n344}, n342);
	defparam lut_267.LUT_SIZE = 4;
	defparam lut_267.mask = 16'HC8FA;

	lut_sub lut_268 ({i_8_, n326}, n346);
	defparam lut_268.LUT_SIZE = 2;
	defparam lut_268.mask = 4'b1110;

	lut_sub lut_269 ({n185, n197, n344, n346}, n345);
	defparam lut_269.LUT_SIZE = 4;
	defparam lut_269.mask = 16'HE0EE;

	lut_sub lut_270 ({i_6_, n342, n345}, n349);
	defparam lut_270.LUT_SIZE = 3;
	defparam lut_270.mask = 8'HAC;

	lut_sub lut_271 ({i_8_, n657, n920}, n348);
	defparam lut_271.LUT_SIZE = 3;
	defparam lut_271.mask = 8'HAC;

	lut_sub lut_272 ({n349, i_13_, n348}, n347);
	defparam lut_272.LUT_SIZE = 3;
	defparam lut_272.mask = 8'HE0;

	lut_sub lut_273 ({i_7_, n704, n705}, n352);
	defparam lut_273.LUT_SIZE = 3;
	defparam lut_273.mask = 8'HCA;

	lut_sub lut_274 ({i_7_, n542}, n351);
	defparam lut_274.LUT_SIZE = 2;
	defparam lut_274.mask = 4'b1110;

	lut_sub lut_275 ({i_6_, i_11_, n352, n351}, n350);
	defparam lut_275.LUT_SIZE = 4;
	defparam lut_275.mask = 16'H8CCC;

	lut_sub lut_276 ({n340, i_12_, n306}, n353);
	defparam lut_276.LUT_SIZE = 3;
	defparam lut_276.mask = 8'HE0;

	lut_sub lut_277 ({i_2_, i_6_, n353, n951}, n354);
	defparam lut_277.LUT_SIZE = 4;
	defparam lut_277.mask = 16'H0051;

	lut_sub lut_278 ({i_4_, n354, n719}, n357);
	defparam lut_278.LUT_SIZE = 3;
	defparam lut_278.mask = 8'H13;

	lut_sub lut_279 ({i_2_, i_4_, n738}, n362);
	defparam lut_279.LUT_SIZE = 3;
	defparam lut_279.mask = 8'HFB;

	lut_sub lut_280 ({n199, n357, n362, n453}, n360);
	defparam lut_280.LUT_SIZE = 4;
	defparam lut_280.mask = 16'HC040;

	lut_sub lut_281 ({i_7_, n335}, n365);
	defparam lut_281.LUT_SIZE = 2;
	defparam lut_281.mask = 4'b1011;

	lut_sub lut_282 ({i_6_, i_7_}, n364);
	defparam lut_282.LUT_SIZE = 2;
	defparam lut_282.mask = 4'b1110;

	lut_sub lut_283 ({i_9_, i_10_, n365, n364}, n363);
	defparam lut_283.LUT_SIZE = 4;
	defparam lut_283.mask = 16'H0C8C;

	lut_sub lut_284 ({i_6_, n317, n674}, n367);
	defparam lut_284.LUT_SIZE = 3;
	defparam lut_284.mask = 8'H53;

	lut_sub lut_285 ({i_4_, i_11_, n367, n718}, n366);
	defparam lut_285.LUT_SIZE = 4;
	defparam lut_285.mask = 16'H00D5;

	lut_sub lut_286 ({i_3_, n347, n350}, n370);
	defparam lut_286.LUT_SIZE = 3;
	defparam lut_286.mask = 8'HAC;

	lut_sub lut_287 ({i_13_, n334, n360}, n371);
	defparam lut_287.LUT_SIZE = 3;
	defparam lut_287.mask = 8'HCA;

	lut_sub lut_288 ({i_2_, n363, n366, n816}, n372);
	defparam lut_288.LUT_SIZE = 4;
	defparam lut_288.mask = 16'H2022;

	lut_sub lut_289 ({n370, n336, n371, n372}, n369);
	defparam lut_289.LUT_SIZE = 4;
	defparam lut_289.mask = 16'H8000;

	lut_sub lut_290 ({i_3_, i_4_}, n376);
	defparam lut_290.LUT_SIZE = 2;
	defparam lut_290.mask = 4'b1011;

	lut_sub lut_291 ({n338, n376, n479, n506}, n373);
	defparam lut_291.LUT_SIZE = 4;
	defparam lut_291.mask = 16'HF531;

	lut_sub lut_292 ({i_3_, i_4_, n125, n406}, n377);
	defparam lut_292.LUT_SIZE = 4;
	defparam lut_292.mask = 16'H5F4C;

	lut_sub lut_293 ({i_3_, n287, n506, n685}, n380);
	defparam lut_293.LUT_SIZE = 4;
	defparam lut_293.mask = 16'H0B0F;

	lut_sub lut_294 ({i_2_, i_7_, n373, n664}, n381);
	defparam lut_294.LUT_SIZE = 4;
	defparam lut_294.mask = 16'H8ACF;

	lut_sub lut_295 ({n380, n381, n377, n197}, n379);
	defparam lut_295.LUT_SIZE = 4;
	defparam lut_295.mask = 16'HE000;

	lut_sub lut_296 ({i_4_, n421}, n384);
	defparam lut_296.LUT_SIZE = 2;
	defparam lut_296.mask = 4'b1000;

	lut_sub lut_297 ({i_11_, n421}, n383);
	defparam lut_297.LUT_SIZE = 2;
	defparam lut_297.mask = 4'b0010;

	lut_sub lut_298 ({i_3_, n196, n384, n383}, n382);
	defparam lut_298.LUT_SIZE = 4;
	defparam lut_298.mask = 16'H0C0E;

	lut_sub lut_299 ({i_2_, i_7_, n499}, n387);
	defparam lut_299.LUT_SIZE = 3;
	defparam lut_299.mask = 8'HDF;

	lut_sub lut_300 ({n383, n702}, n388);
	defparam lut_300.LUT_SIZE = 2;
	defparam lut_300.mask = 4'b1011;

	lut_sub lut_301 ({i_3_, n317, n479}, n389);
	defparam lut_301.LUT_SIZE = 3;
	defparam lut_301.mask = 8'HDF;

	lut_sub lut_302 ({i_2_, i_8_, n307}, n390);
	defparam lut_302.LUT_SIZE = 3;
	defparam lut_302.mask = 8'HEF;

	lut_sub lut_303 ({i_7_, n50, n376, n479}, n391);
	defparam lut_303.LUT_SIZE = 4;
	defparam lut_303.mask = 16'H0F0D;

	lut_sub lut_304 ({n382, n387, n388, n389, n390, n391}, n385);
	defparam lut_304.LUT_SIZE = 6;
	defparam lut_304.mask = 64'H0000000080000000;

	lut_sub lut_305 ({i_11_, n626, n697, n702}, n393);
	defparam lut_305.LUT_SIZE = 4;
	defparam lut_305.mask = 16'HFFDF;

	lut_sub lut_306 ({i_6_, n379, n385}, n394);
	defparam lut_306.LUT_SIZE = 3;
	defparam lut_306.mask = 8'HAC;

	lut_sub lut_307 ({n393, n394, n90, n307}, n392);
	defparam lut_307.LUT_SIZE = 4;
	defparam lut_307.mask = 16'HE000;

	lut_sub lut_308 ({i_11_, n648}, n396);
	defparam lut_308.LUT_SIZE = 2;
	defparam lut_308.mask = 4'b1011;

	lut_sub lut_309 ({n185, n604}, n397);
	defparam lut_309.LUT_SIZE = 2;
	defparam lut_309.mask = 4'b0111;

	lut_sub lut_310 ({i_4_, i_9_}, n398);
	defparam lut_310.LUT_SIZE = 2;
	defparam lut_310.mask = 4'b1011;

	lut_sub lut_311 ({n396, n397, n398, n73}, n395);
	defparam lut_311.LUT_SIZE = 4;
	defparam lut_311.mask = 16'HEEE0;

	lut_sub lut_312 ({i_3_, i_12_, n651}, n399);
	defparam lut_312.LUT_SIZE = 3;
	defparam lut_312.mask = 8'H40;

	lut_sub lut_313 ({i_1_, n45}, n402);
	defparam lut_313.LUT_SIZE = 2;
	defparam lut_313.mask = 4'b1110;

	lut_sub lut_314 ({i_11_, n185}, n403);
	defparam lut_314.LUT_SIZE = 2;
	defparam lut_314.mask = 4'b0111;

	lut_sub lut_315 ({n205, n268, n402, n403}, n401);
	defparam lut_315.LUT_SIZE = 4;
	defparam lut_315.mask = 16'HEE0E;

	lut_sub lut_316 ({i_11_, i_13_}, n406);
	defparam lut_316.LUT_SIZE = 2;
	defparam lut_316.mask = 4'b0100;

	lut_sub lut_317 ({i_4_, n402, n406, n809}, n404);
	defparam lut_317.LUT_SIZE = 4;
	defparam lut_317.mask = 16'H5D00;

	lut_sub lut_318 ({i_1_, n453}, n409);
	defparam lut_318.LUT_SIZE = 2;
	defparam lut_318.mask = 4'b0010;

	lut_sub lut_319 ({i_7_, n399, n409, n268}, n408);
	defparam lut_319.LUT_SIZE = 4;
	defparam lut_319.mask = 16'HF800;

	lut_sub lut_320 ({i_8_, n401, n921}, n411);
	defparam lut_320.LUT_SIZE = 3;
	defparam lut_320.mask = 8'H8A;

	lut_sub lut_321 ({n500, n433, n228, n700}, n412);
	defparam lut_321.LUT_SIZE = 4;
	defparam lut_321.mask = 16'HEEE0;

	lut_sub lut_322 ({n24, n42, n651, n696}, n415);
	defparam lut_322.LUT_SIZE = 4;
	defparam lut_322.mask = 16'HE0EE;

	lut_sub lut_323 ({n395, n404, n408, n411, n412, n415}, n410);
	defparam lut_323.LUT_SIZE = 6;
	defparam lut_323.mask = 64'H0000008000000000;

	lut_sub lut_324 ({i_2_, i_12_}, n417);
	defparam lut_324.LUT_SIZE = 2;
	defparam lut_324.mask = 4'b1011;

	lut_sub lut_325 ({i_8_, n42, n417, n488}, n416);
	defparam lut_325.LUT_SIZE = 4;
	defparam lut_325.mask = 16'HD0DD;

	lut_sub lut_326 ({i_12_, i_13_}, n421);
	defparam lut_326.LUT_SIZE = 2;
	defparam lut_326.mask = 4'b0100;

	lut_sub lut_327 ({i_4_, n402, n421, n813}, n419);
	defparam lut_327.LUT_SIZE = 4;
	defparam lut_327.mask = 16'H4C44;

	lut_sub lut_328 ({i_8_, n499, n700, n814}, n424);
	defparam lut_328.LUT_SIZE = 4;
	defparam lut_328.mask = 16'HAA8A;

	lut_sub lut_329 ({i_9_, n416, n419, n424}, n422);
	defparam lut_329.LUT_SIZE = 4;
	defparam lut_329.mask = 16'H2022;

	lut_sub lut_330 ({i_8_, i_9_}, n426);
	defparam lut_330.LUT_SIZE = 2;
	defparam lut_330.mask = 4'b1011;

	lut_sub lut_331 ({n205, n312, n409, n426}, n425);
	defparam lut_331.LUT_SIZE = 4;
	defparam lut_331.mask = 16'H3F2A;

	lut_sub lut_332 ({i_10_, n74}, n428);
	defparam lut_332.LUT_SIZE = 2;
	defparam lut_332.mask = 4'b1110;

	lut_sub lut_333 ({i_6_, n426}, n429);
	defparam lut_333.LUT_SIZE = 2;
	defparam lut_333.mask = 4'b1011;

	lut_sub lut_334 ({i_1_, n376}, n433);
	defparam lut_334.LUT_SIZE = 2;
	defparam lut_334.mask = 4'b1011;

	lut_sub lut_335 ({n308, n365, n433, n445}, n430);
	defparam lut_335.LUT_SIZE = 4;
	defparam lut_335.mask = 16'H54FC;

	lut_sub lut_336 ({i_4_, i_13_, n626, n713}, n434);
	defparam lut_336.LUT_SIZE = 4;
	defparam lut_336.mask = 16'H5155;

	lut_sub lut_337 ({i_6_, i_11_, n647}, n437);
	defparam lut_337.LUT_SIZE = 3;
	defparam lut_337.mask = 8'H54;

	lut_sub lut_338 ({i_3_, n226}, n445);
	defparam lut_338.LUT_SIZE = 2;
	defparam lut_338.mask = 4'b1000;

	lut_sub lut_339 ({i_6_, n522}, n448);
	defparam lut_339.LUT_SIZE = 2;
	defparam lut_339.mask = 4'b0010;

	lut_sub lut_340 ({i_9_, i_11_}, n451);
	defparam lut_340.LUT_SIZE = 2;
	defparam lut_340.mask = 4'b0111;

	lut_sub lut_341 ({i_12_, n451}, n449);
	defparam lut_341.LUT_SIZE = 2;
	defparam lut_341.mask = 4'b1011;

	lut_sub lut_342 ({i_4_, n114}, n455);
	defparam lut_342.LUT_SIZE = 2;
	defparam lut_342.mask = 4'b1011;

	lut_sub lut_343 ({i_3_, i_4_}, n453);
	defparam lut_343.LUT_SIZE = 2;
	defparam lut_343.mask = 4'b0010;

	lut_sub lut_344 ({i_9_, i_12_}, n454);
	defparam lut_344.LUT_SIZE = 2;
	defparam lut_344.mask = 4'b0111;

	lut_sub lut_345 ({n455, n453, n454}, n452);
	defparam lut_345.LUT_SIZE = 3;
	defparam lut_345.mask = 8'HE0;

	lut_sub lut_346 ({i_9_, i_13_, n712}, n457);
	defparam lut_346.LUT_SIZE = 3;
	defparam lut_346.mask = 8'H3A;

	lut_sub lut_347 ({i_3_, n109}, n458);
	defparam lut_347.LUT_SIZE = 2;
	defparam lut_347.mask = 4'b1110;

	lut_sub lut_348 ({i_2_, n99, n185}, n460);
	defparam lut_348.LUT_SIZE = 3;
	defparam lut_348.mask = 8'HFD;

	lut_sub lut_349 ({i_1_, n335, n449, n488}, n461);
	defparam lut_349.LUT_SIZE = 4;
	defparam lut_349.mask = 16'HD0DD;

	lut_sub lut_350 ({i_4_, n53, n449, n452}, n462);
	defparam lut_350.LUT_SIZE = 4;
	defparam lut_350.mask = 16'HAF8C;

	lut_sub lut_351 ({n457, n458, n460, n461, n462, n927}, n456);
	defparam lut_351.LUT_SIZE = 6;
	defparam lut_351.mask = 64'H4000000000000000;

	lut_sub lut_352 ({i_4_, n108, n186, n703}, n463);
	defparam lut_352.LUT_SIZE = 4;
	defparam lut_352.mask = 16'H005D;

	lut_sub lut_353 ({i_10_, i_13_, n226, n923}, n467);
	defparam lut_353.LUT_SIZE = 4;
	defparam lut_353.mask = 16'H0155;

	lut_sub lut_354 ({n108, n323, n463, n852}, n468);
	defparam lut_354.LUT_SIZE = 4;
	defparam lut_354.mask = 16'H2220;

	lut_sub lut_355 ({n467, n468, i_3_, n105}, n466);
	defparam lut_355.LUT_SIZE = 4;
	defparam lut_355.mask = 16'HE000;

	lut_sub lut_356 ({i_7_, n650}, n470);
	defparam lut_356.LUT_SIZE = 2;
	defparam lut_356.mask = 4'b1110;

	lut_sub lut_357 ({i_7_, n236}, n471);
	defparam lut_357.LUT_SIZE = 2;
	defparam lut_357.mask = 4'b1011;

	lut_sub lut_358 ({n470, n118, n114, n471}, n469);
	defparam lut_358.LUT_SIZE = 4;
	defparam lut_358.mask = 16'HEEE0;

	lut_sub lut_359 ({i_2_, n323, n552, n851}, n472);
	defparam lut_359.LUT_SIZE = 4;
	defparam lut_359.mask = 16'H0057;

	lut_sub lut_360 ({i_3_, i_8_, n36}, n476);
	defparam lut_360.LUT_SIZE = 3;
	defparam lut_360.mask = 8'H10;

	lut_sub lut_361 ({i_11_, i_12_}, n479);
	defparam lut_361.LUT_SIZE = 2;
	defparam lut_361.mask = 4'b0100;

	lut_sub lut_362 ({i_0_, i_2_, i_10_, n479}, n478);
	defparam lut_362.LUT_SIZE = 4;
	defparam lut_362.mask = 16'H0080;

	lut_sub lut_363 ({i_0_, n453}, n481);
	defparam lut_363.LUT_SIZE = 2;
	defparam lut_363.mask = 4'b0010;

	lut_sub lut_364 ({i_6_, n61, n478, n481}, n480);
	defparam lut_364.LUT_SIZE = 4;
	defparam lut_364.mask = 16'H00CE;

	lut_sub lut_365 ({n36, n39, n383, n499}, n485);
	defparam lut_365.LUT_SIZE = 4;
	defparam lut_365.mask = 16'HF351;

	lut_sub lut_366 ({i_0_, n21}, n483);
	defparam lut_366.LUT_SIZE = 2;
	defparam lut_366.mask = 4'b1110;

	lut_sub lut_367 ({n307, n480, n485, n483}, n482);
	defparam lut_367.LUT_SIZE = 4;
	defparam lut_367.mask = 16'H0C08;

	lut_sub lut_368 ({i_6_, i_7_, n77, n78}, n486);
	defparam lut_368.LUT_SIZE = 4;
	defparam lut_368.mask = 16'H8CAF;

	lut_sub lut_369 ({i_8_, i_3_}, n488);
	defparam lut_369.LUT_SIZE = 2;
	defparam lut_369.mask = 4'b1000;

	lut_sub lut_370 ({i_7_, n488, n497}, n487);
	defparam lut_370.LUT_SIZE = 3;
	defparam lut_370.mask = 8'H54;

	lut_sub lut_371 ({i_3_, n271, n691}, n490);
	defparam lut_371.LUT_SIZE = 3;
	defparam lut_371.mask = 8'HA3;

	lut_sub lut_372 ({i_4_, n61, n307, n490}, n489);
	defparam lut_372.LUT_SIZE = 4;
	defparam lut_372.mask = 16'H8088;

	lut_sub lut_373 ({i_12_, n712}, n492);
	defparam lut_373.LUT_SIZE = 2;
	defparam lut_373.mask = 4'b1011;

	lut_sub lut_374 ({i_2_, n50, n107, n383}, n493);
	defparam lut_374.LUT_SIZE = 4;
	defparam lut_374.mask = 16'H0F0D;

	lut_sub lut_375 ({n492, n493, n489, n108}, n491);
	defparam lut_375.LUT_SIZE = 4;
	defparam lut_375.mask = 16'HE000;

	lut_sub lut_376 ({i_7_, n451}, n494);
	defparam lut_376.LUT_SIZE = 2;
	defparam lut_376.mask = 4'b1011;

	lut_sub lut_377 ({n226, n197, i_2_, n429}, n495);
	defparam lut_377.LUT_SIZE = 4;
	defparam lut_377.mask = 16'HEEE0;

	lut_sub lut_378 ({i_1_, n557}, n497);
	defparam lut_378.LUT_SIZE = 2;
	defparam lut_378.mask = 4'b1011;

	lut_sub lut_379 ({i_6_, i_8_, n43, n497}, n496);
	defparam lut_379.LUT_SIZE = 4;
	defparam lut_379.mask = 16'H8CAF;

	lut_sub lut_380 ({i_10_, i_12_}, n499);
	defparam lut_380.LUT_SIZE = 2;
	defparam lut_380.mask = 4'b0100;

	lut_sub lut_381 ({i_0_, n226, n476, n499}, n498);
	defparam lut_381.LUT_SIZE = 4;
	defparam lut_381.mask = 16'H88A8;

	lut_sub lut_382 ({i_7_, n186}, n500);
	defparam lut_382.LUT_SIZE = 2;
	defparam lut_382.mask = 4'b1101;

	lut_sub lut_383 ({i_8_, n186, n497, n901}, n502);
	defparam lut_383.LUT_SIZE = 4;
	defparam lut_383.mask = 16'H5070;

	lut_sub lut_384 ({i_11_, i_12_}, n506);
	defparam lut_384.LUT_SIZE = 2;
	defparam lut_384.mask = 4'b0010;

	lut_sub lut_385 ({i_8_, n36, n506, n835}, n504);
	defparam lut_385.LUT_SIZE = 4;
	defparam lut_385.mask = 16'H4C44;

	lut_sub lut_386 ({i_0_, n21}, n508);
	defparam lut_386.LUT_SIZE = 2;
	defparam lut_386.mask = 4'b1011;

	lut_sub lut_387 ({n500, n502, n504, n508}, n507);
	defparam lut_387.LUT_SIZE = 4;
	defparam lut_387.mask = 16'H0302;

	lut_sub lut_388 ({i_1_, i_11_, n287, n335}, n513);
	defparam lut_388.LUT_SIZE = 4;
	defparam lut_388.mask = 16'H3233;

	lut_sub lut_389 ({n53, n529, n834, n833}, n514);
	defparam lut_389.LUT_SIZE = 4;
	defparam lut_389.mask = 16'H08CC;

	lut_sub lut_390 ({n63, n403, n513, n514}, n511);
	defparam lut_390.LUT_SIZE = 4;
	defparam lut_390.mask = 16'H8088;

	lut_sub lut_391 ({i_6_, n268, n481}, n517);
	defparam lut_391.LUT_SIZE = 3;
	defparam lut_391.mask = 8'H7F;

	lut_sub lut_392 ({i_11_, n39, n185}, n518);
	defparam lut_392.LUT_SIZE = 3;
	defparam lut_392.mask = 8'HDF;

	lut_sub lut_393 ({n223, n517, n518, n529}, n515);
	defparam lut_393.LUT_SIZE = 4;
	defparam lut_393.mask = 16'HC040;

	lut_sub lut_394 ({i_4_, i_6_, n196, n264}, n519);
	defparam lut_394.LUT_SIZE = 4;
	defparam lut_394.mask = 16'HA8AA;

	lut_sub lut_395 ({i_7_, n522}, n521);
	defparam lut_395.LUT_SIZE = 2;
	defparam lut_395.mask = 4'b0010;

	lut_sub lut_396 ({i_2_, i_12_, n521}, n520);
	defparam lut_396.LUT_SIZE = 3;
	defparam lut_396.mask = 8'H80;

	lut_sub lut_397 ({i_10_, i_11_}, n522);
	defparam lut_397.LUT_SIZE = 2;
	defparam lut_397.mask = 4'b0100;

	lut_sub lut_398 ({i_4_, i_8_, n118}, n524);
	defparam lut_398.LUT_SIZE = 3;
	defparam lut_398.mask = 8'HEF;

	lut_sub lut_399 ({n32, n276, n524}, n523);
	defparam lut_399.LUT_SIZE = 3;
	defparam lut_399.mask = 8'HA2;

	lut_sub lut_400 ({i_3_, n36, n228, n664}, n525);
	defparam lut_400.LUT_SIZE = 4;
	defparam lut_400.mask = 16'H0705;

	lut_sub lut_401 ({i_4_, n268}, n529);
	defparam lut_401.LUT_SIZE = 2;
	defparam lut_401.mask = 4'b1000;

	lut_sub lut_402 ({i_6_, n46, n520, n529}, n528);
	defparam lut_402.LUT_SIZE = 4;
	defparam lut_402.mask = 16'HCE00;

	lut_sub lut_403 ({i_4_, n507, n651, n42}, n532);
	defparam lut_403.LUT_SIZE = 4;
	defparam lut_403.mask = 16'HEEE0;

	lut_sub lut_404 ({i_0_, i_7_, n511, n515}, n533);
	defparam lut_404.LUT_SIZE = 4;
	defparam lut_404.mask = 16'HAF8C;

	lut_sub lut_405 ({n76, n322, n406, n519}, n534);
	defparam lut_405.LUT_SIZE = 4;
	defparam lut_405.mask = 16'HBBB0;

	lut_sub lut_406 ({i_1_, n448, n529, n832}, n535);
	defparam lut_406.LUT_SIZE = 4;
	defparam lut_406.mask = 16'H0BBB;

	lut_sub lut_407 ({n173, n497, n523, n830}, n537);
	defparam lut_407.LUT_SIZE = 4;
	defparam lut_407.mask = 16'HF5C4;

	lut_sub lut_408 ({n39, n125, n525, n604}, n538);
	defparam lut_408.LUT_SIZE = 4;
	defparam lut_408.mask = 16'H3331;

	lut_sub lut_409 ({n395, n528, n532, n533, n534, n535, n537, n538}, n531);
	defparam lut_409.LUT_SIZE = 8;
	defparam lut_409.mask = 256'H0000000000000000800000000000000000000000000000000000000000000000;

	lut_sub lut_410 ({i_4_, i_10_, n56, n198}, n539);
	defparam lut_410.LUT_SIZE = 4;
	defparam lut_410.mask = 16'HA8AA;

	lut_sub lut_411 ({i_9_, i_11_, i_7_}, n541);
	defparam lut_411.LUT_SIZE = 3;
	defparam lut_411.mask = 8'HFE;

	lut_sub lut_412 ({n207, n235, n541}, n540);
	defparam lut_412.LUT_SIZE = 3;
	defparam lut_412.mask = 8'HE0;

	lut_sub lut_413 ({i_8_, i_9_}, n542);
	defparam lut_413.LUT_SIZE = 2;
	defparam lut_413.mask = 4'b0111;

	lut_sub lut_414 ({i_5_, n674, n697, n708}, n543);
	defparam lut_414.LUT_SIZE = 4;
	defparam lut_414.mask = 16'H1300;

	lut_sub lut_415 ({i_10_, n653}, n548);
	defparam lut_415.LUT_SIZE = 2;
	defparam lut_415.mask = 4'b1000;

	lut_sub lut_416 ({i_4_, n548, n673, n708}, n547);
	defparam lut_416.LUT_SIZE = 4;
	defparam lut_416.mask = 16'H0031;

	lut_sub lut_417 ({i_8_, n236}, n551);
	defparam lut_417.LUT_SIZE = 2;
	defparam lut_417.mask = 4'b1011;

	lut_sub lut_418 ({i_8_, n650}, n552);
	defparam lut_418.LUT_SIZE = 2;
	defparam lut_418.mask = 4'b1110;

	lut_sub lut_419 ({n186, n454, n551, n552}, n550);
	defparam lut_419.LUT_SIZE = 4;
	defparam lut_419.mask = 16'HA8FC;

	lut_sub lut_420 ({i_12_, n174, n521, n664}, n553);
	defparam lut_420.LUT_SIZE = 4;
	defparam lut_420.mask = 16'H00DF;

	lut_sub lut_421 ({i_3_, n113, n542}, n556);
	defparam lut_421.LUT_SIZE = 3;
	defparam lut_421.mask = 8'HEF;

	lut_sub lut_422 ({i_11_, n116, n553, n556}, n554);
	defparam lut_422.LUT_SIZE = 4;
	defparam lut_422.mask = 16'H2220;

	lut_sub lut_423 ({i_0_, i_2_}, n557);
	defparam lut_423.LUT_SIZE = 2;
	defparam lut_423.mask = 4'b0111;

	lut_sub lut_424 ({i_3_, i_5_, i_6_}, n559);
	defparam lut_424.LUT_SIZE = 3;
	defparam lut_424.mask = 8'H40;

	lut_sub lut_425 ({i_7_, n479, n559, n848}, n558);
	defparam lut_425.LUT_SIZE = 4;
	defparam lut_425.mask = 16'H50D0;

	lut_sub lut_426 ({i_7_, n506, n682, n849}, n561);
	defparam lut_426.LUT_SIZE = 4;
	defparam lut_426.mask = 16'H7050;

	lut_sub lut_427 ({i_5_, n453}, n565);
	defparam lut_427.LUT_SIZE = 2;
	defparam lut_427.mask = 4'b1101;

	lut_sub lut_428 ({n104, n406, n421, n565}, n564);
	defparam lut_428.LUT_SIZE = 4;
	defparam lut_428.mask = 16'H23AF;

	lut_sub lut_429 ({i_5_, n656}, n568);
	defparam lut_429.LUT_SIZE = 2;
	defparam lut_429.mask = 4'b1110;

	lut_sub lut_430 ({n78, n568, n77, n552}, n567);
	defparam lut_430.LUT_SIZE = 4;
	defparam lut_430.mask = 16'HEEE0;

	lut_sub lut_431 ({i_5_, n653}, n570);
	defparam lut_431.LUT_SIZE = 2;
	defparam lut_431.mask = 4'b0111;

	lut_sub lut_432 ({n551, n77, n570, n78}, n569);
	defparam lut_432.LUT_SIZE = 4;
	defparam lut_432.mask = 16'HEEE0;

	lut_sub lut_433 ({n149, n508}, n572);
	defparam lut_433.LUT_SIZE = 2;
	defparam lut_433.mask = 4'b1000;

	lut_sub lut_434 ({i_0_, n376}, n573);
	defparam lut_434.LUT_SIZE = 2;
	defparam lut_434.mask = 4'b1011;

	lut_sub lut_435 ({n572, n570, n471, n573}, n571);
	defparam lut_435.LUT_SIZE = 4;
	defparam lut_435.mask = 16'HEEE0;

	lut_sub lut_436 ({i_0_, i_3_, i_5_}, n575);
	defparam lut_436.LUT_SIZE = 3;
	defparam lut_436.mask = 8'H40;

	lut_sub lut_437 ({n108, n186, n575, n823}, n574);
	defparam lut_437.LUT_SIZE = 4;
	defparam lut_437.mask = 16'H50D0;

	lut_sub lut_438 ({i_0_, i_2_, i_4_}, n578);
	defparam lut_438.LUT_SIZE = 3;
	defparam lut_438.mask = 8'H02;

	lut_sub lut_439 ({n268, n578, n709, n824}, n577);
	defparam lut_439.LUT_SIZE = 4;
	defparam lut_439.mask = 16'H3111;

	lut_sub lut_440 ({i_5_, n653}, n584);
	defparam lut_440.LUT_SIZE = 2;
	defparam lut_440.mask = 4'b0010;

	lut_sub lut_441 ({i_0_, i_1_, i_4_}, n582);
	defparam lut_441.LUT_SIZE = 3;
	defparam lut_441.mask = 8'H02;

	lut_sub lut_442 ({n268, n584, n582, n825}, n581);
	defparam lut_442.LUT_SIZE = 4;
	defparam lut_442.mask = 16'HD050;

	lut_sub lut_443 ({n61, n582, n710, n826}, n585);
	defparam lut_443.LUT_SIZE = 4;
	defparam lut_443.mask = 16'H1131;

	lut_sub lut_444 ({n61, n578, n711, n827}, n588);
	defparam lut_444.LUT_SIZE = 4;
	defparam lut_444.mask = 16'H1131;

	lut_sub lut_445 ({n308, n506, n547, n682}, n591);
	defparam lut_445.LUT_SIZE = 4;
	defparam lut_445.mask = 16'HD0C0;

	lut_sub lut_446 ({n351, n479, n543, n559}, n592);
	defparam lut_446.LUT_SIZE = 4;
	defparam lut_446.mask = 16'HC0E0;

	lut_sub lut_447 ({n550, n43, n564, n39}, n596);
	defparam lut_447.LUT_SIZE = 4;
	defparam lut_447.mask = 16'HEEE0;

	lut_sub lut_448 ({i_9_, n174, n497, n581}, n597);
	defparam lut_448.LUT_SIZE = 4;
	defparam lut_448.mask = 16'H5455;

	lut_sub lut_449 ({n874, n872, n567, n32}, n599);
	defparam lut_449.LUT_SIZE = 4;
	defparam lut_449.mask = 16'HE000;

	lut_sub lut_450 ({n871, n869, n571, n454}, n600);
	defparam lut_450.LUT_SIZE = 4;
	defparam lut_450.mask = 16'HE000;

	lut_sub lut_451 ({n876, n878, n879, n882, n884, n885, n932, n933}, n601);
	defparam lut_451.LUT_SIZE = 8;
	defparam lut_451.mask = 256'H1000000000000000000000000000000000000000000000000000000000000000;

	lut_sub lut_452 ({i_5_, n426}, n602);
	defparam lut_452.LUT_SIZE = 2;
	defparam lut_452.mask = 4'b1011;

	lut_sub lut_453 ({i_3_, i_8_}, n604);
	defparam lut_453.LUT_SIZE = 2;
	defparam lut_453.mask = 4'b0010;

	lut_sub lut_454 ({i_7_, n39, n604}, n603);
	defparam lut_454.LUT_SIZE = 3;
	defparam lut_454.mask = 8'H32;

	lut_sub lut_455 ({n736, n197, i_1_, n671}, n607);
	defparam lut_455.LUT_SIZE = 4;
	defparam lut_455.mask = 16'HEEE0;

	lut_sub lut_456 ({n402, n602, n603, n896}, n608);
	defparam lut_456.LUT_SIZE = 4;
	defparam lut_456.mask = 16'H2220;

	lut_sub lut_457 ({i_0_, i_5_, n607, n608}, n606);
	defparam lut_457.LUT_SIZE = 4;
	defparam lut_457.mask = 16'H8808;

	lut_sub lut_458 ({i_7_, n39, n276}, n609);
	defparam lut_458.LUT_SIZE = 3;
	defparam lut_458.mask = 8'H23;

	lut_sub lut_459 ({n357, i_1_, n437}, n610);
	defparam lut_459.LUT_SIZE = 3;
	defparam lut_459.mask = 8'HE0;

	lut_sub lut_460 ({n942, i_5_, n519}, n612);
	defparam lut_460.LUT_SIZE = 3;
	defparam lut_460.mask = 8'HE0;

	lut_sub lut_461 ({n203, i_3_, n348}, n613);
	defparam lut_461.LUT_SIZE = 3;
	defparam lut_461.mask = 8'HE0;

	lut_sub lut_462 ({i_12_, n39, n453, n606}, n614);
	defparam lut_462.LUT_SIZE = 4;
	defparam lut_462.mask = 16'HF3A2;

	lut_sub lut_463 ({n235, n714, n232, n353}, n615);
	defparam lut_463.LUT_SIZE = 4;
	defparam lut_463.mask = 16'HEEE0;

	lut_sub lut_464 ({n898, i_1_, n437, n668}, n616);
	defparam lut_464.LUT_SIZE = 4;
	defparam lut_464.mask = 16'HFE00;

	lut_sub lut_465 ({n899, i_11_, n894, n891}, n617);
	defparam lut_465.LUT_SIZE = 4;
	defparam lut_465.mask = 16'HF800;

	lut_sub lut_466 ({n539, n540, n612, n613, n614, n615, n616, n617}, n611);
	defparam lut_466.LUT_SIZE = 8;
	defparam lut_466.mask = 256'H8000000000000000000000000000000000000000000000000000000000000000;

	lut_sub lut_467 ({i_7_, n454}, n620);
	defparam lut_467.LUT_SIZE = 2;
	defparam lut_467.mask = 4'b1011;

	lut_sub lut_468 ({i_10_, i_12_}, n619);
	defparam lut_468.LUT_SIZE = 2;
	defparam lut_468.mask = 4'b0111;

	lut_sub lut_469 ({i_7_, n620, n619, n626}, n618);
	defparam lut_469.LUT_SIZE = 4;
	defparam lut_469.mask = 16'H5040;

	lut_sub lut_470 ({i_5_, n943, n944}, n622);
	defparam lut_470.LUT_SIZE = 3;
	defparam lut_470.mask = 8'HAC;

	lut_sub lut_471 ({i_0_, n334, n622}, n621);
	defparam lut_471.LUT_SIZE = 3;
	defparam lut_471.mask = 8'H8A;

	lut_sub lut_472 ({i_8_, i_11_}, n624);
	defparam lut_472.LUT_SIZE = 2;
	defparam lut_472.mask = 4'b1101;

	lut_sub lut_473 ({i_3_, n312, n624, n626}, n623);
	defparam lut_473.LUT_SIZE = 4;
	defparam lut_473.mask = 16'H0040;

	lut_sub lut_474 ({i_8_, i_12_}, n626);
	defparam lut_474.LUT_SIZE = 2;
	defparam lut_474.mask = 4'b1000;

	lut_sub lut_475 ({n240, n471, n626}, n625);
	defparam lut_475.LUT_SIZE = 3;
	defparam lut_475.mask = 8'H2A;

	lut_sub lut_476 ({i_1_, n237, n618, n621}, n628);
	defparam lut_476.LUT_SIZE = 4;
	defparam lut_476.mask = 16'HA8FC;

	lut_sub lut_477 ({i_12_, n41, n905, n909}, n629);
	defparam lut_477.LUT_SIZE = 4;
	defparam lut_477.mask = 16'H80AA;

	lut_sub lut_478 ({i_11_, n900, n904, n908}, n630);
	defparam lut_478.LUT_SIZE = 4;
	defparam lut_478.mask = 16'H80AA;

	lut_sub lut_479 ({n906, n624, n250, n470}, n631);
	defparam lut_479.LUT_SIZE = 4;
	defparam lut_479.mask = 16'HF800;

	lut_sub lut_480 ({n628, n629, n630, n631}, n627);
	defparam lut_480.LUT_SIZE = 4;
	defparam lut_480.mask = 16'H8000;

	lut_sub lut_481 ({i_12_, n604}, n633);
	defparam lut_481.LUT_SIZE = 2;
	defparam lut_481.mask = 4'b1101;

	lut_sub lut_482 ({i_11_, n23, n276, n633}, n632);
	defparam lut_482.LUT_SIZE = 4;
	defparam lut_482.mask = 16'H0A02;

	lut_sub lut_483 ({n114, n276, n406, n488}, n635);
	defparam lut_483.LUT_SIZE = 4;
	defparam lut_483.mask = 16'H3F15;

	lut_sub lut_484 ({n50, n276, n287, n604}, n637);
	defparam lut_484.LUT_SIZE = 4;
	defparam lut_484.mask = 16'H153F;

	lut_sub lut_485 ({i_4_, n632, n635}, n638);
	defparam lut_485.LUT_SIZE = 3;
	defparam lut_485.mask = 8'HAC;

	lut_sub lut_486 ({i_13_, n23, n910, n911}, n639);
	defparam lut_486.LUT_SIZE = 4;
	defparam lut_486.mask = 16'H0888;

	lut_sub lut_487 ({n637, n638, n639}, n636);
	defparam lut_487.LUT_SIZE = 3;
	defparam lut_487.mask = 8'H80;

	lut_sub lut_488 ({i_1_, i_2_, n312, n334}, n641);
	defparam lut_488.LUT_SIZE = 4;
	defparam lut_488.mask = 16'H8ACF;

	lut_sub lut_489 ({i_5_, i_9_, i_10_}, n640);
	defparam lut_489.LUT_SIZE = 3;
	defparam lut_489.mask = 8'H35;

	lut_sub lut_490 ({i_6_, i_12_}, n647);
	defparam lut_490.LUT_SIZE = 2;
	defparam lut_490.mask = 4'b0100;

	lut_sub lut_491 ({i_9_, n487, n647, i_1_}, n646);
	defparam lut_491.LUT_SIZE = 4;
	defparam lut_491.mask = 16'HF800;

	lut_sub lut_492 ({i_9_, i_10_}, n648);
	defparam lut_492.LUT_SIZE = 2;
	defparam lut_492.mask = 4'b1110;

	lut_sub lut_493 ({i_3_, i_4_}, n649);
	defparam lut_493.LUT_SIZE = 2;
	defparam lut_493.mask = 4'b1110;

	lut_sub lut_494 ({i_5_, i_6_}, n650);
	defparam lut_494.LUT_SIZE = 2;
	defparam lut_494.mask = 4'b1110;

	lut_sub lut_495 ({i_8_, n522}, n651);
	defparam lut_495.LUT_SIZE = 2;
	defparam lut_495.mask = 4'b1101;

	lut_sub lut_496 ({i_8_, n38}, n652);
	defparam lut_496.LUT_SIZE = 2;
	defparam lut_496.mask = 4'b1011;

	lut_sub lut_497 ({i_8_, i_7_}, n653);
	defparam lut_497.LUT_SIZE = 2;
	defparam lut_497.mask = 4'b1000;

	lut_sub lut_498 ({i_8_, n364}, n654);
	defparam lut_498.LUT_SIZE = 2;
	defparam lut_498.mask = 4'b1011;

	lut_sub lut_499 ({i_0_, i_1_, i_2_}, n655);
	defparam lut_499.LUT_SIZE = 3;
	defparam lut_499.mask = 8'HBF;

	lut_sub lut_500 ({i_8_, i_7_}, n656);
	defparam lut_500.LUT_SIZE = 2;
	defparam lut_500.mask = 4'b1110;

	lut_sub lut_501 ({i_11_, n648}, n657);
	defparam lut_501.LUT_SIZE = 2;
	defparam lut_501.mask = 4'b1110;

	lut_sub lut_502 ({i_5_, n649}, n658);
	defparam lut_502.LUT_SIZE = 2;
	defparam lut_502.mask = 4'b1011;

	lut_sub lut_503 ({n421, n657}, n659);
	defparam lut_503.LUT_SIZE = 2;
	defparam lut_503.mask = 4'b1011;

	lut_sub lut_504 ({i_9_, i_10_}, n660);
	defparam lut_504.LUT_SIZE = 2;
	defparam lut_504.mask = 4'b0111;

	lut_sub lut_505 ({i_7_, n660}, n661);
	defparam lut_505.LUT_SIZE = 2;
	defparam lut_505.mask = 4'b1110;

	lut_sub lut_506 ({i_3_, n660}, n662);
	defparam lut_506.LUT_SIZE = 2;
	defparam lut_506.mask = 4'b1011;

	lut_sub lut_507 ({i_7_, n660}, n663);
	defparam lut_507.LUT_SIZE = 2;
	defparam lut_507.mask = 4'b1011;

	lut_sub lut_508 ({i_11_, n313}, n664);
	defparam lut_508.LUT_SIZE = 2;
	defparam lut_508.mask = 4'b1110;

	lut_sub lut_509 ({i_3_, i_4_, i_5_}, n665);
	defparam lut_509.LUT_SIZE = 3;
	defparam lut_509.mask = 8'H7F;

	lut_sub lut_510 ({i_6_, n398}, n666);
	defparam lut_510.LUT_SIZE = 2;
	defparam lut_510.mask = 4'b1011;

	lut_sub lut_511 ({i_8_, n398}, n667);
	defparam lut_511.LUT_SIZE = 2;
	defparam lut_511.mask = 4'b1011;

	lut_sub lut_512 ({i_5_, i_10_}, n668);
	defparam lut_512.LUT_SIZE = 2;
	defparam lut_512.mask = 4'b1110;

	lut_sub lut_513 ({i_7_, n668}, n669);
	defparam lut_513.LUT_SIZE = 2;
	defparam lut_513.mask = 4'b1110;

	lut_sub lut_514 ({i_2_, n453}, n670);
	defparam lut_514.LUT_SIZE = 2;
	defparam lut_514.mask = 4'b0010;

	lut_sub lut_515 ({i_9_, n236}, n671);
	defparam lut_515.LUT_SIZE = 2;
	defparam lut_515.mask = 4'b1110;

	lut_sub lut_516 ({i_5_, n398}, n672);
	defparam lut_516.LUT_SIZE = 2;
	defparam lut_516.mask = 4'b1011;

	lut_sub lut_517 ({i_5_, i_6_}, n673);
	defparam lut_517.LUT_SIZE = 2;
	defparam lut_517.mask = 4'b1101;

	lut_sub lut_518 ({i_9_, n656}, n674);
	defparam lut_518.LUT_SIZE = 2;
	defparam lut_518.mask = 4'b1011;

	lut_sub lut_519 ({n287, n674}, n675);
	defparam lut_519.LUT_SIZE = 2;
	defparam lut_519.mask = 4'b1011;

	lut_sub lut_520 ({n50, n308}, n677);
	defparam lut_520.LUT_SIZE = 2;
	defparam lut_520.mask = 4'b0111;

	lut_sub lut_521 ({n268, n565}, n680);
	defparam lut_521.LUT_SIZE = 2;
	defparam lut_521.mask = 4'b1011;

	lut_sub lut_522 ({n287, n351}, n681);
	defparam lut_522.LUT_SIZE = 2;
	defparam lut_522.mask = 4'b1011;

	lut_sub lut_523 ({i_3_, n673}, n682);
	defparam lut_523.LUT_SIZE = 2;
	defparam lut_523.mask = 4'b1011;

	lut_sub lut_524 ({i_3_, n650}, n683);
	defparam lut_524.LUT_SIZE = 2;
	defparam lut_524.mask = 4'b1011;

	lut_sub lut_525 ({i_3_, n236}, n684);
	defparam lut_525.LUT_SIZE = 2;
	defparam lut_525.mask = 4'b1011;

	lut_sub lut_526 ({i_7_, n542}, n685);
	defparam lut_526.LUT_SIZE = 2;
	defparam lut_526.mask = 4'b1011;

	lut_sub lut_527 ({n287, n685}, n686);
	defparam lut_527.LUT_SIZE = 2;
	defparam lut_527.mask = 4'b1011;

	lut_sub lut_528 ({n50, n317}, n687);
	defparam lut_528.LUT_SIZE = 2;
	defparam lut_528.mask = 4'b1011;

	lut_sub lut_529 ({n287, n318}, n688);
	defparam lut_529.LUT_SIZE = 2;
	defparam lut_529.mask = 4'b1011;

	lut_sub lut_530 ({i_13_, n116}, n690);
	defparam lut_530.LUT_SIZE = 2;
	defparam lut_530.mask = 4'b1110;

	lut_sub lut_531 ({i_11_, n499}, n691);
	defparam lut_531.LUT_SIZE = 2;
	defparam lut_531.mask = 4'b0111;

	lut_sub lut_532 ({i_13_, n174}, n692);
	defparam lut_532.LUT_SIZE = 2;
	defparam lut_532.mask = 4'b1110;

	lut_sub lut_533 ({i_9_, n506}, n693);
	defparam lut_533.LUT_SIZE = 2;
	defparam lut_533.mask = 4'b0111;

	lut_sub lut_534 ({n112, n662}, n695);
	defparam lut_534.LUT_SIZE = 2;
	defparam lut_534.mask = 4'b1000;

	lut_sub lut_535 ({i_2_, i_3_}, n696);
	defparam lut_535.LUT_SIZE = 2;
	defparam lut_535.mask = 4'b0111;

	lut_sub lut_536 ({i_4_, i_6_}, n697);
	defparam lut_536.LUT_SIZE = 2;
	defparam lut_536.mask = 4'b1110;

	lut_sub lut_537 ({i_3_, i_12_}, n698);
	defparam lut_537.LUT_SIZE = 2;
	defparam lut_537.mask = 4'b1011;

	lut_sub lut_538 ({i_4_, n247}, n699);
	defparam lut_538.LUT_SIZE = 2;
	defparam lut_538.mask = 4'b1110;

	lut_sub lut_539 ({i_1_, n696}, n700);
	defparam lut_539.LUT_SIZE = 2;
	defparam lut_539.mask = 4'b1110;

	lut_sub lut_540 ({i_1_, n45}, n701);
	defparam lut_540.LUT_SIZE = 2;
	defparam lut_540.mask = 4'b1011;

	lut_sub lut_541 ({i_7_, i_2_}, n702);
	defparam lut_541.LUT_SIZE = 2;
	defparam lut_541.mask = 4'b1110;

	lut_sub lut_542 ({i_11_, n619}, n703);
	defparam lut_542.LUT_SIZE = 2;
	defparam lut_542.mask = 4'b1011;

	lut_sub lut_543 ({i_9_, n619}, n704);
	defparam lut_543.LUT_SIZE = 2;
	defparam lut_543.mask = 4'b1011;

	lut_sub lut_544 ({i_9_, n186}, n705);
	defparam lut_544.LUT_SIZE = 2;
	defparam lut_544.mask = 4'b0111;

	lut_sub lut_545 ({i_8_, n341}, n707);
	defparam lut_545.LUT_SIZE = 2;
	defparam lut_545.mask = 4'b1011;

	lut_sub lut_546 ({i_0_, n696}, n708);
	defparam lut_546.LUT_SIZE = 2;
	defparam lut_546.mask = 4'b1110;

	lut_sub lut_547 ({i_8_, n673}, n709);
	defparam lut_547.LUT_SIZE = 2;
	defparam lut_547.mask = 4'b1011;

	lut_sub lut_548 ({i_5_, n656}, n710);
	defparam lut_548.LUT_SIZE = 2;
	defparam lut_548.mask = 4'b1011;

	lut_sub lut_549 ({i_5_, n74}, n711);
	defparam lut_549.LUT_SIZE = 2;
	defparam lut_549.mask = 4'b1011;

	lut_sub lut_550 ({n241, n344}, n712);
	defparam lut_550.LUT_SIZE = 2;
	defparam lut_550.mask = 4'b1011;

	lut_sub lut_551 ({n276, n383}, n713);
	defparam lut_551.LUT_SIZE = 2;
	defparam lut_551.mask = 4'b1000;

	lut_sub lut_552 ({i_12_, n326}, n714);
	defparam lut_552.LUT_SIZE = 2;
	defparam lut_552.mask = 4'b1110;

	lut_sub lut_553 ({i_5_, n499, n522}, n716);
	defparam lut_553.LUT_SIZE = 3;
	defparam lut_553.mask = 8'HCA;

	lut_sub lut_554 ({i_4_, n82, n912}, n717);
	defparam lut_554.LUT_SIZE = 3;
	defparam lut_554.mask = 8'HCA;

	lut_sub lut_555 ({i_6_, n449, n703}, n718);
	defparam lut_555.LUT_SIZE = 3;
	defparam lut_555.mask = 8'HCA;

	lut_sub lut_556 ({i_6_, n196, n197}, n719);
	defparam lut_556.LUT_SIZE = 3;
	defparam lut_556.mask = 8'H53;

	lut_sub lut_557 ({i_10_, i_13_, n479, n654}, n722);
	defparam lut_557.LUT_SIZE = 4;
	defparam lut_557.mask = 16'HFFFB;

	lut_sub lut_558 ({n256, n280, n722}, n720);
	defparam lut_558.LUT_SIZE = 3;
	defparam lut_558.mask = 8'HA2;

	lut_sub lut_559 ({i_9_, i_13_, n98, n506}, n725);
	defparam lut_559.LUT_SIZE = 4;
	defparam lut_559.mask = 16'HFFFD;

	lut_sub lut_560 ({n95, n271, n725}, n723);
	defparam lut_560.LUT_SIZE = 3;
	defparam lut_560.mask = 8'HA2;

	lut_sub lut_561 ({i_3_, n251, n661}, n727);
	defparam lut_561.LUT_SIZE = 3;
	defparam lut_561.mask = 8'HEF;

	lut_sub lut_562 ({n727, i_8_, n250, n660}, n726);
	defparam lut_562.LUT_SIZE = 4;
	defparam lut_562.mask = 16'HFE00;

	lut_sub lut_563 ({n231, n232, n448, n651}, n728);
	defparam lut_563.LUT_SIZE = 4;
	defparam lut_563.mask = 16'HFA32;

	lut_sub lut_564 ({n228, n235, n243, n728}, n730);
	defparam lut_564.LUT_SIZE = 4;
	defparam lut_564.mask = 16'H2220;

	lut_sub lut_565 ({n20, n224, n508, n684}, n733);
	defparam lut_565.LUT_SIZE = 4;
	defparam lut_565.mask = 16'H8000;

	lut_sub lut_566 ({i_0_, n227, n733, n663}, n732);
	defparam lut_566.LUT_SIZE = 4;
	defparam lut_566.mask = 16'HEEE0;

	lut_sub lut_567 ({n223, n218, n215}, n736);
	defparam lut_567.LUT_SIZE = 3;
	defparam lut_567.mask = 8'H80;

	lut_sub lut_568 ({n221, n521, n664, n736}, n734);
	defparam lut_568.LUT_SIZE = 4;
	defparam lut_568.mask = 16'HEE0E;

	lut_sub lut_569 ({n429, n428}, n738);
	defparam lut_569.LUT_SIZE = 2;
	defparam lut_569.mask = 4'b1000;

	lut_sub lut_570 ({n46, n666, n324, n223}, n740);
	defparam lut_570.LUT_SIZE = 4;
	defparam lut_570.mask = 16'HEEE0;

	lut_sub lut_571 ({n675, n217}, n742);
	defparam lut_571.LUT_SIZE = 2;
	defparam lut_571.mask = 4'b1110;

	lut_sub lut_572 ({n168, n174, n114}, n743);
	defparam lut_572.LUT_SIZE = 3;
	defparam lut_572.mask = 8'HFE;

	lut_sub lut_573 ({n108, n174, n499}, n744);
	defparam lut_573.LUT_SIZE = 3;
	defparam lut_573.mask = 8'HFD;

	lut_sub lut_574 ({n559, n687}, n745);
	defparam lut_574.LUT_SIZE = 2;
	defparam lut_574.mask = 4'b1011;

	lut_sub lut_575 ({n559, n686}, n746);
	defparam lut_575.LUT_SIZE = 2;
	defparam lut_575.mask = 4'b1011;

	lut_sub lut_576 ({n140, n174, n114}, n747);
	defparam lut_576.LUT_SIZE = 3;
	defparam lut_576.mask = 8'HFE;

	lut_sub lut_577 ({n217, n308, n653, n684}, n748);
	defparam lut_577.LUT_SIZE = 4;
	defparam lut_577.mask = 16'HAF23;

	lut_sub lut_578 ({n662, n683, n317}, n749);
	defparam lut_578.LUT_SIZE = 3;
	defparam lut_578.mask = 8'HE0;

	lut_sub lut_579 ({n53, n114, n665}, n751);
	defparam lut_579.LUT_SIZE = 3;
	defparam lut_579.mask = 8'HEF;

	lut_sub lut_580 ({n751, n115, n108}, n750);
	defparam lut_580.LUT_SIZE = 3;
	defparam lut_580.mask = 8'HE0;

	lut_sub lut_581 ({n220, n165, n98, n145}, n752);
	defparam lut_581.LUT_SIZE = 4;
	defparam lut_581.mask = 16'HEEE0;

	lut_sub lut_582 ({n750, n752, n217, n688}, n753);
	defparam lut_582.LUT_SIZE = 4;
	defparam lut_582.mask = 16'HE000;

	lut_sub lut_583 ({n109, n658, n105, n124}, n754);
	defparam lut_583.LUT_SIZE = 4;
	defparam lut_583.mask = 16'HEEE0;

	lut_sub lut_584 ({i_4_, n119, n695, n754}, n755);
	defparam lut_584.LUT_SIZE = 4;
	defparam lut_584.mask = 16'H0A08;

	lut_sub lut_585 ({n36, n654, n652, n40}, n757);
	defparam lut_585.LUT_SIZE = 4;
	defparam lut_585.mask = 16'HEEE0;

	lut_sub lut_586 ({n89, n92, n181, n565}, n758);
	defparam lut_586.LUT_SIZE = 4;
	defparam lut_586.mask = 16'HFA32;

	lut_sub lut_587 ({n97, n100, n665, n758}, n759);
	defparam lut_587.LUT_SIZE = 4;
	defparam lut_587.mask = 16'H0A08;

	lut_sub lut_588 ({n602, n259, n671, n260}, n761);
	defparam lut_588.LUT_SIZE = 4;
	defparam lut_588.mask = 16'HEEE0;

	lut_sub lut_589 ({n672, n42, n324, n508}, n762);
	defparam lut_589.LUT_SIZE = 4;
	defparam lut_589.mask = 16'HEEE0;

	lut_sub lut_590 ({i_6_, i_11_, n44}, n764);
	defparam lut_590.LUT_SIZE = 3;
	defparam lut_590.mask = 8'HEF;

	lut_sub lut_591 ({i_10_, n41, n764}, n763);
	defparam lut_591.LUT_SIZE = 3;
	defparam lut_591.mask = 8'H8A;

	lut_sub lut_592 ({i_10_, n102, n383, n654}, n766);
	defparam lut_592.LUT_SIZE = 4;
	defparam lut_592.mask = 16'HFFBF;

	lut_sub lut_593 ({n766, n37, n179}, n765);
	defparam lut_593.LUT_SIZE = 3;
	defparam lut_593.mask = 8'HE0;

	lut_sub lut_594 ({i_10_, n173, n383, n652}, n768);
	defparam lut_594.LUT_SIZE = 4;
	defparam lut_594.mask = 16'HFFFB;

	lut_sub lut_595 ({n768, n26, n40, n125}, n767);
	defparam lut_595.LUT_SIZE = 4;
	defparam lut_595.mask = 16'HFE00;

	lut_sub lut_596 ({n767, n654, n655, n32}, n769);
	defparam lut_596.LUT_SIZE = 4;
	defparam lut_596.mask = 16'HFE00;

	lut_sub lut_597 ({n30, n34, n53, n101}, n770);
	defparam lut_597.LUT_SIZE = 4;
	defparam lut_597.mask = 16'HF351;

	lut_sub lut_598 ({n101, n125, n178, n668}, n772);
	defparam lut_598.LUT_SIZE = 4;
	defparam lut_598.mask = 16'HFEFF;

	lut_sub lut_599 ({i_4_, n42, n716, n772}, n771);
	defparam lut_599.LUT_SIZE = 4;
	defparam lut_599.mask = 16'HAAA2;

	lut_sub lut_600 ({n51, n116, n769, n770}, n773);
	defparam lut_600.LUT_SIZE = 4;
	defparam lut_600.mask = 16'H00F8;

	lut_sub lut_601 ({i_10_, n402, i_2_, n428}, n775);
	defparam lut_601.LUT_SIZE = 4;
	defparam lut_601.mask = 16'HEEE0;

	lut_sub lut_602 ({n42, n697, i_11_, n317}, n777);
	defparam lut_602.LUT_SIZE = 4;
	defparam lut_602.mask = 16'HFFFE;

	lut_sub lut_603 ({n777, i_9_, n258, n73}, n776);
	defparam lut_603.LUT_SIZE = 4;
	defparam lut_603.mask = 16'HFE00;

	lut_sub lut_604 ({i_2_, n61, n429}, n779);
	defparam lut_604.LUT_SIZE = 3;
	defparam lut_604.mask = 8'HEF;

	lut_sub lut_605 ({n779, n241, n61, n197}, n778);
	defparam lut_605.LUT_SIZE = 4;
	defparam lut_605.mask = 16'HFE00;

	lut_sub lut_606 ({i_10_, n296, n398}, n781);
	defparam lut_606.LUT_SIZE = 3;
	defparam lut_606.mask = 8'HFB;

	lut_sub lut_607 ({n185, n253, n396, n781}, n780);
	defparam lut_607.LUT_SIZE = 4;
	defparam lut_607.mask = 16'HA8AA;

	lut_sub lut_608 ({i_13_, n470, n651, n780}, n782);
	defparam lut_608.LUT_SIZE = 4;
	defparam lut_608.mask = 16'HA8AA;

	lut_sub lut_609 ({n212, n268, n665}, n785);
	defparam lut_609.LUT_SIZE = 3;
	defparam lut_609.mask = 8'HFB;

	lut_sub lut_610 ({n102, n192, n292, n785}, n783);
	defparam lut_610.LUT_SIZE = 4;
	defparam lut_610.mask = 16'H2022;

	lut_sub lut_611 ({n187, n173, n169, n655}, n788);
	defparam lut_611.LUT_SIZE = 4;
	defparam lut_611.mask = 16'HEEE0;

	lut_sub lut_612 ({n788, n163, n36}, n789);
	defparam lut_612.LUT_SIZE = 3;
	defparam lut_612.mask = 8'HE0;

	lut_sub lut_613 ({n156, n40, n143, n31}, n790);
	defparam lut_613.LUT_SIZE = 4;
	defparam lut_613.mask = 16'HEEE0;

	lut_sub lut_614 ({n790, n789, n131, n39}, n791);
	defparam lut_614.LUT_SIZE = 4;
	defparam lut_614.mask = 16'HE000;

	lut_sub lut_615 ({n297, n497, n753, n755}, n792);
	defparam lut_615.LUT_SIZE = 4;
	defparam lut_615.mask = 16'H00F8;

	lut_sub lut_616 ({i_7_, n320, n914}, n794);
	defparam lut_616.LUT_SIZE = 3;
	defparam lut_616.mask = 8'H8A;

	lut_sub lut_617 ({i_4_, n73, n542}, n796);
	defparam lut_617.LUT_SIZE = 3;
	defparam lut_617.mask = 8'HDF;

	lut_sub lut_618 ({n796, i_8_, i_13_, n260}, n795);
	defparam lut_618.LUT_SIZE = 4;
	defparam lut_618.mask = 16'HFE00;

	lut_sub lut_619 ({i_11_, n178, n406, n670}, n797);
	defparam lut_619.LUT_SIZE = 4;
	defparam lut_619.mask = 16'H7770;

	lut_sub lut_620 ({i_8_, i_13_, n260}, n799);
	defparam lut_620.LUT_SIZE = 3;
	defparam lut_620.mask = 8'HEF;

	lut_sub lut_621 ({n421, n667, n670, n799}, n798);
	defparam lut_621.LUT_SIZE = 4;
	defparam lut_621.mask = 16'H20AA;

	lut_sub lut_622 ({i_2_, n312, n376}, n802);
	defparam lut_622.LUT_SIZE = 3;
	defparam lut_622.mask = 8'HEF;

	lut_sub lut_623 ({i_7_, n795, n797, n916}, n803);
	defparam lut_623.LUT_SIZE = 4;
	defparam lut_623.mask = 16'H5540;

	lut_sub lut_624 ({n448, n626, n702}, n805);
	defparam lut_624.LUT_SIZE = 3;
	defparam lut_624.mask = 8'H7F;

	lut_sub lut_625 ({n805, n437, n700}, n804);
	defparam lut_625.LUT_SIZE = 3;
	defparam lut_625.mask = 8'HE0;

	lut_sub lut_626 ({n185, n344, n428, n429}, n806);
	defparam lut_626.LUT_SIZE = 4;
	defparam lut_626.mask = 16'HA8FC;

	lut_sub lut_627 ({i_3_, i_6_, i_8_, i_10_, n185, n945}, n808);
	defparam lut_627.LUT_SIZE = 6;
	defparam lut_627.mask = 64'HFFFFFFFFFFFFFBFF;

	lut_sub lut_628 ({n421, n425, n808}, n807);
	defparam lut_628.LUT_SIZE = 3;
	defparam lut_628.mask = 8'H8A;

	lut_sub lut_629 ({n945, n624, i_10_, i_13_}, n810);
	defparam lut_629.LUT_SIZE = 4;
	defparam lut_629.mask = 16'HFFFE;

	lut_sub lut_630 ({n810, n118, n701}, n809);
	defparam lut_630.LUT_SIZE = 3;
	defparam lut_630.mask = 8'HE0;

	lut_sub lut_631 ({i_10_, i_8_}, n812);
	defparam lut_631.LUT_SIZE = 2;
	defparam lut_631.mask = 4'b1110;

	lut_sub lut_632 ({n205, n341, n409, n812}, n813);
	defparam lut_632.LUT_SIZE = 4;
	defparam lut_632.mask = 16'HF3A2;

	lut_sub lut_633 ({i_8_, n383, n402}, n814);
	defparam lut_633.LUT_SIZE = 3;
	defparam lut_633.mask = 8'HFB;

	lut_sub lut_634 ({i_6_, i_12_, n453, n685}, n816);
	defparam lut_634.LUT_SIZE = 4;
	defparam lut_634.mask = 16'HEFFF;

	lut_sub lut_635 ({i_3_, i_9_, n479, n652}, n818);
	defparam lut_635.LUT_SIZE = 4;
	defparam lut_635.mask = 16'HBFFF;

	lut_sub lut_636 ({n334, n626, n699, n818}, n817);
	defparam lut_636.LUT_SIZE = 4;
	defparam lut_636.mask = 16'HAA8A;

	lut_sub lut_637 ({n417, n365, n434, n99}, n819);
	defparam lut_637.LUT_SIZE = 4;
	defparam lut_637.mask = 16'HEEE0;

	lut_sub lut_638 ({i_6_, n410, n422}, n821);
	defparam lut_638.LUT_SIZE = 3;
	defparam lut_638.mask = 8'HAC;

	lut_sub lut_639 ({i_1_, n369, n392}, n822);
	defparam lut_639.LUT_SIZE = 3;
	defparam lut_639.mask = 8'HCA;

	lut_sub lut_640 ({i_12_, n430, n821, n822}, n820);
	defparam lut_640.LUT_SIZE = 4;
	defparam lut_640.mask = 16'H8088;

	lut_sub lut_641 ({n572, n568, n470, n573}, n823);
	defparam lut_641.LUT_SIZE = 4;
	defparam lut_641.mask = 16'HEEE0;

	lut_sub lut_642 ({n46, n280, n693, n708}, n824);
	defparam lut_642.LUT_SIZE = 4;
	defparam lut_642.mask = 16'HEE0E;

	lut_sub lut_643 ({n223, n280, n483, n693}, n825);
	defparam lut_643.LUT_SIZE = 4;
	defparam lut_643.mask = 16'HEE0E;

	lut_sub lut_644 ({n223, n271, n483, n691}, n826);
	defparam lut_644.LUT_SIZE = 4;
	defparam lut_644.mask = 16'HEE0E;

	lut_sub lut_645 ({n46, n271, n691, n708}, n827);
	defparam lut_645.LUT_SIZE = 4;
	defparam lut_645.mask = 16'HEE0E;

	lut_sub lut_646 ({n185, n209, n344, n669}, n828);
	defparam lut_646.LUT_SIZE = 4;
	defparam lut_646.mask = 16'HE0EE;

	lut_sub lut_647 ({n104, n114, n118, n565}, n829);
	defparam lut_647.LUT_SIZE = 4;
	defparam lut_647.mask = 16'HE0EE;

	lut_sub lut_648 ({i_3_, i_7_, i_8_, i_10_}, n830);
	defparam lut_648.LUT_SIZE = 4;
	defparam lut_648.mask = 16'H2A0A;

	lut_sub lut_649 ({i_8_, n39}, n832);
	defparam lut_649.LUT_SIZE = 2;
	defparam lut_649.mask = 4'b1011;

	lut_sub lut_650 ({i_2_, n365, n506, n934}, n834);
	defparam lut_650.LUT_SIZE = 4;
	defparam lut_650.mask = 16'HA2AA;

	lut_sub lut_651 ({i_3_, n280, n693}, n833);
	defparam lut_651.LUT_SIZE = 3;
	defparam lut_651.mask = 8'HA3;

	lut_sub lut_652 ({i_0_, i_7_, n53, n483}, n835);
	defparam lut_652.LUT_SIZE = 4;
	defparam lut_652.mask = 16'HAF23;

	lut_sub lut_653 ({i_8_, n36, n479}, n838);
	defparam lut_653.LUT_SIZE = 3;
	defparam lut_653.mask = 8'HFD;

	lut_sub lut_654 ({n838, n496, n454}, n837);
	defparam lut_654.LUT_SIZE = 3;
	defparam lut_654.mask = 8'HE0;

	lut_sub lut_655 ({i_8_, n114, n173}, n841);
	defparam lut_655.LUT_SIZE = 3;
	defparam lut_655.mask = 8'HEF;

	lut_sub lut_656 ({n421, n495, n841}, n840);
	defparam lut_656.LUT_SIZE = 3;
	defparam lut_656.mask = 8'H8A;

	lut_sub lut_657 ({i_6_, n494, n417}, n844);
	defparam lut_657.LUT_SIZE = 3;
	defparam lut_657.mask = 8'HFE;

	lut_sub lut_658 ({n844, n486, n455}, n843);
	defparam lut_658.LUT_SIZE = 3;
	defparam lut_658.mask = 8'HE0;

	lut_sub lut_659 ({n173, n276, n320, n659}, n845);
	defparam lut_659.LUT_SIZE = 4;
	defparam lut_659.mask = 16'HAF8C;

	lut_sub lut_660 ({n39, n713, n843, n845}, n846);
	defparam lut_660.LUT_SIZE = 4;
	defparam lut_660.mask = 16'H8808;

	lut_sub lut_661 ({i_0_, n491, i_7_, n482}, n847);
	defparam lut_661.LUT_SIZE = 4;
	defparam lut_661.mask = 16'HEEE0;

	lut_sub lut_662 ({i_1_, i_2_, n710, n711}, n848);
	defparam lut_662.LUT_SIZE = 4;
	defparam lut_662.mask = 16'H8CAF;

	lut_sub lut_663 ({i_1_, i_2_, n584, n709}, n849);
	defparam lut_663.LUT_SIZE = 4;
	defparam lut_663.mask = 16'H23AF;

	lut_sub lut_664 ({n106, n671, n455, n551}, n851);
	defparam lut_664.LUT_SIZE = 4;
	defparam lut_664.mask = 16'HEEE0;

	lut_sub lut_665 ({i_2_, n107, n344}, n852);
	defparam lut_665.LUT_SIZE = 3;
	defparam lut_665.mask = 8'HFE;

	lut_sub lut_666 ({n455, n570, n568, n323}, n854);
	defparam lut_666.LUT_SIZE = 4;
	defparam lut_666.mask = 16'HEEE0;

	lut_sub lut_667 ({i_10_, n106, n234}, n857);
	defparam lut_667.LUT_SIZE = 3;
	defparam lut_667.mask = 8'HFE;

	lut_sub lut_668 ({i_9_, n670, n703, n857}, n856);
	defparam lut_668.LUT_SIZE = 4;
	defparam lut_668.mask = 16'HA8AA;

	lut_sub lut_669 ({n453, n469, n472, n856}, n858);
	defparam lut_669.LUT_SIZE = 4;
	defparam lut_669.mask = 16'H2022;

	lut_sub lut_670 ({i_13_, n348, i_3_}, n863);
	defparam lut_670.LUT_SIZE = 3;
	defparam lut_670.mask = 8'HFE;

	lut_sub lut_671 ({i_6_, i_12_, n663, n922}, n862);
	defparam lut_671.LUT_SIZE = 4;
	defparam lut_671.mask = 16'H8AAA;

	lut_sub lut_672 ({i_3_, n336, n863, n862}, n861);
	defparam lut_672.LUT_SIZE = 4;
	defparam lut_672.mask = 16'H80C0;

	lut_sub lut_673 ({i_5_, n456, n466}, n867);
	defparam lut_673.LUT_SIZE = 3;
	defparam lut_673.mask = 8'HCA;

	lut_sub lut_674 ({i_1_, n660, n867, n930}, n865);
	defparam lut_674.LUT_SIZE = 4;
	defparam lut_674.mask = 16'H4044;

	lut_sub lut_675 ({i_8_, n575, n703}, n870);
	defparam lut_675.LUT_SIZE = 3;
	defparam lut_675.mask = 8'HFB;

	lut_sub lut_676 ({n870, n232, n306, n403}, n869);
	defparam lut_676.LUT_SIZE = 4;
	defparam lut_676.mask = 16'HFE00;

	lut_sub lut_677 ({i_10_, n116, n497}, n871);
	defparam lut_677.LUT_SIZE = 3;
	defparam lut_677.mask = 8'HEF;

	lut_sub lut_678 ({n219, n125, n707}, n873);
	defparam lut_678.LUT_SIZE = 3;
	defparam lut_678.mask = 8'HFE;

	lut_sub lut_679 ({n873, n569, n110}, n872);
	defparam lut_679.LUT_SIZE = 3;
	defparam lut_679.mask = 8'HE0;

	lut_sub lut_680 ({n215, n346, n383}, n874);
	defparam lut_680.LUT_SIZE = 3;
	defparam lut_680.mask = 8'HFD;

	lut_sub lut_681 ({n173, n588, n828, n829}, n876);
	defparam lut_681.LUT_SIZE = 4;
	defparam lut_681.mask = 16'H0F08;

	lut_sub lut_682 ({n239, n704, n554, n36}, n878);
	defparam lut_682.LUT_SIZE = 4;
	defparam lut_682.mask = 16'HEEE0;

	lut_sub lut_683 ({n151, n550, n591, n592}, n879);
	defparam lut_683.LUT_SIZE = 4;
	defparam lut_683.mask = 16'H1110;

	lut_sub lut_684 ({n296, n421, n539, n540}, n882);
	defparam lut_684.LUT_SIZE = 4;
	defparam lut_684.mask = 16'H8CAF;

	lut_sub lut_685 ({n705, n249, n672, n61}, n884);
	defparam lut_685.LUT_SIZE = 4;
	defparam lut_685.mask = 16'HEEE0;

	lut_sub lut_686 ({n647, n500, n557, i_5_}, n886);
	defparam lut_686.LUT_SIZE = 4;
	defparam lut_686.mask = 16'HFFFE;

	lut_sub lut_687 ({i_5_, n531, n886, n940}, n885);
	defparam lut_687.LUT_SIZE = 4;
	defparam lut_687.mask = 16'H4440;

	lut_sub lut_688 ({n221, n196, n736, n346}, n890);
	defparam lut_688.LUT_SIZE = 4;
	defparam lut_688.mask = 16'HEEE0;

	lut_sub lut_689 ({n46, n428, n609, n890}, n891);
	defparam lut_689.LUT_SIZE = 4;
	defparam lut_689.mask = 16'H2220;

	lut_sub lut_690 ({n231, n428, n204, n402}, n893);
	defparam lut_690.LUT_SIZE = 4;
	defparam lut_690.mask = 16'HEEE0;

	lut_sub lut_691 ({i_5_, i_9_, n241}, n895);
	defparam lut_691.LUT_SIZE = 3;
	defparam lut_691.mask = 8'HDF;

	lut_sub lut_692 ({n895, n893, i_0_, i_5_}, n894);
	defparam lut_692.LUT_SIZE = 4;
	defparam lut_692.mask = 16'HE000;

	lut_sub lut_693 ({n44, n429, n221, n707}, n896);
	defparam lut_693.LUT_SIZE = 4;
	defparam lut_693.mask = 16'HEEE0;

	lut_sub lut_694 ({i_10_, n398}, n898);
	defparam lut_694.LUT_SIZE = 2;
	defparam lut_694.mask = 4'b1110;

	lut_sub lut_695 ({i_0_, n610, i_2_, n337}, n899);
	defparam lut_695.LUT_SIZE = 4;
	defparam lut_695.mask = 16'HEEE0;

	lut_sub lut_696 ({i_6_, n43}, n901);
	defparam lut_696.LUT_SIZE = 2;
	defparam lut_696.mask = 4'b1110;

	lut_sub lut_697 ({i_5_, i_12_, n42, n901}, n900);
	defparam lut_697.LUT_SIZE = 4;
	defparam lut_697.mask = 16'H0A08;

	lut_sub lut_698 ({i_3_, i_7_, n251}, n903);
	defparam lut_698.LUT_SIZE = 3;
	defparam lut_698.mask = 8'HEF;

	lut_sub lut_699 ({n903, i_7_, n508}, n902);
	defparam lut_699.LUT_SIZE = 3;
	defparam lut_699.mask = 8'HE0;

	lut_sub lut_700 ({i_2_, i_7_, n683, n902}, n904);
	defparam lut_700.LUT_SIZE = 4;
	defparam lut_700.mask = 16'H88A8;

	lut_sub lut_701 ({i_2_, i_7_, n684, n733}, n905);
	defparam lut_701.LUT_SIZE = 4;
	defparam lut_701.mask = 16'H8CAF;

	lut_sub lut_702 ({n246, n494, n500, n625}, n906);
	defparam lut_702.LUT_SIZE = 4;
	defparam lut_702.mask = 16'H5540;

	lut_sub lut_703 ({i_0_, n640}, n908);
	defparam lut_703.LUT_SIZE = 2;
	defparam lut_703.mask = 4'b1011;

	lut_sub lut_704 ({n623, n497}, n909);
	defparam lut_704.LUT_SIZE = 2;
	defparam lut_704.mask = 4'b1110;

	lut_sub lut_705 ({i_3_, n323, n542}, n910);
	defparam lut_705.LUT_SIZE = 3;
	defparam lut_705.mask = 8'HDF;

	lut_sub lut_706 ({i_8_, n421, n453}, n911);
	defparam lut_706.LUT_SIZE = 3;
	defparam lut_706.mask = 8'H7F;

	lut_sub lut_707 ({i_5_, n42, n647, n685}, n912);
	defparam lut_707.LUT_SIZE = 4;
	defparam lut_707.mask = 16'HFBFF;

	lut_sub lut_708 ({i_7_, n32, n276}, n914);
	defparam lut_708.LUT_SIZE = 3;
	defparam lut_708.mask = 8'HFD;

	lut_sub lut_709 ({i_7_, n713, n50}, n915);
	defparam lut_709.LUT_SIZE = 3;
	defparam lut_709.mask = 8'HE0;

	lut_sub lut_710 ({i_7_, i_12_, n178, n798}, n916);
	defparam lut_710.LUT_SIZE = 4;
	defparam lut_710.mask = 16'H5700;

	lut_sub lut_711 ({i_12_, n648}, n920);
	defparam lut_711.LUT_SIZE = 2;
	defparam lut_711.mask = 4'b1110;

	lut_sub lut_712 ({i_8_, n186, n699}, n921);
	defparam lut_712.LUT_SIZE = 3;
	defparam lut_712.mask = 8'HFB;

	lut_sub lut_713 ({i_6_, i_11_, n661}, n922);
	defparam lut_713.LUT_SIZE = 3;
	defparam lut_713.mask = 8'HFB;

	lut_sub lut_714 ({i_10_, n63, n185, n712}, n923);
	defparam lut_714.LUT_SIZE = 4;
	defparam lut_714.mask = 16'H00D5;

	lut_sub lut_715 ({i_2_, i_12_, n365, n494}, n927);
	defparam lut_715.LUT_SIZE = 4;
	defparam lut_715.mask = 16'H7000;

	lut_sub lut_716 ({i_1_, n185, n671, n854}, n930);
	defparam lut_716.LUT_SIZE = 4;
	defparam lut_716.mask = 16'H0075;

	lut_sub lut_717 ({i_0_, i_4_, n558, n561}, n932);
	defparam lut_717.LUT_SIZE = 4;
	defparam lut_717.mask = 16'H000E;

	lut_sub lut_718 ({i_0_, n858, n861, n865}, n933);
	defparam lut_718.LUT_SIZE = 4;
	defparam lut_718.mask = 16'H7F00;

	lut_sub lut_719 ({n99, n125, i_2_}, n934);
	defparam lut_719.LUT_SIZE = 3;
	defparam lut_719.mask = 8'HFE;

	lut_sub lut_720 ({i_4_, n56, n61, n840}, n935);
	defparam lut_720.LUT_SIZE = 4;
	defparam lut_720.mask = 16'H5700;

	lut_sub lut_721 ({i_4_, n508, n620, n837}, n937);
	defparam lut_721.LUT_SIZE = 4;
	defparam lut_721.mask = 16'H0057;

	lut_sub lut_722 ({n498, n646, n846, n847, n935, n937}, n941);
	defparam lut_722.LUT_SIZE = 6;
	defparam lut_722.mask = 64'HFFFFFFFFFFFFEFFF;

	lut_sub lut_723 ({i_5_, n941}, n940);
	defparam lut_723.LUT_SIZE = 2;
	defparam lut_723.mask = 4'b1000;

	lut_sub lut_724 ({i_4_, i_5_, n495}, n942);
	defparam lut_724.LUT_SIZE = 3;
	defparam lut_724.mask = 8'HBF;

	lut_sub lut_725 ({i_6_, n186, n451}, n943);
	defparam lut_725.LUT_SIZE = 3;
	defparam lut_725.mask = 8'HA3;

	lut_sub lut_726 ({i_6_, n454, n619}, n944);
	defparam lut_726.LUT_SIZE = 3;
	defparam lut_726.mask = 8'HCA;

	lut_sub lut_727 ({i_2_, i_7_}, n945);
	defparam lut_727.LUT_SIZE = 2;
	defparam lut_727.mask = 4'b1000;

	lut_sub lut_728 ({n667, i_3_, n521}, n946);
	defparam lut_728.LUT_SIZE = 3;
	defparam lut_728.mask = 8'H80;

	lut_sub lut_729 ({n714, n541, i_6_}, n951);
	defparam lut_729.LUT_SIZE = 3;
	defparam lut_729.mask = 8'H80;

endmodule


module lut_sub (din, out);
	parameter LUT_SIZE = 4;
	parameter NUM_BITS = 2**LUT_SIZE;

	input[LUT_SIZE - 1:0] din;

	oupput out;

	wire out;

	// buffer the LUT inputs...
	wire[LUT_SIZE - 1:0] din_w;

	genvar i;
	generate
		for (i = 0; i < LUT_SIZE; i = i + 1)
			begin: liloop
			lut_input li_buf(din[i], din_w[i]);
		end
	endgenerate

	// build up the pterms for the LUT
	wire[NUM_BITS - 1:0] pterms;
	generate
		for (i = 0; i < NUM_BITS; i = i + 1)
			begin: ploop
			assign pterms[i] = ((din_w == i) & mask[i]);
		end
	endgenerate

	// assign the pterms to the LUT function
	wire result;
	assign result = | pterms;
	lut_output lo_buf (result, out);
endmodule