module clma (
	Pi416, Pi415, Pi414, Pi413, Pi412, Pi411, Pi410, Pi409, 
	Pi408, Pi407, Pi406, Pi405, Pi404, Pi403, Pi402, Pi401, Pi400, Pi399, 
	Pi398, Pi397, Pi396, Pi395, Pi394, Pi393, Pi392, Pi391, Pi390, Pi389, 
	Pi388, Pi387, Pi386, Pi385, Pi384, Pi383, Pi382, Pi381, Pi380, Pi379, 
	Pi378, Pi377, Pi376, Pi375, Pi374, Pi373, Pi372, Pi371, Pi370, Pi369, 
	Pi368, Pi367, Pi366, Pi365, Pi364, Pi363, Pi362, Pi361, Pi360, Pi359, 
	Pi358, Pi357, Pi356, Pi355, Pi354, Pi353, Pi352, Pi351, Pi350, Pi349, 
	Pi348, Pi347, Pi346, Pi345, Pi344, Pi343, Pi342, Pi341, Pi340, Pi339, 
	Pi338, Pi337, Pi336, Pi335, Pi334, Pi333, Pi332, Pi331, Pi330, Pi329, 
	Pi328, Pi327, Pi326, Pi325, Pi324, Pi323, Pi322, Pi321, Pi320, Pi319, 
	Pi318, Pi317, Pi316, Pi315, Pi314, Pi313, Pi312, Pi311, Pi310, Pi309, 
	Pi308, Pi307, Pi306, Pi305, Pi304, Pi303, Pi302, Pi301, Pi300, Pi299, 
	Pi298, Pi297, Pi296, Pi295, Pi294, Pi293, Pi292, Pi291, Pi290, Pi289, 
	Pi288, Pi287, Pi286, Pi285, Pi284, Pi283, Pi282, Pi281, Pi280, Pi279, 
	Pi278, Pi277, Pi276, Pi275, Pi274, Pi273, Pi272, Pi271, Pi270, Pi269, 
	Pi268, Pi267, Pi266, Pi265, Pi264, Pi263, Pi262, Pi261, Pi260, Pi259, 
	Pi258, Pi257, Pi256, Pi255, Pi254, Pi253, Pi252, Pi251, Pi250, Pi249, 
	Pi248, Pi247, Pi246, Pi245, Pi244, Pi243, Pi242, Pi241, Pi240, Pi239, 
	Pi238, Pi237, Pi236, Pi235, Pi234, Pi233, Pi232, Pi231, Pi230, Pi229, 
	Pi228, Pi227, Pi226, Pi225, Pi224, Pi223, Pi222, Pi221, Pi220, Pi219, 
	Pi218, Pi217, Pi216, Pi215, Pi214, Pi213, Pi212, Pi211, Pi210, Pi209, 
	Pi208, Pi207, Pi206, Pi205, Pi204, Pi203, Pi202, Pi201, Pi200, Pi199, 
	Pi198, Pi197, Pi196, Pi195, Pi194, Pi193, Pi192, Pi191, Pi190, Pi189, 
	Pi188, Pi187, Pi186, Pi185, Pi184, Pi183, Pi182, Pi181, Pi180, Pi179, 
	Pi178, Pi177, Pi176, Pi175, Pi174, Pi173, Pi172, Pi171, Pi170, Pi169, 
	Pi168, Pi167, Pi166, Pi165, Pi164, Pi163, Pi162, Pi161, Pi160, Pi159, 
	Pi158, Pi157, Pi156, Pi155, Pi154, Pi153, Pi152, Pi151, Pi150, Pi149, 
	Pi148, Pi147, Pi146, Pi145, Pi144, Pi143, Pi142, Pi141, Pi140, Pi139, 
	Pi138, Pi137, Pi136, Pi135, Pi134, Pi133, Pi132, Pi131, Pi130, Pi129, 
	Pi128, Pi127, Pi126, Pi125, Pi124, Pi123, Pi122, Pi121, Pi120, Pi119, 
	Pi118, Pi117, Pi116, Pi115, Pi114, Pi113, Pi112, Pi111, Pi110, Pi109, 
	Pi108, Pi107, Pi106, Pi105, Pi104, Pi103, Pi102, Pi101, Pi100, Pi99, 
	Pi98, Pi97, Pi96, Pi95, Pi94, Pi93, Pi92, Pi91, Pi90, Pi89, 
	Pi88, Pi87, Pi86, Pi85, Pi84, Pi83, Pi82, Pi81, Pi80, Pi79, 
	Pi78, Pi77, Pi76, Pi75, Pi74, Pi73, Pi72, Pi71, Pi70, Pi69, 
	Pi68, Pi67, Pi66, Pi65, Pi64, Pi63, Pi62, Pi61, Pi60, Pi59, 
	Pi58, Pi57, Pi56, Pi55, Pi54, Pi53, Pi52, Pi51, Pi50, Pi49, 
	Pi28, Pi27, Pi26, Pi25, Pi24, Pi23, Pi22, Pi21, Pi20, Pi19, 
	Pi18, Pi17, Pi16, Pi15, PCLK, P__cmxir_1, P__cmxir_0, P__cmxig_1, P__cmxig_0, P__cmxcl_1, 
	P__cmxcl_0, P__cmx1ad_35, P__cmx1ad_34, P__cmx1ad_33, P__cmx1ad_32, P__cmx1ad_31, P__cmx1ad_30, P__cmx1ad_29, P__cmx1ad_28, P__cmx1ad_27, 
	P__cmx1ad_26, P__cmx1ad_25, P__cmx1ad_24, P__cmx1ad_23, P__cmx1ad_22, P__cmx1ad_21, P__cmx1ad_20, P__cmx1ad_19, P__cmx1ad_18, P__cmx1ad_17, 
	P__cmx1ad_16, P__cmx1ad_15, P__cmx1ad_14, P__cmx1ad_13, P__cmx1ad_12, P__cmx1ad_11, P__cmx1ad_10, P__cmx1ad_9, P__cmx1ad_8, P__cmx1ad_7, 
	P__cmx1ad_6, P__cmx1ad_5, P__cmx1ad_4, P__cmx1ad_3, P__cmx1ad_2, P__cmx1ad_1, P__cmx1ad_0, P__cmx0ad_35, P__cmx0ad_34, P__cmx0ad_33, 
	P__cmx0ad_32, P__cmx0ad_31, P__cmx0ad_30, P__cmx0ad_29, P__cmx0ad_28, P__cmx0ad_27, P__cmx0ad_26, P__cmx0ad_25, P__cmx0ad_24, P__cmx0ad_23, 
	P__cmx0ad_22, P__cmx0ad_21, P__cmx0ad_20, P__cmx0ad_19, P__cmx0ad_18, P__cmx0ad_17, P__cmx0ad_16, P__cmx0ad_15, P__cmx0ad_14, P__cmx0ad_13, 
	P__cmx0ad_12, P__cmx0ad_11, P__cmx0ad_10, P__cmx0ad_9, P__cmx0ad_8, P__cmx0ad_7, P__cmx0ad_6, P__cmx0ad_5, P__cmx0ad_4, P__cmx0ad_3, 
	P__cmx0ad_2, P__cmx0ad_1, P__cmx0ad_0, P__cmnxcp_1, P__cmnxcp_0, P__cmndst1p0, P__cmndst0p0);

input Pi416, Pi415, Pi414, Pi413, Pi412, Pi411, Pi410, Pi409, Pi408, Pi407, Pi406, Pi405, Pi404, Pi403, Pi402, Pi401, Pi400, Pi399, Pi398, Pi397, Pi396, Pi395, Pi394, Pi393, Pi392, Pi391, Pi390, Pi389, Pi388, Pi387, Pi386, Pi385, Pi384, Pi383, Pi382, Pi381, Pi380, Pi379, Pi378, Pi377, Pi376, Pi375, Pi374, Pi373, Pi372, Pi371, Pi370, Pi369, Pi368, Pi367, Pi366, Pi365, Pi364, Pi363, Pi362, Pi361, Pi360, Pi359, Pi358, Pi357, Pi356, Pi355, Pi354, Pi353, Pi352, Pi351, Pi350, Pi349, Pi348, Pi347, Pi346, Pi345, Pi344, Pi343, Pi342, Pi341, Pi340, Pi339, Pi338, Pi337, Pi336, Pi335, Pi334, Pi333, Pi332, Pi331, Pi330, Pi329, Pi328, Pi327, Pi326, Pi325, Pi324, Pi323, Pi322, Pi321, Pi320, Pi319, Pi318, Pi317, Pi316, Pi315, Pi314, Pi313, Pi312, Pi311, Pi310, Pi309, Pi308, Pi307, Pi306, Pi305, Pi304, Pi303, Pi302, Pi301, Pi300, Pi299, Pi298, Pi297, Pi296, Pi295, Pi294, Pi293, Pi292, Pi291, Pi290, Pi289, Pi288, Pi287, Pi286, Pi285, Pi284, Pi283, Pi282, Pi281, Pi280, Pi279, Pi278, Pi277, Pi276, Pi275, Pi274, Pi273, Pi272, Pi271, Pi270, Pi269, Pi268, Pi267, Pi266, Pi265, Pi264, Pi263, Pi262, Pi261, Pi260, Pi259, Pi258, Pi257, Pi256, Pi255, Pi254, Pi253, Pi252, Pi251, Pi250, Pi249, Pi248, Pi247, Pi246, Pi245, Pi244, Pi243, Pi242, Pi241, Pi240, Pi239, Pi238, Pi237, Pi236, Pi235, Pi234, Pi233, Pi232, Pi231, Pi230, Pi229, Pi228, Pi227, Pi226, Pi225, Pi224, Pi223, Pi222, Pi221, Pi220, Pi219, Pi218, Pi217, Pi216, Pi215, Pi214, Pi213, Pi212, Pi211, Pi210, Pi209, Pi208, Pi207, Pi206, Pi205, Pi204, Pi203, Pi202, Pi201, Pi200, Pi199, Pi198, Pi197, Pi196, Pi195, Pi194, Pi193, Pi192, Pi191, Pi190, Pi189, Pi188, Pi187, Pi186, Pi185, Pi184, Pi183, Pi182, Pi181, Pi180, Pi179, Pi178, Pi177, Pi176, Pi175, Pi174, Pi173, Pi172, Pi171, Pi170, Pi169, Pi168, Pi167, Pi166, Pi165, Pi164, Pi163, Pi162, Pi161, Pi160, Pi159, Pi158, Pi157, Pi156, Pi155, Pi154, Pi153, Pi152, Pi151, Pi150, Pi149, Pi148, Pi147, Pi146, Pi145, Pi144, Pi143, Pi142, Pi141, Pi140, Pi139, Pi138, Pi137, Pi136, Pi135, Pi134, Pi133, Pi132, Pi131, Pi130, Pi129, Pi128, Pi127, Pi126, Pi125, Pi124, Pi123, Pi122, Pi121, Pi120, Pi119, Pi118, Pi117, Pi116, Pi115, Pi114, Pi113, Pi112, Pi111, Pi110, Pi109, Pi108, Pi107, Pi106, Pi105, Pi104, Pi103, Pi102, Pi101, Pi100, Pi99, Pi98, Pi97, Pi96, Pi95, Pi94, Pi93, Pi92, Pi91, Pi90, Pi89, Pi88, Pi87, Pi86, Pi85, Pi84, Pi83, Pi82, Pi81, Pi80, Pi79, Pi78, Pi77, Pi76, Pi75, Pi74, Pi73, Pi72, Pi71, Pi70, Pi69, Pi68, Pi67, Pi66, Pi65, Pi64, Pi63, Pi62, Pi61, Pi60, Pi59, Pi58, Pi57, Pi56, Pi55, Pi54, Pi53, Pi52, Pi51, Pi50, Pi49, Pi28, Pi27, Pi26, Pi25, Pi24, Pi23, Pi22, Pi21, Pi20, Pi19, Pi18, Pi17, Pi16, Pi15, PCLK;

output P__cmxir_1, P__cmxir_0, P__cmxig_1, P__cmxig_0, P__cmxcl_1, P__cmxcl_0, P__cmx1ad_35, P__cmx1ad_34, P__cmx1ad_33, P__cmx1ad_32, P__cmx1ad_31, P__cmx1ad_30, P__cmx1ad_29, P__cmx1ad_28, P__cmx1ad_27, P__cmx1ad_26, P__cmx1ad_25, P__cmx1ad_24, P__cmx1ad_23, P__cmx1ad_22, P__cmx1ad_21, P__cmx1ad_20, P__cmx1ad_19, P__cmx1ad_18, P__cmx1ad_17, P__cmx1ad_16, P__cmx1ad_15, P__cmx1ad_14, P__cmx1ad_13, P__cmx1ad_12, P__cmx1ad_11, P__cmx1ad_10, P__cmx1ad_9, P__cmx1ad_8, P__cmx1ad_7, P__cmx1ad_6, P__cmx1ad_5, P__cmx1ad_4, P__cmx1ad_3, P__cmx1ad_2, P__cmx1ad_1, P__cmx1ad_0, P__cmx0ad_35, P__cmx0ad_34, P__cmx0ad_33, P__cmx0ad_32, P__cmx0ad_31, P__cmx0ad_30, P__cmx0ad_29, P__cmx0ad_28, P__cmx0ad_27, P__cmx0ad_26, P__cmx0ad_25, P__cmx0ad_24, P__cmx0ad_23, P__cmx0ad_22, P__cmx0ad_21, P__cmx0ad_20, P__cmx0ad_19, P__cmx0ad_18, P__cmx0ad_17, P__cmx0ad_16, P__cmx0ad_15, P__cmx0ad_14, P__cmx0ad_13, P__cmx0ad_12, P__cmx0ad_11, P__cmx0ad_10, P__cmx0ad_9, P__cmx0ad_8, P__cmx0ad_7, P__cmx0ad_6, P__cmx0ad_5, P__cmx0ad_4, P__cmx0ad_3, P__cmx0ad_2, P__cmx0ad_1, P__cmx0ad_0, P__cmnxcp_1, P__cmnxcp_0, P__cmndst1p0, P__cmndst0p0;

wire n19, Nv2, n20, n21, Nv31, n22, Nv59, n25, n24, n23, n26, Nv243, n27, Nv294, n28, Nv345, n29, n30, n31, n32, n34, Nv349, n35, Nv499, n36, Nv550, n37, Nv601, n38, n42, n44, n45, n43, n46, Nv2153, n47, Nv3888, n48, n49, Nv6425, n50, Nv6437, n55, n52, n53, n51, n60, n59, n58, n64, n65, n62, n63, n61, n68, n69, n67, n66, n72, n73, n71, n70, n76, n77, n75, n74, n80, n79, n78, n83, n82, n81, n86, n85, n84, n89, n90, n88, n87, n93, n94, n92, n91, n97, n98, n96, n95, n101, n102, n100, n99, n105, n104, n103, n108, n107, n106, n109, n111, n110, n114, n113, n116, n115, n118, n117, n119, n120, n122, n121, n124, n123, n126, n125, n128, n127, n130, n129, n133, n132, n134, n135, n136, Nv10056, n137, Nv10068, n140, n138, n142, Nv10112, n143, Nv10126, n144, Nv10143, n145, n149, Nv10247, n150, n153, n157, n158, n159, n160, n161, n162, N_N13960, n163, n166, n164, n168, n167, n171, n169, n173, n177, n178, n176, n180, n179, n183, n184, n188, n190, n193, n192, n195, n196, n194, n200, n198, n197, n202, n201, n203, n206, n205, n207, n212, n210, n211, n209, n214, n213, n216, n215, n218, n217, n220, n221, n219, n223, n222, n225, n224, n227, n226, n229, n230, n228, n231, n234, n233, n232, n236, n235, n238, n237, n240, n239, n241, n243, n242, n244, n247, n246, n249, n248, n251, n250, n252, n254, n255, n253, n257, n256, n259, n258, n260, n262, n263, n261, n264, n266, n265, n267, n269, n268, n272, n271, n273, n275, n276, n274, n278, n277, n281, n279, n282, n290, n287, n288, n286, n291, n294, n292, n295, n297, n296, n299, n298, n301, n300, n304, n303, n308, n307, n311, n312, n310, n309, n313, n315, n314, n316, n317, n319, n318, n320, n322, n321, n323, n324, n326, n327, n325, n329, n328, n330, n331, n333, n334, n332, n335, n337, n336, n338, n340, n339, n341, n342, n344, n343, n346, n345, n347, n348, n350, n351, n349, n353, n352, n354, n355, n357, n358, n356, n359, n361, n360, n362, n363, n364, n366, n367, n368, n370, n371, n377, n375, n374, n378, n379, n381, n384, n383, n386, n387, n385, n388, n390, n391, n389, n394, n393, n392, n396, n397, n395, n399, n400, n398, n401, n403, n402, n404, n405, n407, n406, n408, n409, n410, n412, n411, n413, n415, n416, n414, n417, n418, n420, n423, n422, n425, n426, n424, n427, n428, n429, n430, n432, n431, n433, n434, n435, n436, n437, n439, n438, n440, n442, n443, n441, n444, n445, n447, n450, n449, n452, n453, n451, n455, n454, n457, n456, n458, n463, n464, n462, n466, n470, n471, n469, n473, n478, n476, n479, n481, n480, n483, n482, n484, n488, n487, n490, n494, n493, n496, n501, n499, n502, n504, n503, n505, n506, n508, n507, n510, n511, n509, n513, n512, n514, n515, n517, n518, n516, n520, n519, n521, n522, n524, n525, n523, n526, n528, n527, n529, n531, n530, n532, n533, n535, n534, n536, n538, n537, n539, n540, n542, n543, n541, n545, n544, n546, n547, n549, n550, n548, n551, n553, n552, n554, n555, n557, n559, n560, n562, n561, n564, n563, n565, n568, n567, n570, n573, n572, n575, n580, n578, n581, n583, n582, n585, n584, n586, n589, n588, n591, n594, n593, n596, n601, n599, n602, n604, n603, n605, n606, n608, n607, n610, n609, n611, n612, n614, n615, n613, n617, n616, n618, n619, n621, n622, n620, n623, n625, n624, n626, n628, n627, n629, n630, n632, n631, n634, n633, n635, n636, n638, n639, n637, n641, n640, n642, n643, n645, n646, n644, n647, n649, n648, n650, n651, n653, n655, n656, n658, n660, n661, n657, n663, n662, n666, n665, n664, n669, n668, n667, n670, n675, n673, n676, n677, n678, n679, n680, n685, n683, n686, n687, n688, n690, n691, n689, n693, n694, n692, n695, n697, n696, n698, n699, n700, n701, n702, n703, n705, n704, n706, n707, n709, n711, n712, n713, n714, n715, n716, n721, n719, n722, n723, n724, n725, n726, n731, n729, n732, n733, n734, n735, n736, n738, n737, n739, n740, n741, n742, n743, n745, n744, n746, n747, n749, n751, n752, n754, n756, n757, n753, n759, n758, n764, n763, n769, n768, n774, n775, n776, n777, n773, n779, n778, n782, n783, n784, n785, n781, n788, n787, n786, n791, n789, n794, n792, n797, n798, n796, n795, n801, n799, n804, n802, n807, n805, n809, n810, n808, n812, n811, n815, n813, n818, n816, n820, n821, n819, n824, n822, n827, n825, n830, n828, n832, n833, n831, n835, n834, n837, n836, n841, n840, n839, n843, n842, n845, n844, n848, n849, n847, n846, n851, n850, n853, n852, n855, n854, n858, n857, n856, n860, n859, n862, n861, n864, n863, n867, n866, n865, n869, n868, n871, n870, n873, n872, n876, n875, n874, n878, n879, n877, n881, n880, n882, n884, n883, n886, n885, n888, n887, n892, n893, n890, n891, n889, n895, n894, n897, n896, n899, n898, n901, n900, n904, n905, n903, n902, n907, n906, n909, n908, n911, n910, n913, n912, n916, n917, n915, n914, n919, n918, n921, n920, n923, n922, n925, n924, n928, n929, n927, n926, n931, n933, n934, n930, n935, n941, n940, n939, n943, n942, n945, n946, n944, n949, n950, n948, n947, n953, n954, n952, n951, n957, n956, n955, n960, n958, n963, n961, n966, n964, n969, n967, n972, n970, n975, n973, n978, n976, n981, n979, n984, n982, n987, n985, n990, n988, n993, n991, n995, n996, n997, n998, n994, n999, n1003, n1007, n1008, n1009, n1010, n1006, n1013, n1011, n1016, n1014, n1019, n1017, n1022, n1020, n1025, n1023, n1028, n1026, n1031, n1029, n1034, n1032, n1037, n1035, n1040, n1038, n1043, n1041, n1046, n1044, n1049, n1047, n1052, n1050, n1054, n1055, n1053, n1056, n1059, n1063, n1062, n1066, n1069, n1068, n1067, n1074, n1071, n1075, n1079, n1084, n1088, n1089, n1087, n1090, n1093, n1094, n1092, n1091, n1096, n1097, n1095, n1099, n1100, n1098, n1102, n1103, n1101, n1105, n1106, n1104, n1108, n1109, n1107, n1111, n1112, n1110, n1114, n1115, n1113, n1117, n1118, n1116, n1120, n1121, n1119, n1123, n1124, n1122, n1126, n1127, n1125, n1129, n1130, n1128, n1132, n1133, n1131, n1135, n1136, n1134, n1138, n1139, n1137, n1141, n1142, n1140, n1145, n1144, n1146, n1152, n1150, n1149, n1153, n1158, n1159, n1157, n1156, n1161, n1162, n1160, n1164, n1165, n1163, n1167, n1168, n1166, n1170, n1171, n1169, n1173, n1174, n1172, n1176, n1177, n1175, n1179, n1180, n1178, n1182, n1183, n1181, n1185, n1186, n1184, n1188, n1189, n1187, n1191, n1192, n1190, n1194, n1195, n1193, n1197, n1198, n1196, n1200, n1201, n1199, n1203, n1204, n1202, n1206, n1207, n1205, n1210, n1209, n1211, n1214, n1212, n1215, n1218, n1221, n1220, n1219, n1224, n1223, n1222, n1227, n1226, n1225, n1230, n1229, n1228, n1233, n1234, n1232, n1231, n1237, n1238, n1236, n1235, n1241, n1242, n1240, n1239, n1245, n1246, n1244, n1243, n1248, n1249, n1250, n1247, n1252, n1251, n1254, n1253, n1256, n1257, n1255, n1259, n1260, n1258, n1262, n1263, n1261, n1266, n1265, n1264, n1269, n1268, n1267, n1272, n1271, n1270, n1276, n1277, n1274, n1275, n1273, n1280, n1279, n1278, n1283, n1282, n1281, n1285, n1286, n1284, n1289, n1288, n1287, n1292, n1291, n1290, n1295, n1296, n1294, n1293, n1299, n1298, n1297, n1301, n1302, n1300, n1305, n1304, n1303, n1308, n1307, n1306, n1311, n1312, n1310, n1309, n1315, n1314, n1313, n1318, n1317, n1316, n1320, n1321, n1319, n1324, n1323, n1322, n1327, n1326, n1325, n1330, n1331, n1329, n1328, n1334, n1333, n1332, n1336, n1337, n1335, n1340, n1339, n1338, n1343, n1342, n1341, n1346, n1347, n1345, n1344, n1350, n1349, n1348, n1353, n1352, n1351, n1355, n1356, n1354, n1359, n1358, n1357, n1362, n1361, n1360, n1365, n1366, n1364, n1363, n1369, n1368, n1367, n1371, n1372, n1370, n1375, n1374, n1373, n1378, n1377, n1376, n1381, n1382, n1380, n1379, n1385, n1384, n1383, n1388, n1387, n1386, n1390, n1391, n1389, n1394, n1393, n1392, n1397, n1396, n1395, n1400, n1401, n1399, n1398, n1404, n1403, n1402, n1406, n1407, n1405, n1408, n1411, n1415, n1416, n1414, n1419, n1420, n1418, n1417, n1422, n1423, n1421, n1425, n1426, n1424, n1428, n1429, n1427, n1431, n1432, n1430, n1434, n1435, n1433, n1437, n1438, n1436, n1440, n1441, n1439, n1443, n1444, n1442, n1446, n1447, n1445, n1449, n1450, n1448, n1452, n1453, n1451, n1455, n1456, n1454, n1458, n1459, n1457, n1461, n1462, n1460, n1464, n1465, n1463, n1467, n1468, n1466, n1470, n1471, n1469, n1475, n1473, n1474, n1472, n1478, n1477, n1476, n1481, n1480, n1479, n1482, n1487, n1490, n1494, n1498, n1504, n1503, n1502, n1505, n1508, n1511, n1514, n1517, n1522, n1520, n1523, n1526, n1525, n1524, n1528, n1527, n1530, n1529, n1532, n1533, n1531, n1536, n1535, n1534, n1539, n1538, n1537, n1541, n1540, n1543, n1544, n1542, n1546, n1545, n1548, n1547, n1550, n1549, n1552, n1553, n1551, n1555, n1554, n1557, n1556, n1559, n1558, n1561, n1562, n1560, n1564, n1563, n1567, n1566, n1565, n1569, n1568, n1571, n1570, n1573, n1574, n1572, n1576, n1575, n1578, n1577, n1580, n1579, n1582, n1583, n1581, n1585, n1584, n1587, n1586, n1589, n1588, n1591, n1592, n1590, n1594, n1593, n1596, n1595, n1598, n1597, n1600, n1601, n1599, n1603, n1602, n1607, n1606, n1605, n1609, n1608, n1611, n1610, n1613, n1614, n1612, n1616, n1615, n1618, n1617, n1620, n1619, n1622, n1623, n1621, n1625, n1624, n1627, n1626, n1629, n1628, n1631, n1632, n1630, n1634, n1633, n1636, n1635, n1638, n1637, n1640, n1641, n1639, n1645, n1646, n1644, n1642, n1647, n1651, n1650, n1649, n1655, n1653, n1654, n1652, n1657, n1658, n1660, n1662, n1663, n1661, n1665, n1667, n1668, n1670, n1671, n1669, n1672, n1673, n1674, n1676, n1675, n1677, n1678, n1679, n1681, n1680, n1682, n1683, n1684, n1686, n1685, n1687, n1688, n1689, n1690, n1693, n1694, n1692, n1691, n1695, n1696, n1697, n1698, n1700, n1701, n1699, n1702, n1703, n1704, n1705, n1707, n1708, n1706, n1709, n1710, n1711, n1712, n1714, n1715, n1713, n1716, n1721, n1719, n1718, n1722, n1726, n1725, n1724, n1727, n1731, n1730, n1729, n1733, n1732, n1734, n1738, n1737, n1736, n1739, n1743, n1742, n1741, n1744, n1748, n1747, n1746, n1750, n1749, n1751, n1755, n1754, n1753, n1756, n1760, n1759, n1758, n1761, n1765, n1764, n1763, n1767, n1766, n1768, n1772, n1771, n1770, n1773, n1777, n1776, n1775, n1778, n1782, n1781, n1780, n1784, n1783, n1785, n1789, n1788, n1787, n1790, n1794, n1793, n1792, n1795, n1797, n1801, n1800, n1799, n1803, n1804, n1802, n1805, n1809, n1808, n1807, n1810, n1814, n1813, n1812, n1815, n1817, n1821, n1820, n1819, n1823, n1824, n1822, n1825, n1829, n1828, n1827, n1830, n1834, n1833, n1832, n1835, n1837, n1841, n1840, n1839, n1843, n1844, n1842, n1845, n1849, n1848, n1847, n1850, n1854, n1853, n1852, n1855, n1857, n1861, n1860, n1859, n1863, n1864, n1862, n1867, n1868, n1866, n1865, n1870, n1869, n1872, n1871, n1874, n1873, n1876, n1875, n1878, n1877, n1880, n1879, n1882, n1881, n1885, n1886, n1884, n1883, n1888, n1887, n1891, n1890, n1889, n1893, n1892, n1895, n1894, n1898, n1897, n1896, n1900, n1899, n1902, n1903, n1901, n1905, n1904, n1907, n1906, n1909, n1908, n1911, n1910, n1913, n1912, n1915, n1914, n1917, n1916, n1919, n1918, n1921, n1922, n1920, n1924, n1923, n1927, n1926, n1925, n1929, n1928, n1931, n1930, n1934, n1933, n1932, n1936, n1935, n1938, n1939, n1937, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1951, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1961, n1965, n1963, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1976, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1986, n1988, n1994, n1993, n1991, n1992, n1990, n1995, n1997, n1996, n1998, n1999, n2000, n2001, n2002, n2003, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2017, n2016, n2025, n2024, n2028, n2026, n2031, n2029, n2032, n2036, n2042, n2040, n2045, n2043, n2046, n2050, n2049, n2048, n2052, n2055, n2053, n2056, n2058, n2059, n2060, n2061, n2057, n2062, n2063, n2065, n2064, n2066, n2069, n2068, n2073, n2071, n2070, n2074, n2079, n2078, n2076, n2081, n2082, n2083, n2084, n2080, n2086, n2087, n2085, n2088, n2091, n2094, n2093, n2092, n2096, n2095, n2098, n2099, n2097, n2100, n2101, n2103, n2105, n2104, n2106, n2108, n2107, n2109, n2111, n2113, n2112, n2116, n2115, n2114, n2118, n2117, n2119, n2120, n2122, n2124, n2123, n2126, n2125, n2127, n2128, n2130, n2132, n2131, n2134, n2133, n2135, n2137, n2139, n2138, n2142, n2141, n2140, n2143, n2145, n2147, n2149, n2148, n2150, n2151, n2153, n2155, n2154, n2156, n2158, n2160, n2159, n2163, n2162, n2161, n2164, n2165, n2167, n2169, n2168, n2170, n2171, n2173, n2175, n2174, n2176, n2178, n2180, n2179, n2183, n2182, n2181, n2184, n2185, n2187, n2189, n2188, n2190, n2191, n2193, n2195, n2194, n2197, n2196, n2199, n2198, n2200, n2202, n2204, n2203, n2206, n2205, n2207, n2208, n2210, n2212, n2211, n2215, n2216, n2214, n2213, n2217, n2219, n2221, n2220, n2222, n2224, n2226, n2225, n2228, n2227, n2229, n2230, n2232, n2234, n2233, n2236, n2235, n2237, n2238, n2240, n2242, n2241, n2245, n2246, n2244, n2243, n2248, n2247, n2249, n2251, n2250, n2253, n2252, n2254, n2256, n2255, n2257, n2259, n2261, n2263, n2262, n2264, n2265, n2267, n2269, n2268, n2272, n2273, n2271, n2270, n2275, n2274, n2276, n2278, n2277, n2280, n2279, n2281, n2283, n2282, n2284, n2285, n2287, n2289, n2288, n2290, n2291, n2293, n2295, n2294, n2298, n2299, n2297, n2296, n2302, n2300, n2303, n2306, n2305, n2304, n2307, n2310, n2309, n2308, n2313, n2312, n2311, n2316, n2315, n2314, n2317, n2323, n2321, n2326, n2325, n2324, n2328, n2327, n2331, n2332, n2330, n2329, n2333, n2335, n2334, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2351, n2352, n2350, n2353, n2356, n2360, n2361, n2362, n2359, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2378, n2379, n2377, n2380, n2383, n2386, n2391, n2392, n2390, n2393, n2394, n2396, n2397, n2401, n2404, n2407, n2412, n2410, n2411, n2409, n2415, n2414, n2413, n2417, n2416, n2419, n2420, n2418, n2423, n2422, n2421, n2426, n2425, n2424, n2428, n2427, n2430, n2431, n2429, n2434, n2433, n2432, n2437, n2436, n2435, n2439, n2438, n2441, n2442, n2440, n2445, n2444, n2443, n2448, n2447, n2446, n2450, n2449, n2452, n2453, n2451, n2456, n2454, n2458, n2461, n2462, n2464, n2467, n2466, n2465, n2469, n2468, n2471, n2470, n2473, n2474, n2472, n2476, n2475, n2478, n2477, n2480, n2479, n2482, n2483, n2481, n2485, n2484, n2487, n2486, n2489, n2488, n2491, n2492, n2490, n2494, n2493, n2496, n2495, n2498, n2497, n2500, n2501, n2499, n2502, n2504, n2506, n2508, n2509, n2512, n2511, n2510, n2513, n2514, n2515, n2518, n2517, n2516, n2519, n2520, n2521, n2524, n2523, n2522, n2525, n2526, n2527, n2530, n2529, n2528, n2531, n2532, n2533, n2534, n2537, n2538, n2536, n2535, n2539, n2540, n2541, n2542, n2545, n2546, n2544, n2543, n2547, n2548, n2549, n2550, n2553, n2554, n2552, n2551, n2555, n2556, n2557, n2558, n2561, n2562, n2560, n2559, n2564, n2563, n2566, n2565, n2568, n2567, n2570, n2571, n2569, n2573, n2574, n2572, n2576, n2577, n2575, n2580, n2579, n2578, n2582, n2581, n2584, n2583, n2587, n2588, n2586, n2585, n2590, n2589, n2592, n2591, n2594, n2595, n2593, n2597, n2596, n2599, n2598, n2602, n2603, n2601, n2600, n2605, n2604, n2607, n2608, n2606, n2610, n2609, n2612, n2611, n2615, n2616, n2614, n2613, n2618, n2617, n2620, n2619, n2622, n2623, n2621, n2625, n2624, n2627, n2626, n2630, n2631, n2629, n2628, n2633, n2632, n2635, n2636, n2634, n2638, n2637, n2640, n2639, n2643, n2644, n2642, n2641, n2646, n2645, n2648, n2647, n2650, n2651, n2649, n2653, n2652, n2655, n2654, n2658, n2659, n2657, n2656, n2661, n2660, n2663, n2664, n2662, n2666, n2665, n2668, n2667, n2671, n2672, n2670, n2669, n2674, n2673, n2676, n2675, n2678, n2679, n2677, n2681, n2680, n2683, n2682, n2686, n2687, n2685, n2684, n2689, n2688, n2691, n2692, n2690, n2693, n2696, n2700, n2701, n2699, n2703, n2704, n2702, n2706, n2707, n2705, n2709, n2710, n2708, n2712, n2713, n2711, n2715, n2716, n2714, n2718, n2719, n2717, n2721, n2722, n2720, n2724, n2725, n2723, n2727, n2728, n2726, n2730, n2731, n2729, n2733, n2734, n2732, n2736, n2737, n2735, n2739, n2740, n2738, n2742, n2743, n2741, n2745, n2746, n2744, n2748, n2749, n2747, n2751, n2752, n2750, n2754, n2753, n2757, n2756, n2755, n2760, n2759, n2758, n2763, n2762, n2761, n2764, n2767, n2770, n2773, n2776, n2781, n2780, n2782, n2785, n2788, n2791, n2794, n2799, n2797, n2800, n2802, n2801, n2804, n2803, n2806, n2805, n2808, n2809, n2807, n2811, n2810, n2813, n2812, n2815, n2814, n2817, n2818, n2816, n2820, n2819, n2822, n2821, n2824, n2823, n2826, n2827, n2825, n2830, n2829, n2828, n2833, n2832, n2831, n2835, n2834, n2837, n2838, n2836, n2839, n2841, n2840, n2843, n2842, n2845, n2844, n2847, n2848, n2846, n2850, n2849, n2852, n2851, n2854, n2853, n2856, n2857, n2855, n2859, n2858, n2861, n2860, n2863, n2862, n2865, n2866, n2864, n2868, n2867, n2870, n2869, n2872, n2871, n2874, n2875, n2873, n2876, n2878, n2877, n2880, n2879, n2882, n2881, n2884, n2885, n2883, n2887, n2886, n2889, n2888, n2891, n2890, n2893, n2894, n2892, n2896, n2895, n2898, n2897, n2900, n2899, n2902, n2903, n2901, n2905, n2904, n2907, n2906, n2909, n2908, n2911, n2912, n2910, n2913, n2916, n2920, n2923, n2926, n2931, n2932, n2936, n2937, n2939, n2947, n2946, n2950, n2952, n2953, n2954, n2955, n2959, n2958, n2961, n2962, n2960, n2965, n2964, n2963, n2967, n2966, n2968, n2971, n2970, n2972, n2973, n2975, n2976, n2974, n2979, n2978, n2977, n2980, n2981, n2986, n2985, n2989, n2990, n2988, n2992, n2991, n2993, n2995, n2996, n2994, n2997, n3001, n2999, n2998, n3003, n3002, n3005, n3004, n3006, n3007, n3009, n3008, n3011, n3010, n3012, n3013, n3014, n3015, n3018, n3017, n3021, n3020, n3019, n3023, n3022, n3025, n3024, n3026, n3028, n3027, n3029, n3031, n3030, n3033, n3032, n3034, n3035, n3039, n3040, n3038, n3043, n3042, n3044, n3046, n3045, n3048, n3047, n3049, n3051, n3050, n3053, n3052, n3055, n3054, n3057, n3056, n3058, n3060, n3059, n3062, n3063, n3061, n3065, n3064, n3068, n3072, n3071, n3074, n3073, n3075, n3077, n3076, n3078, n3081, n3080, n3083, n3082, n3084, n3086, n3085, n3087, n3089, n3091, n3090, n3092, n3094, n3093, n3096, n3097, n3095, n3098, n3100, n3099, n3101, n3103, n3102, n3105, n3106, n3104, n3107, n3109, n3113, n3111, n3114, n3116, n3120, n3119, n3122, n3121, n3125, n3124, n3127, n3126, n3129, n3130, n3128, n3132, n3131, n3134, n3133, n3136, n3135, n3138, n3137, n3140, n3139, n3141, n3143, n3142, n3144, n3145, n3147, n3146, n3149, n3148, n3151, n3150, n3153, n3152, n3154, n3156, n3155, n3158, n3157, n3160, n3159, n3161, n3162, n3163, n3164, n3166, n3165, n3167, n3168, n3169, n3170, n3171, n3173, n3172, n3174, n3175, n3176, n3177, n3178, n3180, n3179, n3182, n3183, n3181, n3185, n3184, n3186, n3188, n3189, n3187, n3191, n3190, n3192, n3194, n3193, n3196, n3195, n3198, n3197, n3199, n3201, n3200, n3203, n3202, n3205, n3204, n3206, n3208, n3209, n3207, n3211, n3210, n3213, n3212, n3214, n3216, n3215, n3218, n3217, n3219, n3221, n3220, n3223, n3222, n3225, n3224, n3226, n3228, n3227, n3230, n3229, n3232, n3231, n3233, n3235, n3236, n3234, n3238, n3237, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3247, n3248, n3246, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3258, n3259, n3257, n3261, n3260, n3262, n3265, n3268, n3270, n3271, n3273, n3275, n3279, n3278, n3277, n3281, n3280, n3282, n3283, n3285, n3284, n3286, n3287, n3288, n3290, n3289, n3291, n3292, n3293, n3295, n3294, n3296, n3297, n3298, n3300, n3299, n3301, n3302, n3303, n3304, n3306, n3307, n3305, n3308, n3309, n3310, n3311, n3313, n3314, n3312, n3315, n3316, n3317, n3318, n3320, n3321, n3319, n3322, n3323, n3324, n3325, n3327, n3328, n3326, n3329, n3330, n3332, n3334, n3335, n3337, n3339, n3342, n3341, n3344, n3343, n3346, n3345, n3348, n3347, n3350, n3349, n3353, n3352, n3351, n3355, n3354, n3357, n3356, n3359, n3358, n3361, n3360, n3363, n3362, n3365, n3364, n3367, n3366, n3369, n3368, n3371, n3370, n3373, n3372, n3375, n3374, n3377, n3376, n3379, n3378, n3381, n3380, n3383, n3382, n3385, n3386, n3384, n3388, n3387, n3390, n3389, n3392, n3391, n3394, n3393, n3396, n3397, n3395, n3399, n3398, n3401, n3400, n3403, n3402, n3405, n3404, n3407, n3408, n3406, n3410, n3409, n3412, n3411, n3414, n3413, n3416, n3415, n3418, n3419, n3417, n3421, n3420, n3424, n3425, n3423, n3428, n3427, n3426, n3431, n3430, n3429, n3432, n3433, n3438, n3437, n3439, n3440, n3442, n3441, n3444, n3446, n3448, n3450, n3452, n3451, n3453, n3455, n3454, n3456, n3457, n3460, n3459, n3461, n3462, n3463, n3465, n3467, n3469, n3472, n3471, n3477, n3476, n3474, n3480, n3478, n3482, n3486, n3487, n3489, n3490, n3488, n3492, n3495, n3496, n3494, n3493, n3500, n3501, n3498, n3499, n3497, n3503, n3502, n3504, n3510, n3508, n3507, n3511, n3514, n3512, n3516, n3515, n3518, n3519, n3517, n3520, n3526, n3524, n3525, n3523, n3528, n3529, n3527, n3530, n3531, n3533, n3535, n3534, n3538, n3540, n3539, n3542, n3543, n3545, n3544, n3548, n3550, n3549, n3554, n3553, n3555, n3556, n3557, n3558, n3560, n3559, n3563, n3561, n3564, n3568, n3566, n3567, n3565, n3569, n3573, n3572, n3571, n3574, n3577, n3576, n3575, n3580, n3579, n3578, n3583, n3582, n3581, n3585, n3584, n3586, n3587, n3589, n3588, n3592, n3590, n3591, n3593, n3595, n3594, n3596, n3597, N_N13958, n3598, n3603, n3601, n3604, n3608, n3610, n3612, n3613, n3614, n3611, n3615, n3616, n3618, n3617, Nv437, n3620, Nv43, n3621, Nv14, n3622, n3623, n3624, N_N13959, n3626, n3627, n3628, n3629, n3631, n3632, n3630, n3634, n3635, n3633, n3638, n3639, n3640, n3641, n3643, n3646, n3647, n3645, n3649, n3650, n3653, n3655, n3659, n3657, n3662, n3660, n3663, n3665, n3666, n3667, n3668, n3671, n3670, n3669, n3672, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3685, n3684, n3687, n3686, n3691, n3690, n3692, n3695, n3696, n3697, n3698, n3699, n3701, n3700, n3702, n3703, n3705, n3706, n3708, n3712, n3713, n3716, n3718, n3719, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3731, n3733, n3734, n3732, n3735, n3736, n3737, n3738, n3739, n3740, n3742, n3747, n3748, n3746, n3749, n3750, n3751, n3754, n3757, n3758, n3756, n3760, n3761, n3759, n3763, n3767, n3768, n3766, n3770, n3771, n3769, n3774, n3775, n3776, n3777, n3778, n3779, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3842, n3841, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3851, n3852, n3854, n3855, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3869, n3870, n3871, n3874, n3875, n3876, n3877, n3879, n3880, n3881, n3882, Nv8909, n3886, n3887, n3888, n3890, n3891, n3893, n3894, n3898, n3899, n3900, n3901, n3905, n3908, n3906, n3910, n3912, n3914, n3916, n3918, n3920, n3922, n3923, n3926, n3925, n3928, n3930, n3932, n3931, n3934, n3936, n3938, n3939, n3940, n3941, n3937, n3943, n3944, n3945, n3946, n3942, n3948, n3949, n3950, n3951, n3953, n3952, n3955, Nv10316, n3957, n3958, n3956, n3959, Nv10135, n3960, Nv10099, n3962, n3961, n3963, Nv10091, n3964, Nv10082, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3984, n3983, n3985, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3997, n3996, n3998, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4053, n4055, n4057, n4056, n4059, n4058, n4061, n4062, n4060, n4064, n4063, n4066, n4067, n4065, n4068, n4069, n4071, n4070, n4073, n4072, n4075, n4076, n4074, n4078, n4077, n4080, n4081, n4079, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4093, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4117, n4116, n4120, n4119, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4141, n4140, n4142, n4143, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4161, n4160, n4162, n4163, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4177, n4176, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4202, n4203, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4221, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4233, n4236, n4238, n4239, n4240, n4241, n4244, n4245, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4269, n4270, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4281, n4283, n4285, n4287, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4299, n4300, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4311, n4313, n4315, n4317, n4319, n4320, n4321, n4322, n4323, n4325, n4324, n4326, n4328, n4330, n4331, n4332, n4333, n4334, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4361, n4363, n4365, n4364, n4366, n4368, n4367, n4369, n4371, n4370, n4372, n4373, n4375, n4374, n4376, n4378, n4377, n4379, n4381, n4380, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4391, n4394, n4395, n4396, n4398, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4414, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4442, n4441, n4443, n4444, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4462, n4461, n4463, n4464, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4484, n4483, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4500, n4499, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4516, n4517, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4536, n4539, n4540, n4541, n4542, n4544, n4543, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4560, n4559, n4561, n4562, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4574, n4573, n4575, n4577, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4599, n4598, n4600, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4612, n4613, n4614, n4615, n4616, n4617, n4619, n4620, n4621, n4622, n4623, n4625, n4627, n4628, n4629, n4631, n4632, n4633, n4635, n4636, n4637, n4638, n4639, n4641, n4643, n4644, n4645, n4647, n4648, n4649, n4650, n4652, n4654, n4657, n4658, n4659, n4665, n4666, n4667, n4669, n4670, n4671, n4672, n4673, n4675, n4676, n4677, n4678, n4682, n4686, n4685, n4688, n4687, n4689, n4691, n4692, n4693, n4696, n4699, n4698, n4701, n4702, n4703, n4704, n4705, n4706, n4708, n4709, n4711, n4712, n4713, n4714, n4716, n4717, n4718, n4719, n4720, n4722, n4724, n4730, n4733, n4735, n4737, n4738, n4740, n4743, n4747, n4746, n4749, n4748, n4750, n4752, n4753, n4754, n4755, n4756, n4759, n4760, n4761, n4763, n4764, n4766, n4767, n4769, n4770, n4772, n4773, n4775, n4776, n4777, n4779, n4780, n4783, n4784, n4785, n4786, n4787, n4790, n4791, n4792, n4797, n4798, n4799, n4800, n4801, n4803, n4805, n4808, n4810, n4811, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4822, n4823, n4825, n4827, n4832, n4833, n4835, n4836;

reg Ni48, Ni47, Ni46, Ni45, Ni44, Ni43, Ni42, Ni41, Ni40, Ni39, Ni38, Ni37, Ni36, Ni35, Ni34, Ni33, Ni32, Ni31, Ni30, n18, Ni14, Ni13, Ni12, Ni11, Ni10, Ni9, Ni8, Ni7, Ni6, Ni5, Ni4, Ni3, Ni2;

always  @(posedge PCLK)
	Ni48<=Nv2;

 always  @(posedge PCLK)
	Ni47<=Nv14;

 always  @(posedge PCLK)
	Ni46<=Nv31;

 always  @(posedge PCLK)
	Ni45<=Nv43;

 always  @(posedge PCLK)
	Ni44<=Nv59;

 always  @(posedge PCLK)
	Ni43<=N_N13960;

 always  @(posedge PCLK)
	Ni42<=N_N13959;

 always  @(posedge PCLK)
	Ni41<=Nv243;

 always  @(posedge PCLK)
	Ni40<=Nv294;

 always  @(posedge PCLK)
	Ni39<=Nv345;

 always  @(posedge PCLK)
	Ni38<=Nv349;

 always  @(posedge PCLK)
	Ni37<=Nv437;

 always  @(posedge PCLK)
	Ni36<=Nv499;

 always  @(posedge PCLK)
	Ni35<=Nv550;

 always  @(posedge PCLK)
	Ni34<=Nv601;

 always  @(posedge PCLK)
	Ni33<=Nv2153;

 always  @(posedge PCLK)
	Ni32<=Nv3888;

 always  @(posedge PCLK)
	Ni31<=Nv6425;

 always  @(posedge PCLK)
	Ni30<=Nv6437;

 always  @(posedge PCLK)
	n18<=Nv8909;

 always  @(posedge PCLK)
	Ni14<=Nv10056;

 always  @(posedge PCLK)
	Ni13<=Nv10068;

 always  @(posedge PCLK)
	Ni12<=Nv10082;

 always  @(posedge PCLK)
	Ni11<=Nv10091;

 always  @(posedge PCLK)
	Ni10<=Nv10099;

 always  @(posedge PCLK)
	Ni9<=Nv10112;

 always  @(posedge PCLK)
	Ni8<=Nv10126;

 always  @(posedge PCLK)
	Ni7<=Nv10135;

 always  @(posedge PCLK)
	Ni6<=Nv10143;

 always  @(posedge PCLK)
	Ni5<=Nv10247;

 always  @(posedge PCLK)
	Ni4<=Nv10316;

 always  @(posedge PCLK)
	Ni3<=P__cmxcl_0;

 always  @(posedge PCLK)
	Ni2<=N_N13958;

 assign P__cmxir_1 = ( n157  &  (~ n3113)  &  (~ n3540) ) ;
 assign P__cmxir_0 = ( (~ n138)  &  (~ n3476) ) ;
 assign P__cmxig_1 = ( (~ n157) ) ;
 assign P__cmxig_0 = ( (~ n3837) ) ;
 assign P__cmxcl_1 = ( (~ n3540) ) ;
 assign P__cmxcl_0 = ( (~ n3540) ) ;
 assign P__cmx1ad_35 =((~ Pi416) & Pi416);
 assign P__cmx1ad_34 =((~ Pi416) & Pi416);
 assign P__cmx1ad_33 =((~ Pi416) & Pi416);
 assign P__cmx1ad_32 =((~ Pi416) & Pi416);
 assign P__cmx1ad_31 = ( Pi255  &  (~ n3880) ) ;
 assign P__cmx1ad_30 = ( Pi254  &  (~ n3880) ) ;
 assign P__cmx1ad_29 = ( Pi253  &  (~ n3880) ) ;
 assign P__cmx1ad_28 = ( Pi252  &  (~ n3880) ) ;
 assign P__cmx1ad_27 = ( Pi251  &  (~ n3880) ) ;
 assign P__cmx1ad_26 = ( Pi250  &  (~ n3880) ) ;
 assign P__cmx1ad_25 = ( Pi249  &  (~ n3880) ) ;
 assign P__cmx1ad_24 = ( Pi248  &  (~ n3880) ) ;
 assign P__cmx1ad_23 = ( Pi247  &  (~ n3880) ) ;
 assign P__cmx1ad_22 = ( Pi246  &  (~ n3880) ) ;
 assign P__cmx1ad_21 = ( Pi245  &  (~ n3880) ) ;
 assign P__cmx1ad_20 = ( Pi244  &  (~ n3880) ) ;
 assign P__cmx1ad_19 = ( Pi243  &  (~ n3880) ) ;
 assign P__cmx1ad_18 = ( Pi242  &  (~ n3880) ) ;
 assign P__cmx1ad_17 = ( Pi241  &  (~ n3880) ) ;
 assign P__cmx1ad_16 = ( Pi240  &  (~ n3880) ) ;
 assign P__cmx1ad_15 = ( Pi27  &  Pi26  &  (~ n3880) ) ;
 assign P__cmx1ad_14 = ( (~ n3966) ) ;
 assign P__cmx1ad_13 = ( n161  &  (~ n3880) ) ;
 assign P__cmx1ad_12 = ( (~ n4813) ) ;
 assign P__cmx1ad_11 =((~ Pi416) & Pi416);
 assign P__cmx1ad_10 =((~ Pi416) & Pi416);
 assign P__cmx1ad_9 = ( (~ n3880) ) ;
 assign P__cmx1ad_8 =((~ Pi416) & Pi416);
 assign P__cmx1ad_7 = ( Pi239  &  (~ n3880) ) ;
 assign P__cmx1ad_6 = ( Pi238  &  (~ n3880) ) ;
 assign P__cmx1ad_5 = ( Pi237  &  (~ n3880) ) ;
 assign P__cmx1ad_4 = ( Pi236  &  (~ n3880) ) ;
 assign P__cmx1ad_3 = ( Pi235  &  (~ n3880) ) ;
 assign P__cmx1ad_2 = ( Pi234  &  (~ n3880) ) ;
 assign P__cmx1ad_1 = ( Pi233  &  (~ n3880) ) ;
 assign P__cmx1ad_0 = ( Pi232  &  (~ n3880) ) ;
 assign P__cmx0ad_35 =((~ Pi416) & Pi416);
 assign P__cmx0ad_34 =((~ Pi416) & Pi416);
 assign P__cmx0ad_33 =((~ Pi416) & Pi416);
 assign P__cmx0ad_32 =((~ Pi416) & Pi416);
 assign P__cmx0ad_31 = ( Pi72  &  (~ n3881) ) ;
 assign P__cmx0ad_30 = ( Pi71  &  (~ n3881) ) ;
 assign P__cmx0ad_29 = ( Pi70  &  (~ n3881) ) ;
 assign P__cmx0ad_28 = ( Pi69  &  (~ n3881) ) ;
 assign P__cmx0ad_27 = ( Pi68  &  (~ n3881) ) ;
 assign P__cmx0ad_26 = ( Pi67  &  (~ n3881) ) ;
 assign P__cmx0ad_25 = ( Pi66  &  (~ n3881) ) ;
 assign P__cmx0ad_24 = ( Pi65  &  (~ n3881) ) ;
 assign P__cmx0ad_23 = ( Pi64  &  (~ n3881) ) ;
 assign P__cmx0ad_22 = ( Pi63  &  (~ n3881) ) ;
 assign P__cmx0ad_21 = ( Pi62  &  (~ n3881) ) ;
 assign P__cmx0ad_20 = ( Pi61  &  (~ n3881) ) ;
 assign P__cmx0ad_19 = ( Pi60  &  (~ n3881) ) ;
 assign P__cmx0ad_18 = ( Pi59  &  (~ n3881) ) ;
 assign P__cmx0ad_17 = ( Pi58  &  (~ n3881) ) ;
 assign P__cmx0ad_16 = ( Pi57  &  (~ n3881) ) ;
 assign P__cmx0ad_15 = ( Pi24  &  Pi23  &  (~ n3881) ) ;
 assign P__cmx0ad_14 = ( (~ n3967) ) ;
 assign P__cmx0ad_13 = ( n160  &  (~ n3881) ) ;
 assign P__cmx0ad_12 = ( (~ n4815) ) ;
 assign P__cmx0ad_11 =((~ Pi416) & Pi416);
 assign P__cmx0ad_10 =((~ Pi416) & Pi416);
 assign P__cmx0ad_9 = ( (~ n3881) ) ;
 assign P__cmx0ad_8 =((~ Pi416) & Pi416);
 assign P__cmx0ad_7 = ( Pi56  &  (~ n3881) ) ;
 assign P__cmx0ad_6 = ( Pi55  &  (~ n3881) ) ;
 assign P__cmx0ad_5 = ( Pi54  &  (~ n3881) ) ;
 assign P__cmx0ad_4 = ( Pi53  &  (~ n3881) ) ;
 assign P__cmx0ad_3 = ( Pi52  &  (~ n3881) ) ;
 assign P__cmx0ad_2 = ( Pi51  &  (~ n3881) ) ;
 assign P__cmx0ad_1 = ( Pi50  &  (~ n3881) ) ;
 assign P__cmx0ad_0 = ( Pi49  &  (~ n3881) ) ;
 assign P__cmnxcp_1 = ( (~ n159) ) ;
 assign P__cmnxcp_0 = ( (~ n158) ) ;
 assign P__cmndst1p0 = ( n153  &  (~ n3593) ) ;
 assign P__cmndst0p0 = ( n150  &  (~ n3879) ) ;
 assign n19 = ( (~ n3478)  &  (~ Ni48) ) | ( (~ Pi22)  &  (~ n3478)  &  n3482 ) ;
 assign Nv2 = ( (~ n19) ) ;
 assign n20 = ( Pi20  &  (~ n299)  &  n2947 ) | ( (~ n299)  &  n2947  &  n2946 ) ;
 assign n21 = ( Pi21  &  Ni46 ) | ( (~ Ni32)  &  (~ n2065)  &  Ni46 ) ;
 assign Nv31 = ( n20 ) | ( n21 ) ;
 assign n22 = ( (~ Ni44)  &  (~ n3687) ) | ( (~ n3592)  &  (~ n3687) ) ;
 assign Nv59 = ( (~ n22) ) ;
 assign n25 = ( Ni44  &  Ni39 ) | ( (~ Ni44)  &  (~ Ni39) ) ;
 assign n24 = ( n25  &  Ni38 ) ;
 assign n23 = ( n25  &  Ni32  &  Ni37 ) | ( n25  &  Ni32  &  n24 ) ;
 assign n26 = ( n2040  &  n2954 ) | ( n2954  &  (~ Ni41) ) ;
 assign Nv243 = ( (~ n26) ) ;
 assign n27 = ( n2040  &  n2952 ) | ( n2952  &  (~ Ni40) ) ;
 assign Nv294 = ( (~ n27) ) ;
 assign n28 = ( n32  &  n2028 ) | ( n2028  &  (~ Ni39) ) ;
 assign Nv345 = ( (~ n28) ) ;
 assign n29 = ( (~ n694)  &  (~ n2937)  &  (~ n3735) ) | ( (~ n2025)  &  (~ n2937)  &  (~ n3735) ) ;
 assign n30 = ( n190  &  (~ n796)  &  (~ n2937) ) | ( (~ n400)  &  (~ n796)  &  (~ n2937) ) ;
 assign n31 = ( Pi15  &  (~ n107)  &  (~ n3879) ) ;
 assign n32 = ( (~ Ni32)  &  n2055 ) ;
 assign n34 = ( (~ n2937)  &  n2939  &  (~ n3879) ) ;
 assign Nv349 = ( n29 ) | ( n30 ) | ( n31 ) | ( n32 ) | ( n34 ) | ( (~ n4835) ) ;
 assign n35 = ( (~ Ni36)  &  (~ n2048)  &  n2052 ) | ( n2040  &  (~ n2048)  &  n2052 ) ;
 assign Nv499 = ( (~ n35) ) ;
 assign n36 = ( (~ Ni35)  &  (~ n2036)  &  n2042 ) | ( (~ n2036)  &  n2042  &  n2040 ) ;
 assign Nv550 = ( (~ n36) ) ;
 assign n37 = ( (~ Ni34)  &  (~ n2016)  &  (~ n3657) ) | ( (~ n2016)  &  (~ n3540)  &  (~ n3657) ) ;
 assign Nv601 = ( (~ n37) ) ;
 assign n38 = ( (~ Ni44)  &  (~ Ni42) ) | ( (~ n104)  &  (~ Ni42) ) ;
 assign n42 = ( Ni44  &  (~ Ni42) ) | ( (~ n104)  &  (~ Ni42) ) ;
 assign n44 = ( (~ Ni47)  &  (~ Ni45) ) ;
 assign n45 = ( (~ Ni42) ) | ( Ni43 ) ;
 assign n43 = ( n44  &  n45 ) ;
 assign n46 = ( n3477  &  n3476 ) | ( (~ n3471)  &  n3477  &  n3474 ) ;
 assign Nv2153 = ( (~ n46) ) ;
 assign n47 = ( (~ n1653)  &  (~ n2932)  &  n2936 ) | ( (~ n2932)  &  n2936  &  (~ n4391) ) ;
 assign Nv3888 = ( (~ n47) ) ;
 assign n48 = ( (~ n43)  &  n1660  &  (~ n3540) ) | ( (~ n200)  &  n1660  &  (~ n3540) ) ;
 assign n49 = ( (~ Ni32)  &  (~ Ni30)  &  n1866  &  (~ n3540) ) ;
 assign Nv6425 = ( n48 ) | ( n49 ) | ( Ni31 ) ;
 assign n50 = ( (~ Ni30)  &  n1657  &  n1658 ) | ( n1657  &  n1658  &  (~ n3540) ) ;
 assign Nv6437 = ( (~ n50) ) ;
 assign n55 = ( n878  &  n879  &  n52 ) | ( n878  &  n879  &  n877 ) ;
 assign n52 = ( n4823  &  n79 ) ;
 assign n53 = ( (~ n200) ) | ( (~ Ni36) ) ;
 assign n51 = ( n55  &  n52  &  (~ n1063) ) | ( n55  &  n53  &  (~ n1063) ) ;
 assign n60 = ( n878  &  n879  &  n59 ) | ( n878  &  n879  &  n882 ) ;
 assign n59 = ( n4825  &  n79 ) ;
 assign n58 = ( n53  &  n60  &  (~ n1063) ) | ( n60  &  n59  &  (~ n1063) ) ;
 assign n64 = ( n62  &  n390 ) | ( n390  &  (~ Ni38) ) ;
 assign n65 = ( n111  &  (~ n1063) ) | ( (~ Ni35)  &  (~ n1063) ) ;
 assign n62 = ( n52  &  n79 ) | ( n79  &  (~ Ni40) ) ;
 assign n63 = ( Ni37 ) | ( (~ Ni36) ) ;
 assign n61 = ( n64  &  n65  &  n62 ) | ( n64  &  n65  &  n63 ) ;
 assign n68 = ( n67  &  n390 ) | ( n390  &  (~ Ni38) ) ;
 assign n69 = ( n114  &  (~ n1063) ) | ( (~ Ni35)  &  (~ n1063) ) ;
 assign n67 = ( n59  &  n79 ) | ( n79  &  (~ Ni40) ) ;
 assign n66 = ( n68  &  n69  &  n67 ) | ( n68  &  n69  &  n63 ) ;
 assign n72 = ( n71  &  n390 ) | ( n390  &  (~ Ni38) ) ;
 assign n73 = ( Ni35  &  (~ n1063) ) | ( n116  &  (~ n1063) ) ;
 assign n71 = ( n79  &  Ni40 ) | ( n79  &  n52 ) ;
 assign n70 = ( n72  &  n73  &  n71 ) | ( n72  &  n73  &  n63 ) ;
 assign n76 = ( n75  &  n390 ) | ( n390  &  (~ Ni38) ) ;
 assign n77 = ( Ni35  &  (~ n1063) ) | ( n118  &  (~ n1063) ) ;
 assign n75 = ( n79  &  Ni40 ) | ( n79  &  n59 ) ;
 assign n74 = ( n76  &  n77  &  n75 ) | ( n76  &  n77  &  n63 ) ;
 assign n80 = ( n79  &  n390 ) | ( n390  &  (~ Ni38) ) ;
 assign n79 = ( n104  &  n835 ) | ( n104  &  (~ Ni41) ) ;
 assign n78 = ( n63  &  n80  &  (~ n1063) ) | ( n80  &  n79  &  (~ n1063) ) ;
 assign n83 = ( n878  &  n879  &  n82 ) | ( n878  &  n879  &  n877 ) ;
 assign n82 = ( n104  &  n4823 ) ;
 assign n81 = ( n53  &  n83  &  (~ n1063) ) | ( n83  &  n82  &  (~ n1063) ) ;
 assign n86 = ( n878  &  n879  &  n85 ) | ( n878  &  n879  &  n882 ) ;
 assign n85 = ( n104  &  n4825 ) ;
 assign n84 = ( n53  &  n86  &  (~ n1063) ) | ( n86  &  n85  &  (~ n1063) ) ;
 assign n89 = ( n88  &  n390 ) | ( n390  &  (~ Ni38) ) ;
 assign n90 = ( (~ Ni35)  &  (~ n1063) ) | ( n122  &  (~ n1063) ) ;
 assign n88 = ( n82  &  n104 ) | ( n104  &  (~ Ni40) ) ;
 assign n87 = ( n89  &  n90  &  n88 ) | ( n89  &  n90  &  n63 ) ;
 assign n93 = ( n92  &  n390 ) | ( n390  &  (~ Ni38) ) ;
 assign n94 = ( (~ Ni35)  &  (~ n1063) ) | ( n124  &  (~ n1063) ) ;
 assign n92 = ( n85  &  n104 ) | ( n104  &  (~ Ni40) ) ;
 assign n91 = ( n93  &  n94  &  n92 ) | ( n93  &  n94  &  n63 ) ;
 assign n97 = ( n96  &  n390 ) | ( n390  &  (~ Ni38) ) ;
 assign n98 = ( Ni35  &  (~ n1063) ) | ( n126  &  (~ n1063) ) ;
 assign n96 = ( n104  &  Ni40 ) | ( n104  &  n82 ) ;
 assign n95 = ( n97  &  n98  &  n96 ) | ( n97  &  n98  &  n63 ) ;
 assign n101 = ( n100  &  n390 ) | ( n390  &  (~ Ni38) ) ;
 assign n102 = ( Ni35  &  (~ n1063) ) | ( n128  &  (~ n1063) ) ;
 assign n100 = ( n104  &  Ni40 ) | ( n104  &  n85 ) ;
 assign n99 = ( n101  &  n102  &  n100 ) | ( n101  &  n102  &  n63 ) ;
 assign n105 = ( n104  &  n390 ) | ( n390  &  (~ Ni38) ) ;
 assign n104 = ( n44  &  (~ Ni43) ) ;
 assign n103 = ( n63  &  n105  &  (~ n1063) ) | ( n105  &  n104  &  (~ n1063) ) ;
 assign n108 = ( n390  &  (~ n1063) ) ;
 assign n107 = ( (~ Ni36) ) | ( (~ Ni38) ) ;
 assign n106 = ( n55  &  n108  &  n52 ) | ( n55  &  n108  &  n107 ) ;
 assign n109 = ( n60  &  n108  &  n59 ) | ( n60  &  n108  &  n107 ) ;
 assign n111 = ( n62 ) | ( n202 ) ;
 assign n110 = ( n64  &  n111  &  (~ n1063) ) | ( n64  &  (~ Ni35)  &  (~ n1063) ) ;
 assign n114 = ( n67 ) | ( n240 ) ;
 assign n113 = ( n68  &  n114  &  (~ n1063) ) | ( n68  &  (~ Ni35)  &  (~ n1063) ) ;
 assign n116 = ( n71 ) | ( n202 ) ;
 assign n115 = ( n72  &  Ni35  &  (~ n1063) ) | ( n72  &  n116  &  (~ n1063) ) ;
 assign n118 = ( n75 ) | ( n240 ) ;
 assign n117 = ( n76  &  Ni35  &  (~ n1063) ) | ( n76  &  n118  &  (~ n1063) ) ;
 assign n119 = ( n108  &  n83  &  n82 ) | ( n108  &  n83  &  n107 ) ;
 assign n120 = ( n108  &  n86  &  n85 ) | ( n108  &  n86  &  n107 ) ;
 assign n122 = ( n88 ) | ( n202 ) ;
 assign n121 = ( n89  &  (~ Ni35)  &  (~ n1063) ) | ( n89  &  n122  &  (~ n1063) ) ;
 assign n124 = ( n92 ) | ( n240 ) ;
 assign n123 = ( n93  &  (~ Ni35)  &  (~ n1063) ) | ( n93  &  n124  &  (~ n1063) ) ;
 assign n126 = ( n96 ) | ( n202 ) ;
 assign n125 = ( n97  &  Ni35  &  (~ n1063) ) | ( n97  &  n126  &  (~ n1063) ) ;
 assign n128 = ( n100 ) | ( n240 ) ;
 assign n127 = ( n101  &  Ni35  &  (~ n1063) ) | ( n101  &  n128  &  (~ n1063) ) ;
 assign n130 = ( Ni47 ) | ( n320 ) ;
 assign n129 = ( (~ Ni44)  &  (~ Ni41) ) | ( n130  &  (~ Ni41) ) ;
 assign n133 = ( Ni45 ) | ( n320 ) ;
 assign n132 = ( (~ Ni44)  &  (~ Ni41) ) | ( n133  &  (~ Ni41) ) ;
 assign n134 = ( Ni44  &  (~ Ni41) ) | ( n130  &  (~ Ni41) ) ;
 assign n135 = ( Ni44  &  (~ Ni41) ) | ( n133  &  (~ Ni41) ) ;
 assign n136 = ( (~ Ni14)  &  (~ n3569) ) | ( n3545  &  (~ n3569)  &  (~ Ni2) ) ;
 assign Nv10056 = ( (~ n136) ) ;
 assign n137 = ( (~ Ni13)  &  n3564 ) | ( (~ n3540)  &  n3564  &  (~ n3568) ) ;
 assign Nv10068 = ( (~ n137) ) ;
 assign n140 = ( (~ Pi25) ) | ( Ni10 ) ;
 assign n138 = ( n140  &  (~ Ni10)  &  (~ Ni9) ) | ( n140  &  (~ Ni9)  &  (~ n3837) ) ;
 assign n142 = ( n3555  &  (~ Ni9) ) | ( (~ n3540)  &  n3555  &  (~ n3844) ) ;
 assign Nv10112 = ( (~ n142) ) ;
 assign n143 = ( n2049  &  (~ Ni8) ) | ( (~ Ni8)  &  n3540 ) | ( n2049  &  n3549 ) | ( n3540  &  n3549 ) ;
 assign Nv10126 = ( (~ n143) ) ;
 assign n144 = ( Ni6  &  n3548  &  (~ n4805) ) | ( n3544  &  n3548  &  (~ n4805) ) ;
 assign Nv10143 = ( (~ n144) ) ;
 assign n145 = ( Ni6  &  (~ n3488)  &  (~ n3705) ) | ( Ni6  &  (~ n3705)  &  (~ n3876) ) ;
 assign n149 = ( n3542  &  n3543  &  n2066 ) | ( n3542  &  n3543  &  n3539 ) ;
 assign Nv10247 = ( (~ n149) ) ;
 assign n150 = ( (~ Ni37)  &  Ni38 ) ;
 assign n153 = ( (~ Ni32) ) | ( (~ Ni30) ) ;
 assign n157 = ( (~ n18) ) | ( (~ Ni33) ) ;
 assign n158 = ( n3615  &  n3616  &  n3611 ) | ( n3615  &  n3616  &  n3540 ) ;
 assign n159 = ( n3540  &  (~ n3604)  &  n3608 ) | ( n3601  &  (~ n3604)  &  n3608 ) ;
 assign n160 = ( Pi23 ) | ( Pi24 ) ;
 assign n161 = ( Pi26 ) | ( Pi27 ) ;
 assign n162 = ( (~ n153)  &  n3592 ) | ( n3592  &  n3590  &  n3591 ) ;
 assign N_N13960 = ( (~ n162) ) ;
 assign n163 = ( Ni34  &  Ni30 ) | ( Ni34  &  Ni32 ) | ( Ni34  &  Ni31 ) ;
 assign n166 = ( (~ Pi21) ) | ( (~ n2328) ) ;
 assign n164 = ( n160  &  Ni30  &  n166 ) | ( Ni30  &  n166  &  (~ n953) ) ;
 assign n168 = ( Pi24 ) | ( (~ Pi23) ) ;
 assign n167 = ( Ni30  &  n166  &  n168 ) | ( Ni30  &  n166  &  (~ n953) ) ;
 assign n171 = ( (~ n3640) ) | ( n3843 ) | ( n3863 ) ;
 assign n169 = ( n171  &  (~ n1471) ) | ( (~ n1471)  &  (~ n4827) ) ;
 assign n173 = ( n171  &  (~ n1866) ) | ( (~ n1866)  &  (~ n3342) ) | ( (~ n1866)  &  (~ n4827) ) ;
 assign n177 = ( n3843 ) | ( n3592 ) ;
 assign n178 = ( (~ Ni32) ) | ( (~ Ni31) ) ;
 assign n176 = ( n177  &  n178 ) ;
 assign n180 = ( n3666  &  n2083 ) ;
 assign n179 = ( n180  &  (~ n2068) ) | ( (~ Ni33)  &  (~ n2068) ) ;
 assign n183 = ( n180  &  (~ n2068) ) | ( Ni33  &  (~ n2068) ) ;
 assign n184 = ( (~ n23)  &  (~ n153) ) | ( Ni31  &  (~ n153) ) ;
 assign n188 = ( (~ Pi20)  &  n3060 ) | ( n3060  &  (~ n3869) ) ;
 assign n190 = ( (~ Ni35)  &  (~ Ni30) ) ;
 assign n193 = ( n171 ) | ( (~ n4827) ) ;
 assign n192 = ( Pi22  &  n193 ) | ( Pi22  &  (~ n3342) ) ;
 assign n195 = ( n2069  &  Ni45 ) | ( n2069  &  n2068 ) ;
 assign n196 = ( n178  &  (~ n3687) ) ;
 assign n194 = ( n195  &  n196 ) ;
 assign n200 = ( (~ Ni37) ) | ( Ni38 ) ;
 assign n198 = ( n269  &  Ni40 ) | ( n269  &  n457 ) ;
 assign n197 = ( (~ Ni37)  &  n200 ) | ( n200  &  n198 ) ;
 assign n202 = ( (~ n2961) ) | ( n3722 ) ;
 assign n201 = ( n43  &  n198 ) | ( n43  &  n202 ) ;
 assign n203 = ( n43  &  (~ n150)  &  n197 ) | ( n43  &  n198  &  n197 ) ;
 assign n206 = ( n198  &  n203 ) | ( n63  &  n203 ) | ( n198  &  n2087 ) | ( n63  &  n2087 ) ;
 assign n205 = ( n197  &  n206  &  Ni35 ) | ( n197  &  n206  &  n201 ) ;
 assign n207 = ( (~ Ni37)  &  Ni36 ) | ( (~ Ni37)  &  n44  &  (~ n2961) ) ;
 assign n212 = ( n510 ) | ( n511 ) ;
 assign n210 = ( (~ Ni36)  &  n207 ) ;
 assign n211 = ( Ni35 ) | ( n2094 ) ;
 assign n209 = ( n212  &  n210 ) | ( n212  &  n211 ) ;
 assign n214 = ( n272  &  Ni40 ) | ( n272  &  n463 ) ;
 assign n213 = ( (~ Ni37)  &  n200 ) | ( n200  &  n214 ) ;
 assign n216 = ( n3718 ) | ( n3724 ) ;
 assign n215 = ( n216  &  n213  &  n214 ) | ( n216  &  n213  &  n202 ) ;
 assign n218 = ( Ni38 ) | ( n3718 ) ;
 assign n217 = ( (~ n150)  &  n213  &  n218 ) | ( n214  &  n213  &  n218 ) ;
 assign n220 = ( n214  &  n213 ) | ( n464  &  n213 ) | ( n214  &  n275 ) | ( n464  &  n275 ) ;
 assign n221 = ( n217  &  n215 ) | ( n3726  &  n215 ) | ( n217  &  n397 ) | ( n3726  &  n397 ) ;
 assign n219 = ( n220  &  n221 ) ;
 assign n223 = ( n278  &  Ni40 ) | ( n278  &  n470 ) ;
 assign n222 = ( (~ Ni37)  &  n200 ) | ( n200  &  n223 ) ;
 assign n225 = ( n3749 ) | ( n3724 ) ;
 assign n224 = ( n225  &  n222  &  n223 ) | ( n225  &  n222  &  n202 ) ;
 assign n227 = ( Ni38 ) | ( n3749 ) ;
 assign n226 = ( (~ n150)  &  n222  &  n227 ) | ( n223  &  n222  &  n227 ) ;
 assign n229 = ( n224  &  n222 ) | ( n400  &  n222 ) | ( n224  &  n281 ) | ( n400  &  n281 ) ;
 assign n230 = ( n226  &  n223 ) | ( n3721  &  n223 ) | ( n226  &  n471 ) | ( n3721  &  n471 ) ;
 assign n228 = ( n229  &  n230 ) ;
 assign n231 = ( n219  &  n228 ) ;
 assign n234 = ( n231  &  n205 ) | ( n3719  &  n205 ) | ( n231  &  n288 ) | ( n3719  &  n288 ) ;
 assign n233 = ( Ni32 ) | ( n841 ) ;
 assign n232 = ( n209  &  n234  &  n198 ) | ( n209  &  n234  &  n233 ) ;
 assign n236 = ( n18 ) | ( (~ n1063) ) ;
 assign n235 = ( n236  &  n232  &  n18 ) | ( n236  &  n232  &  n205 ) ;
 assign n238 = ( n269  &  Ni40 ) | ( n269  &  n483 ) ;
 assign n237 = ( (~ Ni37)  &  n200 ) | ( n200  &  n238 ) ;
 assign n240 = ( (~ n2962) ) | ( n3722 ) ;
 assign n239 = ( n43  &  n238 ) | ( n43  &  n240 ) ;
 assign n241 = ( n43  &  (~ n150)  &  n237 ) | ( n43  &  n238  &  n237 ) ;
 assign n243 = ( n238  &  n241 ) | ( n63  &  n241 ) | ( n238  &  n2087 ) | ( n63  &  n2087 ) ;
 assign n242 = ( n237  &  n243  &  Ni35 ) | ( n237  &  n243  &  n239 ) ;
 assign n244 = ( (~ Ni37)  &  Ni36 ) | ( (~ Ni37)  &  n44  &  (~ n2962) ) ;
 assign n247 = ( (~ Ni36)  &  n244 ) ;
 assign n246 = ( n212  &  n247 ) | ( n212  &  n211 ) ;
 assign n249 = ( n272  &  Ni40 ) | ( n272  &  n488 ) ;
 assign n248 = ( (~ Ni37)  &  n200 ) | ( n200  &  n249 ) ;
 assign n251 = ( n3718 ) | ( n3725 ) ;
 assign n250 = ( n251  &  n248  &  n249 ) | ( n251  &  n248  &  n240 ) ;
 assign n252 = ( (~ n150)  &  n218  &  n248 ) | ( n218  &  n249  &  n248 ) ;
 assign n254 = ( n249  &  n248 ) | ( n464  &  n248 ) | ( n249  &  n275 ) | ( n464  &  n275 ) ;
 assign n255 = ( n252  &  n250 ) | ( n3726  &  n250 ) | ( n252  &  n397 ) | ( n3726  &  n397 ) ;
 assign n253 = ( n254  &  n255 ) ;
 assign n257 = ( n278  &  Ni40 ) | ( n278  &  n494 ) ;
 assign n256 = ( (~ Ni37)  &  n200 ) | ( n200  &  n257 ) ;
 assign n259 = ( n3749 ) | ( n3725 ) ;
 assign n258 = ( n259  &  n256  &  n257 ) | ( n259  &  n256  &  n240 ) ;
 assign n260 = ( (~ n150)  &  n227  &  n256 ) | ( n227  &  n257  &  n256 ) ;
 assign n262 = ( n258  &  n256 ) | ( n400  &  n256 ) | ( n258  &  n281 ) | ( n400  &  n281 ) ;
 assign n263 = ( n260  &  n257 ) | ( n3721  &  n257 ) | ( n260  &  n471 ) | ( n3721  &  n471 ) ;
 assign n261 = ( n262  &  n263 ) ;
 assign n264 = ( n253  &  n261 ) ;
 assign n266 = ( n264  &  n242 ) | ( n3719  &  n242 ) | ( n264  &  n288 ) | ( n3719  &  n288 ) ;
 assign n265 = ( n246  &  n266  &  n238 ) | ( n246  &  n266  &  n233 ) ;
 assign n267 = ( n236  &  n265  &  n18 ) | ( n236  &  n265  &  n242 ) ;
 assign n269 = ( n313  &  (~ Ni41) ) ;
 assign n268 = ( n43  &  n200  &  n269 ) | ( n43  &  n200  &  (~ Ni38) ) ;
 assign n272 = ( (~ n130)  &  (~ Ni41) ) ;
 assign n271 = ( n200  &  n218  &  n272 ) | ( n200  &  n218  &  (~ Ni38) ) ;
 assign n273 = ( n272  &  n200 ) ;
 assign n275 = ( Ni32 ) | ( (~ Ni36) ) ;
 assign n276 = ( Ni32 ) | ( Ni36 ) ;
 assign n274 = ( n273  &  n271 ) | ( n275  &  n271 ) | ( n273  &  n276 ) | ( n275  &  n276 ) ;
 assign n278 = ( (~ n133)  &  (~ Ni41) ) ;
 assign n277 = ( n200  &  n227  &  n278 ) | ( n200  &  n227  &  (~ Ni38) ) ;
 assign n281 = ( (~ Ni32) ) | ( (~ Ni36) ) ;
 assign n279 = ( (~ Ni32)  &  n278 ) | ( n278  &  n277 ) | ( (~ Ni32)  &  n281 ) | ( n277  &  n281 ) ;
 assign n282 = ( (~ n274)  &  (~ n3719) ) | ( (~ n279)  &  (~ n3719) ) ;
 assign n290 = ( n269  &  n510 ) | ( n233  &  n510 ) | ( n269  &  n2094 ) | ( n233  &  n2094 ) ;
 assign n287 = ( (~ Ni36)  &  n268 ) | ( n269  &  n268 ) ;
 assign n288 = ( (~ n18) ) | ( n2068 ) ;
 assign n286 = ( (~ n282)  &  n290  &  n287 ) | ( (~ n282)  &  n290  &  n288 ) ;
 assign n291 = ( n236  &  n286  &  n18 ) | ( n236  &  n286  &  n287 ) ;
 assign n294 = ( Pi22 ) | ( (~ Ni30) ) ;
 assign n292 = ( Pi22  &  n294 ) | ( (~ n178)  &  n294 ) ;
 assign n295 = ( n292  &  Pi22 ) | ( n292  &  n18 ) ;
 assign n297 = ( Pi21 ) | ( (~ Ni30) ) ;
 assign n296 = ( n297  &  Ni31 ) | ( n297  &  Pi21 ) ;
 assign n299 = ( n2073  &  n296 ) ;
 assign n298 = ( n299  &  Pi21 ) | ( n299  &  n18 ) ;
 assign n301 = ( Pi21  &  (~ Pi20) ) ;
 assign n300 = ( (~ n228)  &  n301 ) ;
 assign n304 = ( Pi20  &  Pi21 ) ;
 assign n303 = ( (~ Pi22)  &  n300 ) | ( (~ Pi22)  &  (~ n261)  &  n304 ) ;
 assign n308 = ( n295  &  Pi22 ) | ( n295  &  n279 ) ;
 assign n307 = ( n298  &  n308  &  Pi21 ) | ( n298  &  n308  &  n274 ) ;
 assign n311 = ( Pi19  &  n307 ) | ( (~ Pi19)  &  (~ n3732) ) | ( n307  &  (~ n3732) ) ;
 assign n312 = ( n291  &  n235 ) | ( n1250  &  n235 ) | ( n291  &  n891 ) | ( n1250  &  n891 ) ;
 assign n310 = ( Pi19 ) | ( n3729 ) ;
 assign n309 = ( n311  &  n312  &  n267 ) | ( n311  &  n312  &  n310 ) ;
 assign n313 = ( n104  &  (~ Ni42) ) ;
 assign n315 = ( n313  &  Ni40 ) | ( n313  &  n564 ) ;
 assign n314 = ( (~ Ni37)  &  n200 ) | ( n200  &  n315 ) ;
 assign n316 = ( n43  &  n315 ) | ( n43  &  n202 ) ;
 assign n317 = ( n43  &  (~ n150)  &  n314 ) | ( n43  &  n315  &  n314 ) ;
 assign n319 = ( n315  &  n317 ) | ( n63  &  n317 ) | ( n315  &  n2087 ) | ( n63  &  n2087 ) ;
 assign n318 = ( n314  &  n319  &  Ni35 ) | ( n314  &  n319  &  n316 ) ;
 assign n320 = ( Ni43 ) | ( Ni42 ) ;
 assign n322 = ( (~ n130)  &  n568 ) | ( (~ n130)  &  Ni40 ) ;
 assign n321 = ( (~ Ni37)  &  n200 ) | ( n200  &  n322 ) ;
 assign n323 = ( n216  &  n321  &  n322 ) | ( n216  &  n321  &  n202 ) ;
 assign n324 = ( (~ n150)  &  n218  &  n321 ) | ( n218  &  n322  &  n321 ) ;
 assign n326 = ( n322  &  n321 ) | ( n464  &  n321 ) | ( n322  &  n275 ) | ( n464  &  n275 ) ;
 assign n327 = ( n324  &  n323 ) | ( n3726  &  n323 ) | ( n324  &  n397 ) | ( n3726  &  n397 ) ;
 assign n325 = ( n326  &  n327 ) ;
 assign n329 = ( (~ n133)  &  n573 ) | ( (~ n133)  &  Ni40 ) ;
 assign n328 = ( (~ Ni37)  &  n200 ) | ( n200  &  n329 ) ;
 assign n330 = ( n225  &  n328  &  n329 ) | ( n225  &  n328  &  n202 ) ;
 assign n331 = ( (~ n150)  &  n227  &  n328 ) | ( n227  &  n329  &  n328 ) ;
 assign n333 = ( n330  &  n328 ) | ( n400  &  n328 ) | ( n330  &  n281 ) | ( n400  &  n281 ) ;
 assign n334 = ( n331  &  n329 ) | ( n3721  &  n329 ) | ( n331  &  n471 ) | ( n3721  &  n471 ) ;
 assign n332 = ( n333  &  n334 ) ;
 assign n335 = ( n325  &  n332 ) ;
 assign n337 = ( n335  &  n318 ) | ( n3719  &  n318 ) | ( n335  &  n288 ) | ( n3719  &  n288 ) ;
 assign n336 = ( n209  &  n337  &  n315 ) | ( n209  &  n337  &  n233 ) ;
 assign n338 = ( n236  &  n336  &  n18 ) | ( n236  &  n336  &  n318 ) ;
 assign n340 = ( n313  &  Ni40 ) | ( n313  &  n585 ) ;
 assign n339 = ( (~ Ni37)  &  n200 ) | ( n200  &  n340 ) ;
 assign n341 = ( n43  &  n340 ) | ( n43  &  n240 ) ;
 assign n342 = ( n43  &  (~ n150)  &  n339 ) | ( n43  &  n340  &  n339 ) ;
 assign n344 = ( n340  &  n342 ) | ( n63  &  n342 ) | ( n340  &  n2087 ) | ( n63  &  n2087 ) ;
 assign n343 = ( n339  &  n344  &  Ni35 ) | ( n339  &  n344  &  n341 ) ;
 assign n346 = ( (~ n130)  &  n589 ) | ( (~ n130)  &  Ni40 ) ;
 assign n345 = ( (~ Ni37)  &  n200 ) | ( n200  &  n346 ) ;
 assign n347 = ( n251  &  n345  &  n346 ) | ( n251  &  n345  &  n240 ) ;
 assign n348 = ( (~ n150)  &  n218  &  n345 ) | ( n218  &  n346  &  n345 ) ;
 assign n350 = ( n346  &  n345 ) | ( n464  &  n345 ) | ( n346  &  n275 ) | ( n464  &  n275 ) ;
 assign n351 = ( n348  &  n347 ) | ( n3726  &  n347 ) | ( n348  &  n397 ) | ( n3726  &  n397 ) ;
 assign n349 = ( n350  &  n351 ) ;
 assign n353 = ( (~ n133)  &  n594 ) | ( (~ n133)  &  Ni40 ) ;
 assign n352 = ( (~ Ni37)  &  n200 ) | ( n200  &  n353 ) ;
 assign n354 = ( n259  &  n352  &  n353 ) | ( n259  &  n352  &  n240 ) ;
 assign n355 = ( (~ n150)  &  n227  &  n352 ) | ( n227  &  n353  &  n352 ) ;
 assign n357 = ( n354  &  n352 ) | ( n400  &  n352 ) | ( n354  &  n281 ) | ( n400  &  n281 ) ;
 assign n358 = ( n355  &  n353 ) | ( n3721  &  n353 ) | ( n355  &  n471 ) | ( n3721  &  n471 ) ;
 assign n356 = ( n357  &  n358 ) ;
 assign n359 = ( n349  &  n356 ) ;
 assign n361 = ( n359  &  n343 ) | ( n3719  &  n343 ) | ( n359  &  n288 ) | ( n3719  &  n288 ) ;
 assign n360 = ( n246  &  n361  &  n340 ) | ( n246  &  n361  &  n233 ) ;
 assign n362 = ( n236  &  n360  &  n18 ) | ( n236  &  n360  &  n343 ) ;
 assign n363 = ( n43  &  n200  &  n313 ) | ( n43  &  n200  &  (~ Ni38) ) ;
 assign n364 = ( (~ n130)  &  n200  &  n218 ) | ( n200  &  n218  &  (~ Ni38) ) ;
 assign n366 = ( (~ n130)  &  n200 ) ;
 assign n367 = ( n366  &  n364 ) | ( n275  &  n364 ) | ( n366  &  n276 ) | ( n275  &  n276 ) ;
 assign n368 = ( (~ n133)  &  n200  &  n227 ) | ( n200  &  n227  &  (~ Ni38) ) ;
 assign n370 = ( (~ Ni32)  &  (~ n133) ) | ( (~ Ni32)  &  n281 ) | ( (~ n133)  &  n368 ) | ( n281  &  n368 ) ;
 assign n371 = ( (~ n367)  &  (~ n3719) ) | ( (~ n370)  &  (~ n3719) ) ;
 assign n377 = ( n313  &  n510 ) | ( n233  &  n510 ) | ( n313  &  n2094 ) | ( n233  &  n2094 ) ;
 assign n375 = ( (~ Ni36)  &  n363 ) | ( n313  &  n363 ) ;
 assign n374 = ( n288  &  (~ n371)  &  n377 ) | ( (~ n371)  &  n377  &  n375 ) ;
 assign n378 = ( n236  &  n374  &  n18 ) | ( n236  &  n374  &  n375 ) ;
 assign n379 = ( n301  &  (~ n332) ) ;
 assign n381 = ( (~ Pi22)  &  n379 ) | ( (~ Pi22)  &  n304  &  (~ n356) ) ;
 assign n384 = ( n295  &  Pi22 ) | ( n295  &  n370 ) ;
 assign n383 = ( n298  &  n384  &  Pi21 ) | ( n298  &  n384  &  n367 ) ;
 assign n386 = ( Pi19  &  n383 ) | ( (~ Pi19)  &  (~ n3756) ) | ( n383  &  (~ n3756) ) ;
 assign n387 = ( n378  &  n338 ) | ( n1250  &  n338 ) | ( n378  &  n891 ) | ( n1250  &  n891 ) ;
 assign n385 = ( n386  &  n387  &  n362 ) | ( n386  &  n387  &  n310 ) ;
 assign n388 = ( n203  &  Ni35 ) | ( n203  &  n201 ) ;
 assign n390 = ( Ni38 ) | ( n44 ) ;
 assign n391 = ( (~ Ni37)  &  (~ Ni38) ) ;
 assign n389 = ( n390  &  n391 ) ;
 assign n394 = ( n389 ) | ( n511 ) ;
 assign n393 = ( n389  &  n207 ) ;
 assign n392 = ( n394  &  n393 ) | ( n394  &  n211 ) ;
 assign n396 = ( Ni32 ) | ( (~ n2199) ) ;
 assign n397 = ( Ni32 ) | ( Ni35 ) ;
 assign n395 = ( n217  &  n215 ) | ( n396  &  n215 ) | ( n217  &  n397 ) | ( n396  &  n397 ) ;
 assign n399 = ( n694  &  n281 ) ;
 assign n400 = ( (~ Ni32) ) | ( Ni35 ) ;
 assign n398 = ( n226  &  n224 ) | ( n399  &  n224 ) | ( n226  &  n400 ) | ( n399  &  n400 ) ;
 assign n401 = ( n395  &  n398 ) ;
 assign n403 = ( n401  &  n388 ) | ( n3719  &  n388 ) | ( n401  &  n288 ) | ( n3719  &  n288 ) ;
 assign n402 = ( n392  &  n403  &  n198 ) | ( n392  &  n403  &  n233 ) ;
 assign n404 = ( n236  &  n402  &  n18 ) | ( n236  &  n402  &  n388 ) ;
 assign n405 = ( n241  &  Ni35 ) | ( n241  &  n239 ) ;
 assign n407 = ( n389  &  n244 ) ;
 assign n406 = ( n394  &  n407 ) | ( n394  &  n211 ) ;
 assign n408 = ( n252  &  n250 ) | ( n396  &  n250 ) | ( n252  &  n397 ) | ( n396  &  n397 ) ;
 assign n409 = ( n260  &  n258 ) | ( n399  &  n258 ) | ( n260  &  n400 ) | ( n399  &  n400 ) ;
 assign n410 = ( n408  &  n409 ) ;
 assign n412 = ( n410  &  n405 ) | ( n3719  &  n405 ) | ( n410  &  n288 ) | ( n3719  &  n288 ) ;
 assign n411 = ( n406  &  n412  &  n238 ) | ( n406  &  n412  &  n233 ) ;
 assign n413 = ( n236  &  n411  &  n18 ) | ( n236  &  n411  &  n405 ) ;
 assign n415 = ( n3987  &  n277 ) | ( n3987  &  n3482 ) ;
 assign n416 = ( n269  &  n389 ) | ( n233  &  n389 ) | ( n269  &  n2094 ) | ( n233  &  n2094 ) ;
 assign n414 = ( n415  &  n416  &  n268 ) | ( n415  &  n416  &  n288 ) ;
 assign n417 = ( n236  &  n414  &  n18 ) | ( n236  &  n414  &  n268 ) ;
 assign n418 = ( n301  &  (~ n398) ) ;
 assign n420 = ( (~ Pi22)  &  n418 ) | ( (~ Pi22)  &  n304  &  (~ n409) ) ;
 assign n423 = ( n295  &  Pi22 ) | ( n295  &  n277 ) ;
 assign n422 = ( n298  &  n423  &  Pi21 ) | ( n298  &  n423  &  n271 ) ;
 assign n425 = ( Pi19  &  n422 ) | ( (~ Pi19)  &  (~ n3746) ) | ( n422  &  (~ n3746) ) ;
 assign n426 = ( n417  &  n404 ) | ( n1250  &  n404 ) | ( n417  &  n891 ) | ( n1250  &  n891 ) ;
 assign n424 = ( n425  &  n426  &  n413 ) | ( n425  &  n426  &  n310 ) ;
 assign n427 = ( n317  &  Ni35 ) | ( n317  &  n316 ) ;
 assign n428 = ( n324  &  n323 ) | ( n396  &  n323 ) | ( n324  &  n397 ) | ( n396  &  n397 ) ;
 assign n429 = ( n331  &  n330 ) | ( n399  &  n330 ) | ( n331  &  n400 ) | ( n399  &  n400 ) ;
 assign n430 = ( n428  &  n429 ) ;
 assign n432 = ( n430  &  n427 ) | ( n3719  &  n427 ) | ( n430  &  n288 ) | ( n3719  &  n288 ) ;
 assign n431 = ( n392  &  n432  &  n315 ) | ( n392  &  n432  &  n233 ) ;
 assign n433 = ( n236  &  n431  &  n18 ) | ( n236  &  n431  &  n427 ) ;
 assign n434 = ( n342  &  Ni35 ) | ( n342  &  n341 ) ;
 assign n435 = ( n348  &  n347 ) | ( n396  &  n347 ) | ( n348  &  n397 ) | ( n396  &  n397 ) ;
 assign n436 = ( n355  &  n354 ) | ( n399  &  n354 ) | ( n355  &  n400 ) | ( n399  &  n400 ) ;
 assign n437 = ( n435  &  n436 ) ;
 assign n439 = ( n437  &  n434 ) | ( n3719  &  n434 ) | ( n437  &  n288 ) | ( n3719  &  n288 ) ;
 assign n438 = ( n406  &  n439  &  n340 ) | ( n406  &  n439  &  n233 ) ;
 assign n440 = ( n236  &  n438  &  n18 ) | ( n236  &  n438  &  n434 ) ;
 assign n442 = ( n3988  &  n368 ) | ( n3988  &  n3482 ) ;
 assign n443 = ( n313  &  n389 ) | ( n233  &  n389 ) | ( n313  &  n2094 ) | ( n233  &  n2094 ) ;
 assign n441 = ( n442  &  n443  &  n363 ) | ( n442  &  n443  &  n288 ) ;
 assign n444 = ( n236  &  n441  &  n18 ) | ( n236  &  n441  &  n363 ) ;
 assign n445 = ( n301  &  (~ n429) ) ;
 assign n447 = ( (~ Pi22)  &  n445 ) | ( (~ Pi22)  &  n304  &  (~ n436) ) ;
 assign n450 = ( n295  &  Pi22 ) | ( n295  &  n368 ) ;
 assign n449 = ( n298  &  n450  &  Pi21 ) | ( n298  &  n450  &  n364 ) ;
 assign n452 = ( Pi19  &  n449 ) | ( (~ Pi19)  &  (~ n3766) ) | ( n449  &  (~ n3766) ) ;
 assign n453 = ( n444  &  n433 ) | ( n1250  &  n433 ) | ( n444  &  n891 ) | ( n1250  &  n891 ) ;
 assign n451 = ( n452  &  n453  &  n440 ) | ( n452  &  n453  &  n310 ) ;
 assign n455 = ( n457 ) | ( (~ Ni37)  &  n202 ) ;
 assign n454 = ( n200  &  n43  &  n455 ) ;
 assign n457 = ( (~ n38)  &  (~ n2078) ) ;
 assign n456 = ( n454  &  n457 ) | ( n454  &  n63 ) ;
 assign n458 = ( (~ Ni32)  &  (~ n200) ) | ( (~ Ni32)  &  (~ n216) ) | ( (~ Ni32)  &  (~ n3971) ) ;
 assign n463 = ( (~ n129)  &  (~ Ni41) ) ;
 assign n464 = ( Ni32 ) | ( n63 ) ;
 assign n462 = ( (~ n458)  &  n463 ) | ( (~ n458)  &  n464 ) ;
 assign n466 = ( Ni32  &  (~ n200) ) | ( Ni32  &  (~ n225) ) | ( Ni32  &  (~ n3970) ) ;
 assign n470 = ( (~ n132)  &  (~ Ni41) ) ;
 assign n471 = ( Ni37 ) | ( n281 ) ;
 assign n469 = ( (~ n466)  &  n470 ) | ( (~ n466)  &  n471 ) ;
 assign n473 = ( (~ n462)  &  (~ n3719) ) | ( (~ n469)  &  (~ n3719) ) ;
 assign n478 = ( n457  &  n210 ) | ( n233  &  n210 ) | ( n457  &  n2094 ) | ( n233  &  n2094 ) ;
 assign n476 = ( n288  &  (~ n473)  &  n478 ) | ( n456  &  (~ n473)  &  n478 ) ;
 assign n479 = ( n236  &  n476  &  n18 ) | ( n236  &  n476  &  n456 ) ;
 assign n481 = ( n483 ) | ( (~ Ni37)  &  n240 ) ;
 assign n480 = ( n200  &  n43  &  n481 ) ;
 assign n483 = ( (~ n42)  &  (~ n2078) ) ;
 assign n482 = ( n480  &  n483 ) | ( n480  &  n63 ) ;
 assign n484 = ( (~ Ni32)  &  (~ n200) ) | ( (~ Ni32)  &  (~ n251) ) | ( (~ Ni32)  &  (~ n3973) ) ;
 assign n488 = ( (~ n134)  &  (~ Ni41) ) ;
 assign n487 = ( n464  &  (~ n484) ) | ( (~ n484)  &  n488 ) ;
 assign n490 = ( Ni32  &  (~ n200) ) | ( Ni32  &  (~ n259) ) | ( Ni32  &  (~ n3972) ) ;
 assign n494 = ( (~ n135)  &  (~ Ni41) ) ;
 assign n493 = ( n471  &  (~ n490) ) | ( (~ n490)  &  n494 ) ;
 assign n496 = ( (~ n487)  &  (~ n3719) ) | ( (~ n493)  &  (~ n3719) ) ;
 assign n501 = ( n483  &  n247 ) | ( n233  &  n247 ) | ( n483  &  n2094 ) | ( n233  &  n2094 ) ;
 assign n499 = ( n288  &  (~ n496)  &  n501 ) | ( n482  &  (~ n496)  &  n501 ) ;
 assign n502 = ( n236  &  n499  &  n18 ) | ( n236  &  n499  &  n482 ) ;
 assign n504 = ( n269  &  n457 ) | ( n269  &  (~ Ni40) ) ;
 assign n503 = ( (~ Ni37)  &  n200 ) | ( n200  &  n504 ) ;
 assign n505 = ( n43  &  (~ n150)  &  n503 ) | ( n43  &  n504  &  n503 ) ;
 assign n506 = ( n43  &  n504 ) | ( n43  &  n202 ) ;
 assign n508 = ( n504  &  n505 ) | ( n63  &  n505 ) | ( n504  &  n2199 ) | ( n63  &  n2199 ) ;
 assign n507 = ( (~ Ni35)  &  n503  &  n508 ) | ( n503  &  n506  &  n508 ) ;
 assign n510 = ( (~ Ni36)  &  n389 ) ;
 assign n511 = ( (~ Ni35) ) | ( n2094 ) ;
 assign n509 = ( n510  &  n210 ) | ( n211  &  n210 ) | ( n510  &  n511 ) | ( n211  &  n511 ) ;
 assign n513 = ( n272  &  n463 ) | ( n272  &  (~ Ni40) ) ;
 assign n512 = ( (~ Ni37)  &  n200 ) | ( n200  &  n513 ) ;
 assign n514 = ( (~ n150)  &  n218  &  n512 ) | ( n218  &  n513  &  n512 ) ;
 assign n515 = ( n216  &  n512  &  n513 ) | ( n216  &  n512  &  n202 ) ;
 assign n517 = ( n513  &  n512 ) | ( n464  &  n512 ) | ( n513  &  n275 ) | ( n464  &  n275 ) ;
 assign n518 = ( n514  &  n515 ) | ( n3740  &  n515 ) | ( n514  &  n691 ) | ( n3740  &  n691 ) ;
 assign n516 = ( n517  &  n518 ) ;
 assign n520 = ( n278  &  n470 ) | ( n278  &  (~ Ni40) ) ;
 assign n519 = ( (~ Ni37)  &  n200 ) | ( n200  &  n520 ) ;
 assign n521 = ( (~ n150)  &  n227  &  n519 ) | ( n227  &  n520  &  n519 ) ;
 assign n522 = ( n225  &  n519  &  n520 ) | ( n225  &  n519  &  n202 ) ;
 assign n524 = ( n522  &  n519 ) | ( n694  &  n519 ) | ( n522  &  n281 ) | ( n694  &  n281 ) ;
 assign n525 = ( n521  &  n520 ) | ( n3739  &  n520 ) | ( n521  &  n471 ) | ( n3739  &  n471 ) ;
 assign n523 = ( n524  &  n525 ) ;
 assign n526 = ( n516  &  n523 ) ;
 assign n528 = ( n526  &  n507 ) | ( n3719  &  n507 ) | ( n526  &  n288 ) | ( n3719  &  n288 ) ;
 assign n527 = ( n509  &  n528  &  n504 ) | ( n509  &  n528  &  n233 ) ;
 assign n529 = ( n236  &  n527  &  n18 ) | ( n236  &  n527  &  n507 ) ;
 assign n531 = ( n269  &  n483 ) | ( n269  &  (~ Ni40) ) ;
 assign n530 = ( (~ Ni37)  &  n200 ) | ( n200  &  n531 ) ;
 assign n532 = ( n43  &  (~ n150)  &  n530 ) | ( n43  &  n531  &  n530 ) ;
 assign n533 = ( n43  &  n531 ) | ( n43  &  n240 ) ;
 assign n535 = ( n531  &  n532 ) | ( n63  &  n532 ) | ( n531  &  n2199 ) | ( n63  &  n2199 ) ;
 assign n534 = ( (~ Ni35)  &  n530  &  n535 ) | ( n530  &  n533  &  n535 ) ;
 assign n536 = ( n510  &  n247 ) | ( n211  &  n247 ) | ( n510  &  n511 ) | ( n211  &  n511 ) ;
 assign n538 = ( n272  &  n488 ) | ( n272  &  (~ Ni40) ) ;
 assign n537 = ( (~ Ni37)  &  n200 ) | ( n200  &  n538 ) ;
 assign n539 = ( (~ n150)  &  n218  &  n537 ) | ( n218  &  n538  &  n537 ) ;
 assign n540 = ( n251  &  n537  &  n538 ) | ( n251  &  n537  &  n240 ) ;
 assign n542 = ( n538  &  n537 ) | ( n464  &  n537 ) | ( n538  &  n275 ) | ( n464  &  n275 ) ;
 assign n543 = ( n539  &  n540 ) | ( n3740  &  n540 ) | ( n539  &  n691 ) | ( n3740  &  n691 ) ;
 assign n541 = ( n542  &  n543 ) ;
 assign n545 = ( n278  &  n494 ) | ( n278  &  (~ Ni40) ) ;
 assign n544 = ( (~ Ni37)  &  n200 ) | ( n200  &  n545 ) ;
 assign n546 = ( (~ n150)  &  n227  &  n544 ) | ( n227  &  n545  &  n544 ) ;
 assign n547 = ( n259  &  n544  &  n545 ) | ( n259  &  n544  &  n240 ) ;
 assign n549 = ( n547  &  n544 ) | ( n694  &  n544 ) | ( n547  &  n281 ) | ( n694  &  n281 ) ;
 assign n550 = ( n546  &  n545 ) | ( n3739  &  n545 ) | ( n546  &  n471 ) | ( n3739  &  n471 ) ;
 assign n548 = ( n549  &  n550 ) ;
 assign n551 = ( n541  &  n548 ) ;
 assign n553 = ( n551  &  n534 ) | ( n3719  &  n534 ) | ( n551  &  n288 ) | ( n3719  &  n288 ) ;
 assign n552 = ( n536  &  n553  &  n531 ) | ( n536  &  n553  &  n233 ) ;
 assign n554 = ( n236  &  n552  &  n18 ) | ( n236  &  n552  &  n534 ) ;
 assign n555 = ( n301  &  (~ n523) ) ;
 assign n557 = ( (~ Pi22)  &  n555 ) | ( (~ Pi22)  &  n304  &  (~ n548) ) ;
 assign n559 = ( n301  &  (~ n469) ) ;
 assign n560 = ( (~ Pi22)  &  n559 ) | ( (~ Pi22)  &  n304  &  (~ n493) ) ;
 assign n562 = ( n564 ) | ( (~ Ni37)  &  n202 ) ;
 assign n561 = ( n200  &  n43  &  n562 ) ;
 assign n564 = ( n4823  &  n313 ) ;
 assign n563 = ( n561  &  n564 ) | ( n561  &  n63 ) ;
 assign n565 = ( (~ Ni32)  &  (~ n200) ) | ( (~ Ni32)  &  (~ n216) ) | ( (~ Ni32)  &  (~ n3977) ) ;
 assign n568 = ( (~ n130)  &  (~ n129) ) ;
 assign n567 = ( n464  &  (~ n565) ) | ( (~ n565)  &  n568 ) ;
 assign n570 = ( Ni32  &  (~ n200) ) | ( Ni32  &  (~ n225) ) | ( Ni32  &  (~ n3976) ) ;
 assign n573 = ( (~ n133)  &  (~ n132) ) ;
 assign n572 = ( n471  &  (~ n570) ) | ( (~ n570)  &  n573 ) ;
 assign n575 = ( (~ n567)  &  (~ n3719) ) | ( (~ n572)  &  (~ n3719) ) ;
 assign n580 = ( n564  &  n210 ) | ( n233  &  n210 ) | ( n564  &  n2094 ) | ( n233  &  n2094 ) ;
 assign n578 = ( n288  &  (~ n575)  &  n580 ) | ( n563  &  (~ n575)  &  n580 ) ;
 assign n581 = ( n236  &  n578  &  n18 ) | ( n236  &  n578  &  n563 ) ;
 assign n583 = ( n585 ) | ( (~ Ni37)  &  n240 ) ;
 assign n582 = ( n200  &  n43  &  n583 ) ;
 assign n585 = ( n4825  &  n313 ) ;
 assign n584 = ( n582  &  n585 ) | ( n582  &  n63 ) ;
 assign n586 = ( (~ Ni32)  &  (~ n200) ) | ( (~ Ni32)  &  (~ n251) ) | ( (~ Ni32)  &  (~ n3979) ) ;
 assign n589 = ( (~ n130)  &  (~ n134) ) ;
 assign n588 = ( n464  &  (~ n586) ) | ( (~ n586)  &  n589 ) ;
 assign n591 = ( Ni32  &  (~ n200) ) | ( Ni32  &  (~ n259) ) | ( Ni32  &  (~ n3978) ) ;
 assign n594 = ( (~ n133)  &  (~ n135) ) ;
 assign n593 = ( n471  &  (~ n591) ) | ( (~ n591)  &  n594 ) ;
 assign n596 = ( (~ n588)  &  (~ n3719) ) | ( (~ n593)  &  (~ n3719) ) ;
 assign n601 = ( n585  &  n247 ) | ( n233  &  n247 ) | ( n585  &  n2094 ) | ( n233  &  n2094 ) ;
 assign n599 = ( n288  &  (~ n596)  &  n601 ) | ( n584  &  (~ n596)  &  n601 ) ;
 assign n602 = ( n236  &  n599  &  n18 ) | ( n236  &  n599  &  n584 ) ;
 assign n604 = ( n313  &  n564 ) | ( n313  &  (~ Ni40) ) ;
 assign n603 = ( (~ Ni37)  &  n200 ) | ( n200  &  n604 ) ;
 assign n605 = ( n43  &  (~ n150)  &  n603 ) | ( n43  &  n604  &  n603 ) ;
 assign n606 = ( n43  &  n604 ) | ( n43  &  n202 ) ;
 assign n608 = ( n604  &  n605 ) | ( n63  &  n605 ) | ( n604  &  n2199 ) | ( n63  &  n2199 ) ;
 assign n607 = ( (~ Ni35)  &  n603  &  n608 ) | ( n603  &  n606  &  n608 ) ;
 assign n610 = ( (~ n130)  &  n568 ) | ( (~ n130)  &  (~ Ni40) ) ;
 assign n609 = ( (~ Ni37)  &  n200 ) | ( n200  &  n610 ) ;
 assign n611 = ( (~ n150)  &  n218  &  n609 ) | ( n218  &  n610  &  n609 ) ;
 assign n612 = ( n216  &  n609  &  n610 ) | ( n216  &  n609  &  n202 ) ;
 assign n614 = ( n610  &  n609 ) | ( n464  &  n609 ) | ( n610  &  n275 ) | ( n464  &  n275 ) ;
 assign n615 = ( n611  &  n612 ) | ( n3740  &  n612 ) | ( n611  &  n691 ) | ( n3740  &  n691 ) ;
 assign n613 = ( n614  &  n615 ) ;
 assign n617 = ( (~ n133)  &  n573 ) | ( (~ n133)  &  (~ Ni40) ) ;
 assign n616 = ( (~ Ni37)  &  n200 ) | ( n200  &  n617 ) ;
 assign n618 = ( (~ n150)  &  n227  &  n616 ) | ( n227  &  n617  &  n616 ) ;
 assign n619 = ( n225  &  n616  &  n617 ) | ( n225  &  n616  &  n202 ) ;
 assign n621 = ( n619  &  n616 ) | ( n694  &  n616 ) | ( n619  &  n281 ) | ( n694  &  n281 ) ;
 assign n622 = ( n618  &  n617 ) | ( n3739  &  n617 ) | ( n618  &  n471 ) | ( n3739  &  n471 ) ;
 assign n620 = ( n621  &  n622 ) ;
 assign n623 = ( n613  &  n620 ) ;
 assign n625 = ( n623  &  n607 ) | ( n3719  &  n607 ) | ( n623  &  n288 ) | ( n3719  &  n288 ) ;
 assign n624 = ( n509  &  n625  &  n604 ) | ( n509  &  n625  &  n233 ) ;
 assign n626 = ( n236  &  n624  &  n18 ) | ( n236  &  n624  &  n607 ) ;
 assign n628 = ( n313  &  n585 ) | ( n313  &  (~ Ni40) ) ;
 assign n627 = ( (~ Ni37)  &  n200 ) | ( n200  &  n628 ) ;
 assign n629 = ( n43  &  (~ n150)  &  n627 ) | ( n43  &  n628  &  n627 ) ;
 assign n630 = ( n43  &  n628 ) | ( n43  &  n240 ) ;
 assign n632 = ( n628  &  n629 ) | ( n63  &  n629 ) | ( n628  &  n2199 ) | ( n63  &  n2199 ) ;
 assign n631 = ( (~ Ni35)  &  n627  &  n632 ) | ( n627  &  n630  &  n632 ) ;
 assign n634 = ( (~ n130)  &  n589 ) | ( (~ n130)  &  (~ Ni40) ) ;
 assign n633 = ( (~ Ni37)  &  n200 ) | ( n200  &  n634 ) ;
 assign n635 = ( (~ n150)  &  n218  &  n633 ) | ( n218  &  n634  &  n633 ) ;
 assign n636 = ( n251  &  n633  &  n634 ) | ( n251  &  n633  &  n240 ) ;
 assign n638 = ( n634  &  n633 ) | ( n464  &  n633 ) | ( n634  &  n275 ) | ( n464  &  n275 ) ;
 assign n639 = ( n635  &  n636 ) | ( n3740  &  n636 ) | ( n635  &  n691 ) | ( n3740  &  n691 ) ;
 assign n637 = ( n638  &  n639 ) ;
 assign n641 = ( (~ n133)  &  n594 ) | ( (~ n133)  &  (~ Ni40) ) ;
 assign n640 = ( (~ Ni37)  &  n200 ) | ( n200  &  n641 ) ;
 assign n642 = ( (~ n150)  &  n227  &  n640 ) | ( n227  &  n641  &  n640 ) ;
 assign n643 = ( n259  &  n640  &  n641 ) | ( n259  &  n640  &  n240 ) ;
 assign n645 = ( n643  &  n640 ) | ( n694  &  n640 ) | ( n643  &  n281 ) | ( n694  &  n281 ) ;
 assign n646 = ( n642  &  n641 ) | ( n3739  &  n641 ) | ( n642  &  n471 ) | ( n3739  &  n471 ) ;
 assign n644 = ( n645  &  n646 ) ;
 assign n647 = ( n637  &  n644 ) ;
 assign n649 = ( n647  &  n631 ) | ( n3719  &  n631 ) | ( n647  &  n288 ) | ( n3719  &  n288 ) ;
 assign n648 = ( n536  &  n649  &  n628 ) | ( n536  &  n649  &  n233 ) ;
 assign n650 = ( n236  &  n648  &  n18 ) | ( n236  &  n648  &  n631 ) ;
 assign n651 = ( n301  &  (~ n620) ) ;
 assign n653 = ( (~ Pi22)  &  n651 ) | ( (~ Pi22)  &  n304  &  (~ n644) ) ;
 assign n655 = ( n301  &  (~ n572) ) ;
 assign n656 = ( (~ Pi22)  &  n655 ) | ( (~ Pi22)  &  n304  &  (~ n593) ) ;
 assign n658 = ( Pi19  &  n310 ) | ( Pi19  &  n602 ) | ( n310  &  (~ n3759) ) | ( n602  &  (~ n3759) ) ;
 assign n660 = ( n626  &  n650 ) | ( n3776  &  n650 ) | ( n626  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n661 = ( n581 ) | ( n891 ) ;
 assign n657 = ( n658  &  n660  &  n661  &  (~ n3630) ) ;
 assign n663 = ( n63 ) | ( (~ Ni38) ) ;
 assign n662 = ( n454  &  n457 ) | ( n454  &  n663 ) ;
 assign n666 = ( n218 ) | ( n464 ) ;
 assign n665 = ( Ni32 ) | ( n663 ) ;
 assign n664 = ( (~ n458)  &  n463  &  n666 ) | ( (~ n458)  &  n666  &  n665 ) ;
 assign n669 = ( n281 ) | ( n227 ) ;
 assign n668 = ( (~ n150) ) | ( n281 ) ;
 assign n667 = ( (~ n466)  &  n470  &  n669 ) | ( (~ n466)  &  n669  &  n668 ) ;
 assign n670 = ( (~ n664)  &  (~ n3719) ) | ( (~ n667)  &  (~ n3719) ) ;
 assign n675 = ( n457  &  n393 ) | ( n233  &  n393 ) | ( n457  &  n2094 ) | ( n233  &  n2094 ) ;
 assign n673 = ( n288  &  (~ n670)  &  n675 ) | ( n662  &  (~ n670)  &  n675 ) ;
 assign n676 = ( n236  &  n673  &  n18 ) | ( n236  &  n673  &  n662 ) ;
 assign n677 = ( n480  &  n483 ) | ( n480  &  n663 ) ;
 assign n678 = ( (~ n484)  &  n488  &  n666 ) | ( (~ n484)  &  n666  &  n665 ) ;
 assign n679 = ( (~ n490)  &  n494  &  n669 ) | ( (~ n490)  &  n669  &  n668 ) ;
 assign n680 = ( (~ n678)  &  (~ n3719) ) | ( (~ n679)  &  (~ n3719) ) ;
 assign n685 = ( n483  &  n407 ) | ( n233  &  n407 ) | ( n483  &  n2094 ) | ( n233  &  n2094 ) ;
 assign n683 = ( n288  &  (~ n680)  &  n685 ) | ( n677  &  (~ n680)  &  n685 ) ;
 assign n686 = ( n236  &  n683  &  n18 ) | ( n236  &  n683  &  n677 ) ;
 assign n687 = ( (~ Ni35)  &  n505 ) | ( n505  &  n506 ) ;
 assign n688 = ( n389  &  n393 ) | ( n211  &  n393 ) | ( n389  &  n511 ) | ( n211  &  n511 ) ;
 assign n690 = ( Ni32 ) | ( (~ n2087) ) ;
 assign n691 = ( Ni32 ) | ( (~ Ni35) ) ;
 assign n689 = ( n514  &  n515 ) | ( n690  &  n515 ) | ( n514  &  n691 ) | ( n690  &  n691 ) ;
 assign n693 = ( n400  &  n281 ) ;
 assign n694 = ( (~ Ni32) ) | ( (~ Ni35) ) ;
 assign n692 = ( n521  &  n522 ) | ( n693  &  n522 ) | ( n521  &  n694 ) | ( n693  &  n694 ) ;
 assign n695 = ( n689  &  n692 ) ;
 assign n697 = ( n695  &  n687 ) | ( n3719  &  n687 ) | ( n695  &  n288 ) | ( n3719  &  n288 ) ;
 assign n696 = ( n688  &  n697  &  n504 ) | ( n688  &  n697  &  n233 ) ;
 assign n698 = ( n236  &  n696  &  n18 ) | ( n236  &  n696  &  n687 ) ;
 assign n699 = ( (~ Ni35)  &  n532 ) | ( n532  &  n533 ) ;
 assign n700 = ( n389  &  n407 ) | ( n211  &  n407 ) | ( n389  &  n511 ) | ( n211  &  n511 ) ;
 assign n701 = ( n539  &  n540 ) | ( n690  &  n540 ) | ( n539  &  n691 ) | ( n690  &  n691 ) ;
 assign n702 = ( n546  &  n547 ) | ( n693  &  n547 ) | ( n546  &  n694 ) | ( n693  &  n694 ) ;
 assign n703 = ( n701  &  n702 ) ;
 assign n705 = ( n703  &  n699 ) | ( n3719  &  n699 ) | ( n703  &  n288 ) | ( n3719  &  n288 ) ;
 assign n704 = ( n700  &  n705  &  n531 ) | ( n700  &  n705  &  n233 ) ;
 assign n706 = ( n236  &  n704  &  n18 ) | ( n236  &  n704  &  n699 ) ;
 assign n707 = ( n301  &  (~ n692) ) ;
 assign n709 = ( (~ Pi22)  &  n707 ) | ( (~ Pi22)  &  n304  &  (~ n702) ) ;
 assign n711 = ( n301  &  (~ n667) ) ;
 assign n712 = ( (~ Pi22)  &  n711 ) | ( (~ Pi22)  &  n304  &  (~ n679) ) ;
 assign n713 = ( n561  &  n564 ) | ( n561  &  n663 ) ;
 assign n714 = ( (~ n565)  &  n568  &  n666 ) | ( (~ n565)  &  n666  &  n665 ) ;
 assign n715 = ( (~ n570)  &  n573  &  n669 ) | ( (~ n570)  &  n669  &  n668 ) ;
 assign n716 = ( (~ n714)  &  (~ n3719) ) | ( (~ n715)  &  (~ n3719) ) ;
 assign n721 = ( n564  &  n393 ) | ( n233  &  n393 ) | ( n564  &  n2094 ) | ( n233  &  n2094 ) ;
 assign n719 = ( n288  &  (~ n716)  &  n721 ) | ( n713  &  (~ n716)  &  n721 ) ;
 assign n722 = ( n236  &  n719  &  n18 ) | ( n236  &  n719  &  n713 ) ;
 assign n723 = ( n582  &  n585 ) | ( n582  &  n663 ) ;
 assign n724 = ( (~ n586)  &  n589  &  n666 ) | ( (~ n586)  &  n666  &  n665 ) ;
 assign n725 = ( (~ n591)  &  n594  &  n669 ) | ( (~ n591)  &  n669  &  n668 ) ;
 assign n726 = ( (~ n724)  &  (~ n3719) ) | ( (~ n725)  &  (~ n3719) ) ;
 assign n731 = ( n585  &  n407 ) | ( n233  &  n407 ) | ( n585  &  n2094 ) | ( n233  &  n2094 ) ;
 assign n729 = ( n288  &  (~ n726)  &  n731 ) | ( n723  &  (~ n726)  &  n731 ) ;
 assign n732 = ( n236  &  n729  &  n18 ) | ( n236  &  n729  &  n723 ) ;
 assign n733 = ( (~ Ni35)  &  n605 ) | ( n605  &  n606 ) ;
 assign n734 = ( n611  &  n612 ) | ( n690  &  n612 ) | ( n611  &  n691 ) | ( n690  &  n691 ) ;
 assign n735 = ( n618  &  n619 ) | ( n693  &  n619 ) | ( n618  &  n694 ) | ( n693  &  n694 ) ;
 assign n736 = ( n734  &  n735 ) ;
 assign n738 = ( n736  &  n733 ) | ( n3719  &  n733 ) | ( n736  &  n288 ) | ( n3719  &  n288 ) ;
 assign n737 = ( n688  &  n738  &  n604 ) | ( n688  &  n738  &  n233 ) ;
 assign n739 = ( n236  &  n737  &  n18 ) | ( n236  &  n737  &  n733 ) ;
 assign n740 = ( (~ Ni35)  &  n629 ) | ( n629  &  n630 ) ;
 assign n741 = ( n635  &  n636 ) | ( n690  &  n636 ) | ( n635  &  n691 ) | ( n690  &  n691 ) ;
 assign n742 = ( n642  &  n643 ) | ( n693  &  n643 ) | ( n642  &  n694 ) | ( n693  &  n694 ) ;
 assign n743 = ( n741  &  n742 ) ;
 assign n745 = ( n743  &  n740 ) | ( n3719  &  n740 ) | ( n743  &  n288 ) | ( n3719  &  n288 ) ;
 assign n744 = ( n700  &  n745  &  n628 ) | ( n700  &  n745  &  n233 ) ;
 assign n746 = ( n236  &  n744  &  n18 ) | ( n236  &  n744  &  n740 ) ;
 assign n747 = ( n301  &  (~ n735) ) ;
 assign n749 = ( (~ Pi22)  &  n747 ) | ( (~ Pi22)  &  n304  &  (~ n742) ) ;
 assign n751 = ( n301  &  (~ n715) ) ;
 assign n752 = ( (~ Pi22)  &  n751 ) | ( (~ Pi22)  &  n304  &  (~ n725) ) ;
 assign n754 = ( Pi19  &  n310 ) | ( Pi19  &  n732 ) | ( n310  &  (~ n3769) ) | ( n732  &  (~ n3769) ) ;
 assign n756 = ( n739  &  n746 ) | ( n3776  &  n746 ) | ( n739  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n757 = ( n722 ) | ( n891 ) ;
 assign n753 = ( n754  &  n756  &  n757  &  (~ n3633) ) ;
 assign n759 = ( (~ n295) ) | ( n557 ) | ( n3626 ) | ( n3627 ) ;
 assign n758 = ( n759  &  (~ n3742) ) | ( (~ n3742)  &  (~ n4001) ) | ( (~ n3742)  &  (~ n4002) ) ;
 assign n764 = ( (~ n295) ) | ( n709 ) | ( n3628 ) | ( n3629 ) ;
 assign n763 = ( n764  &  (~ n3754) ) | ( (~ n3754)  &  (~ n4004) ) | ( (~ n3754)  &  (~ n4005) ) ;
 assign n769 = ( (~ n295) ) | ( n712 ) | ( n3750 ) | ( n3751 ) ;
 assign n768 = ( n769  &  (~ n1884) ) | ( (~ n1884)  &  (~ n3991) ) ;
 assign n774 = ( n18  &  n3576 ) | ( n18  &  (~ n3633)  &  n3994 ) ;
 assign n775 = ( n3582  &  n3998 ) | ( (~ n3769)  &  n3993  &  n3998 ) ;
 assign n776 = ( n3579  &  n3996 ) | ( (~ n3766)  &  n3990  &  n3996 ) ;
 assign n777 = ( n3995  &  n414 ) | ( n3995  &  n996 ) ;
 assign n773 = ( n774  &  n775  &  n776  &  n777 ) ;
 assign n779 = ( (~ n295) ) | ( n560 ) | ( n3736 ) | ( n3737 ) ;
 assign n778 = ( n779  &  (~ n1884) ) | ( (~ n1884)  &  (~ n3974) ) ;
 assign n782 = ( n18  &  n3576 ) | ( n18  &  (~ n3630)  &  n3981 ) ;
 assign n783 = ( n3582  &  n3985 ) | ( (~ n3759)  &  n3980  &  n3985 ) ;
 assign n784 = ( n3579  &  n3983 ) | ( (~ n3756)  &  n3969  &  n3983 ) ;
 assign n785 = ( n3982  &  n286 ) | ( n3982  &  n996 ) ;
 assign n781 = ( n782  &  n783  &  n784  &  n785 ) ;
 assign n788 = ( n4021  &  n626 ) | ( n4021  &  n1997 ) ;
 assign n787 = ( (~ Pi25) ) | ( n3729 ) ;
 assign n786 = ( n650  &  n788  &  (~ n3630) ) | ( n788  &  n787  &  (~ n3630) ) ;
 assign n791 = ( n4020  &  n581 ) | ( n4020  &  n1997 ) ;
 assign n789 = ( n602  &  n791  &  (~ n3759) ) | ( n787  &  n791  &  (~ n3759) ) ;
 assign n794 = ( n4019  &  n338 ) | ( n4019  &  n1997 ) ;
 assign n792 = ( n362  &  n794  &  (~ n3756) ) | ( n787  &  n794  &  (~ n3756) ) ;
 assign n797 = ( n792  &  n789 ) | ( n3735  &  n789 ) | ( n792  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n798 = ( n4014  &  n4022  &  n374 ) | ( n4014  &  n4022  &  n3716 ) ;
 assign n796 = ( (~ Pi19) ) | ( Pi17 ) ;
 assign n795 = ( n797  &  n798  &  n786 ) | ( n797  &  n798  &  n796 ) ;
 assign n801 = ( n4012  &  n529 ) | ( n4012  &  n1997 ) ;
 assign n799 = ( n554  &  (~ n759)  &  n801 ) | ( (~ n759)  &  n787  &  n801 ) ;
 assign n804 = ( n4011  &  n479 ) | ( n4011  &  n1997 ) ;
 assign n802 = ( n502  &  (~ n779)  &  n804 ) | ( (~ n779)  &  n787  &  n804 ) ;
 assign n807 = ( n4010  &  n235 ) | ( n4010  &  n1997 ) ;
 assign n805 = ( n267  &  n807  &  (~ n3732) ) | ( n787  &  n807  &  (~ n3732) ) ;
 assign n809 = ( n805  &  n802 ) | ( n3735  &  n802 ) | ( n805  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n810 = ( n4014  &  n4013  &  n286 ) | ( n4014  &  n4013  &  n3716 ) ;
 assign n808 = ( n809  &  n810  &  n799 ) | ( n809  &  n810  &  n796 ) ;
 assign n812 = ( n4025  &  n739 ) | ( n4025  &  n1997 ) ;
 assign n811 = ( n746  &  n812  &  (~ n3633) ) | ( n787  &  n812  &  (~ n3633) ) ;
 assign n815 = ( n4024  &  n722 ) | ( n4024  &  n1997 ) ;
 assign n813 = ( n732  &  n815  &  (~ n3769) ) | ( n787  &  n815  &  (~ n3769) ) ;
 assign n818 = ( n4023  &  n433 ) | ( n4023  &  n1997 ) ;
 assign n816 = ( n440  &  n818  &  (~ n3766) ) | ( n787  &  n818  &  (~ n3766) ) ;
 assign n820 = ( n816  &  n813 ) | ( n3735  &  n813 ) | ( n816  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n821 = ( n4014  &  n4026  &  n441 ) | ( n4014  &  n4026  &  n3716 ) ;
 assign n819 = ( n820  &  n821  &  n811 ) | ( n820  &  n821  &  n796 ) ;
 assign n824 = ( n4017  &  n698 ) | ( n4017  &  n1997 ) ;
 assign n822 = ( n706  &  (~ n764)  &  n824 ) | ( (~ n764)  &  n787  &  n824 ) ;
 assign n827 = ( n4016  &  n676 ) | ( n4016  &  n1997 ) ;
 assign n825 = ( n686  &  (~ n769)  &  n827 ) | ( (~ n769)  &  n787  &  n827 ) ;
 assign n830 = ( n4015  &  n404 ) | ( n4015  &  n1997 ) ;
 assign n828 = ( n413  &  n830  &  (~ n3746) ) | ( n787  &  n830  &  (~ n3746) ) ;
 assign n832 = ( n828  &  n825 ) | ( n3735  &  n825 ) | ( n828  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n833 = ( n4014  &  n4018  &  n414 ) | ( n4014  &  n4018  &  n3716 ) ;
 assign n831 = ( n832  &  n833  &  n822 ) | ( n832  &  n833  &  n796 ) ;
 assign n835 = ( n104  &  Ni42 ) ;
 assign n834 = ( (~ n200)  &  n390 ) | ( n390  &  n835 ) ;
 assign n837 = ( (~ Ni31) ) | ( (~ Ni30) ) ;
 assign n836 = ( (~ Ni30)  &  n837 ) | ( Ni33  &  n837 ) ;
 assign n841 = ( (~ n18) ) | ( (~ Ni30) ) ;
 assign n840 = ( (~ n70)  &  (~ Ni30) ) ;
 assign n839 = ( n841  &  n18 ) | ( n841  &  n840 ) ;
 assign n843 = ( (~ n74)  &  (~ Ni30) ) ;
 assign n842 = ( n841  &  n18 ) | ( n841  &  n843 ) ;
 assign n845 = ( (~ n78)  &  (~ Ni30) ) ;
 assign n844 = ( n841  &  n18 ) | ( n841  &  n845 ) ;
 assign n848 = ( n294  &  n297 ) ;
 assign n849 = ( n1054  &  n4055 ) | ( n1250  &  n4055 ) | ( n1054  &  n891 ) | ( n1250  &  n891 ) ;
 assign n847 = ( n1034  &  n842 ) ;
 assign n846 = ( n848  &  n849  &  n847 ) | ( n848  &  n849  &  n310 ) ;
 assign n851 = ( (~ n95)  &  (~ Ni30) ) ;
 assign n850 = ( n841  &  n18 ) | ( n841  &  n851 ) ;
 assign n853 = ( (~ n99)  &  (~ Ni30) ) ;
 assign n852 = ( n841  &  n18 ) | ( n841  &  n853 ) ;
 assign n855 = ( (~ n103)  &  (~ Ni30) ) ;
 assign n854 = ( n841  &  n18 ) | ( n841  &  n855 ) ;
 assign n858 = ( n1055  &  n4057 ) | ( n1250  &  n4057 ) | ( n1055  &  n891 ) | ( n1250  &  n891 ) ;
 assign n857 = ( n1052  &  n852 ) ;
 assign n856 = ( n848  &  n858  &  n857 ) | ( n848  &  n858  &  n310 ) ;
 assign n860 = ( (~ n115)  &  (~ Ni30) ) ;
 assign n859 = ( n841  &  n18 ) | ( n841  &  n860 ) ;
 assign n862 = ( (~ n117)  &  (~ Ni30) ) ;
 assign n861 = ( n841  &  n18 ) | ( n841  &  n862 ) ;
 assign n864 = ( (~ Ni30)  &  n952 ) ;
 assign n863 = ( n841  &  n18 ) | ( n841  &  n864 ) ;
 assign n867 = ( n995  &  n4069 ) | ( n1250  &  n4069 ) | ( n995  &  n891 ) | ( n1250  &  n891 ) ;
 assign n866 = ( n975  &  n861 ) ;
 assign n865 = ( n848  &  n867  &  n866 ) | ( n848  &  n867  &  n310 ) ;
 assign n869 = ( (~ n125)  &  (~ Ni30) ) ;
 assign n868 = ( n841  &  n18 ) | ( n841  &  n869 ) ;
 assign n871 = ( (~ n127)  &  (~ Ni30) ) ;
 assign n870 = ( n841  &  n18 ) | ( n841  &  n871 ) ;
 assign n873 = ( (~ Ni30)  &  n956 ) ;
 assign n872 = ( n841  &  n18 ) | ( n841  &  n873 ) ;
 assign n876 = ( n997  &  n4071 ) | ( n1250  &  n4071 ) | ( n997  &  n891 ) | ( n1250  &  n891 ) ;
 assign n875 = ( n993  &  n870 ) ;
 assign n874 = ( n848  &  n876  &  n875 ) | ( n848  &  n876  &  n310 ) ;
 assign n878 = ( (~ Ni37) ) | ( n390 ) ;
 assign n879 = ( n44 ) | ( n3723 ) ;
 assign n877 = ( n3846  &  n2937 ) ;
 assign n881 = ( (~ n51)  &  (~ Ni30) ) ;
 assign n880 = ( n841  &  n18 ) | ( n841  &  n881 ) ;
 assign n882 = ( n3848  &  n2937 ) ;
 assign n884 = ( (~ n58)  &  (~ Ni30) ) ;
 assign n883 = ( n841  &  n18 ) | ( n841  &  n884 ) ;
 assign n886 = ( (~ n61)  &  (~ Ni30) ) ;
 assign n885 = ( n841  &  n18 ) | ( n841  &  n886 ) ;
 assign n888 = ( (~ n66)  &  (~ Ni30) ) ;
 assign n887 = ( n841  &  n18 ) | ( n841  &  n888 ) ;
 assign n892 = ( n4061  &  n4062 ) | ( n3776  &  n4062 ) | ( n4061  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n893 = ( n848  &  n4059 ) | ( n848  &  n310 ) ;
 assign n890 = ( n1025  &  n880 ) ;
 assign n891 = ( Pi19 ) | ( n3727 ) ;
 assign n889 = ( n892  &  n893  &  n890 ) | ( n892  &  n893  &  n891 ) ;
 assign n895 = ( (~ n81)  &  (~ Ni30) ) ;
 assign n894 = ( n841  &  n18 ) | ( n841  &  n895 ) ;
 assign n897 = ( (~ n84)  &  (~ Ni30) ) ;
 assign n896 = ( n841  &  n18 ) | ( n841  &  n897 ) ;
 assign n899 = ( (~ n87)  &  (~ Ni30) ) ;
 assign n898 = ( n841  &  n18 ) | ( n841  &  n899 ) ;
 assign n901 = ( (~ n91)  &  (~ Ni30) ) ;
 assign n900 = ( n841  &  n18 ) | ( n841  &  n901 ) ;
 assign n904 = ( n4066  &  n4067 ) | ( n3776  &  n4067 ) | ( n4066  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n905 = ( n848  &  n4064 ) | ( n848  &  n310 ) ;
 assign n903 = ( n1043  &  n894 ) ;
 assign n902 = ( n904  &  n905  &  n903 ) | ( n904  &  n905  &  n891 ) ;
 assign n907 = ( (~ n106)  &  (~ Ni30) ) ;
 assign n906 = ( n841  &  n18 ) | ( n841  &  n907 ) ;
 assign n909 = ( (~ n109)  &  (~ Ni30) ) ;
 assign n908 = ( n841  &  n18 ) | ( n841  &  n909 ) ;
 assign n911 = ( (~ n110)  &  (~ Ni30) ) ;
 assign n910 = ( n841  &  n18 ) | ( n841  &  n911 ) ;
 assign n913 = ( (~ n113)  &  (~ Ni30) ) ;
 assign n912 = ( n841  &  n18 ) | ( n841  &  n913 ) ;
 assign n916 = ( n4075  &  n4076 ) | ( n3776  &  n4076 ) | ( n4075  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n917 = ( n848  &  n4073 ) | ( n848  &  n310 ) ;
 assign n915 = ( n966  &  n906 ) ;
 assign n914 = ( n916  &  n917  &  n915 ) | ( n916  &  n917  &  n891 ) ;
 assign n919 = ( (~ n119)  &  (~ Ni30) ) ;
 assign n918 = ( n841  &  n18 ) | ( n841  &  n919 ) ;
 assign n921 = ( (~ n120)  &  (~ Ni30) ) ;
 assign n920 = ( n841  &  n18 ) | ( n841  &  n921 ) ;
 assign n923 = ( (~ n121)  &  (~ Ni30) ) ;
 assign n922 = ( n841  &  n18 ) | ( n841  &  n923 ) ;
 assign n925 = ( (~ n123)  &  (~ Ni30) ) ;
 assign n924 = ( n841  &  n18 ) | ( n841  &  n925 ) ;
 assign n928 = ( n4080  &  n4081 ) | ( n3776  &  n4081 ) | ( n4080  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n929 = ( n848  &  n4078 ) | ( n848  &  n310 ) ;
 assign n927 = ( n984  &  n918 ) ;
 assign n926 = ( n928  &  n929  &  n927 ) | ( n928  &  n929  &  n891 ) ;
 assign n931 = ( Ni12 ) | ( n2456 ) ;
 assign n933 = ( n948  &  n848 ) ;
 assign n934 = ( Ni12 ) | ( (~ n2456) ) ;
 assign n930 = ( n931  &  n933 ) | ( n931  &  n934 ) | ( n933  &  (~ n3888) ) | ( n934  &  (~ n3888) ) ;
 assign n935 = ( (~ n1087)  &  (~ n3525) ) | ( (~ n1564)  &  (~ n1866)  &  (~ n3525) ) ;
 assign n941 = ( (~ n935)  &  n2312 ) | ( (~ n935)  &  (~ n3804)  &  n4233 ) ;
 assign n940 = ( (~ Ni12) ) | ( (~ Ni13) ) ;
 assign n939 = ( n930  &  n941  &  n933 ) | ( n930  &  n941  &  n940 ) ;
 assign n943 = ( (~ Ni30)  &  n836 ) | ( n836  &  (~ n3603) ) ;
 assign n942 = ( n943 ) | ( Pi22  &  Pi21 ) ;
 assign n945 = ( n942 ) | ( n3499 ) ;
 assign n946 = ( n933  &  n1066 ) | ( n933  &  n1150 ) | ( n1066  &  (~ n3784) ) | ( n1150  &  (~ n3784) ) ;
 assign n944 = ( n945  &  n946  &  Ni11 ) | ( n945  &  n946  &  n939 ) ;
 assign n949 = ( n4832 ) | ( n1866 ) ;
 assign n950 = ( Pi24  &  (~ n166) ) | ( (~ n166)  &  n848 ) | ( Pi24  &  n953 ) | ( n848  &  n953 ) ;
 assign n948 = ( n1470 ) | ( n1866 ) ;
 assign n947 = ( n949  &  n950  &  Pi24 ) | ( n949  &  n950  &  n948 ) ;
 assign n953 = ( n837  &  n3640 ) ;
 assign n954 = ( n4819 ) | ( n952 ) ;
 assign n952 = ( (~ n80) ) | ( n1063 ) ;
 assign n951 = ( n953  &  n954  &  n18 ) | ( n953  &  n954  &  n952 ) ;
 assign n957 = ( n4819 ) | ( n956 ) ;
 assign n956 = ( (~ n105) ) | ( n1063 ) ;
 assign n955 = ( n953  &  n957  &  n18 ) | ( n953  &  n957  &  n956 ) ;
 assign n960 = ( (~ n110) ) | ( n4819 ) ;
 assign n958 = ( n18  &  n953  &  n960 ) | ( (~ n110)  &  n953  &  n960 ) ;
 assign n963 = ( (~ n113) ) | ( n4819 ) ;
 assign n961 = ( n18  &  n953  &  n963 ) | ( (~ n113)  &  n953  &  n963 ) ;
 assign n966 = ( (~ n106) ) | ( n4819 ) ;
 assign n964 = ( n18  &  n953  &  n966 ) | ( (~ n106)  &  n953  &  n966 ) ;
 assign n969 = ( (~ n109) ) | ( n4819 ) ;
 assign n967 = ( n18  &  n953  &  n969 ) | ( (~ n109)  &  n953  &  n969 ) ;
 assign n972 = ( (~ n115) ) | ( n4819 ) ;
 assign n970 = ( n18  &  n953  &  n972 ) | ( (~ n115)  &  n953  &  n972 ) ;
 assign n975 = ( (~ n117) ) | ( n4819 ) ;
 assign n973 = ( n18  &  n953  &  n975 ) | ( (~ n117)  &  n953  &  n975 ) ;
 assign n978 = ( (~ n121) ) | ( n4819 ) ;
 assign n976 = ( n18  &  n953  &  n978 ) | ( (~ n121)  &  n953  &  n978 ) ;
 assign n981 = ( (~ n123) ) | ( n4819 ) ;
 assign n979 = ( n18  &  n953  &  n981 ) | ( (~ n123)  &  n953  &  n981 ) ;
 assign n984 = ( (~ n119) ) | ( n4819 ) ;
 assign n982 = ( n18  &  n953  &  n984 ) | ( (~ n119)  &  n953  &  n984 ) ;
 assign n987 = ( (~ n120) ) | ( n4819 ) ;
 assign n985 = ( n18  &  n953  &  n987 ) | ( (~ n120)  &  n953  &  n987 ) ;
 assign n990 = ( (~ n125) ) | ( n4819 ) ;
 assign n988 = ( n18  &  n953  &  n990 ) | ( (~ n125)  &  n953  &  n990 ) ;
 assign n993 = ( (~ n127) ) | ( n4819 ) ;
 assign n991 = ( n18  &  n953  &  n993 ) | ( (~ n127)  &  n953  &  n993 ) ;
 assign n995 = ( n954  &  n863 ) ;
 assign n996 = ( Pi16 ) | ( n3716 ) ;
 assign n997 = ( n957  &  n872 ) ;
 assign n998 = ( (~ Pi16) ) | ( n3716 ) ;
 assign n994 = ( n995  &  n997 ) | ( n996  &  n997 ) | ( n995  &  n998 ) | ( n996  &  n998 ) ;
 assign n999 = ( (~ n3777)  &  (~ n4207) ) | ( (~ n3777)  &  (~ n4208) ) ;
 assign n1003 = ( (~ n1884)  &  (~ n4211) ) | ( (~ n1884)  &  (~ n4212) ) ;
 assign n1007 = ( n950  &  n3576 ) | ( n950  &  n4218  &  n4217 ) ;
 assign n1008 = ( n4221  &  n3582 ) | ( n4221  &  n4216  &  n4215 ) ;
 assign n1009 = ( (~ n999)  &  n3579 ) | ( (~ n999)  &  n4209  &  n4210 ) ;
 assign n1010 = ( n4219  &  Pi24 ) | ( n4219  &  n994 ) ;
 assign n1006 = ( n1007  &  n1008  &  n1009  &  n1010 ) ;
 assign n1013 = ( (~ n78) ) | ( n4819 ) ;
 assign n1011 = ( n18  &  n953  &  n1013 ) | ( (~ n78)  &  n953  &  n1013 ) ;
 assign n1016 = ( (~ n103) ) | ( n4819 ) ;
 assign n1014 = ( n18  &  n953  &  n1016 ) | ( (~ n103)  &  n953  &  n1016 ) ;
 assign n1019 = ( (~ n61) ) | ( n4819 ) ;
 assign n1017 = ( n18  &  n953  &  n1019 ) | ( (~ n61)  &  n953  &  n1019 ) ;
 assign n1022 = ( (~ n66) ) | ( n4819 ) ;
 assign n1020 = ( n18  &  n953  &  n1022 ) | ( (~ n66)  &  n953  &  n1022 ) ;
 assign n1025 = ( (~ n51) ) | ( n4819 ) ;
 assign n1023 = ( n18  &  n953  &  n1025 ) | ( (~ n51)  &  n953  &  n1025 ) ;
 assign n1028 = ( (~ n58) ) | ( n4819 ) ;
 assign n1026 = ( n18  &  n953  &  n1028 ) | ( (~ n58)  &  n953  &  n1028 ) ;
 assign n1031 = ( (~ n70) ) | ( n4819 ) ;
 assign n1029 = ( n18  &  n953  &  n1031 ) | ( (~ n70)  &  n953  &  n1031 ) ;
 assign n1034 = ( (~ n74) ) | ( n4819 ) ;
 assign n1032 = ( n18  &  n953  &  n1034 ) | ( (~ n74)  &  n953  &  n1034 ) ;
 assign n1037 = ( (~ n87) ) | ( n4819 ) ;
 assign n1035 = ( n18  &  n953  &  n1037 ) | ( (~ n87)  &  n953  &  n1037 ) ;
 assign n1040 = ( (~ n91) ) | ( n4819 ) ;
 assign n1038 = ( n18  &  n953  &  n1040 ) | ( (~ n91)  &  n953  &  n1040 ) ;
 assign n1043 = ( (~ n81) ) | ( n4819 ) ;
 assign n1041 = ( n18  &  n953  &  n1043 ) | ( (~ n81)  &  n953  &  n1043 ) ;
 assign n1046 = ( (~ n84) ) | ( n4819 ) ;
 assign n1044 = ( n18  &  n953  &  n1046 ) | ( (~ n84)  &  n953  &  n1046 ) ;
 assign n1049 = ( (~ n95) ) | ( n4819 ) ;
 assign n1047 = ( n18  &  n953  &  n1049 ) | ( (~ n95)  &  n953  &  n1049 ) ;
 assign n1052 = ( (~ n99) ) | ( n4819 ) ;
 assign n1050 = ( n18  &  n953  &  n1052 ) | ( (~ n99)  &  n953  &  n1052 ) ;
 assign n1054 = ( n1013  &  n844 ) ;
 assign n1055 = ( n1016  &  n854 ) ;
 assign n1053 = ( n1054  &  n1055 ) | ( n996  &  n1055 ) | ( n1054  &  n998 ) | ( n996  &  n998 ) ;
 assign n1056 = ( (~ n3777)  &  (~ n4187) ) | ( (~ n3777)  &  (~ n4188) ) ;
 assign n1059 = ( (~ n1884)  &  (~ n4191) ) | ( (~ n1884)  &  (~ n4192) ) ;
 assign n1063 = ( Ni32 ) | ( n2068 ) ;
 assign n1062 = ( (~ n834) ) | ( n1063 ) ;
 assign n1066 = ( n3639  &  Pi26 ) | ( n3639  &  n1470 ) ;
 assign n1069 = ( (~ Ni11) ) | ( (~ Ni12) ) ;
 assign n1068 = ( Ni12 ) | ( Ni11 ) ;
 assign n1067 = ( n1069  &  Ni14  &  (~ Ni13) ) | ( n1069  &  n1068  &  (~ Ni13) ) ;
 assign n1074 = ( Ni11  &  (~ Ni12) ) ;
 assign n1071 = ( (~ n947)  &  (~ n1066)  &  n1074 ) | ( (~ n947)  &  (~ Ni14)  &  n1074 ) ;
 assign n1075 = ( Ni14  &  (~ n3814)  &  (~ n4675) ) | ( (~ n3814)  &  (~ n3891)  &  (~ n4675) ) ;
 assign n1079 = ( (~ n3831)  &  (~ n4202) ) | ( (~ n3831)  &  (~ n4205) ) | ( (~ n3831)  &  (~ n4206) ) ;
 assign n1084 = ( (~ n160)  &  (~ n164)  &  n949 ) | ( (~ n164)  &  n949  &  n948 ) ;
 assign n1088 = ( Pi21 ) | ( n3649 ) ;
 assign n1089 = ( Pi22 ) | ( n3649 ) ;
 assign n1087 = ( n1088  &  n1089 ) ;
 assign n1090 = ( Ni14  &  (~ Ni13) ) | ( Ni12  &  (~ Ni13) ) ;
 assign n1093 = ( (~ n164)  &  n1035 ) | ( (~ n164)  &  n3822 ) ;
 assign n1094 = ( n4066  &  n4067 ) | ( n3823  &  n4067 ) | ( n4066  &  n2411 ) | ( n3823  &  n2411 ) ;
 assign n1092 = ( n3729 ) | ( n160 ) ;
 assign n1091 = ( n1093  &  n1094  &  n1038 ) | ( n1093  &  n1094  &  n1092 ) ;
 assign n1096 = ( (~ n164)  &  n1041 ) | ( (~ n164)  &  n3822 ) ;
 assign n1097 = ( n903  &  n4064 ) | ( n3823  &  n4064 ) | ( n903  &  n2411 ) | ( n3823  &  n2411 ) ;
 assign n1095 = ( n1096  &  n1097  &  n1044 ) | ( n1096  &  n1097  &  n1092 ) ;
 assign n1099 = ( (~ n164)  &  n1047 ) | ( (~ n164)  &  n3822 ) ;
 assign n1100 = ( n4057  &  n857 ) | ( n3823  &  n857 ) | ( n4057  &  n2411 ) | ( n3823  &  n2411 ) ;
 assign n1098 = ( n1099  &  n1100  &  n1050 ) | ( n1099  &  n1100  &  n1092 ) ;
 assign n1102 = ( n1098  &  n1095 ) | ( n3735  &  n1095 ) | ( n1098  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1103 = ( n4181  &  n4179  &  n1055 ) | ( n4181  &  n4179  &  n3821 ) ;
 assign n1101 = ( n1102  &  n1103  &  n1091 ) | ( n1102  &  n1103  &  n796 ) ;
 assign n1105 = ( (~ n164)  &  n1017 ) | ( (~ n164)  &  n3822 ) ;
 assign n1106 = ( n4061  &  n4062 ) | ( n3823  &  n4062 ) | ( n4061  &  n2411 ) | ( n3823  &  n2411 ) ;
 assign n1104 = ( n1105  &  n1106  &  n1020 ) | ( n1105  &  n1106  &  n1092 ) ;
 assign n1108 = ( (~ n164)  &  n1023 ) | ( (~ n164)  &  n3822 ) ;
 assign n1109 = ( n890  &  n4059 ) | ( n3823  &  n4059 ) | ( n890  &  n2411 ) | ( n3823  &  n2411 ) ;
 assign n1107 = ( n1108  &  n1109  &  n1026 ) | ( n1108  &  n1109  &  n1092 ) ;
 assign n1111 = ( (~ n164)  &  n1029 ) | ( (~ n164)  &  n3822 ) ;
 assign n1112 = ( n4055  &  n847 ) | ( n3823  &  n847 ) | ( n4055  &  n2411 ) | ( n3823  &  n2411 ) ;
 assign n1110 = ( n1111  &  n1112  &  n1032 ) | ( n1111  &  n1112  &  n1092 ) ;
 assign n1114 = ( n1110  &  n1107 ) | ( n3735  &  n1107 ) | ( n1110  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1115 = ( n4178  &  n4179  &  n1054 ) | ( n4178  &  n4179  &  n3821 ) ;
 assign n1113 = ( n1114  &  n1115  &  n1104 ) | ( n1114  &  n1115  &  n796 ) ;
 assign n1117 = ( (~ n164)  &  n976 ) | ( (~ n164)  &  n3822 ) ;
 assign n1118 = ( n4080  &  n4081 ) | ( n3823  &  n4081 ) | ( n4080  &  n2411 ) | ( n3823  &  n2411 ) ;
 assign n1116 = ( n1117  &  n1118  &  n979 ) | ( n1117  &  n1118  &  n1092 ) ;
 assign n1120 = ( (~ n164)  &  n982 ) | ( (~ n164)  &  n3822 ) ;
 assign n1121 = ( n927  &  n4078 ) | ( n3823  &  n4078 ) | ( n927  &  n2411 ) | ( n3823  &  n2411 ) ;
 assign n1119 = ( n1120  &  n1121  &  n985 ) | ( n1120  &  n1121  &  n1092 ) ;
 assign n1123 = ( (~ n164)  &  n988 ) | ( (~ n164)  &  n3822 ) ;
 assign n1124 = ( n4071  &  n875 ) | ( n3823  &  n875 ) | ( n4071  &  n2411 ) | ( n3823  &  n2411 ) ;
 assign n1122 = ( n1123  &  n1124  &  n991 ) | ( n1123  &  n1124  &  n1092 ) ;
 assign n1126 = ( n1122  &  n1119 ) | ( n3735  &  n1119 ) | ( n1122  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1127 = ( n4182  &  n4179  &  n997 ) | ( n4182  &  n4179  &  n3821 ) ;
 assign n1125 = ( n1126  &  n1127  &  n1116 ) | ( n1126  &  n1127  &  n796 ) ;
 assign n1129 = ( (~ n164)  &  n958 ) | ( (~ n164)  &  n3822 ) ;
 assign n1130 = ( n4075  &  n4076 ) | ( n3823  &  n4076 ) | ( n4075  &  n2411 ) | ( n3823  &  n2411 ) ;
 assign n1128 = ( n1129  &  n1130  &  n961 ) | ( n1129  &  n1130  &  n1092 ) ;
 assign n1132 = ( (~ n164)  &  n964 ) | ( (~ n164)  &  n3822 ) ;
 assign n1133 = ( n915  &  n4073 ) | ( n3823  &  n4073 ) | ( n915  &  n2411 ) | ( n3823  &  n2411 ) ;
 assign n1131 = ( n1132  &  n1133  &  n967 ) | ( n1132  &  n1133  &  n1092 ) ;
 assign n1135 = ( (~ n164)  &  n970 ) | ( (~ n164)  &  n3822 ) ;
 assign n1136 = ( n4069  &  n866 ) | ( n3823  &  n866 ) | ( n4069  &  n2411 ) | ( n3823  &  n2411 ) ;
 assign n1134 = ( n1135  &  n1136  &  n973 ) | ( n1135  &  n1136  &  n1092 ) ;
 assign n1138 = ( n1134  &  n1131 ) | ( n3735  &  n1131 ) | ( n1134  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1139 = ( n4180  &  n4179  &  n995 ) | ( n4180  &  n4179  &  n3821 ) ;
 assign n1137 = ( n1138  &  n1139  &  n1128 ) | ( n1138  &  n1139  &  n796 ) ;
 assign n1141 = ( n160  &  (~ Ni14)  &  (~ n3641) ) | ( (~ Ni14)  &  (~ n3641)  &  (~ n3643) ) ;
 assign n1142 = ( n160  &  Ni14  &  (~ n1564)  &  (~ n1866) ) ;
 assign n1140 = ( Ni12  &  n1141 ) | ( Ni12  &  n1142 ) | ( Ni12  &  (~ n4176) ) ;
 assign n1145 = ( n931  &  (~ n1140) ) | ( (~ n1140)  &  n4183  &  n4184 ) ;
 assign n1144 = ( n1145  &  n1084 ) | ( n1145  &  n1090 ) ;
 assign n1146 = ( n160  &  (~ n943)  &  (~ n3499) ) | ( (~ n943)  &  (~ n953)  &  (~ n3499) ) ;
 assign n1152 = ( Ni11  &  n1084 ) | ( n1084  &  n1144 ) | ( Ni11  &  (~ n3784) ) | ( n1144  &  (~ n3784) ) ;
 assign n1150 = ( n1866 ) | ( n3499 ) ;
 assign n1149 = ( n1062  &  (~ n1146)  &  n1152 ) | ( (~ n1146)  &  n1152  &  n1150 ) ;
 assign n1153 = ( (~ n168)  &  (~ n167)  &  n949 ) | ( (~ n167)  &  n949  &  n948 ) ;
 assign n1158 = ( (~ n167)  &  n1035 ) | ( (~ n167)  &  n3834 ) ;
 assign n1159 = ( n4066  &  n4067 ) | ( n3835  &  n4067 ) | ( n4066  &  n2466 ) | ( n3835  &  n2466 ) ;
 assign n1157 = ( n3729 ) | ( n168 ) ;
 assign n1156 = ( n1158  &  n1159  &  n1038 ) | ( n1158  &  n1159  &  n1157 ) ;
 assign n1161 = ( (~ n167)  &  n1041 ) | ( (~ n167)  &  n3834 ) ;
 assign n1162 = ( n903  &  n4064 ) | ( n3835  &  n4064 ) | ( n903  &  n2466 ) | ( n3835  &  n2466 ) ;
 assign n1160 = ( n1161  &  n1162  &  n1044 ) | ( n1161  &  n1162  &  n1157 ) ;
 assign n1164 = ( (~ n167)  &  n1047 ) | ( (~ n167)  &  n3834 ) ;
 assign n1165 = ( n4057  &  n857 ) | ( n3835  &  n857 ) | ( n4057  &  n2466 ) | ( n3835  &  n2466 ) ;
 assign n1163 = ( n1164  &  n1165  &  n1050 ) | ( n1164  &  n1165  &  n1157 ) ;
 assign n1167 = ( n1163  &  n1160 ) | ( n3735  &  n1160 ) | ( n1163  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1168 = ( n4228  &  n4226  &  n1055 ) | ( n4228  &  n4226  &  n3833 ) ;
 assign n1166 = ( n1167  &  n1168  &  n1156 ) | ( n1167  &  n1168  &  n796 ) ;
 assign n1170 = ( (~ n167)  &  n1017 ) | ( (~ n167)  &  n3834 ) ;
 assign n1171 = ( n4061  &  n4062 ) | ( n3835  &  n4062 ) | ( n4061  &  n2466 ) | ( n3835  &  n2466 ) ;
 assign n1169 = ( n1170  &  n1171  &  n1020 ) | ( n1170  &  n1171  &  n1157 ) ;
 assign n1173 = ( (~ n167)  &  n1023 ) | ( (~ n167)  &  n3834 ) ;
 assign n1174 = ( n890  &  n4059 ) | ( n3835  &  n4059 ) | ( n890  &  n2466 ) | ( n3835  &  n2466 ) ;
 assign n1172 = ( n1173  &  n1174  &  n1026 ) | ( n1173  &  n1174  &  n1157 ) ;
 assign n1176 = ( (~ n167)  &  n1029 ) | ( (~ n167)  &  n3834 ) ;
 assign n1177 = ( n4055  &  n847 ) | ( n3835  &  n847 ) | ( n4055  &  n2466 ) | ( n3835  &  n2466 ) ;
 assign n1175 = ( n1176  &  n1177  &  n1032 ) | ( n1176  &  n1177  &  n1157 ) ;
 assign n1179 = ( n1175  &  n1172 ) | ( n3735  &  n1172 ) | ( n1175  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1180 = ( n4225  &  n4226  &  n1054 ) | ( n4225  &  n4226  &  n3833 ) ;
 assign n1178 = ( n1179  &  n1180  &  n1169 ) | ( n1179  &  n1180  &  n796 ) ;
 assign n1182 = ( (~ n167)  &  n976 ) | ( (~ n167)  &  n3834 ) ;
 assign n1183 = ( n4080  &  n4081 ) | ( n3835  &  n4081 ) | ( n4080  &  n2466 ) | ( n3835  &  n2466 ) ;
 assign n1181 = ( n1182  &  n1183  &  n979 ) | ( n1182  &  n1183  &  n1157 ) ;
 assign n1185 = ( (~ n167)  &  n982 ) | ( (~ n167)  &  n3834 ) ;
 assign n1186 = ( n927  &  n4078 ) | ( n3835  &  n4078 ) | ( n927  &  n2466 ) | ( n3835  &  n2466 ) ;
 assign n1184 = ( n1185  &  n1186  &  n985 ) | ( n1185  &  n1186  &  n1157 ) ;
 assign n1188 = ( (~ n167)  &  n988 ) | ( (~ n167)  &  n3834 ) ;
 assign n1189 = ( n4071  &  n875 ) | ( n3835  &  n875 ) | ( n4071  &  n2466 ) | ( n3835  &  n2466 ) ;
 assign n1187 = ( n1188  &  n1189  &  n991 ) | ( n1188  &  n1189  &  n1157 ) ;
 assign n1191 = ( n1187  &  n1184 ) | ( n3735  &  n1184 ) | ( n1187  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1192 = ( n4229  &  n4226  &  n997 ) | ( n4229  &  n4226  &  n3833 ) ;
 assign n1190 = ( n1191  &  n1192  &  n1181 ) | ( n1191  &  n1192  &  n796 ) ;
 assign n1194 = ( (~ n167)  &  n958 ) | ( (~ n167)  &  n3834 ) ;
 assign n1195 = ( n4075  &  n4076 ) | ( n3835  &  n4076 ) | ( n4075  &  n2466 ) | ( n3835  &  n2466 ) ;
 assign n1193 = ( n1194  &  n1195  &  n961 ) | ( n1194  &  n1195  &  n1157 ) ;
 assign n1197 = ( (~ n167)  &  n964 ) | ( (~ n167)  &  n3834 ) ;
 assign n1198 = ( n915  &  n4073 ) | ( n3835  &  n4073 ) | ( n915  &  n2466 ) | ( n3835  &  n2466 ) ;
 assign n1196 = ( n1197  &  n1198  &  n967 ) | ( n1197  &  n1198  &  n1157 ) ;
 assign n1200 = ( (~ n167)  &  n970 ) | ( (~ n167)  &  n3834 ) ;
 assign n1201 = ( n4069  &  n866 ) | ( n3835  &  n866 ) | ( n4069  &  n2466 ) | ( n3835  &  n2466 ) ;
 assign n1199 = ( n1200  &  n1201  &  n973 ) | ( n1200  &  n1201  &  n1157 ) ;
 assign n1203 = ( n1199  &  n1196 ) | ( n3735  &  n1196 ) | ( n1199  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1204 = ( n4227  &  n4226  &  n995 ) | ( n4227  &  n4226  &  n3833 ) ;
 assign n1202 = ( n1203  &  n1204  &  n1193 ) | ( n1203  &  n1204  &  n796 ) ;
 assign n1206 = ( n168  &  (~ Ni14)  &  (~ n3641) ) | ( (~ Ni14)  &  (~ n3641)  &  (~ n3643) ) ;
 assign n1207 = ( n168  &  Ni14  &  (~ n1564)  &  (~ n1866) ) ;
 assign n1205 = ( Ni12  &  n1206 ) | ( Ni12  &  n1207 ) | ( Ni12  &  (~ n4224) ) ;
 assign n1210 = ( n931  &  (~ n1205) ) | ( (~ n1205)  &  n4230  &  n4231 ) ;
 assign n1209 = ( n1210  &  n1090 ) | ( n1210  &  n1153 ) ;
 assign n1211 = ( n168  &  (~ n943)  &  (~ n3499) ) | ( (~ n943)  &  (~ n953)  &  (~ n3499) ) ;
 assign n1214 = ( Ni11  &  n1153 ) | ( n1153  &  n1209 ) | ( Ni11  &  (~ n3784) ) | ( n1209  &  (~ n3784) ) ;
 assign n1212 = ( n1062  &  (~ n1211)  &  n1214 ) | ( n1150  &  (~ n1211)  &  n1214 ) ;
 assign n1215 = ( (~ Ni8)  &  (~ Ni9) ) | ( (~ Ni9)  &  (~ Ni7) ) ;
 assign n1218 = ( n1215  &  Ni10 ) | ( n1215  &  (~ Ni7) ) ;
 assign n1221 = ( n4047  &  n1329 ) | ( n1250  &  n1329 ) | ( n4047  &  n891 ) | ( n1250  &  n891 ) ;
 assign n1220 = ( n1327  &  n842 ) ;
 assign n1219 = ( n848  &  n1221  &  n1220 ) | ( n848  &  n1221  &  n310 ) ;
 assign n1224 = ( n4049  &  n1294 ) | ( n1250  &  n1294 ) | ( n4049  &  n891 ) | ( n1250  &  n891 ) ;
 assign n1223 = ( n1292  &  n852 ) ;
 assign n1222 = ( n848  &  n1224  &  n1223 ) | ( n848  &  n1224  &  n310 ) ;
 assign n1227 = ( n4048  &  n1399 ) | ( n1250  &  n1399 ) | ( n4048  &  n891 ) | ( n1250  &  n891 ) ;
 assign n1226 = ( n1397  &  n861 ) ;
 assign n1225 = ( n848  &  n1227  &  n1226 ) | ( n848  &  n1227  &  n310 ) ;
 assign n1230 = ( n4050  &  n1364 ) | ( n1250  &  n1364 ) | ( n4050  &  n891 ) | ( n1250  &  n891 ) ;
 assign n1229 = ( n1362  &  n870 ) ;
 assign n1228 = ( n848  &  n1230  &  n1229 ) | ( n848  &  n1230  &  n310 ) ;
 assign n1233 = ( n1310  &  n4037 ) | ( n3776  &  n4037 ) | ( n1310  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n1234 = ( n848  &  n4038 ) | ( n848  &  n310 ) ;
 assign n1232 = ( n1315  &  n880 ) ;
 assign n1231 = ( n1233  &  n1234  &  n1232 ) | ( n1233  &  n1234  &  n891 ) ;
 assign n1237 = ( n1274  &  n4041 ) | ( n3776  &  n4041 ) | ( n1274  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n1238 = ( n848  &  n4042 ) | ( n848  &  n310 ) ;
 assign n1236 = ( n1280  &  n894 ) ;
 assign n1235 = ( n1237  &  n1238  &  n1236 ) | ( n1237  &  n1238  &  n891 ) ;
 assign n1241 = ( n1380  &  n4039 ) | ( n3776  &  n4039 ) | ( n1380  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n1242 = ( n848  &  n4040 ) | ( n848  &  n310 ) ;
 assign n1240 = ( n1385  &  n906 ) ;
 assign n1239 = ( n1241  &  n1242  &  n1240 ) | ( n1241  &  n1242  &  n891 ) ;
 assign n1245 = ( n1345  &  n4043 ) | ( n3776  &  n4043 ) | ( n1345  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n1246 = ( n848  &  n4044 ) | ( n848  &  n310 ) ;
 assign n1244 = ( n1350  &  n918 ) ;
 assign n1243 = ( n1245  &  n1246  &  n1244 ) | ( n1245  &  n1246  &  n891 ) ;
 assign n1248 = ( (~ Pi20)  &  n851 ) | ( Pi20  &  n853 ) | ( n851  &  n853 ) ;
 assign n1249 = ( Pi19 ) | ( n1866 ) ;
 assign n1250 = ( (~ Pi19) ) | ( n1866 ) ;
 assign n1247 = ( n1248  &  n855 ) | ( n1249  &  n855 ) | ( n1248  &  n1250 ) | ( n1249  &  n1250 ) ;
 assign n1252 = ( (~ Pi20)  &  n860 ) | ( Pi20  &  n862 ) | ( n860  &  n862 ) ;
 assign n1251 = ( n1252  &  n864 ) | ( n1249  &  n864 ) | ( n1252  &  n1250 ) | ( n1249  &  n1250 ) ;
 assign n1254 = ( (~ Pi20)  &  n869 ) | ( Pi20  &  n871 ) | ( n869  &  n871 ) ;
 assign n1253 = ( n1254  &  n873 ) | ( n1249  &  n873 ) | ( n1254  &  n1250 ) | ( n1249  &  n1250 ) ;
 assign n1256 = ( (~ Pi20)  &  n895 ) | ( Pi20  &  n897 ) | ( n895  &  n897 ) ;
 assign n1257 = ( (~ Pi20)  &  n899 ) | ( Pi20  &  n901 ) | ( n899  &  n901 ) ;
 assign n1255 = ( n1256  &  n1257 ) | ( n1249  &  n1257 ) | ( n1256  &  n1250 ) | ( n1249  &  n1250 ) ;
 assign n1259 = ( (~ Pi20)  &  n907 ) | ( Pi20  &  n909 ) | ( n907  &  n909 ) ;
 assign n1260 = ( (~ Pi20)  &  n911 ) | ( Pi20  &  n913 ) | ( n911  &  n913 ) ;
 assign n1258 = ( n1259  &  n1260 ) | ( n1249  &  n1260 ) | ( n1259  &  n1250 ) | ( n1249  &  n1250 ) ;
 assign n1262 = ( (~ Pi20)  &  n919 ) | ( Pi20  &  n921 ) | ( n919  &  n921 ) ;
 assign n1263 = ( (~ Pi20)  &  n923 ) | ( Pi20  &  n925 ) | ( n923  &  n925 ) ;
 assign n1261 = ( n1262  &  n1263 ) | ( n1249  &  n1263 ) | ( n1262  &  n1250 ) | ( n1249  &  n1250 ) ;
 assign n1266 = ( n4691 ) | ( n4692 ) | ( n931 ) ;
 assign n1265 = ( Pi17  &  (~ n4689) ) | ( n4045  &  n4046  &  (~ n4689) ) ;
 assign n1264 = ( n1266  &  n1265 ) | ( n1266  &  n934 ) ;
 assign n1269 = ( (~ n87) ) | ( n4820 ) ;
 assign n1268 = ( (~ n87)  &  n836 ) ;
 assign n1267 = ( n836  &  n1269  &  n18 ) | ( n836  &  n1269  &  n1268 ) ;
 assign n1272 = ( (~ n91) ) | ( n4820 ) ;
 assign n1271 = ( (~ n91)  &  n836 ) ;
 assign n1270 = ( n836  &  n1272  &  n18 ) | ( n836  &  n1272  &  n1271 ) ;
 assign n1276 = ( n1267  &  n1270 ) | ( n3801  &  n1270 ) | ( n1267  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n1277 = ( n3803  &  (~ n3804) ) | ( (~ n3804)  &  n4041 ) ;
 assign n1274 = ( n1269  &  n898 ) ;
 assign n1275 = ( (~ n161) ) | ( n3727 ) ;
 assign n1273 = ( n1276  &  n1277  &  n1274 ) | ( n1276  &  n1277  &  n1275 ) ;
 assign n1280 = ( (~ n81) ) | ( n4820 ) ;
 assign n1279 = ( (~ n81)  &  n836 ) ;
 assign n1278 = ( n836  &  n1280  &  n18 ) | ( n836  &  n1280  &  n1279 ) ;
 assign n1283 = ( (~ n84) ) | ( n4820 ) ;
 assign n1282 = ( (~ n84)  &  n836 ) ;
 assign n1281 = ( n836  &  n1283  &  n18 ) | ( n836  &  n1283  &  n1282 ) ;
 assign n1285 = ( n1278  &  n1281 ) | ( n3801  &  n1281 ) | ( n1278  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n1286 = ( n3803  &  (~ n3804) ) | ( (~ n3804)  &  n4042 ) ;
 assign n1284 = ( n1285  &  n1286  &  n1236 ) | ( n1285  &  n1286  &  n1275 ) ;
 assign n1289 = ( (~ n95) ) | ( n4820 ) ;
 assign n1288 = ( (~ n95)  &  n836 ) ;
 assign n1287 = ( n836  &  n1289  &  n18 ) | ( n836  &  n1289  &  n1288 ) ;
 assign n1292 = ( (~ n99) ) | ( n4820 ) ;
 assign n1291 = ( (~ n99)  &  n836 ) ;
 assign n1290 = ( n836  &  n1292  &  n18 ) | ( n836  &  n1292  &  n1291 ) ;
 assign n1295 = ( n1287  &  n1290 ) | ( n3801  &  n1290 ) | ( n1287  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n1296 = ( n1223  &  (~ n3804) ) | ( n3803  &  (~ n3804) ) ;
 assign n1294 = ( n1289  &  n850 ) ;
 assign n1293 = ( n1295  &  n1296  &  n1294 ) | ( n1295  &  n1296  &  n1275 ) ;
 assign n1299 = ( (~ n103) ) | ( n4820 ) ;
 assign n1298 = ( (~ n103)  &  n836 ) ;
 assign n1297 = ( n836  &  n1299  &  n18 ) | ( n836  &  n1299  &  n1298 ) ;
 assign n1301 = ( n1293  &  n1284 ) | ( n3735  &  n1284 ) | ( n1293  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1302 = ( n4170  &  n4168  &  n4049 ) | ( n4170  &  n4168  &  n3800 ) ;
 assign n1300 = ( n1301  &  n1302  &  n1273 ) | ( n1301  &  n1302  &  n796 ) ;
 assign n1305 = ( (~ n61) ) | ( n4820 ) ;
 assign n1304 = ( (~ n61)  &  n836 ) ;
 assign n1303 = ( n836  &  n1305  &  n18 ) | ( n836  &  n1305  &  n1304 ) ;
 assign n1308 = ( (~ n66) ) | ( n4820 ) ;
 assign n1307 = ( (~ n66)  &  n836 ) ;
 assign n1306 = ( n836  &  n1308  &  n18 ) | ( n836  &  n1308  &  n1307 ) ;
 assign n1311 = ( n1303  &  n1306 ) | ( n3801  &  n1306 ) | ( n1303  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n1312 = ( n3803  &  (~ n3804) ) | ( (~ n3804)  &  n4037 ) ;
 assign n1310 = ( n1305  &  n885 ) ;
 assign n1309 = ( n1311  &  n1312  &  n1310 ) | ( n1311  &  n1312  &  n1275 ) ;
 assign n1315 = ( (~ n51) ) | ( n4820 ) ;
 assign n1314 = ( (~ n51)  &  n836 ) ;
 assign n1313 = ( n836  &  n1315  &  n18 ) | ( n836  &  n1315  &  n1314 ) ;
 assign n1318 = ( (~ n58) ) | ( n4820 ) ;
 assign n1317 = ( (~ n58)  &  n836 ) ;
 assign n1316 = ( n836  &  n1318  &  n18 ) | ( n836  &  n1318  &  n1317 ) ;
 assign n1320 = ( n1313  &  n1316 ) | ( n3801  &  n1316 ) | ( n1313  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n1321 = ( n3803  &  (~ n3804) ) | ( (~ n3804)  &  n4038 ) ;
 assign n1319 = ( n1320  &  n1321  &  n1232 ) | ( n1320  &  n1321  &  n1275 ) ;
 assign n1324 = ( (~ n70) ) | ( n4820 ) ;
 assign n1323 = ( (~ n70)  &  n836 ) ;
 assign n1322 = ( n18  &  n836  &  n1324 ) | ( n836  &  n1324  &  n1323 ) ;
 assign n1327 = ( (~ n74) ) | ( n4820 ) ;
 assign n1326 = ( (~ n74)  &  n836 ) ;
 assign n1325 = ( n18  &  n836  &  n1327 ) | ( n836  &  n1327  &  n1326 ) ;
 assign n1330 = ( n1322  &  n1325 ) | ( n3801  &  n1325 ) | ( n1322  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n1331 = ( n1220  &  (~ n3804) ) | ( n3803  &  (~ n3804) ) ;
 assign n1329 = ( n1324  &  n839 ) ;
 assign n1328 = ( n1330  &  n1331  &  n1329 ) | ( n1330  &  n1331  &  n1275 ) ;
 assign n1334 = ( (~ n78) ) | ( n4820 ) ;
 assign n1333 = ( (~ n78)  &  n836 ) ;
 assign n1332 = ( n18  &  n836  &  n1334 ) | ( n836  &  n1334  &  n1333 ) ;
 assign n1336 = ( n1328  &  n1319 ) | ( n3735  &  n1319 ) | ( n1328  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1337 = ( n4167  &  n4168  &  n4047 ) | ( n4167  &  n4168  &  n3800 ) ;
 assign n1335 = ( n1336  &  n1337  &  n1309 ) | ( n1336  &  n1337  &  n796 ) ;
 assign n1340 = ( (~ n121) ) | ( n4820 ) ;
 assign n1339 = ( (~ n121)  &  n836 ) ;
 assign n1338 = ( n18  &  n836  &  n1340 ) | ( n836  &  n1340  &  n1339 ) ;
 assign n1343 = ( (~ n123) ) | ( n4820 ) ;
 assign n1342 = ( (~ n123)  &  n836 ) ;
 assign n1341 = ( n18  &  n836  &  n1343 ) | ( n836  &  n1343  &  n1342 ) ;
 assign n1346 = ( n1338  &  n1341 ) | ( n3801  &  n1341 ) | ( n1338  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n1347 = ( n3803  &  (~ n3804) ) | ( (~ n3804)  &  n4043 ) ;
 assign n1345 = ( n1340  &  n922 ) ;
 assign n1344 = ( n1346  &  n1347  &  n1345 ) | ( n1346  &  n1347  &  n1275 ) ;
 assign n1350 = ( (~ n119) ) | ( n4820 ) ;
 assign n1349 = ( (~ n119)  &  n836 ) ;
 assign n1348 = ( n18  &  n836  &  n1350 ) | ( n836  &  n1350  &  n1349 ) ;
 assign n1353 = ( (~ n120) ) | ( n4820 ) ;
 assign n1352 = ( (~ n120)  &  n836 ) ;
 assign n1351 = ( n18  &  n836  &  n1353 ) | ( n836  &  n1353  &  n1352 ) ;
 assign n1355 = ( n1348  &  n1351 ) | ( n3801  &  n1351 ) | ( n1348  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n1356 = ( n3803  &  (~ n3804) ) | ( (~ n3804)  &  n4044 ) ;
 assign n1354 = ( n1355  &  n1356  &  n1244 ) | ( n1355  &  n1356  &  n1275 ) ;
 assign n1359 = ( (~ n125) ) | ( n4820 ) ;
 assign n1358 = ( (~ n125)  &  n836 ) ;
 assign n1357 = ( n18  &  n836  &  n1359 ) | ( n836  &  n1359  &  n1358 ) ;
 assign n1362 = ( (~ n127) ) | ( n4820 ) ;
 assign n1361 = ( (~ n127)  &  n836 ) ;
 assign n1360 = ( n18  &  n836  &  n1362 ) | ( n836  &  n1362  &  n1361 ) ;
 assign n1365 = ( n1357  &  n1360 ) | ( n3801  &  n1360 ) | ( n1357  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n1366 = ( n1229  &  (~ n3804) ) | ( n3803  &  (~ n3804) ) ;
 assign n1364 = ( n1359  &  n868 ) ;
 assign n1363 = ( n1365  &  n1366  &  n1364 ) | ( n1365  &  n1366  &  n1275 ) ;
 assign n1369 = ( n4820 ) | ( n956 ) ;
 assign n1368 = ( n956  &  n836 ) ;
 assign n1367 = ( n18  &  n836  &  n1369 ) | ( n836  &  n1369  &  n1368 ) ;
 assign n1371 = ( n1363  &  n1354 ) | ( n3735  &  n1354 ) | ( n1363  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1372 = ( n4171  &  n4168  &  n4050 ) | ( n4171  &  n4168  &  n3800 ) ;
 assign n1370 = ( n1371  &  n1372  &  n1344 ) | ( n1371  &  n1372  &  n796 ) ;
 assign n1375 = ( (~ n110) ) | ( n4820 ) ;
 assign n1374 = ( (~ n110)  &  n836 ) ;
 assign n1373 = ( n18  &  n836  &  n1375 ) | ( n836  &  n1375  &  n1374 ) ;
 assign n1378 = ( (~ n113) ) | ( n4820 ) ;
 assign n1377 = ( (~ n113)  &  n836 ) ;
 assign n1376 = ( n18  &  n836  &  n1378 ) | ( n836  &  n1378  &  n1377 ) ;
 assign n1381 = ( n1373  &  n1376 ) | ( n3801  &  n1376 ) | ( n1373  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n1382 = ( n3803  &  (~ n3804) ) | ( (~ n3804)  &  n4039 ) ;
 assign n1380 = ( n1375  &  n910 ) ;
 assign n1379 = ( n1381  &  n1382  &  n1380 ) | ( n1381  &  n1382  &  n1275 ) ;
 assign n1385 = ( (~ n106) ) | ( n4820 ) ;
 assign n1384 = ( (~ n106)  &  n836 ) ;
 assign n1383 = ( n18  &  n836  &  n1385 ) | ( n836  &  n1385  &  n1384 ) ;
 assign n1388 = ( (~ n109) ) | ( n4820 ) ;
 assign n1387 = ( (~ n109)  &  n836 ) ;
 assign n1386 = ( n18  &  n836  &  n1388 ) | ( n836  &  n1388  &  n1387 ) ;
 assign n1390 = ( n1383  &  n1386 ) | ( n3801  &  n1386 ) | ( n1383  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n1391 = ( n3803  &  (~ n3804) ) | ( (~ n3804)  &  n4040 ) ;
 assign n1389 = ( n1390  &  n1391  &  n1240 ) | ( n1390  &  n1391  &  n1275 ) ;
 assign n1394 = ( (~ n115) ) | ( n4820 ) ;
 assign n1393 = ( (~ n115)  &  n836 ) ;
 assign n1392 = ( n18  &  n836  &  n1394 ) | ( n836  &  n1394  &  n1393 ) ;
 assign n1397 = ( (~ n117) ) | ( n4820 ) ;
 assign n1396 = ( (~ n117)  &  n836 ) ;
 assign n1395 = ( n18  &  n836  &  n1397 ) | ( n836  &  n1397  &  n1396 ) ;
 assign n1400 = ( n1392  &  n1395 ) | ( n3801  &  n1395 ) | ( n1392  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n1401 = ( n1226  &  (~ n3804) ) | ( n3803  &  (~ n3804) ) ;
 assign n1399 = ( n1394  &  n859 ) ;
 assign n1398 = ( n1400  &  n1401  &  n1399 ) | ( n1400  &  n1401  &  n1275 ) ;
 assign n1404 = ( n4820 ) | ( n952 ) ;
 assign n1403 = ( n952  &  n836 ) ;
 assign n1402 = ( n18  &  n836  &  n1404 ) | ( n836  &  n1404  &  n1403 ) ;
 assign n1406 = ( n1398  &  n1389 ) | ( n3735  &  n1389 ) | ( n1398  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1407 = ( n4169  &  n4168  &  n4048 ) | ( n4169  &  n4168  &  n3800 ) ;
 assign n1405 = ( n1406  &  n1407  &  n1379 ) | ( n1406  &  n1407  &  n796 ) ;
 assign n1408 = ( (~ n1884)  &  (~ n4151) ) | ( (~ n1884)  &  (~ n4152) ) ;
 assign n1411 = ( (~ n1884)  &  (~ n4131) ) | ( (~ n1884)  &  (~ n4132) ) ;
 assign n1415 = ( n4685 ) | ( n4687 ) | ( n3525 ) ;
 assign n1416 = ( n1264  &  n2312 ) | ( n1264  &  n4173  &  n4172 ) ;
 assign n1414 = ( n1415  &  n1416  &  n1265 ) | ( n1415  &  n1416  &  n940 ) ;
 assign n1419 = ( n1267  &  n1270 ) | ( n3787  &  n1270 ) | ( n1267  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n1420 = ( n942  &  n4041 ) | ( n942  &  n3789 ) ;
 assign n1418 = ( (~ n3603) ) | ( n3727 ) ;
 assign n1417 = ( n1419  &  n1420  &  n1274 ) | ( n1419  &  n1420  &  n1418 ) ;
 assign n1422 = ( n1278  &  n1281 ) | ( n3787  &  n1281 ) | ( n1278  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n1423 = ( n942  &  n4042 ) | ( n942  &  n3789 ) ;
 assign n1421 = ( n1422  &  n1423  &  n1236 ) | ( n1422  &  n1423  &  n1418 ) ;
 assign n1425 = ( n1287  &  n1290 ) | ( n3787  &  n1290 ) | ( n1287  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n1426 = ( n942  &  n1223 ) | ( n942  &  n3789 ) ;
 assign n1424 = ( n1425  &  n1426  &  n1294 ) | ( n1425  &  n1426  &  n1418 ) ;
 assign n1428 = ( n1424  &  n1421 ) | ( n3735  &  n1421 ) | ( n1424  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1429 = ( n4125  &  n4123  &  n4049 ) | ( n4125  &  n4123  &  n3786 ) ;
 assign n1427 = ( n1428  &  n1429  &  n1417 ) | ( n1428  &  n1429  &  n796 ) ;
 assign n1431 = ( n1303  &  n1306 ) | ( n3787  &  n1306 ) | ( n1303  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n1432 = ( n942  &  n4037 ) | ( n942  &  n3789 ) ;
 assign n1430 = ( n1431  &  n1432  &  n1310 ) | ( n1431  &  n1432  &  n1418 ) ;
 assign n1434 = ( n1313  &  n1316 ) | ( n3787  &  n1316 ) | ( n1313  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n1435 = ( n942  &  n4038 ) | ( n942  &  n3789 ) ;
 assign n1433 = ( n1434  &  n1435  &  n1232 ) | ( n1434  &  n1435  &  n1418 ) ;
 assign n1437 = ( n1322  &  n1325 ) | ( n3787  &  n1325 ) | ( n1322  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n1438 = ( n942  &  n1220 ) | ( n942  &  n3789 ) ;
 assign n1436 = ( n1437  &  n1438  &  n1329 ) | ( n1437  &  n1438  &  n1418 ) ;
 assign n1440 = ( n1436  &  n1433 ) | ( n3735  &  n1433 ) | ( n1436  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1441 = ( n4122  &  n4123  &  n4047 ) | ( n4122  &  n4123  &  n3786 ) ;
 assign n1439 = ( n1440  &  n1441  &  n1430 ) | ( n1440  &  n1441  &  n796 ) ;
 assign n1443 = ( n1338  &  n1341 ) | ( n3787  &  n1341 ) | ( n1338  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n1444 = ( n942  &  n4043 ) | ( n942  &  n3789 ) ;
 assign n1442 = ( n1443  &  n1444  &  n1345 ) | ( n1443  &  n1444  &  n1418 ) ;
 assign n1446 = ( n1348  &  n1351 ) | ( n3787  &  n1351 ) | ( n1348  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n1447 = ( n942  &  n4044 ) | ( n942  &  n3789 ) ;
 assign n1445 = ( n1446  &  n1447  &  n1244 ) | ( n1446  &  n1447  &  n1418 ) ;
 assign n1449 = ( n1357  &  n1360 ) | ( n3787  &  n1360 ) | ( n1357  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n1450 = ( n942  &  n1229 ) | ( n942  &  n3789 ) ;
 assign n1448 = ( n1449  &  n1450  &  n1364 ) | ( n1449  &  n1450  &  n1418 ) ;
 assign n1452 = ( n1448  &  n1445 ) | ( n3735  &  n1445 ) | ( n1448  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1453 = ( n4126  &  n4123  &  n4050 ) | ( n4126  &  n4123  &  n3786 ) ;
 assign n1451 = ( n1452  &  n1453  &  n1442 ) | ( n1452  &  n1453  &  n796 ) ;
 assign n1455 = ( n1373  &  n1376 ) | ( n3787  &  n1376 ) | ( n1373  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n1456 = ( n942  &  n4039 ) | ( n942  &  n3789 ) ;
 assign n1454 = ( n1455  &  n1456  &  n1380 ) | ( n1455  &  n1456  &  n1418 ) ;
 assign n1458 = ( n1383  &  n1386 ) | ( n3787  &  n1386 ) | ( n1383  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n1459 = ( n942  &  n4040 ) | ( n942  &  n3789 ) ;
 assign n1457 = ( n1458  &  n1459  &  n1240 ) | ( n1458  &  n1459  &  n1418 ) ;
 assign n1461 = ( n1392  &  n1395 ) | ( n3787  &  n1395 ) | ( n1392  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n1462 = ( n942  &  n1226 ) | ( n942  &  n3789 ) ;
 assign n1460 = ( n1461  &  n1462  &  n1399 ) | ( n1461  &  n1462  &  n1418 ) ;
 assign n1464 = ( n1460  &  n1457 ) | ( n3735  &  n1457 ) | ( n1460  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1465 = ( n4124  &  n4123  &  n4048 ) | ( n4124  &  n4123  &  n3786 ) ;
 assign n1463 = ( n1464  &  n1465  &  n1454 ) | ( n1464  &  n1465  &  n796 ) ;
 assign n1467 = ( n1427  &  n1451 ) | ( n3763  &  n1451 ) | ( n1427  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n1468 = ( n1439  &  n1463 ) | ( n3742  &  n1463 ) | ( n1439  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n1466 = ( n1467  &  n1468 ) ;
 assign n1470 = ( (~ Ni30)  &  n1062 ) ;
 assign n1471 = ( Pi25 ) | ( n1866 ) ;
 assign n1469 = ( n848  &  n1470 ) | ( n848  &  n1471 ) ;
 assign n1475 = ( n1469  &  n1480 ) | ( n1469  &  n4036  &  n4034 ) ;
 assign n1473 = ( (~ Pi16)  &  n864 ) | ( n864  &  n873 ) ;
 assign n1474 = ( (~ Pi25) ) | ( n3716 ) ;
 assign n1472 = ( n1475  &  n1473 ) | ( n1475  &  n1474 ) ;
 assign n1478 = ( n1469  &  n1480 ) | ( n1469  &  n4032  &  n4030 ) ;
 assign n1477 = ( (~ Pi16)  &  n845 ) | ( n845  &  n855 ) ;
 assign n1476 = ( n1478  &  n1477 ) | ( n1478  &  n1474 ) ;
 assign n1481 = ( n4069  &  n866 ) | ( n3728  &  n866 ) | ( n4069  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n1480 = ( (~ Pi25) ) | ( n1866 ) ;
 assign n1479 = ( n1481  &  n1252 ) | ( n1481  &  n1480 ) ;
 assign n1482 = ( (~ n3579)  &  (~ n4070) ) | ( (~ n1254)  &  (~ n1480)  &  (~ n3579) ) ;
 assign n1487 = ( (~ n1884)  &  (~ n4072) ) | ( (~ n1259)  &  (~ n1480)  &  (~ n1884) ) ;
 assign n1490 = ( (~ n3778)  &  (~ n4074) ) | ( (~ n1260)  &  (~ n1480)  &  (~ n3778) ) ;
 assign n1494 = ( (~ n3582)  &  (~ n4077) ) | ( (~ n1262)  &  (~ n1480)  &  (~ n3582) ) ;
 assign n1498 = ( (~ n3576)  &  (~ n4079) ) | ( (~ n1263)  &  (~ n1480)  &  (~ n3576) ) ;
 assign n1504 = ( n4055  &  n847 ) | ( n3728  &  n847 ) | ( n4055  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n1503 = ( (~ Pi20)  &  n840 ) | ( Pi20  &  n843 ) | ( n840  &  n843 ) ;
 assign n1502 = ( n1504  &  n1503 ) | ( n1504  &  n1480 ) ;
 assign n1505 = ( (~ n3579)  &  (~ n4056) ) | ( (~ n1248)  &  (~ n1480)  &  (~ n3579) ) ;
 assign n1508 = ( (~ n1884)  &  (~ n4058) ) | ( (~ n1480)  &  (~ n1538)  &  (~ n1884) ) ;
 assign n1511 = ( (~ n3778)  &  (~ n4060) ) | ( (~ n1480)  &  (~ n1535)  &  (~ n3778) ) ;
 assign n1514 = ( (~ n3582)  &  (~ n4063) ) | ( (~ n1256)  &  (~ n1480)  &  (~ n3582) ) ;
 assign n1517 = ( (~ n3576)  &  (~ n4065) ) | ( (~ n1257)  &  (~ n1480)  &  (~ n3576) ) ;
 assign n1522 = ( Pi15  &  n1472 ) | ( (~ Pi15)  &  n1476 ) | ( n1472  &  n1476 ) ;
 assign n1520 = ( n931  &  n934 ) | ( n931  &  n1522 ) | ( n934  &  (~ n3887) ) | ( n1522  &  (~ n3887) ) ;
 assign n1523 = ( n942  &  n1066 ) | ( n942  &  n1471 ) ;
 assign n1526 = ( n1268  &  n1271 ) | ( n3817  &  n1271 ) | ( n1268  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n1525 = ( n1480 ) | ( (~ n3603) ) ;
 assign n1524 = ( n1523  &  n1526  &  n1257 ) | ( n1523  &  n1526  &  n1525 ) ;
 assign n1528 = ( n1279  &  n1282 ) | ( n3817  &  n1282 ) | ( n1279  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n1527 = ( n1523  &  n1528  &  n1256 ) | ( n1523  &  n1528  &  n1525 ) ;
 assign n1530 = ( n1288  &  n1291 ) | ( n3817  &  n1291 ) | ( n1288  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n1529 = ( n1523  &  n1530  &  n1248 ) | ( n1523  &  n1530  &  n1525 ) ;
 assign n1532 = ( n1529  &  n1527 ) | ( n3735  &  n1527 ) | ( n1529  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1533 = ( n4112  &  n4110  &  n855 ) | ( n4112  &  n4110  &  n3816 ) ;
 assign n1531 = ( n1532  &  n1533  &  n1524 ) | ( n1532  &  n1533  &  n796 ) ;
 assign n1536 = ( n1304  &  n1307 ) | ( n3817  &  n1307 ) | ( n1304  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n1535 = ( (~ Pi20)  &  n886 ) | ( Pi20  &  n888 ) | ( n886  &  n888 ) ;
 assign n1534 = ( n1523  &  n1536  &  n1535 ) | ( n1523  &  n1536  &  n1525 ) ;
 assign n1539 = ( n1314  &  n1317 ) | ( n3817  &  n1317 ) | ( n1314  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n1538 = ( (~ Pi20)  &  n881 ) | ( Pi20  &  n884 ) | ( n881  &  n884 ) ;
 assign n1537 = ( n1523  &  n1539  &  n1538 ) | ( n1523  &  n1539  &  n1525 ) ;
 assign n1541 = ( n1323  &  n1326 ) | ( n3817  &  n1326 ) | ( n1323  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n1540 = ( n1523  &  n1541  &  n1503 ) | ( n1523  &  n1541  &  n1525 ) ;
 assign n1543 = ( n1540  &  n1537 ) | ( n3735  &  n1537 ) | ( n1540  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1544 = ( n4109  &  n4110  &  n845 ) | ( n4109  &  n4110  &  n3816 ) ;
 assign n1542 = ( n1543  &  n1544  &  n1534 ) | ( n1543  &  n1544  &  n796 ) ;
 assign n1546 = ( n1339  &  n1342 ) | ( n3817  &  n1342 ) | ( n1339  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n1545 = ( n1523  &  n1546  &  n1263 ) | ( n1523  &  n1546  &  n1525 ) ;
 assign n1548 = ( n1349  &  n1352 ) | ( n3817  &  n1352 ) | ( n1349  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n1547 = ( n1523  &  n1548  &  n1262 ) | ( n1523  &  n1548  &  n1525 ) ;
 assign n1550 = ( n1358  &  n1361 ) | ( n3817  &  n1361 ) | ( n1358  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n1549 = ( n1523  &  n1550  &  n1254 ) | ( n1523  &  n1550  &  n1525 ) ;
 assign n1552 = ( n1549  &  n1547 ) | ( n3735  &  n1547 ) | ( n1549  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1553 = ( n4113  &  n4110  &  n873 ) | ( n4113  &  n4110  &  n3816 ) ;
 assign n1551 = ( n1552  &  n1553  &  n1545 ) | ( n1552  &  n1553  &  n796 ) ;
 assign n1555 = ( n1374  &  n1377 ) | ( n3817  &  n1377 ) | ( n1374  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n1554 = ( n1523  &  n1555  &  n1260 ) | ( n1523  &  n1555  &  n1525 ) ;
 assign n1557 = ( n1384  &  n1387 ) | ( n3817  &  n1387 ) | ( n1384  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n1556 = ( n1523  &  n1557  &  n1259 ) | ( n1523  &  n1557  &  n1525 ) ;
 assign n1559 = ( n1393  &  n1396 ) | ( n3817  &  n1396 ) | ( n1393  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n1558 = ( n1523  &  n1559  &  n1252 ) | ( n1523  &  n1559  &  n1525 ) ;
 assign n1561 = ( n1558  &  n1556 ) | ( n3735  &  n1556 ) | ( n1558  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1562 = ( n4111  &  n4110  &  n864 ) | ( n4111  &  n4110  &  n3816 ) ;
 assign n1560 = ( n1561  &  n1562  &  n1554 ) | ( n1561  &  n1562  &  n796 ) ;
 assign n1564 = ( n3638  &  Pi27 ) | ( n3638  &  n1470 ) ;
 assign n1563 = ( n1087  &  n1564 ) | ( n1087  &  n1471 ) ;
 assign n1567 = ( n1257  &  n1268 ) | ( n3808  &  n1268 ) | ( n1257  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n1566 = ( (~ Pi27) ) | ( n787 ) ;
 assign n1565 = ( n1563  &  n1567  &  n1271 ) | ( n1563  &  n1567  &  n1566 ) ;
 assign n1569 = ( n1256  &  n1279 ) | ( n3808  &  n1279 ) | ( n1256  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n1568 = ( n1563  &  n1569  &  n1282 ) | ( n1563  &  n1569  &  n1566 ) ;
 assign n1571 = ( n1248  &  n1288 ) | ( n3808  &  n1288 ) | ( n1248  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n1570 = ( n1563  &  n1571  &  n1291 ) | ( n1563  &  n1571  &  n1566 ) ;
 assign n1573 = ( n1570  &  n1568 ) | ( n3735  &  n1568 ) | ( n1570  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1574 = ( n4105  &  n4103  &  n1298 ) | ( n4105  &  n4103  &  n3807 ) ;
 assign n1572 = ( n1573  &  n1574  &  n1565 ) | ( n1573  &  n1574  &  n796 ) ;
 assign n1576 = ( n1535  &  n1304 ) | ( n3808  &  n1304 ) | ( n1535  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n1575 = ( n1563  &  n1576  &  n1307 ) | ( n1563  &  n1576  &  n1566 ) ;
 assign n1578 = ( n1538  &  n1314 ) | ( n3808  &  n1314 ) | ( n1538  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n1577 = ( n1563  &  n1578  &  n1317 ) | ( n1563  &  n1578  &  n1566 ) ;
 assign n1580 = ( n1503  &  n1323 ) | ( n3808  &  n1323 ) | ( n1503  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n1579 = ( n1563  &  n1580  &  n1326 ) | ( n1563  &  n1580  &  n1566 ) ;
 assign n1582 = ( n1579  &  n1577 ) | ( n3735  &  n1577 ) | ( n1579  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1583 = ( n4102  &  n4103  &  n1333 ) | ( n4102  &  n4103  &  n3807 ) ;
 assign n1581 = ( n1582  &  n1583  &  n1575 ) | ( n1582  &  n1583  &  n796 ) ;
 assign n1585 = ( n1263  &  n1339 ) | ( n3808  &  n1339 ) | ( n1263  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n1584 = ( n1563  &  n1585  &  n1342 ) | ( n1563  &  n1585  &  n1566 ) ;
 assign n1587 = ( n1262  &  n1349 ) | ( n3808  &  n1349 ) | ( n1262  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n1586 = ( n1563  &  n1587  &  n1352 ) | ( n1563  &  n1587  &  n1566 ) ;
 assign n1589 = ( n1254  &  n1358 ) | ( n3808  &  n1358 ) | ( n1254  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n1588 = ( n1563  &  n1589  &  n1361 ) | ( n1563  &  n1589  &  n1566 ) ;
 assign n1591 = ( n1588  &  n1586 ) | ( n3735  &  n1586 ) | ( n1588  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1592 = ( n4106  &  n4103  &  n1368 ) | ( n4106  &  n4103  &  n3807 ) ;
 assign n1590 = ( n1591  &  n1592  &  n1584 ) | ( n1591  &  n1592  &  n796 ) ;
 assign n1594 = ( n1260  &  n1374 ) | ( n3808  &  n1374 ) | ( n1260  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n1593 = ( n1563  &  n1594  &  n1377 ) | ( n1563  &  n1594  &  n1566 ) ;
 assign n1596 = ( n1259  &  n1384 ) | ( n3808  &  n1384 ) | ( n1259  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n1595 = ( n1563  &  n1596  &  n1387 ) | ( n1563  &  n1596  &  n1566 ) ;
 assign n1598 = ( n1252  &  n1393 ) | ( n3808  &  n1393 ) | ( n1252  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n1597 = ( n1563  &  n1598  &  n1396 ) | ( n1563  &  n1598  &  n1566 ) ;
 assign n1600 = ( n1597  &  n1595 ) | ( n3735  &  n1595 ) | ( n1597  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1601 = ( n4104  &  n4103  &  n1403 ) | ( n4104  &  n4103  &  n3807 ) ;
 assign n1599 = ( n1600  &  n1601  &  n1593 ) | ( n1600  &  n1601  &  n796 ) ;
 assign n1603 = ( (~ Pi26)  &  n3639 ) | ( n1470  &  n3639 ) ;
 assign n1602 = ( n1471  &  (~ n3804) ) | ( n1603  &  (~ n3804) ) ;
 assign n1607 = ( n1268  &  n1271 ) | ( n3812  &  n1271 ) | ( n1268  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n1606 = ( (~ n161) ) | ( n1480 ) ;
 assign n1605 = ( n1602  &  n1607  &  n1257 ) | ( n1602  &  n1607  &  n1606 ) ;
 assign n1609 = ( n1279  &  n1282 ) | ( n3812  &  n1282 ) | ( n1279  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n1608 = ( n1602  &  n1609  &  n1256 ) | ( n1602  &  n1609  &  n1606 ) ;
 assign n1611 = ( n1288  &  n1291 ) | ( n3812  &  n1291 ) | ( n1288  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n1610 = ( n1602  &  n1611  &  n1248 ) | ( n1602  &  n1611  &  n1606 ) ;
 assign n1613 = ( n1610  &  n1608 ) | ( n3735  &  n1608 ) | ( n1610  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1614 = ( n4098  &  n4096  &  n855 ) | ( n4098  &  n4096  &  n3811 ) ;
 assign n1612 = ( n1613  &  n1614  &  n1605 ) | ( n1613  &  n1614  &  n796 ) ;
 assign n1616 = ( n1304  &  n1307 ) | ( n3812  &  n1307 ) | ( n1304  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n1615 = ( n1602  &  n1616  &  n1535 ) | ( n1602  &  n1616  &  n1606 ) ;
 assign n1618 = ( n1314  &  n1317 ) | ( n3812  &  n1317 ) | ( n1314  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n1617 = ( n1602  &  n1618  &  n1538 ) | ( n1602  &  n1618  &  n1606 ) ;
 assign n1620 = ( n1323  &  n1326 ) | ( n3812  &  n1326 ) | ( n1323  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n1619 = ( n1602  &  n1620  &  n1503 ) | ( n1602  &  n1620  &  n1606 ) ;
 assign n1622 = ( n1619  &  n1617 ) | ( n3735  &  n1617 ) | ( n1619  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1623 = ( n4095  &  n4096  &  n845 ) | ( n4095  &  n4096  &  n3811 ) ;
 assign n1621 = ( n1622  &  n1623  &  n1615 ) | ( n1622  &  n1623  &  n796 ) ;
 assign n1625 = ( n1339  &  n1342 ) | ( n3812  &  n1342 ) | ( n1339  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n1624 = ( n1602  &  n1625  &  n1263 ) | ( n1602  &  n1625  &  n1606 ) ;
 assign n1627 = ( n1349  &  n1352 ) | ( n3812  &  n1352 ) | ( n1349  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n1626 = ( n1602  &  n1627  &  n1262 ) | ( n1602  &  n1627  &  n1606 ) ;
 assign n1629 = ( n1358  &  n1361 ) | ( n3812  &  n1361 ) | ( n1358  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n1628 = ( n1602  &  n1629  &  n1254 ) | ( n1602  &  n1629  &  n1606 ) ;
 assign n1631 = ( n1628  &  n1626 ) | ( n3735  &  n1626 ) | ( n1628  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1632 = ( n4099  &  n4096  &  n873 ) | ( n4099  &  n4096  &  n3811 ) ;
 assign n1630 = ( n1631  &  n1632  &  n1624 ) | ( n1631  &  n1632  &  n796 ) ;
 assign n1634 = ( n1374  &  n1377 ) | ( n3812  &  n1377 ) | ( n1374  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n1633 = ( n1602  &  n1634  &  n1260 ) | ( n1602  &  n1634  &  n1606 ) ;
 assign n1636 = ( n1384  &  n1387 ) | ( n3812  &  n1387 ) | ( n1384  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n1635 = ( n1602  &  n1636  &  n1259 ) | ( n1602  &  n1636  &  n1606 ) ;
 assign n1638 = ( n1393  &  n1396 ) | ( n3812  &  n1396 ) | ( n1393  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n1637 = ( n1602  &  n1638  &  n1252 ) | ( n1602  &  n1638  &  n1606 ) ;
 assign n1640 = ( n1637  &  n1635 ) | ( n3735  &  n1635 ) | ( n1637  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n1641 = ( n4097  &  n4096  &  n864 ) | ( n4097  &  n4096  &  n3811 ) ;
 assign n1639 = ( n1640  &  n1641  &  n1633 ) | ( n1640  &  n1641  &  n796 ) ;
 assign n1645 = ( n1149  &  n3659 ) | ( n3659  &  n3824 ) | ( n1149  &  (~ n3890) ) | ( n3824  &  (~ n3890) ) ;
 assign n1646 = ( n1212  &  n944 ) | ( n3612  &  n944 ) | ( n1212  &  n1218 ) | ( n3612  &  n1218 ) ;
 assign n1644 = ( (~ Ni10) ) | ( n3614 ) ;
 assign n1642 = ( n1645  &  n1646  &  n1644 ) | ( n1645  &  n1646  &  (~ n4833) ) ;
 assign n1647 = ( n933  &  n930 ) | ( n933  &  Ni11 ) | ( n930  &  (~ n1068) ) | ( Ni11  &  (~ n1068) ) ;
 assign n1651 = ( (~ n1068)  &  n1520 ) | ( (~ n1068)  &  n3783 ) | ( n1520  &  (~ n3886) ) | ( n3783  &  (~ n3886) ) ;
 assign n1650 = ( Ni11 ) | ( (~ Ni10) ) ;
 assign n1649 = ( n1651  &  n1264 ) | ( n1651  &  n1650 ) ;
 assign n1655 = ( Ni7  &  n2040 ) ;
 assign n1653 = ( n2040  &  (~ Ni7) ) ;
 assign n1654 = ( Ni9 ) | ( Ni8 ) ;
 assign n1652 = ( (~ n1647)  &  n1655 ) | ( (~ n1647)  &  n1653  &  n1654 ) ;
 assign n1657 = ( n1642 ) | ( n3540 ) | ( (~ n3779) ) ;
 assign n1658 = ( n1649  &  (~ n1652) ) | ( (~ n1653)  &  (~ n1652) ) | ( n1654  &  (~ n1652) ) ;
 assign n1660 = ( (~ Ni32)  &  (~ Ni30) ) ;
 assign n1662 = ( (~ n18) ) | ( n1063 ) ;
 assign n1663 = ( (~ Ni34) ) | ( (~ Ni33) ) ;
 assign n1661 = ( (~ n163)  &  n1662 ) | ( (~ n163)  &  n1663 ) ;
 assign n1665 = ( (~ Ni34)  &  n1661 ) | ( n205  &  n1661 ) ;
 assign n1667 = ( (~ Ni34)  &  n1661 ) | ( n242  &  n1661 ) ;
 assign n1668 = ( (~ Ni34)  &  n1661 ) | ( n287  &  n1661 ) ;
 assign n1670 = ( (~ Ni34) ) | ( (~ n166) ) ;
 assign n1671 = ( n1665  &  n1667 ) | ( n891  &  n1667 ) | ( n1665  &  n310 ) | ( n891  &  n310 ) ;
 assign n1669 = ( n1670  &  n1671  &  n1668 ) | ( n1670  &  n1671  &  n1250 ) ;
 assign n1672 = ( (~ Ni34)  &  n1661 ) | ( n318  &  n1661 ) ;
 assign n1673 = ( (~ Ni34)  &  n1661 ) | ( n343  &  n1661 ) ;
 assign n1674 = ( (~ Ni34)  &  n1661 ) | ( n375  &  n1661 ) ;
 assign n1676 = ( n1672  &  n1673 ) | ( n891  &  n1673 ) | ( n1672  &  n310 ) | ( n891  &  n310 ) ;
 assign n1675 = ( n1670  &  n1676  &  n1674 ) | ( n1670  &  n1676  &  n1250 ) ;
 assign n1677 = ( (~ Ni34)  &  n1661 ) | ( n388  &  n1661 ) ;
 assign n1678 = ( (~ Ni34)  &  n1661 ) | ( n405  &  n1661 ) ;
 assign n1679 = ( (~ Ni34)  &  n1661 ) | ( n268  &  n1661 ) ;
 assign n1681 = ( n1677  &  n1678 ) | ( n891  &  n1678 ) | ( n1677  &  n310 ) | ( n891  &  n310 ) ;
 assign n1680 = ( n1670  &  n1681  &  n1679 ) | ( n1670  &  n1681  &  n1250 ) ;
 assign n1682 = ( (~ Ni34)  &  n1661 ) | ( n427  &  n1661 ) ;
 assign n1683 = ( (~ Ni34)  &  n1661 ) | ( n434  &  n1661 ) ;
 assign n1684 = ( (~ Ni34)  &  n1661 ) | ( n363  &  n1661 ) ;
 assign n1686 = ( n1682  &  n1683 ) | ( n891  &  n1683 ) | ( n1682  &  n310 ) | ( n891  &  n310 ) ;
 assign n1685 = ( n1670  &  n1686  &  n1684 ) | ( n1670  &  n1686  &  n1250 ) ;
 assign n1687 = ( (~ Ni34)  &  n1661 ) | ( n456  &  n1661 ) ;
 assign n1688 = ( (~ Ni34)  &  n1661 ) | ( n482  &  n1661 ) ;
 assign n1689 = ( (~ Ni34)  &  n1661 ) | ( n507  &  n1661 ) ;
 assign n1690 = ( (~ Ni34)  &  n1661 ) | ( n534  &  n1661 ) ;
 assign n1693 = ( n1670  &  n1689 ) | ( n1670  &  n3776 ) ;
 assign n1694 = ( n1687  &  n1688 ) | ( n891  &  n1688 ) | ( n1687  &  n310 ) | ( n891  &  n310 ) ;
 assign n1692 = ( (~ Pi19) ) | ( n3729 ) ;
 assign n1691 = ( n1693  &  n1694  &  n1690 ) | ( n1693  &  n1694  &  n1692 ) ;
 assign n1695 = ( (~ Ni34)  &  n1661 ) | ( n563  &  n1661 ) ;
 assign n1696 = ( (~ Ni34)  &  n1661 ) | ( n584  &  n1661 ) ;
 assign n1697 = ( (~ Ni34)  &  n1661 ) | ( n607  &  n1661 ) ;
 assign n1698 = ( (~ Ni34)  &  n1661 ) | ( n631  &  n1661 ) ;
 assign n1700 = ( n1670  &  n1697 ) | ( n1670  &  n3776 ) ;
 assign n1701 = ( n1695  &  n1696 ) | ( n891  &  n1696 ) | ( n1695  &  n310 ) | ( n891  &  n310 ) ;
 assign n1699 = ( n1700  &  n1701  &  n1698 ) | ( n1700  &  n1701  &  n1692 ) ;
 assign n1702 = ( (~ Ni34)  &  n1661 ) | ( n662  &  n1661 ) ;
 assign n1703 = ( (~ Ni34)  &  n1661 ) | ( n677  &  n1661 ) ;
 assign n1704 = ( (~ Ni34)  &  n1661 ) | ( n687  &  n1661 ) ;
 assign n1705 = ( (~ Ni34)  &  n1661 ) | ( n699  &  n1661 ) ;
 assign n1707 = ( n1670  &  n1704 ) | ( n1670  &  n3776 ) ;
 assign n1708 = ( n1702  &  n1703 ) | ( n891  &  n1703 ) | ( n1702  &  n310 ) | ( n891  &  n310 ) ;
 assign n1706 = ( n1707  &  n1708  &  n1705 ) | ( n1707  &  n1708  &  n1692 ) ;
 assign n1709 = ( (~ Ni34)  &  n1661 ) | ( n713  &  n1661 ) ;
 assign n1710 = ( (~ Ni34)  &  n1661 ) | ( n723  &  n1661 ) ;
 assign n1711 = ( (~ Ni34)  &  n1661 ) | ( n733  &  n1661 ) ;
 assign n1712 = ( (~ Ni34)  &  n1661 ) | ( n740  &  n1661 ) ;
 assign n1714 = ( n1670  &  n1711 ) | ( n1670  &  n3776 ) ;
 assign n1715 = ( n1709  &  n1710 ) | ( n891  &  n1710 ) | ( n1709  &  n310 ) | ( n891  &  n310 ) ;
 assign n1713 = ( n1714  &  n1715  &  n1712 ) | ( n1714  &  n1715  &  n1692 ) ;
 assign n1716 = ( (~ Ni33)  &  n1663 ) | ( (~ n205)  &  n1663 ) ;
 assign n1721 = ( (~ n205)  &  n1716 ) | ( (~ n205)  &  n3836 ) | ( n1716  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1719 = ( (~ n205)  &  n4701 ) | ( n205  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1718 = ( (~ Pi25)  &  n1665  &  n1721 ) | ( n1665  &  n1721  &  n1719 ) ;
 assign n1722 = ( (~ Ni33)  &  n1663 ) | ( (~ n242)  &  n1663 ) ;
 assign n1726 = ( (~ n242)  &  n1722 ) | ( (~ n242)  &  n3836 ) | ( n1722  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1725 = ( (~ n242)  &  n4701 ) | ( n242  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1724 = ( (~ Pi25)  &  n1667  &  n1726 ) | ( n1667  &  n1726  &  n1725 ) ;
 assign n1727 = ( (~ Ni33)  &  n1663 ) | ( (~ n287)  &  n1663 ) ;
 assign n1731 = ( (~ n287)  &  n1727 ) | ( (~ n287)  &  n3836 ) | ( n1727  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1730 = ( (~ n287)  &  n4701 ) | ( n287  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1729 = ( (~ Pi25)  &  n1668  &  n1731 ) | ( n1668  &  n1731  &  n1730 ) ;
 assign n1733 = ( n1718  &  n1724 ) | ( n891  &  n1724 ) | ( n1718  &  n310 ) | ( n891  &  n310 ) ;
 assign n1732 = ( n1670  &  n1733  &  n1729 ) | ( n1670  &  n1733  &  n1250 ) ;
 assign n1734 = ( (~ Ni33)  &  n1663 ) | ( (~ n318)  &  n1663 ) ;
 assign n1738 = ( (~ n318)  &  n1734 ) | ( (~ n318)  &  n3836 ) | ( n1734  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1737 = ( (~ n318)  &  n4701 ) | ( n318  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1736 = ( (~ Pi25)  &  n1672  &  n1738 ) | ( n1672  &  n1738  &  n1737 ) ;
 assign n1739 = ( (~ Ni33)  &  n1663 ) | ( (~ n343)  &  n1663 ) ;
 assign n1743 = ( (~ n343)  &  n1739 ) | ( (~ n343)  &  n3836 ) | ( n1739  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1742 = ( (~ n343)  &  n4701 ) | ( n343  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1741 = ( (~ Pi25)  &  n1673  &  n1743 ) | ( n1673  &  n1743  &  n1742 ) ;
 assign n1744 = ( (~ Ni33)  &  n1663 ) | ( (~ n375)  &  n1663 ) ;
 assign n1748 = ( (~ n375)  &  n1744 ) | ( (~ n375)  &  n3836 ) | ( n1744  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1747 = ( (~ n375)  &  n4701 ) | ( n375  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1746 = ( (~ Pi25)  &  n1674  &  n1748 ) | ( n1674  &  n1748  &  n1747 ) ;
 assign n1750 = ( n1736  &  n1741 ) | ( n891  &  n1741 ) | ( n1736  &  n310 ) | ( n891  &  n310 ) ;
 assign n1749 = ( n1670  &  n1750  &  n1746 ) | ( n1670  &  n1750  &  n1250 ) ;
 assign n1751 = ( (~ Ni33)  &  n1663 ) | ( (~ n388)  &  n1663 ) ;
 assign n1755 = ( (~ n388)  &  n1751 ) | ( (~ n388)  &  n3836 ) | ( n1751  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1754 = ( (~ n388)  &  n4701 ) | ( n388  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1753 = ( (~ Pi25)  &  n1677  &  n1755 ) | ( n1677  &  n1755  &  n1754 ) ;
 assign n1756 = ( (~ Ni33)  &  n1663 ) | ( (~ n405)  &  n1663 ) ;
 assign n1760 = ( (~ n405)  &  n1756 ) | ( (~ n405)  &  n3836 ) | ( n1756  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1759 = ( (~ n405)  &  n4701 ) | ( n405  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1758 = ( (~ Pi25)  &  n1678  &  n1760 ) | ( n1678  &  n1760  &  n1759 ) ;
 assign n1761 = ( (~ Ni33)  &  n1663 ) | ( (~ n268)  &  n1663 ) ;
 assign n1765 = ( (~ n268)  &  n1761 ) | ( (~ n268)  &  n3836 ) | ( n1761  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1764 = ( (~ n268)  &  n4701 ) | ( n268  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1763 = ( (~ Pi25)  &  n1679  &  n1765 ) | ( n1679  &  n1765  &  n1764 ) ;
 assign n1767 = ( n1753  &  n1758 ) | ( n891  &  n1758 ) | ( n1753  &  n310 ) | ( n891  &  n310 ) ;
 assign n1766 = ( n1670  &  n1767  &  n1763 ) | ( n1670  &  n1767  &  n1250 ) ;
 assign n1768 = ( (~ Ni33)  &  n1663 ) | ( (~ n427)  &  n1663 ) ;
 assign n1772 = ( (~ n427)  &  n1768 ) | ( (~ n427)  &  n3836 ) | ( n1768  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1771 = ( (~ n427)  &  n4701 ) | ( n427  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1770 = ( (~ Pi25)  &  n1682  &  n1772 ) | ( n1682  &  n1772  &  n1771 ) ;
 assign n1773 = ( (~ Ni33)  &  n1663 ) | ( (~ n434)  &  n1663 ) ;
 assign n1777 = ( (~ n434)  &  n1773 ) | ( (~ n434)  &  n3836 ) | ( n1773  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1776 = ( (~ n434)  &  n4701 ) | ( n434  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1775 = ( (~ Pi25)  &  n1683  &  n1777 ) | ( n1683  &  n1777  &  n1776 ) ;
 assign n1778 = ( (~ Ni33)  &  n1663 ) | ( (~ n363)  &  n1663 ) ;
 assign n1782 = ( (~ n363)  &  n1778 ) | ( (~ n363)  &  n3836 ) | ( n1778  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1781 = ( (~ n363)  &  n4701 ) | ( n363  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1780 = ( (~ Pi25)  &  n1684  &  n1782 ) | ( n1684  &  n1782  &  n1781 ) ;
 assign n1784 = ( n1770  &  n1775 ) | ( n891  &  n1775 ) | ( n1770  &  n310 ) | ( n891  &  n310 ) ;
 assign n1783 = ( n1670  &  n1784  &  n1780 ) | ( n1670  &  n1784  &  n1250 ) ;
 assign n1785 = ( (~ Ni33)  &  n1663 ) | ( (~ n456)  &  n1663 ) ;
 assign n1789 = ( (~ n456)  &  n1785 ) | ( (~ n456)  &  n3836 ) | ( n1785  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1788 = ( (~ n456)  &  n4701 ) | ( n456  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1787 = ( (~ Pi25)  &  n1687  &  n1789 ) | ( n1687  &  n1789  &  n1788 ) ;
 assign n1790 = ( (~ Ni33)  &  n1663 ) | ( (~ n482)  &  n1663 ) ;
 assign n1794 = ( (~ n482)  &  n1790 ) | ( (~ n482)  &  n3836 ) | ( n1790  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1793 = ( (~ n482)  &  n4701 ) | ( n482  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1792 = ( (~ Pi25)  &  n1688  &  n1794 ) | ( n1688  &  n1794  &  n1793 ) ;
 assign n1795 = ( (~ Ni33)  &  n1663 ) | ( (~ n507)  &  n1663 ) ;
 assign n1797 = ( (~ Ni33)  &  n1663 ) | ( (~ n534)  &  n1663 ) ;
 assign n1801 = ( (~ n534)  &  n1797 ) | ( (~ n534)  &  n3836 ) | ( n1797  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1800 = ( (~ n534)  &  n4701 ) | ( n534  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1799 = ( (~ Pi25)  &  n1690  &  n1801 ) | ( n1690  &  n1801  &  n1800 ) ;
 assign n1803 = ( n1670  &  n3776 ) | ( n1670  &  n4248  &  n4247 ) ;
 assign n1804 = ( n1787  &  n1792 ) | ( n891  &  n1792 ) | ( n1787  &  n310 ) | ( n891  &  n310 ) ;
 assign n1802 = ( n1803  &  n1804  &  n1799 ) | ( n1803  &  n1804  &  n1692 ) ;
 assign n1805 = ( (~ Ni33)  &  n1663 ) | ( (~ n563)  &  n1663 ) ;
 assign n1809 = ( (~ n563)  &  n1805 ) | ( (~ n563)  &  n3836 ) | ( n1805  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1808 = ( (~ n563)  &  n4701 ) | ( n563  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1807 = ( (~ Pi25)  &  n1695  &  n1809 ) | ( n1695  &  n1809  &  n1808 ) ;
 assign n1810 = ( (~ Ni33)  &  n1663 ) | ( (~ n584)  &  n1663 ) ;
 assign n1814 = ( (~ n584)  &  n1810 ) | ( (~ n584)  &  n3836 ) | ( n1810  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1813 = ( (~ n584)  &  n4701 ) | ( n584  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1812 = ( (~ Pi25)  &  n1696  &  n1814 ) | ( n1696  &  n1814  &  n1813 ) ;
 assign n1815 = ( (~ Ni33)  &  n1663 ) | ( (~ n607)  &  n1663 ) ;
 assign n1817 = ( (~ Ni33)  &  n1663 ) | ( (~ n631)  &  n1663 ) ;
 assign n1821 = ( (~ n631)  &  n1817 ) | ( (~ n631)  &  n3836 ) | ( n1817  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1820 = ( (~ n631)  &  n4701 ) | ( n631  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1819 = ( (~ Pi25)  &  n1698  &  n1821 ) | ( n1698  &  n1821  &  n1820 ) ;
 assign n1823 = ( n1670  &  n3776 ) | ( n1670  &  n4252  &  n4251 ) ;
 assign n1824 = ( n1807  &  n1812 ) | ( n891  &  n1812 ) | ( n1807  &  n310 ) | ( n891  &  n310 ) ;
 assign n1822 = ( n1823  &  n1824  &  n1819 ) | ( n1823  &  n1824  &  n1692 ) ;
 assign n1825 = ( (~ Ni33)  &  n1663 ) | ( (~ n662)  &  n1663 ) ;
 assign n1829 = ( (~ n662)  &  n1825 ) | ( (~ n662)  &  n3836 ) | ( n1825  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1828 = ( (~ n662)  &  n4701 ) | ( n662  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1827 = ( (~ Pi25)  &  n1702  &  n1829 ) | ( n1702  &  n1829  &  n1828 ) ;
 assign n1830 = ( (~ Ni33)  &  n1663 ) | ( (~ n677)  &  n1663 ) ;
 assign n1834 = ( (~ n677)  &  n1830 ) | ( (~ n677)  &  n3836 ) | ( n1830  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1833 = ( (~ n677)  &  n4701 ) | ( n677  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1832 = ( (~ Pi25)  &  n1703  &  n1834 ) | ( n1703  &  n1834  &  n1833 ) ;
 assign n1835 = ( (~ Ni33)  &  n1663 ) | ( (~ n687)  &  n1663 ) ;
 assign n1837 = ( (~ Ni33)  &  n1663 ) | ( (~ n699)  &  n1663 ) ;
 assign n1841 = ( (~ n699)  &  n1837 ) | ( (~ n699)  &  n3836 ) | ( n1837  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1840 = ( (~ n699)  &  n4701 ) | ( n699  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1839 = ( (~ Pi25)  &  n1705  &  n1841 ) | ( n1705  &  n1841  &  n1840 ) ;
 assign n1843 = ( n1670  &  n3776 ) | ( n1670  &  n4250  &  n4249 ) ;
 assign n1844 = ( n1827  &  n1832 ) | ( n891  &  n1832 ) | ( n1827  &  n310 ) | ( n891  &  n310 ) ;
 assign n1842 = ( n1843  &  n1844  &  n1839 ) | ( n1843  &  n1844  &  n1692 ) ;
 assign n1845 = ( (~ Ni33)  &  n1663 ) | ( (~ n713)  &  n1663 ) ;
 assign n1849 = ( (~ n713)  &  n1845 ) | ( (~ n713)  &  n3836 ) | ( n1845  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1848 = ( (~ n713)  &  n4701 ) | ( n713  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1847 = ( (~ Pi25)  &  n1709  &  n1849 ) | ( n1709  &  n1849  &  n1848 ) ;
 assign n1850 = ( (~ Ni33)  &  n1663 ) | ( (~ n723)  &  n1663 ) ;
 assign n1854 = ( (~ n723)  &  n1850 ) | ( (~ n723)  &  n3836 ) | ( n1850  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1853 = ( (~ n723)  &  n4701 ) | ( n723  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1852 = ( (~ Pi25)  &  n1710  &  n1854 ) | ( n1710  &  n1854  &  n1853 ) ;
 assign n1855 = ( (~ Ni33)  &  n1663 ) | ( (~ n733)  &  n1663 ) ;
 assign n1857 = ( (~ Ni33)  &  n1663 ) | ( (~ n740)  &  n1663 ) ;
 assign n1861 = ( (~ n740)  &  n1857 ) | ( (~ n740)  &  n3836 ) | ( n1857  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n1860 = ( (~ n740)  &  n4701 ) | ( n740  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1859 = ( (~ Pi25)  &  n1712  &  n1861 ) | ( n1712  &  n1861  &  n1860 ) ;
 assign n1863 = ( n1670  &  n3776 ) | ( n1670  &  n4254  &  n4253 ) ;
 assign n1864 = ( n1847  &  n1852 ) | ( n891  &  n1852 ) | ( n1847  &  n310 ) | ( n891  &  n310 ) ;
 assign n1862 = ( n1863  &  n1864  &  n1859 ) | ( n1863  &  n1864  &  n1692 ) ;
 assign n1867 = ( (~ n163)  &  n1670 ) ;
 assign n1868 = ( n268  &  n1761 ) | ( n3842  &  n1761 ) | ( n268  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1866 = ( (~ Pi22) ) | ( (~ Pi21) ) ;
 assign n1865 = ( n1867  &  n1868  &  n1764 ) | ( n1867  &  n1868  &  n1866 ) ;
 assign n1870 = ( n363  &  n1778 ) | ( n3842  &  n1778 ) | ( n363  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1869 = ( n1867  &  n1870  &  n1781 ) | ( n1867  &  n1870  &  n1866 ) ;
 assign n1872 = ( n677  &  n1830 ) | ( n3842  &  n1830 ) | ( n677  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1871 = ( n1867  &  n1872  &  n1833 ) | ( n1867  &  n1872  &  n1866 ) ;
 assign n1874 = ( n699  &  n1837 ) | ( n3842  &  n1837 ) | ( n699  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1873 = ( n1867  &  n1874  &  n1840 ) | ( n1867  &  n1874  &  n1866 ) ;
 assign n1876 = ( n405  &  n1756 ) | ( n3842  &  n1756 ) | ( n405  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1875 = ( n1867  &  n1876  &  n1759 ) | ( n1867  &  n1876  &  n1866 ) ;
 assign n1878 = ( n723  &  n1850 ) | ( n3842  &  n1850 ) | ( n723  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1877 = ( n1867  &  n1878  &  n1853 ) | ( n1867  &  n1878  &  n1866 ) ;
 assign n1880 = ( n740  &  n1857 ) | ( n3842  &  n1857 ) | ( n740  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1879 = ( n1867  &  n1880  &  n1860 ) | ( n1867  &  n1880  &  n1866 ) ;
 assign n1882 = ( n434  &  n1773 ) | ( n3842  &  n1773 ) | ( n434  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1881 = ( n1867  &  n1882  &  n1776 ) | ( n1867  &  n1882  &  n1866 ) ;
 assign n1885 = ( n1875  &  n1881 ) | ( n3777  &  n1881 ) | ( n1875  &  n3579 ) | ( n3777  &  n3579 ) ;
 assign n1886 = ( n4323  &  n1879 ) | ( n4323  &  n3576 ) ;
 assign n1884 = ( Pi16 ) | ( n3738 ) ;
 assign n1883 = ( n1885  &  n1886  &  n1871 ) | ( n1885  &  n1886  &  n1884 ) ;
 assign n1888 = ( n662  &  n1825 ) | ( n3842  &  n1825 ) | ( n662  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1887 = ( n1867  &  n1888  &  n1828 ) | ( n1867  &  n1888  &  n1866 ) ;
 assign n1891 = ( n687  &  n1835 ) | ( n3842  &  n1835 ) | ( n687  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1890 = ( (~ n687)  &  n4701 ) | ( n687  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1889 = ( n1867  &  n1891  &  n1890 ) | ( n1867  &  n1891  &  n1866 ) ;
 assign n1893 = ( n388  &  n1751 ) | ( n3842  &  n1751 ) | ( n388  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1892 = ( n1867  &  n1893  &  n1754 ) | ( n1867  &  n1893  &  n1866 ) ;
 assign n1895 = ( n713  &  n1845 ) | ( n3842  &  n1845 ) | ( n713  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1894 = ( n1867  &  n1895  &  n1848 ) | ( n1867  &  n1895  &  n1866 ) ;
 assign n1898 = ( n733  &  n1855 ) | ( n3842  &  n1855 ) | ( n733  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1897 = ( (~ n733)  &  n4701 ) | ( n733  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1896 = ( n1867  &  n1898  &  n1897 ) | ( n1867  &  n1898  &  n1866 ) ;
 assign n1900 = ( n427  &  n1768 ) | ( n3842  &  n1768 ) | ( n427  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1899 = ( n1867  &  n1900  &  n1771 ) | ( n1867  &  n1900  &  n1866 ) ;
 assign n1902 = ( n1892  &  n1899 ) | ( n3777  &  n1899 ) | ( n1892  &  n3579 ) | ( n3777  &  n3579 ) ;
 assign n1903 = ( n4322  &  n1896 ) | ( n4322  &  n3576 ) ;
 assign n1901 = ( n1902  &  n1903  &  n1887 ) | ( n1902  &  n1903  &  n1884 ) ;
 assign n1905 = ( n287  &  n1727 ) | ( n3842  &  n1727 ) | ( n287  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1904 = ( n1867  &  n1905  &  n1730 ) | ( n1867  &  n1905  &  n1866 ) ;
 assign n1907 = ( n375  &  n1744 ) | ( n3842  &  n1744 ) | ( n375  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1906 = ( n1867  &  n1907  &  n1747 ) | ( n1867  &  n1907  &  n1866 ) ;
 assign n1909 = ( n482  &  n1790 ) | ( n3842  &  n1790 ) | ( n482  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1908 = ( n1867  &  n1909  &  n1793 ) | ( n1867  &  n1909  &  n1866 ) ;
 assign n1911 = ( n534  &  n1797 ) | ( n3842  &  n1797 ) | ( n534  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1910 = ( n1867  &  n1911  &  n1800 ) | ( n1867  &  n1911  &  n1866 ) ;
 assign n1913 = ( n242  &  n1722 ) | ( n3842  &  n1722 ) | ( n242  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1912 = ( n1867  &  n1913  &  n1725 ) | ( n1867  &  n1913  &  n1866 ) ;
 assign n1915 = ( n584  &  n1810 ) | ( n3842  &  n1810 ) | ( n584  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1914 = ( n1867  &  n1915  &  n1813 ) | ( n1867  &  n1915  &  n1866 ) ;
 assign n1917 = ( n631  &  n1817 ) | ( n3842  &  n1817 ) | ( n631  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1916 = ( n1867  &  n1917  &  n1820 ) | ( n1867  &  n1917  &  n1866 ) ;
 assign n1919 = ( n343  &  n1739 ) | ( n3842  &  n1739 ) | ( n343  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1918 = ( n1867  &  n1919  &  n1742 ) | ( n1867  &  n1919  &  n1866 ) ;
 assign n1921 = ( n1912  &  n1918 ) | ( n3777  &  n1918 ) | ( n1912  &  n3579 ) | ( n3777  &  n3579 ) ;
 assign n1922 = ( n4320  &  n1916 ) | ( n4320  &  n3576 ) ;
 assign n1920 = ( n1921  &  n1922  &  n1908 ) | ( n1921  &  n1922  &  n1884 ) ;
 assign n1924 = ( n456  &  n1785 ) | ( n3842  &  n1785 ) | ( n456  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1923 = ( n1867  &  n1924  &  n1788 ) | ( n1867  &  n1924  &  n1866 ) ;
 assign n1927 = ( n507  &  n1795 ) | ( n3842  &  n1795 ) | ( n507  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1926 = ( (~ n507)  &  n4701 ) | ( n507  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1925 = ( n1867  &  n1927  &  n1926 ) | ( n1867  &  n1927  &  n1866 ) ;
 assign n1929 = ( n205  &  n1716 ) | ( n3842  &  n1716 ) | ( n205  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1928 = ( n1867  &  n1929  &  n1719 ) | ( n1867  &  n1929  &  n1866 ) ;
 assign n1931 = ( n563  &  n1805 ) | ( n3842  &  n1805 ) | ( n563  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1930 = ( n1867  &  n1931  &  n1808 ) | ( n1867  &  n1931  &  n1866 ) ;
 assign n1934 = ( n607  &  n1815 ) | ( n3842  &  n1815 ) | ( n607  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1933 = ( (~ n607)  &  n4701 ) | ( n607  &  n4702 ) | ( n4701  &  n4702 ) ;
 assign n1932 = ( n1867  &  n1934  &  n1933 ) | ( n1867  &  n1934  &  n1866 ) ;
 assign n1936 = ( n318  &  n1734 ) | ( n3842  &  n1734 ) | ( n318  &  n3839 ) | ( n3842  &  n3839 ) ;
 assign n1935 = ( n1867  &  n1936  &  n1737 ) | ( n1867  &  n1936  &  n1866 ) ;
 assign n1938 = ( n1928  &  n1935 ) | ( n3777  &  n1935 ) | ( n1928  &  n3579 ) | ( n3777  &  n3579 ) ;
 assign n1939 = ( n4319  &  n1932 ) | ( n4319  &  n3576 ) ;
 assign n1937 = ( n1938  &  n1939  &  n1923 ) | ( n1938  &  n1939  &  n1884 ) ;
 assign n1940 = ( (~ Ni34)  &  (~ n268) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1941 = ( (~ Ni34)  &  (~ n363) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1942 = ( (~ Ni34)  &  (~ n677) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1943 = ( (~ Ni34)  &  (~ n699) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1944 = ( (~ Ni34)  &  (~ n405) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1945 = ( (~ Ni34)  &  (~ n723) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1946 = ( (~ Ni34)  &  (~ n740) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1947 = ( (~ Ni34)  &  (~ n434) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1948 = ( (~ n3777)  &  (~ n3841) ) | ( (~ n3777)  &  (~ n4303) ) ;
 assign n1951 = ( (~ n3582)  &  (~ n3841) ) | ( (~ n3582)  &  (~ n4307) ) ;
 assign n1953 = ( (~ Ni34)  &  (~ n662) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1954 = ( (~ Ni34)  &  (~ n687) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1955 = ( (~ Ni34)  &  (~ n388) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1956 = ( (~ Ni34)  &  (~ n713) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1957 = ( (~ Ni34)  &  (~ n733) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1958 = ( (~ Ni34)  &  (~ n427) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1959 = ( (~ n3777)  &  (~ n3841) ) | ( (~ n3777)  &  (~ n4291) ) ;
 assign n1961 = ( (~ n3582)  &  (~ n3841) ) | ( (~ n3582)  &  (~ n4295) ) ;
 assign n1965 = ( n2939  &  Pi16 ) ;
 assign n1963 = ( n1965  &  (~ n3841) ) | ( n1965  &  (~ n4290) ) ;
 assign n1966 = ( (~ Ni34)  &  (~ n287) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1967 = ( (~ Ni34)  &  (~ n375) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1968 = ( (~ Ni34)  &  (~ n482) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1969 = ( (~ Ni34)  &  (~ n534) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1970 = ( (~ Ni34)  &  (~ n242) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1971 = ( (~ Ni34)  &  (~ n584) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1972 = ( (~ Ni34)  &  (~ n631) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1973 = ( (~ Ni34)  &  (~ n343) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1974 = ( (~ n3777)  &  (~ n3841) ) | ( (~ n3777)  &  (~ n4273) ) ;
 assign n1976 = ( (~ n3582)  &  (~ n3841) ) | ( (~ n3582)  &  (~ n4277) ) ;
 assign n1978 = ( (~ Ni34)  &  (~ n456) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1979 = ( (~ Ni34)  &  (~ n507) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1980 = ( (~ Ni34)  &  (~ n205) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1981 = ( (~ Ni34)  &  (~ n563) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1982 = ( (~ Ni34)  &  (~ n607) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1983 = ( (~ Ni34)  &  (~ n318) ) | ( (~ Ni34)  &  n1063 ) ;
 assign n1984 = ( (~ n3777)  &  (~ n3841) ) | ( (~ n3777)  &  (~ n4261) ) ;
 assign n1986 = ( (~ n3582)  &  (~ n3841) ) | ( (~ n3582)  &  (~ n4265) ) ;
 assign n1988 = ( n1965  &  (~ n3841) ) | ( n1965  &  (~ n4260) ) ;
 assign n1994 = ( n4325  &  n3831 ) | ( n4325  &  n4321  &  n4324 ) ;
 assign n1993 = ( (~ Pi15) ) | ( n3113 ) ;
 assign n1991 = ( n1865  &  n1869 ) | ( n1865  &  (~ n1965) ) | ( n1869  &  (~ n3618) ) | ( (~ n1965)  &  (~ n3618) ) ;
 assign n1992 = ( Pi20  &  n1883 ) | ( (~ Pi20)  &  n1901 ) | ( n1883  &  n1901 ) ;
 assign n1990 = ( n1994  &  n1993 ) | ( n1994  &  n1991  &  n1992 ) ;
 assign n1995 = ( (~ Ni34)  &  n1670 ) | ( n1471  &  n1670 ) ;
 assign n1997 = ( (~ Pi25) ) | ( n3727 ) ;
 assign n1996 = ( n1954  &  n1943 ) | ( n1997  &  n1943 ) | ( n1954  &  n787 ) | ( n1997  &  n787 ) ;
 assign n1998 = ( n1953  &  n1942 ) | ( n1997  &  n1942 ) | ( n1953  &  n787 ) | ( n1997  &  n787 ) ;
 assign n1999 = ( n1955  &  n1944 ) | ( n1997  &  n1944 ) | ( n1955  &  n787 ) | ( n1997  &  n787 ) ;
 assign n2000 = ( n1957  &  n1946 ) | ( n1997  &  n1946 ) | ( n1957  &  n787 ) | ( n1997  &  n787 ) ;
 assign n2001 = ( n1956  &  n1945 ) | ( n1997  &  n1945 ) | ( n1956  &  n787 ) | ( n1997  &  n787 ) ;
 assign n2002 = ( n1958  &  n1947 ) | ( n1997  &  n1947 ) | ( n1958  &  n787 ) | ( n1997  &  n787 ) ;
 assign n2003 = ( Pi16  &  (~ n1474)  &  (~ n1941) ) | ( (~ n1474)  &  (~ n1940)  &  (~ n1941) ) ;
 assign n2007 = ( n1979  &  n1969 ) | ( n1997  &  n1969 ) | ( n1979  &  n787 ) | ( n1997  &  n787 ) ;
 assign n2008 = ( n1978  &  n1968 ) | ( n1997  &  n1968 ) | ( n1978  &  n787 ) | ( n1997  &  n787 ) ;
 assign n2009 = ( n1980  &  n1970 ) | ( n1997  &  n1970 ) | ( n1980  &  n787 ) | ( n1997  &  n787 ) ;
 assign n2010 = ( n1982  &  n1972 ) | ( n1997  &  n1972 ) | ( n1982  &  n787 ) | ( n1997  &  n787 ) ;
 assign n2011 = ( n1981  &  n1971 ) | ( n1997  &  n1971 ) | ( n1981  &  n787 ) | ( n1997  &  n787 ) ;
 assign n2012 = ( n1983  &  n1973 ) | ( n1997  &  n1973 ) | ( n1983  &  n787 ) | ( n1997  &  n787 ) ;
 assign n2013 = ( Pi16  &  (~ n1474)  &  (~ n1967) ) | ( (~ n1474)  &  (~ n1966)  &  (~ n1967) ) ;
 assign n2017 = ( (~ Pi15)  &  (~ n4698) ) | ( (~ n4241)  &  (~ n4698) ) | ( (~ n4245)  &  (~ n4698) ) ;
 assign n2016 = ( (~ n3476)  &  (~ n3893) ) | ( n2017  &  (~ n3476)  &  (~ n3775) ) ;
 assign n2025 = ( (~ Ni35) ) | ( Ni30 ) ;
 assign n2024 = ( (~ Ni35)  &  n694  &  n2025 ) | ( n694  &  n837  &  n2025 ) ;
 assign n2028 = ( Ni32 ) | ( n3845 ) ;
 assign n2026 = ( (~ Pi26)  &  n2024 ) | ( n2024  &  n2028 ) ;
 assign n2031 = ( n1068 ) | ( n3568 ) ;
 assign n2029 = ( Ni35  &  n2031 ) | ( Ni35  &  (~ n3662) ) ;
 assign n2032 = ( (~ n1655)  &  (~ n1653) ) | ( (~ n1655)  &  (~ n2049) ) ;
 assign n2036 = ( n2029  &  (~ n2032) ) | ( (~ n2026)  &  (~ n2031)  &  (~ n2032) ) ;
 assign n2042 = ( (~ n1653) ) | ( n2049 ) | ( n4716 ) | ( n4717 ) ;
 assign n2040 = ( (~ n3540)  &  (~ n3779) ) ;
 assign n2045 = ( (~ Ni31) ) | ( (~ Ni36) ) ;
 assign n2043 = ( Ni30  &  n281  &  n2045 ) | ( (~ Ni36)  &  n281  &  n2045 ) ;
 assign n2046 = ( (~ Pi27)  &  n2043 ) | ( n2028  &  n2043 ) ;
 assign n2050 = ( Ni36  &  (~ n4720) ) | ( (~ n2031)  &  (~ n4720) ) ;
 assign n2049 = ( Ni8 ) | ( n3844 ) ;
 assign n2048 = ( n2050  &  n1655 ) | ( n2050  &  n1653  &  n2049 ) ;
 assign n2052 = ( (~ n1653) ) | ( n2049 ) | ( n4718 ) | ( n4719 ) ;
 assign n2055 = ( (~ Ni31)  &  Ni30 ) ;
 assign n2053 = ( (~ Ni32)  &  n2055  &  (~ n4724) ) ;
 assign n2056 = ( (~ Ni30)  &  (~ n200) ) | ( Ni37  &  (~ Ni30)  &  (~ n4724) ) ;
 assign n2058 = ( (~ Pi20) ) | ( n3848 ) | ( n3849 ) ;
 assign n2059 = ( n3846 ) | ( n3849 ) | ( Pi20 ) ;
 assign n2060 = ( n3846 ) | ( n3847 ) | ( Pi20 ) ;
 assign n2061 = ( (~ Pi20) ) | ( n3847 ) | ( n3848 ) ;
 assign n2057 = ( n2058  &  n2059  &  n2060  &  n2061 ) ;
 assign n2062 = ( n663 ) | ( n153  &  Ni30 ) ;
 assign n2063 = ( (~ n153)  &  (~ n200) ) | ( Ni37  &  n24  &  (~ n153) ) ;
 assign n2065 = ( (~ Ni31) ) | ( Ni30 ) ;
 assign n2064 = ( Ni45  &  Ni32 ) | ( Ni45  &  n2065 ) ;
 assign n2066 = ( (~ Ni6) ) | ( Ni5 ) ;
 assign n2069 = ( (~ Ni32) ) | ( Ni30 ) ;
 assign n2068 = ( Ni30 ) | ( Ni31 ) ;
 assign n2073 = ( Pi21 ) | ( (~ Ni32) ) ;
 assign n2071 = ( Pi22 ) | ( n3667 ) ;
 assign n2070 = ( (~ Pi21)  &  n2073 ) | ( n2073  &  n2071 ) ;
 assign n2074 = ( (~ n180)  &  n2069 ) | ( n2069  &  n2068 ) ;
 assign n2079 = ( Ni47  &  (~ Ni45) ) | ( (~ Ni45)  &  (~ Ni43) ) ;
 assign n2078 = ( Ni41 ) | ( Ni42 ) ;
 assign n2076 = ( Ni47  &  n2079 ) | ( n2079  &  n2078 ) | ( n2079  &  (~ n3120) ) ;
 assign n2081 = ( n2079  &  n2106 ) ;
 assign n2082 = ( n2184 ) | ( Ni40 ) ;
 assign n2083 = ( (~ Ni37) ) | ( Ni47 ) | ( Ni38 ) ;
 assign n2084 = ( n3666 ) | ( n3724 ) ;
 assign n2080 = ( n2081  &  n2082  &  n2083  &  n2084 ) ;
 assign n2086 = ( Ni38 ) | ( n3666 ) ;
 assign n2087 = ( (~ Ni35) ) | ( Ni36 ) ;
 assign n2085 = ( n2080  &  n2086 ) | ( n2080  &  n2087 ) ;
 assign n2088 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2085) ) ;
 assign n2091 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2085) ) ;
 assign n2094 = ( (~ n18) ) | ( n153 ) ;
 assign n2093 = ( n153  &  n2091 ) ;
 assign n2092 = ( n18  &  n2094 ) | ( n2094  &  n2093 ) ;
 assign n2096 = ( (~ Ni44)  &  (~ Ni43) ) ;
 assign n2095 = ( n2079  &  Ni47 ) | ( n2079  &  n2096 ) | ( n2079  &  n2078 ) ;
 assign n2098 = ( n2190 ) | ( Ni40 ) ;
 assign n2099 = ( n3666 ) | ( n3725 ) ;
 assign n2097 = ( n2081  &  n2098  &  n2083  &  n2099 ) ;
 assign n2100 = ( n2097  &  n2086 ) | ( n2097  &  n2087 ) ;
 assign n2101 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2100) ) ;
 assign n2103 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2100) ) ;
 assign n2105 = ( n153  &  n2103 ) ;
 assign n2104 = ( n18  &  n2094 ) | ( n2094  &  n2105 ) ;
 assign n2106 = ( (~ Ni41) ) | ( n3666 ) ;
 assign n2108 = ( n2086  &  n2083  &  n2081 ) ;
 assign n2107 = ( n2081  &  n2083  &  Ni36 ) | ( n2081  &  n2083  &  n2108 ) ;
 assign n2109 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2107) ) ;
 assign n2111 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2107) ) ;
 assign n2113 = ( n153  &  n2111 ) ;
 assign n2112 = ( n18  &  n2094 ) | ( n2094  &  n2113 ) ;
 assign n2116 = ( n2378  &  n4363 ) | ( n1250  &  n4363 ) | ( n2378  &  n891 ) | ( n1250  &  n891 ) ;
 assign n2115 = ( n2101  &  n2104 ) ;
 assign n2114 = ( n2070  &  n2116  &  n2115 ) | ( n2070  &  n2116  &  n310 ) ;
 assign n2118 = ( n2076 ) | ( Ni40 ) ;
 assign n2117 = ( n2079  &  n2118  &  n2083  &  n2084 ) ;
 assign n2119 = ( n2117  &  n2086 ) | ( n2117  &  n2087 ) ;
 assign n2120 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2119) ) ;
 assign n2122 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2119) ) ;
 assign n2124 = ( n153  &  n2122 ) ;
 assign n2123 = ( n18  &  n2094 ) | ( n2094  &  n2124 ) ;
 assign n2126 = ( n2095 ) | ( Ni40 ) ;
 assign n2125 = ( n2079  &  n2126  &  n2083  &  n2099 ) ;
 assign n2127 = ( n2125  &  n2086 ) | ( n2125  &  n2087 ) ;
 assign n2128 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2127) ) ;
 assign n2130 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2127) ) ;
 assign n2132 = ( n153  &  n2130 ) ;
 assign n2131 = ( n18  &  n2094 ) | ( n2094  &  n2132 ) ;
 assign n2134 = ( n2086  &  n2083  &  n2079 ) ;
 assign n2133 = ( n2079  &  n2083  &  Ni36 ) | ( n2079  &  n2083  &  n2134 ) ;
 assign n2135 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2133) ) ;
 assign n2137 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2133) ) ;
 assign n2139 = ( n153  &  n2137 ) ;
 assign n2138 = ( n18  &  n2094 ) | ( n2094  &  n2139 ) ;
 assign n2142 = ( n2379  &  n4365 ) | ( n1250  &  n4365 ) | ( n2379  &  n891 ) | ( n1250  &  n891 ) ;
 assign n2141 = ( n2128  &  n2131 ) ;
 assign n2140 = ( n2070  &  n2142  &  n2141 ) | ( n2070  &  n2142  &  n310 ) ;
 assign n2143 = ( n2080  &  n2086 ) | ( n2080  &  (~ n2199) ) ;
 assign n2145 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2143) ) ;
 assign n2147 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2143) ) ;
 assign n2149 = ( n153  &  n2147 ) ;
 assign n2148 = ( n18  &  n2094 ) | ( n2094  &  n2149 ) ;
 assign n2150 = ( n2086  &  n2097 ) | ( n2097  &  (~ n2199) ) ;
 assign n2151 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2150) ) ;
 assign n2153 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2150) ) ;
 assign n2155 = ( n153  &  n2153 ) ;
 assign n2154 = ( n18  &  n2094 ) | ( n2094  &  n2155 ) ;
 assign n2156 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2108) ) ;
 assign n2158 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2108) ) ;
 assign n2160 = ( n153  &  n2158 ) ;
 assign n2159 = ( n18  &  n2094 ) | ( n2094  &  n2160 ) ;
 assign n2163 = ( n2351  &  n4373 ) | ( n1250  &  n4373 ) | ( n2351  &  n891 ) | ( n1250  &  n891 ) ;
 assign n2162 = ( n2151  &  n2154 ) ;
 assign n2161 = ( n2070  &  n2163  &  n2162 ) | ( n2070  &  n2163  &  n310 ) ;
 assign n2164 = ( n2086  &  n2117 ) | ( n2117  &  (~ n2199) ) ;
 assign n2165 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2164) ) ;
 assign n2167 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2164) ) ;
 assign n2169 = ( n153  &  n2167 ) ;
 assign n2168 = ( n18  &  n2094 ) | ( n2094  &  n2169 ) ;
 assign n2170 = ( n2086  &  n2125 ) | ( n2125  &  (~ n2199) ) ;
 assign n2171 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2170) ) ;
 assign n2173 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2170) ) ;
 assign n2175 = ( n153  &  n2173 ) ;
 assign n2174 = ( n18  &  n2094 ) | ( n2094  &  n2175 ) ;
 assign n2176 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2134) ) ;
 assign n2178 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2134) ) ;
 assign n2180 = ( n153  &  n2178 ) ;
 assign n2179 = ( n18  &  n2094 ) | ( n2094  &  n2180 ) ;
 assign n2183 = ( n2352  &  n4375 ) | ( n1250  &  n4375 ) | ( n2352  &  n891 ) | ( n1250  &  n891 ) ;
 assign n2182 = ( n2171  &  n2174 ) ;
 assign n2181 = ( n2070  &  n2183  &  n2182 ) | ( n2070  &  n2183  &  n310 ) ;
 assign n2184 = ( n2106  &  n2076 ) ;
 assign n2185 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n3851) ) ;
 assign n2187 = ( n2069  &  n2068 ) | ( n2069  &  (~ n3851) ) ;
 assign n2189 = ( n153  &  n2187 ) ;
 assign n2188 = ( n18  &  n2094 ) | ( n2094  &  n2189 ) ;
 assign n2190 = ( n2106  &  n2095 ) ;
 assign n2191 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n3852) ) ;
 assign n2193 = ( n2069  &  n2068 ) | ( n2069  &  (~ n3852) ) ;
 assign n2195 = ( n153  &  n2193 ) ;
 assign n2194 = ( n18  &  n2094 ) | ( n2094  &  n2195 ) ;
 assign n2197 = ( n2184 ) | ( (~ Ni40) ) ;
 assign n2196 = ( n2081  &  n2197  &  n2083  &  n2084 ) ;
 assign n2199 = ( Ni35 ) | ( Ni36 ) ;
 assign n2198 = ( n2196  &  n2086 ) | ( n2196  &  n2199 ) ;
 assign n2200 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2198) ) ;
 assign n2202 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2198) ) ;
 assign n2204 = ( n153  &  n2202 ) ;
 assign n2203 = ( n18  &  n2094 ) | ( n2094  &  n2204 ) ;
 assign n2206 = ( n2190 ) | ( (~ Ni40) ) ;
 assign n2205 = ( n2081  &  n2206  &  n2083  &  n2099 ) ;
 assign n2207 = ( n2205  &  n2086 ) | ( n2205  &  n2199 ) ;
 assign n2208 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2207) ) ;
 assign n2210 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2207) ) ;
 assign n2212 = ( n153  &  n2210 ) ;
 assign n2211 = ( n18  &  n2094 ) | ( n2094  &  n2212 ) ;
 assign n2215 = ( n4368  &  n2422 ) | ( n3776  &  n2422 ) | ( n4368  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n2216 = ( n2070  &  n2425 ) | ( n2070  &  n310 ) ;
 assign n2214 = ( n2185  &  n2188 ) ;
 assign n2213 = ( n2215  &  n2216  &  n2214 ) | ( n2215  &  n2216  &  n891 ) ;
 assign n2217 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n3854) ) ;
 assign n2219 = ( n2069  &  n2068 ) | ( n2069  &  (~ n3854) ) ;
 assign n2221 = ( n153  &  n2219 ) ;
 assign n2220 = ( n18  &  n2094 ) | ( n2094  &  n2221 ) ;
 assign n2222 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n3855) ) ;
 assign n2224 = ( n2069  &  n2068 ) | ( n2069  &  (~ n3855) ) ;
 assign n2226 = ( n153  &  n2224 ) ;
 assign n2225 = ( n18  &  n2094 ) | ( n2094  &  n2226 ) ;
 assign n2228 = ( n2076 ) | ( (~ Ni40) ) ;
 assign n2227 = ( n2079  &  n2228  &  n2083  &  n2084 ) ;
 assign n2229 = ( n2227  &  n2086 ) | ( n2227  &  n2199 ) ;
 assign n2230 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2229) ) ;
 assign n2232 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2229) ) ;
 assign n2234 = ( n153  &  n2232 ) ;
 assign n2233 = ( n18  &  n2094 ) | ( n2094  &  n2234 ) ;
 assign n2236 = ( n2095 ) | ( (~ Ni40) ) ;
 assign n2235 = ( n2079  &  n2236  &  n2083  &  n2099 ) ;
 assign n2237 = ( n2235  &  n2086 ) | ( n2235  &  n2199 ) ;
 assign n2238 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2237) ) ;
 assign n2240 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2237) ) ;
 assign n2242 = ( n153  &  n2240 ) ;
 assign n2241 = ( n18  &  n2094 ) | ( n2094  &  n2242 ) ;
 assign n2245 = ( n4371  &  n2410 ) | ( n3776  &  n2410 ) | ( n4371  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n2246 = ( n2070  &  n2414 ) | ( n2070  &  n310 ) ;
 assign n2244 = ( n2217  &  n2220 ) ;
 assign n2243 = ( n2245  &  n2246  &  n2244 ) | ( n2245  &  n2246  &  n891 ) ;
 assign n2248 = ( (~ n3851) ) | ( (~ n4822) ) ;
 assign n2247 = ( (~ n179)  &  n2069 ) | ( n2069  &  n2248 ) ;
 assign n2249 = ( n2069  &  n2068 ) | ( n2069  &  n2248 ) ;
 assign n2251 = ( n153  &  n2249 ) ;
 assign n2250 = ( n18  &  n2094 ) | ( n2094  &  n2251 ) ;
 assign n2253 = ( (~ n3852) ) | ( (~ n4822) ) ;
 assign n2252 = ( (~ n179)  &  n2069 ) | ( n2069  &  n2253 ) ;
 assign n2254 = ( n2069  &  n2068 ) | ( n2069  &  n2253 ) ;
 assign n2256 = ( n153  &  n2254 ) ;
 assign n2255 = ( n18  &  n2094 ) | ( n2094  &  n2256 ) ;
 assign n2257 = ( n2086  &  n2196 ) | ( (~ n2087)  &  n2196 ) ;
 assign n2259 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2257) ) ;
 assign n2261 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2257) ) ;
 assign n2263 = ( n153  &  n2261 ) ;
 assign n2262 = ( n18  &  n2094 ) | ( n2094  &  n2263 ) ;
 assign n2264 = ( n2086  &  n2205 ) | ( (~ n2087)  &  n2205 ) ;
 assign n2265 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2264) ) ;
 assign n2267 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2264) ) ;
 assign n2269 = ( n153  &  n2267 ) ;
 assign n2268 = ( n18  &  n2094 ) | ( n2094  &  n2269 ) ;
 assign n2272 = ( n4378  &  n2444 ) | ( n3776  &  n2444 ) | ( n4378  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n2273 = ( n2070  &  n2447 ) | ( n2070  &  n310 ) ;
 assign n2271 = ( n2247  &  n2250 ) ;
 assign n2270 = ( n2272  &  n2273  &  n2271 ) | ( n2272  &  n2273  &  n891 ) ;
 assign n2275 = ( (~ n3854) ) | ( (~ n4822) ) ;
 assign n2274 = ( (~ n179)  &  n2069 ) | ( n2069  &  n2275 ) ;
 assign n2276 = ( n2069  &  n2068 ) | ( n2069  &  n2275 ) ;
 assign n2278 = ( n153  &  n2276 ) ;
 assign n2277 = ( n18  &  n2094 ) | ( n2094  &  n2278 ) ;
 assign n2280 = ( (~ n3855) ) | ( (~ n4822) ) ;
 assign n2279 = ( (~ n179)  &  n2069 ) | ( n2069  &  n2280 ) ;
 assign n2281 = ( n2069  &  n2068 ) | ( n2069  &  n2280 ) ;
 assign n2283 = ( n153  &  n2281 ) ;
 assign n2282 = ( n18  &  n2094 ) | ( n2094  &  n2283 ) ;
 assign n2284 = ( n2086  &  n2227 ) | ( (~ n2087)  &  n2227 ) ;
 assign n2285 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2284) ) ;
 assign n2287 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2284) ) ;
 assign n2289 = ( n153  &  n2287 ) ;
 assign n2288 = ( n18  &  n2094 ) | ( n2094  &  n2289 ) ;
 assign n2290 = ( n2086  &  n2235 ) | ( (~ n2087)  &  n2235 ) ;
 assign n2291 = ( (~ n179)  &  n2069 ) | ( n2069  &  (~ n2290) ) ;
 assign n2293 = ( n2069  &  n2068 ) | ( n2069  &  (~ n2290) ) ;
 assign n2295 = ( n153  &  n2293 ) ;
 assign n2294 = ( n18  &  n2094 ) | ( n2094  &  n2295 ) ;
 assign n2298 = ( n4381  &  n2433 ) | ( n3776  &  n2433 ) | ( n4381  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n2299 = ( n2070  &  n2436 ) | ( n2070  &  n310 ) ;
 assign n2297 = ( n2274  &  n2277 ) ;
 assign n2296 = ( n2298  &  n2299  &  n2297 ) | ( n2298  &  n2299  &  n891 ) ;
 assign n2302 = ( n2325  &  n2070 ) ;
 assign n2300 = ( n931  &  n934 ) | ( n931  &  n2302 ) | ( n934  &  (~ n3900) ) | ( n2302  &  (~ n3900) ) ;
 assign n2303 = ( (~ Pi27)  &  n176  &  n2069 ) | ( (~ Ni32)  &  n176  &  n2069 ) ;
 assign n2306 = ( Pi22  &  n4730 ) | ( (~ Pi21)  &  n4730 ) | ( n3677  &  n4730 ) ;
 assign n2305 = ( (~ Pi26)  &  n3672 ) | ( n2754  &  n3672 ) ;
 assign n2304 = ( n2306  &  n2305 ) | ( n2306  &  n1866 ) ;
 assign n2307 = ( Pi27  &  n176  &  n2069 ) | ( (~ Ni32)  &  n176  &  n2069 ) ;
 assign n2310 = ( (~ Pi21)  &  n2307 ) | ( Pi21  &  (~ n3901) ) | ( n2307  &  (~ n3901) ) ;
 assign n2309 = ( n3668  &  Pi27 ) | ( n3668  &  n2754 ) ;
 assign n2308 = ( n2310  &  n2309 ) | ( n2310  &  n1866 ) ;
 assign n2313 = ( n2302  &  n2308 ) | ( n940  &  n2308 ) | ( n2302  &  n3525 ) | ( n940  &  n3525 ) ;
 assign n2312 = ( (~ Ni12) ) | ( n3798 ) ;
 assign n2311 = ( n2300  &  n2313  &  n2304 ) | ( n2300  &  n2313  &  n2312 ) ;
 assign n2316 = ( Pi22  &  (~ n4735) ) | ( (~ Pi21)  &  (~ n4735) ) | ( n3682  &  (~ n4735) ) ;
 assign n2315 = ( n3672  &  Pi26 ) | ( n3672  &  n2754 ) ;
 assign n2314 = ( n2316  &  n2315 ) | ( n2316  &  n1866 ) ;
 assign n2317 = ( (~ Pi24)  &  Pi21  &  (~ n2071) ) | ( Pi21  &  (~ n194)  &  (~ n2071) ) ;
 assign n2323 = ( Pi21 ) | ( n3678 ) ;
 assign n2321 = ( Pi24  &  (~ n2317)  &  n2323 ) | ( n2073  &  (~ n2317)  &  n2323 ) ;
 assign n2326 = ( n3681 ) | ( n1866 ) ;
 assign n2325 = ( n2754 ) | ( n1866 ) ;
 assign n2324 = ( n2326  &  n2321  &  Pi24 ) | ( n2326  &  n2321  &  n2325 ) ;
 assign n2328 = ( Pi22 ) | ( (~ Pi21) ) ;
 assign n2327 = ( n2326  &  n2323  &  n194 ) | ( n2326  &  n2323  &  n2328 ) ;
 assign n2331 = ( n3679 ) | ( n2328 ) ;
 assign n2332 = ( (~ Pi27)  &  n2333 ) | ( n2333  &  n3678 ) ;
 assign n2330 = ( (~ Pi27)  &  n3680 ) | ( n3680  &  n3681 ) ;
 assign n2329 = ( n2331  &  n2332  &  n2330 ) | ( n2331  &  n2332  &  n1866 ) ;
 assign n2333 = ( n2069  &  n178 ) ;
 assign n2335 = ( n2456  &  n3798 ) | ( n3798  &  (~ n3914) ) | ( n2456  &  (~ n3916) ) | ( (~ n3914)  &  (~ n3916) ) ;
 assign n2334 = ( n2324  &  n2335 ) | ( n2335  &  (~ Ni13) ) ;
 assign n2336 = ( n18  &  n196  &  n2156 ) | ( n196  &  n2156  &  n2158 ) ;
 assign n2337 = ( n18  &  n196  &  n2176 ) | ( n196  &  n2176  &  n2178 ) ;
 assign n2338 = ( n18  &  n196  &  n2259 ) | ( n196  &  n2259  &  n2261 ) ;
 assign n2339 = ( n18  &  n196  &  n2265 ) | ( n196  &  n2265  &  n2267 ) ;
 assign n2340 = ( n18  &  n196  &  n2247 ) | ( n196  &  n2247  &  n2249 ) ;
 assign n2341 = ( n18  &  n196  &  n2252 ) | ( n196  &  n2252  &  n2254 ) ;
 assign n2342 = ( n18  &  n196  &  n2145 ) | ( n196  &  n2145  &  n2147 ) ;
 assign n2343 = ( n18  &  n196  &  n2151 ) | ( n196  &  n2151  &  n2153 ) ;
 assign n2344 = ( n18  &  n196  &  n2285 ) | ( n196  &  n2285  &  n2287 ) ;
 assign n2345 = ( n18  &  n196  &  n2291 ) | ( n196  &  n2291  &  n2293 ) ;
 assign n2346 = ( n18  &  n196  &  n2274 ) | ( n196  &  n2274  &  n2276 ) ;
 assign n2347 = ( n18  &  n196  &  n2279 ) | ( n196  &  n2279  &  n2281 ) ;
 assign n2348 = ( n18  &  n196  &  n2165 ) | ( n196  &  n2165  &  n2167 ) ;
 assign n2349 = ( n18  &  n196  &  n2171 ) | ( n196  &  n2171  &  n2173 ) ;
 assign n2351 = ( n2156  &  n2159 ) ;
 assign n2352 = ( n2176  &  n2179 ) ;
 assign n2350 = ( n2351  &  n2352 ) | ( n996  &  n2352 ) | ( n2351  &  n998 ) | ( n996  &  n998 ) ;
 assign n2353 = ( (~ n3579)  &  (~ n4523) ) | ( (~ n3579)  &  (~ n4524) ) ;
 assign n2356 = ( (~ n1884)  &  (~ n4525) ) | ( (~ n1884)  &  (~ n4526) ) ;
 assign n2360 = ( n2321  &  n3576 ) | ( n2321  &  n4532  &  n4531 ) ;
 assign n2361 = ( n4536  &  n3582 ) | ( n4536  &  n4530  &  n4529 ) ;
 assign n2362 = ( n4533  &  n4534  &  Pi24 ) | ( n4533  &  n4534  &  n2350 ) ;
 assign n2359 = ( n2360  &  n2361  &  n2362 ) ;
 assign n2363 = ( n18  &  n196  &  n2109 ) | ( n196  &  n2109  &  n2111 ) ;
 assign n2364 = ( n18  &  n196  &  n2135 ) | ( n196  &  n2135  &  n2137 ) ;
 assign n2365 = ( n18  &  n196  &  n2200 ) | ( n196  &  n2200  &  n2202 ) ;
 assign n2366 = ( n18  &  n196  &  n2208 ) | ( n196  &  n2208  &  n2210 ) ;
 assign n2367 = ( n18  &  n196  &  n2185 ) | ( n196  &  n2185  &  n2187 ) ;
 assign n2368 = ( n18  &  n196  &  n2191 ) | ( n196  &  n2191  &  n2193 ) ;
 assign n2369 = ( n18  &  n196  &  n2088 ) | ( n196  &  n2088  &  n2091 ) ;
 assign n2370 = ( n18  &  n196  &  n2101 ) | ( n196  &  n2101  &  n2103 ) ;
 assign n2371 = ( n18  &  n196  &  n2230 ) | ( n196  &  n2230  &  n2232 ) ;
 assign n2372 = ( n18  &  n196  &  n2238 ) | ( n196  &  n2238  &  n2240 ) ;
 assign n2373 = ( n18  &  n196  &  n2217 ) | ( n196  &  n2217  &  n2219 ) ;
 assign n2374 = ( n18  &  n196  &  n2222 ) | ( n196  &  n2222  &  n2224 ) ;
 assign n2375 = ( n18  &  n196  &  n2120 ) | ( n196  &  n2120  &  n2122 ) ;
 assign n2376 = ( n18  &  n196  &  n2128 ) | ( n196  &  n2128  &  n2130 ) ;
 assign n2378 = ( n2109  &  n2112 ) ;
 assign n2379 = ( n2135  &  n2138 ) ;
 assign n2377 = ( n2378  &  n2379 ) | ( n996  &  n2379 ) | ( n2378  &  n998 ) | ( n996  &  n998 ) ;
 assign n2380 = ( (~ n3579)  &  (~ n4503) ) | ( (~ n3579)  &  (~ n4504) ) ;
 assign n2383 = ( (~ n1884)  &  (~ n4505) ) | ( (~ n1884)  &  (~ n4506) ) ;
 assign n2386 = ( (~ n3831)  &  (~ n4516) ) | ( (~ n3831)  &  (~ n4519) ) | ( (~ n3831)  &  (~ n4520) ) ;
 assign n2391 = ( n2324  &  (~ n2386) ) | ( n934  &  n1069  &  (~ n2386) ) ;
 assign n2392 = ( n2334  &  n3499 ) | ( n3499  &  n3805 ) | ( n2334  &  (~ n3918) ) | ( n3805  &  (~ n3918) ) ;
 assign n2390 = ( n2391  &  n2392  &  n2359 ) | ( n2391  &  n2392  &  n1993 ) ;
 assign n2393 = ( Pi21  &  n160  &  (~ n2071) ) | ( Pi21  &  (~ n194)  &  (~ n2071) ) ;
 assign n2394 = ( (~ n160)  &  n2323  &  (~ n2393) ) | ( n2073  &  n2323  &  (~ n2393) ) ;
 assign n2396 = ( (~ n160)  &  n2326  &  n2394 ) | ( n2326  &  n2325  &  n2394 ) ;
 assign n2397 = ( (~ n2328)  &  (~ n4476) ) | ( Pi24  &  (~ n2328)  &  (~ n3677) ) ;
 assign n2401 = ( (~ n1866)  &  (~ n4477) ) | ( Pi24  &  (~ n1866)  &  (~ n2305) ) ;
 assign n2404 = ( (~ Pi21)  &  (~ n4478) ) | ( Pi24  &  (~ Pi21)  &  (~ n3674) ) ;
 assign n2407 = ( n1069  &  n1068 ) | ( n1069  &  (~ n2456) ) ;
 assign n2412 = ( n4491  &  n4371 ) | ( n4491  &  n3823 ) ;
 assign n2410 = ( n2238  &  n2241 ) ;
 assign n2411 = ( (~ n160) ) | ( n3729 ) ;
 assign n2409 = ( n2394  &  n2412  &  n2410 ) | ( n2394  &  n2412  &  n2411 ) ;
 assign n2415 = ( n4490  &  n2244 ) | ( n4490  &  n3823 ) ;
 assign n2414 = ( n2222  &  n2225 ) ;
 assign n2413 = ( n2394  &  n2415  &  n2414 ) | ( n2394  &  n2415  &  n2411 ) ;
 assign n2417 = ( n4489  &  n4365 ) | ( n4489  &  n3823 ) ;
 assign n2416 = ( n2394  &  n2417  &  n2141 ) | ( n2394  &  n2417  &  n2411 ) ;
 assign n2419 = ( n2416  &  n2413 ) | ( n3735  &  n2413 ) | ( n2416  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2420 = ( n4492  &  n2379 ) | ( n4492  &  n3821 ) ;
 assign n2418 = ( n2419  &  n2420  &  n2409 ) | ( n2419  &  n2420  &  n796 ) ;
 assign n2423 = ( n4482  &  n4368 ) | ( n4482  &  n3823 ) ;
 assign n2422 = ( n2208  &  n2211 ) ;
 assign n2421 = ( n2394  &  n2423  &  n2422 ) | ( n2394  &  n2423  &  n2411 ) ;
 assign n2426 = ( n4481  &  n2214 ) | ( n4481  &  n3823 ) ;
 assign n2425 = ( n2191  &  n2194 ) ;
 assign n2424 = ( n2394  &  n2426  &  n2425 ) | ( n2394  &  n2426  &  n2411 ) ;
 assign n2428 = ( n4480  &  n4363 ) | ( n4480  &  n3823 ) ;
 assign n2427 = ( n2394  &  n2428  &  n2115 ) | ( n2394  &  n2428  &  n2411 ) ;
 assign n2430 = ( n2427  &  n2424 ) | ( n3735  &  n2424 ) | ( n2427  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2431 = ( n4483  &  n2378 ) | ( n4483  &  n3821 ) ;
 assign n2429 = ( n2430  &  n2431  &  n2421 ) | ( n2430  &  n2431  &  n796 ) ;
 assign n2434 = ( n4495  &  n4381 ) | ( n4495  &  n3823 ) ;
 assign n2433 = ( n2291  &  n2294 ) ;
 assign n2432 = ( n2394  &  n2434  &  n2433 ) | ( n2394  &  n2434  &  n2411 ) ;
 assign n2437 = ( n4494  &  n2297 ) | ( n4494  &  n3823 ) ;
 assign n2436 = ( n2279  &  n2282 ) ;
 assign n2435 = ( n2394  &  n2437  &  n2436 ) | ( n2394  &  n2437  &  n2411 ) ;
 assign n2439 = ( n4493  &  n4375 ) | ( n4493  &  n3823 ) ;
 assign n2438 = ( n2394  &  n2439  &  n2182 ) | ( n2394  &  n2439  &  n2411 ) ;
 assign n2441 = ( n2438  &  n2435 ) | ( n3735  &  n2435 ) | ( n2438  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2442 = ( n4496  &  n4484  &  n2352 ) | ( n4496  &  n4484  &  n3821 ) ;
 assign n2440 = ( n2441  &  n2442  &  n2432 ) | ( n2441  &  n2442  &  n796 ) ;
 assign n2445 = ( n4487  &  n4378 ) | ( n4487  &  n3823 ) ;
 assign n2444 = ( n2265  &  n2268 ) ;
 assign n2443 = ( n2394  &  n2445  &  n2444 ) | ( n2394  &  n2445  &  n2411 ) ;
 assign n2448 = ( n4486  &  n2271 ) | ( n4486  &  n3823 ) ;
 assign n2447 = ( n2252  &  n2255 ) ;
 assign n2446 = ( n2394  &  n2448  &  n2447 ) | ( n2394  &  n2448  &  n2411 ) ;
 assign n2450 = ( n4485  &  n4373 ) | ( n4485  &  n3823 ) ;
 assign n2449 = ( n2394  &  n2450  &  n2162 ) | ( n2394  &  n2450  &  n2411 ) ;
 assign n2452 = ( n2449  &  n2446 ) | ( n3735  &  n2446 ) | ( n2449  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2453 = ( n4488  &  n2351 ) | ( n4488  &  n3821 ) ;
 assign n2451 = ( n2452  &  n2453  &  n2443 ) | ( n2452  &  n2453  &  n796 ) ;
 assign n2456 = ( (~ Ni14) ) | ( Ni13 ) ;
 assign n2454 = ( n1074  &  (~ n2314)  &  (~ n2396) ) | ( n1074  &  (~ n2396)  &  n2456 ) ;
 assign n2458 = ( (~ n3805)  &  (~ n4479) ) | ( (~ n2396)  &  Ni13  &  (~ n3805) ) ;
 assign n2461 = ( Pi21  &  n168  &  (~ n2071) ) | ( Pi21  &  (~ n194)  &  (~ n2071) ) ;
 assign n2462 = ( (~ n168)  &  n2323  &  (~ n2461) ) | ( n2073  &  n2323  &  (~ n2461) ) ;
 assign n2464 = ( (~ n168)  &  n2326  &  n2462 ) | ( n2326  &  n2325  &  n2462 ) ;
 assign n2467 = ( n4551  &  n4371 ) | ( n4551  &  n3835 ) ;
 assign n2466 = ( (~ n168) ) | ( n3729 ) ;
 assign n2465 = ( n2462  &  n2467  &  n2410 ) | ( n2462  &  n2467  &  n2466 ) ;
 assign n2469 = ( n4550  &  n2244 ) | ( n4550  &  n3835 ) ;
 assign n2468 = ( n2462  &  n2469  &  n2414 ) | ( n2462  &  n2469  &  n2466 ) ;
 assign n2471 = ( n4549  &  n4365 ) | ( n4549  &  n3835 ) ;
 assign n2470 = ( n2462  &  n2471  &  n2141 ) | ( n2462  &  n2471  &  n2466 ) ;
 assign n2473 = ( n2470  &  n2468 ) | ( n3735  &  n2468 ) | ( n2470  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2474 = ( n4552  &  n2379 ) | ( n4552  &  n3833 ) ;
 assign n2472 = ( n2473  &  n2474  &  n2465 ) | ( n2473  &  n2474  &  n796 ) ;
 assign n2476 = ( n4542  &  n4368 ) | ( n4542  &  n3835 ) ;
 assign n2475 = ( n2462  &  n2476  &  n2422 ) | ( n2462  &  n2476  &  n2466 ) ;
 assign n2478 = ( n4541  &  n2214 ) | ( n4541  &  n3835 ) ;
 assign n2477 = ( n2462  &  n2478  &  n2425 ) | ( n2462  &  n2478  &  n2466 ) ;
 assign n2480 = ( n4540  &  n4363 ) | ( n4540  &  n3835 ) ;
 assign n2479 = ( n2462  &  n2480  &  n2115 ) | ( n2462  &  n2480  &  n2466 ) ;
 assign n2482 = ( n2479  &  n2477 ) | ( n3735  &  n2477 ) | ( n2479  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2483 = ( n4543  &  n2378 ) | ( n4543  &  n3833 ) ;
 assign n2481 = ( n2482  &  n2483  &  n2475 ) | ( n2482  &  n2483  &  n796 ) ;
 assign n2485 = ( n4555  &  n4381 ) | ( n4555  &  n3835 ) ;
 assign n2484 = ( n2462  &  n2485  &  n2433 ) | ( n2462  &  n2485  &  n2466 ) ;
 assign n2487 = ( n4554  &  n2297 ) | ( n4554  &  n3835 ) ;
 assign n2486 = ( n2462  &  n2487  &  n2436 ) | ( n2462  &  n2487  &  n2466 ) ;
 assign n2489 = ( n4553  &  n4375 ) | ( n4553  &  n3835 ) ;
 assign n2488 = ( n2462  &  n2489  &  n2182 ) | ( n2462  &  n2489  &  n2466 ) ;
 assign n2491 = ( n2488  &  n2486 ) | ( n3735  &  n2486 ) | ( n2488  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2492 = ( n4556  &  n4544  &  n2352 ) | ( n4556  &  n4544  &  n3833 ) ;
 assign n2490 = ( n2491  &  n2492  &  n2484 ) | ( n2491  &  n2492  &  n796 ) ;
 assign n2494 = ( n4547  &  n4378 ) | ( n4547  &  n3835 ) ;
 assign n2493 = ( n2462  &  n2494  &  n2444 ) | ( n2462  &  n2494  &  n2466 ) ;
 assign n2496 = ( n4546  &  n2271 ) | ( n4546  &  n3835 ) ;
 assign n2495 = ( n2462  &  n2496  &  n2447 ) | ( n2462  &  n2496  &  n2466 ) ;
 assign n2498 = ( n4545  &  n4373 ) | ( n4545  &  n3835 ) ;
 assign n2497 = ( n2462  &  n2498  &  n2162 ) | ( n2462  &  n2498  &  n2466 ) ;
 assign n2500 = ( n2497  &  n2495 ) | ( n3735  &  n2495 ) | ( n2497  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2501 = ( n4548  &  n2351 ) | ( n4548  &  n3833 ) ;
 assign n2499 = ( n2500  &  n2501  &  n2493 ) | ( n2500  &  n2501  &  n796 ) ;
 assign n2502 = ( n1074  &  (~ n2314)  &  (~ n2464) ) | ( n1074  &  n2456  &  (~ n2464) ) ;
 assign n2504 = ( (~ n3805)  &  (~ n4539) ) | ( Ni13  &  (~ n2464)  &  (~ n3805) ) ;
 assign n2506 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2085) ) ;
 assign n2508 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2100) ) ;
 assign n2509 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2107) ) ;
 assign n2512 = ( n4355  &  n2629 ) | ( n1250  &  n2629 ) | ( n4355  &  n891 ) | ( n1250  &  n891 ) ;
 assign n2511 = ( n2508  &  n2104 ) ;
 assign n2510 = ( n2070  &  n2512  &  n2511 ) | ( n2070  &  n2512  &  n310 ) ;
 assign n2513 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2119) ) ;
 assign n2514 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2127) ) ;
 assign n2515 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2133) ) ;
 assign n2518 = ( n4357  &  n2601 ) | ( n1250  &  n2601 ) | ( n4357  &  n891 ) | ( n1250  &  n891 ) ;
 assign n2517 = ( n2514  &  n2131 ) ;
 assign n2516 = ( n2070  &  n2518  &  n2517 ) | ( n2070  &  n2518  &  n310 ) ;
 assign n2519 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2143) ) ;
 assign n2520 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2150) ) ;
 assign n2521 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2108) ) ;
 assign n2524 = ( n4356  &  n2685 ) | ( n1250  &  n2685 ) | ( n4356  &  n891 ) | ( n1250  &  n891 ) ;
 assign n2523 = ( n2520  &  n2154 ) ;
 assign n2522 = ( n2070  &  n2524  &  n2523 ) | ( n2070  &  n2524  &  n310 ) ;
 assign n2525 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2164) ) ;
 assign n2526 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2170) ) ;
 assign n2527 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2134) ) ;
 assign n2530 = ( n4358  &  n2657 ) | ( n1250  &  n2657 ) | ( n4358  &  n891 ) | ( n1250  &  n891 ) ;
 assign n2529 = ( n2526  &  n2174 ) ;
 assign n2528 = ( n2070  &  n2530  &  n2529 ) | ( n2070  &  n2530  &  n310 ) ;
 assign n2531 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n3851) ) ;
 assign n2532 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n3852) ) ;
 assign n2533 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2198) ) ;
 assign n2534 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2207) ) ;
 assign n2537 = ( n2614  &  n4345 ) | ( n3776  &  n4345 ) | ( n2614  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n2538 = ( n2070  &  n4346 ) | ( n2070  &  n310 ) ;
 assign n2536 = ( n2531  &  n2188 ) ;
 assign n2535 = ( n2537  &  n2538  &  n2536 ) | ( n2537  &  n2538  &  n891 ) ;
 assign n2539 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n3854) ) ;
 assign n2540 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n3855) ) ;
 assign n2541 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2229) ) ;
 assign n2542 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2237) ) ;
 assign n2545 = ( n2586  &  n4349 ) | ( n3776  &  n4349 ) | ( n2586  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n2546 = ( n2070  &  n4350 ) | ( n2070  &  n310 ) ;
 assign n2544 = ( n2539  &  n2220 ) ;
 assign n2543 = ( n2545  &  n2546  &  n2544 ) | ( n2545  &  n2546  &  n891 ) ;
 assign n2547 = ( (~ n183)  &  n2069 ) | ( n2069  &  n2248 ) ;
 assign n2548 = ( (~ n183)  &  n2069 ) | ( n2069  &  n2253 ) ;
 assign n2549 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2257) ) ;
 assign n2550 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2264) ) ;
 assign n2553 = ( n2670  &  n4347 ) | ( n3776  &  n4347 ) | ( n2670  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n2554 = ( n2070  &  n4348 ) | ( n2070  &  n310 ) ;
 assign n2552 = ( n2547  &  n2250 ) ;
 assign n2551 = ( n2553  &  n2554  &  n2552 ) | ( n2553  &  n2554  &  n891 ) ;
 assign n2555 = ( (~ n183)  &  n2069 ) | ( n2069  &  n2275 ) ;
 assign n2556 = ( (~ n183)  &  n2069 ) | ( n2069  &  n2280 ) ;
 assign n2557 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2284) ) ;
 assign n2558 = ( (~ n183)  &  n2069 ) | ( n2069  &  (~ n2290) ) ;
 assign n2561 = ( n2642  &  n4351 ) | ( n3776  &  n4351 ) | ( n2642  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n2562 = ( n2070  &  n4352 ) | ( n2070  &  n310 ) ;
 assign n2560 = ( n2555  &  n2277 ) ;
 assign n2559 = ( n2561  &  n2562  &  n2560 ) | ( n2561  &  n2562  &  n891 ) ;
 assign n2564 = ( (~ Pi20)  &  n2093 ) | ( Pi20  &  n2105 ) | ( n2093  &  n2105 ) ;
 assign n2563 = ( n2564  &  n2113 ) | ( n1249  &  n2113 ) | ( n2564  &  n1250 ) | ( n1249  &  n1250 ) ;
 assign n2566 = ( (~ Pi20)  &  n2124 ) | ( Pi20  &  n2132 ) | ( n2124  &  n2132 ) ;
 assign n2565 = ( n2566  &  n2139 ) | ( n1249  &  n2139 ) | ( n2566  &  n1250 ) | ( n1249  &  n1250 ) ;
 assign n2568 = ( (~ Pi20)  &  n2169 ) | ( Pi20  &  n2175 ) | ( n2169  &  n2175 ) ;
 assign n2567 = ( n2568  &  n2180 ) | ( n1249  &  n2180 ) | ( n2568  &  n1250 ) | ( n1249  &  n1250 ) ;
 assign n2570 = ( (~ Pi20)  &  n2189 ) | ( Pi20  &  n2195 ) | ( n2189  &  n2195 ) ;
 assign n2571 = ( (~ Pi20)  &  n2204 ) | ( Pi20  &  n2212 ) | ( n2204  &  n2212 ) ;
 assign n2569 = ( n2570  &  n2571 ) | ( n1249  &  n2571 ) | ( n2570  &  n1250 ) | ( n1249  &  n1250 ) ;
 assign n2573 = ( (~ Pi20)  &  n2221 ) | ( Pi20  &  n2226 ) | ( n2221  &  n2226 ) ;
 assign n2574 = ( (~ Pi20)  &  n2234 ) | ( Pi20  &  n2242 ) | ( n2234  &  n2242 ) ;
 assign n2572 = ( n2573  &  n2574 ) | ( n1249  &  n2574 ) | ( n2573  &  n1250 ) | ( n1249  &  n1250 ) ;
 assign n2576 = ( (~ Pi20)  &  n2278 ) | ( Pi20  &  n2283 ) | ( n2278  &  n2283 ) ;
 assign n2577 = ( (~ Pi20)  &  n2289 ) | ( Pi20  &  n2295 ) | ( n2289  &  n2295 ) ;
 assign n2575 = ( n2576  &  n2577 ) | ( n1249  &  n2577 ) | ( n2576  &  n1250 ) | ( n1249  &  n1250 ) ;
 assign n2580 = ( n4752 ) | ( n4753 ) | ( n931 ) ;
 assign n2579 = ( Pi17  &  (~ n4750) ) | ( n4353  &  n4354  &  (~ n4750) ) ;
 assign n2578 = ( n2580  &  n2579 ) | ( n2580  &  n934 ) ;
 assign n2582 = ( n176  &  n2232 ) ;
 assign n2581 = ( n18  &  n176  &  n2541 ) | ( n176  &  n2541  &  n2582 ) ;
 assign n2584 = ( n176  &  n2240 ) ;
 assign n2583 = ( n18  &  n176  &  n2542 ) | ( n176  &  n2542  &  n2584 ) ;
 assign n2587 = ( n2581  &  n2583 ) | ( n3801  &  n2583 ) | ( n2581  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n2588 = ( n2306  &  n4349 ) | ( n2306  &  n3803 ) ;
 assign n2586 = ( n2541  &  n2233 ) ;
 assign n2585 = ( n2587  &  n2588  &  n2586 ) | ( n2587  &  n2588  &  n1275 ) ;
 assign n2590 = ( n176  &  n2219 ) ;
 assign n2589 = ( n18  &  n176  &  n2539 ) | ( n176  &  n2539  &  n2590 ) ;
 assign n2592 = ( n176  &  n2224 ) ;
 assign n2591 = ( n18  &  n176  &  n2540 ) | ( n176  &  n2540  &  n2592 ) ;
 assign n2594 = ( n2589  &  n2591 ) | ( n3801  &  n2591 ) | ( n2589  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n2595 = ( n2306  &  n4350 ) | ( n2306  &  n3803 ) ;
 assign n2593 = ( n2594  &  n2595  &  n2544 ) | ( n2594  &  n2595  &  n1275 ) ;
 assign n2597 = ( n176  &  n2122 ) ;
 assign n2596 = ( n18  &  n176  &  n2513 ) | ( n176  &  n2513  &  n2597 ) ;
 assign n2599 = ( n176  &  n2130 ) ;
 assign n2598 = ( n18  &  n176  &  n2514 ) | ( n176  &  n2514  &  n2599 ) ;
 assign n2602 = ( n2596  &  n2598 ) | ( n3801  &  n2598 ) | ( n2596  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n2603 = ( n2306  &  n2517 ) | ( n2306  &  n3803 ) ;
 assign n2601 = ( n2513  &  n2123 ) ;
 assign n2600 = ( n2602  &  n2603  &  n2601 ) | ( n2602  &  n2603  &  n1275 ) ;
 assign n2605 = ( n176  &  n2137 ) ;
 assign n2604 = ( n18  &  n176  &  n2515 ) | ( n176  &  n2515  &  n2605 ) ;
 assign n2607 = ( n2600  &  n2593 ) | ( n3735  &  n2593 ) | ( n2600  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2608 = ( n4471  &  n4469  &  n4357 ) | ( n4471  &  n4469  &  n3800 ) ;
 assign n2606 = ( n2607  &  n2608  &  n2585 ) | ( n2607  &  n2608  &  n796 ) ;
 assign n2610 = ( n176  &  n2202 ) ;
 assign n2609 = ( n18  &  n176  &  n2533 ) | ( n176  &  n2533  &  n2610 ) ;
 assign n2612 = ( n176  &  n2210 ) ;
 assign n2611 = ( n18  &  n176  &  n2534 ) | ( n176  &  n2534  &  n2612 ) ;
 assign n2615 = ( n2609  &  n2611 ) | ( n3801  &  n2611 ) | ( n2609  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n2616 = ( n2306  &  n4345 ) | ( n2306  &  n3803 ) ;
 assign n2614 = ( n2533  &  n2203 ) ;
 assign n2613 = ( n2615  &  n2616  &  n2614 ) | ( n2615  &  n2616  &  n1275 ) ;
 assign n2618 = ( n176  &  n2187 ) ;
 assign n2617 = ( n18  &  n176  &  n2531 ) | ( n176  &  n2531  &  n2618 ) ;
 assign n2620 = ( n176  &  n2193 ) ;
 assign n2619 = ( n18  &  n176  &  n2532 ) | ( n176  &  n2532  &  n2620 ) ;
 assign n2622 = ( n2617  &  n2619 ) | ( n3801  &  n2619 ) | ( n2617  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n2623 = ( n2306  &  n4346 ) | ( n2306  &  n3803 ) ;
 assign n2621 = ( n2622  &  n2623  &  n2536 ) | ( n2622  &  n2623  &  n1275 ) ;
 assign n2625 = ( n176  &  n2091 ) ;
 assign n2624 = ( n18  &  n176  &  n2506 ) | ( n176  &  n2506  &  n2625 ) ;
 assign n2627 = ( n176  &  n2103 ) ;
 assign n2626 = ( n18  &  n176  &  n2508 ) | ( n176  &  n2508  &  n2627 ) ;
 assign n2630 = ( n2624  &  n2626 ) | ( n3801  &  n2626 ) | ( n2624  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n2631 = ( n2306  &  n2511 ) | ( n2306  &  n3803 ) ;
 assign n2629 = ( n2506  &  n2092 ) ;
 assign n2628 = ( n2630  &  n2631  &  n2629 ) | ( n2630  &  n2631  &  n1275 ) ;
 assign n2633 = ( n176  &  n2111 ) ;
 assign n2632 = ( n18  &  n176  &  n2509 ) | ( n176  &  n2509  &  n2633 ) ;
 assign n2635 = ( n2628  &  n2621 ) | ( n3735  &  n2621 ) | ( n2628  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2636 = ( n4468  &  n4469  &  n4355 ) | ( n4468  &  n4469  &  n3800 ) ;
 assign n2634 = ( n2635  &  n2636  &  n2613 ) | ( n2635  &  n2636  &  n796 ) ;
 assign n2638 = ( n176  &  n2287 ) ;
 assign n2637 = ( n18  &  n176  &  n2557 ) | ( n176  &  n2557  &  n2638 ) ;
 assign n2640 = ( n176  &  n2293 ) ;
 assign n2639 = ( n18  &  n176  &  n2558 ) | ( n176  &  n2558  &  n2640 ) ;
 assign n2643 = ( n2637  &  n2639 ) | ( n3801  &  n2639 ) | ( n2637  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n2644 = ( n2306  &  n4351 ) | ( n2306  &  n3803 ) ;
 assign n2642 = ( n2557  &  n2288 ) ;
 assign n2641 = ( n2643  &  n2644  &  n2642 ) | ( n2643  &  n2644  &  n1275 ) ;
 assign n2646 = ( n176  &  n2276 ) ;
 assign n2645 = ( n18  &  n176  &  n2555 ) | ( n176  &  n2555  &  n2646 ) ;
 assign n2648 = ( n176  &  n2281 ) ;
 assign n2647 = ( n18  &  n176  &  n2556 ) | ( n176  &  n2556  &  n2648 ) ;
 assign n2650 = ( n2645  &  n2647 ) | ( n3801  &  n2647 ) | ( n2645  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n2651 = ( n2306  &  n4352 ) | ( n2306  &  n3803 ) ;
 assign n2649 = ( n2650  &  n2651  &  n2560 ) | ( n2650  &  n2651  &  n1275 ) ;
 assign n2653 = ( n176  &  n2167 ) ;
 assign n2652 = ( n18  &  n176  &  n2525 ) | ( n176  &  n2525  &  n2653 ) ;
 assign n2655 = ( n176  &  n2173 ) ;
 assign n2654 = ( n18  &  n176  &  n2526 ) | ( n176  &  n2526  &  n2655 ) ;
 assign n2658 = ( n2652  &  n2654 ) | ( n3801  &  n2654 ) | ( n2652  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n2659 = ( n2306  &  n2529 ) | ( n2306  &  n3803 ) ;
 assign n2657 = ( n2525  &  n2168 ) ;
 assign n2656 = ( n2658  &  n2659  &  n2657 ) | ( n2658  &  n2659  &  n1275 ) ;
 assign n2661 = ( n176  &  n2178 ) ;
 assign n2660 = ( n18  &  n176  &  n2527 ) | ( n176  &  n2527  &  n2661 ) ;
 assign n2663 = ( n2656  &  n2649 ) | ( n3735  &  n2649 ) | ( n2656  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2664 = ( n4472  &  n4469  &  n4358 ) | ( n4472  &  n4469  &  n3800 ) ;
 assign n2662 = ( n2663  &  n2664  &  n2641 ) | ( n2663  &  n2664  &  n796 ) ;
 assign n2666 = ( n176  &  n2261 ) ;
 assign n2665 = ( n18  &  n176  &  n2549 ) | ( n176  &  n2549  &  n2666 ) ;
 assign n2668 = ( n176  &  n2267 ) ;
 assign n2667 = ( n18  &  n176  &  n2550 ) | ( n176  &  n2550  &  n2668 ) ;
 assign n2671 = ( n2665  &  n2667 ) | ( n3801  &  n2667 ) | ( n2665  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n2672 = ( n2306  &  n4347 ) | ( n2306  &  n3803 ) ;
 assign n2670 = ( n2549  &  n2262 ) ;
 assign n2669 = ( n2671  &  n2672  &  n2670 ) | ( n2671  &  n2672  &  n1275 ) ;
 assign n2674 = ( n176  &  n2249 ) ;
 assign n2673 = ( n18  &  n176  &  n2547 ) | ( n176  &  n2547  &  n2674 ) ;
 assign n2676 = ( n176  &  n2254 ) ;
 assign n2675 = ( n18  &  n176  &  n2548 ) | ( n176  &  n2548  &  n2676 ) ;
 assign n2678 = ( n2673  &  n2675 ) | ( n3801  &  n2675 ) | ( n2673  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n2679 = ( n2306  &  n4348 ) | ( n2306  &  n3803 ) ;
 assign n2677 = ( n2678  &  n2679  &  n2552 ) | ( n2678  &  n2679  &  n1275 ) ;
 assign n2681 = ( n176  &  n2147 ) ;
 assign n2680 = ( n18  &  n176  &  n2519 ) | ( n176  &  n2519  &  n2681 ) ;
 assign n2683 = ( n176  &  n2153 ) ;
 assign n2682 = ( n18  &  n176  &  n2520 ) | ( n176  &  n2520  &  n2683 ) ;
 assign n2686 = ( n2680  &  n2682 ) | ( n3801  &  n2682 ) | ( n2680  &  n3802 ) | ( n3801  &  n3802 ) ;
 assign n2687 = ( n2306  &  n2523 ) | ( n2306  &  n3803 ) ;
 assign n2685 = ( n2519  &  n2148 ) ;
 assign n2684 = ( n2686  &  n2687  &  n2685 ) | ( n2686  &  n2687  &  n1275 ) ;
 assign n2689 = ( n176  &  n2158 ) ;
 assign n2688 = ( n18  &  n176  &  n2521 ) | ( n176  &  n2521  &  n2689 ) ;
 assign n2691 = ( n2684  &  n2677 ) | ( n3735  &  n2677 ) | ( n2684  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2692 = ( n4470  &  n4469  &  n4356 ) | ( n4470  &  n4469  &  n3800 ) ;
 assign n2690 = ( n2691  &  n2692  &  n2669 ) | ( n2691  &  n2692  &  n796 ) ;
 assign n2693 = ( (~ n1884)  &  (~ n4452) ) | ( (~ n1884)  &  (~ n4453) ) ;
 assign n2696 = ( (~ n1884)  &  (~ n4432) ) | ( (~ n1884)  &  (~ n4433) ) ;
 assign n2700 = ( n4746 ) | ( n4748 ) | ( n3525 ) ;
 assign n2701 = ( n2578  &  n2312 ) | ( n2578  &  n4474  &  n4473 ) ;
 assign n2699 = ( n2700  &  n2701  &  n2579 ) | ( n2700  &  n2701  &  n940 ) ;
 assign n2703 = ( n2581  &  n2583 ) | ( n3787  &  n2583 ) | ( n2581  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n2704 = ( n2316  &  n4349 ) | ( n2316  &  n3789 ) ;
 assign n2702 = ( n2703  &  n2704  &  n2586 ) | ( n2703  &  n2704  &  n1418 ) ;
 assign n2706 = ( n2589  &  n2591 ) | ( n3787  &  n2591 ) | ( n2589  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n2707 = ( n2316  &  n4350 ) | ( n2316  &  n3789 ) ;
 assign n2705 = ( n2706  &  n2707  &  n2544 ) | ( n2706  &  n2707  &  n1418 ) ;
 assign n2709 = ( n2596  &  n2598 ) | ( n3787  &  n2598 ) | ( n2596  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n2710 = ( n2316  &  n2517 ) | ( n2316  &  n3789 ) ;
 assign n2708 = ( n2709  &  n2710  &  n2601 ) | ( n2709  &  n2710  &  n1418 ) ;
 assign n2712 = ( n2708  &  n2705 ) | ( n3735  &  n2705 ) | ( n2708  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2713 = ( n4426  &  n4424  &  n4357 ) | ( n4426  &  n4424  &  n3786 ) ;
 assign n2711 = ( n2712  &  n2713  &  n2702 ) | ( n2712  &  n2713  &  n796 ) ;
 assign n2715 = ( n2609  &  n2611 ) | ( n3787  &  n2611 ) | ( n2609  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n2716 = ( n2316  &  n4345 ) | ( n2316  &  n3789 ) ;
 assign n2714 = ( n2715  &  n2716  &  n2614 ) | ( n2715  &  n2716  &  n1418 ) ;
 assign n2718 = ( n2617  &  n2619 ) | ( n3787  &  n2619 ) | ( n2617  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n2719 = ( n2316  &  n4346 ) | ( n2316  &  n3789 ) ;
 assign n2717 = ( n2718  &  n2719  &  n2536 ) | ( n2718  &  n2719  &  n1418 ) ;
 assign n2721 = ( n2624  &  n2626 ) | ( n3787  &  n2626 ) | ( n2624  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n2722 = ( n2316  &  n2511 ) | ( n2316  &  n3789 ) ;
 assign n2720 = ( n2721  &  n2722  &  n2629 ) | ( n2721  &  n2722  &  n1418 ) ;
 assign n2724 = ( n2720  &  n2717 ) | ( n3735  &  n2717 ) | ( n2720  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2725 = ( n4423  &  n4424  &  n4355 ) | ( n4423  &  n4424  &  n3786 ) ;
 assign n2723 = ( n2724  &  n2725  &  n2714 ) | ( n2724  &  n2725  &  n796 ) ;
 assign n2727 = ( n2637  &  n2639 ) | ( n3787  &  n2639 ) | ( n2637  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n2728 = ( n2316  &  n4351 ) | ( n2316  &  n3789 ) ;
 assign n2726 = ( n2727  &  n2728  &  n2642 ) | ( n2727  &  n2728  &  n1418 ) ;
 assign n2730 = ( n2645  &  n2647 ) | ( n3787  &  n2647 ) | ( n2645  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n2731 = ( n2316  &  n4352 ) | ( n2316  &  n3789 ) ;
 assign n2729 = ( n2730  &  n2731  &  n2560 ) | ( n2730  &  n2731  &  n1418 ) ;
 assign n2733 = ( n2652  &  n2654 ) | ( n3787  &  n2654 ) | ( n2652  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n2734 = ( n2316  &  n2529 ) | ( n2316  &  n3789 ) ;
 assign n2732 = ( n2733  &  n2734  &  n2657 ) | ( n2733  &  n2734  &  n1418 ) ;
 assign n2736 = ( n2732  &  n2729 ) | ( n3735  &  n2729 ) | ( n2732  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2737 = ( n4427  &  n4424  &  n4358 ) | ( n4427  &  n4424  &  n3786 ) ;
 assign n2735 = ( n2736  &  n2737  &  n2726 ) | ( n2736  &  n2737  &  n796 ) ;
 assign n2739 = ( n2665  &  n2667 ) | ( n3787  &  n2667 ) | ( n2665  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n2740 = ( n2316  &  n4347 ) | ( n2316  &  n3789 ) ;
 assign n2738 = ( n2739  &  n2740  &  n2670 ) | ( n2739  &  n2740  &  n1418 ) ;
 assign n2742 = ( n2673  &  n2675 ) | ( n3787  &  n2675 ) | ( n2673  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n2743 = ( n2316  &  n4348 ) | ( n2316  &  n3789 ) ;
 assign n2741 = ( n2742  &  n2743  &  n2552 ) | ( n2742  &  n2743  &  n1418 ) ;
 assign n2745 = ( n2680  &  n2682 ) | ( n3787  &  n2682 ) | ( n2680  &  n3788 ) | ( n3787  &  n3788 ) ;
 assign n2746 = ( n2316  &  n2523 ) | ( n2316  &  n3789 ) ;
 assign n2744 = ( n2745  &  n2746  &  n2685 ) | ( n2745  &  n2746  &  n1418 ) ;
 assign n2748 = ( n2744  &  n2741 ) | ( n3735  &  n2741 ) | ( n2744  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2749 = ( n4425  &  n4424  &  n4356 ) | ( n4425  &  n4424  &  n3786 ) ;
 assign n2747 = ( n2748  &  n2749  &  n2738 ) | ( n2748  &  n2749  &  n796 ) ;
 assign n2751 = ( n2711  &  n2735 ) | ( n3763  &  n2735 ) | ( n2711  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n2752 = ( n2723  &  n2747 ) | ( n3742  &  n2747 ) | ( n2723  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n2750 = ( n2751  &  n2752 ) ;
 assign n2754 = ( n153  &  n2074 ) ;
 assign n2753 = ( n2070  &  n2754 ) | ( n2070  &  n1471 ) ;
 assign n2757 = ( n2753  &  n1480 ) | ( n2753  &  n4344  &  n4342 ) ;
 assign n2756 = ( (~ Pi16)  &  n2160 ) | ( n2160  &  n2180 ) ;
 assign n2755 = ( n2757  &  n2756 ) | ( n2757  &  n1474 ) ;
 assign n2760 = ( n2753  &  n1480 ) | ( n2753  &  n4340  &  n4338 ) ;
 assign n2759 = ( (~ Pi16)  &  n2113 ) | ( n2113  &  n2139 ) ;
 assign n2758 = ( n2760  &  n2759 ) | ( n2760  &  n1474 ) ;
 assign n2763 = ( n4373  &  n2162 ) | ( n3728  &  n2162 ) | ( n4373  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n2762 = ( (~ Pi20)  &  n2149 ) | ( Pi20  &  n2155 ) | ( n2149  &  n2155 ) ;
 assign n2761 = ( n2763  &  n2762 ) | ( n2763  &  n1480 ) ;
 assign n2764 = ( (~ n3579)  &  (~ n4374) ) | ( (~ n1480)  &  (~ n2568)  &  (~ n3579) ) ;
 assign n2767 = ( (~ n1884)  &  (~ n4376) ) | ( (~ n1480)  &  (~ n1884)  &  (~ n2832) ) ;
 assign n2770 = ( (~ n3778)  &  (~ n4377) ) | ( (~ n1480)  &  (~ n2829)  &  (~ n3778) ) ;
 assign n2773 = ( (~ n3582)  &  (~ n4379) ) | ( (~ n1480)  &  (~ n2576)  &  (~ n3582) ) ;
 assign n2776 = ( (~ n3576)  &  (~ n4380) ) | ( (~ n1480)  &  (~ n2577)  &  (~ n3576) ) ;
 assign n2781 = ( n4363  &  n2115 ) | ( n3728  &  n2115 ) | ( n4363  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n2780 = ( n2781  &  n2564 ) | ( n2781  &  n1480 ) ;
 assign n2782 = ( (~ n3579)  &  (~ n4364) ) | ( (~ n1480)  &  (~ n2566)  &  (~ n3579) ) ;
 assign n2785 = ( (~ n1884)  &  (~ n4366) ) | ( (~ n1480)  &  (~ n1884)  &  (~ n2570) ) ;
 assign n2788 = ( (~ n3778)  &  (~ n4367) ) | ( (~ n1480)  &  (~ n2571)  &  (~ n3778) ) ;
 assign n2791 = ( (~ n3582)  &  (~ n4369) ) | ( (~ n1480)  &  (~ n2573)  &  (~ n3582) ) ;
 assign n2794 = ( (~ n3576)  &  (~ n4370) ) | ( (~ n1480)  &  (~ n2574)  &  (~ n3576) ) ;
 assign n2799 = ( Pi15  &  n2755 ) | ( (~ Pi15)  &  n2758 ) | ( n2755  &  n2758 ) ;
 assign n2797 = ( n931  &  n934 ) | ( n931  &  n2799 ) | ( n934  &  (~ n3899) ) | ( n2799  &  (~ n3899) ) ;
 assign n2800 = ( n2316  &  n2315 ) | ( n2316  &  n1471 ) ;
 assign n2802 = ( n2582  &  n2584 ) | ( n3817  &  n2584 ) | ( n2582  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n2801 = ( n2800  &  n2802  &  n2574 ) | ( n2800  &  n2802  &  n1525 ) ;
 assign n2804 = ( n2590  &  n2592 ) | ( n3817  &  n2592 ) | ( n2590  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n2803 = ( n2800  &  n2804  &  n2573 ) | ( n2800  &  n2804  &  n1525 ) ;
 assign n2806 = ( n2597  &  n2599 ) | ( n3817  &  n2599 ) | ( n2597  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n2805 = ( n2800  &  n2806  &  n2566 ) | ( n2800  &  n2806  &  n1525 ) ;
 assign n2808 = ( n2805  &  n2803 ) | ( n3735  &  n2803 ) | ( n2805  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2809 = ( n4419  &  n4417  &  n2139 ) | ( n4419  &  n4417  &  n3816 ) ;
 assign n2807 = ( n2808  &  n2809  &  n2801 ) | ( n2808  &  n2809  &  n796 ) ;
 assign n2811 = ( n2610  &  n2612 ) | ( n3817  &  n2612 ) | ( n2610  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n2810 = ( n2800  &  n2811  &  n2571 ) | ( n2800  &  n2811  &  n1525 ) ;
 assign n2813 = ( n2618  &  n2620 ) | ( n3817  &  n2620 ) | ( n2618  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n2812 = ( n2800  &  n2813  &  n2570 ) | ( n2800  &  n2813  &  n1525 ) ;
 assign n2815 = ( n2625  &  n2627 ) | ( n3817  &  n2627 ) | ( n2625  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n2814 = ( n2800  &  n2815  &  n2564 ) | ( n2800  &  n2815  &  n1525 ) ;
 assign n2817 = ( n2814  &  n2812 ) | ( n3735  &  n2812 ) | ( n2814  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2818 = ( n4416  &  n4417  &  n2113 ) | ( n4416  &  n4417  &  n3816 ) ;
 assign n2816 = ( n2817  &  n2818  &  n2810 ) | ( n2817  &  n2818  &  n796 ) ;
 assign n2820 = ( n2638  &  n2640 ) | ( n3817  &  n2640 ) | ( n2638  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n2819 = ( n2800  &  n2820  &  n2577 ) | ( n2800  &  n2820  &  n1525 ) ;
 assign n2822 = ( n2646  &  n2648 ) | ( n3817  &  n2648 ) | ( n2646  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n2821 = ( n2800  &  n2822  &  n2576 ) | ( n2800  &  n2822  &  n1525 ) ;
 assign n2824 = ( n2653  &  n2655 ) | ( n3817  &  n2655 ) | ( n2653  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n2823 = ( n2800  &  n2824  &  n2568 ) | ( n2800  &  n2824  &  n1525 ) ;
 assign n2826 = ( n2823  &  n2821 ) | ( n3735  &  n2821 ) | ( n2823  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2827 = ( n4420  &  n4417  &  n2180 ) | ( n4420  &  n4417  &  n3816 ) ;
 assign n2825 = ( n2826  &  n2827  &  n2819 ) | ( n2826  &  n2827  &  n796 ) ;
 assign n2830 = ( n2666  &  n2668 ) | ( n3817  &  n2668 ) | ( n2666  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n2829 = ( (~ Pi20)  &  n2263 ) | ( Pi20  &  n2269 ) | ( n2263  &  n2269 ) ;
 assign n2828 = ( n2800  &  n2830  &  n2829 ) | ( n2800  &  n2830  &  n1525 ) ;
 assign n2833 = ( n2674  &  n2676 ) | ( n3817  &  n2676 ) | ( n2674  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n2832 = ( (~ Pi20)  &  n2251 ) | ( Pi20  &  n2256 ) | ( n2251  &  n2256 ) ;
 assign n2831 = ( n2800  &  n2833  &  n2832 ) | ( n2800  &  n2833  &  n1525 ) ;
 assign n2835 = ( n2681  &  n2683 ) | ( n3817  &  n2683 ) | ( n2681  &  n3818 ) | ( n3817  &  n3818 ) ;
 assign n2834 = ( n2800  &  n2835  &  n2762 ) | ( n2800  &  n2835  &  n1525 ) ;
 assign n2837 = ( n2834  &  n2831 ) | ( n3735  &  n2831 ) | ( n2834  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2838 = ( n4418  &  n4417  &  n2160 ) | ( n4418  &  n4417  &  n3816 ) ;
 assign n2836 = ( n2837  &  n2838  &  n2828 ) | ( n2837  &  n2838  &  n796 ) ;
 assign n2839 = ( n2310  &  n2309 ) | ( n2310  &  n1471 ) ;
 assign n2841 = ( n2574  &  n2582 ) | ( n3808  &  n2582 ) | ( n2574  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n2840 = ( n2839  &  n2841  &  n2584 ) | ( n2839  &  n2841  &  n1566 ) ;
 assign n2843 = ( n2573  &  n2590 ) | ( n3808  &  n2590 ) | ( n2573  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n2842 = ( n2839  &  n2843  &  n2592 ) | ( n2839  &  n2843  &  n1566 ) ;
 assign n2845 = ( n2566  &  n2597 ) | ( n3808  &  n2597 ) | ( n2566  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n2844 = ( n2839  &  n2845  &  n2599 ) | ( n2839  &  n2845  &  n1566 ) ;
 assign n2847 = ( n2844  &  n2842 ) | ( n3735  &  n2842 ) | ( n2844  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2848 = ( n4410  &  n4408  &  n2605 ) | ( n4410  &  n4408  &  n3807 ) ;
 assign n2846 = ( n2847  &  n2848  &  n2840 ) | ( n2847  &  n2848  &  n796 ) ;
 assign n2850 = ( n2571  &  n2610 ) | ( n3808  &  n2610 ) | ( n2571  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n2849 = ( n2839  &  n2850  &  n2612 ) | ( n2839  &  n2850  &  n1566 ) ;
 assign n2852 = ( n2570  &  n2618 ) | ( n3808  &  n2618 ) | ( n2570  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n2851 = ( n2839  &  n2852  &  n2620 ) | ( n2839  &  n2852  &  n1566 ) ;
 assign n2854 = ( n2564  &  n2625 ) | ( n3808  &  n2625 ) | ( n2564  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n2853 = ( n2839  &  n2854  &  n2627 ) | ( n2839  &  n2854  &  n1566 ) ;
 assign n2856 = ( n2853  &  n2851 ) | ( n3735  &  n2851 ) | ( n2853  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2857 = ( n4407  &  n4408  &  n2633 ) | ( n4407  &  n4408  &  n3807 ) ;
 assign n2855 = ( n2856  &  n2857  &  n2849 ) | ( n2856  &  n2857  &  n796 ) ;
 assign n2859 = ( n2577  &  n2638 ) | ( n3808  &  n2638 ) | ( n2577  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n2858 = ( n2839  &  n2859  &  n2640 ) | ( n2839  &  n2859  &  n1566 ) ;
 assign n2861 = ( n2576  &  n2646 ) | ( n3808  &  n2646 ) | ( n2576  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n2860 = ( n2839  &  n2861  &  n2648 ) | ( n2839  &  n2861  &  n1566 ) ;
 assign n2863 = ( n2568  &  n2653 ) | ( n3808  &  n2653 ) | ( n2568  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n2862 = ( n2839  &  n2863  &  n2655 ) | ( n2839  &  n2863  &  n1566 ) ;
 assign n2865 = ( n2862  &  n2860 ) | ( n3735  &  n2860 ) | ( n2862  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2866 = ( n4411  &  n4408  &  n2661 ) | ( n4411  &  n4408  &  n3807 ) ;
 assign n2864 = ( n2865  &  n2866  &  n2858 ) | ( n2865  &  n2866  &  n796 ) ;
 assign n2868 = ( n2829  &  n2666 ) | ( n3808  &  n2666 ) | ( n2829  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n2867 = ( n2839  &  n2868  &  n2668 ) | ( n2839  &  n2868  &  n1566 ) ;
 assign n2870 = ( n2832  &  n2674 ) | ( n3808  &  n2674 ) | ( n2832  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n2869 = ( n2839  &  n2870  &  n2676 ) | ( n2839  &  n2870  &  n1566 ) ;
 assign n2872 = ( n2762  &  n2681 ) | ( n3808  &  n2681 ) | ( n2762  &  n3809 ) | ( n3808  &  n3809 ) ;
 assign n2871 = ( n2839  &  n2872  &  n2683 ) | ( n2839  &  n2872  &  n1566 ) ;
 assign n2874 = ( n2871  &  n2869 ) | ( n3735  &  n2869 ) | ( n2871  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2875 = ( n4409  &  n4408  &  n2689 ) | ( n4409  &  n4408  &  n3807 ) ;
 assign n2873 = ( n2874  &  n2875  &  n2867 ) | ( n2874  &  n2875  &  n796 ) ;
 assign n2876 = ( n2306  &  n2305 ) | ( n2306  &  n1471 ) ;
 assign n2878 = ( n2582  &  n2584 ) | ( n3812  &  n2584 ) | ( n2582  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n2877 = ( n2876  &  n2878  &  n2574 ) | ( n2876  &  n2878  &  n1606 ) ;
 assign n2880 = ( n2590  &  n2592 ) | ( n3812  &  n2592 ) | ( n2590  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n2879 = ( n2876  &  n2880  &  n2573 ) | ( n2876  &  n2880  &  n1606 ) ;
 assign n2882 = ( n2597  &  n2599 ) | ( n3812  &  n2599 ) | ( n2597  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n2881 = ( n2876  &  n2882  &  n2566 ) | ( n2876  &  n2882  &  n1606 ) ;
 assign n2884 = ( n2881  &  n2879 ) | ( n3735  &  n2879 ) | ( n2881  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2885 = ( n4403  &  n4401  &  n2139 ) | ( n4403  &  n4401  &  n3811 ) ;
 assign n2883 = ( n2884  &  n2885  &  n2877 ) | ( n2884  &  n2885  &  n796 ) ;
 assign n2887 = ( n2610  &  n2612 ) | ( n3812  &  n2612 ) | ( n2610  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n2886 = ( n2876  &  n2887  &  n2571 ) | ( n2876  &  n2887  &  n1606 ) ;
 assign n2889 = ( n2618  &  n2620 ) | ( n3812  &  n2620 ) | ( n2618  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n2888 = ( n2876  &  n2889  &  n2570 ) | ( n2876  &  n2889  &  n1606 ) ;
 assign n2891 = ( n2625  &  n2627 ) | ( n3812  &  n2627 ) | ( n2625  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n2890 = ( n2876  &  n2891  &  n2564 ) | ( n2876  &  n2891  &  n1606 ) ;
 assign n2893 = ( n2890  &  n2888 ) | ( n3735  &  n2888 ) | ( n2890  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2894 = ( n4400  &  n4401  &  n2113 ) | ( n4400  &  n4401  &  n3811 ) ;
 assign n2892 = ( n2893  &  n2894  &  n2886 ) | ( n2893  &  n2894  &  n796 ) ;
 assign n2896 = ( n2638  &  n2640 ) | ( n3812  &  n2640 ) | ( n2638  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n2895 = ( n2876  &  n2896  &  n2577 ) | ( n2876  &  n2896  &  n1606 ) ;
 assign n2898 = ( n2646  &  n2648 ) | ( n3812  &  n2648 ) | ( n2646  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n2897 = ( n2876  &  n2898  &  n2576 ) | ( n2876  &  n2898  &  n1606 ) ;
 assign n2900 = ( n2653  &  n2655 ) | ( n3812  &  n2655 ) | ( n2653  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n2899 = ( n2876  &  n2900  &  n2568 ) | ( n2876  &  n2900  &  n1606 ) ;
 assign n2902 = ( n2899  &  n2897 ) | ( n3735  &  n2897 ) | ( n2899  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2903 = ( n4404  &  n4401  &  n2180 ) | ( n4404  &  n4401  &  n3811 ) ;
 assign n2901 = ( n2902  &  n2903  &  n2895 ) | ( n2902  &  n2903  &  n796 ) ;
 assign n2905 = ( n2666  &  n2668 ) | ( n3812  &  n2668 ) | ( n2666  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n2904 = ( n2876  &  n2905  &  n2829 ) | ( n2876  &  n2905  &  n1606 ) ;
 assign n2907 = ( n2674  &  n2676 ) | ( n3812  &  n2676 ) | ( n2674  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n2906 = ( n2876  &  n2907  &  n2832 ) | ( n2876  &  n2907  &  n1606 ) ;
 assign n2909 = ( n2681  &  n2683 ) | ( n3812  &  n2683 ) | ( n2681  &  n3813 ) | ( n3812  &  n3813 ) ;
 assign n2908 = ( n2876  &  n2909  &  n2762 ) | ( n2876  &  n2909  &  n1606 ) ;
 assign n2911 = ( n2908  &  n2906 ) | ( n3735  &  n2906 ) | ( n2908  &  n3738 ) | ( n3735  &  n3738 ) ;
 assign n2912 = ( n4402  &  n4401  &  n2160 ) | ( n4402  &  n4401  &  n3811 ) ;
 assign n2910 = ( n2911  &  n2912  &  n2904 ) | ( n2911  &  n2912  &  n796 ) ;
 assign n2913 = ( (~ n3499)  &  (~ n4421) ) | ( (~ n3499)  &  (~ n4422) ) ;
 assign n2916 = ( Ni10  &  (~ n3659)  &  (~ n4754) ) | ( (~ n3659)  &  (~ n3906)  &  (~ n4754) ) ;
 assign n2920 = ( n2454  &  (~ n3824) ) | ( n2458  &  (~ n3824) ) | ( (~ n3824)  &  (~ n4499) ) ;
 assign n2923 = ( n2502  &  (~ n3612) ) | ( n2504  &  (~ n3612) ) | ( (~ n3612)  &  (~ n4559) ) ;
 assign n2926 = ( (~ n1218)  &  (~ n4561) ) | ( (~ Ni11)  &  (~ n1218)  &  (~ n2311) ) ;
 assign n2931 = ( Ni11  &  (~ n1068) ) | ( Ni11  &  n2302 ) | ( (~ n1068)  &  n2300 ) | ( n2302  &  n2300 ) ;
 assign n2932 = ( n1655  &  (~ n2931) ) | ( n1653  &  n1654  &  (~ n2931) ) ;
 assign n2936 = ( (~ Ni32)  &  n3540 ) | ( (~ Ni32)  &  (~ n3923) ) | ( (~ n3540)  &  (~ n3923) ) ;
 assign n2937 = ( Ni36 ) | ( (~ Ni38) ) ;
 assign n2939 = ( Pi19  &  Pi17 ) ;
 assign n2947 = ( (~ Ni45) ) | ( n2946 ) ;
 assign n2946 = ( Ni45  &  Ni46 ) ;
 assign n2950 = ( (~ Ni40) ) | ( Ni30  &  n837 ) ;
 assign n2952 = ( (~ n1655)  &  (~ n1653) ) | ( (~ n1653)  &  n3928 ) | ( (~ n1655)  &  (~ n3930) ) | ( n3928  &  (~ n3930) ) ;
 assign n2953 = ( (~ Ni41) ) | ( Ni30  &  n837 ) ;
 assign n2954 = ( (~ n1655)  &  (~ n1653) ) | ( (~ n1653)  &  n3934 ) | ( (~ n1655)  &  (~ n3936) ) | ( n3934  &  (~ n3936) ) ;
 assign n2955 = ( Ni45  &  (~ n2946) ) | ( (~ n2946)  &  (~ n3480) ) ;
 assign n2959 = ( (~ Ni47) ) | ( (~ Ni48) ) ;
 assign n2958 = ( Ni45  &  (~ n2946) ) | ( (~ n2946)  &  n2959 ) ;
 assign n2961 = ( Ni38 ) | ( (~ Ni39) ) ;
 assign n2962 = ( Ni39 ) | ( Ni38 ) ;
 assign n2960 = ( n2955  &  n2958 ) | ( n2961  &  n2958 ) | ( n2955  &  n2962 ) | ( n2961  &  n2962 ) ;
 assign n2965 = ( (~ Ni37) ) | ( n2960 ) ;
 assign n2964 = ( n2958  &  n2971 ) | ( n2958  &  (~ Ni42) ) ;
 assign n2963 = ( (~ n200)  &  n2965 ) | ( n2965  &  n2964 ) ;
 assign n2967 = ( n3122  &  Ni42 ) | ( n3122  &  n2955 ) ;
 assign n2966 = ( (~ n200)  &  n2965 ) | ( n2965  &  n2967 ) ;
 assign n2968 = ( (~ n171)  &  n1063 ) | ( (~ n171)  &  n2958 ) ;
 assign n2971 = ( n2958  &  n2955 ) | ( n2958  &  n3120 ) ;
 assign n2970 = ( n2964  &  Ni41 ) | ( n2964  &  n2971 ) ;
 assign n2972 = ( n2971  &  n2955 ) | ( n2971  &  n320 ) ;
 assign n2973 = ( n2964  &  Ni41 ) | ( n2964  &  n2972 ) ;
 assign n2975 = ( n2967 ) | ( n3724 ) ;
 assign n2976 = ( n2978 ) | ( n202  &  n3858 ) ;
 assign n2974 = ( n2975  &  n2965  &  n2976 ) ;
 assign n2979 = ( Ni37 ) | ( n3866 ) ;
 assign n2978 = ( n2970  &  n2973 ) | ( n2970  &  (~ Ni40) ) ;
 assign n2977 = ( (~ n150)  &  n2979 ) | ( n2979  &  n2978 ) ;
 assign n2980 = ( (~ n2199)  &  n2974 ) | ( n2974  &  n2977 ) ;
 assign n2981 = ( (~ n2078)  &  n2096  &  (~ n2955) ) | ( (~ n2078)  &  (~ n2955)  &  (~ n2958) ) ;
 assign n2986 = ( Ni41 ) | ( (~ Ni42) ) ;
 assign n2985 = ( n2971  &  (~ n2981) ) | ( (~ n2981)  &  n2986 ) ;
 assign n2989 = ( n2967 ) | ( n3725 ) ;
 assign n2990 = ( n2992 ) | ( n240  &  n3858 ) ;
 assign n2988 = ( n2989  &  n2965  &  n2990 ) ;
 assign n2992 = ( n2973  &  n3020 ) | ( n3020  &  (~ Ni40) ) ;
 assign n2991 = ( (~ n150)  &  n2979 ) | ( n2979  &  n2992 ) ;
 assign n2993 = ( (~ n2199)  &  n2988 ) | ( n2988  &  n2991 ) ;
 assign n2995 = ( Pi20 ) | ( Pi19 ) ;
 assign n2996 = ( (~ Pi20) ) | ( Pi19 ) ;
 assign n2994 = ( n2980  &  n2993 ) | ( n2995  &  n2993 ) | ( n2980  &  n2996 ) | ( n2995  &  n2996 ) ;
 assign n2997 = ( n2965  &  n2973  &  n2979 ) | ( n2965  &  n2979  &  (~ Ni38) ) ;
 assign n3001 = ( Pi21  &  Pi19 ) ;
 assign n2999 = ( Pi22  &  (~ n3352) ) ;
 assign n2998 = ( n192  &  n3001 ) | ( (~ n2997)  &  n3001  &  n2999 ) ;
 assign n3003 = ( n3005 ) | ( n202  &  n3858 ) ;
 assign n3002 = ( n2975  &  n2965  &  n3003 ) ;
 assign n3005 = ( n2972  &  n3053 ) | ( n3053  &  (~ Ni40) ) ;
 assign n3004 = ( (~ n150)  &  n2979 ) | ( n2979  &  n3005 ) ;
 assign n3006 = ( (~ n2199)  &  n3002 ) | ( n3002  &  n3004 ) ;
 assign n3007 = ( (~ Ni41)  &  n2985 ) | ( n2972  &  n2985 ) ;
 assign n3009 = ( n3011 ) | ( n240  &  n3858 ) ;
 assign n3008 = ( n2989  &  n2965  &  n3009 ) ;
 assign n3011 = ( n2972  &  n3007 ) | ( n3007  &  (~ Ni40) ) ;
 assign n3010 = ( (~ n150)  &  n2979 ) | ( n2979  &  n3011 ) ;
 assign n3012 = ( (~ n2199)  &  n3008 ) | ( n3008  &  n3010 ) ;
 assign n3013 = ( n3006  &  n3012 ) | ( n2995  &  n3012 ) | ( n3006  &  n2996 ) | ( n2995  &  n2996 ) ;
 assign n3014 = ( n2965  &  n2972  &  n2979 ) | ( n2965  &  n2979  &  (~ Ni38) ) ;
 assign n3015 = ( n192  &  n3001 ) | ( n3001  &  n2999  &  (~ n3014) ) ;
 assign n3018 = ( n3020 ) | ( n240  &  n3858 ) ;
 assign n3017 = ( n2989  &  n2965  &  n3018 ) ;
 assign n3021 = ( n63 ) | ( n3866 ) ;
 assign n3020 = ( n2964  &  n2985 ) ;
 assign n3019 = ( n3021  &  n3017  &  n663 ) | ( n3021  &  n3017  &  n3020 ) ;
 assign n3023 = ( n3020  &  Ni40 ) | ( n3020  &  n2973 ) ;
 assign n3022 = ( (~ n150)  &  n2979 ) | ( n2979  &  n3023 ) ;
 assign n3025 = ( n3023 ) | ( n240  &  n3858 ) ;
 assign n3024 = ( n2989  &  n2965  &  n3025 ) ;
 assign n3026 = ( (~ n2087)  &  n3024 ) | ( n3022  &  n3024 ) ;
 assign n3028 = ( n3007 ) | ( n240  &  n3858 ) ;
 assign n3027 = ( n2989  &  n2965  &  n3028 ) ;
 assign n3029 = ( n3021  &  n3027  &  n663 ) | ( n3021  &  n3027  &  n3007 ) ;
 assign n3031 = ( n3007  &  Ni40 ) | ( n3007  &  n2972 ) ;
 assign n3030 = ( (~ n150)  &  n2979 ) | ( n2979  &  n3031 ) ;
 assign n3033 = ( n3031 ) | ( n240  &  n3858 ) ;
 assign n3032 = ( n2989  &  n2965  &  n3033 ) ;
 assign n3034 = ( (~ n2087)  &  n3032 ) | ( n3030  &  n3032 ) ;
 assign n3035 = ( (~ n173)  &  (~ n3869) ) ;
 assign n3039 = ( n3029  &  n3034 ) | ( n3582  &  n3034 ) | ( n3029  &  n3576 ) | ( n3582  &  n3576 ) ;
 assign n3040 = ( n3019  &  n3026 ) | ( n1884  &  n3026 ) | ( n3019  &  n3778 ) | ( n1884  &  n3778 ) ;
 assign n3038 = ( n3035  &  (~ n3065) ) | ( n3035  &  n3039  &  n3040 ) ;
 assign n3043 = ( n2970 ) | ( n202  &  n3858 ) ;
 assign n3042 = ( n2975  &  n2965  &  n3043 ) ;
 assign n3044 = ( n3021  &  n3042  &  n663 ) | ( n3021  &  n3042  &  n2970 ) ;
 assign n3046 = ( n2970  &  Ni40 ) | ( n2970  &  n2973 ) ;
 assign n3045 = ( (~ n150)  &  n2979 ) | ( n2979  &  n3046 ) ;
 assign n3048 = ( n3046 ) | ( n202  &  n3858 ) ;
 assign n3047 = ( n2975  &  n2965  &  n3048 ) ;
 assign n3049 = ( (~ n2087)  &  n3047 ) | ( n3045  &  n3047 ) ;
 assign n3051 = ( n3053 ) | ( n202  &  n3858 ) ;
 assign n3050 = ( n2975  &  n2965  &  n3051 ) ;
 assign n3053 = ( (~ Ni41)  &  n2971 ) | ( n2971  &  n2972 ) ;
 assign n3052 = ( n3021  &  n3050  &  n663 ) | ( n3021  &  n3050  &  n3053 ) ;
 assign n3055 = ( n3053  &  Ni40 ) | ( n3053  &  n2972 ) ;
 assign n3054 = ( (~ n150)  &  n2979 ) | ( n2979  &  n3055 ) ;
 assign n3057 = ( n3055 ) | ( n202  &  n3858 ) ;
 assign n3056 = ( n2975  &  n2965  &  n3057 ) ;
 assign n3058 = ( (~ n2087)  &  n3056 ) | ( n3054  &  n3056 ) ;
 assign n3060 = ( Pi22  &  (~ n4767) ) | ( (~ Pi21)  &  (~ n4767) ) | ( n2968  &  (~ n4767) ) ;
 assign n3059 = ( (~ n173)  &  n3060 ) ;
 assign n3062 = ( n3052  &  n3058 ) | ( n3582  &  n3058 ) | ( n3052  &  n3576 ) | ( n3582  &  n3576 ) ;
 assign n3063 = ( n3044  &  n3049 ) | ( n1884  &  n3049 ) | ( n3044  &  n3778 ) | ( n1884  &  n3778 ) ;
 assign n3061 = ( n3059  &  (~ n3065) ) | ( n3059  &  n3062  &  n3063 ) ;
 assign n3065 = ( (~ n1866)  &  (~ n3352) ) ;
 assign n3064 = ( n2998  &  (~ n3870) ) | ( (~ n2994)  &  n3065  &  (~ n3870) ) ;
 assign n3068 = ( n3015  &  (~ n3871) ) | ( (~ n3013)  &  n3065  &  (~ n3871) ) ;
 assign n3072 = ( n2978  &  n2977 ) | ( n63  &  n2977 ) | ( n2978  &  n2087 ) | ( n63  &  n2087 ) ;
 assign n3071 = ( n3072  &  n2974 ) ;
 assign n3074 = ( n2992  &  n2991 ) | ( n63  &  n2991 ) | ( n2992  &  n2087 ) | ( n63  &  n2087 ) ;
 assign n3073 = ( n3074  &  n2988 ) ;
 assign n3075 = ( n3071  &  n3073 ) | ( n2995  &  n3073 ) | ( n3071  &  n2996 ) | ( n2995  &  n2996 ) ;
 assign n3077 = ( n2965  &  n2973 ) | ( n2965  &  n53 ) ;
 assign n3076 = ( n3077  &  Ni36 ) | ( n3077  &  n2997 ) ;
 assign n3078 = ( n3001  &  n2999  &  (~ n3076) ) ;
 assign n3081 = ( n3005  &  n3004 ) | ( n63  &  n3004 ) | ( n3005  &  n2087 ) | ( n63  &  n2087 ) ;
 assign n3080 = ( n3081  &  n3002 ) ;
 assign n3083 = ( n3011  &  n3010 ) | ( n63  &  n3010 ) | ( n3011  &  n2087 ) | ( n63  &  n2087 ) ;
 assign n3082 = ( n3083  &  n3008 ) ;
 assign n3084 = ( n3080  &  n3082 ) | ( n2995  &  n3082 ) | ( n3080  &  n2996 ) | ( n2995  &  n2996 ) ;
 assign n3086 = ( n2965  &  n2972 ) | ( n2965  &  n53 ) ;
 assign n3085 = ( n3086  &  Ni36 ) | ( n3086  &  n3014 ) ;
 assign n3087 = ( n192  &  n3001 ) | ( n3001  &  n2999  &  (~ n3085) ) ;
 assign n3089 = ( n3017  &  n3020 ) | ( n3017  &  n63 ) ;
 assign n3091 = ( n3023  &  n3022 ) | ( n63  &  n3022 ) | ( n3023  &  n2199 ) | ( n63  &  n2199 ) ;
 assign n3090 = ( n3091  &  n3024 ) ;
 assign n3092 = ( n3027  &  n3007 ) | ( n3027  &  n63 ) ;
 assign n3094 = ( n3031  &  n3030 ) | ( n63  &  n3030 ) | ( n3031  &  n2199 ) | ( n63  &  n2199 ) ;
 assign n3093 = ( n3094  &  n3032 ) ;
 assign n3096 = ( n3092  &  n3093 ) | ( n3582  &  n3093 ) | ( n3092  &  n3576 ) | ( n3582  &  n3576 ) ;
 assign n3097 = ( n3089  &  n3090 ) | ( n1884  &  n3090 ) | ( n3089  &  n3778 ) | ( n1884  &  n3778 ) ;
 assign n3095 = ( n3035  &  (~ n3065) ) | ( n3035  &  n3096  &  n3097 ) ;
 assign n3098 = ( n3042  &  n2970 ) | ( n3042  &  n63 ) ;
 assign n3100 = ( n3046  &  n3045 ) | ( n63  &  n3045 ) | ( n3046  &  n2199 ) | ( n63  &  n2199 ) ;
 assign n3099 = ( n3100  &  n3047 ) ;
 assign n3101 = ( n3050  &  n3053 ) | ( n3050  &  n63 ) ;
 assign n3103 = ( n3055  &  n3054 ) | ( n63  &  n3054 ) | ( n3055  &  n2199 ) | ( n63  &  n2199 ) ;
 assign n3102 = ( n3103  &  n3056 ) ;
 assign n3105 = ( n3101  &  n3102 ) | ( n3582  &  n3102 ) | ( n3101  &  n3576 ) | ( n3582  &  n3576 ) ;
 assign n3106 = ( n3098  &  n3099 ) | ( n1884  &  n3099 ) | ( n3098  &  n3778 ) | ( n1884  &  n3778 ) ;
 assign n3104 = ( n3059  &  (~ n3065) ) | ( n3059  &  n3105  &  n3106 ) ;
 assign n3107 = ( n3078  &  (~ n3870) ) | ( n3065  &  (~ n3075)  &  (~ n3870) ) ;
 assign n3109 = ( n3087  &  (~ n3871) ) | ( n3065  &  (~ n3084)  &  (~ n3871) ) ;
 assign n3113 = ( Ni11 ) | ( n931 ) ;
 assign n3111 = ( (~ n188)  &  n3113 ) | ( (~ n1866)  &  n3113  &  (~ n3261) ) ;
 assign n3114 = ( n3107  &  (~ n3831) ) | ( n3109  &  (~ n3831) ) | ( (~ n3831)  &  (~ n3949) ) ;
 assign n3116 = ( (~ n1993)  &  n3064 ) | ( (~ n1993)  &  n3068 ) | ( (~ n1993)  &  (~ n3950) ) ;
 assign n3120 = ( (~ Ni44) ) | ( Ni43 ) ;
 assign n3119 = ( (~ n2078)  &  (~ n2955)  &  (~ n2958) ) | ( (~ n2078)  &  (~ n2955)  &  n3120 ) ;
 assign n3122 = ( n2958  &  n2096 ) | ( n2958  &  n2955 ) ;
 assign n3121 = ( n2986  &  (~ n3119) ) | ( (~ n3119)  &  n3122 ) ;
 assign n3125 = ( n2958  &  n2955 ) | ( n2958  &  n3593 ) ;
 assign n3124 = ( n3122  &  n3125 ) | ( n3125  &  (~ Ni42) ) ;
 assign n3127 = ( n3143  &  Ni40 ) | ( n3143  &  n3185 ) ;
 assign n3126 = ( n3127 ) | ( n202 ) ;
 assign n3129 = ( Ni37 ) | ( n3864 ) ;
 assign n3130 = ( n3127 ) | ( (~ n150)  &  n3858 ) ;
 assign n3128 = ( n3129  &  n2965  &  n3130 ) ;
 assign n3132 = ( n3127 ) | ( n63 ) ;
 assign n3131 = ( n3128  &  n3132  &  Ni35 ) | ( n3128  &  n3132  &  n3126 ) ;
 assign n3134 = ( (~ n171)  &  n3279 ) ;
 assign n3133 = ( (~ Ni33)  &  n3134 ) | ( n3131  &  n3134 ) ;
 assign n3136 = ( n3143  &  Ni40 ) | ( n3143  &  n3191 ) ;
 assign n3135 = ( n3136 ) | ( n240 ) ;
 assign n3138 = ( n3136 ) | ( (~ n150)  &  n3858 ) ;
 assign n3137 = ( n3129  &  n2965  &  n3138 ) ;
 assign n3140 = ( n3136 ) | ( n63 ) ;
 assign n3139 = ( n3137  &  n3140  &  Ni35 ) | ( n3137  &  n3140  &  n3135 ) ;
 assign n3141 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3139 ) ;
 assign n3143 = ( n3124  &  n3697 ) ;
 assign n3142 = ( n2965  &  n3129  &  n3143 ) | ( n2965  &  n3129  &  (~ Ni38) ) ;
 assign n3144 = ( n3142  &  n3143 ) | ( n3142  &  n53 ) ;
 assign n3145 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3144 ) ;
 assign n3147 = ( n3133  &  n3141 ) | ( n891  &  n3141 ) | ( n3133  &  n310 ) | ( n891  &  n310 ) ;
 assign n3146 = ( n188  &  n3147  &  n3145 ) | ( n188  &  n3147  &  n1250 ) ;
 assign n3149 = ( n3124  &  Ni40 ) | ( n3124  &  n3213 ) ;
 assign n3148 = ( n3149 ) | ( n202 ) ;
 assign n3151 = ( n3149 ) | ( (~ n150)  &  n3858 ) ;
 assign n3150 = ( n3129  &  n2965  &  n3151 ) ;
 assign n3153 = ( n3149 ) | ( n63 ) ;
 assign n3152 = ( n3150  &  n3153  &  Ni35 ) | ( n3150  &  n3153  &  n3148 ) ;
 assign n3154 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3152 ) ;
 assign n3156 = ( n3124  &  Ni40 ) | ( n3124  &  n3218 ) ;
 assign n3155 = ( n3156 ) | ( n240 ) ;
 assign n3158 = ( n3156 ) | ( (~ n150)  &  n3858 ) ;
 assign n3157 = ( n3129  &  n2965  &  n3158 ) ;
 assign n3160 = ( n3156 ) | ( n63 ) ;
 assign n3159 = ( n3157  &  n3160  &  Ni35 ) | ( n3157  &  n3160  &  n3155 ) ;
 assign n3161 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3159 ) ;
 assign n3162 = ( n2965  &  n3124  &  n3129 ) | ( n2965  &  n3129  &  (~ Ni38) ) ;
 assign n3163 = ( n3162  &  n3124 ) | ( n3162  &  n53 ) ;
 assign n3164 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3163 ) ;
 assign n3166 = ( n3154  &  n3161 ) | ( n891  &  n3161 ) | ( n3154  &  n310 ) | ( n891  &  n310 ) ;
 assign n3165 = ( n188  &  n3166  &  n3164 ) | ( n188  &  n3166  &  n1250 ) ;
 assign n3167 = ( n3128  &  Ni35 ) | ( n3128  &  n3126 ) ;
 assign n3168 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3167 ) ;
 assign n3169 = ( n3137  &  Ni35 ) | ( n3137  &  n3135 ) ;
 assign n3170 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3169 ) ;
 assign n3171 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3142 ) ;
 assign n3173 = ( n3168  &  n3170 ) | ( n891  &  n3170 ) | ( n3168  &  n310 ) | ( n891  &  n310 ) ;
 assign n3172 = ( n188  &  n3173  &  n3171 ) | ( n188  &  n3173  &  n1250 ) ;
 assign n3174 = ( n3150  &  Ni35 ) | ( n3150  &  n3148 ) ;
 assign n3175 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3174 ) ;
 assign n3176 = ( n3157  &  Ni35 ) | ( n3157  &  n3155 ) ;
 assign n3177 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3176 ) ;
 assign n3178 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3162 ) ;
 assign n3180 = ( n3175  &  n3177 ) | ( n891  &  n3177 ) | ( n3175  &  n310 ) | ( n891  &  n310 ) ;
 assign n3179 = ( n188  &  n3180  &  n3178 ) | ( n188  &  n3180  &  n1250 ) ;
 assign n3182 = ( n2964 ) | ( n3724 ) ;
 assign n3183 = ( n3185 ) | ( n202  &  n3858 ) ;
 assign n3181 = ( n3182  &  n2965  &  n3183 ) ;
 assign n3185 = ( n3697  &  n3121 ) ;
 assign n3184 = ( n3181  &  n3185 ) | ( n3181  &  n63 ) ;
 assign n3186 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3184 ) ;
 assign n3188 = ( n2964 ) | ( n3725 ) ;
 assign n3189 = ( n3191 ) | ( n240  &  n3858 ) ;
 assign n3187 = ( n3188  &  n2965  &  n3189 ) ;
 assign n3191 = ( n3122  &  n3697 ) ;
 assign n3190 = ( n3187  &  n3191 ) | ( n3187  &  n63 ) ;
 assign n3192 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3190 ) ;
 assign n3194 = ( n3196 ) | ( (~ n150)  &  n3858 ) ;
 assign n3193 = ( n3129  &  n2965  &  n3194 ) ;
 assign n3196 = ( n3143  &  n3185 ) | ( n3143  &  (~ Ni40) ) ;
 assign n3195 = ( n3196 ) | ( n202 ) ;
 assign n3198 = ( n3196 ) | ( n63 ) ;
 assign n3197 = ( (~ Ni35)  &  n3193  &  n3198 ) | ( n3193  &  n3195  &  n3198 ) ;
 assign n3199 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3197 ) ;
 assign n3201 = ( n3203 ) | ( (~ n150)  &  n3858 ) ;
 assign n3200 = ( n3129  &  n2965  &  n3201 ) ;
 assign n3203 = ( n3143  &  n3191 ) | ( n3143  &  (~ Ni40) ) ;
 assign n3202 = ( n3203 ) | ( n240 ) ;
 assign n3205 = ( n3203 ) | ( n63 ) ;
 assign n3204 = ( (~ Ni35)  &  n3200  &  n3205 ) | ( n3200  &  n3202  &  n3205 ) ;
 assign n3206 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3204 ) ;
 assign n3208 = ( n188  &  n3199 ) | ( n188  &  n3776 ) ;
 assign n3209 = ( n3186  &  n3192 ) | ( n891  &  n3192 ) | ( n3186  &  n310 ) | ( n891  &  n310 ) ;
 assign n3207 = ( n3208  &  n3209  &  n3206 ) | ( n3208  &  n3209  &  n1692 ) ;
 assign n3211 = ( n3213 ) | ( n202  &  n3858 ) ;
 assign n3210 = ( n3182  &  n2965  &  n3211 ) ;
 assign n3213 = ( n3124  &  n3121 ) ;
 assign n3212 = ( n3210  &  n3213 ) | ( n3210  &  n63 ) ;
 assign n3214 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3212 ) ;
 assign n3216 = ( n3218 ) | ( n240  &  n3858 ) ;
 assign n3215 = ( n3188  &  n2965  &  n3216 ) ;
 assign n3218 = ( n3124  &  Ni41 ) | ( n3124  &  n3122 ) ;
 assign n3217 = ( n3215  &  n3218 ) | ( n3215  &  n63 ) ;
 assign n3219 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3217 ) ;
 assign n3221 = ( n3223 ) | ( (~ n150)  &  n3858 ) ;
 assign n3220 = ( n3129  &  n2965  &  n3221 ) ;
 assign n3223 = ( n3124  &  n3213 ) | ( n3124  &  (~ Ni40) ) ;
 assign n3222 = ( n3223 ) | ( n202 ) ;
 assign n3225 = ( n3223 ) | ( n63 ) ;
 assign n3224 = ( (~ Ni35)  &  n3220  &  n3225 ) | ( n3220  &  n3222  &  n3225 ) ;
 assign n3226 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3224 ) ;
 assign n3228 = ( n3230 ) | ( (~ n150)  &  n3858 ) ;
 assign n3227 = ( n3129  &  n2965  &  n3228 ) ;
 assign n3230 = ( n3124  &  n3218 ) | ( n3124  &  (~ Ni40) ) ;
 assign n3229 = ( n3230 ) | ( n240 ) ;
 assign n3232 = ( n3230 ) | ( n63 ) ;
 assign n3231 = ( (~ Ni35)  &  n3227  &  n3232 ) | ( n3227  &  n3229  &  n3232 ) ;
 assign n3233 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3231 ) ;
 assign n3235 = ( n188  &  n3226 ) | ( n188  &  n3776 ) ;
 assign n3236 = ( n3214  &  n3219 ) | ( n891  &  n3219 ) | ( n3214  &  n310 ) | ( n891  &  n310 ) ;
 assign n3234 = ( n3235  &  n3236  &  n3233 ) | ( n3235  &  n3236  &  n1692 ) ;
 assign n3238 = ( n63 ) | ( n3864 ) ;
 assign n3237 = ( n3238  &  n3181  &  n663 ) | ( n3238  &  n3181  &  n3185 ) ;
 assign n3239 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3237 ) ;
 assign n3240 = ( n3238  &  n3187  &  n663 ) | ( n3238  &  n3187  &  n3191 ) ;
 assign n3241 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3240 ) ;
 assign n3242 = ( (~ Ni35)  &  n3193 ) | ( n3193  &  n3195 ) ;
 assign n3243 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3242 ) ;
 assign n3244 = ( (~ Ni35)  &  n3200 ) | ( n3200  &  n3202 ) ;
 assign n3245 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3244 ) ;
 assign n3247 = ( n188  &  n3243 ) | ( n188  &  n3776 ) ;
 assign n3248 = ( n3239  &  n3241 ) | ( n891  &  n3241 ) | ( n3239  &  n310 ) | ( n891  &  n310 ) ;
 assign n3246 = ( n3247  &  n3248  &  n3245 ) | ( n3247  &  n3248  &  n1692 ) ;
 assign n3249 = ( n3238  &  n3210  &  n663 ) | ( n3238  &  n3210  &  n3213 ) ;
 assign n3250 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3249 ) ;
 assign n3251 = ( n3238  &  n3215  &  n663 ) | ( n3238  &  n3215  &  n3218 ) ;
 assign n3252 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3251 ) ;
 assign n3253 = ( (~ Ni35)  &  n3220 ) | ( n3220  &  n3222 ) ;
 assign n3254 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3253 ) ;
 assign n3255 = ( (~ Ni35)  &  n3227 ) | ( n3227  &  n3229 ) ;
 assign n3256 = ( (~ Ni33)  &  n3134 ) | ( n3134  &  n3255 ) ;
 assign n3258 = ( n188  &  n3254 ) | ( n188  &  n3776 ) ;
 assign n3259 = ( n3250  &  n3252 ) | ( n891  &  n3252 ) | ( n3250  &  n310 ) | ( n891  &  n310 ) ;
 assign n3257 = ( n3258  &  n3259  &  n3256 ) | ( n3258  &  n3259  &  n1692 ) ;
 assign n3261 = ( (~ n193)  &  n3279 ) ;
 assign n3260 = ( n188  &  n3261 ) | ( n188  &  n1471 ) ;
 assign n3262 = ( (~ n1965)  &  n3171 ) | ( n3171  &  n3178 ) | ( (~ n1965)  &  (~ n3618) ) | ( n3178  &  (~ n3618) ) ;
 assign n3265 = ( (~ n1884)  &  (~ n3260) ) | ( (~ n1884)  &  (~ n4581) ) ;
 assign n3268 = ( (~ n3260)  &  (~ n3582) ) | ( (~ n3582)  &  (~ n4583) ) ;
 assign n3270 = ( (~ n1965)  &  n3145 ) | ( n3145  &  n3164 ) | ( (~ n1965)  &  (~ n3618) ) | ( n3164  &  (~ n3618) ) ;
 assign n3271 = ( (~ n3260)  &  (~ n3579) ) | ( (~ n3579)  &  (~ n4568) ) ;
 assign n3273 = ( (~ n1884)  &  (~ n3260) ) | ( (~ n1884)  &  (~ n4569) ) ;
 assign n3275 = ( (~ n3260)  &  (~ n3582) ) | ( (~ n3582)  &  (~ n4571) ) ;
 assign n3279 = ( Ni33 ) | ( n2963 ) | ( n1063 ) ;
 assign n3278 = ( (~ Ni34) ) | ( n2966 ) ;
 assign n3277 = ( (~ n171)  &  (~ Ni33)  &  n3279 ) | ( (~ n171)  &  n3279  &  n3278 ) ;
 assign n3281 = ( Ni34 ) | ( (~ Ni33) ) ;
 assign n3280 = ( n3277  &  n3131 ) | ( n3277  &  n3281 ) ;
 assign n3282 = ( n3277  &  n3139 ) | ( n3277  &  n3281 ) ;
 assign n3283 = ( n3277  &  n3144 ) | ( n3277  &  n3281 ) ;
 assign n3285 = ( n3280  &  n3282 ) | ( n891  &  n3282 ) | ( n3280  &  n310 ) | ( n891  &  n310 ) ;
 assign n3284 = ( n188  &  n3285  &  n3283 ) | ( n188  &  n3285  &  n1250 ) ;
 assign n3286 = ( n3277  &  n3152 ) | ( n3277  &  n3281 ) ;
 assign n3287 = ( n3277  &  n3159 ) | ( n3277  &  n3281 ) ;
 assign n3288 = ( n3277  &  n3163 ) | ( n3277  &  n3281 ) ;
 assign n3290 = ( n3286  &  n3287 ) | ( n891  &  n3287 ) | ( n3286  &  n310 ) | ( n891  &  n310 ) ;
 assign n3289 = ( n188  &  n3290  &  n3288 ) | ( n188  &  n3290  &  n1250 ) ;
 assign n3291 = ( n3277  &  n3167 ) | ( n3277  &  n3281 ) ;
 assign n3292 = ( n3277  &  n3169 ) | ( n3277  &  n3281 ) ;
 assign n3293 = ( n3277  &  n3142 ) | ( n3277  &  n3281 ) ;
 assign n3295 = ( n3291  &  n3292 ) | ( n891  &  n3292 ) | ( n3291  &  n310 ) | ( n891  &  n310 ) ;
 assign n3294 = ( n188  &  n3295  &  n3293 ) | ( n188  &  n3295  &  n1250 ) ;
 assign n3296 = ( n3277  &  n3174 ) | ( n3277  &  n3281 ) ;
 assign n3297 = ( n3277  &  n3176 ) | ( n3277  &  n3281 ) ;
 assign n3298 = ( n3277  &  n3162 ) | ( n3277  &  n3281 ) ;
 assign n3300 = ( n3296  &  n3297 ) | ( n891  &  n3297 ) | ( n3296  &  n310 ) | ( n891  &  n310 ) ;
 assign n3299 = ( n188  &  n3300  &  n3298 ) | ( n188  &  n3300  &  n1250 ) ;
 assign n3301 = ( n3277  &  n3184 ) | ( n3277  &  n3281 ) ;
 assign n3302 = ( n3277  &  n3190 ) | ( n3277  &  n3281 ) ;
 assign n3303 = ( n3277  &  n3197 ) | ( n3277  &  n3281 ) ;
 assign n3304 = ( n3277  &  n3204 ) | ( n3277  &  n3281 ) ;
 assign n3306 = ( n188  &  n3303 ) | ( n188  &  n3776 ) ;
 assign n3307 = ( n3301  &  n3302 ) | ( n891  &  n3302 ) | ( n3301  &  n310 ) | ( n891  &  n310 ) ;
 assign n3305 = ( n3306  &  n3307  &  n3304 ) | ( n3306  &  n3307  &  n1692 ) ;
 assign n3308 = ( n3277  &  n3212 ) | ( n3277  &  n3281 ) ;
 assign n3309 = ( n3277  &  n3217 ) | ( n3277  &  n3281 ) ;
 assign n3310 = ( n3277  &  n3224 ) | ( n3277  &  n3281 ) ;
 assign n3311 = ( n3277  &  n3231 ) | ( n3277  &  n3281 ) ;
 assign n3313 = ( n188  &  n3310 ) | ( n188  &  n3776 ) ;
 assign n3314 = ( n3308  &  n3309 ) | ( n891  &  n3309 ) | ( n3308  &  n310 ) | ( n891  &  n310 ) ;
 assign n3312 = ( n3313  &  n3314  &  n3311 ) | ( n3313  &  n3314  &  n1692 ) ;
 assign n3315 = ( n3277  &  n3237 ) | ( n3277  &  n3281 ) ;
 assign n3316 = ( n3277  &  n3240 ) | ( n3277  &  n3281 ) ;
 assign n3317 = ( n3277  &  n3242 ) | ( n3277  &  n3281 ) ;
 assign n3318 = ( n3277  &  n3244 ) | ( n3277  &  n3281 ) ;
 assign n3320 = ( n188  &  n3317 ) | ( n188  &  n3776 ) ;
 assign n3321 = ( n3315  &  n3316 ) | ( n891  &  n3316 ) | ( n3315  &  n310 ) | ( n891  &  n310 ) ;
 assign n3319 = ( n3320  &  n3321  &  n3318 ) | ( n3320  &  n3321  &  n1692 ) ;
 assign n3322 = ( n3277  &  n3249 ) | ( n3277  &  n3281 ) ;
 assign n3323 = ( n3277  &  n3251 ) | ( n3277  &  n3281 ) ;
 assign n3324 = ( n3277  &  n3253 ) | ( n3277  &  n3281 ) ;
 assign n3325 = ( n3277  &  n3255 ) | ( n3277  &  n3281 ) ;
 assign n3327 = ( n188  &  n3324 ) | ( n188  &  n3776 ) ;
 assign n3328 = ( n3322  &  n3323 ) | ( n891  &  n3323 ) | ( n3322  &  n310 ) | ( n891  &  n310 ) ;
 assign n3326 = ( n3327  &  n3328  &  n3325 ) | ( n3327  &  n3328  &  n1692 ) ;
 assign n3329 = ( (~ n1965)  &  n3293 ) | ( n3293  &  n3298 ) | ( (~ n1965)  &  (~ n3618) ) | ( n3298  &  (~ n3618) ) ;
 assign n3330 = ( (~ n1884)  &  (~ n3260) ) | ( (~ n1884)  &  (~ n4605) ) ;
 assign n3332 = ( (~ n3260)  &  (~ n3582) ) | ( (~ n3582)  &  (~ n4607) ) ;
 assign n3334 = ( (~ n1965)  &  n3283 ) | ( n3283  &  n3288 ) | ( (~ n1965)  &  (~ n3618) ) | ( n3288  &  (~ n3618) ) ;
 assign n3335 = ( (~ n3260)  &  (~ n3579) ) | ( (~ n3579)  &  (~ n4593) ) ;
 assign n3337 = ( (~ n1884)  &  (~ n3260) ) | ( (~ n1884)  &  (~ n4594) ) ;
 assign n3339 = ( (~ n3260)  &  (~ n3582) ) | ( (~ n3582)  &  (~ n4596) ) ;
 assign n3342 = ( Ni34 ) | ( n2963 ) | ( n3865 ) ;
 assign n3341 = ( (~ n171)  &  (~ Ni33)  &  n3342 ) | ( (~ n171)  &  n3278  &  n3342 ) ;
 assign n3344 = ( n3071 ) | ( n3352 ) ;
 assign n3343 = ( n3344  &  n3341  &  n3131 ) | ( n3344  &  n3341  &  n3281 ) ;
 assign n3346 = ( n3073 ) | ( n3352 ) ;
 assign n3345 = ( n3346  &  n3341  &  n3139 ) | ( n3346  &  n3341  &  n3281 ) ;
 assign n3348 = ( n3076  &  n3144 ) | ( n3352  &  n3144 ) | ( n3076  &  n3281 ) | ( n3352  &  n3281 ) ;
 assign n3347 = ( n3348  &  n3341 ) ;
 assign n3350 = ( n3343  &  n3345 ) | ( n891  &  n3345 ) | ( n3343  &  n310 ) | ( n891  &  n310 ) ;
 assign n3349 = ( n188  &  n3350  &  n3347 ) | ( n188  &  n3350  &  n1250 ) ;
 assign n3353 = ( n3152 ) | ( n3281 ) ;
 assign n3352 = ( n1063 ) | ( n3840 ) ;
 assign n3351 = ( n3353  &  n3341  &  n3080 ) | ( n3353  &  n3341  &  n3352 ) ;
 assign n3355 = ( n3159 ) | ( n3281 ) ;
 assign n3354 = ( n3355  &  n3341  &  n3082 ) | ( n3355  &  n3341  &  n3352 ) ;
 assign n3357 = ( n3085  &  n3163 ) | ( n3352  &  n3163 ) | ( n3085  &  n3281 ) | ( n3352  &  n3281 ) ;
 assign n3356 = ( n3357  &  n3341 ) ;
 assign n3359 = ( n3351  &  n3354 ) | ( n891  &  n3354 ) | ( n3351  &  n310 ) | ( n891  &  n310 ) ;
 assign n3358 = ( n188  &  n3359  &  n3356 ) | ( n188  &  n3359  &  n1250 ) ;
 assign n3361 = ( n2980 ) | ( n3352 ) ;
 assign n3360 = ( n3361  &  n3341  &  n3167 ) | ( n3361  &  n3341  &  n3281 ) ;
 assign n3363 = ( n2993 ) | ( n3352 ) ;
 assign n3362 = ( n3363  &  n3341  &  n3169 ) | ( n3363  &  n3341  &  n3281 ) ;
 assign n3365 = ( n2997  &  n3142 ) | ( n3352  &  n3142 ) | ( n2997  &  n3281 ) | ( n3352  &  n3281 ) ;
 assign n3364 = ( n3365  &  n3341 ) ;
 assign n3367 = ( n3360  &  n3362 ) | ( n891  &  n3362 ) | ( n3360  &  n310 ) | ( n891  &  n310 ) ;
 assign n3366 = ( n188  &  n3367  &  n3364 ) | ( n188  &  n3367  &  n1250 ) ;
 assign n3369 = ( n3174 ) | ( n3281 ) ;
 assign n3368 = ( n3369  &  n3341  &  n3006 ) | ( n3369  &  n3341  &  n3352 ) ;
 assign n3371 = ( n3176 ) | ( n3281 ) ;
 assign n3370 = ( n3371  &  n3341  &  n3012 ) | ( n3371  &  n3341  &  n3352 ) ;
 assign n3373 = ( n3014  &  n3162 ) | ( n3352  &  n3162 ) | ( n3014  &  n3281 ) | ( n3352  &  n3281 ) ;
 assign n3372 = ( n3373  &  n3341 ) ;
 assign n3375 = ( n3368  &  n3370 ) | ( n891  &  n3370 ) | ( n3368  &  n310 ) | ( n891  &  n310 ) ;
 assign n3374 = ( n188  &  n3375  &  n3372 ) | ( n188  &  n3375  &  n1250 ) ;
 assign n3377 = ( n3098 ) | ( n3352 ) ;
 assign n3376 = ( n3377  &  n3341  &  n3184 ) | ( n3377  &  n3341  &  n3281 ) ;
 assign n3379 = ( n3089 ) | ( n3352 ) ;
 assign n3378 = ( n3379  &  n3341  &  n3190 ) | ( n3379  &  n3341  &  n3281 ) ;
 assign n3381 = ( n3099 ) | ( n3352 ) ;
 assign n3380 = ( n3381  &  n3341  &  n3197 ) | ( n3381  &  n3341  &  n3281 ) ;
 assign n3383 = ( n3090 ) | ( n3352 ) ;
 assign n3382 = ( n3383  &  n3341  &  n3204 ) | ( n3383  &  n3341  &  n3281 ) ;
 assign n3385 = ( n188  &  n3380 ) | ( n188  &  n3776 ) ;
 assign n3386 = ( n3376  &  n3378 ) | ( n891  &  n3378 ) | ( n3376  &  n310 ) | ( n891  &  n310 ) ;
 assign n3384 = ( n3385  &  n3386  &  n3382 ) | ( n3385  &  n3386  &  n1692 ) ;
 assign n3388 = ( n3212 ) | ( n3281 ) ;
 assign n3387 = ( n3388  &  n3341  &  n3101 ) | ( n3388  &  n3341  &  n3352 ) ;
 assign n3390 = ( n3217 ) | ( n3281 ) ;
 assign n3389 = ( n3390  &  n3341  &  n3092 ) | ( n3390  &  n3341  &  n3352 ) ;
 assign n3392 = ( n3224 ) | ( n3281 ) ;
 assign n3391 = ( n3392  &  n3341  &  n3102 ) | ( n3392  &  n3341  &  n3352 ) ;
 assign n3394 = ( n3231 ) | ( n3281 ) ;
 assign n3393 = ( n3394  &  n3341  &  n3093 ) | ( n3394  &  n3341  &  n3352 ) ;
 assign n3396 = ( n188  &  n3391 ) | ( n188  &  n3776 ) ;
 assign n3397 = ( n3387  &  n3389 ) | ( n891  &  n3389 ) | ( n3387  &  n310 ) | ( n891  &  n310 ) ;
 assign n3395 = ( n3396  &  n3397  &  n3393 ) | ( n3396  &  n3397  &  n1692 ) ;
 assign n3399 = ( n3044 ) | ( n3352 ) ;
 assign n3398 = ( n3399  &  n3341  &  n3237 ) | ( n3399  &  n3341  &  n3281 ) ;
 assign n3401 = ( n3019 ) | ( n3352 ) ;
 assign n3400 = ( n3401  &  n3341  &  n3240 ) | ( n3401  &  n3341  &  n3281 ) ;
 assign n3403 = ( n3049 ) | ( n3352 ) ;
 assign n3402 = ( n3403  &  n3341  &  n3242 ) | ( n3403  &  n3341  &  n3281 ) ;
 assign n3405 = ( n3026 ) | ( n3352 ) ;
 assign n3404 = ( n3405  &  n3341  &  n3244 ) | ( n3405  &  n3341  &  n3281 ) ;
 assign n3407 = ( n188  &  n3402 ) | ( n188  &  n3776 ) ;
 assign n3408 = ( n3398  &  n3400 ) | ( n891  &  n3400 ) | ( n3398  &  n310 ) | ( n891  &  n310 ) ;
 assign n3406 = ( n3407  &  n3408  &  n3404 ) | ( n3407  &  n3408  &  n1692 ) ;
 assign n3410 = ( n3249 ) | ( n3281 ) ;
 assign n3409 = ( n3410  &  n3341  &  n3052 ) | ( n3410  &  n3341  &  n3352 ) ;
 assign n3412 = ( n3251 ) | ( n3281 ) ;
 assign n3411 = ( n3412  &  n3341  &  n3029 ) | ( n3412  &  n3341  &  n3352 ) ;
 assign n3414 = ( n3253 ) | ( n3281 ) ;
 assign n3413 = ( n3414  &  n3341  &  n3058 ) | ( n3414  &  n3341  &  n3352 ) ;
 assign n3416 = ( n3255 ) | ( n3281 ) ;
 assign n3415 = ( n3416  &  n3341  &  n3034 ) | ( n3416  &  n3341  &  n3352 ) ;
 assign n3418 = ( n188  &  n3413 ) | ( n188  &  n3776 ) ;
 assign n3419 = ( n3409  &  n3411 ) | ( n891  &  n3411 ) | ( n3409  &  n310 ) | ( n891  &  n310 ) ;
 assign n3417 = ( n3418  &  n3419  &  n3415 ) | ( n3418  &  n3419  &  n1692 ) ;
 assign n3421 = ( n1866 ) | ( n3427 ) ;
 assign n3420 = ( n2993  &  n3362  &  (~ n3442) ) | ( n3362  &  n3421  &  (~ n3442) ) ;
 assign n3424 = ( n2980 ) | ( n3421 ) ;
 assign n3425 = ( (~ n169)  &  n3060 ) ;
 assign n3423 = ( n3424  &  n3425  &  n3360 ) | ( n3424  &  n3425  &  n1480 ) ;
 assign n3428 = ( Pi25 ) | ( (~ n193) ) ;
 assign n3427 = ( Pi25 ) | ( n3865 ) ;
 assign n3426 = ( n3428  &  n3364  &  n2997 ) | ( n3428  &  n3364  &  n3427 ) ;
 assign n3431 = ( n3423  &  n3420 ) | ( n2995  &  n3420 ) | ( n3423  &  n2996 ) | ( n2995  &  n2996 ) ;
 assign n3430 = ( (~ Pi22) ) | ( (~ n3001) ) ;
 assign n3429 = ( n188  &  n3431  &  n3426 ) | ( n188  &  n3431  &  n3430 ) ;
 assign n3432 = ( n3428  &  n3372  &  n3014 ) | ( n3428  &  n3372  &  n3427 ) ;
 assign n3433 = ( (~ n2995)  &  (~ n3425) ) | ( (~ n2995)  &  (~ n4632) ) ;
 assign n3438 = ( n2996  &  (~ n3433) ) | ( (~ n3433)  &  (~ n3442)  &  n4633 ) ;
 assign n3437 = ( n188  &  n3438  &  n3432 ) | ( n188  &  n3438  &  n3430 ) ;
 assign n3439 = ( n3019  &  n3400  &  (~ n3442) ) | ( n3400  &  n3421  &  (~ n3442) ) ;
 assign n3440 = ( n3026  &  n3404  &  (~ n3442) ) | ( n3404  &  n3421  &  (~ n3442) ) ;
 assign n3442 = ( n169 ) | ( n3869 ) ;
 assign n3441 = ( n3442  &  (~ n3582) ) | ( (~ n3582)  &  (~ n4643) ) ;
 assign n3444 = ( n3442  &  (~ n3576) ) | ( (~ n3576)  &  (~ n4644) ) ;
 assign n3446 = ( (~ n1884)  &  (~ n3425) ) | ( (~ n1884)  &  (~ n4635) ) ;
 assign n3448 = ( (~ n3425)  &  (~ n3582) ) | ( (~ n3582)  &  (~ n4637) ) ;
 assign n3450 = ( n3073  &  n3345  &  (~ n3442) ) | ( n3345  &  n3421  &  (~ n3442) ) ;
 assign n3452 = ( n3071 ) | ( n3421 ) ;
 assign n3451 = ( n3452  &  n3425  &  n3343 ) | ( n3452  &  n3425  &  n1480 ) ;
 assign n3453 = ( n3428  &  n3347  &  n3076 ) | ( n3428  &  n3347  &  n3427 ) ;
 assign n3455 = ( n3451  &  n3450 ) | ( n2995  &  n3450 ) | ( n3451  &  n2996 ) | ( n2995  &  n2996 ) ;
 assign n3454 = ( n188  &  n3455  &  n3453 ) | ( n188  &  n3455  &  n3430 ) ;
 assign n3456 = ( n3428  &  n3356  &  n3085 ) | ( n3428  &  n3356  &  n3427 ) ;
 assign n3457 = ( (~ n2995)  &  (~ n3425) ) | ( (~ n2995)  &  (~ n4616) ) ;
 assign n3460 = ( n2996  &  (~ n3457) ) | ( (~ n3442)  &  (~ n3457)  &  n4617 ) ;
 assign n3459 = ( n188  &  n3460  &  n3456 ) | ( n188  &  n3460  &  n3430 ) ;
 assign n3461 = ( n3089  &  n3378  &  (~ n3442) ) | ( n3378  &  n3421  &  (~ n3442) ) ;
 assign n3462 = ( n3090  &  n3382  &  (~ n3442) ) | ( n3382  &  n3421  &  (~ n3442) ) ;
 assign n3463 = ( n3442  &  (~ n3582) ) | ( (~ n3582)  &  (~ n4627) ) ;
 assign n3465 = ( n3442  &  (~ n3576) ) | ( (~ n3576)  &  (~ n4628) ) ;
 assign n3467 = ( (~ n1884)  &  (~ n3425) ) | ( (~ n1884)  &  (~ n4619) ) ;
 assign n3469 = ( (~ n3425)  &  (~ n3582) ) | ( (~ n3582)  &  (~ n4621) ) ;
 assign n3472 = ( (~ Pi17)  &  (~ n4777) ) | ( (~ n4650)  &  (~ n4777) ) | ( (~ n4652)  &  (~ n4777) ) ;
 assign n3471 = ( (~ Ni10)  &  (~ n3113)  &  (~ n4779) ) | ( (~ n3113)  &  n3472  &  (~ n4779) ) ;
 assign n3477 = ( (~ Ni33)  &  n3540 ) | ( (~ Ni33)  &  (~ n3951) ) | ( (~ n3540)  &  (~ n3951) ) ;
 assign n3476 = ( n3540 ) | ( n3659 ) ;
 assign n3474 = ( (~ n3948)  &  n4654 ) | ( (~ n1068)  &  (~ Ni13)  &  n4654 ) ;
 assign n3480 = ( (~ Ni47) ) | ( (~ n2959) ) ;
 assign n3478 = ( Pi20  &  (~ n292)  &  n3480 ) | ( (~ n292)  &  (~ n2959)  &  n3480 ) ;
 assign n3482 = ( Ni30 ) | ( n178 ) ;
 assign n3486 = ( Ni47  &  n178 ) | ( Ni47  &  Ni30 ) ;
 assign n3487 = ( n837  &  Ni30 ) ;
 assign n3489 = ( n953  &  Ni30 ) ;
 assign n3490 = ( Ni12 ) | ( (~ n3568) ) ;
 assign n3488 = ( n3487  &  n3489 ) | ( n3487  &  n3490 ) ;
 assign n3492 = ( n836  &  Ni30 ) ;
 assign n3495 = ( n1069  &  n1068  &  n1090 ) ;
 assign n3496 = ( n4797  &  Ni12 ) | ( n4797  &  n3503 ) ;
 assign n3494 = ( (~ Pi26)  &  n3875 ) ;
 assign n3493 = ( n3495  &  n3496  &  Ni14 ) | ( n3495  &  n3496  &  n3494 ) ;
 assign n3500 = ( n3702  &  n3699 ) | ( n3525  &  n3699 ) | ( n3702  &  n2312 ) | ( n3525  &  n2312 ) ;
 assign n3501 = ( n3495  &  (~ n3703) ) | ( Pi24  &  n3489  &  (~ n3703) ) ;
 assign n3498 = ( n3524  &  Pi26 ) | ( n3524  &  n3489 ) ;
 assign n3499 = ( n931 ) | ( (~ Ni11) ) ;
 assign n3497 = ( n3500  &  n3501  &  n3498 ) | ( n3500  &  n3501  &  n3499 ) ;
 assign n3503 = ( Pi26  &  n3875 ) ;
 assign n3502 = ( n3494  &  n3503 ) | ( n2312  &  n3503 ) | ( n3494  &  n3499 ) | ( n2312  &  n3499 ) ;
 assign n3504 = ( n160  &  (~ n3525)  &  (~ n4836) ) | ( (~ n3525)  &  (~ n3702)  &  (~ n4836) ) ;
 assign n3510 = ( (~ Pi23)  &  n3700 ) | ( n3495  &  n3502  &  n3700 ) ;
 assign n3508 = ( (~ Pi24)  &  n3489 ) ;
 assign n3507 = ( n3495  &  (~ n3504)  &  n3510 ) | ( (~ n3504)  &  n3510  &  n3508 ) ;
 assign n3511 = ( n168  &  (~ n3525)  &  (~ n4836) ) | ( (~ n3525)  &  (~ n3702)  &  (~ n4836) ) ;
 assign n3514 = ( n3700  &  Pi23 ) | ( n3700  &  n3495  &  n3502 ) ;
 assign n3512 = ( n3495  &  (~ n3511)  &  n3514 ) | ( n3508  &  (~ n3511)  &  n3514 ) ;
 assign n3516 = ( Ni7 ) | ( Ni8 ) ;
 assign n3515 = ( n3516  &  n1215  &  Ni8 ) | ( n3516  &  n1215  &  Ni10 ) ;
 assign n3518 = ( n3512  &  n3493 ) | ( n3612  &  n3493 ) | ( n3512  &  n3515 ) | ( n3612  &  n3515 ) ;
 assign n3519 = ( n3507  &  n3497 ) | ( n3824  &  n3497 ) | ( n3507  &  n1644 ) | ( n3824  &  n1644 ) ;
 assign n3517 = ( n3518  &  n3519 ) ;
 assign n3520 = ( (~ Ni6)  &  (~ n3517) ) | ( (~ Ni5)  &  (~ n3517) ) ;
 assign n3526 = ( Pi26 ) | ( n3702 ) | ( n2312 ) ;
 assign n3524 = ( (~ Pi27)  &  n3487 ) | ( n3487  &  n3489 ) ;
 assign n3525 = ( (~ Ni12) ) | ( n2456 ) ;
 assign n3523 = ( n3526  &  n3488  &  n3524 ) | ( n3526  &  n3488  &  n3525 ) ;
 assign n3528 = ( (~ Pi26)  &  n3487 ) | ( n3487  &  n3499 ) | ( n3487  &  n3702 ) ;
 assign n3529 = ( n4657  &  n4658  &  n3492 ) | ( n4657  &  n4658  &  n3876 ) ;
 assign n3527 = ( n3528  &  n3529  &  Ni11 ) | ( n3528  &  n3529  &  n3523 ) ;
 assign n3530 = ( Ni32  &  n178 ) | ( n178  &  n2045 ) | ( Ni32  &  (~ Ni41) ) | ( n2045  &  (~ Ni41) ) ;
 assign n3531 = ( (~ Ni31)  &  (~ Ni5) ) | ( (~ Ni6)  &  (~ Ni5) ) | ( (~ Ni5)  &  (~ n3874) ) ;
 assign n3533 = ( n145  &  (~ n3540) ) | ( (~ Ni6)  &  (~ n3517)  &  (~ n3540) ) ;
 assign n3535 = ( Ni4 ) | ( n3545 ) ;
 assign n3534 = ( Ni31  &  (~ n3533)  &  (~ Ni2) ) | ( (~ n3533)  &  n3535  &  (~ Ni2) ) ;
 assign n3538 = ( n3530  &  Ni30 ) ;
 assign n3540 = ( Ni2 ) | ( Ni3 ) ;
 assign n3539 = ( n837  &  (~ n3527) ) | ( (~ n3527)  &  n3535 ) | ( n837  &  n3540 ) | ( n3535  &  n3540 ) ;
 assign n3542 = ( n3531 ) | ( n3545 ) | ( (~ Ni4) ) | ( (~ n4799) ) ;
 assign n3543 = ( (~ Ni5)  &  n3538 ) | ( n3534  &  n3538 ) | ( (~ Ni5)  &  n3877 ) | ( n3534  &  n3877 ) ;
 assign n3545 = ( Ni2 ) | ( (~ Ni3) ) ;
 assign n3544 = ( (~ n3527)  &  n3545 ) | ( n3540  &  n3545 ) | ( (~ n3527)  &  (~ n4659) ) | ( n3540  &  (~ n4659) ) ;
 assign n3548 = ( (~ n145)  &  n3874 ) | ( n3540  &  n3874 ) | ( (~ n145)  &  n3877 ) | ( n3540  &  n3877 ) ;
 assign n3550 = ( (~ Ni9)  &  (~ Ni7) ) ;
 assign n3549 = ( (~ n3540)  &  (~ n3844) ) | ( (~ n3540)  &  n3550  &  (~ n3613) ) ;
 assign n3554 = ( (~ n168)  &  n3516 ) | ( n3516  &  (~ Ni7) ) | ( (~ n168)  &  n3837 ) | ( (~ Ni7)  &  n3837 ) ;
 assign n3553 = ( Pi24  &  n3554 ) | ( (~ Ni8)  &  n3554 ) ;
 assign n3555 = ( (~ Ni10) ) | ( n3540 ) | ( n3553 ) | ( (~ n3844) ) ;
 assign n3556 = ( (~ n160)  &  (~ Ni9) ) | ( Ni10  &  (~ Ni9) ) ;
 assign n3557 = ( n138  &  (~ Ni8) ) | ( n3516  &  (~ Ni8) ) | ( n138  &  n3556 ) | ( n3516  &  n3556 ) ;
 assign n3558 = ( Ni10  &  n3557 ) | ( n3557  &  (~ Ni7) ) | ( Ni10  &  (~ n3844) ) | ( (~ Ni7)  &  (~ n3844) ) ;
 assign n3560 = ( Pi27  &  (~ n161) ) | ( Pi27  &  Ni14 ) | ( (~ n161)  &  (~ Ni14) ) ;
 assign n3559 = ( (~ Ni11)  &  (~ Ni13)  &  n3560 ) ;
 assign n3563 = ( n157  &  (~ Ni11) ) | ( (~ Ni11)  &  n1068 ) | ( n157  &  (~ n3603) ) | ( n1068  &  (~ n3603) ) ;
 assign n3561 = ( Pi27  &  n3563 ) | ( (~ Ni12)  &  n3563 ) ;
 assign n3564 = ( (~ Ni14) ) | ( n3540 ) | ( n3561 ) | ( (~ n3568) ) ;
 assign n3568 = ( (~ Ni14) ) | ( (~ Ni13) ) ;
 assign n3566 = ( n161  &  (~ Ni14)  &  Ni12 ) ;
 assign n3567 = ( n157  &  Ni14  &  (~ n1068) ) ;
 assign n3565 = ( n3568  &  n3566 ) | ( n3568  &  n3567 ) | ( n3568  &  Ni13 ) ;
 assign n3569 = ( (~ n3540)  &  n3565 ) | ( Ni11  &  (~ Ni14)  &  (~ n3540) ) ;
 assign n3573 = ( (~ Ni42) ) | ( (~ Ni43) ) ;
 assign n3572 = ( Ni44 ) | ( (~ Ni43) ) ;
 assign n3571 = ( n3573  &  n2078 ) | ( n3573  &  n3572 ) ;
 assign n3574 = ( (~ Ni41) ) | ( (~ Ni43) ) ;
 assign n3577 = ( n3579  &  n3706 ) | ( n3706  &  (~ Ni43) ) | ( n3579  &  n3777 ) | ( (~ Ni43)  &  n3777 ) ;
 assign n3576 = ( (~ Pi16) ) | ( n796 ) ;
 assign n3575 = ( n3571  &  n3577  &  n3574 ) | ( n3571  &  n3577  &  n3576 ) ;
 assign n3580 = ( n3576  &  n3706 ) | ( n3706  &  (~ Ni43) ) | ( n3576  &  n3778 ) | ( (~ Ni43)  &  n3778 ) ;
 assign n3579 = ( (~ Pi16) ) | ( n3735 ) ;
 assign n3578 = ( n3571  &  n3580  &  n3574 ) | ( n3571  &  n3580  &  n3579 ) ;
 assign n3583 = ( n3575  &  n3578 ) | ( n3575  &  Ni40 ) | ( n3578  &  (~ Ni40) ) ;
 assign n3582 = ( (~ Pi16) ) | ( n3738 ) ;
 assign n3581 = ( n3583  &  n3574 ) | ( n3583  &  n3582 ) ;
 assign n3585 = ( (~ Ni44) ) | ( (~ Ni43) ) ;
 assign n3584 = ( n3573  &  n2078 ) | ( n3573  &  n3585 ) ;
 assign n3586 = ( n3584  &  n3577  &  n3574 ) | ( n3584  &  n3577  &  n3576 ) ;
 assign n3587 = ( n3584  &  n3580  &  n3574 ) | ( n3584  &  n3580  &  n3579 ) ;
 assign n3589 = ( n3586  &  n3587 ) | ( n3586  &  Ni40 ) | ( n3587  &  (~ Ni40) ) ;
 assign n3588 = ( n3589  &  n3574 ) | ( n3589  &  n3582 ) ;
 assign n3592 = ( Ni31 ) | ( n153 ) ;
 assign n3590 = ( (~ n1965)  &  (~ n3618) ) | ( (~ n1965)  &  n3706 ) | ( (~ n3618)  &  (~ Ni43) ) | ( n3706  &  (~ Ni43) ) ;
 assign n3591 = ( Pi20  &  n3581 ) | ( (~ Pi20)  &  n3588 ) | ( n3581  &  n3588 ) ;
 assign n3593 = ( Ni42 ) | ( (~ Ni43) ) ;
 assign n3595 = ( n2078 ) | ( (~ Ni40) ) ;
 assign n3594 = ( n3572 ) | ( n3595 ) ;
 assign n3596 = ( n3594 ) | ( Ni30  &  (~ n3879) ) ;
 assign n3597 = ( (~ Ni31)  &  n178 ) | ( n178  &  n276 ) | ( (~ Ni31)  &  Ni41 ) | ( n276  &  Ni41 ) ;
 assign N_N13958 = ( (~ n3545) ) ;
 assign n3598 = ( (~ n2066)  &  (~ n3530)  &  (~ n3545)  &  Ni4 ) ;
 assign n3603 = ( Pi27 ) | ( (~ Pi26) ) ;
 assign n3601 = ( (~ Ni12)  &  n3499 ) | ( n3499  &  (~ n3559) ) | ( (~ Ni12)  &  n3603 ) | ( (~ n3559)  &  n3603 ) ;
 assign n3604 = ( n3598  &  (~ n3640) ) | ( (~ n3597)  &  (~ n3640)  &  (~ n3877) ) ;
 assign n3608 = ( Ni30 ) | ( n2066 ) | ( n3535 ) | ( (~ n3863) ) ;
 assign n3610 = ( (~ Ni32)  &  n276 ) | ( n276  &  Ni41 ) ;
 assign n3612 = ( (~ Ni10) ) | ( n1654 ) | ( (~ Ni7) ) ;
 assign n3613 = ( (~ Pi24)  &  n160 ) | ( (~ Pi24)  &  Ni10 ) | ( n160  &  (~ Ni10) ) ;
 assign n3614 = ( (~ Ni8) ) | ( Ni9 ) | ( Ni7 ) ;
 assign n3611 = ( n168  &  n3613 ) | ( n3612  &  n3613 ) | ( n168  &  n3614 ) | ( n3612  &  n3614 ) ;
 assign n3615 = ( n2066 ) | ( n3545 ) | ( n4817 ) | ( n4818 ) ;
 assign n3616 = ( n837 ) | ( n3877 ) | ( Ni33 ) | ( n3610 ) ;
 assign n3618 = ( (~ Pi16)  &  n2939 ) ;
 assign n3617 = ( n1965  &  (~ n3260) ) | ( (~ n3260)  &  n3618 ) ;
 assign Nv437 = ( n2053 ) | ( n2056 ) | ( n2063 ) | ( (~ n4334) ) ;
 assign n3620 = ( Pi21  &  (~ n2064)  &  n3665 ) | ( n178  &  (~ n2064)  &  n3665 ) ;
 assign Nv43 = ( (~ n3620) ) ;
 assign n3621 = ( n292  &  (~ Ni47)  &  n3698 ) | ( n292  &  (~ n3545)  &  n3698 ) ;
 assign Nv14 = ( (~ n3621) ) ;
 assign n3622 = ( n3708  &  (~ n3965) ) | ( n23  &  Ni30  &  n3708 ) ;
 assign n3623 = ( (~ Pi16)  &  (~ n184)  &  Ni41  &  (~ n3593) ) ;
 assign n3624 = ( Pi20  &  n3712  &  (~ n4810) ) | ( (~ n3596)  &  n3712  &  (~ n4810) ) ;
 assign N_N13959 = ( n3622 ) | ( n3623 ) | ( n3624 ) ;
 assign n3626 = ( Pi20  &  (~ n298) ) | ( (~ Pi21)  &  Pi20  &  (~ n541) ) ;
 assign n3627 = ( (~ Pi20)  &  (~ n298) ) | ( (~ Pi21)  &  (~ Pi20)  &  (~ n516) ) ;
 assign n3628 = ( Pi20  &  (~ n298) ) | ( (~ Pi21)  &  Pi20  &  (~ n701) ) ;
 assign n3629 = ( (~ Pi20)  &  (~ n298) ) | ( (~ Pi21)  &  (~ Pi20)  &  (~ n689) ) ;
 assign n3631 = ( Pi20  &  (~ n298) ) | ( (~ Pi21)  &  Pi20  &  (~ n637) ) ;
 assign n3632 = ( (~ Pi20)  &  (~ n298) ) | ( (~ Pi21)  &  (~ Pi20)  &  (~ n613) ) ;
 assign n3630 = ( (~ n295) ) | ( n653 ) | ( n3631 ) | ( n3632 ) ;
 assign n3634 = ( Pi20  &  (~ n298) ) | ( (~ Pi21)  &  Pi20  &  (~ n741) ) ;
 assign n3635 = ( (~ Pi20)  &  (~ n298) ) | ( (~ Pi21)  &  (~ Pi20)  &  (~ n734) ) ;
 assign n3633 = ( (~ n295) ) | ( n749 ) | ( n3634 ) | ( n3635 ) ;
 assign n3638 = ( n1062  &  n836 ) ;
 assign n3639 = ( (~ Pi27)  &  n3638 ) | ( n1470  &  n3638 ) ;
 assign n3640 = ( (~ Ni30) ) | ( (~ Ni33) ) ;
 assign n3641 = ( (~ n161)  &  n836 ) | ( (~ Ni30)  &  n836 ) ;
 assign n3643 = ( (~ n161)  &  n837 ) | ( n837  &  n953 ) ;
 assign n3646 = ( (~ Pi21)  &  (~ n3641) ) ;
 assign n3647 = ( (~ Pi22)  &  (~ n3641) ) ;
 assign n3645 = ( (~ Pi24)  &  n3646 ) | ( (~ Pi24)  &  n3647 ) | ( (~ Pi24)  &  (~ n4233) ) ;
 assign n3649 = ( Pi27  &  n836 ) | ( (~ Ni30)  &  n836 ) ;
 assign n3650 = ( n837  &  Pi27 ) | ( n837  &  n953 ) ;
 assign n3653 = ( Pi24  &  Ni14  &  (~ n3649) ) | ( Ni14  &  (~ n3649)  &  (~ n3650) ) ;
 assign n3655 = ( n1062  &  (~ n3653) ) | ( n1866  &  (~ n3653) ) ;
 assign n3659 = ( Ni7 ) | ( n1654 ) ;
 assign n3657 = ( Ni34  &  n3113  &  n3659 ) | ( Ni34  &  n3659  &  (~ n3894) ) ;
 assign n3662 = ( (~ n32) ) | ( Ni33 ) ;
 assign n3660 = ( (~ Pi26)  &  n2024  &  n3662 ) | ( (~ n32)  &  n2024  &  n3662 ) ;
 assign n3663 = ( (~ Pi27)  &  n2043  &  n3662 ) | ( (~ n32)  &  n2043  &  n3662 ) ;
 assign n3665 = ( n296  &  (~ Ni45) ) | ( n296  &  (~ n2066)  &  (~ n3535) ) ;
 assign n3666 = ( n2079  &  Ni42 ) | ( n2079  &  Ni47 ) ;
 assign n3667 = ( n153  &  n195 ) ;
 assign n3668 = ( n176  &  n2074 ) ;
 assign n3671 = ( n3680  &  Pi27 ) | ( n1866  &  Pi27 ) | ( n3680  &  n3678 ) | ( n1866  &  n3678 ) ;
 assign n3670 = ( n178  &  n195 ) ;
 assign n3669 = ( n2333  &  n3671  &  n3670 ) | ( n2333  &  n3671  &  n2328 ) ;
 assign n3672 = ( (~ Pi27)  &  n3668 ) | ( n2754  &  n3668 ) ;
 assign n3674 = ( (~ Pi26)  &  n2303 ) | ( (~ Ni32)  &  n2303 ) ;
 assign n3675 = ( n176  &  n195 ) ;
 assign n3676 = ( (~ Pi27)  &  n3675 ) | ( n3667  &  n3675 ) ;
 assign n3677 = ( (~ Pi26)  &  n3676 ) | ( n3667  &  n3676 ) ;
 assign n3678 = ( n2069  &  n196 ) ;
 assign n3679 = ( (~ Pi27)  &  n3670 ) | ( n194  &  n3670 ) ;
 assign n3680 = ( n178  &  n2074 ) ;
 assign n3681 = ( n2074  &  n196 ) ;
 assign n3682 = ( n3676  &  Pi26 ) | ( n3676  &  n3667 ) ;
 assign n3685 = ( n3859  &  n2950 ) ;
 assign n3684 = ( (~ Pi26)  &  n177  &  n3685 ) | ( n177  &  n3592  &  n3685 ) ;
 assign n3687 = ( n2055  &  n3843 ) ;
 assign n3686 = ( Pi23  &  (~ n3684) ) | ( (~ n3685)  &  (~ n3684) ) | ( (~ n3684)  &  n3687 ) ;
 assign n3691 = ( n3862  &  n2953 ) ;
 assign n3690 = ( (~ Pi27)  &  n177  &  n3691 ) | ( n177  &  n3592  &  n3691 ) ;
 assign n3692 = ( Pi24  &  (~ n3690) ) | ( n3687  &  (~ n3690) ) | ( (~ n3691)  &  (~ n3690) ) ;
 assign n3695 = ( (~ Pi22)  &  n171 ) | ( (~ Pi22)  &  (~ n1063)  &  (~ n2955) ) ;
 assign n3696 = ( (~ Pi21)  &  n171 ) | ( (~ Pi21)  &  (~ n1063)  &  n2947 ) ;
 assign n3697 = ( n2967 ) | ( (~ Ni41) ) ;
 assign n3698 = ( (~ Ni47)  &  (~ n3486) ) | ( (~ n2066)  &  (~ n3486)  &  (~ Ni4) ) ;
 assign n3699 = ( (~ Pi26)  &  n3524 ) | ( n3489  &  n3524 ) ;
 assign n3701 = ( n3699  &  n3498 ) | ( n2312  &  n3498 ) | ( n3699  &  n3499 ) | ( n2312  &  n3499 ) ;
 assign n3700 = ( (~ Pi24)  &  n3701 ) | ( n3502  &  n3701 ) ;
 assign n3702 = ( n3487  &  Pi27 ) | ( n3487  &  n3489 ) ;
 assign n3703 = ( (~ Pi24)  &  (~ n3502) ) | ( (~ Pi24)  &  (~ n3525)  &  (~ n4836) ) ;
 assign n3705 = ( n3492  &  Ni11 ) | ( n3492  &  n3490 ) ;
 assign n3706 = ( Ni41 ) | ( (~ Ni43) ) ;
 assign n3708 = ( Ni30  &  (~ n184) ) | ( (~ n184)  &  (~ n391) ) | ( (~ n184)  &  n3573 ) ;
 assign n3712 = ( Pi18  &  (~ Pi17) ) ;
 assign n3713 = ( n18 ) | ( n1866 ) ;
 assign n3716 = ( n1866 ) | ( (~ n2939) ) ;
 assign n3718 = ( n45  &  (~ Ni47) ) ;
 assign n3719 = ( (~ n18) ) | ( n2065 ) ;
 assign n3721 = ( Ni36 ) | ( n694 ) ;
 assign n3722 = ( Ni37 ) | ( Ni36 ) ;
 assign n3723 = ( Ni38 ) | ( n3722 ) ;
 assign n3724 = ( n3723 ) | ( (~ Ni39) ) ;
 assign n3725 = ( Ni39 ) | ( n3723 ) ;
 assign n3726 = ( Ni32 ) | ( n2087 ) ;
 assign n3727 = ( Pi20 ) | ( n1866 ) ;
 assign n3728 = ( Pi25 ) | ( n3727 ) ;
 assign n3729 = ( (~ Pi20) ) | ( n1866 ) ;
 assign n3731 = ( Pi25 ) | ( n3729 ) ;
 assign n3733 = ( Pi20  &  (~ n298) ) | ( (~ Pi21)  &  Pi20  &  (~ n253) ) ;
 assign n3734 = ( (~ Pi20)  &  (~ n298) ) | ( (~ Pi21)  &  (~ Pi20)  &  (~ n219) ) ;
 assign n3732 = ( (~ n295) ) | ( n303 ) | ( n3733 ) | ( n3734 ) ;
 assign n3735 = ( Pi19 ) | ( (~ Pi17) ) ;
 assign n3736 = ( Pi20  &  (~ n298) ) | ( (~ Pi21)  &  Pi20  &  (~ n487) ) ;
 assign n3737 = ( (~ Pi20)  &  (~ n298) ) | ( (~ Pi21)  &  (~ Pi20)  &  (~ n462) ) ;
 assign n3738 = ( Pi17 ) | ( Pi19 ) ;
 assign n3739 = ( (~ Ni32) ) | ( n2199 ) ;
 assign n3740 = ( Ni32 ) | ( n2199 ) ;
 assign n3742 = ( Pi16 ) | ( Pi15 ) ;
 assign n3747 = ( Pi20  &  (~ n298) ) | ( (~ Pi21)  &  Pi20  &  (~ n408) ) ;
 assign n3748 = ( (~ Pi20)  &  (~ n298) ) | ( (~ Pi21)  &  (~ Pi20)  &  (~ n395) ) ;
 assign n3746 = ( (~ n295) ) | ( n420 ) | ( n3747 ) | ( n3748 ) ;
 assign n3749 = ( n45  &  (~ Ni45) ) ;
 assign n3750 = ( Pi20  &  (~ n298) ) | ( (~ Pi21)  &  Pi20  &  (~ n678) ) ;
 assign n3751 = ( (~ Pi20)  &  (~ n298) ) | ( (~ Pi21)  &  (~ Pi20)  &  (~ n664) ) ;
 assign n3754 = ( Pi16 ) | ( (~ Pi15) ) ;
 assign n3757 = ( Pi20  &  (~ n298) ) | ( (~ Pi21)  &  Pi20  &  (~ n349) ) ;
 assign n3758 = ( (~ Pi20)  &  (~ n298) ) | ( (~ Pi21)  &  (~ Pi20)  &  (~ n325) ) ;
 assign n3756 = ( (~ n295) ) | ( n381 ) | ( n3757 ) | ( n3758 ) ;
 assign n3760 = ( Pi20  &  (~ n298) ) | ( (~ Pi21)  &  Pi20  &  (~ n588) ) ;
 assign n3761 = ( (~ Pi20)  &  (~ n298) ) | ( (~ Pi21)  &  (~ Pi20)  &  (~ n567) ) ;
 assign n3759 = ( (~ n295) ) | ( n656 ) | ( n3760 ) | ( n3761 ) ;
 assign n3763 = ( (~ Pi16) ) | ( Pi15 ) ;
 assign n3767 = ( Pi20  &  (~ n298) ) | ( (~ Pi21)  &  Pi20  &  (~ n435) ) ;
 assign n3768 = ( (~ Pi20)  &  (~ n298) ) | ( (~ Pi21)  &  (~ Pi20)  &  (~ n428) ) ;
 assign n3766 = ( (~ n295) ) | ( n447 ) | ( n3767 ) | ( n3768 ) ;
 assign n3770 = ( Pi20  &  (~ n298) ) | ( (~ Pi21)  &  Pi20  &  (~ n724) ) ;
 assign n3771 = ( (~ Pi20)  &  (~ n298) ) | ( (~ Pi21)  &  (~ Pi20)  &  (~ n714) ) ;
 assign n3769 = ( (~ n295) ) | ( n752 ) | ( n3770 ) | ( n3771 ) ;
 assign n3774 = ( (~ Pi16) ) | ( (~ Pi15) ) ;
 assign n3775 = ( Ni10 ) | ( (~ n3113) ) ;
 assign n3776 = ( (~ Pi19) ) | ( n3727 ) ;
 assign n3777 = ( Pi16 ) | ( n3735 ) ;
 assign n3778 = ( Pi16 ) | ( n796 ) ;
 assign n3779 = ( Ni4 ) | ( Ni5 ) | ( Ni6 ) ;
 assign n3783 = ( Ni11 ) | ( Ni10 ) ;
 assign n3784 = ( n931  &  Ni11 ) ;
 assign n3785 = ( n3716 ) | ( n3603 ) ;
 assign n3786 = ( (~ n3603) ) | ( n3716 ) ;
 assign n3787 = ( n3727 ) | ( n3603 ) ;
 assign n3788 = ( n3729 ) | ( n3603 ) ;
 assign n3789 = ( (~ n3603) ) | ( n3729 ) ;
 assign n3790 = ( Pi27 ) | ( n996 ) ;
 assign n3791 = ( Pi27 ) | ( n998 ) ;
 assign n3792 = ( (~ Pi27) ) | ( n996 ) ;
 assign n3793 = ( (~ Pi27) ) | ( n998 ) ;
 assign n3794 = ( Pi27 ) | ( n3727 ) ;
 assign n3795 = ( Pi27 ) | ( n3729 ) ;
 assign n3796 = ( (~ Pi27) ) | ( n3727 ) ;
 assign n3797 = ( (~ Pi27) ) | ( n3729 ) ;
 assign n3798 = ( Ni13 ) | ( Ni14 ) ;
 assign n3799 = ( n3716 ) | ( n161 ) ;
 assign n3800 = ( (~ n161) ) | ( n3716 ) ;
 assign n3801 = ( n3727 ) | ( n161 ) ;
 assign n3802 = ( n3729 ) | ( n161 ) ;
 assign n3803 = ( (~ n161) ) | ( n3729 ) ;
 assign n3804 = ( n3647 ) | ( n3646 ) ;
 assign n3805 = ( Ni11 ) | ( (~ Ni12) ) ;
 assign n3806 = ( Pi27 ) | ( n1474 ) ;
 assign n3807 = ( (~ Pi27) ) | ( n1474 ) ;
 assign n3808 = ( Pi27 ) | ( n1480 ) ;
 assign n3809 = ( (~ Pi27) ) | ( n1997 ) ;
 assign n3810 = ( n1474 ) | ( n161 ) ;
 assign n3811 = ( (~ n161) ) | ( n1474 ) ;
 assign n3812 = ( n1997 ) | ( n161 ) ;
 assign n3813 = ( n787 ) | ( n161 ) ;
 assign n3814 = ( Ni13 ) | ( n3805 ) ;
 assign n3815 = ( n1474 ) | ( n3603 ) ;
 assign n3816 = ( n1474 ) | ( (~ n3603) ) ;
 assign n3817 = ( n1997 ) | ( n3603 ) ;
 assign n3818 = ( n787 ) | ( n3603 ) ;
 assign n3820 = ( n3716 ) | ( n160 ) ;
 assign n3821 = ( (~ n160) ) | ( n3716 ) ;
 assign n3822 = ( n3727 ) | ( n160 ) ;
 assign n3823 = ( (~ n160) ) | ( n3727 ) ;
 assign n3824 = ( Ni10 ) | ( n3614 ) ;
 assign n3825 = ( (~ Pi24) ) | ( n996 ) ;
 assign n3826 = ( (~ Pi24) ) | ( n998 ) ;
 assign n3827 = ( Pi24 ) | ( n3727 ) ;
 assign n3828 = ( Pi24 ) | ( n3729 ) ;
 assign n3829 = ( (~ Pi24) ) | ( n3727 ) ;
 assign n3830 = ( (~ Pi24) ) | ( n3729 ) ;
 assign n3831 = ( Pi15 ) | ( n3113 ) ;
 assign n3832 = ( n3716 ) | ( n168 ) ;
 assign n3833 = ( (~ n168) ) | ( n3716 ) ;
 assign n3834 = ( n3727 ) | ( n168 ) ;
 assign n3835 = ( (~ n168) ) | ( n3727 ) ;
 assign n3836 = ( (~ Pi25) ) | ( n1662 ) ;
 assign n3837 = ( (~ n18) ) | ( Ni33 ) ;
 assign n3838 = ( (~ Pi25) ) | ( Ni34 ) | ( n1063 ) | ( n3837 ) ;
 assign n3839 = ( n1866 ) | ( n1662 ) ;
 assign n3840 = ( (~ Ni34) ) | ( Ni33 ) ;
 assign n3842 = ( n3839 ) | ( n3840 ) ;
 assign n3841 = ( (~ n163)  &  n1670  &  n3842 ) ;
 assign n3843 = ( Ni32  &  Ni33 ) ;
 assign n3844 = ( (~ Ni10) ) | ( (~ Ni9) ) ;
 assign n3845 = ( Ni31 ) | ( n3640 ) ;
 assign n3846 = ( Ni39 ) | ( n3722 ) ;
 assign n3847 = ( n694 ) | ( (~ Ni38) ) ;
 assign n3848 = ( n3722 ) | ( (~ Ni39) ) ;
 assign n3849 = ( n2025 ) | ( (~ Ni38) ) ;
 assign n3851 = ( n2083  &  n2084  &  n2184 ) ;
 assign n3852 = ( n2083  &  n2099  &  n2190 ) ;
 assign n3854 = ( n2083  &  n2084  &  n2076 ) ;
 assign n3855 = ( n2083  &  n2099  &  n2095 ) ;
 assign n3857 = ( (~ Pi26) ) | ( Pi24 ) ;
 assign n3858 = ( (~ Ni37) ) | ( (~ Ni38) ) ;
 assign n3859 = ( Ni32 ) | ( (~ Ni40) ) ;
 assign n3860 = ( Ni33 ) | ( n3592 ) ;
 assign n3861 = ( (~ Ni33) ) | ( n3592 ) ;
 assign n3862 = ( Ni32 ) | ( (~ Ni41) ) ;
 assign n3863 = ( Ni31  &  Ni33 ) ;
 assign n3864 = ( Ni38 ) | ( n2964 ) ;
 assign n3865 = ( Ni33 ) | ( n1063 ) ;
 assign n3866 = ( Ni38 ) | ( n2967 ) ;
 assign n3869 = ( n3695 ) | ( n3696 ) ;
 assign n3870 = ( (~ Pi17) ) | ( Pi16 ) ;
 assign n3871 = ( (~ Pi17) ) | ( (~ Pi16) ) ;
 assign n3874 = ( (~ Ni30) ) | ( n3530 ) ;
 assign n3875 = ( (~ Pi27)  &  n3492 ) ;
 assign n3876 = ( n3516 ) | ( (~ n3844) ) ;
 assign n3877 = ( Ni6 ) | ( (~ Ni5) ) | ( n3535 ) ;
 assign n3879 = ( (~ Ni32)  &  Ni30 ) ;
 assign n3880 = ( n3540 ) | ( n2031 ) ;
 assign n3881 = ( Ni7 ) | ( n3540 ) | ( n2049 ) ;
 assign n3882 = ( (~ n18)  &  (~ n4673) ) | ( (~ n3540)  &  (~ n4673) ) ;
 assign Nv8909 = ( (~ n3882) ) ;
 assign n3886 = ( Ni10  &  (~ n1265) ) | ( (~ Ni10)  &  (~ n1522) ) | ( (~ n1265)  &  (~ n1522) ) ;
 assign n3887 = ( (~ Pi15)  &  n4678 ) | ( Pi15  &  n4682 ) | ( n4678  &  n4682 ) ;
 assign n3888 = ( (~ Pi17)  &  (~ n4696) ) | ( (~ n4091)  &  (~ n4696) ) | ( (~ n4093)  &  (~ n4696) ) ;
 assign n3890 = ( Ni10  &  (~ n4693) ) | ( (~ n4116)  &  (~ n4693) ) | ( (~ n4119)  &  (~ n4693) ) ;
 assign n3891 = ( n1062  &  n3643  &  (~ n3645) ) | ( n1866  &  n3643  &  (~ n3645) ) ;
 assign n3893 = ( (~ Ni10)  &  n4713 ) | ( n1990  &  n4713 ) ;
 assign n3894 = ( (~ Pi17)  &  (~ n4714) ) | ( n4330  &  n4331  &  (~ n4714) ) ;
 assign n3898 = ( Ni10  &  (~ n2579) ) | ( (~ Ni10)  &  (~ n2799) ) | ( (~ n2579)  &  (~ n2799) ) ;
 assign n3899 = ( (~ Pi15)  &  n4740 ) | ( Pi15  &  n4743 ) | ( n4740  &  n4743 ) ;
 assign n3900 = ( (~ Pi17)  &  (~ n4756) ) | ( (~ n4396)  &  (~ n4756) ) | ( (~ n4398)  &  (~ n4756) ) ;
 assign n3901 = ( (~ Pi27)  &  (~ Pi22)  &  (~ n3667) ) | ( (~ Pi22)  &  (~ n3667)  &  (~ n3675) ) ;
 assign n3905 = ( (~ Ni14)  &  (~ n4738) ) | ( (~ n4412)  &  (~ n4738) ) | ( (~ n4414)  &  (~ n4738) ) ;
 assign n3908 = ( n4120  &  Ni11 ) | ( n2799  &  Ni11 ) | ( n4120  &  n2797 ) | ( n2799  &  n2797 ) ;
 assign n3906 = ( (~ n2913)  &  n3814  &  n3908 ) | ( (~ n2913)  &  (~ n3905)  &  n3908 ) ;
 assign n3910 = ( Pi23  &  (~ n2304) ) | ( (~ Pi23)  &  n4755 ) | ( (~ n2304)  &  n4755 ) ;
 assign n3912 = ( n160  &  (~ n2308) ) | ( (~ n160)  &  (~ n3669) ) | ( (~ n2308)  &  (~ n3669) ) ;
 assign n3914 = ( (~ Pi24)  &  (~ n2308) ) | ( Pi24  &  (~ n3669) ) | ( (~ n2308)  &  (~ n3669) ) ;
 assign n3916 = ( (~ Pi24)  &  (~ n2304) ) | ( Pi24  &  n4733 ) | ( (~ n2304)  &  n4733 ) ;
 assign n3918 = ( (~ Pi24)  &  (~ n2314) ) | ( Pi24  &  n4737 ) | ( (~ n2314)  &  n4737 ) ;
 assign n3920 = ( (~ Pi23)  &  (~ n2304) ) | ( Pi23  &  n4755 ) | ( (~ n2304)  &  n4755 ) ;
 assign n3922 = ( n168  &  (~ n2308) ) | ( (~ n168)  &  (~ n3669) ) | ( (~ n2308)  &  (~ n3669) ) ;
 assign n3923 = ( n2923  &  n3779 ) | ( n2926  &  n3779 ) | ( n3779  &  (~ n4562) ) ;
 assign n3926 = ( (~ Pi23)  &  n3859 ) | ( n3859  &  n3860 ) ;
 assign n3925 = ( n2950  &  (~ Ni40)  &  n3926 ) | ( n2950  &  n3861  &  n3926 ) ;
 assign n3928 = ( n4761  &  n2031 ) | ( n4761  &  n4565  &  n3685 ) ;
 assign n3930 = ( n2049  &  (~ n3928) ) | ( (~ n2049)  &  n4763 ) | ( (~ n3928)  &  n4763 ) ;
 assign n3932 = ( (~ Pi24)  &  n3862 ) | ( n3860  &  n3862 ) ;
 assign n3931 = ( n2953  &  (~ Ni41)  &  n3932 ) | ( n2953  &  n3861  &  n3932 ) ;
 assign n3934 = ( n4764  &  n2031 ) | ( n4764  &  n4566  &  n3691 ) ;
 assign n3936 = ( n2049  &  (~ n3934) ) | ( (~ n2049)  &  n4766 ) | ( (~ n3934)  &  n4766 ) ;
 assign n3938 = ( n3576  &  (~ n3617) ) | ( n3260  &  (~ n3617)  &  n4584 ) ;
 assign n3939 = ( (~ n3268)  &  n3778 ) | ( n3260  &  (~ n3268)  &  n4582 ) ;
 assign n3940 = ( (~ n3265)  &  n3579 ) | ( n3260  &  (~ n3265)  &  n4580 ) ;
 assign n3941 = ( n4585  &  n3777 ) | ( n4585  &  n4579  &  n3260 ) ;
 assign n3937 = ( n3938  &  n3939  &  n3940  &  n3941 ) ;
 assign n3943 = ( n3576  &  (~ n3617) ) | ( n3260  &  (~ n3617)  &  n4608 ) ;
 assign n3944 = ( (~ n3332)  &  n3778 ) | ( n3260  &  (~ n3332)  &  n4606 ) ;
 assign n3945 = ( (~ n3330)  &  n3579 ) | ( n3260  &  (~ n3330)  &  n4604 ) ;
 assign n3946 = ( n4609  &  n3777 ) | ( n4609  &  n4603  &  n3260 ) ;
 assign n3942 = ( n3943  &  n3944  &  n3945  &  n3946 ) ;
 assign n3948 = ( (~ Ni10)  &  (~ n4792) ) | ( (~ n4790)  &  (~ n4791)  &  (~ n4792) ) ;
 assign n3949 = ( Pi20  &  n3095 ) | ( (~ Pi20)  &  n3104 ) | ( n3095  &  n3104 ) ;
 assign n3950 = ( Pi20  &  n3038 ) | ( (~ Pi20)  &  n3061 ) | ( n3038  &  n3061 ) ;
 assign n3951 = ( n3659  &  n3111 ) | ( n3659  &  n3114 ) | ( n3659  &  n3116 ) ;
 assign n3953 = ( n145 ) | ( n3520 ) | ( (~ Ni4) ) ;
 assign n3952 = ( Ni5  &  n3953  &  (~ n4798) ) | ( (~ n3517)  &  n3953  &  (~ n4798) ) ;
 assign n3955 = ( (~ Ni4)  &  (~ n4803) ) | ( (~ Ni2)  &  (~ n4803) ) ;
 assign Nv10316 = ( (~ n3955) ) ;
 assign n3957 = ( (~ Ni8) ) | ( (~ Ni7) ) | ( n3844 ) ;
 assign n3958 = ( n168  &  n3516 ) | ( (~ Ni10)  &  n3516 ) | ( n1654  &  n3516 ) ;
 assign n3956 = ( Ni7  &  n3957  &  n3958 ) | ( (~ n3844)  &  n3957  &  n3958 ) ;
 assign n3959 = ( n3540  &  (~ Ni7) ) | ( (~ n3540)  &  (~ n3956) ) | ( (~ Ni7)  &  (~ n3956) ) ;
 assign Nv10135 = ( (~ n3959) ) ;
 assign n3960 = ( (~ Ni10)  &  n3540 ) | ( (~ Ni10)  &  n3558 ) | ( (~ n3540)  &  n3558 ) ;
 assign Nv10099 = ( (~ n3960) ) ;
 assign n3962 = ( Ni11  &  n1069 ) | ( Ni11  &  n3568 ) | ( n1069  &  (~ n3568) ) ;
 assign n3961 = ( n1068  &  n3962  &  n931 ) | ( n1068  &  n3962  &  n3603 ) ;
 assign n3963 = ( (~ Ni11)  &  n3540 ) | ( (~ Ni11)  &  (~ n3961) ) | ( (~ n3540)  &  (~ n3961) ) ;
 assign Nv10091 = ( (~ n3963) ) ;
 assign n3964 = ( Ni12  &  (~ n4808) ) | ( n3540  &  (~ n4808) ) | ( n3568  &  (~ n4808) ) ;
 assign Nv10082 = ( (~ n3964) ) ;
 assign n3965 = ( (~ n3572)  &  (~ n4811) ) | ( (~ Ni42)  &  (~ n4811) ) | ( (~ Ni39)  &  (~ n4811) ) ;
 assign n3966 = ( (~ Pi26)  &  n4814 ) | ( n4813  &  n4814 ) ;
 assign n3967 = ( (~ Pi23)  &  n4816 ) | ( n4815  &  n4816 ) ;
 assign n3968 = ( n232  &  n265 ) | ( n3727  &  n265 ) | ( n232  &  n3729 ) | ( n3727  &  n3729 ) ;
 assign n3969 = ( n336  &  n360 ) | ( n3727  &  n360 ) | ( n336  &  n3729 ) | ( n3727  &  n3729 ) ;
 assign n3970 = ( n470 ) | ( (~ Ni37)  &  n202 ) ;
 assign n3971 = ( n463 ) | ( (~ Ni37)  &  n202 ) ;
 assign n3972 = ( n494 ) | ( (~ Ni37)  &  n240 ) ;
 assign n3973 = ( n488 ) | ( (~ Ni37)  &  n240 ) ;
 assign n3974 = ( n476  &  n499 ) | ( n3727  &  n499 ) | ( n476  &  n3729 ) | ( n3727  &  n3729 ) ;
 assign n3975 = ( n527  &  n552 ) | ( n3727  &  n552 ) | ( n527  &  n3729 ) | ( n3727  &  n3729 ) ;
 assign n3976 = ( n573 ) | ( (~ Ni37)  &  n202 ) ;
 assign n3977 = ( n568 ) | ( (~ Ni37)  &  n202 ) ;
 assign n3978 = ( n594 ) | ( (~ Ni37)  &  n240 ) ;
 assign n3979 = ( n589 ) | ( (~ Ni37)  &  n240 ) ;
 assign n3980 = ( n578  &  n599 ) | ( n3727  &  n599 ) | ( n578  &  n3729 ) | ( n3727  &  n3729 ) ;
 assign n3981 = ( n624  &  n648 ) | ( n3727  &  n648 ) | ( n624  &  n3729 ) | ( n3727  &  n3729 ) ;
 assign n3982 = ( n307  &  n383 ) | ( n307  &  (~ n1965) ) | ( n383  &  (~ n3618) ) | ( (~ n1965)  &  (~ n3618) ) ;
 assign n3984 = ( n374 ) | ( n998 ) ;
 assign n3983 = ( n3777  &  n3984 ) | ( (~ n3732)  &  n3968  &  n3984 ) ;
 assign n3985 = ( (~ n778)  &  n3778 ) | ( (~ n759)  &  (~ n778)  &  n3975 ) ;
 assign n3987 = ( Ni32 ) | ( n271 ) | ( n3719 ) ;
 assign n3988 = ( Ni32 ) | ( n364 ) | ( n3719 ) ;
 assign n3989 = ( n402  &  n411 ) | ( n3727  &  n411 ) | ( n402  &  n3729 ) | ( n3727  &  n3729 ) ;
 assign n3990 = ( n431  &  n438 ) | ( n3727  &  n438 ) | ( n431  &  n3729 ) | ( n3727  &  n3729 ) ;
 assign n3991 = ( n673  &  n683 ) | ( n3727  &  n683 ) | ( n673  &  n3729 ) | ( n3727  &  n3729 ) ;
 assign n3992 = ( n696  &  n704 ) | ( n3727  &  n704 ) | ( n696  &  n3729 ) | ( n3727  &  n3729 ) ;
 assign n3993 = ( n719  &  n729 ) | ( n3727  &  n729 ) | ( n719  &  n3729 ) | ( n3727  &  n3729 ) ;
 assign n3994 = ( n737  &  n744 ) | ( n3727  &  n744 ) | ( n737  &  n3729 ) | ( n3727  &  n3729 ) ;
 assign n3995 = ( n422  &  n449 ) | ( n422  &  (~ n1965) ) | ( n449  &  (~ n3618) ) | ( (~ n1965)  &  (~ n3618) ) ;
 assign n3997 = ( n441 ) | ( n998 ) ;
 assign n3996 = ( n3777  &  n3997 ) | ( (~ n3746)  &  n3989  &  n3997 ) ;
 assign n3998 = ( (~ n768)  &  n3778 ) | ( (~ n764)  &  (~ n768)  &  n3992 ) ;
 assign n4000 = ( n529  &  n554 ) | ( n3776  &  n554 ) | ( n529  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n4001 = ( n4000  &  n479 ) | ( n4000  &  n891 ) ;
 assign n4002 = ( Pi19  &  n310 ) | ( Pi19  &  n502 ) | ( n310  &  (~ n779) ) | ( n502  &  (~ n779) ) ;
 assign n4003 = ( n698  &  n706 ) | ( n3776  &  n706 ) | ( n698  &  n1692 ) | ( n3776  &  n1692 ) ;
 assign n4004 = ( n4003  &  n676 ) | ( n4003  &  n891 ) ;
 assign n4005 = ( Pi19  &  n310 ) | ( Pi19  &  n686 ) | ( n310  &  (~ n769) ) | ( n686  &  (~ n769) ) ;
 assign n4006 = ( n657  &  n753 ) | ( n3763  &  n753 ) | ( n657  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4008 = ( n309  &  n424 ) | ( n3742  &  n424 ) | ( n309  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4009 = ( n385  &  n451 ) | ( n3763  &  n451 ) | ( n385  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4010 = ( n232  &  n265 ) | ( n3728  &  n265 ) | ( n232  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4011 = ( n476  &  n499 ) | ( n3728  &  n499 ) | ( n476  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4012 = ( n527  &  n552 ) | ( n3728  &  n552 ) | ( n527  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4013 = ( n291  &  n307 ) | ( n307  &  n1474 ) | ( n291  &  (~ n2939) ) | ( n1474  &  (~ n2939) ) ;
 assign n4014 = ( Pi25 ) | ( n3713 ) ;
 assign n4015 = ( n402  &  n411 ) | ( n3728  &  n411 ) | ( n402  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4016 = ( n673  &  n683 ) | ( n3728  &  n683 ) | ( n673  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4017 = ( n696  &  n704 ) | ( n3728  &  n704 ) | ( n696  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4018 = ( n417  &  n422 ) | ( n422  &  n1474 ) | ( n417  &  (~ n2939) ) | ( n1474  &  (~ n2939) ) ;
 assign n4019 = ( n336  &  n360 ) | ( n3728  &  n360 ) | ( n336  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4020 = ( n578  &  n599 ) | ( n3728  &  n599 ) | ( n578  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4021 = ( n624  &  n648 ) | ( n3728  &  n648 ) | ( n624  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4022 = ( n378  &  n383 ) | ( n383  &  n1474 ) | ( n378  &  (~ n2939) ) | ( n1474  &  (~ n2939) ) ;
 assign n4023 = ( n431  &  n438 ) | ( n3728  &  n438 ) | ( n431  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4024 = ( n719  &  n729 ) | ( n3728  &  n729 ) | ( n719  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4025 = ( n737  &  n744 ) | ( n3728  &  n744 ) | ( n737  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4026 = ( n444  &  n449 ) | ( n449  &  n1474 ) | ( n444  &  (~ n2939) ) | ( n1474  &  (~ n2939) ) ;
 assign n4027 = ( n808  &  n831 ) | ( n3742  &  n831 ) | ( n808  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4028 = ( n795  &  n819 ) | ( n3763  &  n819 ) | ( n795  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4029 = ( n1503  &  n1248 ) | ( n3777  &  n1248 ) | ( n1503  &  n3579 ) | ( n3777  &  n3579 ) ;
 assign n4030 = ( n4029  &  n1538 ) | ( n4029  &  n1884 ) ;
 assign n4031 = ( n1535  &  n1256 ) | ( n3778  &  n1256 ) | ( n1535  &  n3582 ) | ( n3778  &  n3582 ) ;
 assign n4032 = ( n4031  &  n1257 ) | ( n4031  &  n3576 ) ;
 assign n4033 = ( n1252  &  n1254 ) | ( n3777  &  n1254 ) | ( n1252  &  n3579 ) | ( n3777  &  n3579 ) ;
 assign n4034 = ( n4033  &  n1259 ) | ( n4033  &  n1884 ) ;
 assign n4035 = ( n1260  &  n1262 ) | ( n3778  &  n1262 ) | ( n1260  &  n3582 ) | ( n3778  &  n3582 ) ;
 assign n4036 = ( n4035  &  n1263 ) | ( n4035  &  n3576 ) ;
 assign n4037 = ( n1308  &  n887 ) ;
 assign n4038 = ( n1318  &  n883 ) ;
 assign n4039 = ( n1378  &  n912 ) ;
 assign n4040 = ( n1388  &  n908 ) ;
 assign n4041 = ( n1272  &  n900 ) ;
 assign n4042 = ( n1283  &  n896 ) ;
 assign n4043 = ( n1343  &  n924 ) ;
 assign n4044 = ( n1353  &  n920 ) ;
 assign n4045 = ( n1231  &  n1239 ) | ( n3742  &  n1239 ) | ( n1231  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4046 = ( n1235  &  n1243 ) | ( n3763  &  n1243 ) | ( n1235  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4047 = ( n1334  &  n844 ) ;
 assign n4048 = ( n1404  &  n863 ) ;
 assign n4049 = ( n1299  &  n854 ) ;
 assign n4050 = ( n1369  &  n872 ) ;
 assign n4051 = ( n1219  &  n1225 ) | ( n3742  &  n1225 ) | ( n1219  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4053 = ( n1222  &  n1228 ) | ( n3763  &  n1228 ) | ( n1222  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4055 = ( n1031  &  n839 ) ;
 assign n4057 = ( n1049  &  n850 ) ;
 assign n4056 = ( n4057  &  n857 ) | ( n3728  &  n857 ) | ( n4057  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4059 = ( n1028  &  n883 ) ;
 assign n4058 = ( n890  &  n4059 ) | ( n3728  &  n4059 ) | ( n890  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4061 = ( n1019  &  n885 ) ;
 assign n4062 = ( n1022  &  n887 ) ;
 assign n4060 = ( n4061  &  n4062 ) | ( n3728  &  n4062 ) | ( n4061  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4064 = ( n1046  &  n896 ) ;
 assign n4063 = ( n903  &  n4064 ) | ( n3728  &  n4064 ) | ( n903  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4066 = ( n1037  &  n898 ) ;
 assign n4067 = ( n1040  &  n900 ) ;
 assign n4065 = ( n4066  &  n4067 ) | ( n3728  &  n4067 ) | ( n4066  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4068 = ( n1477  &  n1502 ) | ( n1474  &  n1502 ) | ( n1477  &  n3777 ) | ( n1474  &  n3777 ) ;
 assign n4069 = ( n972  &  n859 ) ;
 assign n4071 = ( n990  &  n868 ) ;
 assign n4070 = ( n4071  &  n875 ) | ( n3728  &  n875 ) | ( n4071  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4073 = ( n969  &  n908 ) ;
 assign n4072 = ( n915  &  n4073 ) | ( n3728  &  n4073 ) | ( n915  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4075 = ( n960  &  n910 ) ;
 assign n4076 = ( n963  &  n912 ) ;
 assign n4074 = ( n4075  &  n4076 ) | ( n3728  &  n4076 ) | ( n4075  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4078 = ( n987  &  n920 ) ;
 assign n4077 = ( n927  &  n4078 ) | ( n3728  &  n4078 ) | ( n927  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4080 = ( n978  &  n922 ) ;
 assign n4081 = ( n981  &  n924 ) ;
 assign n4079 = ( n4080  &  n4081 ) | ( n3728  &  n4081 ) | ( n4080  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4082 = ( n1473  &  n1479 ) | ( n1474  &  n1479 ) | ( n1473  &  n3777 ) | ( n1474  &  n3777 ) ;
 assign n4083 = ( n1538  &  n1535 ) | ( n1249  &  n1535 ) | ( n1538  &  n1250 ) | ( n1249  &  n1250 ) ;
 assign n4084 = ( n4083  &  n1258 ) | ( n4083  &  n3754 ) ;
 assign n4085 = ( n1255  &  n1261 ) | ( n3763  &  n1261 ) | ( n1255  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4086 = ( n1503  &  n845 ) | ( n1249  &  n845 ) | ( n1503  &  n1250 ) | ( n1249  &  n1250 ) ;
 assign n4087 = ( n4086  &  n1251 ) | ( n4086  &  n3754 ) ;
 assign n4088 = ( n1247  &  n1253 ) | ( n3763  &  n1253 ) | ( n1247  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4089 = ( n889  &  n914 ) | ( n3742  &  n914 ) | ( n889  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4090 = ( n902  &  n926 ) | ( n3763  &  n926 ) | ( n902  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4091 = ( n846  &  n865 ) | ( n3742  &  n865 ) | ( n846  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4093 = ( n856  &  n874 ) | ( n3763  &  n874 ) | ( n856  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4095 = ( n1333 ) | ( n3810 ) ;
 assign n4096 = ( n1602 ) | ( (~ n2939) ) ;
 assign n4097 = ( n1403 ) | ( n3810 ) ;
 assign n4098 = ( n1298 ) | ( n3810 ) ;
 assign n4099 = ( n1368 ) | ( n3810 ) ;
 assign n4100 = ( n1621  &  n1639 ) | ( n3742  &  n1639 ) | ( n1621  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4101 = ( n1612  &  n1630 ) | ( n3763  &  n1630 ) | ( n1612  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4102 = ( n845 ) | ( n3806 ) ;
 assign n4103 = ( n1563 ) | ( (~ n2939) ) ;
 assign n4104 = ( n864 ) | ( n3806 ) ;
 assign n4105 = ( n855 ) | ( n3806 ) ;
 assign n4106 = ( n873 ) | ( n3806 ) ;
 assign n4107 = ( n1581  &  n1599 ) | ( n3742  &  n1599 ) | ( n1581  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4108 = ( n1572  &  n1590 ) | ( n3763  &  n1590 ) | ( n1572  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4109 = ( n1333 ) | ( n3815 ) ;
 assign n4110 = ( n1523 ) | ( (~ n2939) ) ;
 assign n4111 = ( n1403 ) | ( n3815 ) ;
 assign n4112 = ( n1298 ) | ( n3815 ) ;
 assign n4113 = ( n1368 ) | ( n3815 ) ;
 assign n4114 = ( n1542  &  n1560 ) | ( n3742  &  n1560 ) | ( n1542  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4115 = ( n1531  &  n1551 ) | ( n3763  &  n1551 ) | ( n1531  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4117 = ( n4676 ) | ( n4677 ) | ( n3814 ) ;
 assign n4116 = ( n4117  &  n3499 ) | ( n4117  &  n4115  &  n4114 ) ;
 assign n4120 = ( n940  &  (~ n3784) ) ;
 assign n4119 = ( n4120  &  Ni11 ) | ( n1522  &  Ni11 ) | ( n4120  &  n1520 ) | ( n1522  &  n1520 ) ;
 assign n4122 = ( n1332 ) | ( n3785 ) ;
 assign n4123 = ( n942 ) | ( (~ n2939) ) ;
 assign n4124 = ( n1402 ) | ( n3785 ) ;
 assign n4125 = ( n1297 ) | ( n3785 ) ;
 assign n4126 = ( n1367 ) | ( n3785 ) ;
 assign n4127 = ( n1329  &  n1220 ) | ( n3794  &  n1220 ) | ( n1329  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4128 = ( n1322  &  n1325 ) | ( n3796  &  n1325 ) | ( n1322  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4129 = ( n1294  &  n1223 ) | ( n3794  &  n1223 ) | ( n1294  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4130 = ( n1287  &  n1290 ) | ( n3796  &  n1290 ) | ( n1287  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4131 = ( n1232  &  n4038 ) | ( n3794  &  n4038 ) | ( n1232  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4132 = ( n1313  &  n1316 ) | ( n3796  &  n1316 ) | ( n1313  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4133 = ( n1310  &  n4037 ) | ( n3794  &  n4037 ) | ( n1310  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4134 = ( n1303  &  n1306 ) | ( n3796  &  n1306 ) | ( n1303  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4135 = ( n1236  &  n4042 ) | ( n3794  &  n4042 ) | ( n1236  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4136 = ( n1278  &  n1281 ) | ( n3796  &  n1281 ) | ( n1278  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4137 = ( n1274  &  n4041 ) | ( n3794  &  n4041 ) | ( n1274  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4138 = ( n1267  &  n1270 ) | ( n3796  &  n1270 ) | ( n1267  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4139 = ( n4047  &  n4049 ) | ( n3790  &  n4049 ) | ( n4047  &  n3791 ) | ( n3790  &  n3791 ) ;
 assign n4141 = ( n1297 ) | ( n3793 ) ;
 assign n4140 = ( n4141  &  n3777 ) | ( n4141  &  n4128  &  n4127 ) ;
 assign n4142 = ( n4140  &  n3579 ) | ( n4140  &  n4130  &  n4129 ) ;
 assign n4143 = ( (~ n1411)  &  n3778 ) | ( (~ n1411)  &  n4133  &  n4134 ) ;
 assign n4145 = ( n4143  &  n3582 ) | ( n4143  &  n4136  &  n4135 ) ;
 assign n4146 = ( n1087  &  n3576 ) | ( n1087  &  n4138  &  n4137 ) ;
 assign n4147 = ( n1399  &  n1226 ) | ( n3794  &  n1226 ) | ( n1399  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4148 = ( n1392  &  n1395 ) | ( n3796  &  n1395 ) | ( n1392  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4149 = ( n1364  &  n1229 ) | ( n3794  &  n1229 ) | ( n1364  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4150 = ( n1357  &  n1360 ) | ( n3796  &  n1360 ) | ( n1357  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4151 = ( n1240  &  n4040 ) | ( n3794  &  n4040 ) | ( n1240  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4152 = ( n1383  &  n1386 ) | ( n3796  &  n1386 ) | ( n1383  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4153 = ( n1380  &  n4039 ) | ( n3794  &  n4039 ) | ( n1380  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4154 = ( n1373  &  n1376 ) | ( n3796  &  n1376 ) | ( n1373  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4155 = ( n1244  &  n4044 ) | ( n3794  &  n4044 ) | ( n1244  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4156 = ( n1348  &  n1351 ) | ( n3796  &  n1351 ) | ( n1348  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4157 = ( n1345  &  n4043 ) | ( n3794  &  n4043 ) | ( n1345  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4158 = ( n1338  &  n1341 ) | ( n3796  &  n1341 ) | ( n1338  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4159 = ( n4048  &  n4050 ) | ( n3790  &  n4050 ) | ( n4048  &  n3791 ) | ( n3790  &  n3791 ) ;
 assign n4161 = ( n1367 ) | ( n3793 ) ;
 assign n4160 = ( n4161  &  n3777 ) | ( n4161  &  n4148  &  n4147 ) ;
 assign n4162 = ( n4160  &  n3579 ) | ( n4160  &  n4150  &  n4149 ) ;
 assign n4163 = ( (~ n1408)  &  n3778 ) | ( (~ n1408)  &  n4153  &  n4154 ) ;
 assign n4165 = ( n4163  &  n3582 ) | ( n4163  &  n4156  &  n4155 ) ;
 assign n4166 = ( n1087  &  n3576 ) | ( n1087  &  n4158  &  n4157 ) ;
 assign n4167 = ( n1332 ) | ( n3799 ) ;
 assign n4168 = ( (~ n2939) ) | ( (~ n3804) ) ;
 assign n4169 = ( n1402 ) | ( n3799 ) ;
 assign n4170 = ( n1297 ) | ( n3799 ) ;
 assign n4171 = ( n1367 ) | ( n3799 ) ;
 assign n4172 = ( n1335  &  n1405 ) | ( n3742  &  n1405 ) | ( n1335  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4173 = ( n1300  &  n1370 ) | ( n3763  &  n1370 ) | ( n1300  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4174 = ( n1265  &  n1466 ) | ( n1265  &  n3499 ) | ( n1466  &  (~ n3784) ) | ( n3499  &  (~ n3784) ) ;
 assign n4177 = ( Ni14  &  n1087 ) | ( (~ Ni14)  &  n4233 ) | ( n1087  &  n4233 ) ;
 assign n4176 = ( (~ Pi23)  &  n3655 ) | ( n3655  &  n4177 ) ;
 assign n4178 = ( n1011 ) | ( n3820 ) ;
 assign n4179 = ( (~ n164) ) | ( (~ n2939) ) ;
 assign n4180 = ( n951 ) | ( n3820 ) ;
 assign n4181 = ( n1014 ) | ( n3820 ) ;
 assign n4182 = ( n955 ) | ( n3820 ) ;
 assign n4183 = ( n1113  &  n1137 ) | ( n3742  &  n1137 ) | ( n1113  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4184 = ( n1101  &  n1125 ) | ( n3763  &  n1125 ) | ( n1101  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4186 = ( n1062  &  Pi24 ) | ( n1866  &  Pi24 ) | ( n1062  &  n3649 ) | ( n1866  &  n3649 ) ;
 assign n4187 = ( n4055  &  n847 ) | ( n3827  &  n847 ) | ( n4055  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4188 = ( n1029  &  n1032 ) | ( n3829  &  n1032 ) | ( n1029  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4189 = ( n4057  &  n857 ) | ( n3827  &  n857 ) | ( n4057  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4190 = ( n1047  &  n1050 ) | ( n3829  &  n1050 ) | ( n1047  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4191 = ( n890  &  n4059 ) | ( n3827  &  n4059 ) | ( n890  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4192 = ( n1023  &  n1026 ) | ( n3829  &  n1026 ) | ( n1023  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4193 = ( n4061  &  n4062 ) | ( n3827  &  n4062 ) | ( n4061  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4194 = ( n1017  &  n1020 ) | ( n3829  &  n1020 ) | ( n1017  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4195 = ( n903  &  n4064 ) | ( n3827  &  n4064 ) | ( n903  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4196 = ( n1041  &  n1044 ) | ( n3829  &  n1044 ) | ( n1041  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4197 = ( n4066  &  n4067 ) | ( n3827  &  n4067 ) | ( n4066  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4198 = ( n1035  &  n1038 ) | ( n3829  &  n1038 ) | ( n1035  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4199 = ( n1011  &  n1014 ) | ( n3825  &  n1014 ) | ( n1011  &  n3826 ) | ( n3825  &  n3826 ) ;
 assign n4200 = ( (~ n1056)  &  n3579 ) | ( (~ n1056)  &  n4189  &  n4190 ) ;
 assign n4202 = ( n4199  &  n4200  &  Pi24 ) | ( n4199  &  n4200  &  n1053 ) ;
 assign n4203 = ( (~ n1059)  &  n3778 ) | ( (~ n1059)  &  n4193  &  n4194 ) ;
 assign n4205 = ( n4203  &  n3582 ) | ( n4203  &  n4196  &  n4195 ) ;
 assign n4206 = ( n950  &  n3576 ) | ( n950  &  n4198  &  n4197 ) ;
 assign n4207 = ( n4069  &  n866 ) | ( n3827  &  n866 ) | ( n4069  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4208 = ( n970  &  n973 ) | ( n3829  &  n973 ) | ( n970  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4209 = ( n4071  &  n875 ) | ( n3827  &  n875 ) | ( n4071  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4210 = ( n988  &  n991 ) | ( n3829  &  n991 ) | ( n988  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4211 = ( n915  &  n4073 ) | ( n3827  &  n4073 ) | ( n915  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4212 = ( n964  &  n967 ) | ( n3829  &  n967 ) | ( n964  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4213 = ( n4075  &  n4076 ) | ( n3827  &  n4076 ) | ( n4075  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4214 = ( n958  &  n961 ) | ( n3829  &  n961 ) | ( n958  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4215 = ( n927  &  n4078 ) | ( n3827  &  n4078 ) | ( n927  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4216 = ( n982  &  n985 ) | ( n3829  &  n985 ) | ( n982  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4217 = ( n4080  &  n4081 ) | ( n3827  &  n4081 ) | ( n4080  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4218 = ( n976  &  n979 ) | ( n3829  &  n979 ) | ( n976  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4219 = ( n951  &  n955 ) | ( n3825  &  n955 ) | ( n951  &  n3826 ) | ( n3825  &  n3826 ) ;
 assign n4221 = ( (~ n1003)  &  n3778 ) | ( (~ n1003)  &  n4213  &  n4214 ) ;
 assign n4223 = ( n1006  &  n947 ) | ( n1993  &  n947 ) | ( n1006  &  n1067 ) | ( n1993  &  n1067 ) ;
 assign n4224 = ( n3655  &  Pi23 ) | ( n3655  &  n4177 ) ;
 assign n4225 = ( n1011 ) | ( n3832 ) ;
 assign n4226 = ( (~ n167) ) | ( (~ n2939) ) ;
 assign n4227 = ( n951 ) | ( n3832 ) ;
 assign n4228 = ( n1014 ) | ( n3832 ) ;
 assign n4229 = ( n955 ) | ( n3832 ) ;
 assign n4230 = ( n1178  &  n1202 ) | ( n3742  &  n1202 ) | ( n1178  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4231 = ( n1166  &  n1190 ) | ( n3763  &  n1190 ) | ( n1166  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4233 = ( n1603 ) | ( n1866 ) ;
 assign n4236 = ( n2009  &  (~ n2013) ) | ( (~ n2013)  &  n3777 ) ;
 assign n4238 = ( n2012  &  n2008 ) | ( n3579  &  n2008 ) | ( n2012  &  n1884 ) | ( n3579  &  n1884 ) ;
 assign n4239 = ( n2007  &  n2011 ) | ( n3778  &  n2011 ) | ( n2007  &  n3582 ) | ( n3778  &  n3582 ) ;
 assign n4240 = ( n2002  &  n1998 ) | ( n3579  &  n1998 ) | ( n2002  &  n1884 ) | ( n3579  &  n1884 ) ;
 assign n4241 = ( n1999  &  (~ n2003)  &  n4240 ) | ( (~ n2003)  &  n3777  &  n4240 ) ;
 assign n4244 = ( n1996  &  n2001 ) | ( n3778  &  n2001 ) | ( n1996  &  n3582 ) | ( n3778  &  n3582 ) ;
 assign n4245 = ( n1995  &  n4244  &  n2000 ) | ( n1995  &  n4244  &  n3576 ) ;
 assign n4247 = ( (~ n507)  &  n1795 ) | ( (~ n507)  &  n3836 ) | ( n1795  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n4248 = ( (~ Pi25)  &  n1689 ) | ( n1689  &  n1926 ) ;
 assign n4249 = ( (~ n687)  &  n1835 ) | ( (~ n687)  &  n3836 ) | ( n1835  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n4250 = ( (~ Pi25)  &  n1704 ) | ( n1704  &  n1890 ) ;
 assign n4251 = ( (~ n607)  &  n1815 ) | ( (~ n607)  &  n3836 ) | ( n1815  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n4252 = ( (~ Pi25)  &  n1697 ) | ( n1697  &  n1933 ) ;
 assign n4253 = ( (~ n733)  &  n1855 ) | ( (~ n733)  &  n3836 ) | ( n1855  &  n3838 ) | ( n3836  &  n3838 ) ;
 assign n4254 = ( (~ Pi25)  &  n1711 ) | ( n1711  &  n1897 ) ;
 assign n4255 = ( n1802  &  n1842 ) | ( n3742  &  n1842 ) | ( n1802  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4256 = ( n1822  &  n1862 ) | ( n3763  &  n1862 ) | ( n1822  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4257 = ( n1732  &  n1766 ) | ( n3742  &  n1766 ) | ( n1732  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4258 = ( n1749  &  n1783 ) | ( n3763  &  n1783 ) | ( n1749  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4259 = ( n1966  &  n1727 ) | ( n3713  &  n1727 ) | ( n1966  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4260 = ( n1967  &  n1744 ) | ( n3713  &  n1744 ) | ( n1967  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4261 = ( n1980  &  n1716 ) | ( n3713  &  n1716 ) | ( n1980  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4262 = ( n1983  &  n1734 ) | ( n3713  &  n1734 ) | ( n1983  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4263 = ( n1978  &  n1785 ) | ( n3713  &  n1785 ) | ( n1978  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4264 = ( n1979  &  n1795 ) | ( n3713  &  n1795 ) | ( n1979  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4265 = ( n1981  &  n1805 ) | ( n3713  &  n1805 ) | ( n1981  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4266 = ( n1982  &  n1815 ) | ( n3713  &  n1815 ) | ( n1982  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4267 = ( (~ n1984)  &  n3579 ) | ( (~ n1984)  &  n3841  &  n4262 ) ;
 assign n4269 = ( n4267  &  n1884 ) | ( n4267  &  n4263  &  n3841 ) ;
 assign n4270 = ( (~ n1986)  &  n3778 ) | ( (~ n1986)  &  n3841  &  n4264 ) ;
 assign n4272 = ( n4270  &  n3576 ) | ( n4270  &  n4266  &  n3841 ) ;
 assign n4273 = ( n1970  &  n1722 ) | ( n3713  &  n1722 ) | ( n1970  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4274 = ( n1973  &  n1739 ) | ( n3713  &  n1739 ) | ( n1973  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4275 = ( n1968  &  n1790 ) | ( n3713  &  n1790 ) | ( n1968  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4276 = ( n1969  &  n1797 ) | ( n3713  &  n1797 ) | ( n1969  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4277 = ( n1971  &  n1810 ) | ( n3713  &  n1810 ) | ( n1971  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4278 = ( n1972  &  n1817 ) | ( n3713  &  n1817 ) | ( n1972  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4279 = ( (~ n1974)  &  n3579 ) | ( (~ n1974)  &  n3841  &  n4274 ) ;
 assign n4281 = ( n4279  &  n1884 ) | ( n4279  &  n4275  &  n3841 ) ;
 assign n4283 = ( (~ n1976)  &  n3778 ) | ( (~ n1976)  &  n3841  &  n4276 ) ;
 assign n4285 = ( n4283  &  n3576 ) | ( n4283  &  n4278  &  n3841 ) ;
 assign n4287 = ( (~ n1988)  &  (~ n3618) ) | ( (~ n1988)  &  n3841  &  n4259 ) ;
 assign n4289 = ( n1940  &  n1761 ) | ( n3713  &  n1761 ) | ( n1940  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4290 = ( n1941  &  n1778 ) | ( n3713  &  n1778 ) | ( n1941  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4291 = ( n1955  &  n1751 ) | ( n3713  &  n1751 ) | ( n1955  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4292 = ( n1958  &  n1768 ) | ( n3713  &  n1768 ) | ( n1958  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4293 = ( n1953  &  n1825 ) | ( n3713  &  n1825 ) | ( n1953  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4294 = ( n1954  &  n1835 ) | ( n3713  &  n1835 ) | ( n1954  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4295 = ( n1956  &  n1845 ) | ( n3713  &  n1845 ) | ( n1956  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4296 = ( n1957  &  n1855 ) | ( n3713  &  n1855 ) | ( n1957  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4297 = ( (~ n1959)  &  n3579 ) | ( (~ n1959)  &  n3841  &  n4292 ) ;
 assign n4299 = ( n4297  &  n1884 ) | ( n4297  &  n4293  &  n3841 ) ;
 assign n4300 = ( (~ n1961)  &  n3778 ) | ( (~ n1961)  &  n3841  &  n4294 ) ;
 assign n4302 = ( n4300  &  n3576 ) | ( n4300  &  n4296  &  n3841 ) ;
 assign n4303 = ( n1944  &  n1756 ) | ( n3713  &  n1756 ) | ( n1944  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4304 = ( n1947  &  n1773 ) | ( n3713  &  n1773 ) | ( n1947  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4305 = ( n1942  &  n1830 ) | ( n3713  &  n1830 ) | ( n1942  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4306 = ( n1943  &  n1837 ) | ( n3713  &  n1837 ) | ( n1943  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4307 = ( n1945  &  n1850 ) | ( n3713  &  n1850 ) | ( n1945  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4308 = ( n1946  &  n1857 ) | ( n3713  &  n1857 ) | ( n1946  &  n3839 ) | ( n3713  &  n3839 ) ;
 assign n4309 = ( (~ n1948)  &  n3579 ) | ( (~ n1948)  &  n3841  &  n4304 ) ;
 assign n4311 = ( n4309  &  n1884 ) | ( n4309  &  n4305  &  n3841 ) ;
 assign n4313 = ( (~ n1951)  &  n3778 ) | ( (~ n1951)  &  n3841  &  n4306 ) ;
 assign n4315 = ( n4313  &  n3576 ) | ( n4313  &  n4308  &  n3841 ) ;
 assign n4317 = ( (~ n1963)  &  (~ n3618) ) | ( (~ n1963)  &  n3841  &  n4289 ) ;
 assign n4319 = ( n1925  &  n1930 ) | ( n3778  &  n1930 ) | ( n1925  &  n3582 ) | ( n3778  &  n3582 ) ;
 assign n4320 = ( n1910  &  n1914 ) | ( n3778  &  n1914 ) | ( n1910  &  n3582 ) | ( n3778  &  n3582 ) ;
 assign n4321 = ( n1904  &  n1906 ) | ( n1904  &  (~ n1965) ) | ( n1906  &  (~ n3618) ) | ( (~ n1965)  &  (~ n3618) ) ;
 assign n4322 = ( n1889  &  n1894 ) | ( n3778  &  n1894 ) | ( n1889  &  n3582 ) | ( n3778  &  n3582 ) ;
 assign n4323 = ( n1873  &  n1877 ) | ( n3778  &  n1877 ) | ( n1873  &  n3582 ) | ( n3778  &  n3582 ) ;
 assign n4325 = ( (~ n3113) ) | ( n4711 ) | ( n4712 ) ;
 assign n4324 = ( Pi20  &  n1920 ) | ( (~ Pi20)  &  n1937 ) | ( n1920  &  n1937 ) ;
 assign n4326 = ( n1691  &  n1706 ) | ( n3742  &  n1706 ) | ( n1691  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4328 = ( n1699  &  n1713 ) | ( n3763  &  n1713 ) | ( n1699  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4330 = ( n1669  &  n1680 ) | ( n3742  &  n1680 ) | ( n1669  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4331 = ( n1675  &  n1685 ) | ( n3763  &  n1685 ) | ( n1675  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4332 = ( (~ Pi23)  &  n691 ) | ( n691  &  n3662 ) | ( (~ Pi23)  &  n3845 ) | ( n3662  &  n3845 ) ;
 assign n4333 = ( (~ Pi24)  &  n275 ) | ( n275  &  n3662 ) | ( (~ Pi24)  &  n3845 ) | ( n3662  &  n3845 ) ;
 assign n4334 = ( Pi15  &  n2057 ) | ( n2057  &  n2062 ) | ( Pi15  &  (~ n3712) ) | ( n2062  &  (~ n3712) ) ;
 assign n4337 = ( n2564  &  n2566 ) | ( n3777  &  n2566 ) | ( n2564  &  n3579 ) | ( n3777  &  n3579 ) ;
 assign n4338 = ( n4337  &  n2570 ) | ( n4337  &  n1884 ) ;
 assign n4339 = ( n2571  &  n2573 ) | ( n3778  &  n2573 ) | ( n2571  &  n3582 ) | ( n3778  &  n3582 ) ;
 assign n4340 = ( n4339  &  n2574 ) | ( n4339  &  n3576 ) ;
 assign n4341 = ( n2762  &  n2568 ) | ( n3777  &  n2568 ) | ( n2762  &  n3579 ) | ( n3777  &  n3579 ) ;
 assign n4342 = ( n4341  &  n2832 ) | ( n4341  &  n1884 ) ;
 assign n4343 = ( n2829  &  n2576 ) | ( n3778  &  n2576 ) | ( n2829  &  n3582 ) | ( n3778  &  n3582 ) ;
 assign n4344 = ( n4343  &  n2577 ) | ( n4343  &  n3576 ) ;
 assign n4345 = ( n2534  &  n2211 ) ;
 assign n4346 = ( n2532  &  n2194 ) ;
 assign n4347 = ( n2550  &  n2268 ) ;
 assign n4348 = ( n2548  &  n2255 ) ;
 assign n4349 = ( n2542  &  n2241 ) ;
 assign n4350 = ( n2540  &  n2225 ) ;
 assign n4351 = ( n2558  &  n2294 ) ;
 assign n4352 = ( n2556  &  n2282 ) ;
 assign n4353 = ( n2535  &  n2551 ) | ( n3742  &  n2551 ) | ( n2535  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4354 = ( n2543  &  n2559 ) | ( n3763  &  n2559 ) | ( n2543  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4355 = ( n2509  &  n2112 ) ;
 assign n4356 = ( n2521  &  n2159 ) ;
 assign n4357 = ( n2515  &  n2138 ) ;
 assign n4358 = ( n2527  &  n2179 ) ;
 assign n4359 = ( n2510  &  n2522 ) | ( n3742  &  n2522 ) | ( n2510  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4361 = ( n2516  &  n2528 ) | ( n3763  &  n2528 ) | ( n2516  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4363 = ( n2088  &  n2092 ) ;
 assign n4365 = ( n2120  &  n2123 ) ;
 assign n4364 = ( n4365  &  n2141 ) | ( n3728  &  n2141 ) | ( n4365  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4366 = ( n2214  &  n2425 ) | ( n3728  &  n2425 ) | ( n2214  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4368 = ( n2200  &  n2203 ) ;
 assign n4367 = ( n4368  &  n2422 ) | ( n3728  &  n2422 ) | ( n4368  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4369 = ( n2244  &  n2414 ) | ( n3728  &  n2414 ) | ( n2244  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4371 = ( n2230  &  n2233 ) ;
 assign n4370 = ( n4371  &  n2410 ) | ( n3728  &  n2410 ) | ( n4371  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4372 = ( n2759  &  n2780 ) | ( n1474  &  n2780 ) | ( n2759  &  n3777 ) | ( n1474  &  n3777 ) ;
 assign n4373 = ( n2145  &  n2148 ) ;
 assign n4375 = ( n2165  &  n2168 ) ;
 assign n4374 = ( n4375  &  n2182 ) | ( n3728  &  n2182 ) | ( n4375  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4376 = ( n2271  &  n2447 ) | ( n3728  &  n2447 ) | ( n2271  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4378 = ( n2259  &  n2262 ) ;
 assign n4377 = ( n4378  &  n2444 ) | ( n3728  &  n2444 ) | ( n4378  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4379 = ( n2297  &  n2436 ) | ( n3728  &  n2436 ) | ( n2297  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4381 = ( n2285  &  n2288 ) ;
 assign n4380 = ( n4381  &  n2433 ) | ( n3728  &  n2433 ) | ( n4381  &  n3731 ) | ( n3728  &  n3731 ) ;
 assign n4382 = ( n2756  &  n2761 ) | ( n1474  &  n2761 ) | ( n2756  &  n3777 ) | ( n1474  &  n3777 ) ;
 assign n4383 = ( n2832  &  n2829 ) | ( n1249  &  n2829 ) | ( n2832  &  n1250 ) | ( n1249  &  n1250 ) ;
 assign n4384 = ( n4383  &  n2569 ) | ( n4383  &  n3742 ) ;
 assign n4385 = ( n2572  &  n2575 ) | ( n3763  &  n2575 ) | ( n2572  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4386 = ( n2762  &  n2160 ) | ( n1249  &  n2160 ) | ( n2762  &  n1250 ) | ( n1249  &  n1250 ) ;
 assign n4387 = ( n4386  &  n2563 ) | ( n4386  &  n3742 ) ;
 assign n4388 = ( n2565  &  n2567 ) | ( n3763  &  n2567 ) | ( n2565  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4389 = ( (~ n1068)  &  n2797 ) | ( (~ n1068)  &  n3783 ) | ( n2797  &  (~ n3898) ) | ( n3783  &  (~ n3898) ) ;
 assign n4391 = ( (~ n1654)  &  (~ n4389) ) | ( (~ n1650)  &  (~ n1654)  &  (~ n2578) ) ;
 assign n4394 = ( n2213  &  n2270 ) | ( n3742  &  n2270 ) | ( n2213  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4395 = ( n2243  &  n2296 ) | ( n3763  &  n2296 ) | ( n2243  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4396 = ( n2114  &  n2161 ) | ( n3742  &  n2161 ) | ( n2114  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4398 = ( n2140  &  n2181 ) | ( n3763  &  n2181 ) | ( n2140  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4400 = ( n2633 ) | ( n3810 ) ;
 assign n4401 = ( n2876 ) | ( (~ n2939) ) ;
 assign n4402 = ( n2689 ) | ( n3810 ) ;
 assign n4403 = ( n2605 ) | ( n3810 ) ;
 assign n4404 = ( n2661 ) | ( n3810 ) ;
 assign n4405 = ( n2892  &  n2910 ) | ( n3742  &  n2910 ) | ( n2892  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4406 = ( n2883  &  n2901 ) | ( n3763  &  n2901 ) | ( n2883  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4407 = ( n2113 ) | ( n3806 ) ;
 assign n4408 = ( n2839 ) | ( (~ n2939) ) ;
 assign n4409 = ( n2160 ) | ( n3806 ) ;
 assign n4410 = ( n2139 ) | ( n3806 ) ;
 assign n4411 = ( n2180 ) | ( n3806 ) ;
 assign n4412 = ( n2855  &  n2873 ) | ( n3742  &  n2873 ) | ( n2855  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4414 = ( n2846  &  n2864 ) | ( n3763  &  n2864 ) | ( n2846  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4416 = ( n2633 ) | ( n3815 ) ;
 assign n4417 = ( n2800 ) | ( (~ n2939) ) ;
 assign n4418 = ( n2689 ) | ( n3815 ) ;
 assign n4419 = ( n2605 ) | ( n3815 ) ;
 assign n4420 = ( n2661 ) | ( n3815 ) ;
 assign n4421 = ( n2816  &  n2836 ) | ( n3742  &  n2836 ) | ( n2816  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4422 = ( n2807  &  n2825 ) | ( n3763  &  n2825 ) | ( n2807  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4423 = ( n2632 ) | ( n3785 ) ;
 assign n4424 = ( n2316 ) | ( (~ n2939) ) ;
 assign n4425 = ( n2688 ) | ( n3785 ) ;
 assign n4426 = ( n2604 ) | ( n3785 ) ;
 assign n4427 = ( n2660 ) | ( n3785 ) ;
 assign n4428 = ( n2629  &  n2511 ) | ( n3794  &  n2511 ) | ( n2629  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4429 = ( n2624  &  n2626 ) | ( n3796  &  n2626 ) | ( n2624  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4430 = ( n2601  &  n2517 ) | ( n3794  &  n2517 ) | ( n2601  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4431 = ( n2596  &  n2598 ) | ( n3796  &  n2598 ) | ( n2596  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4432 = ( n2536  &  n4346 ) | ( n3794  &  n4346 ) | ( n2536  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4433 = ( n2617  &  n2619 ) | ( n3796  &  n2619 ) | ( n2617  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4434 = ( n2614  &  n4345 ) | ( n3794  &  n4345 ) | ( n2614  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4435 = ( n2609  &  n2611 ) | ( n3796  &  n2611 ) | ( n2609  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4436 = ( n2544  &  n4350 ) | ( n3794  &  n4350 ) | ( n2544  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4437 = ( n2589  &  n2591 ) | ( n3796  &  n2591 ) | ( n2589  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4438 = ( n2586  &  n4349 ) | ( n3794  &  n4349 ) | ( n2586  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4439 = ( n2581  &  n2583 ) | ( n3796  &  n2583 ) | ( n2581  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4440 = ( n4355  &  n4357 ) | ( n3790  &  n4357 ) | ( n4355  &  n3791 ) | ( n3790  &  n3791 ) ;
 assign n4442 = ( n2604 ) | ( n3793 ) ;
 assign n4441 = ( n4442  &  n3777 ) | ( n4442  &  n4429  &  n4428 ) ;
 assign n4443 = ( n4441  &  n3579 ) | ( n4441  &  n4431  &  n4430 ) ;
 assign n4444 = ( (~ n2696)  &  n3778 ) | ( (~ n2696)  &  n4434  &  n4435 ) ;
 assign n4446 = ( n4444  &  n3582 ) | ( n4444  &  n4437  &  n4436 ) ;
 assign n4447 = ( n2310  &  n3576 ) | ( n2310  &  n4439  &  n4438 ) ;
 assign n4448 = ( n2685  &  n2523 ) | ( n3794  &  n2523 ) | ( n2685  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4449 = ( n2680  &  n2682 ) | ( n3796  &  n2682 ) | ( n2680  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4450 = ( n2657  &  n2529 ) | ( n3794  &  n2529 ) | ( n2657  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4451 = ( n2652  &  n2654 ) | ( n3796  &  n2654 ) | ( n2652  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4452 = ( n2552  &  n4348 ) | ( n3794  &  n4348 ) | ( n2552  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4453 = ( n2673  &  n2675 ) | ( n3796  &  n2675 ) | ( n2673  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4454 = ( n2670  &  n4347 ) | ( n3794  &  n4347 ) | ( n2670  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4455 = ( n2665  &  n2667 ) | ( n3796  &  n2667 ) | ( n2665  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4456 = ( n2560  &  n4352 ) | ( n3794  &  n4352 ) | ( n2560  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4457 = ( n2645  &  n2647 ) | ( n3796  &  n2647 ) | ( n2645  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4458 = ( n2642  &  n4351 ) | ( n3794  &  n4351 ) | ( n2642  &  n3795 ) | ( n3794  &  n3795 ) ;
 assign n4459 = ( n2637  &  n2639 ) | ( n3796  &  n2639 ) | ( n2637  &  n3797 ) | ( n3796  &  n3797 ) ;
 assign n4460 = ( n4356  &  n4358 ) | ( n3790  &  n4358 ) | ( n4356  &  n3791 ) | ( n3790  &  n3791 ) ;
 assign n4462 = ( n2660 ) | ( n3793 ) ;
 assign n4461 = ( n4462  &  n3777 ) | ( n4462  &  n4449  &  n4448 ) ;
 assign n4463 = ( n4461  &  n3579 ) | ( n4461  &  n4451  &  n4450 ) ;
 assign n4464 = ( (~ n2693)  &  n3778 ) | ( (~ n2693)  &  n4454  &  n4455 ) ;
 assign n4466 = ( n4464  &  n3582 ) | ( n4464  &  n4457  &  n4456 ) ;
 assign n4467 = ( n2310  &  n3576 ) | ( n2310  &  n4459  &  n4458 ) ;
 assign n4468 = ( n2632 ) | ( n3799 ) ;
 assign n4469 = ( n2306 ) | ( (~ n2939) ) ;
 assign n4470 = ( n2688 ) | ( n3799 ) ;
 assign n4471 = ( n2604 ) | ( n3799 ) ;
 assign n4472 = ( n2660 ) | ( n3799 ) ;
 assign n4473 = ( n2634  &  n2690 ) | ( n3742  &  n2690 ) | ( n2634  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4474 = ( n2606  &  n2662 ) | ( n3763  &  n2662 ) | ( n2606  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4475 = ( n2579  &  n2750 ) | ( n2579  &  n3499 ) | ( n2750  &  (~ n3784) ) | ( n3499  &  (~ n3784) ) ;
 assign n4476 = ( n3679  &  n194 ) | ( n3679  &  n3857 ) ;
 assign n4477 = ( n2330  &  n3681 ) | ( n2330  &  n3857 ) ;
 assign n4478 = ( n2332  &  n3678 ) | ( n2332  &  n3857 ) ;
 assign n4479 = ( n2456  &  n3798 ) | ( n2456  &  (~ n3910) ) | ( n3798  &  (~ n3912) ) | ( (~ n3910)  &  (~ n3912) ) ;
 assign n4480 = ( n2369  &  n2370 ) | ( n3822  &  n2370 ) | ( n2369  &  n1092 ) | ( n3822  &  n1092 ) ;
 assign n4481 = ( n2367  &  n2368 ) | ( n3822  &  n2368 ) | ( n2367  &  n1092 ) | ( n3822  &  n1092 ) ;
 assign n4482 = ( n2365  &  n2366 ) | ( n3822  &  n2366 ) | ( n2365  &  n1092 ) | ( n3822  &  n1092 ) ;
 assign n4484 = ( n2394 ) | ( (~ n2939) ) ;
 assign n4483 = ( n4484  &  n2363 ) | ( n4484  &  n3820 ) ;
 assign n4485 = ( n2342  &  n2343 ) | ( n3822  &  n2343 ) | ( n2342  &  n1092 ) | ( n3822  &  n1092 ) ;
 assign n4486 = ( n2340  &  n2341 ) | ( n3822  &  n2341 ) | ( n2340  &  n1092 ) | ( n3822  &  n1092 ) ;
 assign n4487 = ( n2338  &  n2339 ) | ( n3822  &  n2339 ) | ( n2338  &  n1092 ) | ( n3822  &  n1092 ) ;
 assign n4488 = ( n4484  &  n2336 ) | ( n4484  &  n3820 ) ;
 assign n4489 = ( n2375  &  n2376 ) | ( n3822  &  n2376 ) | ( n2375  &  n1092 ) | ( n3822  &  n1092 ) ;
 assign n4490 = ( n2373  &  n2374 ) | ( n3822  &  n2374 ) | ( n2373  &  n1092 ) | ( n3822  &  n1092 ) ;
 assign n4491 = ( n2371  &  n2372 ) | ( n3822  &  n2372 ) | ( n2371  &  n1092 ) | ( n3822  &  n1092 ) ;
 assign n4492 = ( n4484  &  n2364 ) | ( n4484  &  n3820 ) ;
 assign n4493 = ( n2348  &  n2349 ) | ( n3822  &  n2349 ) | ( n2348  &  n1092 ) | ( n3822  &  n1092 ) ;
 assign n4494 = ( n2346  &  n2347 ) | ( n3822  &  n2347 ) | ( n2346  &  n1092 ) | ( n3822  &  n1092 ) ;
 assign n4495 = ( n2344  &  n2345 ) | ( n3822  &  n2345 ) | ( n2344  &  n1092 ) | ( n3822  &  n1092 ) ;
 assign n4496 = ( n2337 ) | ( n3820 ) ;
 assign n4497 = ( n2429  &  n2451 ) | ( n3742  &  n2451 ) | ( n2429  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4498 = ( n2418  &  n2440 ) | ( n3763  &  n2440 ) | ( n2418  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4500 = ( n2396 ) | ( n2407 ) ;
 assign n4499 = ( n4500  &  n3113 ) | ( n4500  &  n4498  &  n4497 ) ;
 assign n4501 = ( n4363  &  n2115 ) | ( n3827  &  n2115 ) | ( n4363  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4502 = ( n2369  &  n2370 ) | ( n3829  &  n2370 ) | ( n2369  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4503 = ( n4365  &  n2141 ) | ( n3827  &  n2141 ) | ( n4365  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4504 = ( n2375  &  n2376 ) | ( n3829  &  n2376 ) | ( n2375  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4505 = ( n2214  &  n2425 ) | ( n3827  &  n2425 ) | ( n2214  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4506 = ( n2367  &  n2368 ) | ( n3829  &  n2368 ) | ( n2367  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4507 = ( n4368  &  n2422 ) | ( n3827  &  n2422 ) | ( n4368  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4508 = ( n2365  &  n2366 ) | ( n3829  &  n2366 ) | ( n2365  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4509 = ( n2244  &  n2414 ) | ( n3827  &  n2414 ) | ( n2244  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4510 = ( n2373  &  n2374 ) | ( n3829  &  n2374 ) | ( n2373  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4511 = ( n4371  &  n2410 ) | ( n3827  &  n2410 ) | ( n4371  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4512 = ( n2371  &  n2372 ) | ( n3829  &  n2372 ) | ( n2371  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4513 = ( n2363  &  n2364 ) | ( n3825  &  n2364 ) | ( n2363  &  n3826 ) | ( n3825  &  n3826 ) ;
 assign n4514 = ( (~ n2380)  &  n3777 ) | ( (~ n2380)  &  n4501  &  n4502 ) ;
 assign n4516 = ( n4513  &  n4514  &  Pi24 ) | ( n4513  &  n4514  &  n2377 ) ;
 assign n4517 = ( (~ n2383)  &  n3778 ) | ( (~ n2383)  &  n4507  &  n4508 ) ;
 assign n4519 = ( n4517  &  n3582 ) | ( n4517  &  n4510  &  n4509 ) ;
 assign n4520 = ( n2321  &  n3576 ) | ( n2321  &  n4512  &  n4511 ) ;
 assign n4521 = ( n4373  &  n2162 ) | ( n3827  &  n2162 ) | ( n4373  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4522 = ( n2342  &  n2343 ) | ( n3829  &  n2343 ) | ( n2342  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4523 = ( n4375  &  n2182 ) | ( n3827  &  n2182 ) | ( n4375  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4524 = ( n2348  &  n2349 ) | ( n3829  &  n2349 ) | ( n2348  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4525 = ( n2271  &  n2447 ) | ( n3827  &  n2447 ) | ( n2271  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4526 = ( n2340  &  n2341 ) | ( n3829  &  n2341 ) | ( n2340  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4527 = ( n4378  &  n2444 ) | ( n3827  &  n2444 ) | ( n4378  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4528 = ( n2338  &  n2339 ) | ( n3829  &  n2339 ) | ( n2338  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4529 = ( n2297  &  n2436 ) | ( n3827  &  n2436 ) | ( n2297  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4530 = ( n2346  &  n2347 ) | ( n3829  &  n2347 ) | ( n2346  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4531 = ( n4381  &  n2433 ) | ( n3827  &  n2433 ) | ( n4381  &  n3828 ) | ( n3827  &  n3828 ) ;
 assign n4532 = ( n2344  &  n2345 ) | ( n3829  &  n2345 ) | ( n2344  &  n3830 ) | ( n3829  &  n3830 ) ;
 assign n4533 = ( n2336  &  n2337 ) | ( n3825  &  n2337 ) | ( n2336  &  n3826 ) | ( n3825  &  n3826 ) ;
 assign n4534 = ( (~ n2353)  &  n3777 ) | ( (~ n2353)  &  n4521  &  n4522 ) ;
 assign n4536 = ( (~ n2356)  &  n3778 ) | ( (~ n2356)  &  n4527  &  n4528 ) ;
 assign n4539 = ( n2456  &  n3798 ) | ( n2456  &  (~ n3920) ) | ( n3798  &  (~ n3922) ) | ( (~ n3920)  &  (~ n3922) ) ;
 assign n4540 = ( n2369  &  n2370 ) | ( n3834  &  n2370 ) | ( n2369  &  n1157 ) | ( n3834  &  n1157 ) ;
 assign n4541 = ( n2367  &  n2368 ) | ( n3834  &  n2368 ) | ( n2367  &  n1157 ) | ( n3834  &  n1157 ) ;
 assign n4542 = ( n2365  &  n2366 ) | ( n3834  &  n2366 ) | ( n2365  &  n1157 ) | ( n3834  &  n1157 ) ;
 assign n4544 = ( n2462 ) | ( (~ n2939) ) ;
 assign n4543 = ( n4544  &  n2363 ) | ( n4544  &  n3832 ) ;
 assign n4545 = ( n2342  &  n2343 ) | ( n3834  &  n2343 ) | ( n2342  &  n1157 ) | ( n3834  &  n1157 ) ;
 assign n4546 = ( n2340  &  n2341 ) | ( n3834  &  n2341 ) | ( n2340  &  n1157 ) | ( n3834  &  n1157 ) ;
 assign n4547 = ( n2338  &  n2339 ) | ( n3834  &  n2339 ) | ( n2338  &  n1157 ) | ( n3834  &  n1157 ) ;
 assign n4548 = ( n4544  &  n2336 ) | ( n4544  &  n3832 ) ;
 assign n4549 = ( n2375  &  n2376 ) | ( n3834  &  n2376 ) | ( n2375  &  n1157 ) | ( n3834  &  n1157 ) ;
 assign n4550 = ( n2373  &  n2374 ) | ( n3834  &  n2374 ) | ( n2373  &  n1157 ) | ( n3834  &  n1157 ) ;
 assign n4551 = ( n2371  &  n2372 ) | ( n3834  &  n2372 ) | ( n2371  &  n1157 ) | ( n3834  &  n1157 ) ;
 assign n4552 = ( n4544  &  n2364 ) | ( n4544  &  n3832 ) ;
 assign n4553 = ( n2348  &  n2349 ) | ( n3834  &  n2349 ) | ( n2348  &  n1157 ) | ( n3834  &  n1157 ) ;
 assign n4554 = ( n2346  &  n2347 ) | ( n3834  &  n2347 ) | ( n2346  &  n1157 ) | ( n3834  &  n1157 ) ;
 assign n4555 = ( n2344  &  n2345 ) | ( n3834  &  n2345 ) | ( n2344  &  n1157 ) | ( n3834  &  n1157 ) ;
 assign n4556 = ( n2337 ) | ( n3832 ) ;
 assign n4557 = ( n2481  &  n2499 ) | ( n3742  &  n2499 ) | ( n2481  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4558 = ( n2472  &  n2490 ) | ( n3763  &  n2490 ) | ( n2472  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4560 = ( n2407 ) | ( n2464 ) ;
 assign n4559 = ( n4560  &  n3113 ) | ( n4560  &  n4558  &  n4557 ) ;
 assign n4561 = ( n2302  &  n2314 ) | ( n2302  &  n3499 ) | ( n2314  &  (~ n3784) ) | ( n3499  &  (~ n3784) ) ;
 assign n4562 = ( n1644  &  (~ n2916)  &  (~ n2920) ) | ( n2390  &  (~ n2916)  &  (~ n2920) ) ;
 assign n4565 = ( (~ Pi26)  &  (~ Ni40) ) | ( (~ Pi26)  &  n3860 ) | ( (~ Ni40)  &  n3861 ) | ( n3860  &  n3861 ) ;
 assign n4566 = ( (~ Pi27)  &  (~ Ni41) ) | ( (~ Pi27)  &  n3860 ) | ( (~ Ni41)  &  n3861 ) | ( n3860  &  n3861 ) ;
 assign n4567 = ( n3133  &  n3141 ) | ( n1997  &  n3141 ) | ( n3133  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4568 = ( n3154  &  n3161 ) | ( n1997  &  n3161 ) | ( n3154  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4569 = ( n3186  &  n3192 ) | ( n1997  &  n3192 ) | ( n3186  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4570 = ( n3199  &  n3206 ) | ( n1997  &  n3206 ) | ( n3199  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4571 = ( n3214  &  n3219 ) | ( n1997  &  n3219 ) | ( n3214  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4572 = ( n3226  &  n3233 ) | ( n1997  &  n3233 ) | ( n3226  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4574 = ( n3270 ) | ( n1480 ) ;
 assign n4573 = ( n4574  &  n3777 ) | ( n4574  &  n4567  &  n3260 ) ;
 assign n4575 = ( (~ n3275)  &  n3778 ) | ( n3260  &  (~ n3275)  &  n4570 ) ;
 assign n4577 = ( n3576  &  (~ n3617) ) | ( n3260  &  (~ n3617)  &  n4572 ) ;
 assign n4579 = ( n3168  &  n3170 ) | ( n1997  &  n3170 ) | ( n3168  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4580 = ( n3175  &  n3177 ) | ( n1997  &  n3177 ) | ( n3175  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4581 = ( n3239  &  n3241 ) | ( n1997  &  n3241 ) | ( n3239  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4582 = ( n3243  &  n3245 ) | ( n1997  &  n3245 ) | ( n3243  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4583 = ( n3250  &  n3252 ) | ( n1997  &  n3252 ) | ( n3250  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4584 = ( n3254  &  n3256 ) | ( n1997  &  n3256 ) | ( n3254  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4585 = ( n3262 ) | ( n1480 ) ;
 assign n4588 = ( n3207  &  n3246 ) | ( n3742  &  n3246 ) | ( n3207  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4589 = ( n3234  &  n3257 ) | ( n3763  &  n3257 ) | ( n3234  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4590 = ( n3146  &  n3172 ) | ( n3742  &  n3172 ) | ( n3146  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4591 = ( n3165  &  n3179 ) | ( n3763  &  n3179 ) | ( n3165  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4592 = ( n3280  &  n3282 ) | ( n1997  &  n3282 ) | ( n3280  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4593 = ( n3286  &  n3287 ) | ( n1997  &  n3287 ) | ( n3286  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4594 = ( n3301  &  n3302 ) | ( n1997  &  n3302 ) | ( n3301  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4595 = ( n3303  &  n3304 ) | ( n1997  &  n3304 ) | ( n3303  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4596 = ( n3308  &  n3309 ) | ( n1997  &  n3309 ) | ( n3308  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4597 = ( n3310  &  n3311 ) | ( n1997  &  n3311 ) | ( n3310  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4599 = ( n3334 ) | ( n1480 ) ;
 assign n4598 = ( n4599  &  n3777 ) | ( n4599  &  n4592  &  n3260 ) ;
 assign n4600 = ( (~ n3339)  &  n3778 ) | ( n3260  &  (~ n3339)  &  n4595 ) ;
 assign n4602 = ( n3576  &  (~ n3617) ) | ( n3260  &  (~ n3617)  &  n4597 ) ;
 assign n4603 = ( n3291  &  n3292 ) | ( n1997  &  n3292 ) | ( n3291  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4604 = ( n3296  &  n3297 ) | ( n1997  &  n3297 ) | ( n3296  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4605 = ( n3315  &  n3316 ) | ( n1997  &  n3316 ) | ( n3315  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4606 = ( n3317  &  n3318 ) | ( n1997  &  n3318 ) | ( n3317  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4607 = ( n3322  &  n3323 ) | ( n1997  &  n3323 ) | ( n3322  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4608 = ( n3324  &  n3325 ) | ( n1997  &  n3325 ) | ( n3324  &  n787 ) | ( n1997  &  n787 ) ;
 assign n4609 = ( n3329 ) | ( n1480 ) ;
 assign n4612 = ( n3305  &  n3319 ) | ( n3742  &  n3319 ) | ( n3305  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4613 = ( n3312  &  n3326 ) | ( n3763  &  n3326 ) | ( n3312  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4614 = ( n3284  &  n3294 ) | ( n3742  &  n3294 ) | ( n3284  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4615 = ( n3289  &  n3299 ) | ( n3763  &  n3299 ) | ( n3289  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4616 = ( n3080  &  n3351 ) | ( n3421  &  n3351 ) | ( n3080  &  n1480 ) | ( n3421  &  n1480 ) ;
 assign n4617 = ( n3082  &  n3354 ) | ( n3421  &  n3354 ) | ( n3082  &  n1480 ) | ( n3421  &  n1480 ) ;
 assign n4619 = ( n3098  &  n3376 ) | ( n3421  &  n3376 ) | ( n3098  &  n1480 ) | ( n3421  &  n1480 ) ;
 assign n4620 = ( n3099  &  n3380 ) | ( n3421  &  n3380 ) | ( n3099  &  n1480 ) | ( n3421  &  n1480 ) ;
 assign n4621 = ( n3101  &  n3387 ) | ( n3421  &  n3387 ) | ( n3101  &  n1480 ) | ( n3421  &  n1480 ) ;
 assign n4622 = ( n3102  &  n3391 ) | ( n3421  &  n3391 ) | ( n3102  &  n1480 ) | ( n3421  &  n1480 ) ;
 assign n4623 = ( (~ n3467)  &  n3778 ) | ( n3425  &  (~ n3467)  &  n4620 ) ;
 assign n4625 = ( (~ n3469)  &  n3576 ) | ( n3425  &  (~ n3469)  &  n4622 ) ;
 assign n4627 = ( n3092  &  n3389 ) | ( n3421  &  n3389 ) | ( n3092  &  n1480 ) | ( n3421  &  n1480 ) ;
 assign n4628 = ( n3093  &  n3393 ) | ( n3421  &  n3393 ) | ( n3093  &  n1480 ) | ( n3421  &  n1480 ) ;
 assign n4629 = ( n3461  &  n3462 ) | ( n1884  &  n3462 ) | ( n3461  &  n3778 ) | ( n1884  &  n3778 ) ;
 assign n4631 = ( n3454  &  n3459 ) | ( n3870  &  n3459 ) | ( n3454  &  n3871 ) | ( n3870  &  n3871 ) ;
 assign n4632 = ( n3006  &  n3368 ) | ( n3421  &  n3368 ) | ( n3006  &  n1480 ) | ( n3421  &  n1480 ) ;
 assign n4633 = ( n3012  &  n3370 ) | ( n3421  &  n3370 ) | ( n3012  &  n1480 ) | ( n3421  &  n1480 ) ;
 assign n4635 = ( n3044  &  n3398 ) | ( n3421  &  n3398 ) | ( n3044  &  n1480 ) | ( n3421  &  n1480 ) ;
 assign n4636 = ( n3049  &  n3402 ) | ( n3421  &  n3402 ) | ( n3049  &  n1480 ) | ( n3421  &  n1480 ) ;
 assign n4637 = ( n3052  &  n3409 ) | ( n3421  &  n3409 ) | ( n3052  &  n1480 ) | ( n3421  &  n1480 ) ;
 assign n4638 = ( n3058  &  n3413 ) | ( n3421  &  n3413 ) | ( n3058  &  n1480 ) | ( n3421  &  n1480 ) ;
 assign n4639 = ( (~ n3446)  &  n3778 ) | ( n3425  &  (~ n3446)  &  n4636 ) ;
 assign n4641 = ( (~ n3448)  &  n3576 ) | ( n3425  &  (~ n3448)  &  n4638 ) ;
 assign n4643 = ( n3029  &  n3411 ) | ( n3421  &  n3411 ) | ( n3029  &  n1480 ) | ( n3421  &  n1480 ) ;
 assign n4644 = ( n3034  &  n3415 ) | ( n3421  &  n3415 ) | ( n3034  &  n1480 ) | ( n3421  &  n1480 ) ;
 assign n4645 = ( n3439  &  n3440 ) | ( n1884  &  n3440 ) | ( n3439  &  n3778 ) | ( n1884  &  n3778 ) ;
 assign n4647 = ( n3429  &  n3437 ) | ( n3870  &  n3437 ) | ( n3429  &  n3871 ) | ( n3870  &  n3871 ) ;
 assign n4648 = ( n3384  &  n3406 ) | ( n3742  &  n3406 ) | ( n3384  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4649 = ( n3395  &  n3417 ) | ( n3763  &  n3417 ) | ( n3395  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4650 = ( n3349  &  n3366 ) | ( n3742  &  n3366 ) | ( n3349  &  n3754 ) | ( n3742  &  n3754 ) ;
 assign n4652 = ( n3358  &  n3374 ) | ( n3763  &  n3374 ) | ( n3358  &  n3774 ) | ( n3763  &  n3774 ) ;
 assign n4654 = ( n3798 ) | ( n1068 ) | ( n4785 ) | ( n4786 ) ;
 assign n4657 = ( n168 ) | ( (~ Ni10) ) | ( n1654 ) | ( n3492 ) ;
 assign n4658 = ( n3492 ) | ( n3613 ) | ( n3614 ) ;
 assign n4659 = ( Ni31  &  (~ Ni30) ) | ( Ni31  &  (~ Ni5) ) | ( Ni31  &  Ni4 ) ;
 assign n4665 = ( Pi15  &  n773 ) | ( (~ Pi15)  &  n781 ) | ( n773  &  n781 ) ;
 assign n4666 = ( (~ Pi17)  &  n758 ) | ( (~ Pi17)  &  n763 ) | ( (~ Pi17)  &  (~ n4006) ) ;
 assign n4667 = ( (~ Pi17)  &  (~ n4666) ) | ( n4008  &  n4009  &  (~ n4666) ) ;
 assign n4669 = ( n3113  &  n4665 ) | ( (~ n3113)  &  n4667 ) | ( n4665  &  n4667 ) ;
 assign n4670 = ( (~ n3775)  &  n4027  &  n4028 ) ;
 assign n4671 = ( (~ n1654)  &  n4670 ) | ( (~ n1654)  &  n3775  &  n4667 ) ;
 assign n4672 = ( (~ Ni7)  &  n4671 ) | ( n1654  &  (~ Ni7)  &  n4669 ) ;
 assign n4673 = ( (~ n3540)  &  n4672 ) | ( (~ n3540)  &  Ni7  &  n4669 ) ;
 assign n4675 = ( n4186  &  n3650  &  Ni14 ) ;
 assign n4676 = ( (~ Ni14)  &  n4100  &  n4101 ) ;
 assign n4677 = ( n4108  &  n4107  &  Ni14 ) ;
 assign n4678 = ( (~ n848) ) | ( (~ n1053) ) | ( n1505 ) | ( n1508 ) | ( n1511 ) | ( n1514 ) | ( n1517 ) | ( (~ n4068) ) ;
 assign n4682 = ( (~ n848) ) | ( (~ n994) ) | ( n1482 ) | ( n1487 ) | ( n1490 ) | ( n1494 ) | ( n1498 ) | ( (~ n4082) ) ;
 assign n4686 = ( n1332 ) | ( n3792 ) ;
 assign n4685 = ( (~ Pi15)  &  n4139  &  n4142  &  n4145  &  n4146  &  n4686 ) ;
 assign n4688 = ( n1402 ) | ( n3792 ) ;
 assign n4687 = ( n4159  &  n4688  &  n4162  &  n4166  &  n4165  &  Pi15 ) ;
 assign n4689 = ( Pi17  &  (~ n4051) ) | ( Pi17  &  (~ n4053) ) ;
 assign n4691 = ( (~ Pi17)  &  n848  &  n4084  &  n4085 ) ;
 assign n4692 = ( n4088  &  n848  &  n4087  &  Pi17 ) ;
 assign n4693 = ( n4174  &  Ni10  &  Ni11 ) | ( n4174  &  Ni10  &  n1414 ) ;
 assign n4696 = ( (~ Pi17)  &  n4089  &  n4090 ) ;
 assign n4699 = ( n2010 ) | ( n3576 ) ;
 assign n4698 = ( (~ Pi15)  &  n1995  &  n4236  &  n4238  &  n4239  &  n4699 ) ;
 assign n4701 = ( n18 ) | ( (~ Ni34) ) ;
 assign n4702 = ( Ni34 ) | ( n18 ) | ( n1063 ) ;
 assign n4703 = ( (~ Pi17)  &  n4255  &  n4256 ) ;
 assign n4704 = ( n4258  &  n4257  &  Pi17 ) ;
 assign n4705 = ( Pi20  &  (~ n4281) ) | ( Pi20  &  (~ n4285) ) ;
 assign n4706 = ( Pi20  &  (~ n4705) ) | ( n4269  &  n4272  &  (~ n4705) ) ;
 assign n4708 = ( Pi20  &  (~ n4311) ) | ( Pi20  &  (~ n4315) ) ;
 assign n4709 = ( Pi20  &  (~ n4708) ) | ( n4299  &  n4302  &  (~ n4708) ) ;
 assign n4711 = ( (~ Pi15)  &  n4287  &  n4706 ) ;
 assign n4712 = ( n4317  &  n4709  &  Pi15 ) ;
 assign n4713 = ( n4703 ) | ( n4704 ) | ( n3113 ) | ( Ni10 ) ;
 assign n4714 = ( (~ Pi17)  &  (~ n4326) ) | ( (~ Pi17)  &  (~ n4328) ) ;
 assign n4716 = ( n4332  &  n2024  &  n2031 ) ;
 assign n4717 = ( (~ n2031)  &  n3660 ) | ( (~ Pi23)  &  n2026  &  (~ n2031) ) ;
 assign n4718 = ( n4333  &  n2043  &  n2031 ) ;
 assign n4719 = ( (~ n2031)  &  n3663 ) | ( (~ Pi24)  &  (~ n2031)  &  n2046 ) ;
 assign n4720 = ( Ni33  &  (~ n2031)  &  n2046 ) | ( n275  &  (~ n2031)  &  n2046 ) ;
 assign n4722 = ( (~ Ni44)  &  (~ n3572)  &  (~ Ni39) ) | ( (~ Ni44)  &  Ni42  &  (~ Ni39) ) ;
 assign n4724 = ( (~ Ni44)  &  (~ n4722) ) | ( (~ n320)  &  (~ n4722) ) | ( (~ Ni39)  &  (~ n4722) ) ;
 assign n4730 = ( Pi21 ) | ( n3674 ) ;
 assign n4733 = ( Pi26  &  (~ n2327) ) | ( (~ Pi26)  &  (~ n2329) ) | ( (~ n2327)  &  (~ n2329) ) ;
 assign n4735 = ( (~ Pi21)  &  (~ n2303) ) | ( (~ Pi26)  &  (~ Pi21)  &  Ni32 ) ;
 assign n4737 = ( (~ Pi26)  &  (~ n2327) ) | ( Pi26  &  (~ n2329) ) | ( (~ n2327)  &  (~ n2329) ) ;
 assign n4738 = ( (~ Ni14)  &  n4405  &  n4406 ) ;
 assign n4740 = ( (~ n2070) ) | ( (~ n2377) ) | ( n2782 ) | ( n2785 ) | ( n2788 ) | ( n2791 ) | ( n2794 ) | ( (~ n4372) ) ;
 assign n4743 = ( (~ n2070) ) | ( (~ n2350) ) | ( n2764 ) | ( n2767 ) | ( n2770 ) | ( n2773 ) | ( n2776 ) | ( (~ n4382) ) ;
 assign n4747 = ( n2632 ) | ( n3792 ) ;
 assign n4746 = ( (~ Pi15)  &  n4440  &  n4443  &  n4446  &  n4447  &  n4747 ) ;
 assign n4749 = ( n2688 ) | ( n3792 ) ;
 assign n4748 = ( n4460  &  n4749  &  n4463  &  n4467  &  n4466  &  Pi15 ) ;
 assign n4750 = ( Pi17  &  (~ n4359) ) | ( Pi17  &  (~ n4361) ) ;
 assign n4752 = ( (~ Pi17)  &  n2070  &  n4384  &  n4385 ) ;
 assign n4753 = ( n4388  &  n2070  &  n4387  &  Pi17 ) ;
 assign n4754 = ( n4475  &  Ni10  &  Ni11 ) | ( n4475  &  Ni10  &  n2699 ) ;
 assign n4755 = ( n2397 ) | ( n2401 ) | ( n2404 ) ;
 assign n4756 = ( (~ Pi17)  &  n4394  &  n4395 ) ;
 assign n4759 = ( (~ Pi20)  &  n2937  &  n3858 ) | ( (~ Pi20)  &  (~ Ni39)  &  n3858 ) ;
 assign n4760 = ( n3858  &  Pi20  &  Ni39 ) | ( n3858  &  Pi20  &  n2937 ) ;
 assign n4761 = ( (~ n2031) ) | ( (~ Ni40) ) ;
 assign n4763 = ( (~ n2031)  &  n3686 ) | ( n2031  &  (~ n3925) ) | ( n3686  &  (~ n3925) ) ;
 assign n4764 = ( (~ n2031) ) | ( (~ Ni41) ) ;
 assign n4766 = ( (~ n2031)  &  n3692 ) | ( n2031  &  (~ n3931) ) | ( n3692  &  (~ n3931) ) ;
 assign n4767 = ( (~ Pi21)  &  n171 ) | ( (~ Pi21)  &  (~ n1063)  &  n2946 ) ;
 assign n4769 = ( Pi20  &  n3463 ) | ( Pi20  &  n3465 ) | ( Pi20  &  (~ n4629) ) ;
 assign n4770 = ( Pi20  &  (~ n4769) ) | ( n4623  &  n4625  &  (~ n4769) ) ;
 assign n4772 = ( Pi20  &  n3441 ) | ( Pi20  &  n3444 ) | ( Pi20  &  (~ n4645) ) ;
 assign n4773 = ( Pi20  &  (~ n4772) ) | ( n4639  &  n4641  &  (~ n4772) ) ;
 assign n4775 = ( (~ Pi15)  &  n4631  &  n4770 ) ;
 assign n4776 = ( n4647  &  n4773  &  Pi15 ) ;
 assign n4777 = ( (~ Pi17)  &  n4648  &  n4649 ) ;
 assign n4779 = ( (~ Ni10)  &  n4775 ) | ( (~ Ni10)  &  n4776 ) ;
 assign n4780 = ( (~ Pi15)  &  (~ n3271)  &  (~ n3273)  &  n4573  &  n4575  &  n4577 ) ;
 assign n4783 = ( (~ Pi17)  &  n4588  &  n4589 ) ;
 assign n4784 = ( n4591  &  n4590  &  Pi17 ) ;
 assign n4785 = ( (~ Ni10)  &  n4780 ) | ( Pi15  &  (~ Ni10)  &  n3937 ) ;
 assign n4786 = ( Ni10  &  n4783 ) | ( Ni10  &  n4784 ) ;
 assign n4787 = ( (~ Pi15)  &  (~ n3335)  &  (~ n3337)  &  n4598  &  n4600  &  n4602 ) ;
 assign n4790 = ( (~ Pi17)  &  n4612  &  n4613 ) ;
 assign n4791 = ( n4615  &  n4614  &  Pi17 ) ;
 assign n4792 = ( (~ Ni10)  &  n4787 ) | ( Pi15  &  (~ Ni10)  &  n3942 ) ;
 assign n4797 = ( (~ Ni14) ) | ( (~ Ni12) ) | ( n4836 ) ;
 assign n4798 = ( (~ Ni6)  &  (~ Ni4) ) | ( (~ Ni5)  &  (~ Ni4) ) | ( (~ n3527)  &  (~ Ni4) ) ;
 assign n4799 = ( (~ Ni31) ) | ( (~ Ni6) ) | ( (~ Ni5) ) ;
 assign n4800 = ( n4799  &  Ni4  &  n2066 ) | ( n4799  &  Ni4  &  n3874 ) ;
 assign n4801 = ( Ni3  &  n4800 ) | ( (~ Ni4)  &  Ni3  &  (~ n4799) ) ;
 assign n4803 = ( (~ Ni2)  &  n4801 ) | ( (~ Ni2)  &  (~ Ni3)  &  n3952 ) ;
 assign n4805 = ( Ni6  &  Ni2 ) | ( (~ Ni31)  &  Ni6  &  Ni3 ) ;
 assign n4808 = ( Ni12  &  n3540 ) | ( Ni12  &  (~ n3559)  &  n3568 ) ;
 assign n4810 = ( Pi20  &  n184 ) | ( Pi20  &  n3585 ) | ( Pi20  &  n3595 ) ;
 assign n4811 = ( (~ Ni44)  &  Ni42  &  (~ Ni39) ) | ( n3573  &  Ni42  &  (~ Ni39) ) ;
 assign n4813 = ( Pi27 ) | ( n3880 ) ;
 assign n4814 = ( (~ Pi27) ) | ( Pi26 ) | ( n3880 ) ;
 assign n4815 = ( Pi24 ) | ( n3881 ) ;
 assign n4816 = ( (~ Pi24) ) | ( Pi23 ) | ( n3881 ) ;
 assign n4817 = ( n2065  &  (~ Ni4) ) | ( (~ Ni4)  &  n3863 ) ;
 assign n4818 = ( Ni4  &  Ni33 ) | ( Ni4  &  n3874 ) ;
 assign n4819 = ( Ni33  &  (~ n834) ) ;
 assign n4820 = ( (~ Ni33)  &  (~ n834) ) ;
 assign n4822 = ( n63 ) | ( n2086 ) ;
 assign n4823 = ( (~ n38) ) | ( Ni41 ) ;
 assign n4825 = ( (~ n42) ) | ( Ni41 ) ;
 assign n4827 = ( (~ Ni33) ) | ( n2966 ) ;
 assign n4832 = ( n1062  &  n953 ) ;
 assign n4833 = ( n1071 ) | ( n1075 ) | ( n1079 ) | ( (~ n4223) ) ;
 assign n4835 = ( n4759 ) | ( n4760 ) | ( n3879 ) ;
 assign n4836 = ( n3492  &  Pi27 ) ;


endmodule

