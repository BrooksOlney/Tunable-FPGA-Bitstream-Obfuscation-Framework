module apex2_qmap_map (sk, i_36_, i_34_, i_28_, i_29_, i_35_, i_27_, i_23_, i_24_, i_16_, i_13_, i_7_, i_8_, i_12_, i_6_, i_2_, i_4_, i_5_, i_9_, i_17_, i_11_, i_19_, i_3_, i_18_, i_14_, i_10_, i_32_, i_1_, i_31_, i_30_, i_21_, i_26_, i_25_, i_22_, i_33_, i_20_, i_0_, i_37_, i_38_, o_0_, o_1_, o_2_);

	input i_36_;
	input i_34_;
	input i_28_;
	input i_29_;
	input i_35_;
	input i_27_;
	input i_23_;
	input i_24_;
	input i_16_;
	input i_13_;
	input i_7_;
	input i_8_;
	input i_12_;
	input i_6_;
	input i_2_;
	input i_4_;
	input i_5_;
	input i_9_;
	input i_17_;
	input i_11_;
	input i_19_;
	input i_3_;
	input i_18_;
	input i_14_;
	input i_10_;
	input i_32_;
	input i_1_;
	input i_31_;
	input i_30_;
	input i_21_;
	input i_26_;
	input i_25_;
	input i_22_;
	input i_33_;
	input i_20_;
	input i_0_;
	input i_37_;
	input i_38_;
	output o_0_;
	output o_1_;
	output o_2_;



	wire g427, g661, g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19;
	wire g20, g21, g22, g23, g24, g25, g26, g27, g28, g29, g30, g31, g32, g33, g34, g35, g36, g37, g38, g39, g40;
	wire g41, g42, g43, g44, g45, g46, g47, g48, g49, g50, g51, g52, g53, g54, g55, g56, g57, g58, g59, g60, g61;
	wire g62, g63, g64, g65, g66, g67, g68, g69, g70, g71, g72, g73, g74, g75, g76, g77, g78, g79, g80, g81, g82;
	wire g83, g84, g85, g86, g87, g88, g89, g90, g91, g92, g93, g94, g95, g96, g97, g98, g99, g100, g101, g102, g103;
	wire g104, g105, g106, g107, g108, g109, g110, g111, g112, g113, g114, g115, g116, g117, g118, g119, g120, g121, g122, g123, g124;
	wire g125, g126, g127, g128, g129, g130, g131, g132, g133, g134, g135, g136, g137, g138, g139, g140, g141, g142, g143, g144, g145;
	wire g146, g147, g148, g149, g150, g151, g152, g153, g154, g155, g156, g157, g158, g159, g160, g161, g162, g163, g164, g165, g166;
	wire g167, g168, g169, g170, g171, g172, g173, g174, g175, g176, g177, g178, g179, g180, g181, g182, g183, g712, g184, g185, g186;
	wire g187, g188, g189, g190, g191, g192, g193, g194, g195, g196, g197, g198, g199, g200, g201, g202, g203, g204, g205, g206, g207;
	wire g208, g209, g210, g211, g212, g213, g214, g215, g216, g217, g218, g219, g220, g702, g221, g222, g223, g224, g225, g226, g227;
	wire g228, g229, g230, g231, g232, g233, g234, g235, g236, g237, g238, g239, g240, g241, g242, g243, g244, g245, g247, g248, g249;
	wire g250, g251, g252, g253, g254, g255, g256, g257, g258, g259, g260, g261, g262, g263, g264, g265, g266, g267, g268, g269, g270;
	wire g271, g272, g273, g274, g275, g276, g277, g278, g279, g280, g281, g282, g283, g284, g285, g286, g287, g288, g289, g290, g291;
	wire g292, g293, g294, g295, g296, g297, g298, g299, g300, g301, g302, g303, g304, g305, g306, g307, g308, g309, g310, g311, g312;
	wire g313, g314, g315, g316, g317, g318, g319, g320, g321, g322, g323, g324, g325, g326, g327, g328, g329, g330, g331, g332, g333;
	wire g334, g335, g336, g337, g338, g339, g340, g341, g342, g343, g344, g345, g346, g347, g348, g349, g350, g351, g352, g353, g354;
	wire g355, g356, g357, g358, g359, g360, g361, g362, g363, g364, g365, g366, g367, g368, g369, g370, g371, g372, g373, g374, g375;
	wire g376, g377, g378, g379, g380, g381, g382, g383, g384, g385, g386, g387, g388, g389, g390, g391, g392, g393, g394, g395, g396;
	wire g397, g398, g399, g400, g401, g402, g403, g404, g405, g406, g407, g408, g409, g410, g411, g412, g413, g414, g415, g416, g417;
	wire g418, g419, g420, g421, g422, g423, g424, g425, g426, g428, g429, g430, g431, g432, g433, g434, g435, g436, g437, g438, g439;
	wire g440, g441, g442, g443, g444, g445, g446, g447, g448, g449, g450, g451, g452, g453, g454, g455, g456, g457, g458, g459, g460;
	wire g461, g462, g463, g464, g465, g466, g467, g468, g469, g470, g471, g472, g473, g474, g475, g696, g476, g477, g478, g479, g480;
	wire g481, g482, g483, g484, g485, g486, g487, g488, g489, g490, g491, g492, g493, g494, g495, g496, g497, g498, g499, g500, g501;
	wire g502, g503, g504, g505, g506, g507, g508, g509, g510, g511, g512, g513, g514, g515, g516, g517, g518, g519, g520, g521, g522;
	wire g523, g524, g525, g526, g527, g528, g529, g530, g531, g532, g533, g534, g535, g536, g537, g538, g539, g540, g541, g542, g543;
	wire g544, g545, g546, g547, g548, g549, g550, g551, g552, g553, g554, g555, g556, g557, g558, g559, g560, g561, g562, g563, g564;
	wire g565, g566, g567, g568, g569, g570, g571, g572, g573, g574, g575, g576, g577, g578, g579, g580, g685, g581, g582, g583, g584;
	wire g585, g586, g587, g588, g589, g590, g591, g592, g593, g594, g595, g596, g597, g598, g599, g600, g601, g602, g603, g604, g605;
	wire g606, g607, g608, g609, g610, g611, g612, g613, g614, g615, g616, g617, g618, g619, g620, g621, g672, g622, g623, g624, g625;
	wire g626, g627, g628, g629, g630, g631, g632, g633, g634, g635, g636, g637, g638, g639, g640, g641, g642, g643, g644, g645, g646;
	wire g647, g648, g649, g662, g650, g651, g652, g653, g654, g655, g656, g657, g658, g659, g660, g663, g664, g665, g666, g669, g667;
	wire g668, g670, g671, g673, g674, g675, g678, g676, g677, g681, g682, g679, g680, g683, g684, g686, g687, g688, g691, g689, g690;
	wire g693, g694, g692, g695, g697, g698, g699, g700, g701, g703, g704, g705, g706, g709, g707, g708, g710, g711, g713, g714, g715;
	wire g716, g717, g718;

	lut_sub lut_5 ({g427}, o_1_);
	defparam lut_5.LUT_SIZE = 1;
	defparam lut_5.mask = 2'b10;

	lut_sub lut_9 ({g661}, o_2_);
	defparam lut_9.LUT_SIZE = 1;
	defparam lut_9.mask = 2'b10;

	lut_sub lut_13 ({i_28_, i_29_}, g1);
	defparam lut_13.LUT_SIZE = 2;
	defparam lut_13.mask = 4'b1000;

	lut_sub lut_17 ({i_34_, i_35_}, g2);
	defparam lut_17.LUT_SIZE = 2;
	defparam lut_17.mask = 4'b0100;

	lut_sub lut_21 ({i_27_, i_28_, i_23_}, g3);
	defparam lut_21.LUT_SIZE = 3;
	defparam lut_21.mask = 8'h80;

	lut_sub lut_27 ({g2, g3, i_29_}, g4);
	defparam lut_27.LUT_SIZE = 3;
	defparam lut_27.mask = 8'h02;

	lut_sub lut_31 ({i_24_, i_27_, i_23_}, g5);
	defparam lut_31.LUT_SIZE = 3;
	defparam lut_31.mask = 8'h7f;

	lut_sub lut_44 ({i_34_, g1, g4, g5}, g6);
	defparam lut_44.LUT_SIZE = 4;
	defparam lut_44.mask = 16'hccc4;

	lut_sub lut_54 ({i_7_, i_8_}, g7);
	defparam lut_54.LUT_SIZE = 2;
	defparam lut_54.mask = 4'b1000;

	lut_sub lut_58 ({i_2_, i_4_, i_5_}, g8);
	defparam lut_58.LUT_SIZE = 3;
	defparam lut_58.mask = 8'h80;

	lut_sub lut_63 ({i_12_, i_6_, g8}, g9);
	defparam lut_63.LUT_SIZE = 3;
	defparam lut_63.mask = 8'h40;

	lut_sub lut_67 ({i_2_, i_9_, i_6_, i_4_, i_5_}, g10);
	defparam lut_67.LUT_SIZE = 5;
	defparam lut_67.mask = 32'h80000000;

	lut_sub lut_73 ({g7, g10}, g11);
	defparam lut_73.LUT_SIZE = 2;
	defparam lut_73.mask = 4'b0001;

	lut_sub lut_77 ({i_11_, i_19_}, g12);
	defparam lut_77.LUT_SIZE = 2;
	defparam lut_77.mask = 4'b1000;

	lut_sub lut_82 ({i_17_, g12}, g13);
	defparam lut_82.LUT_SIZE = 2;
	defparam lut_82.mask = 4'b0100;

	lut_sub lut_86 ({i_6_, i_4_, i_5_}, g14);
	defparam lut_86.LUT_SIZE = 3;
	defparam lut_86.mask = 8'h80;

	lut_sub lut_90 ({i_17_, i_9_, i_18_}, g15);
	defparam lut_90.LUT_SIZE = 3;
	defparam lut_90.mask = 8'h80;

	lut_sub lut_96 ({i_2_, i_7_, i_3_, g14, g15}, g16);
	defparam lut_96.LUT_SIZE = 5;
	defparam lut_96.mask = 32'h01000000;

	lut_sub lut_103 ({i_16_, i_8_, g11, g13, g16}, g17);
	defparam lut_103.LUT_SIZE = 5;
	defparam lut_103.mask = 32'h57030000;

	lut_sub lut_116 ({i_16_, i_13_, g7, g9, g17}, g18);
	defparam lut_116.LUT_SIZE = 5;
	defparam lut_116.mask = 32'h57005500;

	lut_sub lut_128 ({i_27_, i_28_}, g19);
	defparam lut_128.LUT_SIZE = 2;
	defparam lut_128.mask = 4'b1000;

	lut_sub lut_133 ({i_24_, g19}, g20);
	defparam lut_133.LUT_SIZE = 2;
	defparam lut_133.mask = 4'b0100;

	lut_sub lut_138 ({g20, i_29_}, g21);
	defparam lut_138.LUT_SIZE = 2;
	defparam lut_138.mask = 4'b0010;

	lut_sub lut_142 ({i_13_, i_14_}, g22);
	defparam lut_142.LUT_SIZE = 2;
	defparam lut_142.mask = 4'b0001;

	lut_sub lut_146 ({i_16_, i_17_, i_23_}, g23);
	defparam lut_146.LUT_SIZE = 3;
	defparam lut_146.mask = 8'h80;

	lut_sub lut_150 ({i_13_, i_10_}, g24);
	defparam lut_150.LUT_SIZE = 2;
	defparam lut_150.mask = 4'b0100;

	lut_sub lut_156 ({g11, g24}, g25);
	defparam lut_156.LUT_SIZE = 2;
	defparam lut_156.mask = 4'b0010;

	lut_sub lut_163 ({g22, g23, g25}, g26);
	defparam lut_163.LUT_SIZE = 3;
	defparam lut_163.mask = 8'h10;

	lut_sub lut_167 ({i_16_, i_13_, i_14_, i_10_}, g27);
	defparam lut_167.LUT_SIZE = 4;
	defparam lut_167.mask = 16'hac00;

	lut_sub lut_174 ({i_16_, i_13_, i_14_}, g28);
	defparam lut_174.LUT_SIZE = 3;
	defparam lut_174.mask = 8'he0;

	lut_sub lut_181 ({i_2_, g14, i_1_}, g29);
	defparam lut_181.LUT_SIZE = 3;
	defparam lut_181.mask = 8'h20;

	lut_sub lut_187 ({g28, i_7_, i_8_, g29}, g30);
	defparam lut_187.LUT_SIZE = 4;
	defparam lut_187.mask = 16'h0040;

	lut_sub lut_191 ({i_7_, i_9_, i_6_}, g31);
	defparam lut_191.LUT_SIZE = 3;
	defparam lut_191.mask = 8'h80;

	lut_sub lut_197 ({g8, g31}, g32);
	defparam lut_197.LUT_SIZE = 2;
	defparam lut_197.mask = 4'b0001;

	lut_sub lut_201 ({i_24_, i_23_}, g33);
	defparam lut_201.LUT_SIZE = 2;
	defparam lut_201.mask = 4'b1000;

	lut_sub lut_205 ({i_27_, i_28_, i_29_}, g34);
	defparam lut_205.LUT_SIZE = 3;
	defparam lut_205.mask = 8'h80;

	lut_sub lut_211 ({i_17_, g33, g34}, g35);
	defparam lut_211.LUT_SIZE = 3;
	defparam lut_211.mask = 8'h10;

	lut_sub lut_219 ({i_32_, g27, g30, g32, g35}, g36);
	defparam lut_219.LUT_SIZE = 5;
	defparam lut_219.mask = 32'h05150505;

	lut_sub lut_232 ({i_32_, g1}, g37);
	defparam lut_232.LUT_SIZE = 2;
	defparam lut_232.mask = 4'b0100;

	lut_sub lut_236 ({i_27_, i_17_, i_23_}, g38);
	defparam lut_236.LUT_SIZE = 3;
	defparam lut_236.mask = 8'h80;

	lut_sub lut_244 ({g37, g27, g32, g38}, g39);
	defparam lut_244.LUT_SIZE = 4;
	defparam lut_244.mask = 16'h0001;

	lut_sub lut_251 ({i_34_, i_35_, g34, g26, g39}, g40);
	defparam lut_251.LUT_SIZE = 5;
	defparam lut_251.mask = 32'hffa80000;

	lut_sub lut_267 ({i_17_, g28, i_7_, g29}, g41);
	defparam lut_267.LUT_SIZE = 4;
	defparam lut_267.mask = 16'h0400;

	lut_sub lut_273 ({g5, g37}, g42);
	defparam lut_273.LUT_SIZE = 2;
	defparam lut_273.mask = 4'b0100;

	lut_sub lut_279 ({i_34_, g41, g42}, g43);
	defparam lut_279.LUT_SIZE = 3;
	defparam lut_279.mask = 8'h0e;

	lut_sub lut_290 ({g21, g26, g36, g40, g43}, g44);
	defparam lut_290.LUT_SIZE = 5;
	defparam lut_290.mask = 32'h8c8c8ccc;

	lut_sub lut_306 ({i_16_, i_13_}, g45);
	defparam lut_306.LUT_SIZE = 2;
	defparam lut_306.mask = 4'b1000;

	lut_sub lut_310 ({i_2_, i_8_}, g46);
	defparam lut_310.LUT_SIZE = 2;
	defparam lut_310.mask = 4'b1000;

	lut_sub lut_317 ({i_3_, g14, g15, g46}, g47);
	defparam lut_317.LUT_SIZE = 4;
	defparam lut_317.mask = 16'h0001;

	lut_sub lut_321 ({i_9_, i_6_, i_8_}, g48);
	defparam lut_321.LUT_SIZE = 3;
	defparam lut_321.mask = 8'h80;

	lut_sub lut_327 ({g8, g48}, g49);
	defparam lut_327.LUT_SIZE = 2;
	defparam lut_327.mask = 4'b0001;

	lut_sub lut_335 ({i_23_, g45, g13, g47, g49}, g50);
	defparam lut_335.LUT_SIZE = 5;
	defparam lut_335.mask = 32'h00370000;

	lut_sub lut_344 ({i_8_, g9}, g51);
	defparam lut_344.LUT_SIZE = 2;
	defparam lut_344.mask = 4'b0100;

	lut_sub lut_351 ({i_23_, g28, i_31_, g50, g51}, g52);
	defparam lut_351.LUT_SIZE = 5;
	defparam lut_351.mask = 32'hcc8ccccc;

	lut_sub lut_370 ({i_17_, g45}, g53);
	defparam lut_370.LUT_SIZE = 2;
	defparam lut_370.mask = 4'b0100;

	lut_sub lut_374 ({i_16_, i_14_}, g54);
	defparam lut_374.LUT_SIZE = 2;
	defparam lut_374.mask = 4'b1000;

	lut_sub lut_379 ({i_17_, g54}, g55);
	defparam lut_379.LUT_SIZE = 2;
	defparam lut_379.mask = 4'b0100;

	lut_sub lut_386 ({i_13_, g53, g10, i_10_, g55}, g56);
	defparam lut_386.LUT_SIZE = 5;
	defparam lut_386.mask = 32'h000c050d;

	lut_sub lut_396 ({i_32_, i_31_}, g57);
	defparam lut_396.LUT_SIZE = 2;
	defparam lut_396.mask = 4'b1000;

	lut_sub lut_402 ({g29, g23}, g58);
	defparam lut_402.LUT_SIZE = 2;
	defparam lut_402.mask = 4'b0001;

	lut_sub lut_410 ({g20, g22, g57, i_29_, g58}, g59);
	defparam lut_410.LUT_SIZE = 5;
	defparam lut_410.mask = 32'h00000400;

	lut_sub lut_415 ({i_31_, g1}, g60);
	defparam lut_415.LUT_SIZE = 2;
	defparam lut_415.mask = 4'b0100;

	lut_sub lut_421 ({i_17_, g28, i_8_, g29}, g61);
	defparam lut_421.LUT_SIZE = 4;
	defparam lut_421.mask = 16'h0400;

	lut_sub lut_431 ({g5, g27, g60, g61, g49, g35}, g62);
	defparam lut_431.LUT_SIZE = 6;
	defparam lut_431.mask = 64'h000f111f00001111;

	lut_sub lut_453 ({g42, g56, g59, g62}, g63);
	defparam lut_453.LUT_SIZE = 4;
	defparam lut_453.mask = 16'h8880;

	lut_sub lut_462 ({i_34_, i_35_, g52, g21, g63}, g64);
	defparam lut_462.LUT_SIZE = 5;
	defparam lut_462.mask = 32'h0000ba00;

	lut_sub lut_470 ({i_35_, i_32_}, g65);
	defparam lut_470.LUT_SIZE = 2;
	defparam lut_470.mask = 4'b1000;

	lut_sub lut_475 ({i_34_, g65}, g66);
	defparam lut_475.LUT_SIZE = 2;
	defparam lut_475.mask = 4'b0001;

	lut_sub lut_480 ({i_2_, i_9_, i_3_, g14}, g67);
	defparam lut_480.LUT_SIZE = 4;
	defparam lut_480.mask = 16'h1000;

	lut_sub lut_487 ({g33, i_18_, i_11_, i_19_, g67, g10}, g68);
	defparam lut_487.LUT_SIZE = 6;
	defparam lut_487.mask = 64'h0000000073335000;

	lut_sub lut_503 ({g53, g68}, g69);
	defparam lut_503.LUT_SIZE = 2;
	defparam lut_503.mask = 4'b0001;

	lut_sub lut_507 ({i_30_, i_32_}, g70);
	defparam lut_507.LUT_SIZE = 2;
	defparam lut_507.mask = 4'b0111;

	lut_sub lut_513 ({i_24_, i_26_}, g71);
	defparam lut_513.LUT_SIZE = 2;
	defparam lut_513.mask = 4'b0111;

	lut_sub lut_520 ({i_27_, i_23_, i_21_, g71}, g72);
	defparam lut_520.LUT_SIZE = 4;
	defparam lut_520.mask = 16'h8000;

	lut_sub lut_525 ({i_12_, g22, i_7_}, g73);
	defparam lut_525.LUT_SIZE = 3;
	defparam lut_525.mask = 8'h80;

	lut_sub lut_531 ({i_16_, g72, g73}, g74);
	defparam lut_531.LUT_SIZE = 3;
	defparam lut_531.mask = 8'h10;

	lut_sub lut_537 ({i_28_, g70, g74}, g75);
	defparam lut_537.LUT_SIZE = 3;
	defparam lut_537.mask = 8'h40;

	lut_sub lut_542 ({i_24_, i_34_, i_35_, i_32_, g34}, g76);
	defparam lut_542.LUT_SIZE = 5;
	defparam lut_542.mask = 32'h04440400;

	lut_sub lut_550 ({i_7_, g9}, g77);
	defparam lut_550.LUT_SIZE = 2;
	defparam lut_550.mask = 4'b0100;

	lut_sub lut_556 ({g13, g32}, g78);
	defparam lut_556.LUT_SIZE = 2;
	defparam lut_556.mask = 4'b0001;

	lut_sub lut_564 ({i_23_, g45, g77, g16, g78}, g79);
	defparam lut_564.LUT_SIZE = 5;
	defparam lut_564.mask = 32'h007f0000;

	lut_sub lut_580 ({g66, g34, g69, g75, g76, g79}, g80);
	defparam lut_580.LUT_SIZE = 6;
	defparam lut_580.mask = 64'he0e0e0e0e0e0e000;

	lut_sub lut_606 ({i_28_, i_17_, g72, g30}, g81);
	defparam lut_606.LUT_SIZE = 4;
	defparam lut_606.mask = 16'h1000;

	lut_sub lut_611 ({i_28_, g2, i_29_}, g82);
	defparam lut_611.LUT_SIZE = 3;
	defparam lut_611.mask = 8'h20;

	lut_sub lut_618 ({g30, g38, g82}, g83);
	defparam lut_618.LUT_SIZE = 3;
	defparam lut_618.mask = 8'h01;

	lut_sub lut_622 ({i_28_, i_30_, i_29_}, g84);
	defparam lut_622.LUT_SIZE = 3;
	defparam lut_622.mask = 8'h80;

	lut_sub lut_629 ({i_34_, g57, g33, g84}, g85);
	defparam lut_629.LUT_SIZE = 4;
	defparam lut_629.mask = 16'h0001;

	lut_sub lut_634 ({i_31_, g70}, g86);
	defparam lut_634.LUT_SIZE = 2;
	defparam lut_634.mask = 4'b0111;

	lut_sub lut_643 ({i_7_, g85, g82, g86}, g87);
	defparam lut_643.LUT_SIZE = 4;
	defparam lut_643.mask = 16'h2f00;

	lut_sub lut_651 ({i_28_, i_29_}, g88);
	defparam lut_651.LUT_SIZE = 2;
	defparam lut_651.mask = 4'b0100;

	lut_sub lut_656 ({i_32_, g88}, g89);
	defparam lut_656.LUT_SIZE = 2;
	defparam lut_656.mask = 4'b0100;

	lut_sub lut_660 ({i_16_, i_27_, i_23_}, g90);
	defparam lut_660.LUT_SIZE = 3;
	defparam lut_660.mask = 8'h7f;

	lut_sub lut_673 ({g2, i_32_, g84, g90}, g91);
	defparam lut_673.LUT_SIZE = 4;
	defparam lut_673.mask = 16'h0020;

	lut_sub lut_682 ({g14, g73, g74, g89, g91}, g92);
	defparam lut_682.LUT_SIZE = 5;
	defparam lut_682.mask = 32'h00550357;

	lut_sub lut_696 ({i_24_, i_23_, i_26_}, g93);
	defparam lut_696.LUT_SIZE = 3;
	defparam lut_696.mask = 8'h80;

	lut_sub lut_702 ({g19, g93, i_30_}, g94);
	defparam lut_702.LUT_SIZE = 3;
	defparam lut_702.mask = 8'h02;

	lut_sub lut_708 ({i_17_, i_21_, i_2_, g94, g28}, g95);
	defparam lut_708.LUT_SIZE = 5;
	defparam lut_708.mask = 32'h10000000;

	lut_sub lut_712 ({i_30_, i_31_}, g96);
	defparam lut_712.LUT_SIZE = 2;
	defparam lut_712.mask = 4'b1000;

	lut_sub lut_717 ({i_28_, i_29_, g96}, g97);
	defparam lut_717.LUT_SIZE = 3;
	defparam lut_717.mask = 8'h40;

	lut_sub lut_723 ({g33, g97}, g98);
	defparam lut_723.LUT_SIZE = 2;
	defparam lut_723.mask = 4'b0001;

	lut_sub lut_730 ({i_7_, i_32_, g95, g66, g98}, g99);
	defparam lut_730.LUT_SIZE = 5;
	defparam lut_730.mask = 32'h1f111111;

	lut_sub lut_746 ({g93, g34}, g100);
	defparam lut_746.LUT_SIZE = 2;
	defparam lut_746.mask = 4'b0001;

	lut_sub lut_751 ({g19, i_26_}, g101);
	defparam lut_751.LUT_SIZE = 2;
	defparam lut_751.mask = 4'b0010;

	lut_sub lut_758 ({i_21_, g33, g100, g101}, g102);
	defparam lut_758.LUT_SIZE = 4;
	defparam lut_758.mask = 16'hc8cc;

	lut_sub lut_771 ({i_32_, g4, g102, g41}, g103);
	defparam lut_771.LUT_SIZE = 4;
	defparam lut_771.mask = 16'h4500;

	lut_sub lut_782 ({g83, g87, g92, g99, g103}, g104);
	defparam lut_782.LUT_SIZE = 5;
	defparam lut_782.mask = 32'h80000000;

	lut_sub lut_789 ({g88, g7, g27}, g105);
	defparam lut_789.LUT_SIZE = 3;
	defparam lut_789.mask = 8'h01;

	lut_sub lut_796 ({i_17_, i_9_, g14, g72, g105}, g106);
	defparam lut_796.LUT_SIZE = 5;
	defparam lut_796.mask = 32'h01000000;

	lut_sub lut_801 ({i_23_, g54}, g107);
	defparam lut_801.LUT_SIZE = 2;
	defparam lut_801.mask = 4'b0100;

	lut_sub lut_806 ({i_27_, g71}, g108);
	defparam lut_806.LUT_SIZE = 2;
	defparam lut_806.mask = 4'b0111;

	lut_sub lut_816 ({i_23_, g28, g37, g77, g108}, g109);
	defparam lut_816.LUT_SIZE = 5;
	defparam lut_816.mask = 32'h00020000;

	lut_sub lut_824 ({g7, g54, g6, g9}, g110);
	defparam lut_824.LUT_SIZE = 4;
	defparam lut_824.mask = 16'h0004;

	lut_sub lut_830 ({i_27_, g93, g88}, g111);
	defparam lut_830.LUT_SIZE = 3;
	defparam lut_830.mask = 8'h10;

	lut_sub lut_836 ({i_3_, i_18_, g14, g12}, g112);
	defparam lut_836.LUT_SIZE = 4;
	defparam lut_836.mask = 16'h1131;

	lut_sub lut_847 ({g111, i_9_, g112, g53}, g113);
	defparam lut_847.LUT_SIZE = 4;
	defparam lut_847.mask = 16'h0010;

	lut_sub lut_856 ({i_21_, g28, g7, g9, g100, g113}, g114);
	defparam lut_856.LUT_SIZE = 6;
	defparam lut_856.mask = 64'h0055005700000003;

	lut_sub lut_876 ({g77, g76, g107, g109, g110, g114}, g115);
	defparam lut_876.LUT_SIZE = 6;
	defparam lut_876.mask = 64'h8080808080808000;

	lut_sub lut_891 ({g80, g81, g104, g106, g115}, g116);
	defparam lut_891.LUT_SIZE = 5;
	defparam lut_891.mask = 32'h00000400;

	lut_sub lut_900 ({g6, g18, g44, g64, g116}, g117);
	defparam lut_900.LUT_SIZE = 5;
	defparam lut_900.mask = 32'h40004040;

	lut_sub lut_906 ({i_35_, i_36_}, g118);
	defparam lut_906.LUT_SIZE = 2;
	defparam lut_906.mask = 4'b0100;

	lut_sub lut_911 ({i_32_, g118}, g119);
	defparam lut_911.LUT_SIZE = 2;
	defparam lut_911.mask = 4'b0100;

	lut_sub lut_919 ({g22, g108, g60, g58}, g120);
	defparam lut_919.LUT_SIZE = 4;
	defparam lut_919.mask = 16'h1000;

	lut_sub lut_924 ({i_28_, g71}, g121);
	defparam lut_924.LUT_SIZE = 2;
	defparam lut_924.mask = 4'b1000;

	lut_sub lut_930 ({i_34_, i_29_, g96, g121}, g122);
	defparam lut_930.LUT_SIZE = 4;
	defparam lut_930.mask = 16'h1000;

	lut_sub lut_939 ({g100, g56, g119, g120, g122}, g123);
	defparam lut_939.LUT_SIZE = 5;
	defparam lut_939.mask = 32'h0707070f;

	lut_sub lut_958 ({g95, i_31_, i_8_, g102, g61}, g124);
	defparam lut_958.LUT_SIZE = 5;
	defparam lut_958.mask = 32'h4400f400;

	lut_sub lut_971 ({i_16_, g22, g33, g9}, g125);
	defparam lut_971.LUT_SIZE = 4;
	defparam lut_971.mask = 16'h1000;

	lut_sub lut_978 ({i_34_, g57, g34, g125}, g126);
	defparam lut_978.LUT_SIZE = 4;
	defparam lut_978.mask = 16'h0001;

	lut_sub lut_987 ({g1, g108, g50, g124, g126}, g127);
	defparam lut_987.LUT_SIZE = 5;
	defparam lut_987.mask = 32'h88888088;

	lut_sub lut_997 ({i_7_, i_10_}, g128);
	defparam lut_997.LUT_SIZE = 2;
	defparam lut_997.mask = 4'b0001;

	lut_sub lut_1003 ({i_17_, i_12_, i_13_, g54, g128}, g129);
	defparam lut_1003.LUT_SIZE = 5;
	defparam lut_1003.mask = 32'h01010100;

	lut_sub lut_1010 ({i_27_, g88}, g130);
	defparam lut_1010.LUT_SIZE = 2;
	defparam lut_1010.mask = 4'b0100;

	lut_sub lut_1016 ({g33, g130, i_22_}, g131);
	defparam lut_1016.LUT_SIZE = 3;
	defparam lut_1016.mask = 8'h01;

	lut_sub lut_1021 ({i_33_, g57}, g132);
	defparam lut_1021.LUT_SIZE = 2;
	defparam lut_1021.mask = 4'b0001;

	lut_sub lut_1028 ({g33, g84, g132}, g133);
	defparam lut_1028.LUT_SIZE = 3;
	defparam lut_1028.mask = 8'h01;

	lut_sub lut_1033 ({i_17_, i_12_, g54}, g134);
	defparam lut_1033.LUT_SIZE = 3;
	defparam lut_1033.mask = 8'h54;

	lut_sub lut_1043 ({i_12_, g45, i_25_, g131, g133, g134}, g135);
	defparam lut_1043.LUT_SIZE = 6;
	defparam lut_1043.mask = 64'h05370f3f05370537;

	lut_sub lut_1078 ({i_28_, i_31_, i_29_, g5}, g136);
	defparam lut_1078.LUT_SIZE = 4;
	defparam lut_1078.mask = 16'h0800;

	lut_sub lut_1083 ({i_21_, i_30_, g33}, g137);
	defparam lut_1083.LUT_SIZE = 3;
	defparam lut_1083.mask = 8'h04;

	lut_sub lut_1090 ({i_28_, i_14_, g132, i_25_, g133, g137}, g138);
	defparam lut_1090.LUT_SIZE = 6;
	defparam lut_1090.mask = 64'h0005337700003333;

	lut_sub lut_1117 ({i_34_, g129, g135, g136, g138}, g139);
	defparam lut_1117.LUT_SIZE = 5;
	defparam lut_1117.mask = 32'h00005f7f;

	lut_sub lut_1133 ({i_24_, i_28_, i_26_, i_30_}, g140);
	defparam lut_1133.LUT_SIZE = 4;
	defparam lut_1133.mask = 16'h8000;

	lut_sub lut_1139 ({i_33_, i_28_, g2, g86}, g141);
	defparam lut_1139.LUT_SIZE = 4;
	defparam lut_1139.mask = 16'h0020;

	lut_sub lut_1146 ({i_34_, g132, g140, g141}, g142);
	defparam lut_1146.LUT_SIZE = 4;
	defparam lut_1146.mask = 16'ha8aa;

	lut_sub lut_1158 ({i_33_, g2, g1}, g143);
	defparam lut_1158.LUT_SIZE = 3;
	defparam lut_1158.mask = 8'h01;

	lut_sub lut_1165 ({i_34_, g71, g84, g132}, g144);
	defparam lut_1165.LUT_SIZE = 4;
	defparam lut_1165.mask = 16'h1000;

	lut_sub lut_1172 ({g86, g143, g144}, g145);
	defparam lut_1172.LUT_SIZE = 3;
	defparam lut_1172.mask = 8'h8a;

	lut_sub lut_1180 ({i_14_, i_21_, g142, i_25_, g145}, g146);
	defparam lut_1180.LUT_SIZE = 5;
	defparam lut_1180.mask = 32'h2232aafa;

	lut_sub lut_1200 ({g2, g86, i_22_}, g147);
	defparam lut_1200.LUT_SIZE = 3;
	defparam lut_1200.mask = 8'h04;

	lut_sub lut_1205 ({i_34_, i_35_, g71, i_30_, i_32_, i_31_}, g148);
	defparam lut_1205.LUT_SIZE = 6;
	defparam lut_1205.mask = 64'h8000808000000000;

	lut_sub lut_1214 ({i_21_, g88, i_20_, g147, g148}, g149);
	defparam lut_1214.LUT_SIZE = 5;
	defparam lut_1214.mask = 32'h00370033;

	lut_sub lut_1227 ({i_17_, i_12_, g45}, g150);
	defparam lut_1227.LUT_SIZE = 3;
	defparam lut_1227.mask = 8'h54;

	lut_sub lut_1237 ({g33, i_29_, g101, g55, i_22_, g150}, g151);
	defparam lut_1237.LUT_SIZE = 6;
	defparam lut_1237.mask = 64'h0000000000000013;

	lut_sub lut_1244 ({i_12_, g28}, g152);
	defparam lut_1244.LUT_SIZE = 2;
	defparam lut_1244.mask = 4'b0100;

	lut_sub lut_1250 ({i_21_, i_2_, g111, g152, i_20_}, g153);
	defparam lut_1250.LUT_SIZE = 5;
	defparam lut_1250.mask = 32'h00020000;

	lut_sub lut_1255 ({i_34_, i_23_, i_26_, g88, i_22_}, g154);
	defparam lut_1255.LUT_SIZE = 5;
	defparam lut_1255.mask = 32'h10101100;

	lut_sub lut_1265 ({i_24_, i_30_, g57, g153, g154}, g155);
	defparam lut_1265.LUT_SIZE = 5;
	defparam lut_1265.mask = 32'hc8cccccc;

	lut_sub lut_1287 ({i_34_, g53, g131, g151, g155}, g156);
	defparam lut_1287.LUT_SIZE = 5;
	defparam lut_1287.mask = 32'h44444440;

	lut_sub lut_1298 ({i_17_, i_12_, g28}, g157);
	defparam lut_1298.LUT_SIZE = 3;
	defparam lut_1298.mask = 8'h54;

	lut_sub lut_1306 ({i_16_, i_12_, i_13_, i_14_, g90, g38}, g158);
	defparam lut_1306.LUT_SIZE = 6;
	defparam lut_1306.mask = 64'h0c0004000c000000;

	lut_sub lut_1314 ({i_21_, i_22_, i_20_}, g159);
	defparam lut_1314.LUT_SIZE = 3;
	defparam lut_1314.mask = 8'h40;

	lut_sub lut_1323 ({g111, g143, g157, g158, g159}, g160);
	defparam lut_1323.LUT_SIZE = 5;
	defparam lut_1323.mask = 32'h00330537;

	lut_sub lut_1340 ({i_16_, i_36_, g33, g70, g73}, g161);
	defparam lut_1340.LUT_SIZE = 5;
	defparam lut_1340.mask = 32'h00040000;

	lut_sub lut_1346 ({g33, i_8_, g157}, g162);
	defparam lut_1346.LUT_SIZE = 3;
	defparam lut_1346.mask = 8'h04;

	lut_sub lut_1355 ({i_34_, g96, g34, g161, g118, g162}, g163);
	defparam lut_1355.LUT_SIZE = 6;
	defparam lut_1355.mask = 64'h00000000000f001f;

	lut_sub lut_1367 ({i_33_, i_25_}, g164);
	defparam lut_1367.LUT_SIZE = 2;
	defparam lut_1367.mask = 4'b0001;

	lut_sub lut_1373 ({g134, g164}, g165);
	defparam lut_1373.LUT_SIZE = 2;
	defparam lut_1373.mask = 4'b0001;

	lut_sub lut_1379 ({i_27_, i_28_, i_31_, g129, g165}, g166);
	defparam lut_1379.LUT_SIZE = 5;
	defparam lut_1379.mask = 32'h57000000;

	lut_sub lut_1387 ({i_24_, i_34_, i_35_, i_23_, i_21_}, g167);
	defparam lut_1387.LUT_SIZE = 5;
	defparam lut_1387.mask = 32'h04440400;

	lut_sub lut_1396 ({i_27_, i_28_, g93, i_31_, g4}, g168);
	defparam lut_1396.LUT_SIZE = 5;
	defparam lut_1396.mask = 32'h13111111;

	lut_sub lut_1408 ({i_16_, i_33_, i_17_, i_12_, i_13_, i_14_}, g169);
	defparam lut_1408.LUT_SIZE = 6;
	defparam lut_1408.mask = 64'h0000444000000000;

	lut_sub lut_1415 ({g20, i_34_, i_35_, i_21_}, g170);
	defparam lut_1415.LUT_SIZE = 4;
	defparam lut_1415.mask = 16'h1015;

	lut_sub lut_1427 ({g3, g168, g129, g169, g170}, g171);
	defparam lut_1427.LUT_SIZE = 5;
	defparam lut_1427.mask = 32'h000f111f;

	lut_sub lut_1446 ({g160, g163, g166, g167, g171}, g172);
	defparam lut_1446.LUT_SIZE = 5;
	defparam lut_1446.mask = 32'ha8000000;

	lut_sub lut_1453 ({i_3_, i_18_, i_4_, i_5_, g31}, g173);
	defparam lut_1453.LUT_SIZE = 5;
	defparam lut_1453.mask = 32'h00004000;

	lut_sub lut_1459 ({i_7_, i_9_, g14, g12}, g174);
	defparam lut_1459.LUT_SIZE = 4;
	defparam lut_1459.mask = 16'h1000;

	lut_sub lut_1466 ({i_36_, g89, g173, g174}, g175);
	defparam lut_1466.LUT_SIZE = 4;
	defparam lut_1466.mask = 16'h0007;

	lut_sub lut_1474 ({i_2_, g14, i_8_, g118}, g176);
	defparam lut_1474.LUT_SIZE = 4;
	defparam lut_1474.mask = 16'hfb00;

	lut_sub lut_1487 ({g88, i_9_, g12, g176}, g177);
	defparam lut_1487.LUT_SIZE = 4;
	defparam lut_1487.mask = 16'h0020;

	lut_sub lut_1493 ({i_4_, i_5_, g48, g118}, g178);
	defparam lut_1493.LUT_SIZE = 4;
	defparam lut_1493.mask = 16'h1000;

	lut_sub lut_1499 ({i_2_, g88, i_9_, i_3_, i_18_, g178}, g179);
	defparam lut_1499.LUT_SIZE = 6;
	defparam lut_1499.mask = 64'h0000040400000c04;

	lut_sub lut_1512 ({g53, g72, g175, g177, g179}, g180);
	defparam lut_1512.LUT_SIZE = 5;
	defparam lut_1512.mask = 32'h0000007f;

	lut_sub lut_1522 ({i_24_, i_34_, i_35_, i_26_}, g181);
	defparam lut_1522.LUT_SIZE = 4;
	defparam lut_1522.mask = 16'h40cf;

	lut_sub lut_1534 ({i_27_, i_36_, g84, g181}, g182);
	defparam lut_1534.LUT_SIZE = 4;
	defparam lut_1534.mask = 16'h0200;

	lut_sub lut_1540 ({i_23_, i_7_, i_8_, g152, g182}, g183);
	defparam lut_1540.LUT_SIZE = 5;
	defparam lut_1540.mask = 32'h10330000;

	lut_sub lut_1551 ({i_7_, i_9_, g712, g180, g183}, g184);
	defparam lut_1551.LUT_SIZE = 5;
	defparam lut_1551.mask = 32'h88888ccc;

	lut_sub lut_1570 ({g146, g149, g156, g172, g184}, g185);
	defparam lut_1570.LUT_SIZE = 5;
	defparam lut_1570.mask = 32'h01000000;

	lut_sub lut_1579 ({g118, g123, g127, g139, g185}, g186);
	defparam lut_1579.LUT_SIZE = 5;
	defparam lut_1579.mask = 32'h44000400;

	lut_sub lut_1589 ({g27, g30, g49, g118}, g187);
	defparam lut_1589.LUT_SIZE = 4;
	defparam lut_1589.mask = 16'hf0e0;

	lut_sub lut_1600 ({i_17_, i_36_, g33}, g188);
	defparam lut_1600.LUT_SIZE = 3;
	defparam lut_1600.mask = 8'h10;

	lut_sub lut_1608 ({i_29_, g69, g119, g187, g188}, g189);
	defparam lut_1608.LUT_SIZE = 5;
	defparam lut_1608.mask = 32'h444f0000;

	lut_sub lut_1620 ({i_3_, g14, g15}, g190);
	defparam lut_1620.LUT_SIZE = 3;
	defparam lut_1620.mask = 8'h01;

	lut_sub lut_1624 ({i_16_, i_17_, i_13_, i_14_, i_10_}, g191);
	defparam lut_1624.LUT_SIZE = 5;
	defparam lut_1624.mask = 32'hac000000;

	lut_sub lut_1634 ({i_31_, g14, g119, g152}, g192);
	defparam lut_1634.LUT_SIZE = 4;
	defparam lut_1634.mask = 16'h0100;

	lut_sub lut_1639 ({i_36_, i_7_, i_32_, g14}, g193);
	defparam lut_1639.LUT_SIZE = 4;
	defparam lut_1639.mask = 16'h0040;

	lut_sub lut_1647 ({i_9_, g14, g45, g13, g119}, g194);
	defparam lut_1647.LUT_SIZE = 5;
	defparam lut_1647.mask = 32'h00010000;

	lut_sub lut_1656 ({i_9_, g176, g191, g192, g193, g194}, g195);
	defparam lut_1656.LUT_SIZE = 6;
	defparam lut_1656.mask = 64'ha000a080a0a0a0a0;

	lut_sub lut_1676 ({i_29_, g45, g119, g190, g195}, g196);
	defparam lut_1676.LUT_SIZE = 5;
	defparam lut_1676.mask = 32'h0000aaab;

	lut_sub lut_1689 ({i_30_, g7}, g197);
	defparam lut_1689.LUT_SIZE = 2;
	defparam lut_1689.mask = 4'b0100;

	lut_sub lut_1695 ({i_17_, i_36_, i_2_, g28, g197}, g198);
	defparam lut_1695.LUT_SIZE = 5;
	defparam lut_1695.mask = 32'h00100000;

	lut_sub lut_1703 ({g86, g118, g152, g198}, g199);
	defparam lut_1703.LUT_SIZE = 4;
	defparam lut_1703.mask = 16'ha8aa;

	lut_sub lut_1717 ({i_21_, g33, g189, g196, g199}, g200);
	defparam lut_1717.LUT_SIZE = 5;
	defparam lut_1717.mask = 32'hf040f0f0;

	lut_sub lut_1737 ({g57, i_29_, g96, g125, g162}, g201);
	defparam lut_1737.LUT_SIZE = 5;
	defparam lut_1737.mask = 32'h05003700;

	lut_sub lut_1749 ({i_12_, g33, i_29_, g54, i_22_}, g202);
	defparam lut_1749.LUT_SIZE = 5;
	defparam lut_1749.mask = 32'h00010000;

	lut_sub lut_1757 ({i_29_, g161, g118, g201, g202}, g203);
	defparam lut_1757.LUT_SIZE = 5;
	defparam lut_1757.mask = 32'ha800a8a8;

	lut_sub lut_1771 ({g2, i_21_, g130, i_22_, i_20_}, g204);
	defparam lut_1771.LUT_SIZE = 5;
	defparam lut_1771.mask = 32'h00000703;

	lut_sub lut_1781 ({i_24_, i_27_, i_28_, i_29_, g86, g157}, g205);
	defparam lut_1781.LUT_SIZE = 6;
	defparam lut_1781.mask = 64'h0d000c0000000000;

	lut_sub lut_1790 ({i_34_, i_21_, i_20_, g205}, g206);
	defparam lut_1790.LUT_SIZE = 4;
	defparam lut_1790.mask = 16'h0010;

	lut_sub lut_1796 ({i_34_, g34, g101}, g207);
	defparam lut_1796.LUT_SIZE = 3;
	defparam lut_1796.mask = 8'ha8;

	lut_sub lut_1802 ({i_33_, i_24_, i_13_, i_14_, i_25_}, g208);
	defparam lut_1802.LUT_SIZE = 5;
	defparam lut_1802.mask = 32'h00007400;

	lut_sub lut_1811 ({i_16_, i_17_, i_12_, g207, g208}, g209);
	defparam lut_1811.LUT_SIZE = 5;
	defparam lut_1811.mask = 32'h44400000;

	lut_sub lut_1818 ({i_3_, i_18_, i_11_, i_19_, g128}, g210);
	defparam lut_1818.LUT_SIZE = 5;
	defparam lut_1818.mask = 32'h40405540;

	lut_sub lut_1829 ({i_27_, i_28_, g2, i_31_, i_29_}, g211);
	defparam lut_1829.LUT_SIZE = 5;
	defparam lut_1829.mask = 32'h02000000;

	lut_sub lut_1837 ({g150, g209, g210, g211}, g212);
	defparam lut_1837.LUT_SIZE = 4;
	defparam lut_1837.mask = 16'hf0e0;

	lut_sub lut_1852 ({g28, g108, g60, g51, g118}, g213);
	defparam lut_1852.LUT_SIZE = 5;
	defparam lut_1852.mask = 32'h00000100;

	lut_sub lut_1860 ({i_27_, g2, g1, g165, g213}, g214);
	defparam lut_1860.LUT_SIZE = 5;
	defparam lut_1860.mask = 32'haaa8aaaa;

	lut_sub lut_1883 ({g157, g204, g206, g212, g214}, g215);
	defparam lut_1883.LUT_SIZE = 5;
	defparam lut_1883.mask = 32'h10101000;

	lut_sub lut_1893 ({i_23_, g101, g200, g203, g215}, g216);
	defparam lut_1893.LUT_SIZE = 5;
	defparam lut_1893.mask = 32'h5501ff03;

	lut_sub lut_1914 ({g2, i_32_, g84, g38}, g217);
	defparam lut_1914.LUT_SIZE = 4;
	defparam lut_1914.mask = 16'h0010;

	lut_sub lut_1921 ({i_17_, g33, i_29_, g70, g101}, g218);
	defparam lut_1921.LUT_SIZE = 5;
	defparam lut_1921.mask = 32'h00400000;

	lut_sub lut_1929 ({i_34_, g70, g35, g217, g218}, g219);
	defparam lut_1929.LUT_SIZE = 5;
	defparam lut_1929.mask = 32'h88888088;

	lut_sub lut_1942 ({g19, i_30_, g130, g14}, g220);
	defparam lut_1942.LUT_SIZE = 4;
	defparam lut_1942.mask = 16'h11f1;

	lut_sub lut_1953 ({i_12_, i_7_, i_9_, g702}, g221);
	defparam lut_1953.LUT_SIZE = 4;
	defparam lut_1953.mask = 16'h0400;

	lut_sub lut_1959 ({i_12_, i_21_, i_36_, g93, g7}, g222);
	defparam lut_1959.LUT_SIZE = 5;
	defparam lut_1959.mask = 32'h01000000;

	lut_sub lut_1964 ({i_28_, g96}, g223);
	defparam lut_1964.LUT_SIZE = 2;
	defparam lut_1964.mask = 4'b0100;

	lut_sub lut_1971 ({i_2_, g88, g119, i_0_, g223}, g224);
	defparam lut_1971.LUT_SIZE = 5;
	defparam lut_1971.mask = 32'h05370033;

	lut_sub lut_1988 ({g7, g23, g182}, g225);
	defparam lut_1988.LUT_SIZE = 3;
	defparam lut_1988.mask = 8'h01;

	lut_sub lut_1993 ({i_12_, g88, i_0_}, g226);
	defparam lut_1993.LUT_SIZE = 3;
	defparam lut_1993.mask = 8'h10;

	lut_sub lut_2001 ({i_17_, g72, g224, g225, g226}, g227);
	defparam lut_2001.LUT_SIZE = 5;
	defparam lut_2001.mask = 32'hcc80cc88;

	lut_sub lut_2019 ({g220, g221, g222, g227}, g228);
	defparam lut_2019.LUT_SIZE = 4;
	defparam lut_2019.mask = 16'h5040;

	lut_sub lut_2027 ({i_16_, i_36_, i_7_, g219, g228}, g229);
	defparam lut_2027.LUT_SIZE = 5;
	defparam lut_2027.mask = 32'haaea0000;

	lut_sub lut_2040 ({i_16_, i_17_, g702}, g230);
	defparam lut_2040.LUT_SIZE = 3;
	defparam lut_2040.mask = 8'h40;

	lut_sub lut_2047 ({i_7_, i_9_, g23, g230, g712}, g231);
	defparam lut_2047.LUT_SIZE = 5;
	defparam lut_2047.mask = 32'h00003b00;

	lut_sub lut_2056 ({i_28_, i_12_, i_30_, i_31_, i_29_, g14}, g232);
	defparam lut_2056.LUT_SIZE = 6;
	defparam lut_2056.mask = 64'hf010000000000000;

	lut_sub lut_2067 ({i_23_, i_8_, g108, g118, g232}, g233);
	defparam lut_2067.LUT_SIZE = 5;
	defparam lut_2067.mask = 32'h10000000;

	lut_sub lut_2074 ({g111, i_9_, g14, g24}, g234);
	defparam lut_2074.LUT_SIZE = 4;
	defparam lut_2074.mask = 16'h0020;

	lut_sub lut_2080 ({g19, g93, i_31_}, g235);
	defparam lut_2080.LUT_SIZE = 3;
	defparam lut_2080.mask = 8'h02;

	lut_sub lut_2088 ({i_17_, g29, g119, g234, g235}, g236);
	defparam lut_2088.LUT_SIZE = 5;
	defparam lut_2088.mask = 32'h03070000;

	lut_sub lut_2098 ({i_16_, i_21_, g233, g236}, g237);
	defparam lut_2098.LUT_SIZE = 4;
	defparam lut_2098.mask = 16'h7000;

	lut_sub lut_2105 ({i_3_, i_18_, i_11_, i_19_, g128}, g238);
	defparam lut_2105.LUT_SIZE = 5;
	defparam lut_2105.mask = 32'hcc40dd40;

	lut_sub lut_2122 ({i_31_, g33, i_18_, i_19_, g207}, g239);
	defparam lut_2122.LUT_SIZE = 5;
	defparam lut_2122.mask = 32'h000000a8;

	lut_sub lut_2129 ({i_24_, i_34_, i_35_, g3, i_21_, i_31_}, g240);
	defparam lut_2129.LUT_SIZE = 6;
	defparam lut_2129.mask = 64'h0001010100010000;

	lut_sub lut_2137 ({i_3_, i_11_, g128}, g241);
	defparam lut_2137.LUT_SIZE = 3;
	defparam lut_2137.mask = 8'h04;

	lut_sub lut_2146 ({g33, g238, g239, g240, g241}, g242);
	defparam lut_2146.LUT_SIZE = 5;
	defparam lut_2146.mask = 32'h0537053f;

	lut_sub lut_2164 ({i_16_, i_17_, i_12_, i_13_}, g243);
	defparam lut_2164.LUT_SIZE = 4;
	defparam lut_2164.mask = 16'ha800;

	lut_sub lut_2173 ({i_3_, i_11_, g128, g242, g243}, g244);
	defparam lut_2173.LUT_SIZE = 5;
	defparam lut_2173.mask = 32'h01000101;

	lut_sub lut_2184 ({g22, g229, g231, g237, g244}, g245);
	defparam lut_2184.LUT_SIZE = 5;
	defparam lut_2184.mask = 32'h8000aaff;

	lut_sub lut_2204 ({i_36_, g117, g186, g216, g245}, o_0_);
	defparam lut_2204.LUT_SIZE = 5;
	defparam lut_2204.mask = 32'hfefefffe;

	lut_sub lut_2239 ({i_23_, g45, g50, g51}, g247);
	defparam lut_2239.LUT_SIZE = 4;
	defparam lut_2239.mask = 16'hc8cc;

	lut_sub lut_2249 ({i_4_, i_5_, i_0_}, g248);
	defparam lut_2249.LUT_SIZE = 3;
	defparam lut_2249.mask = 8'h80;

	lut_sub lut_2255 ({g54, g24}, g249);
	defparam lut_2255.LUT_SIZE = 2;
	defparam lut_2255.mask = 4'b0010;

	lut_sub lut_2261 ({i_33_, g45, i_10_, g249}, g250);
	defparam lut_2261.LUT_SIZE = 4;
	defparam lut_2261.mask = 16'ha2aa;

	lut_sub lut_2271 ({i_17_, i_23_, i_20_, i_37_}, g251);
	defparam lut_2271.LUT_SIZE = 4;
	defparam lut_2271.mask = 16'h4000;

	lut_sub lut_2280 ({g31, g89, g248, g250, g251}, g252);
	defparam lut_2280.LUT_SIZE = 5;
	defparam lut_2280.mask = 32'h00000004;

	lut_sub lut_2285 ({i_17_, i_23_, g88, i_20_}, g253);
	defparam lut_2285.LUT_SIZE = 4;
	defparam lut_2285.mask = 16'h2000;

	lut_sub lut_2289 ({i_35_, i_37_}, g254);
	defparam lut_2289.LUT_SIZE = 2;
	defparam lut_2289.mask = 4'b0100;

	lut_sub lut_2295 ({i_33_, g45, i_10_, g254}, g255);
	defparam lut_2295.LUT_SIZE = 4;
	defparam lut_2295.mask = 16'h0400;

	lut_sub lut_2304 ({g48, g254, g249, g248, g255}, g256);
	defparam lut_2304.LUT_SIZE = 5;
	defparam lut_2304.mask = 32'h00000013;

	lut_sub lut_2313 ({i_2_, g28, g253, g256}, g257);
	defparam lut_2313.LUT_SIZE = 4;
	defparam lut_2313.mask = 16'h1113;

	lut_sub lut_2323 ({i_23_, i_21_, g88, i_22_, g157}, g258);
	defparam lut_2323.LUT_SIZE = 5;
	defparam lut_2323.mask = 32'h00040000;

	lut_sub lut_2328 ({i_33_, i_13_, i_14_, g254}, g259);
	defparam lut_2328.LUT_SIZE = 4;
	defparam lut_2328.mask = 16'h5444;

	lut_sub lut_2337 ({i_16_, i_23_, i_20_, g259}, g260);
	defparam lut_2337.LUT_SIZE = 4;
	defparam lut_2337.mask = 16'h4000;

	lut_sub lut_2341 ({i_17_, i_12_, i_23_, i_20_, i_0_}, g261);
	defparam lut_2341.LUT_SIZE = 5;
	defparam lut_2341.mask = 32'haa80aa00;

	lut_sub lut_2357 ({i_28_, g70, g258, g260, g261}, g262);
	defparam lut_2357.LUT_SIZE = 5;
	defparam lut_2357.mask = 32'he0f0f0f0;

	lut_sub lut_2376 ({g14, i_1_, i_0_}, g263);
	defparam lut_2376.LUT_SIZE = 3;
	defparam lut_2376.mask = 8'h08;

	lut_sub lut_2382 ({i_7_, i_8_, i_37_, g263, g253}, g264);
	defparam lut_2382.LUT_SIZE = 5;
	defparam lut_2382.mask = 32'h01000000;

	lut_sub lut_2389 ({i_33_, g45, g54, g264}, g265);
	defparam lut_2389.LUT_SIZE = 4;
	defparam lut_2389.mask = 16'h1511;

	lut_sub lut_2400 ({i_33_, i_13_, i_14_, g37, g58, g254}, g266);
	defparam lut_2400.LUT_SIZE = 6;
	defparam lut_2400.mask = 64'h0101010001000100;

	lut_sub lut_2411 ({i_33_, i_17_, g28, g54, g254}, g267);
	defparam lut_2411.LUT_SIZE = 5;
	defparam lut_2411.mask = 32'h05000100;

	lut_sub lut_2419 ({i_23_, i_9_, g89, i_20_, g267}, g268);
	defparam lut_2419.LUT_SIZE = 5;
	defparam lut_2419.mask = 32'h04000000;

	lut_sub lut_2424 ({i_3_, i_18_, g14, i_0_}, g269);
	defparam lut_2424.LUT_SIZE = 4;
	defparam lut_2424.mask = 16'h0020;

	lut_sub lut_2432 ({i_6_, g12, g248, g268, g269}, g270);
	defparam lut_2432.LUT_SIZE = 5;
	defparam lut_2432.mask = 32'h11131111;

	lut_sub lut_2449 ({g257, g262, g265, g266, g270}, g271);
	defparam lut_2449.LUT_SIZE = 5;
	defparam lut_2449.mask = 32'h00800000;

	lut_sub lut_2455 ({i_33_, g1, g254}, g272);
	defparam lut_2455.LUT_SIZE = 3;
	defparam lut_2455.mask = 8'h10;

	lut_sub lut_2464 ({g13, g107, g47, g49, g51}, g273);
	defparam lut_2464.LUT_SIZE = 5;
	defparam lut_2464.mask = 32'h005f007f;

	lut_sub lut_2482 ({i_12_, i_6_, g248, g260}, g274);
	defparam lut_2482.LUT_SIZE = 4;
	defparam lut_2482.mask = 16'h1000;

	lut_sub lut_2491 ({g1, g89, g254, g273, g274}, g275);
	defparam lut_2491.LUT_SIZE = 5;
	defparam lut_2491.mask = 32'h00550357;

	lut_sub lut_2510 ({g247, g252, g271, g272, g275}, g276);
	defparam lut_2510.LUT_SIZE = 5;
	defparam lut_2510.mask = 32'h08000a00;

	lut_sub lut_2516 ({i_33_, i_34_, i_32_}, g277);
	defparam lut_2516.LUT_SIZE = 3;
	defparam lut_2516.mask = 8'h20;

	lut_sub lut_2523 ({i_16_, i_13_, g33, g9, g69}, g278);
	defparam lut_2523.LUT_SIZE = 5;
	defparam lut_2523.mask = 32'ha8aaaaaa;

	lut_sub lut_2542 ({i_33_, g2, i_37_}, g279);
	defparam lut_2542.LUT_SIZE = 3;
	defparam lut_2542.mask = 8'h10;

	lut_sub lut_2547 ({i_16_, i_17_, i_12_, i_13_, i_23_, g7}, g280);
	defparam lut_2547.LUT_SIZE = 6;
	defparam lut_2547.mask = 64'h4040400000000000;

	lut_sub lut_2554 ({i_16_, i_34_, i_12_, i_13_, g33}, g281);
	defparam lut_2554.LUT_SIZE = 5;
	defparam lut_2554.mask = 32'h00400000;

	lut_sub lut_2560 ({i_33_, i_8_, g254, g281}, g282);
	defparam lut_2560.LUT_SIZE = 4;
	defparam lut_2560.mask = 16'h1000;

	lut_sub lut_2567 ({i_30_, g279, g280, g282}, g283);
	defparam lut_2567.LUT_SIZE = 4;
	defparam lut_2567.mask = 16'h5700;

	lut_sub lut_2578 ({g93, g53, g10, i_10_, i_37_}, g284);
	defparam lut_2578.LUT_SIZE = 5;
	defparam lut_2578.mask = 32'h00000004;

	lut_sub lut_2584 ({i_13_, i_10_, g11, g23}, g285);
	defparam lut_2584.LUT_SIZE = 4;
	defparam lut_2584.mask = 16'h1000;

	lut_sub lut_2588 ({i_33_, i_32_, i_37_}, g286);
	defparam lut_2588.LUT_SIZE = 3;
	defparam lut_2588.mask = 8'h40;

	lut_sub lut_2595 ({g93, i_30_, i_31_, g150, g286}, g287);
	defparam lut_2595.LUT_SIZE = 5;
	defparam lut_2595.mask = 32'h00000100;

	lut_sub lut_2602 ({i_33_, g93, g55, g254}, g288);
	defparam lut_2602.LUT_SIZE = 4;
	defparam lut_2602.mask = 16'h0501;

	lut_sub lut_2613 ({g61, g279, g285, g287, g288}, g289);
	defparam lut_2613.LUT_SIZE = 5;
	defparam lut_2613.mask = 32'hccc08880;

	lut_sub lut_2629 ({i_33_, g65, g283, g284, g289}, g290);
	defparam lut_2629.LUT_SIZE = 5;
	defparam lut_2629.mask = 32'h50405050;

	lut_sub lut_2641 ({i_32_, g79, g279}, g291);
	defparam lut_2641.LUT_SIZE = 3;
	defparam lut_2641.mask = 8'h10;

	lut_sub lut_2650 ({g254, g277, g278, g290, g291}, g292);
	defparam lut_2650.LUT_SIZE = 5;
	defparam lut_2650.mask = 32'h22222202;

	lut_sub lut_2664 ({i_27_, g71, g1, g276, g292}, g293);
	defparam lut_2664.LUT_SIZE = 5;
	defparam lut_2664.mask = 32'hce0a0000;

	lut_sub lut_2675 ({i_7_, g29}, g294);
	defparam lut_2675.LUT_SIZE = 2;
	defparam lut_2675.mask = 4'b0100;

	lut_sub lut_2681 ({g32, g249}, g295);
	defparam lut_2681.LUT_SIZE = 2;
	defparam lut_2681.mask = 4'b0001;

	lut_sub lut_2687 ({g45, i_8_, g294}, g296);
	defparam lut_2687.LUT_SIZE = 3;
	defparam lut_2687.mask = 8'h04;

	lut_sub lut_2693 ({i_33_, g2, i_32_, g1, i_37_}, g297);
	defparam lut_2693.LUT_SIZE = 5;
	defparam lut_2693.mask = 32'h00110010;

	lut_sub lut_2703 ({i_33_, g37, g295, g296, g297}, g298);
	defparam lut_2703.LUT_SIZE = 5;
	defparam lut_2703.mask = 32'h11150105;

	lut_sub lut_2717 ({g2, g1, g54, i_37_}, g299);
	defparam lut_2717.LUT_SIZE = 4;
	defparam lut_2717.mask = 16'h0001;

	lut_sub lut_2725 ({i_8_, g294, g38, g298, g299}, g300);
	defparam lut_2725.LUT_SIZE = 5;
	defparam lut_2725.mask = 32'h03070303;

	lut_sub lut_2739 ({i_33_, i_17_, g45, i_8_, g294}, g301);
	defparam lut_2739.LUT_SIZE = 5;
	defparam lut_2739.mask = 32'h05040000;

	lut_sub lut_2750 ({g53, g42, g35, g296, g301}, g302);
	defparam lut_2750.LUT_SIZE = 5;
	defparam lut_2750.mask = 32'h01050155;

	lut_sub lut_2765 ({i_8_, g294, g42, g55, g35}, g303);
	defparam lut_2765.LUT_SIZE = 5;
	defparam lut_2765.mask = 32'h00130003;

	lut_sub lut_2776 ({i_33_, i_7_, g57, g33, g84}, g304);
	defparam lut_2776.LUT_SIZE = 5;
	defparam lut_2776.mask = 32'h01000000;

	lut_sub lut_2783 ({i_33_, i_30_, g21, g304, g280}, g305);
	defparam lut_2783.LUT_SIZE = 5;
	defparam lut_2783.mask = 32'hc8cccccc;

	lut_sub lut_2804 ({i_34_, i_37_, g302, g303, g305}, g306);
	defparam lut_2804.LUT_SIZE = 5;
	defparam lut_2804.mask = 32'h000000bf;

	lut_sub lut_2816 ({g142, i_25_, g144, i_20_}, g307);
	defparam lut_2816.LUT_SIZE = 4;
	defparam lut_2816.mask = 16'h0703;

	lut_sub lut_2826 ({i_13_, g10, i_10_, g55}, g308);
	defparam lut_2826.LUT_SIZE = 4;
	defparam lut_2826.mask = 16'h0405;

	lut_sub lut_2837 ({i_34_, g42, g21, g254, g308, g273}, g309);
	defparam lut_2837.LUT_SIZE = 6;
	defparam lut_2837.mask = 64'h0000000000050307;

	lut_sub lut_2848 ({i_24_, i_34_, i_35_, g34, i_37_}, g310);
	defparam lut_2848.LUT_SIZE = 5;
	defparam lut_2848.mask = 32'h01110100;

	lut_sub lut_2858 ({i_34_, i_29_, g34, g101, g254}, g311);
	defparam lut_2858.LUT_SIZE = 5;
	defparam lut_2858.mask = 32'h11001505;

	lut_sub lut_2869 ({i_16_, i_17_, i_12_, i_14_, g33, i_8_}, g312);
	defparam lut_2869.LUT_SIZE = 6;
	defparam lut_2869.mask = 64'h2020200000000000;

	lut_sub lut_2877 ({i_12_, g7, g107}, g313);
	defparam lut_2877.LUT_SIZE = 3;
	defparam lut_2877.mask = 8'h10;

	lut_sub lut_2885 ({i_30_, g310, g311, g312, g313}, g314);
	defparam lut_2885.LUT_SIZE = 5;
	defparam lut_2885.mask = 32'h03570000;

	lut_sub lut_2897 ({i_32_, i_29_, g101, g254}, g315);
	defparam lut_2897.LUT_SIZE = 4;
	defparam lut_2897.mask = 16'h1000;

	lut_sub lut_2904 ({g66, g34, i_37_, g315}, g316);
	defparam lut_2904.LUT_SIZE = 4;
	defparam lut_2904.mask = 16'haaa8;

	lut_sub lut_2916 ({i_16_, i_14_, g33, g9}, g317);
	defparam lut_2916.LUT_SIZE = 4;
	defparam lut_2916.mask = 16'h1000;

	lut_sub lut_2925 ({g68, g55, g314, g316, g317}, g318);
	defparam lut_2925.LUT_SIZE = 5;
	defparam lut_2925.mask = 32'hb0b0b030;

	lut_sub lut_2944 ({g300, g306, g307, g309, g318}, g319);
	defparam lut_2944.LUT_SIZE = 5;
	defparam lut_2944.mask = 32'h40000000;

	lut_sub lut_2950 ({i_33_, i_17_, i_12_, g45, g54}, g320);
	defparam lut_2950.LUT_SIZE = 5;
	defparam lut_2950.mask = 32'h77705550;

	lut_sub lut_2971 ({i_31_, g84, g5, g320}, g321);
	defparam lut_2971.LUT_SIZE = 4;
	defparam lut_2971.mask = 16'h0004;

	lut_sub lut_2978 ({i_34_, g35, g295, g321}, g322);
	defparam lut_2978.LUT_SIZE = 4;
	defparam lut_2978.mask = 16'h0057;

	lut_sub lut_2986 ({i_16_, i_17_, i_20_}, g323);
	defparam lut_2986.LUT_SIZE = 3;
	defparam lut_2986.mask = 8'h80;

	lut_sub lut_2992 ({g19, i_14_, i_7_, i_0_, g323}, g324);
	defparam lut_2992.LUT_SIZE = 5;
	defparam lut_2992.mask = 32'h00004000;

	lut_sub lut_2999 ({i_31_, g34, g134, g324}, g325);
	defparam lut_2999.LUT_SIZE = 4;
	defparam lut_2999.mask = 16'haaa8;

	lut_sub lut_3013 ({g111, g13, g31, i_20_, g248}, g326);
	defparam lut_3013.LUT_SIZE = 5;
	defparam lut_3013.mask = 32'h00000004;

	lut_sub lut_3019 ({g111, g190, i_20_}, g327);
	defparam lut_3019.LUT_SIZE = 3;
	defparam lut_3019.mask = 8'h02;

	lut_sub lut_3024 ({i_7_, i_0_, g327}, g328);
	defparam lut_3024.LUT_SIZE = 3;
	defparam lut_3024.mask = 8'h40;

	lut_sub lut_3030 ({i_12_, i_7_, g130, i_6_, g248}, g329);
	defparam lut_3030.LUT_SIZE = 5;
	defparam lut_3030.mask = 32'h04000000;

	lut_sub lut_3035 ({g19, i_12_, i_30_, i_7_, i_0_}, g330);
	defparam lut_3035.LUT_SIZE = 5;
	defparam lut_3035.mask = 32'h00008000;

	lut_sub lut_3042 ({g93, i_20_, g329, g330}, g331);
	defparam lut_3042.LUT_SIZE = 4;
	defparam lut_3042.mask = 16'h0070;

	lut_sub lut_3052 ({g54, g326, g328, g331}, g332);
	defparam lut_3052.LUT_SIZE = 4;
	defparam lut_3052.mask = 16'h007f;

	lut_sub lut_3065 ({g93, i_30_, g325, g332}, g333);
	defparam lut_3065.LUT_SIZE = 4;
	defparam lut_3065.mask = 16'haa2a;

	lut_sub lut_3075 ({i_29_, i_20_}, g334);
	defparam lut_3075.LUT_SIZE = 2;
	defparam lut_3075.mask = 4'b0010;

	lut_sub lut_3079 ({i_9_, i_6_}, g335);
	defparam lut_3079.LUT_SIZE = 2;
	defparam lut_3079.mask = 4'b1000;

	lut_sub lut_3085 ({g335, i_10_, g248}, g336);
	defparam lut_3085.LUT_SIZE = 3;
	defparam lut_3085.mask = 8'h04;

	lut_sub lut_3092 ({i_33_, g53, g254, g336}, g337);
	defparam lut_3092.LUT_SIZE = 4;
	defparam lut_3092.mask = 16'h0100;

	lut_sub lut_3100 ({g335, g24, g254, g248}, g338);
	defparam lut_3100.LUT_SIZE = 4;
	defparam lut_3100.mask = 16'h0010;

	lut_sub lut_3106 ({i_7_, i_37_, g263, g338}, g339);
	defparam lut_3106.LUT_SIZE = 4;
	defparam lut_3106.mask = 16'ha8aa;

	lut_sub lut_3122 ({g33, g101, g55, g334, g337, g339}, g340);
	defparam lut_3122.LUT_SIZE = 6;
	defparam lut_3122.mask = 64'h000000000000030b;

	lut_sub lut_3132 ({g2, i_7_, g29, i_37_}, g341);
	defparam lut_3132.LUT_SIZE = 4;
	defparam lut_3132.mask = 16'h0010;

	lut_sub lut_3139 ({g3, i_29_, g55, g341}, g342);
	defparam lut_3139.LUT_SIZE = 4;
	defparam lut_3139.mask = 16'h0010;

	lut_sub lut_3147 ({i_14_, g111, g254, g263, g323}, g343);
	defparam lut_3147.LUT_SIZE = 5;
	defparam lut_3147.mask = 32'h00010000;

	lut_sub lut_3155 ({i_14_, i_21_, g84, g88, g223, g254}, g344);
	defparam lut_3155.LUT_SIZE = 6;
	defparam lut_3155.mask = 64'h0011131300000303;

	lut_sub lut_3174 ({i_34_, g71, g342, g343, g344}, g345);
	defparam lut_3174.LUT_SIZE = 5;
	defparam lut_3174.mask = 32'h80c0c0c0;

	lut_sub lut_3189 ({g100, g254, g308, g340, g345}, g346);
	defparam lut_3189.LUT_SIZE = 5;
	defparam lut_3189.mask = 32'h44444440;

	lut_sub lut_3202 ({g53, g10, i_10_, g42}, g347);
	defparam lut_3202.LUT_SIZE = 4;
	defparam lut_3202.mask = 16'h0004;

	lut_sub lut_3209 ({g45, i_10_, g49, g35}, g348);
	defparam lut_3209.LUT_SIZE = 4;
	defparam lut_3209.mask = 16'h0010;

	lut_sub lut_3215 ({i_33_, i_34_, i_35_, g347, g348}, g349);
	defparam lut_3215.LUT_SIZE = 5;
	defparam lut_3215.mask = 32'h00700000;

	lut_sub lut_3225 ({g77, g16, g78, g107}, g350);
	defparam lut_3225.LUT_SIZE = 4;
	defparam lut_3225.mask = 16'h1555;

	lut_sub lut_3237 ({g197, i_20_, i_0_, g320}, g351);
	defparam lut_3237.LUT_SIZE = 4;
	defparam lut_3237.mask = 16'h0040;

	lut_sub lut_3243 ({i_33_, i_34_, g21, g285}, g352);
	defparam lut_3243.LUT_SIZE = 4;
	defparam lut_3243.mask = 16'h0100;

	lut_sub lut_3250 ({i_33_, g2, g37, g38}, g353);
	defparam lut_3250.LUT_SIZE = 4;
	defparam lut_3250.mask = 16'h0100;

	lut_sub lut_3259 ({g45, i_10_, g32, g35, g277, g353}, g354);
	defparam lut_3259.LUT_SIZE = 6;
	defparam lut_3259.mask = 64'h0000000000570000;

	lut_sub lut_3272 ({g33, g101, g351, g352, g354}, g355);
	defparam lut_3272.LUT_SIZE = 5;
	defparam lut_3272.mask = 32'h88888880;

	lut_sub lut_3287 ({g76, g110, g349, g350, g355}, g356);
	defparam lut_3287.LUT_SIZE = 5;
	defparam lut_3287.mask = 32'h50004000;

	lut_sub lut_3297 ({i_32_, i_37_, g322, g333, g346, g356}, g357);
	defparam lut_3297.LUT_SIZE = 6;
	defparam lut_3297.mask = 64'hccccfeff0000aaaa;

	lut_sub lut_3333 ({g23, g310}, g358);
	defparam lut_3333.LUT_SIZE = 2;
	defparam lut_3333.mask = 4'b0001;

	lut_sub lut_3341 ({g7, g335, g248, g323}, g359);
	defparam lut_3341.LUT_SIZE = 4;
	defparam lut_3341.mask = 16'h0001;

	lut_sub lut_3347 ({g2, i_7_, i_32_, g97}, g360);
	defparam lut_3347.LUT_SIZE = 4;
	defparam lut_3347.mask = 16'h0040;

	lut_sub lut_3355 ({g111, g24, g359, g360}, g361);
	defparam lut_3355.LUT_SIZE = 4;
	defparam lut_3355.mask = 16'haa8a;

	lut_sub lut_3368 ({g6, g17, i_37_, g361}, g362);
	defparam lut_3368.LUT_SIZE = 4;
	defparam lut_3368.mask = 16'h2322;

	lut_sub lut_3378 ({i_10_, g11, g197}, g363);
	defparam lut_3378.LUT_SIZE = 3;
	defparam lut_3378.mask = 8'h8a;

	lut_sub lut_3385 ({i_24_, i_34_, i_23_, g1, i_37_}, g364);
	defparam lut_3385.LUT_SIZE = 5;
	defparam lut_3385.mask = 32'h00100000;

	lut_sub lut_3393 ({i_7_, g85, g86, g254, g364}, g365);
	defparam lut_3393.LUT_SIZE = 5;
	defparam lut_3393.mask = 32'h50730033;

	lut_sub lut_3411 ({i_14_, g358, g362, g363, g365}, g366);
	defparam lut_3411.LUT_SIZE = 5;
	defparam lut_3411.mask = 32'h5fdf0000;

	lut_sub lut_3427 ({i_33_, i_32_, i_29_}, g367);
	defparam lut_3427.LUT_SIZE = 3;
	defparam lut_3427.mask = 8'h80;

	lut_sub lut_3431 ({i_24_, i_23_, i_30_, i_8_}, g368);
	defparam lut_3431.LUT_SIZE = 4;
	defparam lut_3431.mask = 16'h8000;

	lut_sub lut_3437 ({i_33_, i_29_, g243, g368}, g369);
	defparam lut_3437.LUT_SIZE = 4;
	defparam lut_3437.mask = 16'h1000;

	lut_sub lut_3445 ({g254, g367, g369, g278}, g370);
	defparam lut_3445.LUT_SIZE = 4;
	defparam lut_3445.mask = 16'h003b;

	lut_sub lut_3454 ({i_3_, i_18_, g12}, g371);
	defparam lut_3454.LUT_SIZE = 3;
	defparam lut_3454.mask = 8'ha2;

	lut_sub lut_3461 ({i_17_, i_9_, g371}, g372);
	defparam lut_3461.LUT_SIZE = 3;
	defparam lut_3461.mask = 8'h80;

	lut_sub lut_3465 ({i_16_, i_7_, i_8_, i_0_, i_37_}, g373);
	defparam lut_3465.LUT_SIZE = 5;
	defparam lut_3465.mask = 32'h40000000;

	lut_sub lut_3471 ({i_33_, i_13_, i_14_, g14, g373}, g374);
	defparam lut_3471.LUT_SIZE = 5;
	defparam lut_3471.mask = 32'h11101010;

	lut_sub lut_3482 ({i_7_, g53, g286, g263}, g375);
	defparam lut_3482.LUT_SIZE = 4;
	defparam lut_3482.mask = 16'h0100;

	lut_sub lut_3489 ({i_29_, i_8_, g263, g267, g375}, g376);
	defparam lut_3489.LUT_SIZE = 5;
	defparam lut_3489.mask = 32'h0000a8aa;

	lut_sub lut_3501 ({i_17_, g33, g49}, g377);
	defparam lut_3501.LUT_SIZE = 3;
	defparam lut_3501.mask = 8'h10;

	lut_sub lut_3508 ({g33, i_29_, i_20_, g377, g255}, g378);
	defparam lut_3508.LUT_SIZE = 5;
	defparam lut_3508.mask = 32'h110011f0;

	lut_sub lut_3523 ({i_12_, g372, g374, g376, g378}, g379);
	defparam lut_3523.LUT_SIZE = 5;
	defparam lut_3523.mask = 32'h45454445;

	lut_sub lut_3542 ({g101, g202, g366, g370, g379}, g380);
	defparam lut_3542.LUT_SIZE = 5;
	defparam lut_3542.mask = 32'hf0f08000;

	lut_sub lut_3559 ({g45, g286, g326, g328, g331}, g381);
	defparam lut_3559.LUT_SIZE = 5;
	defparam lut_3559.mask = 32'h0000007f;

	lut_sub lut_3571 ({i_34_, i_13_, g58, g254}, g382);
	defparam lut_3571.LUT_SIZE = 4;
	defparam lut_3571.mask = 16'h0010;

	lut_sub lut_3579 ({g20, i_34_, g79, i_37_, g367, g382}, g383);
	defparam lut_3579.LUT_SIZE = 6;
	defparam lut_3579.mask = 64'h0000000000000103;

	lut_sub lut_3588 ({i_34_, g53, i_8_, g29, g254}, g384);
	defparam lut_3588.LUT_SIZE = 5;
	defparam lut_3588.mask = 32'h00000010;

	lut_sub lut_3593 ({i_33_, i_34_, g5}, g385);
	defparam lut_3593.LUT_SIZE = 3;
	defparam lut_3593.mask = 8'h20;

	lut_sub lut_3601 ({g1, g18, i_37_, g384, g385}, g386);
	defparam lut_3601.LUT_SIZE = 5;
	defparam lut_3601.mask = 32'h00000105;

	lut_sub lut_3611 ({i_33_, g7, g65, g263, g336}, g387);
	defparam lut_3611.LUT_SIZE = 5;
	defparam lut_3611.mask = 32'h03570000;

	lut_sub lut_3623 ({g94, i_7_, i_0_, g286}, g388);
	defparam lut_3623.LUT_SIZE = 4;
	defparam lut_3623.mask = 16'h0040;

	lut_sub lut_3630 ({g111, i_37_, g387, g388}, g389);
	defparam lut_3630.LUT_SIZE = 4;
	defparam lut_3630.mask = 16'haaa8;

	lut_sub lut_3643 ({i_33_, g54, g152, i_20_, g254}, g390);
	defparam lut_3643.LUT_SIZE = 5;
	defparam lut_3643.mask = 32'h04040004;

	lut_sub lut_3653 ({i_33_, g28, g54, g48, g254}, g391);
	defparam lut_3653.LUT_SIZE = 5;
	defparam lut_3653.mask = 32'h00110001;

	lut_sub lut_3662 ({g111, g13, i_20_, g391}, g392);
	defparam lut_3662.LUT_SIZE = 4;
	defparam lut_3662.mask = 16'h0004;

	lut_sub lut_3669 ({g111, i_6_, i_8_, g390, g392}, g393);
	defparam lut_3669.LUT_SIZE = 5;
	defparam lut_3669.mask = 32'haaaa8aaa;

	lut_sub lut_3691 ({i_13_, g248, g323, g389, g393}, g394);
	defparam lut_3691.LUT_SIZE = 5;
	defparam lut_3691.mask = 32'h0cae00aa;

	lut_sub lut_3708 ({i_33_, g45, i_8_, g35, g254}, g395);
	defparam lut_3708.LUT_SIZE = 5;
	defparam lut_3708.mask = 32'h00100000;

	lut_sub lut_3714 ({i_28_, g33, g132, i_25_, i_20_}, g396);
	defparam lut_3714.LUT_SIZE = 5;
	defparam lut_3714.mask = 32'h00010000;

	lut_sub lut_3720 ({i_34_, i_30_, g395, g396}, g397);
	defparam lut_3720.LUT_SIZE = 4;
	defparam lut_3720.mask = 16'h0070;

	lut_sub lut_3726 ({i_34_, i_35_, i_21_, i_29_, i_22_}, g398);
	defparam lut_3726.LUT_SIZE = 5;
	defparam lut_3726.mask = 32'h00130303;

	lut_sub lut_3736 ({i_24_, i_34_, i_26_, i_22_}, g399);
	defparam lut_3736.LUT_SIZE = 4;
	defparam lut_3736.mask = 16'h23ab;

	lut_sub lut_3748 ({i_21_, i_29_, i_20_, g399}, g400);
	defparam lut_3748.LUT_SIZE = 4;
	defparam lut_3748.mask = 16'h0400;

	lut_sub lut_3753 ({i_24_, i_34_, i_35_, i_26_, g157}, g401);
	defparam lut_3753.LUT_SIZE = 5;
	defparam lut_3753.mask = 32'h45550500;

	lut_sub lut_3770 ({g3, g164, g398, g400, g401}, g402);
	defparam lut_3770.LUT_SIZE = 5;
	defparam lut_3770.mask = 32'h00000444;

	lut_sub lut_3778 ({g2, i_21_, g88, i_22_}, g403);
	defparam lut_3778.LUT_SIZE = 4;
	defparam lut_3778.mask = 16'h0013;

	lut_sub lut_3787 ({i_7_, g1, g279, g403}, g404);
	defparam lut_3787.LUT_SIZE = 4;
	defparam lut_3787.mask = 16'ha8aa;

	lut_sub lut_3800 ({g86, g143, i_25_, g404}, g405);
	defparam lut_3800.LUT_SIZE = 4;
	defparam lut_3800.mask = 16'hab00;

	lut_sub lut_3811 ({i_33_, g28, g54, g254}, g406);
	defparam lut_3811.LUT_SIZE = 4;
	defparam lut_3811.mask = 16'h0501;

	lut_sub lut_3819 ({i_8_, i_0_, g327, g406}, g407);
	defparam lut_3819.LUT_SIZE = 4;
	defparam lut_3819.mask = 16'h1000;

	lut_sub lut_3827 ({g94, i_8_, i_0_, g323, g390, g259}, g408);
	defparam lut_3827.LUT_SIZE = 6;
	defparam lut_3827.mask = 64'h0000000037000000;

	lut_sub lut_3836 ({i_24_, i_34_, i_35_, i_26_, g334}, g409);
	defparam lut_3836.LUT_SIZE = 5;
	defparam lut_3836.mask = 32'hceee0a00;

	lut_sub lut_3855 ({g3, i_7_, i_31_, g157, g409}, g410);
	defparam lut_3855.LUT_SIZE = 5;
	defparam lut_3855.mask = 32'h00000001;

	lut_sub lut_3863 ({i_34_, g57, g88, g137, g410}, g411);
	defparam lut_3863.LUT_SIZE = 5;
	defparam lut_3863.mask = 32'haaaaaaa8;

	lut_sub lut_3882 ({i_13_, i_14_, g11}, g412);
	defparam lut_3882.LUT_SIZE = 3;
	defparam lut_3882.mask = 8'h04;

	lut_sub lut_3891 ({g358, g311, g377, g249, g412}, g413);
	defparam lut_3891.LUT_SIZE = 5;
	defparam lut_3891.mask = 32'h00035557;

	lut_sub lut_3910 ({g405, g407, g408, g411, g413}, g414);
	defparam lut_3910.LUT_SIZE = 5;
	defparam lut_3910.mask = 32'h20000000;

	lut_sub lut_3919 ({i_34_, g135, g156, g397, g402, g414}, g415);
	defparam lut_3919.LUT_SIZE = 6;
	defparam lut_3919.mask = 64'h0040004000400000;

	lut_sub lut_3926 ({i_14_, i_32_, g58}, g416);
	defparam lut_3926.LUT_SIZE = 3;
	defparam lut_3926.mask = 8'h40;

	lut_sub lut_3933 ({i_33_, i_34_, g21, g247, g416}, g417);
	defparam lut_3933.LUT_SIZE = 5;
	defparam lut_3933.mask = 32'h000d0005;

	lut_sub lut_3944 ({i_34_, g1, i_8_, g5, g29}, g418);
	defparam lut_3944.LUT_SIZE = 5;
	defparam lut_3944.mask = 32'h00000040;

	lut_sub lut_3952 ({g98, g55, g277, g418}, g419);
	defparam lut_3952.LUT_SIZE = 4;
	defparam lut_3952.mask = 16'h0537;

	lut_sub lut_3964 ({i_33_, i_32_, g122, g419}, g420);
	defparam lut_3964.LUT_SIZE = 4;
	defparam lut_3964.mask = 16'h8aaa;

	lut_sub lut_3977 ({i_33_, g2, i_32_, g150, g134}, g421);
	defparam lut_3977.LUT_SIZE = 5;
	defparam lut_3977.mask = 32'h00700050;

	lut_sub lut_3986 ({i_30_, i_31_, i_29_, i_37_, g421}, g422);
	defparam lut_3986.LUT_SIZE = 5;
	defparam lut_3986.mask = 32'h00100000;

	lut_sub lut_3993 ({g53, g367, g341}, g423);
	defparam lut_3993.LUT_SIZE = 3;
	defparam lut_3993.mask = 8'h01;

	lut_sub lut_4001 ({i_29_, g18, g279, g422, g423}, g424);
	defparam lut_4001.LUT_SIZE = 5;
	defparam lut_4001.mask = 32'h88808888;

	lut_sub lut_4016 ({g3, g254, g417, g420, g424}, g425);
	defparam lut_4016.LUT_SIZE = 5;
	defparam lut_4016.mask = 32'hff305510;

	lut_sub lut_4040 ({g381, g383, g386, g394, g415, g425}, g426);
	defparam lut_4040.LUT_SIZE = 6;
	defparam lut_4040.mask = 64'h1000000000000000;

	lut_sub lut_4049 ({g293, g319, g357, g380, g426}, g427);
	defparam lut_4049.LUT_SIZE = 5;
	defparam lut_4049.mask = 32'h00100000;

	lut_sub lut_4053 ({i_35_, i_38_}, g428);
	defparam lut_4053.LUT_SIZE = 2;
	defparam lut_4053.mask = 4'b0100;

	lut_sub lut_4058 ({i_33_, g428}, g429);
	defparam lut_4058.LUT_SIZE = 2;
	defparam lut_4058.mask = 4'b0100;

	lut_sub lut_4064 ({i_9_, i_8_, g9, i_10_, g29}, g430);
	defparam lut_4064.LUT_SIZE = 5;
	defparam lut_4064.mask = 32'h00004c00;

	lut_sub lut_4071 ({i_33_, i_7_, g70, i_38_}, g431);
	defparam lut_4071.LUT_SIZE = 4;
	defparam lut_4071.mask = 16'h4000;

	lut_sub lut_4078 ({i_2_, i_8_, g96, g429, g431}, g432);
	defparam lut_4078.LUT_SIZE = 5;
	defparam lut_4078.mask = 32'h57550000;

	lut_sub lut_4094 ({i_33_, g57, g9, g29, g428}, g433);
	defparam lut_4094.LUT_SIZE = 5;
	defparam lut_4094.mask = 32'h00150000;

	lut_sub lut_4102 ({i_23_, i_29_, g157, g433}, g434);
	defparam lut_4102.LUT_SIZE = 4;
	defparam lut_4102.mask = 16'ha2a0;

	lut_sub lut_4111 ({i_31_, g428}, g435);
	defparam lut_4111.LUT_SIZE = 2;
	defparam lut_4111.mask = 4'b0100;

	lut_sub lut_4116 ({i_2_, i_7_, i_9_, i_3_, i_18_, g14}, g436);
	defparam lut_4116.LUT_SIZE = 6;
	defparam lut_4116.mask = 64'h0400000000000000;

	lut_sub lut_4123 ({g12, g32, g436}, g437);
	defparam lut_4123.LUT_SIZE = 3;
	defparam lut_4123.mask = 8'ha8;

	lut_sub lut_4131 ({i_32_, g25, g437}, g438);
	defparam lut_4131.LUT_SIZE = 3;
	defparam lut_4131.mask = 8'h4c;

	lut_sub lut_4139 ({i_9_, i_3_, i_18_, g14, g46}, g439);
	defparam lut_4139.LUT_SIZE = 5;
	defparam lut_4139.mask = 32'h00100000;

	lut_sub lut_4146 ({g12, g49, g439}, g440);
	defparam lut_4146.LUT_SIZE = 3;
	defparam lut_4146.mask = 8'ha8;

	lut_sub lut_4155 ({i_33_, i_38_, g435, g438, g440}, g441);
	defparam lut_4155.LUT_SIZE = 5;
	defparam lut_4155.mask = 32'h0ace0000;

	lut_sub lut_4171 ({g121, g429, g430, g432, g434, g441}, g442);
	defparam lut_4171.LUT_SIZE = 6;
	defparam lut_4171.mask = 64'h00000000dfdfdfff;

	lut_sub lut_4204 ({g71, i_25_}, g443);
	defparam lut_4204.LUT_SIZE = 2;
	defparam lut_4204.mask = 4'b1000;

	lut_sub lut_4210 ({i_35_, i_31_, g438, g440}, g444);
	defparam lut_4210.LUT_SIZE = 4;
	defparam lut_4210.mask = 16'h1333;

	lut_sub lut_4223 ({i_32_, i_31_, g9, g29, g428}, g445);
	defparam lut_4223.LUT_SIZE = 5;
	defparam lut_4223.mask = 32'h15000000;

	lut_sub lut_4231 ({i_2_, i_7_, g70, i_38_, g445}, g446);
	defparam lut_4231.LUT_SIZE = 5;
	defparam lut_4231.mask = 32'h8aaaaaaa;

	lut_sub lut_4254 ({g46, g223, g428, g430, g446}, g447);
	defparam lut_4254.LUT_SIZE = 5;
	defparam lut_4254.mask = 32'h54545450;

	lut_sub lut_4271 ({i_28_, i_38_, g443, g444, g447}, g448);
	defparam lut_4271.LUT_SIZE = 5;
	defparam lut_4271.mask = 32'h0a0e0000;

	lut_sub lut_4281 ({i_18_, i_11_, i_19_, g67, g10}, g449);
	defparam lut_4281.LUT_SIZE = 5;
	defparam lut_4281.mask = 32'h73335000;

	lut_sub lut_4297 ({i_32_, i_25_, g449, g435}, g450);
	defparam lut_4297.LUT_SIZE = 4;
	defparam lut_4297.mask = 16'h1000;

	lut_sub lut_4303 ({i_7_, i_8_, g9, g29}, g451);
	defparam lut_4303.LUT_SIZE = 4;
	defparam lut_4303.mask = 16'h7000;

	lut_sub lut_4311 ({i_9_, g65, g9, i_10_}, g452);
	defparam lut_4311.LUT_SIZE = 4;
	defparam lut_4311.mask = 16'h0002;

	lut_sub lut_4317 ({i_33_, i_31_, g65, g449}, g453);
	defparam lut_4317.LUT_SIZE = 4;
	defparam lut_4317.mask = 16'h1000;

	lut_sub lut_4325 ({g164, i_38_, g451, g452, g453}, g454);
	defparam lut_4325.LUT_SIZE = 5;
	defparam lut_4325.mask = 32'h007f0055;

	lut_sub lut_4341 ({i_8_, g9, g29}, g455);
	defparam lut_4341.LUT_SIZE = 3;
	defparam lut_4341.mask = 8'h70;

	lut_sub lut_4347 ({i_13_, i_9_, i_18_}, g456);
	defparam lut_4347.LUT_SIZE = 3;
	defparam lut_4347.mask = 8'h10;

	lut_sub lut_4353 ({i_11_, g455, g456}, g457);
	defparam lut_4353.LUT_SIZE = 3;
	defparam lut_4353.mask = 8'h01;

	lut_sub lut_4359 ({i_12_, i_9_, i_3_, g14, i_1_, g46}, g458);
	defparam lut_4359.LUT_SIZE = 6;
	defparam lut_4359.mask = 64'h0000050000000400;

	lut_sub lut_4366 ({i_13_, i_11_, g458}, g459);
	defparam lut_4366.LUT_SIZE = 3;
	defparam lut_4366.mask = 8'h10;

	lut_sub lut_4370 ({i_33_, i_30_, i_32_, i_31_, i_25_}, g460);
	defparam lut_4370.LUT_SIZE = 5;
	defparam lut_4370.mask = 32'hc0008000;

	lut_sub lut_4381 ({i_2_, g164, g428, g457, g459, g460}, g461);
	defparam lut_4381.LUT_SIZE = 6;
	defparam lut_4381.mask = 64'h007f0055003f0000;

	lut_sub lut_4404 ({i_24_, i_28_, i_26_, g450, g454, g461}, g462);
	defparam lut_4404.LUT_SIZE = 6;
	defparam lut_4404.mask = 64'h7f00000000000000;

	lut_sub lut_4417 ({i_32_, g223, g443, g428}, g463);
	defparam lut_4417.LUT_SIZE = 4;
	defparam lut_4417.mask = 16'h0100;

	lut_sub lut_4425 ({i_12_, g86, g121, g429, g463}, g464);
	defparam lut_4425.LUT_SIZE = 5;
	defparam lut_4425.mask = 32'h00005755;

	lut_sub lut_4437 ({i_35_, i_31_, i_8_, i_38_}, g465);
	defparam lut_4437.LUT_SIZE = 4;
	defparam lut_4437.mask = 16'h4000;

	lut_sub lut_4443 ({i_7_, i_32_, g335, i_38_, g465}, g466);
	defparam lut_4443.LUT_SIZE = 5;
	defparam lut_4443.mask = 32'h07050505;

	lut_sub lut_4456 ({i_28_, i_26_, i_25_, g466}, g467);
	defparam lut_4456.LUT_SIZE = 4;
	defparam lut_4456.mask = 16'h4000;

	lut_sub lut_4461 ({i_28_, i_26_, i_31_, g48}, g468);
	defparam lut_4461.LUT_SIZE = 4;
	defparam lut_4461.mask = 16'h4000;

	lut_sub lut_4466 ({i_28_, i_26_, i_32_, g31}, g469);
	defparam lut_4466.LUT_SIZE = 4;
	defparam lut_4466.mask = 16'h4000;

	lut_sub lut_4472 ({i_33_, i_35_, i_38_, g468, g469}, g470);
	defparam lut_4472.LUT_SIZE = 5;
	defparam lut_4472.mask = 32'h07050000;

	lut_sub lut_4483 ({i_24_, g8, g467, g470}, g471);
	defparam lut_4483.LUT_SIZE = 4;
	defparam lut_4483.mask = 16'h0700;

	lut_sub lut_4489 ({i_35_, i_30_, i_32_, i_38_}, g472);
	defparam lut_4489.LUT_SIZE = 4;
	defparam lut_4489.mask = 16'h4000;

	lut_sub lut_4495 ({i_33_, i_28_, g71, i_25_, g472}, g473);
	defparam lut_4495.LUT_SIZE = 5;
	defparam lut_4495.mask = 32'h50004000;

	lut_sub lut_4501 ({i_13_, i_3_, i_11_}, g474);
	defparam lut_4501.LUT_SIZE = 3;
	defparam lut_4501.mask = 8'h40;

	lut_sub lut_4507 ({i_2_, i_9_, g473, g474}, g475);
	defparam lut_4507.LUT_SIZE = 4;
	defparam lut_4507.mask = 16'hfeff;

	lut_sub lut_4529 ({i_13_, i_9_, g160, g464, g471, g696}, g476);
	defparam lut_4529.LUT_SIZE = 6;
	defparam lut_4529.mask = 64'h5500500044004000;

	lut_sub lut_4546 ({i_22_, g160, g442, g448, g462, g476}, g477);
	defparam lut_4546.LUT_SIZE = 6;
	defparam lut_4546.mask = 64'h40004000ffff4000;

	lut_sub lut_4568 ({i_24_, i_25_}, g478);
	defparam lut_4568.LUT_SIZE = 2;
	defparam lut_4568.mask = 4'b1000;

	lut_sub lut_4572 ({i_33_, i_28_, i_32_, i_29_, i_25_}, g479);
	defparam lut_4572.LUT_SIZE = 5;
	defparam lut_4572.mask = 32'hc0008000;

	lut_sub lut_4580 ({i_24_, i_30_, g1, g7, i_25_}, g480);
	defparam lut_4580.LUT_SIZE = 5;
	defparam lut_4580.mask = 32'h02000000;

	lut_sub lut_4588 ({i_24_, g32, g24, g479, g480}, g481);
	defparam lut_4588.LUT_SIZE = 5;
	defparam lut_4588.mask = 32'haa8aaaaa;

	lut_sub lut_4609 ({i_33_, i_24_, g1, g25, g481}, g482);
	defparam lut_4609.LUT_SIZE = 5;
	defparam lut_4609.mask = 32'h54555555;

	lut_sub lut_4630 ({i_7_, i_32_, g84, g478, g482}, g483);
	defparam lut_4630.LUT_SIZE = 5;
	defparam lut_4630.mask = 32'h54555555;

	lut_sub lut_4651 ({i_24_, g12, g32, g436}, g484);
	defparam lut_4651.LUT_SIZE = 4;
	defparam lut_4651.mask = 16'h5700;

	lut_sub lut_4661 ({g37, g484}, g485);
	defparam lut_4661.LUT_SIZE = 2;
	defparam lut_4661.mask = 4'b0001;

	lut_sub lut_4668 ({g12, i_8_, g11, g436}, g486);
	defparam lut_4668.LUT_SIZE = 4;
	defparam lut_4668.mask = 16'h5073;

	lut_sub lut_4681 ({i_24_, i_30_, g1, g7, g486}, g487);
	defparam lut_4681.LUT_SIZE = 5;
	defparam lut_4681.mask = 32'h07050000;

	lut_sub lut_4689 ({i_24_, i_28_}, g488);
	defparam lut_4689.LUT_SIZE = 2;
	defparam lut_4689.mask = 4'b1000;

	lut_sub lut_4695 ({i_7_, i_29_, g70, g488}, g489);
	defparam lut_4695.LUT_SIZE = 4;
	defparam lut_4695.mask = 16'h4000;

	lut_sub lut_4703 ({i_33_, i_38_, g483, g485, g487, g489}, g490);
	defparam lut_4703.LUT_SIZE = 6;
	defparam lut_4703.mask = 64'h0000ff7f0000ff00;

	lut_sub lut_4729 ({i_24_, i_9_, i_10_}, g491);
	defparam lut_4729.LUT_SIZE = 3;
	defparam lut_4729.mask = 8'h20;

	lut_sub lut_4734 ({i_30_, i_32_, g428}, g492);
	defparam lut_4734.LUT_SIZE = 3;
	defparam lut_4734.mask = 8'h40;

	lut_sub lut_4741 ({g1, i_25_, g491, g492}, g493);
	defparam lut_4741.LUT_SIZE = 4;
	defparam lut_4741.mask = 16'h0010;

	lut_sub lut_4746 ({i_28_, g478}, g494);
	defparam lut_4746.LUT_SIZE = 2;
	defparam lut_4746.mask = 4'b0100;

	lut_sub lut_4750 ({i_9_, i_8_, i_10_}, g495);
	defparam lut_4750.LUT_SIZE = 3;
	defparam lut_4750.mask = 8'h08;

	lut_sub lut_4757 ({i_30_, i_29_, g428, g494, g495}, g496);
	defparam lut_4757.LUT_SIZE = 5;
	defparam lut_4757.mask = 32'h01000000;

	lut_sub lut_4766 ({g84, g478, g465, g493, g496}, g497);
	defparam lut_4766.LUT_SIZE = 5;
	defparam lut_4766.mask = 32'h88888880;

	lut_sub lut_4779 ({i_24_, g12, g49, g439}, g498);
	defparam lut_4779.LUT_SIZE = 4;
	defparam lut_4779.mask = 16'h5700;

	lut_sub lut_4789 ({i_24_, i_35_, i_31_, g25, g498}, g499);
	defparam lut_4789.LUT_SIZE = 5;
	defparam lut_4789.mask = 32'h73335000;

	lut_sub lut_4804 ({g1, i_25_, i_38_}, g500);
	defparam lut_4804.LUT_SIZE = 3;
	defparam lut_4804.mask = 8'h04;

	lut_sub lut_4810 ({i_29_, g494, g435}, g501);
	defparam lut_4810.LUT_SIZE = 3;
	defparam lut_4810.mask = 8'h10;

	lut_sub lut_4818 ({i_24_, g60, g429, g455, g501}, g502);
	defparam lut_4818.LUT_SIZE = 5;
	defparam lut_4818.mask = 32'h11131111;

	lut_sub lut_4834 ({i_32_, g484, g499, g500, g502}, g503);
	defparam lut_4834.LUT_SIZE = 5;
	defparam lut_4834.mask = 32'ha888a8a8;

	lut_sub lut_4849 ({i_24_, i_17_, i_12_, g22}, g504);
	defparam lut_4849.LUT_SIZE = 4;
	defparam lut_4849.mask = 16'h5700;

	lut_sub lut_4858 ({i_28_, i_31_, i_29_, g504}, g505);
	defparam lut_4858.LUT_SIZE = 4;
	defparam lut_4858.mask = 16'h0400;

	lut_sub lut_4865 ({i_24_, i_30_, g1, g429, g495}, g506);
	defparam lut_4865.LUT_SIZE = 5;
	defparam lut_4865.mask = 32'h01000000;

	lut_sub lut_4871 ({i_17_, i_12_, g22, g86}, g507);
	defparam lut_4871.LUT_SIZE = 4;
	defparam lut_4871.mask = 16'h1115;

	lut_sub lut_4881 ({i_23_, i_22_, g488, g507}, g508);
	defparam lut_4881.LUT_SIZE = 4;
	defparam lut_4881.mask = 16'h0103;

	lut_sub lut_4891 ({i_14_, g133, g505, g506, g508}, g509);
	defparam lut_4891.LUT_SIZE = 5;
	defparam lut_4891.mask = 32'h80808000;

	lut_sub lut_4901 ({i_34_, g490, g497, g503, g509}, g510);
	defparam lut_4901.LUT_SIZE = 5;
	defparam lut_4901.mask = 32'h0000feff;

	lut_sub lut_4921 ({i_30_, g121, g495}, g511);
	defparam lut_4921.LUT_SIZE = 3;
	defparam lut_4921.mask = 8'h10;

	lut_sub lut_4926 ({i_34_, i_26_, g488}, g512);
	defparam lut_4926.LUT_SIZE = 3;
	defparam lut_4926.mask = 8'h45;

	lut_sub lut_4936 ({i_33_, i_29_, g457, g459, g511, g512}, g513);
	defparam lut_4936.LUT_SIZE = 6;
	defparam lut_4936.mask = 64'h3777000000000000;

	lut_sub lut_4953 ({i_13_, i_11_, g478, g457, g458}, g514);
	defparam lut_4953.LUT_SIZE = 5;
	defparam lut_4953.mask = 32'h03070000;

	lut_sub lut_4961 ({i_34_, i_26_, i_29_, i_22_}, g515);
	defparam lut_4961.LUT_SIZE = 4;
	defparam lut_4961.mask = 16'he0ec;

	lut_sub lut_4974 ({i_13_, i_19_, g488, g458}, g516);
	defparam lut_4974.LUT_SIZE = 4;
	defparam lut_4974.mask = 16'h0100;

	lut_sub lut_4979 ({i_13_, i_18_, i_19_, g488}, g517);
	defparam lut_4979.LUT_SIZE = 4;
	defparam lut_4979.mask = 16'h0100;

	lut_sub lut_4986 ({i_9_, i_8_, g9, g29, g517}, g518);
	defparam lut_4986.LUT_SIZE = 5;
	defparam lut_4986.mask = 32'h00001500;

	lut_sub lut_4996 ({g164, g515, g516, g518}, g519);
	defparam lut_4996.LUT_SIZE = 4;
	defparam lut_4996.mask = 16'h0700;

	lut_sub lut_5003 ({i_26_, i_29_, i_22_, g488}, g520);
	defparam lut_5003.LUT_SIZE = 4;
	defparam lut_5003.mask = 16'h5400;

	lut_sub lut_5011 ({i_31_, i_25_, g520, g455}, g521);
	defparam lut_5011.LUT_SIZE = 4;
	defparam lut_5011.mask = 16'h1000;

	lut_sub lut_5020 ({g84, g277, g443, g491, g495}, g522);
	defparam lut_5020.LUT_SIZE = 5;
	defparam lut_5020.mask = 32'h00000537;

	lut_sub lut_5031 ({i_34_, i_26_, i_29_, g488}, g523);
	defparam lut_5031.LUT_SIZE = 4;
	defparam lut_5031.mask = 16'h4044;

	lut_sub lut_5038 ({i_12_, i_2_, g14, i_1_}, g524);
	defparam lut_5038.LUT_SIZE = 4;
	defparam lut_5038.mask = 16'h3020;

	lut_sub lut_5048 ({g57, g164, g523, g524}, g525);
	defparam lut_5048.LUT_SIZE = 4;
	defparam lut_5048.mask = 16'h0010;

	lut_sub lut_5055 ({i_9_, i_8_, g9, g70, g29}, g526);
	defparam lut_5055.LUT_SIZE = 5;
	defparam lut_5055.mask = 32'h22332033;

	lut_sub lut_5070 ({i_28_, i_26_, g478}, g527);
	defparam lut_5070.LUT_SIZE = 3;
	defparam lut_5070.mask = 8'h40;

	lut_sub lut_5075 ({i_29_, i_9_, i_10_, g527}, g528);
	defparam lut_5075.LUT_SIZE = 4;
	defparam lut_5075.mask = 16'h0400;

	lut_sub lut_5084 ({g521, g522, g525, g526, g528}, g529);
	defparam lut_5084.LUT_SIZE = 5;
	defparam lut_5084.mask = 32'hb0000000;

	lut_sub lut_5094 ({i_34_, g1, g514, g519, g529}, g530);
	defparam lut_5094.LUT_SIZE = 5;
	defparam lut_5094.mask = 32'h44444440;

	lut_sub lut_5107 ({i_24_, i_30_, i_32_, g7, g484, g499}, g531);
	defparam lut_5107.LUT_SIZE = 6;
	defparam lut_5107.mask = 64'h80a088aa88aa88aa;

	lut_sub lut_5132 ({i_33_, i_34_, g428}, g532);
	defparam lut_5132.LUT_SIZE = 3;
	defparam lut_5132.mask = 8'h10;

	lut_sub lut_5138 ({i_33_, i_26_, g84, g65, i_38_}, g533);
	defparam lut_5138.LUT_SIZE = 5;
	defparam lut_5138.mask = 32'h01000000;

	lut_sub lut_5146 ({g1, g70, g532, g533}, g534);
	defparam lut_5146.LUT_SIZE = 4;
	defparam lut_5146.mask = 16'haa8a;

	lut_sub lut_5157 ({i_26_, g1}, g535);
	defparam lut_5157.LUT_SIZE = 2;
	defparam lut_5157.mask = 4'b0100;

	lut_sub lut_5165 ({g84, g66, i_38_, g535, g492}, g536);
	defparam lut_5165.LUT_SIZE = 5;
	defparam lut_5165.mask = 32'h1111111f;

	lut_sub lut_5181 ({g478, g536}, g537);
	defparam lut_5181.LUT_SIZE = 2;
	defparam lut_5181.mask = 4'b0001;

	lut_sub lut_5188 ({i_24_, i_11_, g456, g534, g537}, g538);
	defparam lut_5188.LUT_SIZE = 5;
	defparam lut_5188.mask = 32'h000d0005;

	lut_sub lut_5196 ({i_28_, i_26_, i_29_, i_25_, i_38_}, g539);
	defparam lut_5196.LUT_SIZE = 5;
	defparam lut_5196.mask = 32'h40000000;

	lut_sub lut_5206 ({g428, g513, g530, g531, g538, g539}, g540);
	defparam lut_5206.LUT_SIZE = 6;
	defparam lut_5206.mask = 64'h8c8c8c8c008c0000;

	lut_sub lut_5226 ({i_24_, i_9_, i_8_, g9, i_10_, g29}, g541);
	defparam lut_5226.LUT_SIZE = 6;
	defparam lut_5226.mask = 64'h00004c0000000000;

	lut_sub lut_5235 ({i_33_, g428, g541, g514}, g542);
	defparam lut_5235.LUT_SIZE = 4;
	defparam lut_5235.mask = 16'h0705;

	lut_sub lut_5245 ({i_9_, g9, i_10_, g29}, g543);
	defparam lut_5245.LUT_SIZE = 4;
	defparam lut_5245.mask = 16'h004c;

	lut_sub lut_5253 ({i_32_, g428, g543}, g544);
	defparam lut_5253.LUT_SIZE = 3;
	defparam lut_5253.mask = 8'h10;

	lut_sub lut_5259 ({i_30_, i_32_, i_8_, g449, g435}, g545);
	defparam lut_5259.LUT_SIZE = 5;
	defparam lut_5259.mask = 32'h51501100;

	lut_sub lut_5275 ({g8, g24, g478, g466, g544, g545}, g546);
	defparam lut_5275.LUT_SIZE = 6;
	defparam lut_5275.mask = 64'h00770077007f0077;

	lut_sub lut_5306 ({i_33_, i_38_, g472, g491, g531}, g547);
	defparam lut_5306.LUT_SIZE = 5;
	defparam lut_5306.mask = 32'h03ab0000;

	lut_sub lut_5317 ({i_28_, i_26_, i_30_, i_22_, g478}, g548);
	defparam lut_5317.LUT_SIZE = 5;
	defparam lut_5317.mask = 32'h40000000;

	lut_sub lut_5323 ({i_33_, g71, g428}, g549);
	defparam lut_5323.LUT_SIZE = 3;
	defparam lut_5323.mask = 8'h40;

	lut_sub lut_5331 ({i_22_, g223, g548, g435, g549}, g550);
	defparam lut_5331.LUT_SIZE = 5;
	defparam lut_5331.mask = 32'h03570303;

	lut_sub lut_5345 ({i_33_, i_25_, i_22_, i_38_}, g551);
	defparam lut_5345.LUT_SIZE = 4;
	defparam lut_5345.mask = 16'h4440;

	lut_sub lut_5353 ({i_26_, i_30_, i_7_, i_32_, g488, g551}, g552);
	defparam lut_5353.LUT_SIZE = 6;
	defparam lut_5353.mask = 64'h1000000000000000;

	lut_sub lut_5359 ({i_8_, g550, g552}, g553);
	defparam lut_5359.LUT_SIZE = 3;
	defparam lut_5359.mask = 8'h8a;

	lut_sub lut_5365 ({i_33_, i_12_, i_25_, i_22_, i_38_}, g554);
	defparam lut_5365.LUT_SIZE = 5;
	defparam lut_5365.mask = 32'h00440040;

	lut_sub lut_5373 ({i_24_, i_28_, i_26_, g197, g554}, g555);
	defparam lut_5373.LUT_SIZE = 5;
	defparam lut_5373.mask = 32'h10000000;

	lut_sub lut_5378 ({i_13_, i_18_, i_19_, g555}, g556);
	defparam lut_5378.LUT_SIZE = 4;
	defparam lut_5378.mask = 16'h0100;

	lut_sub lut_5384 ({i_22_, g474, g464}, g557);
	defparam lut_5384.LUT_SIZE = 3;
	defparam lut_5384.mask = 8'h10;

	lut_sub lut_5388 ({i_12_, i_13_, i_18_, i_11_}, g558);
	defparam lut_5388.LUT_SIZE = 4;
	defparam lut_5388.mask = 16'h0010;

	lut_sub lut_5396 ({i_10_, g553, g556, g557, g558}, g559);
	defparam lut_5396.LUT_SIZE = 5;
	defparam lut_5396.mask = 32'h00007f3f;

	lut_sub lut_5415 ({g57, i_29_, i_8_, g96, g449}, g560);
	defparam lut_5415.LUT_SIZE = 5;
	defparam lut_5415.mask = 32'h30007500;

	lut_sub lut_5426 ({i_34_, g428}, g561);
	defparam lut_5426.LUT_SIZE = 2;
	defparam lut_5426.mask = 4'b0001;

	lut_sub lut_5433 ({g479, g561, g543}, g562);
	defparam lut_5433.LUT_SIZE = 3;
	defparam lut_5433.mask = 8'h01;

	lut_sub lut_5438 ({i_16_, i_27_, i_32_, g96}, g563);
	defparam lut_5438.LUT_SIZE = 4;
	defparam lut_5438.mask = 16'hf444;

	lut_sub lut_5449 ({i_28_, i_34_, i_23_, i_29_, i_22_, g563}, g564);
	defparam lut_5449.LUT_SIZE = 6;
	defparam lut_5449.mask = 64'h0000a2f200000000;

	lut_sub lut_5464 ({i_24_, i_28_, g532, g560, g562, g564}, g565);
	defparam lut_5464.LUT_SIZE = 6;
	defparam lut_5464.mask = 64'h777f777700000000;

	lut_sub lut_5498 ({g535, g542, g546, g547, g559, g565}, g566);
	defparam lut_5498.LUT_SIZE = 6;
	defparam lut_5498.mask = 64'h8888888880000000;

	lut_sub lut_5510 ({i_13_, i_3_, i_19_, i_22_}, g567);
	defparam lut_5510.LUT_SIZE = 4;
	defparam lut_5510.mask = 16'h2000;

	lut_sub lut_5515 ({i_13_, i_18_, g12, i_22_}, g568);
	defparam lut_5515.LUT_SIZE = 4;
	defparam lut_5515.mask = 16'h0800;

	lut_sub lut_5521 ({g567, g568}, g569);
	defparam lut_5521.LUT_SIZE = 2;
	defparam lut_5521.mask = 4'b1000;

	lut_sub lut_5528 ({i_12_, g473, g552, g569}, g570);
	defparam lut_5528.LUT_SIZE = 4;
	defparam lut_5528.mask = 16'h003b;

	lut_sub lut_5538 ({i_12_, i_2_, i_22_, g474, g568}, g571);
	defparam lut_5538.LUT_SIZE = 5;
	defparam lut_5538.mask = 32'h55007530;

	lut_sub lut_5556 ({i_28_, g70, g527, g549, g492}, g572);
	defparam lut_5556.LUT_SIZE = 5;
	defparam lut_5556.mask = 32'h37050505;

	lut_sub lut_5571 ({i_12_, i_2_, i_10_, i_22_, g572}, g573);
	defparam lut_5571.LUT_SIZE = 5;
	defparam lut_5571.mask = 32'h40004040;

	lut_sub lut_5579 ({i_35_, i_26_, i_30_, g488, g551}, g574);
	defparam lut_5579.LUT_SIZE = 5;
	defparam lut_5579.mask = 32'h10000000;

	lut_sub lut_5585 ({i_13_, i_3_, i_19_, g46, g574}, g575);
	defparam lut_5585.LUT_SIZE = 5;
	defparam lut_5585.mask = 32'h01000000;

	lut_sub lut_5594 ({g473, g555, g571, g573, g575}, g576);
	defparam lut_5594.LUT_SIZE = 5;
	defparam lut_5594.mask = 32'h88008000;

	lut_sub lut_5602 ({i_24_, i_19_, i_25_, g534, g536}, g577);
	defparam lut_5602.LUT_SIZE = 5;
	defparam lut_5602.mask = 32'h00dc0000;

	lut_sub lut_5613 ({i_24_, g474, g534, g537}, g578);
	defparam lut_5613.LUT_SIZE = 4;
	defparam lut_5613.mask = 16'h0d00;

	lut_sub lut_5621 ({i_13_, i_3_, g577, g578}, g579);
	defparam lut_5621.LUT_SIZE = 4;
	defparam lut_5621.mask = 16'h8aaa;

	lut_sub lut_5632 ({i_33_, g71, i_38_}, g580);
	defparam lut_5632.LUT_SIZE = 3;
	defparam lut_5632.mask = 8'h40;

	lut_sub lut_5641 ({g37, g31, g48, g580, g685}, g581);
	defparam lut_5641.LUT_SIZE = 5;
	defparam lut_5641.mask = 32'h0a0a0a3b;

	lut_sub lut_5657 ({i_32_, i_31_, i_25_, g520, g428}, g582);
	defparam lut_5657.LUT_SIZE = 5;
	defparam lut_5657.mask = 32'h10000000;

	lut_sub lut_5664 ({i_33_, i_34_, g121, g428, g494}, g583);
	defparam lut_5664.LUT_SIZE = 5;
	defparam lut_5664.mask = 32'h03330011;

	lut_sub lut_5677 ({i_26_, i_25_, g488, g583}, g584);
	defparam lut_5677.LUT_SIZE = 4;
	defparam lut_5677.mask = 16'h1110;

	lut_sub lut_5686 ({i_33_, i_24_, g57, g1, g561}, g585);
	defparam lut_5686.LUT_SIZE = 5;
	defparam lut_5686.mask = 32'h01000000;

	lut_sub lut_5693 ({i_28_, g57, i_22_, g549, g585}, g586);
	defparam lut_5693.LUT_SIZE = 5;
	defparam lut_5693.mask = 32'haa8aaaaa;

	lut_sub lut_5715 ({g57, i_29_, g582, g584, g586}, g587);
	defparam lut_5715.LUT_SIZE = 5;
	defparam lut_5715.mask = 32'h50504050;

	lut_sub lut_5730 ({g8, g335, g24, g581, g587}, g588);
	defparam lut_5730.LUT_SIZE = 5;
	defparam lut_5730.mask = 32'h000030b0;

	lut_sub lut_5742 ({i_9_, g570, g576, g579, g588}, g589);
	defparam lut_5742.LUT_SIZE = 5;
	defparam lut_5742.mask = 32'haaaa0200;

	lut_sub lut_5756 ({i_16_, i_33_, i_34_, g33, g34}, g590);
	defparam lut_5756.LUT_SIZE = 5;
	defparam lut_5756.mask = 32'h00010000;

	lut_sub lut_5762 ({i_33_, i_34_, i_14_, g45, g35}, g591);
	defparam lut_5762.LUT_SIZE = 5;
	defparam lut_5762.mask = 32'h00000001;

	lut_sub lut_5768 ({i_12_, i_13_, i_14_, g590, g591}, g592);
	defparam lut_5768.LUT_SIZE = 5;
	defparam lut_5768.mask = 32'ha8aaaaaa;

	lut_sub lut_5788 ({i_7_, g70, g451}, g593);
	defparam lut_5788.LUT_SIZE = 3;
	defparam lut_5788.mask = 8'h2a;

	lut_sub lut_5800 ({g66, g60, g478, g449, g535, g593}, g594);
	defparam lut_5800.LUT_SIZE = 6;
	defparam lut_5800.mask = 64'h002200220022002f;

	lut_sub lut_5815 ({i_26_, i_29_, i_22_, g478}, g595);
	defparam lut_5815.LUT_SIZE = 4;
	defparam lut_5815.mask = 16'h0b0f;

	lut_sub lut_5827 ({i_7_, i_32_, g9, g29}, g596);
	defparam lut_5827.LUT_SIZE = 4;
	defparam lut_5827.mask = 16'h7000;

	lut_sub lut_5834 ({i_28_, i_34_, i_35_, i_26_, g164}, g597);
	defparam lut_5834.LUT_SIZE = 5;
	defparam lut_5834.mask = 32'h8aaa0000;

	lut_sub lut_5848 ({i_24_, g2, g595, g596, g597}, g598);
	defparam lut_5848.LUT_SIZE = 5;
	defparam lut_5848.mask = 32'h10100010;

	lut_sub lut_5855 ({i_33_, i_34_, i_29_, g96}, g599);
	defparam lut_5855.LUT_SIZE = 4;
	defparam lut_5855.mask = 16'h4404;

	lut_sub lut_5864 ({i_33_, i_34_, g65, g121, g494}, g600);
	defparam lut_5864.LUT_SIZE = 5;
	defparam lut_5864.mask = 32'h030f0105;

	lut_sub lut_5879 ({i_26_, i_25_, g488, g599, g600}, g601);
	defparam lut_5879.LUT_SIZE = 5;
	defparam lut_5879.mask = 32'h01010100;

	lut_sub lut_5889 ({i_33_, g71, g65, g60, g449}, g602);
	defparam lut_5889.LUT_SIZE = 5;
	defparam lut_5889.mask = 32'h01000000;

	lut_sub lut_5896 ({g2, g84, g7, i_25_}, g603);
	defparam lut_5896.LUT_SIZE = 4;
	defparam lut_5896.mask = 16'h0002;

	lut_sub lut_5902 ({i_33_, g2, g1}, g604);
	defparam lut_5902.LUT_SIZE = 3;
	defparam lut_5902.mask = 8'h10;

	lut_sub lut_5909 ({i_2_, i_30_, g7, g604, g548}, g605);
	defparam lut_5909.LUT_SIZE = 5;
	defparam lut_5909.mask = 32'h07050300;

	lut_sub lut_5924 ({g2, g479, g437, g603, g605}, g606);
	defparam lut_5924.LUT_SIZE = 5;
	defparam lut_5924.mask = 32'h88888808;

	lut_sub lut_5939 ({g592, g598, g601, g602, g606}, g607);
	defparam lut_5939.LUT_SIZE = 5;
	defparam lut_5939.mask = 32'h00004000;

	lut_sub lut_5946 ({i_32_, g1, g11, g32}, g608);
	defparam lut_5946.LUT_SIZE = 4;
	defparam lut_5946.mask = 16'h0703;

	lut_sub lut_5957 ({i_33_, g2, g24, g608}, g609);
	defparam lut_5957.LUT_SIZE = 4;
	defparam lut_5957.mask = 16'h0400;

	lut_sub lut_5964 ({i_32_, g11, g32, g24}, g610);
	defparam lut_5964.LUT_SIZE = 4;
	defparam lut_5964.mask = 16'h2a0a;

	lut_sub lut_5974 ({i_34_, g1, g478}, g611);
	defparam lut_5974.LUT_SIZE = 3;
	defparam lut_5974.mask = 8'h01;

	lut_sub lut_5983 ({g82, i_25_, g451, g604, g610, g611}, g612);
	defparam lut_5983.LUT_SIZE = 6;
	defparam lut_5983.mask = 64'h005f005f33ff005f;

	lut_sub lut_6020 ({i_33_, g451, g523, g609, g612}, g613);
	defparam lut_6020.LUT_SIZE = 5;
	defparam lut_6020.mask = 32'h88808888;

	lut_sub lut_6033 ({g2, i_7_, g1, g70}, g614);
	defparam lut_6033.LUT_SIZE = 4;
	defparam lut_6033.mask = 16'h0020;

	lut_sub lut_6038 ({i_34_, i_26_, i_29_, i_22_, g494}, g615);
	defparam lut_6038.LUT_SIZE = 5;
	defparam lut_6038.mask = 32'h44005450;

	lut_sub lut_6054 ({g2, g1, g164, g486, g443, g615}, g616);
	defparam lut_6054.LUT_SIZE = 6;
	defparam lut_6054.mask = 64'h0505070705050f07;

	lut_sub lut_6080 ({i_33_, i_25_, g614, g616}, g617);
	defparam lut_6080.LUT_SIZE = 4;
	defparam lut_6080.mask = 16'h888a;

	lut_sub lut_6093 ({i_38_, g592, g594, g607, g613, g617}, g618);
	defparam lut_6093.LUT_SIZE = 6;
	defparam lut_6093.mask = 64'h0100ffff01000100;

	lut_sub lut_6118 ({g1, g541, g561}, g619);
	defparam lut_6118.LUT_SIZE = 3;
	defparam lut_6118.mask = 8'h01;

	lut_sub lut_6123 ({i_12_, i_9_, i_8_, g550}, g620);
	defparam lut_6123.LUT_SIZE = 4;
	defparam lut_6123.mask = 16'h0004;

	lut_sub lut_6132 ({g108, g164, g258, g619, g620}, g621);
	defparam lut_6132.LUT_SIZE = 5;
	defparam lut_6132.mask = 32'h80a088aa;

	lut_sub lut_6146 ({i_28_, i_22_, g672, g621}, g622);
	defparam lut_6146.LUT_SIZE = 4;
	defparam lut_6146.mask = 16'h5455;

	lut_sub lut_6158 ({i_24_, g70, g498}, g623);
	defparam lut_6158.LUT_SIZE = 3;
	defparam lut_6158.mask = 8'h2a;

	lut_sub lut_6169 ({g60, g456, g532, g577, g623}, g624);
	defparam lut_6169.LUT_SIZE = 5;
	defparam lut_6169.mask = 32'h00330a3b;

	lut_sub lut_6183 ({i_12_, i_13_, i_18_, i_19_, i_10_}, g625);
	defparam lut_6183.LUT_SIZE = 5;
	defparam lut_6183.mask = 32'h00000100;

	lut_sub lut_6191 ({i_10_, g464, g553, g569, g625}, g626);
	defparam lut_6191.LUT_SIZE = 5;
	defparam lut_6191.mask = 32'h505050dc;

	lut_sub lut_6208 ({i_34_, g1, g70, g504}, g627);
	defparam lut_6208.LUT_SIZE = 4;
	defparam lut_6208.mask = 16'h0001;

	lut_sub lut_6215 ({i_14_, g86, g143, g627}, g628);
	defparam lut_6215.LUT_SIZE = 4;
	defparam lut_6215.mask = 16'haa8a;

	lut_sub lut_6226 ({i_24_, i_28_, i_26_, g65, i_10_}, g629);
	defparam lut_6226.LUT_SIZE = 5;
	defparam lut_6226.mask = 32'h20000000;

	lut_sub lut_6233 ({i_9_, g29, g551, g629}, g630);
	defparam lut_6233.LUT_SIZE = 4;
	defparam lut_6233.mask = 16'h0001;

	lut_sub lut_6237 ({i_7_, i_3_, i_18_, i_11_, i_19_, i_8_}, g631);
	defparam lut_6237.LUT_SIZE = 6;
	defparam lut_6237.mask = 64'h2a2a000a00000000;

	lut_sub lut_6252 ({i_12_, g24, g140, g551, g631}, g632);
	defparam lut_6252.LUT_SIZE = 5;
	defparam lut_6252.mask = 32'h00000001;

	lut_sub lut_6257 ({i_12_, i_2_, i_22_, g495}, g633);
	defparam lut_6257.LUT_SIZE = 4;
	defparam lut_6257.mask = 16'h4044;

	lut_sub lut_6266 ({i_33_, g140, i_25_, g428, g633}, g634);
	defparam lut_6266.LUT_SIZE = 5;
	defparam lut_6266.mask = 32'h00110010;

	lut_sub lut_6276 ({g90, g70, g121, g634}, g635);
	defparam lut_6276.LUT_SIZE = 4;
	defparam lut_6276.mask = 16'haaa8;

	lut_sub lut_6288 ({i_12_, i_2_, g12, i_8_, g456}, g636);
	defparam lut_6288.LUT_SIZE = 5;
	defparam lut_6288.mask = 32'h40004040;

	lut_sub lut_6298 ({i_9_, g46, g474, g574, g636}, g637);
	defparam lut_6298.LUT_SIZE = 5;
	defparam lut_6298.mask = 32'h11111113;

	lut_sub lut_6313 ({i_13_, i_9_, g164, g488, g428}, g638);
	defparam lut_6313.LUT_SIZE = 5;
	defparam lut_6313.mask = 32'h00100000;

	lut_sub lut_6317 ({i_34_, i_26_, i_30_, i_29_, i_8_}, g639);
	defparam lut_6317.LUT_SIZE = 5;
	defparam lut_6317.mask = 32'h80008080;

	lut_sub lut_6323 ({i_34_, i_26_, i_32_, i_29_, i_22_}, g640);
	defparam lut_6323.LUT_SIZE = 5;
	defparam lut_6323.mask = 32'he000e0c0;

	lut_sub lut_6339 ({g371, g524, g638, g639, g640}, g641);
	defparam lut_6339.LUT_SIZE = 5;
	defparam lut_6339.mask = 32'h00000307;

	lut_sub lut_6350 ({i_33_, g486, g520, i_38_, g641}, g642);
	defparam lut_6350.LUT_SIZE = 5;
	defparam lut_6350.mask = 32'haaa8aaaa;

	lut_sub lut_6373 ({g630, g632, g635, g637, g642}, g643);
	defparam lut_6373.LUT_SIZE = 5;
	defparam lut_6373.mask = 32'h04000000;

	lut_sub lut_6380 ({i_31_, g520, g429, g455}, g644);
	defparam lut_6380.LUT_SIZE = 4;
	defparam lut_6380.mask = 16'h0100;

	lut_sub lut_6387 ({g37, g549, g543}, g645);
	defparam lut_6387.LUT_SIZE = 3;
	defparam lut_6387.mask = 8'h01;

	lut_sub lut_6394 ({i_28_, i_2_, i_22_, g197, g596, g580}, g646);
	defparam lut_6394.LUT_SIZE = 6;
	defparam lut_6394.mask = 64'h1500110000000000;

	lut_sub lut_6404 ({i_2_, i_9_, g473, g567}, g647);
	defparam lut_6404.LUT_SIZE = 4;
	defparam lut_6404.mask = 16'h0100;

	lut_sub lut_6410 ({i_27_, g71, g88, i_22_}, g648);
	defparam lut_6410.LUT_SIZE = 4;
	defparam lut_6410.mask = 16'h0020;

	lut_sub lut_6417 ({i_33_, i_14_, g121, g647, g648}, g649);
	defparam lut_6417.LUT_SIZE = 5;
	defparam lut_6417.mask = 32'h88888880;

	lut_sub lut_6432 ({g644, g645, g662, g646, g649}, g650);
	defparam lut_6432.LUT_SIZE = 5;
	defparam lut_6432.mask = 32'h40000000;

	lut_sub lut_6439 ({i_7_, i_32_, g443, g435, g580}, g651);
	defparam lut_6439.LUT_SIZE = 5;
	defparam lut_6439.mask = 32'h57000300;

	lut_sub lut_6453 ({i_33_, g71, g84, g465, g651}, g652);
	defparam lut_6453.LUT_SIZE = 5;
	defparam lut_6453.mask = 32'h07050505;

	lut_sub lut_6466 ({g2, i_29_, i_22_}, g653);
	defparam lut_6466.LUT_SIZE = 3;
	defparam lut_6466.mask = 8'h0d;

	lut_sub lut_6475 ({i_28_, i_26_, g504, g507, g653}, g654);
	defparam lut_6475.LUT_SIZE = 5;
	defparam lut_6475.mask = 32'h13110000;

	lut_sub lut_6486 ({i_10_, i_22_, g471, g652, g654}, g655);
	defparam lut_6486.LUT_SIZE = 5;
	defparam lut_6486.mask = 32'h80888888;

	lut_sub lut_6497 ({i_9_, i_3_, i_8_, g574}, g656);
	defparam lut_6497.LUT_SIZE = 4;
	defparam lut_6497.mask = 16'h0040;

	lut_sub lut_6504 ({i_3_, i_8_, i_10_, g550, g552, g656}, g657);
	defparam lut_6504.LUT_SIZE = 6;
	defparam lut_6504.mask = 64'haa80aa88aaaaaaaa;

	lut_sub lut_6535 ({i_12_, i_13_, i_11_, i_19_, g657}, g658);
	defparam lut_6535.LUT_SIZE = 5;
	defparam lut_6535.mask = 32'h00002a00;

	lut_sub lut_6546 ({g628, g643, g650, g655, g658}, g659);
	defparam lut_6546.LUT_SIZE = 5;
	defparam lut_6546.mask = 32'h00000002;

	lut_sub lut_6555 ({g618, g622, g624, g626, g659}, g660);
	defparam lut_6555.LUT_SIZE = 5;
	defparam lut_6555.mask = 32'h00000040;

	lut_sub lut_6565 ({g477, g510, g540, g566, g589, g660}, g661);
	defparam lut_6565.LUT_SIZE = 6;
	defparam lut_6565.mask = 64'h0000000000010000;

	lut_sub lut_6571 ({g663, g664}, g662);
	defparam lut_6571.LUT_SIZE = 2;
	defparam lut_6571.mask = 4'b1000;

	lut_sub lut_6577 ({g2, g665}, g663);
	defparam lut_6577.LUT_SIZE = 2;
	defparam lut_6577.mask = 4'b0100;

	lut_sub lut_6583 ({g2, g666}, g664);
	defparam lut_6583.LUT_SIZE = 2;
	defparam lut_6583.mask = 4'b0001;

	lut_sub lut_6588 ({i_31_, g669}, g665);
	defparam lut_6588.LUT_SIZE = 2;
	defparam lut_6588.mask = 4'b0001;

	lut_sub lut_6594 ({g667, g668}, g666);
	defparam lut_6594.LUT_SIZE = 2;
	defparam lut_6594.mask = 4'b1000;

	lut_sub lut_6599 ({i_31_, g670}, g667);
	defparam lut_6599.LUT_SIZE = 2;
	defparam lut_6599.mask = 4'b0100;

	lut_sub lut_6604 ({i_31_, g671}, g668);
	defparam lut_6604.LUT_SIZE = 2;
	defparam lut_6604.mask = 4'b0001;

	lut_sub lut_6610 ({g90, g71, i_28_}, g669);
	defparam lut_6610.LUT_SIZE = 3;
	defparam lut_6610.mask = 8'h08;

	lut_sub lut_6616 ({g90, i_29_, g70, i_28_}, g670);
	defparam lut_6616.LUT_SIZE = 4;
	defparam lut_6616.mask = 16'h0020;

	lut_sub lut_6622 ({g90, i_29_, g71, i_28_}, g671);
	defparam lut_6622.LUT_SIZE = 4;
	defparam lut_6622.mask = 16'h00a8;

	lut_sub lut_6630 ({g673, g674}, g672);
	defparam lut_6630.LUT_SIZE = 2;
	defparam lut_6630.mask = 4'b1000;

	lut_sub lut_6636 ({g90, g675}, g673);
	defparam lut_6636.LUT_SIZE = 2;
	defparam lut_6636.mask = 4'b0100;

	lut_sub lut_6642 ({g90, g678}, g674);
	defparam lut_6642.LUT_SIZE = 2;
	defparam lut_6642.mask = 4'b0001;

	lut_sub lut_6648 ({g676, g677}, g675);
	defparam lut_6648.LUT_SIZE = 2;
	defparam lut_6648.mask = 4'b1000;

	lut_sub lut_6653 ({i_34_, g681}, g676);
	defparam lut_6653.LUT_SIZE = 2;
	defparam lut_6653.mask = 4'b0100;

	lut_sub lut_6658 ({i_34_, g682}, g677);
	defparam lut_6658.LUT_SIZE = 2;
	defparam lut_6658.mask = 4'b0001;

	lut_sub lut_6664 ({g679, g680}, g678);
	defparam lut_6664.LUT_SIZE = 2;
	defparam lut_6664.mask = 4'b1000;

	lut_sub lut_6669 ({i_34_, g683}, g679);
	defparam lut_6669.LUT_SIZE = 2;
	defparam lut_6669.mask = 4'b0100;

	lut_sub lut_6674 ({i_34_, g684}, g680);
	defparam lut_6674.LUT_SIZE = 2;
	defparam lut_6674.mask = 4'b0001;

	lut_sub lut_6678 ({i_14_, i_33_, i_35_}, g681);
	defparam lut_6678.LUT_SIZE = 3;
	defparam lut_6678.mask = 8'h01;

	lut_sub lut_6682 ({i_14_, i_33_, i_24_}, g682);
	defparam lut_6682.LUT_SIZE = 3;
	defparam lut_6682.mask = 8'h02;

	lut_sub lut_6687 ({i_14_, i_33_, g86, i_35_}, g683);
	defparam lut_6687.LUT_SIZE = 4;
	defparam lut_6687.mask = 16'h1115;

	lut_sub lut_6695 ({i_14_, i_33_, i_24_}, g684);
	defparam lut_6695.LUT_SIZE = 3;
	defparam lut_6695.mask = 8'h02;

	lut_sub lut_6701 ({g686, g687}, g685);
	defparam lut_6701.LUT_SIZE = 2;
	defparam lut_6701.mask = 4'b1000;

	lut_sub lut_6706 ({i_33_, g688}, g686);
	defparam lut_6706.LUT_SIZE = 2;
	defparam lut_6706.mask = 4'b0100;

	lut_sub lut_6711 ({i_33_, g691}, g687);
	defparam lut_6711.LUT_SIZE = 2;
	defparam lut_6711.mask = 4'b0001;

	lut_sub lut_6717 ({g689, g690}, g688);
	defparam lut_6717.LUT_SIZE = 2;
	defparam lut_6717.mask = 4'b1000;

	lut_sub lut_6722 ({i_34_, g693}, g689);
	defparam lut_6722.LUT_SIZE = 2;
	defparam lut_6722.mask = 4'b0100;

	lut_sub lut_6727 ({i_34_, g694}, g690);
	defparam lut_6727.LUT_SIZE = 2;
	defparam lut_6727.mask = 4'b0001;

	lut_sub lut_6732 ({i_34_, g692}, g691);
	defparam lut_6732.LUT_SIZE = 2;
	defparam lut_6732.mask = 4'b0010;

	lut_sub lut_6737 ({i_34_, g695}, g692);
	defparam lut_6737.LUT_SIZE = 2;
	defparam lut_6737.mask = 4'b0001;

	lut_sub lut_6743 ({g428, g60, i_26_, i_24_}, g693);
	defparam lut_6743.LUT_SIZE = 4;
	defparam lut_6743.mask = 16'hfff7;

	lut_sub lut_6763 ({g428, g60, i_24_}, g694);
	defparam lut_6763.LUT_SIZE = 3;
	defparam lut_6763.mask = 8'hfd;

	lut_sub lut_6775 ({g428, g60, i_25_, i_24_}, g695);
	defparam lut_6775.LUT_SIZE = 4;
	defparam lut_6775.mask = 16'hfff7;

	lut_sub lut_6795 ({g475, g697}, g696);
	defparam lut_6795.LUT_SIZE = 2;
	defparam lut_6795.mask = 4'b0001;

	lut_sub lut_6801 ({g698, g699}, g697);
	defparam lut_6801.LUT_SIZE = 2;
	defparam lut_6801.mask = 4'b1000;

	lut_sub lut_6806 ({i_34_, g700}, g698);
	defparam lut_6806.LUT_SIZE = 2;
	defparam lut_6806.mask = 4'b0100;

	lut_sub lut_6811 ({i_34_, g701}, g699);
	defparam lut_6811.LUT_SIZE = 2;
	defparam lut_6811.mask = 4'b0001;

	lut_sub lut_6816 ({i_20_, g88, i_35_, i_21_}, g700);
	defparam lut_6816.LUT_SIZE = 4;
	defparam lut_6816.mask = 16'hfefc;

	lut_sub lut_6833 ({i_20_, g88, i_24_, i_21_}, g701);
	defparam lut_6833.LUT_SIZE = 4;
	defparam lut_6833.mask = 16'hfbf3;

	lut_sub lut_6851 ({g703, g704}, g702);
	defparam lut_6851.LUT_SIZE = 2;
	defparam lut_6851.mask = 4'b1000;

	lut_sub lut_6857 ({g3, g705}, g703);
	defparam lut_6857.LUT_SIZE = 2;
	defparam lut_6857.mask = 4'b0100;

	lut_sub lut_6863 ({g3, g706}, g704);
	defparam lut_6863.LUT_SIZE = 2;
	defparam lut_6863.mask = 4'b0001;

	lut_sub lut_6868 ({i_34_, g709}, g705);
	defparam lut_6868.LUT_SIZE = 2;
	defparam lut_6868.mask = 4'b0001;

	lut_sub lut_6874 ({g707, g708}, g706);
	defparam lut_6874.LUT_SIZE = 2;
	defparam lut_6874.mask = 4'b1000;

	lut_sub lut_6879 ({i_34_, g710}, g707);
	defparam lut_6879.LUT_SIZE = 2;
	defparam lut_6879.mask = 4'b0100;

	lut_sub lut_6884 ({i_34_, g711}, g708);
	defparam lut_6884.LUT_SIZE = 2;
	defparam lut_6884.mask = 4'b0001;

	lut_sub lut_6889 ({g5, i_31_, i_28_, i_21_}, g709);
	defparam lut_6889.LUT_SIZE = 4;
	defparam lut_6889.mask = 16'h0400;

	lut_sub lut_6893 ({i_31_, i_35_, i_21_}, g710);
	defparam lut_6893.LUT_SIZE = 3;
	defparam lut_6893.mask = 8'h01;

	lut_sub lut_6898 ({g5, i_31_, i_28_, i_21_}, g711);
	defparam lut_6898.LUT_SIZE = 4;
	defparam lut_6898.mask = 16'h0400;

	lut_sub lut_6903 ({i_31_, g713}, g712);
	defparam lut_6903.LUT_SIZE = 2;
	defparam lut_6903.mask = 4'b0010;

	lut_sub lut_6908 ({i_31_, g714}, g713);
	defparam lut_6908.LUT_SIZE = 2;
	defparam lut_6908.mask = 4'b0001;

	lut_sub lut_6914 ({g715, g716}, g714);
	defparam lut_6914.LUT_SIZE = 2;
	defparam lut_6914.mask = 4'b1000;

	lut_sub lut_6919 ({i_34_, g717}, g715);
	defparam lut_6919.LUT_SIZE = 2;
	defparam lut_6919.mask = 4'b0100;

	lut_sub lut_6924 ({i_34_, g718}, g716);
	defparam lut_6924.LUT_SIZE = 2;
	defparam lut_6924.mask = 4'b0001;

	lut_sub lut_6930 ({g108, g34, i_35_, i_28_}, g717);
	defparam lut_6930.LUT_SIZE = 4;
	defparam lut_6930.mask = 16'h54fc;

	lut_sub lut_6944 ({g108, g21, i_28_}, g718);
	defparam lut_6944.LUT_SIZE = 3;
	defparam lut_6944.mask = 8'h4c;


endmodule