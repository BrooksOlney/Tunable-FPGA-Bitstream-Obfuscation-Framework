module alu4x6xv (i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_3_, i_13_, i_4_, i_12_, i_1_, i_11_, i_2_, i_0_, o_1_, o_2_, o_0_, o_7_, o_5_, o_6_, o_3_, o_4_);

	input i_9_;
	input i_10_;
	input i_7_;
	input i_8_;
	input i_5_;
	input i_6_;
	input i_3_;
	input i_13_;
	input i_4_;
	input i_12_;
	input i_1_;
	input i_11_;
	input i_2_;
	input i_0_;
	output o_1_;
	output o_2_;
	output o_0_;
	output o_7_;
	output o_5_;
	output o_6_;
	output o_3_;
	output o_4_;

	wire [911 : 0] sk /* synthesis noprune */;

	lut_sub lut_3 ({sk[0], i_4_, n_n861, n_n860, x415x, x6485x}, o_1_);
	defparam lut_3.LUT_SIZE = 6;
	defparam lut_3.mask = 64'h0f3fffff7fff5fff;

	lut_sub lut_8 ({sk[1], x6530x, x6520x, n_n872, n_n879, x6513x, x6514x}, o_2_);
	defparam lut_8.LUT_SIZE = 7;
	defparam lut_8.mask = 128'h00ffffff00ffffff7fffffffffffffff;

	lut_sub lut_15 ({sk[2], x6538x, x6536x, x6537x}, o_0_);
	defparam lut_15.LUT_SIZE = 4;
	defparam lut_15.mask = 16'h777f;

	lut_sub lut_19 ({sk[3], x6829x, x6825x, x6826x, x6827x}, o_7_);
	defparam lut_19.LUT_SIZE = 5;
	defparam lut_19.mask = 32'h77ff7fff;

	lut_sub lut_24 ({sk[4], x6951x, x6869x, x6870x, x6948x}, o_5_);
	defparam lut_24.LUT_SIZE = 5;
	defparam lut_24.mask = 32'h77ff7fff;

	lut_sub lut_29 ({sk[5], n_n1185, x6975x, n_n1184, n_n1187, x6999x}, o_6_);
	defparam lut_29.LUT_SIZE = 6;
	defparam lut_29.mask = 64'h0f0f0f0f7fffffff;

	lut_sub lut_35 ({sk[6], x7076x, n_n910, n_n907, x7054x, x7055x, x7063x}, o_3_);
	defparam lut_35.LUT_SIZE = 7;
	defparam lut_35.mask = 128'h37ffffffffffffff7fffffffffffffff;

	lut_sub lut_42 ({sk[7], n_n955, n_n956, x7336x, x7337x, x7338x}, o_4_);
	defparam lut_42.LUT_SIZE = 6;
	defparam lut_42.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_48 ({sk[8], n_n665, n_n1574, x19x, x295x, x1860x, x1861x}, n_n861);
	defparam lut_48.LUT_SIZE = 7;
	defparam lut_48.mask = 128'h37ffffffffffffff777fffff77ffffff;

	lut_sub lut_54 ({sk[9], n_n761, n_n2368, x318x, x1867x, x1869x, x6474x}, n_n860);
	defparam lut_54.LUT_SIZE = 7;
	defparam lut_54.mask = 128'h37ffffffffffffff7f7fffff7fffffff;

	lut_sub lut_60 ({sk[10], i_9_, i_10_, i_8_, i_3_, i_12_, i_11_}, x415x);
	defparam lut_60.LUT_SIZE = 7;
	defparam lut_60.mask = 128'h37ffffffffffffff00c0aac000ccaacc;

	lut_sub lut_65 ({sk[11], i_9_, i_10_, i_8_, i_3_, i_4_, x6484x}, x6485x);
	defparam lut_65.LUT_SIZE = 7;
	defparam lut_65.mask = 128'h37ffffffffffffff55555d55555d5d5d;

	lut_sub lut_70 ({sk[12], x1842x, x6492x, x6497x, x6498x, x1823x, x6503x}, x6530x);
	defparam lut_70.LUT_SIZE = 7;
	defparam lut_70.mask = 128'h37ffffffffffffff7fffffffffffffff;

	lut_sub lut_77 ({sk[13], i_11_, n_n844, x74x, x665x, x1796x, x6517x}, x6520x);
	defparam lut_77.LUT_SIZE = 7;
	defparam lut_77.mask = 128'h37ffffffffffffff77777f7f77ff7fff;

	lut_sub lut_82 ({sk[14], i_5_, x6528x, x681x}, n_n872);
	defparam lut_82.LUT_SIZE = 4;
	defparam lut_82.mask = 16'h3737;

	lut_sub lut_85 ({sk[15], i_7_, n_n421, n_n197, x385x, x6508x, x6505x}, n_n879);
	defparam lut_85.LUT_SIZE = 7;
	defparam lut_85.mask = 128'h37ffffffffffffff77777f7f777f7f7f;

	lut_sub lut_90 ({sk[16], i_12_, i_0_, n_n36, x28x, x74x, x287x}, x6513x);
	defparam lut_90.LUT_SIZE = 7;
	defparam lut_90.mask = 128'h37ffffffffffffff3333333f7777777f;

	lut_sub lut_94 ({sk[17], i_12_, i_11_, x327x, n_n598, x123x, x662x}, x6514x);
	defparam lut_94.LUT_SIZE = 7;
	defparam lut_94.mask = 128'h37ffffffffffffff050537ff0505ffff;

	lut_sub lut_99 ({sk[18], i_9_, i_10_, i_8_, i_3_, i_2_, x327x}, x6538x);
	defparam lut_99.LUT_SIZE = 7;
	defparam lut_99.mask = 128'h37ffffffffffffff00005500000f7f3f;

	lut_sub lut_104 ({sk[19], i_9_, i_10_, i_6_, i_1_, x126x, x20x}, x6536x);
	defparam lut_104.LUT_SIZE = 7;
	defparam lut_104.mask = 128'h37ffffffffffffff33333f3377777f7f;

	lut_sub lut_109 ({sk[20], i_6_, i_2_, x283x, x285x, x348x, x25x}, x6537x);
	defparam lut_109.LUT_SIZE = 7;
	defparam lut_109.mask = 128'h37ffffffffffffff33337f7f33ff7fff;

	lut_sub lut_114 ({sk[21], x6704x, x6705x, x6792x, x6793x}, x6829x);
	defparam lut_114.LUT_SIZE = 5;
	defparam lut_114.mask = 32'h3f3f7fff;

	lut_sub lut_119 ({sk[22], i_10_, n_n1245, x6567x, x6806x, x1420x, x6804x}, x6825x);
	defparam lut_119.LUT_SIZE = 7;
	defparam lut_119.mask = 128'h37ffffffffffffff0fffffff7fffffff;

	lut_sub lut_125 ({sk[23], n_n1238, n_n1239, x1385x, x1402x, x6813x, x6814x}, x6826x);
	defparam lut_125.LUT_SIZE = 7;
	defparam lut_125.mask = 128'h37ffffffffffffff7fffffffffffffff;

	lut_sub lut_132 ({sk[24], x6605x, x6606x, n_n1240, n_n1241, n_n1236}, x6827x);
	defparam lut_132.LUT_SIZE = 6;
	defparam lut_132.mask = 64'h77ff77ff7fffffff;

	lut_sub lut_138 ({sk[25], n_n1119, x6937x, n_n1108, n_n1123, x6919x, x6936x}, x6951x);
	defparam lut_138.LUT_SIZE = 7;
	defparam lut_138.mask = 128'h5fffffff5fffffff7fffffffffffffff;

	lut_sub lut_145 ({sk[26], i_7_, n_n769, x45x, x295x, x1318x, x6867x}, x6869x);
	defparam lut_145.LUT_SIZE = 7;
	defparam lut_145.mask = 128'h5fffffff5fffffff777f777f777f7f7f;

	lut_sub lut_150 ({sk[27], i_6_, x6857x, x6858x, x472x, x6860x}, x6870x);
	defparam lut_150.LUT_SIZE = 6;
	defparam lut_150.mask = 64'h3333ffff5fff7fff;

	lut_sub lut_155 ({sk[28], x6833x, x6834x, x1366x, x1364x, x1365x, x6839x}, x6948x);
	defparam lut_155.LUT_SIZE = 7;
	defparam lut_155.mask = 128'h77ff77ffffffffff7fffffffffffffff;

	lut_sub lut_162 ({sk[29], i_2_, x340x, x1154x, x6966x, x1165x, x1166x}, n_n1185);
	defparam lut_162.LUT_SIZE = 7;
	defparam lut_162.mask = 128'h77ff77ffffffffff00ff00ff7fffffff;

	lut_sub lut_168 ({sk[30], i_4_, n_n816, x27x, x6969x, x6972x, x6973x}, x6975x);
	defparam lut_168.LUT_SIZE = 7;
	defparam lut_168.mask = 128'h77ff77ffffffffff7f7f7f7f7f7f7fff;

	lut_sub lut_173 ({sk[31], x6992x, x314x, x1132x, x6981x, x365x, x1107x}, n_n1184);
	defparam lut_173.LUT_SIZE = 7;
	defparam lut_173.mask = 128'h77ff77ffffffffff5fff7fffffffffff;

	lut_sub lut_179 ({sk[32], i_7_, x19x, x301x, x630x, x6996x, x6997x}, n_n1187);
	defparam lut_179.LUT_SIZE = 7;
	defparam lut_179.mask = 128'h77ff77ffffffffff777777ff5f5f5f5f;

	lut_sub lut_184 ({sk[33], n_n1189, x1169x, x6962x}, x6999x);
	defparam lut_184.LUT_SIZE = 4;
	defparam lut_184.mask = 16'h377f;

	lut_sub lut_188 ({sk[34], i_10_, x7008x, x658x, x972x, x7072x, x7073x}, x7076x);
	defparam lut_188.LUT_SIZE = 7;
	defparam lut_188.mask = 128'h77ff77ffffffffff7fffffff7f7fffff;

	lut_sub lut_194 ({sk[35], i_11_, x7018x, x7020x, x7997x}, n_n910);
	defparam lut_194.LUT_SIZE = 5;
	defparam lut_194.mask = 32'h55ffbf33;

	lut_sub lut_198 ({sk[36], x7026x, x7027x, x76x, x108x, x403x, x7040x}, n_n907);
	defparam lut_198.LUT_SIZE = 7;
	defparam lut_198.mask = 128'h77ff77ffffffffff7fffffffffffffff;

	lut_sub lut_205 ({sk[37], i_12_, x407x, x105x, x692x, x1023x}, x7054x);
	defparam lut_205.LUT_SIZE = 6;
	defparam lut_205.mask = 64'h337737777fff5fff;

	lut_sub lut_210 ({sk[38], i_12_, x694x, x7052x, x7053x, x1011x, x7048x}, x7055x);
	defparam lut_210.LUT_SIZE = 7;
	defparam lut_210.mask = 128'h77ff77ffffffffff7fffffff77777777;

	lut_sub lut_216 ({sk[39], x41x, x382x, x1076x, x1075x, x7060x, x7061x}, x7063x);
	defparam lut_216.LUT_SIZE = 7;
	defparam lut_216.mask = 128'h77ff77ffffffffff7fff7fff7fffffff;

	lut_sub lut_222 ({sk[40], n_n991, x7198x, x7232x, x7233x, x7242x, x7243x}, n_n955);
	defparam lut_222.LUT_SIZE = 7;
	defparam lut_222.mask = 128'h77ff77ffffffffff7fffffffffffffff;

	lut_sub lut_229 ({sk[41], x7262x, x7263x, x7310x, x7311x, x7318x, x7319x}, n_n956);
	defparam lut_229.LUT_SIZE = 7;
	defparam lut_229.mask = 128'h77ff77ffffffffff7fffffffffffffff;

	lut_sub lut_236 ({sk[42], x7118x, x7107x, x896x, x920x, x7106x, x7333x}, x7336x);
	defparam lut_236.LUT_SIZE = 7;
	defparam lut_236.mask = 128'h77ff77ffffffffff7fffffffffffffff;

	lut_sub lut_243 ({sk[43], n_n972, x7169x, n_n977, n_n984, n_n983}, x7337x);
	defparam lut_243.LUT_SIZE = 6;
	defparam lut_243.mask = 64'h337737777fffffff;

	lut_sub lut_249 ({sk[44], x7151x, n_n957, n_n981, x7149x, x7332x}, x7338x);
	defparam lut_249.LUT_SIZE = 6;
	defparam lut_249.mask = 64'h337737777fffffff;

	lut_sub lut_255 ({sk[45], i_13_, i_12_}, n_n665);
	defparam lut_255.LUT_SIZE = 3;
	defparam lut_255.mask = 8'h32;

	lut_sub lut_257 ({sk[46], i_9_, i_10_, i_13_, i_12_, i_11_}, n_n1574);
	defparam lut_257.LUT_SIZE = 6;
	defparam lut_257.mask = 64'h3377377700000008;

	lut_sub lut_259 ({sk[47], i_8_, i_3_}, x19x);
	defparam lut_259.LUT_SIZE = 3;
	defparam lut_259.mask = 8'h32;

	lut_sub lut_261 ({sk[48], i_13_, i_4_, i_12_}, x295x);
	defparam lut_261.LUT_SIZE = 4;
	defparam lut_261.mask = 16'h3710;

	lut_sub lut_263 ({sk[49], i_3_, i_13_, i_4_, i_12_, i_11_}, x1860x);
	defparam lut_263.LUT_SIZE = 6;
	defparam lut_263.mask = 64'h3377377701880000;

	lut_sub lut_266 ({sk[50], i_9_, i_10_, i_8_, i_3_, i_13_, i_11_}, x1861x);
	defparam lut_266.LUT_SIZE = 7;
	defparam lut_266.mask = 128'h77ff77ffffffffff0000230000032303;

	lut_sub lut_270 ({sk[51], i_7_, i_5_, x33x, n_n36, n_n197, x6490x}, x1842x);
	defparam lut_270.LUT_SIZE = 7;
	defparam lut_270.mask = 128'h77ff77ffffffffff555f0000557f0000;

	lut_sub lut_274 ({sk[52], i_7_, i_5_, x33x, n_n35, x647x, x1840x}, x6492x);
	defparam lut_274.LUT_SIZE = 7;
	defparam lut_274.mask = 128'h77ff77ffffffffff7777555f5555555f;

	lut_sub lut_278 ({sk[53], i_1_, x12x, n_n183, x34x, n_n35, x6496x}, x6497x);
	defparam lut_278.LUT_SIZE = 7;
	defparam lut_278.mask = 128'h77ff77ffffffffff55555555575757ff;

	lut_sub lut_282 ({sk[54], i_2_, x12x, n_n432, n_n35, x316x, x1833x}, x6498x);
	defparam lut_282.LUT_SIZE = 7;
	defparam lut_282.mask = 128'h77ff77ffffffffff5555555555557fff;

	lut_sub lut_287 ({sk[55], i_6_, i_0_, x652x}, x1823x);
	defparam lut_287.LUT_SIZE = 4;
	defparam lut_287.mask = 16'h3701;

	lut_sub lut_289 ({sk[56], i_11_, n_n818, x181x, x384x, x1826x, x6500x}, x6503x);
	defparam lut_289.LUT_SIZE = 7;
	defparam lut_289.mask = 128'h77ff77ffffffffff7777ff777f7fff7f;

	lut_sub lut_294 ({sk[57], i_6_, i_3_, i_2_, i_0_}, x327x);
	defparam lut_294.LUT_SIZE = 5;
	defparam lut_294.mask = 32'h55ff0100;

	lut_sub lut_296 ({sk[58], n_n1250, n_n1256, x6658x, x1609x, x1610x, x6667x}, x6704x);
	defparam lut_296.LUT_SIZE = 7;
	defparam lut_296.mask = 128'h77ff77ffffffffff7fffffffffffffff;

	lut_sub lut_303 ({sk[59], n_n1248, x6695x, x1547x, x1564x, x6691x, x6692x}, x6705x);
	defparam lut_303.LUT_SIZE = 7;
	defparam lut_303.mask = 128'h77ff77ffffffffff7fffffffffffffff;

	lut_sub lut_310 ({sk[60], x1511x, x1512x, x6737x, x6791x}, x6792x);
	defparam lut_310.LUT_SIZE = 5;
	defparam lut_310.mask = 32'h55ff7fff;

	lut_sub lut_315 ({sk[61], x6760x, n_n1265, x6782x, x7982x}, x6793x);
	defparam lut_315.LUT_SIZE = 5;
	defparam lut_315.mask = 32'h55ffbfff;

	lut_sub lut_320 ({sk[62], i_1_, x1353x, x387x, x1350x, x6849x}, n_n1119);
	defparam lut_320.LUT_SIZE = 6;
	defparam lut_320.mask = 64'h3377377777ff7fff;

	lut_sub lut_325 ({sk[63], n_n1126, x1294x, x6882x, x1283x, x6890x, x6935x}, x6937x);
	defparam lut_325.LUT_SIZE = 7;
	defparam lut_325.mask = 128'h0f0fffffffffffff7fffffffffffffff;

	lut_sub lut_332 ({sk[64], i_6_, x526x, x6941x, x634x, x6946x}, n_n1108);
	defparam lut_332.LUT_SIZE = 6;
	defparam lut_332.mask = 64'h333fffff7fff5f5f;

	lut_sub lut_337 ({sk[65], i_6_, x508x, x6903x, x6904x}, n_n1123);
	defparam lut_337.LUT_SIZE = 5;
	defparam lut_337.mask = 32'h5f5f7f77;

	lut_sub lut_341 ({sk[66], n_n638, x511x, x6910x, x6909x, x6916x, x6917x}, x6919x);
	defparam lut_341.LUT_SIZE = 7;
	defparam lut_341.mask = 128'h0f0fffffffffffff7fff7fff7fffffff;

	lut_sub lut_347 ({sk[67], i_6_, x1268x, x6896x, x554x, x1220x, x6926x}, x6936x);
	defparam lut_347.LUT_SIZE = 7;
	defparam lut_347.mask = 128'h0f0fffffffffffff7fffffff77ffffff;

	lut_sub lut_353 ({sk[68], i_3_, i_4_, n_n792, n_n835, n_n791, x109x}, x7008x);
	defparam lut_353.LUT_SIZE = 7;
	defparam lut_353.mask = 128'h0f0fffffffffffff55775f7f55775577;

	lut_sub lut_357 ({sk[69], n_n675, x35x, x30x, n_n685, x1089x, x7972x}, x658x);
	defparam lut_357.LUT_SIZE = 7;
	defparam lut_357.mask = 128'h0f0fffffffffffffbbbfbbbfbbbfffff;

	lut_sub lut_362 ({sk[70], i_9_, i_12_, i_11_, i_2_, x12x, x979x}, x972x);
	defparam lut_362.LUT_SIZE = 7;
	defparam lut_362.mask = 128'h0f0fffffffffffff7555555500000000;

	lut_sub lut_365 ({sk[71], i_8_, i_12_, i_11_, n_n658, x267x, x274x}, x7072x);
	defparam lut_365.LUT_SIZE = 7;
	defparam lut_365.mask = 128'h0f0fffffffffffff5500550003030000;

	lut_sub lut_368 ({sk[72], i_6_, i_1_, n_n741, n_n792, x35x, x7071x}, x7073x);
	defparam lut_368.LUT_SIZE = 7;
	defparam lut_368.mask = 128'h0f0fffffffffffff57ff555557575555;

	lut_sub lut_372 ({sk[73], i_13_, i_11_}, n_n637);
	defparam lut_372.LUT_SIZE = 3;
	defparam lut_372.mask = 8'h52;

	lut_sub lut_374 ({sk[74], i_13_, i_12_}, n_n761);
	defparam lut_374.LUT_SIZE = 3;
	defparam lut_374.mask = 8'h54;

	lut_sub lut_376 ({sk[75], i_9_, i_10_, i_13_, i_4_, i_12_, i_11_}, n_n2368);
	defparam lut_376.LUT_SIZE = 7;
	defparam lut_376.mask = 128'h0f0fffffffffffff0100000000000000;

	lut_sub lut_378 ({sk[76], i_9_, i_8_, i_4_}, x318x);
	defparam lut_378.LUT_SIZE = 4;
	defparam lut_378.mask = 16'h3710;

	lut_sub lut_380 ({sk[77], i_9_, i_10_, i_8_, i_3_, i_13_, i_4_}, x1867x);
	defparam lut_380.LUT_SIZE = 7;
	defparam lut_380.mask = 128'h0f0fffffffffffff0404000404000000;

	lut_sub lut_384 ({sk[78], i_10_, i_8_, i_13_, i_4_, i_11_}, x1869x);
	defparam lut_384.LUT_SIZE = 6;
	defparam lut_384.mask = 64'h333fffff10000000;

	lut_sub lut_386 ({sk[79], i_8_, i_3_, i_13_, i_4_, i_12_, i_11_}, x6474x);
	defparam lut_386.LUT_SIZE = 7;
	defparam lut_386.mask = 128'h0f0fffffffffffffa5a0000080800000;

	lut_sub lut_390 ({sk[80], i_9_, i_10_}, x8x);
	defparam lut_390.LUT_SIZE = 3;
	defparam lut_390.mask = 8'h51;

	lut_sub lut_392 ({sk[81], i_1_, i_2_}, x33x);
	defparam lut_392.LUT_SIZE = 3;
	defparam lut_392.mask = 8'h51;

	lut_sub lut_394 ({sk[82], i_8_, i_11_}, n_n36);
	defparam lut_394.LUT_SIZE = 3;
	defparam lut_394.mask = 8'h54;

	lut_sub lut_396 ({sk[83], i_9_, i_11_}, n_n197);
	defparam lut_396.LUT_SIZE = 3;
	defparam lut_396.mask = 8'h51;

	lut_sub lut_398 ({sk[84], i_9_, i_10_, i_3_, i_1_, i_11_, i_2_}, x6490x);
	defparam lut_398.LUT_SIZE = 7;
	defparam lut_398.mask = 128'h0f0fffffffffffff0001000100010303;

	lut_sub lut_401 ({sk[85], i_8_, i_12_}, n_n35);
	defparam lut_401.LUT_SIZE = 3;
	defparam lut_401.mask = 8'h51;

	lut_sub lut_403 ({sk[86], i_10_, i_8_, i_3_, i_1_, i_11_, i_2_}, x647x);
	defparam lut_403.LUT_SIZE = 7;
	defparam lut_403.mask = 128'h0f0fffffffffffff0303000303030103;

	lut_sub lut_407 ({sk[87], i_9_, i_5_, i_6_, i_1_, i_11_}, x1840x);
	defparam lut_407.LUT_SIZE = 6;
	defparam lut_407.mask = 64'h333fffff00000100;

	lut_sub lut_409 ({sk[88], i_5_, i_6_}, x12x);
	defparam lut_409.LUT_SIZE = 3;
	defparam lut_409.mask = 8'h51;

	lut_sub lut_411 ({sk[89], i_9_, i_12_}, n_n183);
	defparam lut_411.LUT_SIZE = 3;
	defparam lut_411.mask = 8'h51;

	lut_sub lut_413 ({sk[90], i_7_, i_5_}, x34x);
	defparam lut_413.LUT_SIZE = 3;
	defparam lut_413.mask = 8'h51;

	lut_sub lut_415 ({sk[91], i_5_, i_12_, i_1_, i_2_, n_n633, x316x}, x6496x);
	defparam lut_415.LUT_SIZE = 7;
	defparam lut_415.mask = 128'h0f0fffffffffffff0000030300050307;

	lut_sub lut_418 ({sk[92], i_9_, i_10_, i_12_}, n_n432);
	defparam lut_418.LUT_SIZE = 4;
	defparam lut_418.mask = 16'h3701;

	lut_sub lut_420 ({sk[93], i_10_, i_7_, i_12_}, x316x);
	defparam lut_420.LUT_SIZE = 4;
	defparam lut_420.mask = 16'h3704;

	lut_sub lut_422 ({sk[94], i_7_, i_8_, i_5_, i_6_, i_3_, i_12_}, x1833x);
	defparam lut_422.LUT_SIZE = 7;
	defparam lut_422.mask = 128'h0f0fffffffffffff0000000000010005;

	lut_sub lut_425 ({sk[95], i_10_, i_7_, i_8_, i_3_, i_12_, i_2_}, x652x);
	defparam lut_425.LUT_SIZE = 7;
	defparam lut_425.mask = 128'h0f0fffffffffffff0011033311110333;

	lut_sub lut_430 ({sk[96], i_3_, i_2_, i_0_}, n_n818);
	defparam lut_430.LUT_SIZE = 4;
	defparam lut_430.mask = 16'h3701;

	lut_sub lut_432 ({sk[97], i_6_, i_12_}, x181x);
	defparam lut_432.LUT_SIZE = 3;
	defparam lut_432.mask = 8'h5e;

	lut_sub lut_435 ({sk[98], i_5_, i_6_, i_3_, i_2_}, x384x);
	defparam lut_435.LUT_SIZE = 5;
	defparam lut_435.mask = 32'h5f5f1000;

	lut_sub lut_437 ({sk[99], i_10_, i_5_, i_6_, i_1_, i_11_}, x1826x);
	defparam lut_437.LUT_SIZE = 6;
	defparam lut_437.mask = 64'h333fffff00001000;

	lut_sub lut_439 ({sk[100], i_12_, i_2_, i_0_, n_n36, n_n358, x11x}, x6500x);
	defparam lut_439.LUT_SIZE = 7;
	defparam lut_439.mask = 128'h0f0fffffffffffff0000050500000537;

	lut_sub lut_442 ({sk[101], i_1_, i_2_, i_0_}, n_n844);
	defparam lut_442.LUT_SIZE = 4;
	defparam lut_442.mask = 16'h3701;

	lut_sub lut_444 ({sk[102], i_7_, i_8_, i_12_, i_1_, i_0_}, x74x);
	defparam lut_444.LUT_SIZE = 6;
	defparam lut_444.mask = 64'h333fffff00000001;

	lut_sub lut_446 ({sk[103], i_9_, i_10_, i_7_, i_8_, i_12_, i_11_}, x665x);
	defparam lut_446.LUT_SIZE = 7;
	defparam lut_446.mask = 128'h0f0fffffffffffff5353ff5353ffffff;

	lut_sub lut_451 ({sk[104], i_7_, i_8_, i_3_, i_1_, i_11_, i_0_}, x1796x);
	defparam lut_451.LUT_SIZE = 7;
	defparam lut_451.mask = 128'h0f0fffffffffffff0101000100000000;

	lut_sub lut_454 ({sk[105], i_10_, i_6_, i_3_, i_1_, i_2_, i_0_}, x6517x);
	defparam lut_454.LUT_SIZE = 7;
	defparam lut_454.mask = 128'h0f0fffffffffffff0001000105050001;

	lut_sub lut_457 ({sk[106], i_10_, i_12_}, n_n318);
	defparam lut_457.LUT_SIZE = 3;
	defparam lut_457.mask = 8'h51;

	lut_sub lut_459 ({sk[107], i_7_, i_5_, i_3_, i_12_, i_1_}, x1786x);
	defparam lut_459.LUT_SIZE = 6;
	defparam lut_459.mask = 64'h333fffff00000001;

	lut_sub lut_461 ({sk[108], i_7_, i_5_, i_1_, i_11_, i_2_, n_n183}, x6527x);
	defparam lut_461.LUT_SIZE = 7;
	defparam lut_461.mask = 128'h0f0fffffffffffff0000000000000015;

	lut_sub lut_464 ({sk[109], i_5_, i_6_, i_1_, n_n318, x1786x, x6527x}, x6528x);
	defparam lut_464.LUT_SIZE = 7;
	defparam lut_464.mask = 128'h0f0fffffffffffff77777777777f7777;

	lut_sub lut_468 ({sk[110], i_12_, i_1_, n_n638, n_n358, n_n432, x6525x}, x681x);
	defparam lut_468.LUT_SIZE = 7;
	defparam lut_468.mask = 128'h0f0fffffffffffff0000333355557fff;

	lut_sub lut_473 ({sk[111], i_9_, i_8_}, x18x);
	defparam lut_473.LUT_SIZE = 3;
	defparam lut_473.mask = 8'h51;

	lut_sub lut_475 ({sk[112], i_10_, i_8_, i_3_}, x126x);
	defparam lut_475.LUT_SIZE = 4;
	defparam lut_475.mask = 16'h3704;

	lut_sub lut_477 ({sk[113], i_9_, i_1_}, x283x);
	defparam lut_477.LUT_SIZE = 3;
	defparam lut_477.mask = 8'h51;

	lut_sub lut_479 ({sk[114], i_10_, i_7_}, x285x);
	defparam lut_479.LUT_SIZE = 3;
	defparam lut_479.mask = 8'h52;

	lut_sub lut_481 ({sk[115], i_5_, i_0_}, x20x);
	defparam lut_481.LUT_SIZE = 3;
	defparam lut_481.mask = 8'h51;

	lut_sub lut_483 ({sk[116], i_9_, i_5_, i_0_}, x343x);
	defparam lut_483.LUT_SIZE = 4;
	defparam lut_483.mask = 16'h3701;

	lut_sub lut_485 ({sk[117], i_5_, i_0_}, x16x);
	defparam lut_485.LUT_SIZE = 3;
	defparam lut_485.mask = 8'h54;

	lut_sub lut_487 ({sk[118], i_10_, i_5_, i_0_}, x348x);
	defparam lut_487.LUT_SIZE = 4;
	defparam lut_487.mask = 16'h3704;

	lut_sub lut_489 ({sk[119], i_9_, i_7_}, x25x);
	defparam lut_489.LUT_SIZE = 3;
	defparam lut_489.mask = 8'h51;

	lut_sub lut_491 ({sk[120], i_9_, i_7_, i_2_}, x386x);
	defparam lut_491.LUT_SIZE = 4;
	defparam lut_491.mask = 16'h3701;

	lut_sub lut_493 ({sk[121], i_1_, i_0_}, x264x);
	defparam lut_493.LUT_SIZE = 3;
	defparam lut_493.mask = 8'h51;

	lut_sub lut_495 ({sk[122], i_9_, n_n541, n_n746, n_n729, x329x, x6549x}, x1771x);
	defparam lut_495.LUT_SIZE = 7;
	defparam lut_495.mask = 128'h0f0fffffffffffff000011110000111f;

	lut_sub lut_498 ({sk[123], n_n538, n_n453, x341x, n_n575, n_n756, x424x}, x6551x);
	defparam lut_498.LUT_SIZE = 7;
	defparam lut_498.mask = 128'h0f0fffffffffffff0003000300035557;

	lut_sub lut_501 ({sk[124], i_9_, n_n835, n_n748, n_n725, x390x, x7991x}, x1765x);
	defparam lut_501.LUT_SIZE = 7;
	defparam lut_501.mask = 128'h0f0fffffffffffff000000000a0a0a3b;

	lut_sub lut_504 ({sk[125], n_n498, n_n835, n_n725, x341x, x6540x, x6542x}, x6552x);
	defparam lut_504.LUT_SIZE = 7;
	defparam lut_504.mask = 128'h0f0fffffffffffff0003000300035557;

	lut_sub lut_507 ({sk[126], i_2_, x264x, x1771x, x6551x, x1765x, x6552x}, n_n1238);
	defparam lut_507.LUT_SIZE = 7;
	defparam lut_507.mask = 128'h0f0fffffffffffff77777fff77777777;

	lut_sub lut_512 ({sk[127], i_9_, i_10_, i_8_, i_13_, i_11_}, x337x);
	defparam lut_512.LUT_SIZE = 6;
	defparam lut_512.mask = 64'h333fffff00000020;

	lut_sub lut_514 ({sk[128], x12x, n_n665, n_n609, x36x, x433x, x6559x}, x1745x);
	defparam lut_514.LUT_SIZE = 7;
	defparam lut_514.mask = 128'h0f0fffffffffffff0000053700005577;

	lut_sub lut_518 ({sk[129], i_7_, i_5_, i_1_, i_0_, x337x, x1745x}, n_n1245);
	defparam lut_518.LUT_SIZE = 7;
	defparam lut_518.mask = 128'h0f0fffffffffffff5577555755555555;

	lut_sub lut_522 ({sk[130], i_7_, i_6_, i_1_, i_0_, n_n623, n_n619}, x1757x);
	defparam lut_522.LUT_SIZE = 7;
	defparam lut_522.mask = 128'h0f0fffffffffffff0000000030053535;

	lut_sub lut_527 ({sk[131], x12x, n_n638, n_n844, n_n619, n_n612, x1755x}, x6556x);
	defparam lut_527.LUT_SIZE = 7;
	defparam lut_527.mask = 128'h0f0fffffffffffff575f575f575fffff;

	lut_sub lut_532 ({sk[132], i_9_, i_7_, i_8_, i_13_, i_11_}, x353x);
	defparam lut_532.LUT_SIZE = 6;
	defparam lut_532.mask = 64'h333fffff00000200;

	lut_sub lut_534 ({sk[133], i_7_, i_5_, i_1_, n_n623, n_n619, x436x}, x435x);
	defparam lut_534.LUT_SIZE = 7;
	defparam lut_534.mask = 128'h0f0fffffffffffff0505050505050537;

	lut_sub lut_537 ({sk[134], i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x434x);
	defparam lut_537.LUT_SIZE = 7;
	defparam lut_537.mask = 128'h0f0fffffffffffff0000000800000004;

	lut_sub lut_540 ({sk[135], n_n665, x1757x, x6556x, x353x, x435x, x434x}, x6567x);
	defparam lut_540.LUT_SIZE = 7;
	defparam lut_540.mask = 128'h0f0fffffffffffff0505050537ffffff;

	lut_sub lut_545 ({sk[136], i_9_, i_7_, i_8_}, n_n638);
	defparam lut_545.LUT_SIZE = 4;
	defparam lut_545.mask = 16'h3701;

	lut_sub lut_547 ({sk[137], i_10_, i_6_, n_n541, n_n852, x301x, x329x}, x1727x);
	defparam lut_547.LUT_SIZE = 7;
	defparam lut_547.mask = 128'h0f0fffffffffffff0037000500050005;

	lut_sub lut_550 ({sk[138], n_n835, n_n847, n_n197, n_n752, n_n756, x302x}, x1722x);
	defparam lut_550.LUT_SIZE = 7;
	defparam lut_550.mask = 128'h0f0fffffffffffff0000000500110015;

	lut_sub lut_553 ({sk[139], i_6_, i_1_, i_2_, i_0_, x6573x}, x1729x);
	defparam lut_553.LUT_SIZE = 6;
	defparam lut_553.mask = 64'h333fffff00000004;

	lut_sub lut_555 ({sk[140], i_5_, i_6_, i_12_, x294x, x272x, x298x}, x6574x);
	defparam lut_555.LUT_SIZE = 7;
	defparam lut_555.mask = 128'h0f0fffffffffffff0000050500003300;

	lut_sub lut_558 ({sk[141], i_9_, n_n538, n_n844, n_n752, n_n840, x6568x}, x6576x);
	defparam lut_558.LUT_SIZE = 7;
	defparam lut_558.mask = 128'h0f0fffffffffffff010101010101010f;

	lut_sub lut_561 ({sk[142], n_n638, x1727x, x1722x, x1729x, x6574x, x6576x}, n_n1239);
	defparam lut_561.LUT_SIZE = 7;
	defparam lut_561.mask = 128'h0f0fffffffffffff55ff55ff7fffffff;

	lut_sub lut_567 ({sk[143], i_0_, x337x, x28x, n_n598, x385x, x42x}, x1701x);
	defparam lut_567.LUT_SIZE = 7;
	defparam lut_567.mask = 128'h0f0fffffffffffff00007f7f00007fff;

	lut_sub lut_572 ({sk[144], i_13_, i_12_, x1702x, n_n597, x6590x, x7980x}, x6593x);
	defparam lut_572.LUT_SIZE = 7;
	defparam lut_572.mask = 128'h0f0fffffffffffffaaaaaaaaabffaaaa;

	lut_sub lut_576 ({sk[145], i_10_, n_n570, n_n844, x282x, x391x, x6596x}, x6604x);
	defparam lut_576.LUT_SIZE = 7;
	defparam lut_576.mask = 128'h0f0fffffffffffff0505053705050505;

	lut_sub lut_579 ({sk[146], x1701x, x6593x, x6604x}, x6605x);
	defparam lut_579.LUT_SIZE = 4;
	defparam lut_579.mask = 16'h377f;

	lut_sub lut_583 ({sk[147], i_9_, i_7_, i_8_}, n_n581);
	defparam lut_583.LUT_SIZE = 4;
	defparam lut_583.mask = 16'h3708;

	lut_sub lut_585 ({sk[148], i_10_, i_7_, i_8_, n_n665, x462x, x461x}, x1710x);
	defparam lut_585.LUT_SIZE = 7;
	defparam lut_585.mask = 128'h0f0fffffffffffff0000000003000500;

	lut_sub lut_588 ({sk[149], i_13_, n_n844, n_n1574, x6583x, x7979x}, x6587x);
	defparam lut_588.LUT_SIZE = 6;
	defparam lut_588.mask = 64'h333fffffafafafbf;

	lut_sub lut_592 ({sk[150], i_8_, x25x, n_n653, x469x, x6601x, x7978x}, x6603x);
	defparam lut_592.LUT_SIZE = 7;
	defparam lut_592.mask = 128'h0f0fffffffffffffaabbafbfaabbaabb;

	lut_sub lut_596 ({sk[151], i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x467x);
	defparam lut_596.LUT_SIZE = 7;
	defparam lut_596.mask = 128'h0f0fffffffffffff0000080040000400;

	lut_sub lut_600 ({sk[152], n_n637, n_n581, x1710x, x6587x, x6603x, x467x}, x6606x);
	defparam lut_600.LUT_SIZE = 7;
	defparam lut_600.mask = 128'h0f0fffffffffffff0fff0fff3fff7fff;

	lut_sub lut_605 ({sk[153], i_13_, i_12_, i_11_}, n_n545);
	defparam lut_605.LUT_SIZE = 4;
	defparam lut_605.mask = 16'h3740;

	lut_sub lut_607 ({sk[154], i_5_, n_n748, x409x, x277x, x484x, x6613x}, x483x);
	defparam lut_607.LUT_SIZE = 7;
	defparam lut_607.mask = 128'h0f0fffffffffffff000f333f05053737;

	lut_sub lut_611 ({sk[155], i_9_, i_11_, n_n761, n_n538, n_n847, n_n756}, x1672x);
	defparam lut_611.LUT_SIZE = 7;
	defparam lut_611.mask = 128'h0f0fffffffffffff0000000000010000;

	lut_sub lut_613 ({sk[156], x341x, n_n752, n_n852, n_n575, n_n756, n_n729}, x1674x);
	defparam lut_613.LUT_SIZE = 7;
	defparam lut_613.mask = 128'h0f0fffffffffffff000000000011001f;

	lut_sub lut_616 ({sk[157], n_n835, n_n545, x391x, n_n550, n_n732, x6609x}, x6615x);
	defparam lut_616.LUT_SIZE = 7;
	defparam lut_616.mask = 128'h0f0fffffffffffff01010101010101ff;

	lut_sub lut_619 ({sk[158], i_9_, n_n545, x483x, x1672x, x1674x, x6615x}, n_n1240);
	defparam lut_619.LUT_SIZE = 7;
	defparam lut_619.mask = 128'h0f0fffffffffffff7f7f7fff7f7f7f7f;

	lut_sub lut_624 ({sk[159], i_4_, i_2_}, x14x);
	defparam lut_624.LUT_SIZE = 3;
	defparam lut_624.mask = 8'h54;

	lut_sub lut_626 ({sk[160], i_9_, i_10_, i_13_, i_12_, i_11_}, x282x);
	defparam lut_626.LUT_SIZE = 6;
	defparam lut_626.mask = 64'h333fffff40000000;

	lut_sub lut_628 ({sk[161], i_8_, i_5_, i_6_, i_3_}, x317x);
	defparam lut_628.LUT_SIZE = 5;
	defparam lut_628.mask = 32'h5f5f0080;

	lut_sub lut_630 ({sk[162], i_8_, i_5_, i_3_, i_4_, i_1_, i_0_}, x503x);
	defparam lut_630.LUT_SIZE = 7;
	defparam lut_630.mask = 128'h0f0fffffffffffff0000000030001000;

	lut_sub lut_633 ({sk[163], i_5_, i_0_, n_n746, x19x, n_n346, x277x}, x7977x);
	defparam lut_633.LUT_SIZE = 7;
	defparam lut_633.mask = 128'h0f0ffffffffffffffcfcfca8ffffffaa;

	lut_sub lut_643 ({sk[164], i_7_, x14x, x282x, x317x, x503x, x7977x}, x1662x);
	defparam lut_643.LUT_SIZE = 7;
	defparam lut_643.mask = 128'h0f0fffffffffffff00bb00bf00aa00af;

	lut_sub lut_647 ({sk[165], i_9_, i_10_, i_8_, i_3_, i_12_}, x105x);
	defparam lut_647.LUT_SIZE = 6;
	defparam lut_647.mask = 64'h333fffff08000000;

	lut_sub lut_649 ({sk[166], i_8_, x268x, x391x, x284x, x294x, x501x}, x6626x);
	defparam lut_649.LUT_SIZE = 7;
	defparam lut_649.mask = 128'h0f0fffffffffffff0033003300330537;

	lut_sub lut_652 ({sk[167], i_13_, i_4_, x1662x, n_n844, x105x, x6626x}, n_n1241);
	defparam lut_652.LUT_SIZE = 7;
	defparam lut_652.mask = 128'h0f0fffffffffffff57ff55ff55ff55ff;

	lut_sub lut_656 ({sk[168], i_11_, x1637x, x1638x, x6641x}, n_n1250);
	defparam lut_656.LUT_SIZE = 5;
	defparam lut_656.mask = 32'h5f5f7f55;

	lut_sub lut_660 ({sk[169], i_9_, n_n716, n_n732, n_n837, x519x, x6651x}, n_n1256);
	defparam lut_660.LUT_SIZE = 7;
	defparam lut_660.mask = 128'h0f0fffffffffffff5577557f55775577;

	lut_sub lut_664 ({sk[170], n_n835, n_n712, n_n755, n_n837, x6650x, x542x}, x6658x);
	defparam lut_664.LUT_SIZE = 7;
	defparam lut_664.mask = 128'h0f0fffffffffffff0000005503030357;

	lut_sub lut_667 ({sk[171], n_n725, n_n840, n_n755, n_n837, n_n710, x6655x}, x1609x);
	defparam lut_667.LUT_SIZE = 7;
	defparam lut_667.mask = 128'h0f0fffffffffffff0000000305050507;

	lut_sub lut_670 ({sk[172], n_n725, n_n847, n_n832, n_n755, n_n710, x541x}, x1610x);
	defparam lut_670.LUT_SIZE = 7;
	defparam lut_670.mask = 128'h0f0fffffffffffff0000000300550057;

	lut_sub lut_673 ({sk[173], n_n844, x1604x, x6663x, x1596x, x6665x}, x6667x);
	defparam lut_673.LUT_SIZE = 6;
	defparam lut_673.mask = 64'h333fffff77777fff;

	lut_sub lut_678 ({sk[174], x285x, n_n665, x353x, x455x, x453x, x1649x}, n_n1248);
	defparam lut_678.LUT_SIZE = 7;
	defparam lut_678.mask = 128'h0f0fffffffffffff5577557755775f7f;

	lut_sub lut_682 ({sk[175], x1584x, x1570x, x6676x, x6677x, x6681x, x6682x}, x6695x);
	defparam lut_682.LUT_SIZE = 7;
	defparam lut_682.mask = 128'h0f0fffffffffffff7fffffffffffffff;

	lut_sub lut_689 ({sk[176], i_13_, i_12_, x1555x, x6702x}, x1547x);
	defparam lut_689.LUT_SIZE = 5;
	defparam lut_689.mask = 32'h5f5f0070;

	lut_sub lut_692 ({sk[177], n_n853, x117x, x398x, x401x, x108x, x403x}, x1564x);
	defparam lut_692.LUT_SIZE = 7;
	defparam lut_692.mask = 128'h0f0fffffffffffff000000007fffffff;

	lut_sub lut_698 ({sk[178], i_9_, i_7_, x313x, n_n678, n_n685, x6684x}, x6691x);
	defparam lut_698.LUT_SIZE = 7;
	defparam lut_698.mask = 128'h0f0fffffffffffff0505053705050505;

	lut_sub lut_701 ({sk[179], i_3_, x274x, x17x, n_n822, x24x, n_n838}, x6692x);
	defparam lut_701.LUT_SIZE = 7;
	defparam lut_701.mask = 128'h0f0fffffffffffff010101ff000000ff;

	lut_sub lut_704 ({sk[180], i_9_, i_5_, i_6_, x27x, n_n498, x298x}, x1534x);
	defparam lut_704.LUT_SIZE = 7;
	defparam lut_704.mask = 128'h0f0fffffffffffff0000010000000000;

	lut_sub lut_706 ({sk[181], i_10_, i_11_, n_n850, n_n550, x569x, x6709x}, x1535x);
	defparam lut_706.LUT_SIZE = 7;
	defparam lut_706.mask = 128'h0f0fffffffffffff0000000011150005;

	lut_sub lut_709 ({sk[182], n_n538, n_n498, n_n847, n_n843, x302x, x6710x}, x1536x);
	defparam lut_709.LUT_SIZE = 7;
	defparam lut_709.mask = 128'h0f0fffffffffffff001100110011001f;

	lut_sub lut_712 ({sk[183], i_13_, i_12_, n_n633, x314x, x1540x, x1541x}, x1537x);
	defparam lut_712.LUT_SIZE = 7;
	defparam lut_712.mask = 128'h0f0fffffffffffff00000000777f0000;

	lut_sub lut_716 ({sk[184], x1534x, x1535x, x1536x, x1537x}, n_n1236);
	defparam lut_716.LUT_SIZE = 5;
	defparam lut_716.mask = 32'h5f5f7fff;

	lut_sub lut_721 ({sk[185], i_4_, n_n795, n_n822, x1517x, x1519x, x452x}, x1511x);
	defparam lut_721.LUT_SIZE = 7;
	defparam lut_721.mask = 128'h333333333333333300000f0f00003f7f;

	lut_sub lut_725 ({sk[186], i_5_, i_1_, n_n792, n_n853, x9x, x17x}, x1512x);
	defparam lut_725.LUT_SIZE = 7;
	defparam lut_725.mask = 128'h33333333333333330055000300000003;

	lut_sub lut_728 ({sk[187], x17x, x6732x, x370x, x6733x, n_n791, x6734x}, x6737x);
	defparam lut_728.LUT_SIZE = 7;
	defparam lut_728.mask = 128'h0f3f0f3f0f7f0fff111f111f111fffff;

	lut_sub lut_732 ({sk[188], x1425x, x6726x, x6727x, x6728x, x6729x, x6789x}, x6791x);
	defparam lut_732.LUT_SIZE = 7;
	defparam lut_732.mask = 128'h0f3f0f3f0f7f0fff7fffffffffffffff;

	lut_sub lut_739 ({sk[189], x1503x, x1474x, x1475x, x1504x, x6745x, x6757x}, x6760x);
	defparam lut_739.LUT_SIZE = 7;
	defparam lut_739.mask = 128'h0f3f0f3f0f7f0fff7fffffffffffffff;

	lut_sub lut_746 ({sk[190], n_n849, n_n846, n_n851, x6773x, x610x, x609x}, n_n1265);
	defparam lut_746.LUT_SIZE = 7;
	defparam lut_746.mask = 128'h0f3f0f3f0f7f0fff0f0f0f0f0f5f3f7f;

	lut_sub lut_750 ({sk[191], x1438x, x1439x, x6778x, x6779x}, x6782x);
	defparam lut_750.LUT_SIZE = 5;
	defparam lut_750.mask = 32'h01337fff;

	lut_sub lut_755 ({sk[192], n_n764, x495x, x6752x, x6766x, x1466x, x6765x}, x7982x);
	defparam lut_755.LUT_SIZE = 7;
	defparam lut_755.mask = 128'h0f3f0f3f0f7f0fff8000800080000000;

	lut_sub lut_758 ({sk[193], i_1_, i_2_, i_0_, n_n541, n_n550, n_n837}, x1414x);
	defparam lut_758.LUT_SIZE = 7;
	defparam lut_758.mask = 128'h0f3f0f3f0f7f0fff0000000001000000;

	lut_sub lut_760 ({sk[194], i_0_, x265x, n_n538, n_n832, n_n550, x302x}, x1415x);
	defparam lut_760.LUT_SIZE = 7;
	defparam lut_760.mask = 128'h0f3f0f3f0f7f0fff0000050500000003;

	lut_sub lut_763 ({sk[195], i_0_, x33x, x272x, x364x, x6573x, x6795x}, x6805x);
	defparam lut_763.LUT_SIZE = 7;
	defparam lut_763.mask = 128'h0f3f0f3f0f7f0fff0055035700550055;

	lut_sub lut_766 ({sk[196], i_10_, i_11_, x1414x, x1415x, x6805x}, x6806x);
	defparam lut_766.LUT_SIZE = 6;
	defparam lut_766.mask = 64'h3333ffff5555557f;

	lut_sub lut_770 ({sk[197], i_6_, n_n541, n_n545, n_n847, x390x, x1390x}, x6820x);
	defparam lut_770.LUT_SIZE = 7;
	defparam lut_770.mask = 128'h3fff3fff3fffffff575757575555555f;

	lut_sub lut_774 ({sk[198], i_5_, i_2_, n_n665, x15x, n_n633, x287x}, x1388x);
	defparam lut_774.LUT_SIZE = 7;
	defparam lut_774.mask = 128'h3fff3fff3fffffff005500770055007f;

	lut_sub lut_778 ({sk[199], i_13_, i_11_, x30x, x15x, x123x, x7994x}, x1389x);
	defparam lut_778.LUT_SIZE = 7;
	defparam lut_778.mask = 128'h3fff3fff3fffffff00000000bbbf0000;

	lut_sub lut_782 ({sk[200], i_9_, i_10_, x6820x, x1388x, x1389x}, x1385x);
	defparam lut_782.LUT_SIZE = 6;
	defparam lut_782.mask = 64'h7f7f7f7f0000007f;

	lut_sub lut_786 ({sk[201], i_4_, i_1_, i_2_}, n_n779);
	defparam lut_786.LUT_SIZE = 4;
	defparam lut_786.mask = 16'h7708;

	lut_sub lut_788 ({sk[202], i_10_, i_13_, i_12_}, n_n849);
	defparam lut_788.LUT_SIZE = 4;
	defparam lut_788.mask = 16'h7740;

	lut_sub lut_790 ({sk[203], i_13_, i_12_, i_11_}, n_n716);
	defparam lut_790.LUT_SIZE = 4;
	defparam lut_790.mask = 16'h7720;

	lut_sub lut_792 ({sk[204], i_10_, i_7_, i_8_, i_3_, i_1_, i_2_}, x441x);
	defparam lut_792.LUT_SIZE = 7;
	defparam lut_792.mask = 128'h3fff3fff3fffffffc888000088880000;

	lut_sub lut_795 ({sk[205], i_6_, n_n779, n_n849, n_n716, n_n36, x441x}, x6833x);
	defparam lut_795.LUT_SIZE = 7;
	defparam lut_795.mask = 128'h3fff3fff3fffffff0000003305050537;

	lut_sub lut_798 ({sk[206], i_9_, i_7_, i_8_}, n_n764);
	defparam lut_798.LUT_SIZE = 4;
	defparam lut_798.mask = 16'h7710;

	lut_sub lut_800 ({sk[207], i_3_, i_1_, i_2_}, n_n675);
	defparam lut_800.LUT_SIZE = 4;
	defparam lut_800.mask = 16'h7780;

	lut_sub lut_802 ({sk[208], i_10_, i_7_, i_8_}, n_n792);
	defparam lut_802.LUT_SIZE = 4;
	defparam lut_802.mask = 16'h7780;

	lut_sub lut_804 ({sk[209], i_13_, i_4_, i_12_, i_11_}, x17x);
	defparam lut_804.LUT_SIZE = 5;
	defparam lut_804.mask = 32'h00ff0100;

	lut_sub lut_806 ({sk[210], i_9_, i_8_, i_4_, n_n853, x265x, x1381x}, x1378x);
	defparam lut_806.LUT_SIZE = 7;
	defparam lut_806.mask = 128'h3fff3fff3fffffff0505050705050505;

	lut_sub lut_809 ({sk[211], i_1_, n_n764, n_n675, n_n792, x17x, x1378x}, x6834x);
	defparam lut_809.LUT_SIZE = 7;
	defparam lut_809.mask = 128'h3fff3fff3fffffff5777777755775577;

	lut_sub lut_814 ({sk[212], i_9_, i_7_}, x267x);
	defparam lut_814.LUT_SIZE = 3;
	defparam lut_814.mask = 8'h34;

	lut_sub lut_816 ({sk[213], i_3_, i_13_, i_4_, i_12_, i_1_, i_11_}, x445x);
	defparam lut_816.LUT_SIZE = 7;
	defparam lut_816.mask = 128'h3fff3fff3fffffff4044000000440000;

	lut_sub lut_819 ({sk[214], i_8_, i_6_, x267x, n_n675, n_n545, x445x}, x1366x);
	defparam lut_819.LUT_SIZE = 7;
	defparam lut_819.mask = 128'h3fff3fff3fffffff0000000003570000;

	lut_sub lut_822 ({sk[215], i_3_, i_1_}, x328x);
	defparam lut_822.LUT_SIZE = 3;
	defparam lut_822.mask = 8'h34;

	lut_sub lut_824 ({sk[216], i_9_, i_7_, i_8_}, n_n275);
	defparam lut_824.LUT_SIZE = 4;
	defparam lut_824.mask = 16'h7720;

	lut_sub lut_826 ({sk[217], i_13_, i_11_}, n_n274);
	defparam lut_826.LUT_SIZE = 3;
	defparam lut_826.mask = 8'h38;

	lut_sub lut_828 ({sk[218], i_9_, i_7_, i_13_, i_12_, i_1_, i_11_}, x447x);
	defparam lut_828.LUT_SIZE = 7;
	defparam lut_828.mask = 128'h3fff3fff3fffffff2200200000000000;

	lut_sub lut_831 ({sk[219], i_6_, i_2_, x328x, n_n275, n_n274, x447x}, x1353x);
	defparam lut_831.LUT_SIZE = 7;
	defparam lut_831.mask = 128'h3fff3fff3fffffff0000000055570003;

	lut_sub lut_834 ({sk[220], i_9_, i_7_, i_6_, i_13_, i_12_, i_2_}, x387x);
	defparam lut_834.LUT_SIZE = 7;
	defparam lut_834.mask = 128'h3fff3fff3fffffff0000008000000000;

	lut_sub lut_836 ({sk[221], i_6_, i_13_, i_11_, x448x}, x1350x);
	defparam lut_836.LUT_SIZE = 5;
	defparam lut_836.mask = 32'h00ff1000;

	lut_sub lut_838 ({sk[222], i_11_, n_n769, n_n570, n_n819, n_n273, x328x}, x6849x);
	defparam lut_838.LUT_SIZE = 7;
	defparam lut_838.mask = 128'h3fff3fff3fffffff0005003700000033;

	lut_sub lut_841 ({sk[223], i_9_, i_8_, i_6_}, n_n769);
	defparam lut_841.LUT_SIZE = 4;
	defparam lut_841.mask = 16'h7710;

	lut_sub lut_843 ({sk[224], i_9_, i_7_, i_8_, i_6_, i_3_, i_2_}, x45x);
	defparam lut_843.LUT_SIZE = 7;
	defparam lut_843.mask = 128'h3fff3fff3fffffff000a0c0e00000000;

	lut_sub lut_846 ({sk[225], i_6_, x29x, x19x, x282x, x294x, x273x}, x1318x);
	defparam lut_846.LUT_SIZE = 7;
	defparam lut_846.mask = 128'h3fff3fff3fffffff555f777f00000000;

	lut_sub lut_850 ({sk[226], i_10_, i_8_, i_6_, i_3_, x301x, x6866x}, x6867x);
	defparam lut_850.LUT_SIZE = 7;
	defparam lut_850.mask = 128'h3fff3fff3fffffff5555755555555555;

	lut_sub lut_853 ({sk[227], i_13_, i_1_, x407x, x6855x}, x6857x);
	defparam lut_853.LUT_SIZE = 5;
	defparam lut_853.mask = 32'h00ff5755;

	lut_sub lut_856 ({sk[228], x370x, n_n672, x303x, x470x, x6853x, x6854x}, x6858x);
	defparam lut_856.LUT_SIZE = 7;
	defparam lut_856.mask = 128'h3fff3fff3fffffff003355770f3f5f7f;

	lut_sub lut_860 ({sk[229], n_n764, n_n716, n_n570, x328x, x371x, x474x}, x472x);
	defparam lut_860.LUT_SIZE = 7;
	defparam lut_860.mask = 128'h3fff3fff3fffffff00005555333f777f;

	lut_sub lut_864 ({sk[230], n_n716, n_n273, x45x, x371x, x412x, x471x}, x6860x);
	defparam lut_864.LUT_SIZE = 7;
	defparam lut_864.mask = 128'h3fff3fff3fffffff000f555f333f777f;

	lut_sub lut_868 ({sk[231], i_6_, i_1_, n_n665, n_n1574, x6873x, x6872x}, n_n1126);
	defparam lut_868.LUT_SIZE = 7;
	defparam lut_868.mask = 128'h3fff3fff3fffffff7f7f7f7f7fff7f7f;

	lut_sub lut_873 ({sk[232], i_4_, i_1_, i_11_, x490x}, x1294x);
	defparam lut_873.LUT_SIZE = 5;
	defparam lut_873.mask = 32'h00ff0100;

	lut_sub lut_875 ({sk[233], i_9_, i_6_, i_1_, x27x, x297x, x6881x}, x6882x);
	defparam lut_875.LUT_SIZE = 7;
	defparam lut_875.mask = 128'h3fff3fff3fffffff5555575555555757;

	lut_sub lut_879 ({sk[234], i_7_, n_n748, x15x, n_n432, n_n197, x1288x}, x1283x);
	defparam lut_879.LUT_SIZE = 7;
	defparam lut_879.mask = 128'h3fff3fff3fffffff00550077005f007f;

	lut_sub lut_883 ({sk[235], i_3_, n_n183, x1287x, x393x, x6888x, x7976x}, x6890x);
	defparam lut_883.LUT_SIZE = 7;
	defparam lut_883.mask = 128'h3fff3fff3fffffffbbbbbbbbbbffbfff;

	lut_sub lut_888 ({sk[236], i_3_, i_4_, i_1_, x604x, x1204x, x7975x}, x6935x);
	defparam lut_888.LUT_SIZE = 7;
	defparam lut_888.mask = 128'h3fff3fff3fffffff33333333bbbf3333;

	lut_sub lut_892 ({sk[237], n_n792, n_n273, x328x, x371x, n_n274, x49x}, x526x);
	defparam lut_892.LUT_SIZE = 7;
	defparam lut_892.mask = 128'h3fff3fff3fffffff000055550f3f5f7f;

	lut_sub lut_896 ({sk[238], n_n2368, n_n773, n_n273, x43x, x371x, n_n274}, x6941x);
	defparam lut_896.LUT_SIZE = 7;
	defparam lut_896.mask = 128'h3fff3fff3fffffff03030357ffffffff;

	lut_sub lut_900 ({sk[239], i_13_, i_1_, i_2_, x636x, x1193x, x7974x}, x634x);
	defparam lut_900.LUT_SIZE = 7;
	defparam lut_900.mask = 128'h3fff3fff3fffffffbbbbbfbbbbbbbbbb;

	lut_sub lut_904 ({sk[240], i_9_, i_10_, i_13_, i_4_, i_1_, x1185x}, x6946x);
	defparam lut_904.LUT_SIZE = 7;
	defparam lut_904.mask = 128'h3fff3fff3fffffff5755555555555555;

	lut_sub lut_907 ({sk[241], i_7_, i_2_}, x29x);
	defparam lut_907.LUT_SIZE = 3;
	defparam lut_907.mask = 8'h32;

	lut_sub lut_909 ({sk[242], i_9_, i_10_, i_7_, i_8_, i_12_, i_11_}, x595x);
	defparam lut_909.LUT_SIZE = 7;
	defparam lut_909.mask = 128'h3fff3fff3fffffff0000510000515151;

	lut_sub lut_915 ({sk[243], i_8_, i_4_, i_12_, i_11_}, x6952x);
	defparam lut_915.LUT_SIZE = 5;
	defparam lut_915.mask = 32'h00ff4000;

	lut_sub lut_917 ({sk[244], i_9_, i_10_, i_7_, i_3_, i_4_, i_2_}, x1178x);
	defparam lut_917.LUT_SIZE = 7;
	defparam lut_917.mask = 128'h3fff3fff3fffffff0000040000000404;

	lut_sub lut_920 ({sk[245], x25x, x29x, x14x, x595x, x6952x, x1178x}, n_n1189);
	defparam lut_920.LUT_SIZE = 7;
	defparam lut_920.mask = 128'h3fff3fff3fffffff555f777f777f777f;

	lut_sub lut_925 ({sk[246], i_10_, i_7_, i_11_}, n_n656);
	defparam lut_925.LUT_SIZE = 4;
	defparam lut_925.mask = 16'h7708;

	lut_sub lut_927 ({sk[247], i_7_, i_2_}, x275x);
	defparam lut_927.LUT_SIZE = 3;
	defparam lut_927.mask = 8'h38;

	lut_sub lut_929 ({sk[248], i_9_, i_7_, i_12_, i_11_, i_2_}, x6960x);
	defparam lut_929.LUT_SIZE = 6;
	defparam lut_929.mask = 64'h7f7f7f7f80a080f0;

	lut_sub lut_933 ({sk[249], i_3_, i_4_, i_11_, n_n656, x275x, x6960x}, x1169x);
	defparam lut_933.LUT_SIZE = 7;
	defparam lut_933.mask = 128'h3fff3fff3fffffff000000007f5f0000;

	lut_sub lut_937 ({sk[250], i_13_, i_12_, i_11_}, n_n853);
	defparam lut_937.LUT_SIZE = 4;
	defparam lut_937.mask = 16'h7710;

	lut_sub lut_939 ({sk[251], i_8_, i_13_, x25x, n_n822, n_n412, x330x}, x6961x);
	defparam lut_939.LUT_SIZE = 7;
	defparam lut_939.mask = 128'h3fff3fff3fffffff0537003300330033;

	lut_sub lut_942 ({sk[252], i_3_, i_4_, i_2_, n_n853, x318x, x6961x}, x6962x);
	defparam lut_942.LUT_SIZE = 7;
	defparam lut_942.mask = 128'h3fff3fff3fffffff57555f5557555755;

	lut_sub lut_946 ({sk[253], i_9_, i_10_, i_13_, i_4_}, x340x);
	defparam lut_946.LUT_SIZE = 5;
	defparam lut_946.mask = 32'h00ff4000;

	lut_sub lut_948 ({sk[254], i_10_, i_7_, i_3_, i_13_, i_4_, i_11_}, x1154x);
	defparam lut_948.LUT_SIZE = 7;
	defparam lut_948.mask = 128'h3fff3fff3fffffff1000000000000000;

	lut_sub lut_950 ({sk[255], i_3_, i_13_, i_4_, n_n792, x105x, x625x}, x6966x);
	defparam lut_950.LUT_SIZE = 7;
	defparam lut_950.mask = 128'h3fff3fff3fffffff777f5555333f0000;

	lut_sub lut_954 ({sk[256], i_9_, i_10_, i_8_, i_3_, i_13_, i_11_}, x1165x);
	defparam lut_954.LUT_SIZE = 7;
	defparam lut_954.mask = 128'h3fff3fff3fffffff8000000000000000;

	lut_sub lut_956 ({sk[257], i_9_, i_10_, i_3_, i_13_, i_12_, i_11_}, x1166x);
	defparam lut_956.LUT_SIZE = 7;
	defparam lut_956.mask = 128'h3fff3fff3fffffff8000000000000000;

	lut_sub lut_958 ({sk[258], i_10_, i_13_, i_11_}, n_n816);
	defparam lut_958.LUT_SIZE = 4;
	defparam lut_958.mask = 16'h7740;

	lut_sub lut_960 ({sk[259], i_7_, i_8_}, x27x);
	defparam lut_960.LUT_SIZE = 3;
	defparam lut_960.mask = 8'h38;

	lut_sub lut_962 ({sk[260], i_3_, i_4_, n_n849, n_n842, x352x, x351x}, x6969x);
	defparam lut_962.LUT_SIZE = 7;
	defparam lut_962.mask = 128'h3fff3fff3fffffff0055035700550055;

	lut_sub lut_965 ({sk[261], i_7_, i_2_, x618x, x1141x}, x6972x);
	defparam lut_965.LUT_SIZE = 5;
	defparam lut_965.mask = 32'h00ff5557;

	lut_sub lut_968 ({sk[262], i_9_, i_7_, i_8_, n_n2368, x295x, x1142x}, x6973x);
	defparam lut_968.LUT_SIZE = 7;
	defparam lut_968.mask = 128'h3fff3fff3fffffff5f5f5f7f5f5f5f5f;

	lut_sub lut_972 ({sk[263], i_3_, i_13_, i_2_, x8x, n_n638, x6986x}, x6987x);
	defparam lut_972.LUT_SIZE = 7;
	defparam lut_972.mask = 128'h3fff3fff3fffffff5555555f5577557f;

	lut_sub lut_976 ({sk[264], i_9_, i_10_, i_7_, i_12_, i_11_, i_2_}, x621x);
	defparam lut_976.LUT_SIZE = 7;
	defparam lut_976.mask = 128'h3fff3fff3fffffff000000000000ddd5;

	lut_sub lut_980 ({sk[265], i_9_, i_10_, i_7_, i_8_, i_12_, i_11_}, x620x);
	defparam lut_980.LUT_SIZE = 7;
	defparam lut_980.mask = 128'h3fff3fff3fffffff0000030000035353;

	lut_sub lut_984 ({sk[266], i_9_, i_7_, i_8_, i_12_, i_11_, i_2_}, x627x);
	defparam lut_984.LUT_SIZE = 7;
	defparam lut_984.mask = 128'h3fff3fff3fffffff00000000008800f0;

	lut_sub lut_988 ({sk[267], i_3_, x14x, x6987x, x621x, x620x, x627x}, x6992x);
	defparam lut_988.LUT_SIZE = 7;
	defparam lut_988.mask = 128'h3fff3fff3fffffff00ff33ff5fff7fff;

	lut_sub lut_993 ({sk[268], i_9_, i_10_, i_7_}, x314x);
	defparam lut_993.LUT_SIZE = 4;
	defparam lut_993.mask = 16'h7701;

	lut_sub lut_995 ({sk[269], i_3_, i_12_, i_2_, n_n637, n_n609, n_n597}, x1132x);
	defparam lut_995.LUT_SIZE = 7;
	defparam lut_995.mask = 128'h3fff3fff3fffffff0f0000007f000000;

	lut_sub lut_999 ({sk[270], i_8_, i_3_, i_13_, x386x, n_n656, x6980x}, x6981x);
	defparam lut_999.LUT_SIZE = 7;
	defparam lut_999.mask = 128'h3fff3fff3fffffff555f777f555f555f;

	lut_sub lut_1003 ({sk[271], i_3_, i_12_}, x365x);
	defparam lut_1003.LUT_SIZE = 3;
	defparam lut_1003.mask = 8'h32;

	lut_sub lut_1005 ({sk[272], i_8_, i_4_, i_12_, i_11_, n_n656, x275x}, x1107x);
	defparam lut_1005.LUT_SIZE = 7;
	defparam lut_1005.mask = 128'h3fff3fff3fffffff0000000000730000;

	lut_sub lut_1008 ({sk[273], i_13_, i_12_, i_11_, i_2_}, x301x);
	defparam lut_1008.LUT_SIZE = 5;
	defparam lut_1008.mask = 32'h00ff2000;

	lut_sub lut_1010 ({sk[274], i_3_, i_4_, i_2_, n_n761, x335x, x319x}, x630x);
	defparam lut_1010.LUT_SIZE = 7;
	defparam lut_1010.mask = 128'h0fff5fffffffffff00770f7700550055;

	lut_sub lut_1014 ({sk[275], i_9_, i_8_, i_13_, i_11_, n_n672, x330x}, x6996x);
	defparam lut_1014.LUT_SIZE = 7;
	defparam lut_1014.mask = 128'h0fff5fffffffffff0300070003000300;

	lut_sub lut_1017 ({sk[276], i_3_, i_13_, i_12_, i_2_, n_n764, x1095x}, x6997x);
	defparam lut_1017.LUT_SIZE = 7;
	defparam lut_1017.mask = 128'h0fff5fffffffffff5755555555555555;

	lut_sub lut_1020 ({sk[277], i_5_, i_6_, i_3_}, n_n658);
	defparam lut_1020.LUT_SIZE = 4;
	defparam lut_1020.mask = 16'h5f02;

	lut_sub lut_1022 ({sk[278], i_9_, i_10_, i_11_}, n_n741);
	defparam lut_1022.LUT_SIZE = 4;
	defparam lut_1022.mask = 16'h5f80;

	lut_sub lut_1024 ({sk[279], i_12_, i_11_}, n_n526);
	defparam lut_1024.LUT_SIZE = 3;
	defparam lut_1024.mask = 8'h58;

	lut_sub lut_1026 ({sk[280], i_1_, i_2_, i_0_}, n_n835);
	defparam lut_1026.LUT_SIZE = 4;
	defparam lut_1026.mask = 16'h5f80;

	lut_sub lut_1028 ({sk[281], i_4_, i_1_, i_0_}, n_n791);
	defparam lut_1028.LUT_SIZE = 4;
	defparam lut_1028.mask = 16'h5f08;

	lut_sub lut_1030 ({sk[282], i_9_, i_5_, i_3_, i_4_, i_1_, i_2_}, x109x);
	defparam lut_1030.LUT_SIZE = 7;
	defparam lut_1030.mask = 128'h0fff5fffffffffff0000080000000000;

	lut_sub lut_1032 ({sk[283], i_10_, i_5_, i_3_, i_1_, i_2_}, x274x);
	defparam lut_1032.LUT_SIZE = 6;
	defparam lut_1032.mask = 64'h3333333380000000;

	lut_sub lut_1034 ({sk[284], i_5_, i_1_}, x323x);
	defparam lut_1034.LUT_SIZE = 3;
	defparam lut_1034.mask = 8'h58;

	lut_sub lut_1036 ({sk[285], i_6_, i_1_}, x325x);
	defparam lut_1036.LUT_SIZE = 3;
	defparam lut_1036.mask = 8'h52;

	lut_sub lut_1038 ({sk[286], i_6_, i_1_}, x326x);
	defparam lut_1038.LUT_SIZE = 3;
	defparam lut_1038.mask = 8'h58;

	lut_sub lut_1040 ({sk[287], i_10_, i_7_, i_8_, i_5_, i_4_, i_1_}, x378x);
	defparam lut_1040.LUT_SIZE = 7;
	defparam lut_1040.mask = 128'h0fff5fffffffffff2000000000000000;

	lut_sub lut_1042 ({sk[288], i_10_, i_5_, i_6_, i_12_, i_1_, i_11_}, x979x);
	defparam lut_1042.LUT_SIZE = 7;
	defparam lut_1042.mask = 128'h0fff5fffffffffff808080c0000080c0;

	lut_sub lut_1046 ({sk[289], i_9_, i_10_, i_6_, i_12_, i_11_, i_0_}, x529x);
	defparam lut_1046.LUT_SIZE = 7;
	defparam lut_1046.mask = 128'h0fff5fffffffffff4450000000000000;

	lut_sub lut_1049 ({sk[290], i_10_, i_1_, i_0_, n_n570, x305x, x350x}, x7081x);
	defparam lut_1049.LUT_SIZE = 7;
	defparam lut_1049.mask = 128'h0fff5fffffffffff0037000500330000;

	lut_sub lut_1052 ({sk[291], i_13_, i_1_, x529x, x7081x}, x7082x);
	defparam lut_1052.LUT_SIZE = 5;
	defparam lut_1052.mask = 32'h5fff7555;

	lut_sub lut_1055 ({sk[292], i_10_, i_13_}, n_n842);
	defparam lut_1055.LUT_SIZE = 3;
	defparam lut_1055.mask = 8'h58;

	lut_sub lut_1057 ({sk[293], i_5_, i_6_, i_3_, i_2_, i_0_}, x413x);
	defparam lut_1057.LUT_SIZE = 6;
	defparam lut_1057.mask = 64'h3333333340000000;

	lut_sub lut_1059 ({sk[294], i_7_, i_8_, i_5_, i_6_, i_3_, i_2_}, x535x);
	defparam lut_1059.LUT_SIZE = 7;
	defparam lut_1059.mask = 128'h0fff5fffffffffffe000c000a0000000;

	lut_sub lut_1062 ({sk[295], i_7_, i_8_, i_5_, i_6_, i_0_}, x955x);
	defparam lut_1062.LUT_SIZE = 6;
	defparam lut_1062.mask = 64'h3333333340000000;

	lut_sub lut_1064 ({sk[296], i_4_, i_0_, n_n842, x413x, x535x, x955x}, x947x);
	defparam lut_1064.LUT_SIZE = 7;
	defparam lut_1064.mask = 128'h0fff5fffffffffff00000000005f007f;

	lut_sub lut_1068 ({sk[297], i_9_, i_10_, i_13_, i_12_, i_11_}, x303x);
	defparam lut_1068.LUT_SIZE = 6;
	defparam lut_1068.mask = 64'h3333333320000000;

	lut_sub lut_1070 ({sk[298], i_7_, i_8_, i_5_, i_3_, i_2_, x303x}, x937x);
	defparam lut_1070.LUT_SIZE = 7;
	defparam lut_1070.mask = 128'h3f3f3f3f3f3f3f3f0054004400500000;

	lut_sub lut_1073 ({sk[299], i_7_, i_13_, i_2_, n_n741, x407x, x105x}, x939x);
	defparam lut_1073.LUT_SIZE = 7;
	defparam lut_1073.mask = 128'h3f3f3f3f3f3f3f3f7f77000077770000;

	lut_sub lut_1077 ({sk[300], i_3_, i_13_, i_2_, x305x, x392x, x340x}, x7093x);
	defparam lut_1077.LUT_SIZE = 7;
	defparam lut_1077.mask = 128'h3f3f3f3f3f3f3f3f7f7f5f5f7f775f55;

	lut_sub lut_1082 ({sk[301], i_0_, x937x, x939x, x7093x}, n_n972);
	defparam lut_1082.LUT_SIZE = 5;
	defparam lut_1082.mask = 32'h3fff0f7f;

	lut_sub lut_1086 ({sk[302], i_1_, i_2_, i_0_}, n_n838);
	defparam lut_1086.LUT_SIZE = 4;
	defparam lut_1086.mask = 16'h7740;

	lut_sub lut_1088 ({sk[303], i_5_, i_0_, x24x, x387x, n_n752}, x928x);
	defparam lut_1088.LUT_SIZE = 6;
	defparam lut_1088.mask = 64'h55ff55ff00000037;

	lut_sub lut_1091 ({sk[304], i_9_, i_7_, i_5_, n_n838, n_n274, x928x}, x7101x);
	defparam lut_1091.LUT_SIZE = 7;
	defparam lut_1091.mask = 128'h3f3f3f3f3f3f3f3f5557555555555555;

	lut_sub lut_1094 ({sk[305], i_9_, i_13_, i_12_, i_11_}, x335x);
	defparam lut_1094.LUT_SIZE = 5;
	defparam lut_1094.mask = 32'h3fff8000;

	lut_sub lut_1096 ({sk[306], i_9_, i_7_, i_8_, i_13_, i_4_, i_11_}, x7099x);
	defparam lut_1096.LUT_SIZE = 7;
	defparam lut_1096.mask = 128'h3f3f3f3f3f3f3f3fa0b0003000000000;

	lut_sub lut_1099 ({sk[307], i_8_, x12x, x24x, n_n719, n_n670, n_n550}, x7967x);
	defparam lut_1099.LUT_SIZE = 7;
	defparam lut_1099.mask = 128'h3f3f3f3f3f3f3f3ffffffcccffffeecc;

	lut_sub lut_1112 ({sk[308], i_2_, i_0_, x12x, x335x, x7099x, x7967x}, x7102x);
	defparam lut_1112.LUT_SIZE = 7;
	defparam lut_1112.mask = 128'h3f3f3f3f3f3f3f3faaaaaabfaaaaaaaa;

	lut_sub lut_1116 ({sk[309], n_n624, n_n277, x401x, x76x, x403x, x912x}, x670x);
	defparam lut_1116.LUT_SIZE = 7;
	defparam lut_1116.mask = 128'h3f3f3f3f3f3f3f3f7fff7fff7fffffff;

	lut_sub lut_1122 ({sk[310], i_8_, i_13_, i_12_, i_11_, x274x, x908x}, x7113x);
	defparam lut_1122.LUT_SIZE = 7;
	defparam lut_1122.mask = 128'h0f0fffffffffffff5555555557555555;

	lut_sub lut_1125 ({sk[311], i_7_, i_5_, i_2_, x19x, x282x, x273x}, x895x);
	defparam lut_1125.LUT_SIZE = 7;
	defparam lut_1125.mask = 128'h0f0fffffffffffff5757000077570000;

	lut_sub lut_1129 ({sk[312], i_13_, i_11_, i_2_, x35x, n_n773, x894x}, x7115x);
	defparam lut_1129.LUT_SIZE = 7;
	defparam lut_1129.mask = 128'h0f0fffffffffffff5555575555555555;

	lut_sub lut_1132 ({sk[313], i_13_, i_12_, x670x, x7113x, x895x, x7115x}, x7118x);
	defparam lut_1132.LUT_SIZE = 7;
	defparam lut_1132.mask = 128'h0f0fffffffffffff7f7f7fff7f7f7f7f;

	lut_sub lut_1137 ({sk[314], i_9_, i_8_, i_5_, i_4_, i_1_, i_2_}, x406x);
	defparam lut_1137.LUT_SIZE = 7;
	defparam lut_1137.mask = 128'h0f0fffffffffffff0000000800000000;

	lut_sub lut_1139 ({sk[315], i_9_, i_7_, i_5_, i_1_, i_11_, i_2_}, x71x);
	defparam lut_1139.LUT_SIZE = 7;
	defparam lut_1139.mask = 128'h0f0fffffffffffff0080000000000000;

	lut_sub lut_1141 ({sk[316], i_9_, i_7_, i_8_, i_3_, i_4_, i_2_}, x715x);
	defparam lut_1141.LUT_SIZE = 7;
	defparam lut_1141.mask = 128'h0f0fffffffffffff2020203300000000;

	lut_sub lut_1144 ({sk[317], x12x, n_n761, x406x, x71x, x109x, x715x}, x884x);
	defparam lut_1144.LUT_SIZE = 7;
	defparam lut_1144.mask = 128'h0f0fffffffffffff00003fff00007fff;

	lut_sub lut_1149 ({sk[318], i_9_, i_13_, i_11_}, n_n755);
	defparam lut_1149.LUT_SIZE = 4;
	defparam lut_1149.mask = 16'h0f40;

	lut_sub lut_1151 ({sk[319], i_9_, i_7_, i_5_, n_n570, x877x, x7966x}, x639x);
	defparam lut_1151.LUT_SIZE = 7;
	defparam lut_1151.mask = 128'h0f0fffffffffffff33bb33bf33bb33bb;

	lut_sub lut_1155 ({sk[320], i_7_, i_5_, i_4_, n_n683, x7147x, x7145x}, x721x);
	defparam lut_1155.LUT_SIZE = 7;
	defparam lut_1155.mask = 128'h0f0fffffffffffff33773333337f3333;

	lut_sub lut_1159 ({sk[321], i_3_, n_n185, n_n683, n_n752, x284x, x280x}, x868x);
	defparam lut_1159.LUT_SIZE = 7;
	defparam lut_1159.mask = 128'h0f0fffffffffffff0101013300000033;

	lut_sub lut_1162 ({sk[322], i_7_, n_n545, x377x, n_n678, x26x, n_n755}, x869x);
	defparam lut_1162.LUT_SIZE = 7;
	defparam lut_1162.mask = 128'h0f0fffffffffffff0000003301010133;

	lut_sub lut_1165 ({sk[323], n_n838, n_n755, x639x, x721x, x868x, x869x}, x7151x);
	defparam lut_1165.LUT_SIZE = 7;
	defparam lut_1165.mask = 128'h0f0fffffffffffff77777f7f77ff7fff;

	lut_sub lut_1170 ({sk[324], i_7_, i_8_, i_3_, n_n773, n_n835, n_n671}, x725x);
	defparam lut_1170.LUT_SIZE = 7;
	defparam lut_1170.mask = 128'h0f0fffffffffffff3737373737050505;

	lut_sub lut_1174 ({sk[325], i_5_, i_3_, i_0_, x37x, n_n725, n_n843}, x811x);
	defparam lut_1174.LUT_SIZE = 7;
	defparam lut_1174.mask = 128'h0f0fffffffffffff0000000015000500;

	lut_sub lut_1177 ({sk[326], i_8_, n_n849, x37x, n_n771, x13x, n_n671}, x813x);
	defparam lut_1177.LUT_SIZE = 7;
	defparam lut_1177.mask = 128'h0f0fffffffffffff0011031300110011;

	lut_sub lut_1180 ({sk[327], i_13_, i_12_, i_11_, n_n835, n_n712, x398x}, x7166x);
	defparam lut_1180.LUT_SIZE = 7;
	defparam lut_1180.mask = 128'h0f0fffffffffffff0000035700000000;

	lut_sub lut_1183 ({sk[328], i_5_, n_n716, x725x, x811x, x813x, x7166x}, x7169x);
	defparam lut_1183.LUT_SIZE = 7;
	defparam lut_1183.mask = 128'h0f0fffffffffffff7f7f7f7f7f7f7fff;

	lut_sub lut_1188 ({sk[329], i_3_, i_1_, i_0_}, n_n687);
	defparam lut_1188.LUT_SIZE = 4;
	defparam lut_1188.mask = 16'h0f40;

	lut_sub lut_1190 ({sk[330], i_9_, i_8_, i_13_, i_4_, i_12_, i_11_}, x735x);
	defparam lut_1190.LUT_SIZE = 7;
	defparam lut_1190.mask = 128'h0f0fffffffffffffaf00cf0000000000;

	lut_sub lut_1194 ({sk[331], i_7_, i_8_, i_1_, x24x, x335x, x803x}, x732x);
	defparam lut_1194.LUT_SIZE = 7;
	defparam lut_1194.mask = 128'h0f0fffffffffffff7755775577557f55;

	lut_sub lut_1198 ({sk[332], i_1_, i_0_, x24x, x13x, n_n719, x7172x}, x7176x);
	defparam lut_1198.LUT_SIZE = 7;
	defparam lut_1198.mask = 128'h0f0fffffffffffff0055035700550055;

	lut_sub lut_1201 ({sk[333], x20x, n_n687, x34x, x735x, x732x, x7176x}, n_n977);
	defparam lut_1201.LUT_SIZE = 7;
	defparam lut_1201.mask = 128'h0f0fffffffffffff5555555f7777777f;

	lut_sub lut_1205 ({sk[334], i_4_, n_n752, x778x, x7187x, x656x, x7185x}, n_n991);
	defparam lut_1205.LUT_SIZE = 7;
	defparam lut_1205.mask = 128'h0f0fffffffffffff5fff7fff0f0f0f0f;

	lut_sub lut_1210 ({sk[335], x373x, x7192x, x256x, x7196x}, x7198x);
	defparam lut_1210.LUT_SIZE = 5;
	defparam lut_1210.mask = 32'h0fff7fff;

	lut_sub lut_1215 ({sk[336], x7213x, x214x, x7211x, x7212x, x7230x}, x7232x);
	defparam lut_1215.LUT_SIZE = 6;
	defparam lut_1215.mask = 64'h5577ffff7fffffff;

	lut_sub lut_1221 ({sk[337], i_4_, i_1_, x227x, x7222x, x739x}, x7233x);
	defparam lut_1221.LUT_SIZE = 6;
	defparam lut_1221.mask = 64'h5577ffff3f7f3f3f;

	lut_sub lut_1225 ({sk[338], x199x, x201x, x7240x}, x7242x);
	defparam lut_1225.LUT_SIZE = 4;
	defparam lut_1225.mask = 16'h0f7f;

	lut_sub lut_1229 ({sk[339], x785x, x7205x, x784x, x7204x, x7968x}, x7243x);
	defparam lut_1229.LUT_SIZE = 6;
	defparam lut_1229.mask = 64'h5577ffffbfffffff;

	lut_sub lut_1235 ({sk[340], i_2_, n_n432, x168x, x36x, x162x, x7260x}, x7262x);
	defparam lut_1235.LUT_SIZE = 7;
	defparam lut_1235.mask = 128'h0f0fffffffffffff7777777777ff7fff;

	lut_sub lut_1240 ({sk[341], i_10_, x557x, x192x, x177x, x7256x, x7252x}, x7263x);
	defparam lut_1240.LUT_SIZE = 7;
	defparam lut_1240.mask = 128'h0f0fffffffffffff7fff7fff7fffffff;

	lut_sub lut_1246 ({sk[342], i_8_, x596x, x7289x, x7290x, x7291x, x7308x}, x7310x);
	defparam lut_1246.LUT_SIZE = 7;
	defparam lut_1246.mask = 128'h0f0fffffffffffff7fffffff7fff7fff;

	lut_sub lut_1252 ({sk[343], i_8_, n_n213, x705x, x7300x, x750x, x7307x}, x7311x);
	defparam lut_1252.LUT_SIZE = 7;
	defparam lut_1252.mask = 128'h0f0fffffffffffff7f7f7fff5f5f5fff;

	lut_sub lut_1257 ({sk[344], i_5_, x25x, n_n844, x314x, x752x, x7316x}, x7318x);
	defparam lut_1257.LUT_SIZE = 7;
	defparam lut_1257.mask = 128'h0f0fffffffffffff555f777f55557777;

	lut_sub lut_1261 ({sk[345], x7272x, x7278x, x7279x, x7270x, x7271x}, x7319x);
	defparam lut_1261.LUT_SIZE = 6;
	defparam lut_1261.mask = 64'h5577ffff7fffffff;

	lut_sub lut_1267 ({sk[346], i_10_, i_7_, i_6_}, n_n699);
	defparam lut_1267.LUT_SIZE = 4;
	defparam lut_1267.mask = 16'h0f80;

	lut_sub lut_1269 ({sk[347], i_10_, i_13_, i_12_}, n_n575);
	defparam lut_1269.LUT_SIZE = 4;
	defparam lut_1269.mask = 16'h0f80;

	lut_sub lut_1271 ({sk[348], i_3_, i_13_, i_12_, i_11_, i_2_}, x759x);
	defparam lut_1271.LUT_SIZE = 6;
	defparam lut_1271.mask = 64'h5577ffffc8008800;

	lut_sub lut_1274 ({sk[349], i_10_, i_13_, i_4_, i_1_, n_n526, x27x}, x7965x);
	defparam lut_1274.LUT_SIZE = 7;
	defparam lut_1274.mask = 128'h0f0fffffffffffffcf8fffffffffffff;

	lut_sub lut_1280 ({sk[350], x16x, x325x, n_n699, n_n575, x759x, x7965x}, x52x);
	defparam lut_1280.LUT_SIZE = 7;
	defparam lut_1280.mask = 128'h0f0fffffffffffff00000000aabbafbf;

	lut_sub lut_1284 ({sk[351], i_7_, i_8_, i_5_, n_n687, n_n729, x49x}, x50x);
	defparam lut_1284.LUT_SIZE = 7;
	defparam lut_1284.mask = 128'h0f0fffffffffffff0700050000000000;

	lut_sub lut_1287 ({sk[352], i_8_, i_5_, i_4_, n_n838, n_n842, x7329x}, x7330x);
	defparam lut_1287.LUT_SIZE = 7;
	defparam lut_1287.mask = 128'h0f0fffffffffffff5557555555555555;

	lut_sub lut_1290 ({sk[353], x52x, x50x, x7330x}, n_n957);
	defparam lut_1290.LUT_SIZE = 4;
	defparam lut_1290.mask = 16'h0f7f;

	lut_sub lut_1294 ({sk[354], i_1_, i_2_}, x265x);
	defparam lut_1294.LUT_SIZE = 3;
	defparam lut_1294.mask = 8'h38;

	lut_sub lut_1296 ({sk[355], i_10_, i_13_, i_12_, i_11_}, x313x);
	defparam lut_1296.LUT_SIZE = 5;
	defparam lut_1296.mask = 32'h0fff1000;

	lut_sub lut_1298 ({sk[356], i_9_, i_4_}, x9x);
	defparam lut_1298.LUT_SIZE = 3;
	defparam lut_1298.mask = 8'h34;

	lut_sub lut_1300 ({sk[357], i_9_, i_7_, i_8_}, n_n795);
	defparam lut_1300.LUT_SIZE = 4;
	defparam lut_1300.mask = 16'h0f80;

	lut_sub lut_1302 ({sk[358], i_5_, i_4_}, x35x);
	defparam lut_1302.LUT_SIZE = 3;
	defparam lut_1302.mask = 8'h34;

	lut_sub lut_1304 ({sk[359], i_10_, i_13_, i_4_, i_12_}, x37x);
	defparam lut_1304.LUT_SIZE = 5;
	defparam lut_1304.mask = 32'h0fff1000;

	lut_sub lut_1306 ({sk[360], i_10_, i_8_, i_1_, i_2_, i_0_}, x6718x);
	defparam lut_1306.LUT_SIZE = 6;
	defparam lut_1306.mask = 64'h5577ffff80000000;

	lut_sub lut_1308 ({sk[361], i_10_, i_12_, i_11_}, n_n822);
	defparam lut_1308.LUT_SIZE = 4;
	defparam lut_1308.mask = 16'h0f10;

	lut_sub lut_1310 ({sk[362], i_9_, i_13_, i_4_}, x24x);
	defparam lut_1310.LUT_SIZE = 4;
	defparam lut_1310.mask = 16'h0f40;

	lut_sub lut_1312 ({sk[363], i_8_, i_5_}, x288x);
	defparam lut_1312.LUT_SIZE = 3;
	defparam lut_1312.mask = 8'h38;

	lut_sub lut_1314 ({sk[364], i_9_, i_8_, i_5_, i_6_}, x322x);
	defparam lut_1314.LUT_SIZE = 5;
	defparam lut_1314.mask = 32'h0fff0100;

	lut_sub lut_1316 ({sk[365], i_10_, i_8_, i_6_}, n_n773);
	defparam lut_1316.LUT_SIZE = 4;
	defparam lut_1316.mask = 16'h0f80;

	lut_sub lut_1318 ({sk[366], i_4_, i_2_, i_0_}, n_n771);
	defparam lut_1318.LUT_SIZE = 4;
	defparam lut_1318.mask = 16'h0f08;

	lut_sub lut_1320 ({sk[367], i_10_, i_8_, i_6_, i_4_, i_2_, i_0_}, x394x);
	defparam lut_1320.LUT_SIZE = 7;
	defparam lut_1320.mask = 128'h0f0fffffffffffff0800000000000000;

	lut_sub lut_1322 ({sk[368], i_1_, i_2_, i_0_}, n_n833);
	defparam lut_1322.LUT_SIZE = 4;
	defparam lut_1322.mask = 16'h0f04;

	lut_sub lut_1324 ({sk[369], i_5_, i_3_, i_4_}, n_n538);
	defparam lut_1324.LUT_SIZE = 4;
	defparam lut_1324.mask = 16'h0f02;

	lut_sub lut_1326 ({sk[370], i_7_, i_8_, i_6_}, n_n850);
	defparam lut_1326.LUT_SIZE = 4;
	defparam lut_1326.mask = 16'h0f40;

	lut_sub lut_1328 ({sk[371], i_10_, i_11_}, n_n453);
	defparam lut_1328.LUT_SIZE = 3;
	defparam lut_1328.mask = 8'h32;

	lut_sub lut_1330 ({sk[372], i_10_, i_13_, i_12_, i_11_}, n_n498);
	defparam lut_1330.LUT_SIZE = 5;
	defparam lut_1330.mask = 32'h0fff0020;

	lut_sub lut_1332 ({sk[373], i_7_, i_6_}, x269x);
	defparam lut_1332.LUT_SIZE = 3;
	defparam lut_1332.mask = 8'h34;

	lut_sub lut_1334 ({sk[374], i_7_, i_8_, i_6_}, n_n748);
	defparam lut_1334.LUT_SIZE = 4;
	defparam lut_1334.mask = 16'h0f10;

	lut_sub lut_1336 ({sk[375], i_10_, i_13_, i_12_, i_11_}, n_n725);
	defparam lut_1336.LUT_SIZE = 5;
	defparam lut_1336.mask = 32'h0fff2000;

	lut_sub lut_1338 ({sk[376], i_5_, i_3_, i_4_}, n_n541);
	defparam lut_1338.LUT_SIZE = 4;
	defparam lut_1338.mask = 16'h0f20;

	lut_sub lut_1340 ({sk[377], i_9_, i_5_, i_3_, i_4_}, x341x);
	defparam lut_1340.LUT_SIZE = 5;
	defparam lut_1340.mask = 32'h0fff0020;

	lut_sub lut_1342 ({sk[378], i_7_, i_8_, i_6_}, n_n746);
	defparam lut_1342.LUT_SIZE = 4;
	defparam lut_1342.mask = 16'h0f20;

	lut_sub lut_1344 ({sk[379], i_10_, i_13_, i_11_}, n_n729);
	defparam lut_1344.LUT_SIZE = 4;
	defparam lut_1344.mask = 16'h0f80;

	lut_sub lut_1346 ({sk[380], i_10_, i_13_, i_12_, i_11_}, x329x);
	defparam lut_1346.LUT_SIZE = 5;
	defparam lut_1346.mask = 32'h0fff8000;

	lut_sub lut_1348 ({sk[381], i_9_, i_8_, i_6_}, x6549x);
	defparam lut_1348.LUT_SIZE = 4;
	defparam lut_1348.mask = 16'h0f02;

	lut_sub lut_1350 ({sk[382], i_7_, i_8_, i_6_}, n_n756);
	defparam lut_1350.LUT_SIZE = 4;
	defparam lut_1350.mask = 16'h0f02;

	lut_sub lut_1352 ({sk[383], i_9_, i_7_, i_8_, i_6_, i_13_, i_12_}, x424x);
	defparam lut_1352.LUT_SIZE = 7;
	defparam lut_1352.mask = 128'h0f0fffffffffffff0c00080000000000;

	lut_sub lut_1355 ({sk[384], i_9_, i_8_, i_11_}, n_n623);
	defparam lut_1355.LUT_SIZE = 4;
	defparam lut_1355.mask = 16'h0f02;

	lut_sub lut_1357 ({sk[385], i_9_, i_10_, i_8_}, n_n619);
	defparam lut_1357.LUT_SIZE = 4;
	defparam lut_1357.mask = 16'h0f01;

	lut_sub lut_1359 ({sk[386], i_5_, i_1_, i_2_}, n_n612);
	defparam lut_1359.LUT_SIZE = 4;
	defparam lut_1359.mask = 16'h0f01;

	lut_sub lut_1361 ({sk[387], i_9_, i_7_, i_8_, i_5_, i_1_, i_11_}, x1755x);
	defparam lut_1361.LUT_SIZE = 7;
	defparam lut_1361.mask = 128'h0f0fffffffffffff0000000000000008;

	lut_sub lut_1363 ({sk[388], i_7_, i_5_}, x30x);
	defparam lut_1363.LUT_SIZE = 3;
	defparam lut_1363.mask = 8'h38;

	lut_sub lut_1365 ({sk[389], i_10_, i_8_, i_11_}, n_n609);
	defparam lut_1365.LUT_SIZE = 4;
	defparam lut_1365.mask = 16'h0f08;

	lut_sub lut_1367 ({sk[390], i_6_, i_0_}, x36x);
	defparam lut_1367.LUT_SIZE = 3;
	defparam lut_1367.mask = 8'h31;

	lut_sub lut_1369 ({sk[391], i_7_, i_5_, i_6_, i_1_, i_2_, i_0_}, x433x);
	defparam lut_1369.LUT_SIZE = 7;
	defparam lut_1369.mask = 128'h0f0fffffffffffffeec0aa80ccc08880;

	lut_sub lut_1375 ({sk[392], i_9_, i_10_, i_8_, i_2_}, x6559x);
	defparam lut_1375.LUT_SIZE = 5;
	defparam lut_1375.mask = 32'h0fff0001;

	lut_sub lut_1377 ({sk[393], i_5_, i_6_, i_1_, i_2_, i_0_}, x436x);
	defparam lut_1377.LUT_SIZE = 6;
	defparam lut_1377.mask = 64'h5577ffff8088c0cc;

	lut_sub lut_1382 ({sk[394], i_9_, i_10_, i_7_, i_3_, i_4_, i_1_}, x1381x);
	defparam lut_1382.LUT_SIZE = 7;
	defparam lut_1382.mask = 128'h0f0fffffffffffff2020002020000000;

	lut_sub lut_1385 ({sk[395], i_13_, i_12_}, n_n570);
	defparam lut_1385.LUT_SIZE = 3;
	defparam lut_1385.mask = 8'h38;

	lut_sub lut_1387 ({sk[396], i_3_, i_1_}, x31x);
	defparam lut_1387.LUT_SIZE = 3;
	defparam lut_1387.mask = 8'h38;

	lut_sub lut_1389 ({sk[397], i_8_, i_6_}, x289x);
	defparam lut_1389.LUT_SIZE = 3;
	defparam lut_1389.mask = 8'h34;

	lut_sub lut_1391 ({sk[398], i_9_, i_8_}, x309x);
	defparam lut_1391.LUT_SIZE = 3;
	defparam lut_1391.mask = 8'h34;

	lut_sub lut_1393 ({sk[399], i_9_, i_7_, i_6_}, n_n819);
	defparam lut_1393.LUT_SIZE = 4;
	defparam lut_1393.mask = 16'h0f10;

	lut_sub lut_1395 ({sk[400], i_3_, i_1_, i_2_}, n_n273);
	defparam lut_1395.LUT_SIZE = 4;
	defparam lut_1395.mask = 16'h0f20;

	lut_sub lut_1397 ({sk[401], i_3_, i_4_, i_1_, i_2_, x267x, x309x}, x448x);
	defparam lut_1397.LUT_SIZE = 7;
	defparam lut_1397.mask = 128'h0f0fffffffffffff0000f30000005000;

	lut_sub lut_1401 ({sk[402], i_1_, i_0_}, x377x);
	defparam lut_1401.LUT_SIZE = 3;
	defparam lut_1401.mask = 8'h38;

	lut_sub lut_1403 ({sk[403], i_1_, i_2_, i_0_}, n_n847);
	defparam lut_1403.LUT_SIZE = 4;
	defparam lut_1403.mask = 16'h0f20;

	lut_sub lut_1405 ({sk[404], i_3_, i_1_}, x15x);
	defparam lut_1405.LUT_SIZE = 3;
	defparam lut_1405.mask = 8'h31;

	lut_sub lut_1407 ({sk[405], i_3_, i_1_, i_2_}, n_n814);
	defparam lut_1407.LUT_SIZE = 4;
	defparam lut_1407.mask = 16'h0f01;

	lut_sub lut_1409 ({sk[406], i_7_, i_6_}, x28x);
	defparam lut_1409.LUT_SIZE = 3;
	defparam lut_1409.mask = 8'h38;

	lut_sub lut_1411 ({sk[407], i_10_, i_11_}, n_n213);
	defparam lut_1411.LUT_SIZE = 3;
	defparam lut_1411.mask = 8'h31;

	lut_sub lut_1413 ({sk[408], i_9_, i_10_, i_11_}, n_n421);
	defparam lut_1413.LUT_SIZE = 4;
	defparam lut_1413.mask = 16'h0f01;

	lut_sub lut_1415 ({sk[409], i_10_, i_12_, i_11_}, n_n415);
	defparam lut_1415.LUT_SIZE = 4;
	defparam lut_1415.mask = 16'h0f01;

	lut_sub lut_1417 ({sk[410], i_9_, i_7_, i_6_}, n_n358);
	defparam lut_1417.LUT_SIZE = 4;
	defparam lut_1417.mask = 16'h0f01;

	lut_sub lut_1419 ({sk[411], i_3_, i_4_, i_2_}, n_n412);
	defparam lut_1419.LUT_SIZE = 4;
	defparam lut_1419.mask = 16'h0f04;

	lut_sub lut_1421 ({sk[412], i_12_, i_11_}, n_n311);
	defparam lut_1421.LUT_SIZE = 3;
	defparam lut_1421.mask = 8'h34;

	lut_sub lut_1423 ({sk[413], i_5_, i_6_}, x13x);
	defparam lut_1423.LUT_SIZE = 3;
	defparam lut_1423.mask = 8'h32;

	lut_sub lut_1425 ({sk[414], i_5_, i_6_, i_3_}, n_n639);
	defparam lut_1425.LUT_SIZE = 4;
	defparam lut_1425.mask = 16'h0f04;

	lut_sub lut_1427 ({sk[415], i_7_, i_8_, i_5_}, n_n185);
	defparam lut_1427.LUT_SIZE = 4;
	defparam lut_1427.mask = 16'h0f02;

	lut_sub lut_1429 ({sk[416], i_3_, i_1_, i_0_}, n_n826);
	defparam lut_1429.LUT_SIZE = 4;
	defparam lut_1429.mask = 16'h0f01;

	lut_sub lut_1431 ({sk[417], i_3_, i_2_}, x96x);
	defparam lut_1431.LUT_SIZE = 3;
	defparam lut_1431.mask = 8'h3e;

	lut_sub lut_1434 ({sk[418], i_3_, i_4_, i_0_}, n_n153);
	defparam lut_1434.LUT_SIZE = 4;
	defparam lut_1434.mask = 16'h0f04;

	lut_sub lut_1436 ({sk[419], i_12_, i_11_}, n_n316);
	defparam lut_1436.LUT_SIZE = 3;
	defparam lut_1436.mask = 8'h32;

	lut_sub lut_1438 ({sk[420], i_7_, i_8_, i_6_}, n_n843);
	defparam lut_1438.LUT_SIZE = 4;
	defparam lut_1438.mask = 16'h0f80;

	lut_sub lut_1440 ({sk[421], i_3_, i_4_, i_0_}, n_n678);
	defparam lut_1440.LUT_SIZE = 4;
	defparam lut_1440.mask = 16'h0f20;

	lut_sub lut_1442 ({sk[422], i_3_, i_2_, i_0_}, n_n671);
	defparam lut_1442.LUT_SIZE = 4;
	defparam lut_1442.mask = 16'h0f80;

	lut_sub lut_1444 ({sk[423], i_5_, i_6_}, x26x);
	defparam lut_1444.LUT_SIZE = 3;
	defparam lut_1444.mask = 8'h34;

	lut_sub lut_1446 ({sk[424], i_8_, i_5_, i_6_}, n_n176);
	defparam lut_1446.LUT_SIZE = 4;
	defparam lut_1446.mask = 16'h0f04;

	lut_sub lut_1448 ({sk[425], i_5_, i_3_, i_4_}, n_n712);
	defparam lut_1448.LUT_SIZE = 4;
	defparam lut_1448.mask = 16'h0f04;

	lut_sub lut_1450 ({sk[426], i_9_, i_13_, i_11_}, n_n719);
	defparam lut_1450.LUT_SIZE = 4;
	defparam lut_1450.mask = 16'h0f80;

	lut_sub lut_1452 ({sk[427], i_9_, i_7_, i_5_}, n_n827);
	defparam lut_1452.LUT_SIZE = 4;
	defparam lut_1452.mask = 16'h0f10;

	lut_sub lut_1454 ({sk[428], i_3_, i_4_, i_1_}, n_n685);
	defparam lut_1454.LUT_SIZE = 4;
	defparam lut_1454.mask = 16'h0f20;

	lut_sub lut_1456 ({sk[429], i_3_, i_1_, i_0_}, n_n683);
	defparam lut_1456.LUT_SIZE = 4;
	defparam lut_1456.mask = 16'h0f80;

	lut_sub lut_1458 ({sk[430], i_10_, i_7_, i_8_, i_6_, i_0_}, x6732x);
	defparam lut_1458.LUT_SIZE = 6;
	defparam lut_1458.mask = 64'h5577ffff80000000;

	lut_sub lut_1460 ({sk[431], i_13_, i_4_, i_11_}, x370x);
	defparam lut_1460.LUT_SIZE = 4;
	defparam lut_1460.mask = 16'h0f10;

	lut_sub lut_1462 ({sk[432], i_10_, i_7_, i_8_, i_5_, i_6_}, x6733x);
	defparam lut_1462.LUT_SIZE = 6;
	defparam lut_1462.mask = 64'h5577ffff80000000;

	lut_sub lut_1464 ({sk[433], i_10_, i_7_, i_8_, i_13_, i_12_, i_11_}, x6734x);
	defparam lut_1464.LUT_SIZE = 7;
	defparam lut_1464.mask = 128'h0f0fffffffffffff1000000000000000;

	lut_sub lut_1466 ({sk[434], i_10_, i_6_, i_13_, i_4_, i_11_, i_0_}, x1517x);
	defparam lut_1466.LUT_SIZE = 7;
	defparam lut_1466.mask = 128'h0f0fffffffffffff0100000000000000;

	lut_sub lut_1468 ({sk[435], i_10_, i_13_, i_1_, i_11_, i_0_}, x1519x);
	defparam lut_1468.LUT_SIZE = 6;
	defparam lut_1468.mask = 64'h5577ffff01000000;

	lut_sub lut_1470 ({sk[436], i_5_, i_6_, i_13_, i_1_}, x452x);
	defparam lut_1470.LUT_SIZE = 5;
	defparam lut_1470.mask = 32'h0fff00c4;

	lut_sub lut_1473 ({sk[437], i_8_, i_5_, i_6_, i_3_}, x6628x);
	defparam lut_1473.LUT_SIZE = 5;
	defparam lut_1473.mask = 32'h0fff0020;

	lut_sub lut_1475 ({sk[438], i_8_, i_5_, i_6_, i_3_}, x6629x);
	defparam lut_1475.LUT_SIZE = 5;
	defparam lut_1475.mask = 32'h0fff0002;

	lut_sub lut_1477 ({sk[439], i_1_, i_2_, i_0_, x317x, x6628x, x6629x}, x455x);
	defparam lut_1477.LUT_SIZE = 7;
	defparam lut_1477.mask = 128'h0f0fffffffffffff000055330000000f;

	lut_sub lut_1481 ({sk[440], i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x453x);
	defparam lut_1481.LUT_SIZE = 7;
	defparam lut_1481.mask = 128'h0f0fffffffffffff0080000000400000;

	lut_sub lut_1484 ({sk[441], i_5_, i_6_, i_3_}, n_n633);
	defparam lut_1484.LUT_SIZE = 4;
	defparam lut_1484.mask = 16'h0f01;

	lut_sub lut_1486 ({sk[442], i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x456x);
	defparam lut_1486.LUT_SIZE = 7;
	defparam lut_1486.mask = 128'h0f0fffffffffffff0020000200100000;

	lut_sub lut_1490 ({sk[443], i_13_, i_11_, n_n638, n_n844, n_n633, x456x}, x1649x);
	defparam lut_1490.LUT_SIZE = 7;
	defparam lut_1490.mask = 128'h0f0fffffffffffff0000000000570003;

	lut_sub lut_1493 ({sk[444], i_7_, i_8_, i_6_}, n_n752);
	defparam lut_1493.LUT_SIZE = 4;
	defparam lut_1493.mask = 16'h0f01;

	lut_sub lut_1495 ({sk[445], i_1_, i_2_, i_0_}, n_n840);
	defparam lut_1495.LUT_SIZE = 4;
	defparam lut_1495.mask = 16'h0f02;

	lut_sub lut_1497 ({sk[446], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x409x);
	defparam lut_1497.LUT_SIZE = 7;
	defparam lut_1497.mask = 128'h0f0fffffffffffff0000000000000002;

	lut_sub lut_1499 ({sk[447], i_1_, i_2_, i_0_}, n_n852);
	defparam lut_1499.LUT_SIZE = 4;
	defparam lut_1499.mask = 16'h0f10;

	lut_sub lut_1501 ({sk[448], i_5_, i_6_}, x11x);
	defparam lut_1501.LUT_SIZE = 3;
	defparam lut_1501.mask = 8'h38;

	lut_sub lut_1503 ({sk[449], i_7_, i_6_}, x268x);
	defparam lut_1503.LUT_SIZE = 3;
	defparam lut_1503.mask = 8'h32;

	lut_sub lut_1505 ({sk[450], i_7_, i_8_, i_6_}, n_n832);
	defparam lut_1505.LUT_SIZE = 4;
	defparam lut_1505.mask = 16'h0f08;

	lut_sub lut_1507 ({sk[451], i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x462x);
	defparam lut_1507.LUT_SIZE = 7;
	defparam lut_1507.mask = 128'h0f0fffffffffffff0000001000020020;

	lut_sub lut_1511 ({sk[452], i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x461x);
	defparam lut_1511.LUT_SIZE = 7;
	defparam lut_1511.mask = 128'h0f0fffffffffffff0004004000000080;

	lut_sub lut_1515 ({sk[453], i_10_, i_7_, i_8_, i_5_, i_6_, i_3_}, x6583x);
	defparam lut_1515.LUT_SIZE = 7;
	defparam lut_1515.mask = 128'h0f0fffffffffffff0000000040000000;

	lut_sub lut_1517 ({sk[454], i_9_, i_5_, i_3_, n_n637, n_n832, n_n852}, x7979x);
	defparam lut_1517.LUT_SIZE = 7;
	defparam lut_1517.mask = 128'h0f0ffffffffffffffffffffffffffeff;

	lut_sub lut_1533 ({sk[455], i_10_, i_7_, i_8_, i_5_, i_1_, i_11_}, x1702x);
	defparam lut_1533.LUT_SIZE = 7;
	defparam lut_1533.mask = 128'h0f0fffffffffffff0000000080000000;

	lut_sub lut_1535 ({sk[456], i_6_, i_2_, i_0_}, n_n598);
	defparam lut_1535.LUT_SIZE = 4;
	defparam lut_1535.mask = 16'h0f10;

	lut_sub lut_1537 ({sk[457], i_5_, i_6_, i_2_}, x385x);
	defparam lut_1537.LUT_SIZE = 4;
	defparam lut_1537.mask = 16'h0f40;

	lut_sub lut_1539 ({sk[458], i_5_, i_1_, i_2_, i_0_}, x42x);
	defparam lut_1539.LUT_SIZE = 5;
	defparam lut_1539.mask = 32'h0fff0301;

	lut_sub lut_1542 ({sk[459], i_10_, i_7_, i_8_}, n_n597);
	defparam lut_1542.LUT_SIZE = 4;
	defparam lut_1542.mask = 16'h0f02;

	lut_sub lut_1544 ({sk[460], i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x6590x);
	defparam lut_1544.LUT_SIZE = 7;
	defparam lut_1544.mask = 128'h0f0fffffffffffff0000000000080000;

	lut_sub lut_1546 ({sk[461], i_7_, i_13_, i_12_, x377x, x11x, n_n609}, x7980x);
	defparam lut_1546.LUT_SIZE = 7;
	defparam lut_1546.mask = 128'h0f0fffffffffffffffffeaeeffffffff;

	lut_sub lut_1560 ({sk[462], i_6_, i_0_}, x290x);
	defparam lut_1560.LUT_SIZE = 3;
	defparam lut_1560.mask = 8'h34;

	lut_sub lut_1562 ({sk[463], i_5_, i_3_, i_4_}, n_n735);
	defparam lut_1562.LUT_SIZE = 4;
	defparam lut_1562.mask = 16'h0f80;

	lut_sub lut_1564 ({sk[464], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x391x);
	defparam lut_1564.LUT_SIZE = 7;
	defparam lut_1564.mask = 128'h0f0fffffffffffff0000800000000000;

	lut_sub lut_1566 ({sk[465], i_5_, i_6_, i_3_}, n_n653);
	defparam lut_1566.LUT_SIZE = 4;
	defparam lut_1566.mask = 16'h0f80;

	lut_sub lut_1568 ({sk[466], i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x469x);
	defparam lut_1568.LUT_SIZE = 7;
	defparam lut_1568.mask = 128'h0f0fffffffffffff2000000000000100;

	lut_sub lut_1571 ({sk[467], i_7_, i_8_, i_1_, i_2_, i_0_}, x6601x);
	defparam lut_1571.LUT_SIZE = 6;
	defparam lut_1571.mask = 64'h5577ffff80000000;

	lut_sub lut_1573 ({sk[468], i_8_, i_5_, i_6_, i_3_, x25x, n_n840}, x7978x);
	defparam lut_1573.LUT_SIZE = 7;
	defparam lut_1573.mask = 128'h0f0fffffffffffffffefffffffffffff;

	lut_sub lut_1589 ({sk[469], i_3_, i_4_, i_2_}, n_n672);
	defparam lut_1589.LUT_SIZE = 4;
	defparam lut_1589.mask = 16'h0f20;

	lut_sub lut_1591 ({sk[470], i_13_, i_1_}, x32x);
	defparam lut_1591.LUT_SIZE = 3;
	defparam lut_1591.mask = 8'h34;

	lut_sub lut_1593 ({sk[471], i_9_, i_10_, i_13_, i_12_, i_11_}, x305x);
	defparam lut_1593.LUT_SIZE = 6;
	defparam lut_1593.mask = 64'h5577ffff80000000;

	lut_sub lut_1595 ({sk[472], i_9_, i_10_, i_7_, i_12_, i_2_}, x407x);
	defparam lut_1595.LUT_SIZE = 6;
	defparam lut_1595.mask = 64'h5577ffff08000000;

	lut_sub lut_1597 ({sk[473], i_10_, i_7_, i_8_, i_6_, i_3_, i_2_}, x43x);
	defparam lut_1597.LUT_SIZE = 7;
	defparam lut_1597.mask = 128'h0f0fffffffffffffe0c0a00000000000;

	lut_sub lut_1600 ({sk[474], i_10_, i_7_, i_8_, i_6_, i_3_, i_2_}, x470x);
	defparam lut_1600.LUT_SIZE = 7;
	defparam lut_1600.mask = 128'h0f0ffffffffffffff0c0a00000000000;

	lut_sub lut_1604 ({sk[475], i_6_, i_1_, x9x, n_n849, x96x, x305x}, x6855x);
	defparam lut_1604.LUT_SIZE = 7;
	defparam lut_1604.mask = 128'h0f0fffffffffffff00001111000f111f;

	lut_sub lut_1607 ({sk[476], i_8_, i_6_, i_3_}, x6853x);
	defparam lut_1607.LUT_SIZE = 4;
	defparam lut_1607.mask = 16'h0f20;

	lut_sub lut_1609 ({sk[477], i_10_, i_6_, i_13_, i_11_}, x6854x);
	defparam lut_1609.LUT_SIZE = 5;
	defparam lut_1609.mask = 32'h0fff4000;

	lut_sub lut_1611 ({sk[478], i_13_, i_4_, i_1_}, x371x);
	defparam lut_1611.LUT_SIZE = 4;
	defparam lut_1611.mask = 16'h0f10;

	lut_sub lut_1613 ({sk[479], i_9_, i_8_, i_6_, i_3_, i_2_}, x412x);
	defparam lut_1613.LUT_SIZE = 6;
	defparam lut_1613.mask = 64'h5577ffff08000000;

	lut_sub lut_1615 ({sk[480], i_9_, i_7_, i_8_, i_3_, i_2_}, x474x);
	defparam lut_1615.LUT_SIZE = 6;
	defparam lut_1615.mask = 64'h5577ffffaac00000;

	lut_sub lut_1618 ({sk[481], i_9_, i_8_, i_6_, i_13_, i_4_, i_11_}, x471x);
	defparam lut_1618.LUT_SIZE = 7;
	defparam lut_1618.mask = 128'h0f0fffffffffffff00b0003000000000;

	lut_sub lut_1621 ({sk[482], i_9_, i_3_, i_4_, i_2_}, x346x);
	defparam lut_1621.LUT_SIZE = 5;
	defparam lut_1621.mask = 32'h0fff2000;

	lut_sub lut_1623 ({sk[483], i_3_, i_1_, i_2_}, n_n534);
	defparam lut_1623.LUT_SIZE = 4;
	defparam lut_1623.mask = 16'h0f04;

	lut_sub lut_1625 ({sk[484], i_10_, i_7_, i_11_}, n_n242);
	defparam lut_1625.LUT_SIZE = 4;
	defparam lut_1625.mask = 16'h0f80;

	lut_sub lut_1627 ({sk[485], i_4_, i_1_, i_2_}, n_n346);
	defparam lut_1627.LUT_SIZE = 4;
	defparam lut_1627.mask = 16'h0f10;

	lut_sub lut_1629 ({sk[486], i_4_, i_1_}, x281x);
	defparam lut_1629.LUT_SIZE = 3;
	defparam lut_1629.mask = 8'h32;

	lut_sub lut_1631 ({sk[487], i_5_, i_3_, i_4_}, n_n846);
	defparam lut_1631.LUT_SIZE = 4;
	defparam lut_1631.mask = 16'h0f01;

	lut_sub lut_1633 ({sk[488], i_5_, i_3_, i_4_}, n_n851);
	defparam lut_1633.LUT_SIZE = 4;
	defparam lut_1633.mask = 16'h0f10;

	lut_sub lut_1635 ({sk[489], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x479x);
	defparam lut_1635.LUT_SIZE = 7;
	defparam lut_1635.mask = 128'h0f0fffffffffffff0000002000000010;

	lut_sub lut_1638 ({sk[490], i_8_, x409x, x268x, n_n755, n_n851, x479x}, x1503x);
	defparam lut_1638.LUT_SIZE = 7;
	defparam lut_1638.mask = 128'h0f0fffffffffffff0000030300050307;

	lut_sub lut_1641 ({sk[491], i_3_, i_2_, i_0_}, n_n670);
	defparam lut_1641.LUT_SIZE = 4;
	defparam lut_1641.mask = 16'h0f40;

	lut_sub lut_1643 ({sk[492], i_3_, i_1_, i_2_, i_0_}, x6669x);
	defparam lut_1643.LUT_SIZE = 5;
	defparam lut_1643.mask = 32'h0fff8000;

	lut_sub lut_1645 ({sk[493], i_10_, i_6_, i_3_, i_2_, i_0_}, x399x);
	defparam lut_1645.LUT_SIZE = 6;
	defparam lut_1645.mask = 64'h5577ffff80000000;

	lut_sub lut_1647 ({sk[494], i_5_, i_6_, i_3_, i_2_, i_0_}, x480x);
	defparam lut_1647.LUT_SIZE = 6;
	defparam lut_1647.mask = 64'h5577ffffc0008000;

	lut_sub lut_1650 ({sk[495], i_9_, i_6_, i_3_, i_4_, i_2_, i_0_}, x110x);
	defparam lut_1650.LUT_SIZE = 7;
	defparam lut_1650.mask = 128'h0f0fffffffffffff0000080000000000;

	lut_sub lut_1652 ({sk[496], i_10_, i_5_, i_6_, i_3_, i_4_, i_2_}, x111x);
	defparam lut_1652.LUT_SIZE = 7;
	defparam lut_1652.mask = 128'h0f0fffffffffffff2000000000000000;

	lut_sub lut_1654 ({sk[497], x12x, n_n853, x346x, x109x, x110x, x111x}, x1584x);
	defparam lut_1654.LUT_SIZE = 7;
	defparam lut_1654.mask = 128'h0f0fffffffffffff00007f7f00007fff;

	lut_sub lut_1659 ({sk[498], i_9_, i_13_, i_12_}, n_n550);
	defparam lut_1659.LUT_SIZE = 4;
	defparam lut_1659.mask = 16'h0f80;

	lut_sub lut_1661 ({sk[499], i_3_, i_4_}, x277x);
	defparam lut_1661.LUT_SIZE = 3;
	defparam lut_1661.mask = 8'h38;

	lut_sub lut_1663 ({sk[500], i_5_, i_3_, i_4_}, n_n732);
	defparam lut_1663.LUT_SIZE = 4;
	defparam lut_1663.mask = 16'h0f08;

	lut_sub lut_1665 ({sk[501], i_9_, i_13_, i_12_, i_11_}, x284x);
	defparam lut_1665.LUT_SIZE = 5;
	defparam lut_1665.mask = 32'h0fff4000;

	lut_sub lut_1667 ({sk[502], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x484x);
	defparam lut_1667.LUT_SIZE = 7;
	defparam lut_1667.mask = 128'h0f0fffffffffffff0800000004000000;

	lut_sub lut_1670 ({sk[503], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x6613x);
	defparam lut_1670.LUT_SIZE = 7;
	defparam lut_1670.mask = 128'h0f0fffffffffffff0000400000000000;

	lut_sub lut_1672 ({sk[504], i_13_, i_12_, i_11_}, x118x);
	defparam lut_1672.LUT_SIZE = 4;
	defparam lut_1672.mask = 16'h0f08;

	lut_sub lut_1674 ({sk[505], i_9_, i_10_, i_6_, i_13_, i_12_, i_1_}, x6873x);
	defparam lut_1674.LUT_SIZE = 7;
	defparam lut_1674.mask = 128'h0f0fffffffffffff00000500000d050d;

	lut_sub lut_1679 ({sk[506], i_10_, i_6_, i_13_, i_12_, i_1_, i_11_}, x6872x);
	defparam lut_1679.LUT_SIZE = 7;
	defparam lut_1679.mask = 128'h0f0fffffffffffff0088008000aa0080;

	lut_sub lut_1683 ({sk[507], i_4_, i_1_}, x22x);
	defparam lut_1683.LUT_SIZE = 3;
	defparam lut_1683.mask = 8'h34;

	lut_sub lut_1685 ({sk[508], i_4_, i_12_, i_11_}, x297x);
	defparam lut_1685.LUT_SIZE = 4;
	defparam lut_1685.mask = 16'h0f40;

	lut_sub lut_1687 ({sk[509], i_9_, i_10_, i_7_, i_8_, i_6_}, x490x);
	defparam lut_1687.LUT_SIZE = 6;
	defparam lut_1687.mask = 64'h5577ffff008040c0;

	lut_sub lut_1691 ({sk[510], i_9_, i_10_, i_8_, i_6_, i_11_}, x489x);
	defparam lut_1691.LUT_SIZE = 6;
	defparam lut_1691.mask = 64'h5577ffff00401050;

	lut_sub lut_1694 ({sk[511], i_9_, i_1_, x289x, x14x, n_n311, x489x}, x6881x);
	defparam lut_1694.LUT_SIZE = 7;
	defparam lut_1694.mask = 128'h0f0fffffffffffff0003050500030507;

	lut_sub lut_1698 ({sk[512], i_12_, i_2_}, x332x);
	defparam lut_1698.LUT_SIZE = 3;
	defparam lut_1698.mask = 8'h34;

	lut_sub lut_1700 ({sk[513], i_9_, i_7_, i_8_, i_6_, i_12_, i_11_}, x1287x);
	defparam lut_1700.LUT_SIZE = 7;
	defparam lut_1700.mask = 128'h0f0fffffffffffff0000000000040000;

	lut_sub lut_1702 ({sk[514], i_7_, i_8_, i_6_}, n_n837);
	defparam lut_1702.LUT_SIZE = 4;
	defparam lut_1702.mask = 16'h0f04;

	lut_sub lut_1704 ({sk[515], i_10_, i_7_, i_8_}, n_n240);
	defparam lut_1704.LUT_SIZE = 4;
	defparam lut_1704.mask = 16'h0f40;

	lut_sub lut_1706 ({sk[516], i_4_, i_2_}, x330x);
	defparam lut_1706.LUT_SIZE = 3;
	defparam lut_1706.mask = 8'h32;

	lut_sub lut_1708 ({sk[517], i_5_, i_6_, i_2_}, n_n606);
	defparam lut_1708.LUT_SIZE = 4;
	defparam lut_1708.mask = 16'h0f80;

	lut_sub lut_1710 ({sk[518], x12x, n_n853, x17x, n_n791, x295x, x263x}, x7987x);
	defparam lut_1710.LUT_SIZE = 7;
	defparam lut_1710.mask = 128'h0f0fffffffffffff00550f5f33773f7f;

	lut_sub lut_1721 ({sk[519], i_5_, i_1_, x17x, x37x, x36x, x7987x}, x495x);
	defparam lut_1721.LUT_SIZE = 7;
	defparam lut_1721.mask = 128'h0f0fffffffffffff5757575757ff5f5f;

	lut_sub lut_1726 ({sk[520], i_5_, i_1_, i_2_, i_0_, n_n769, x309x}, x7985x);
	defparam lut_1726.LUT_SIZE = 7;
	defparam lut_1726.mask = 128'h0f0ffffffffffffffffcfffcfffcffa8;

	lut_sub lut_1734 ({sk[521], i_10_, i_4_, n_n761, n_n844, x318x, x7985x}, x6752x);
	defparam lut_1734.LUT_SIZE = 7;
	defparam lut_1734.mask = 128'h0f0fffffffffffff000300ab00000000;

	lut_sub lut_1737 ({sk[522], i_10_, i_5_, i_11_}, x360x);
	defparam lut_1737.LUT_SIZE = 4;
	defparam lut_1737.mask = 16'h0f08;

	lut_sub lut_1739 ({sk[523], i_9_, i_6_, i_2_, n_n658, n_n665, n_n671}, x1637x);
	defparam lut_1739.LUT_SIZE = 7;
	defparam lut_1739.mask = 128'h0f0fffffffffffff0000000003001311;

	lut_sub lut_1742 ({sk[524], i_5_, i_6_, i_3_, i_1_, i_0_}, x500x);
	defparam lut_1742.LUT_SIZE = 6;
	defparam lut_1742.mask = 64'h5577ffff8080c0f0;

	lut_sub lut_1746 ({sk[525], i_9_, i_5_, i_3_, i_0_, n_n675, n_n358}, x7989x);
	defparam lut_1746.LUT_SIZE = 7;
	defparam lut_1746.mask = 128'h0f0fffffffffffffafffafffafff8ccc;

	lut_sub lut_1756 ({sk[526], i_9_, i_7_, i_13_, i_12_, x500x, x7989x}, x1638x);
	defparam lut_1756.LUT_SIZE = 7;
	defparam lut_1756.mask = 128'h0f0fffffffffffff00a000a000a000b0;

	lut_sub lut_1759 ({sk[527], i_3_, n_n675, n_n835, n_n665, x118x, x360x}, x6641x);
	defparam lut_1759.LUT_SIZE = 7;
	defparam lut_1759.mask = 128'h0f0fffffffffffff0033053700000505;

	lut_sub lut_1762 ({sk[528], i_10_, i_13_, i_12_, i_11_}, x294x);
	defparam lut_1762.LUT_SIZE = 5;
	defparam lut_1762.mask = 32'h0fff4000;

	lut_sub lut_1764 ({sk[529], i_4_, i_1_, i_2_, i_0_}, x296x);
	defparam lut_1764.LUT_SIZE = 5;
	defparam lut_1764.mask = 32'h0fff0100;

	lut_sub lut_1766 ({sk[530], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x501x);
	defparam lut_1766.LUT_SIZE = 7;
	defparam lut_1766.mask = 128'h0f0fffffffffffff2000000010000000;

	lut_sub lut_1769 ({sk[531], i_3_, i_4_, i_1_, i_2_}, x272x);
	defparam lut_1769.LUT_SIZE = 5;
	defparam lut_1769.mask = 32'h0fff0010;

	lut_sub lut_1771 ({sk[532], i_3_, i_4_, i_1_, i_2_}, x298x);
	defparam lut_1771.LUT_SIZE = 5;
	defparam lut_1771.mask = 32'h0fff0040;

	lut_sub lut_1773 ({sk[533], i_9_, i_3_, i_4_, i_12_, i_1_, i_2_}, x1274x);
	defparam lut_1773.LUT_SIZE = 7;
	defparam lut_1773.mask = 128'h0f0fffffffffffff0000000000005100;

	lut_sub lut_1776 ({sk[534], i_9_, i_10_, i_6_, i_12_, i_11_}, x504x);
	defparam lut_1776.LUT_SIZE = 6;
	defparam lut_1776.mask = 64'h5577ffff00100011;

	lut_sub lut_1779 ({sk[535], i_9_, i_12_, i_11_}, x334x);
	defparam lut_1779.LUT_SIZE = 4;
	defparam lut_1779.mask = 16'h0f01;

	lut_sub lut_1781 ({sk[536], i_6_, i_12_, x22x, x298x, x1274x, x334x}, x1268x);
	defparam lut_1781.LUT_SIZE = 7;
	defparam lut_1781.mask = 128'h0f0fffffffffffff000000003f7f3377;

	lut_sub lut_1785 ({sk[537], i_10_, i_6_, i_3_, i_11_, x14x, x272x}, x7973x);
	defparam lut_1785.LUT_SIZE = 7;
	defparam lut_1785.mask = 128'h0f0fffffffffffffffffffffaa8affff;

	lut_sub lut_1791 ({sk[538], i_4_, i_1_, n_n526, n_n534, x504x, x7973x}, x6896x);
	defparam lut_1791.LUT_SIZE = 7;
	defparam lut_1791.mask = 128'h0f0fffffffffffffaaafbbbfaaaaaaaa;

	lut_sub lut_1795 ({sk[539], i_9_, i_8_, i_12_}, x270x);
	defparam lut_1795.LUT_SIZE = 4;
	defparam lut_1795.mask = 16'h0f01;

	lut_sub lut_1797 ({sk[540], i_10_, i_3_, i_12_, i_1_, i_11_, i_2_}, x509x);
	defparam lut_1797.LUT_SIZE = 7;
	defparam lut_1797.mask = 128'h0f0fffffffffffff0000000000000507;

	lut_sub lut_1800 ({sk[541], i_10_, i_7_, i_8_, i_3_, i_12_, i_1_}, x1262x);
	defparam lut_1800.LUT_SIZE = 7;
	defparam lut_1800.mask = 128'h0f0fffffffffffff0000000000000100;

	lut_sub lut_1802 ({sk[542], i_8_, i_3_, i_2_, n_n453, x509x, x1262x}, x508x);
	defparam lut_1802.LUT_SIZE = 7;
	defparam lut_1802.mask = 128'h0f0fffffffffffff7777777f55555555;

	lut_sub lut_1806 ({sk[543], i_10_, i_3_, x325x, x27x, n_n311, x1256x}, x6903x);
	defparam lut_1806.LUT_SIZE = 7;
	defparam lut_1806.mask = 128'h0f0fffffffffffff5555555555555557;

	lut_sub lut_1809 ({sk[544], i_9_, i_6_, i_11_, x15x, n_n415, x270x}, x6904x);
	defparam lut_1809.LUT_SIZE = 7;
	defparam lut_1809.mask = 128'h0f0fffffffffffff0000000503030307;

	lut_sub lut_1812 ({sk[545], i_10_, i_7_, i_8_, i_6_}, x364x);
	defparam lut_1812.LUT_SIZE = 5;
	defparam lut_1812.mask = 32'h0fff0080;

	lut_sub lut_1814 ({sk[546], i_3_, i_12_, i_1_, i_2_}, x512x);
	defparam lut_1814.LUT_SIZE = 5;
	defparam lut_1814.mask = 32'h0fff0051;

	lut_sub lut_1817 ({sk[547], i_6_, i_3_, i_12_, i_1_, i_11_}, x511x);
	defparam lut_1817.LUT_SIZE = 6;
	defparam lut_1817.mask = 64'h5577ffff00080003;

	lut_sub lut_1820 ({sk[548], i_7_, i_6_, i_3_, i_12_, i_1_}, x510x);
	defparam lut_1820.LUT_SIZE = 6;
	defparam lut_1820.mask = 64'h5577ffff050d0000;

	lut_sub lut_1823 ({sk[549], i_9_, i_10_, i_11_, x15x, x364x, x510x}, x6910x);
	defparam lut_1823.LUT_SIZE = 7;
	defparam lut_1823.mask = 128'h0f0fffffffffffff0003000300030057;

	lut_sub lut_1826 ({sk[550], i_6_, i_12_, i_11_, x18x, n_n534, x512x}, x6909x);
	defparam lut_1826.LUT_SIZE = 7;
	defparam lut_1826.mask = 128'h0f0fffffffffffff0300030007050505;

	lut_sub lut_1830 ({sk[551], i_6_, i_12_, i_1_, i_11_, i_2_, x25x}, x6916x);
	defparam lut_1830.LUT_SIZE = 7;
	defparam lut_1830.mask = 128'h0f0fffffffffffff1000100011110011;

	lut_sub lut_1835 ({sk[552], i_9_, i_10_, x33x, n_n609, x6913x, x1234x}, x6917x);
	defparam lut_1835.LUT_SIZE = 7;
	defparam lut_1835.mask = 128'h0f0fffffffffffff57575757575757ff;

	lut_sub lut_1839 ({sk[553], i_5_, i_3_, i_4_}, n_n710);
	defparam lut_1839.LUT_SIZE = 4;
	defparam lut_1839.mask = 16'h0f40;

	lut_sub lut_1841 ({sk[554], i_5_, i_3_, i_13_, i_4_, i_12_, i_11_}, x6650x);
	defparam lut_1841.LUT_SIZE = 7;
	defparam lut_1841.mask = 128'h0f0fffffffffffff0000000020000000;

	lut_sub lut_1843 ({sk[555], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x520x);
	defparam lut_1843.LUT_SIZE = 7;
	defparam lut_1843.mask = 128'h0f0fffffffffffff0220000000000000;

	lut_sub lut_1846 ({sk[556], i_7_, i_8_, i_1_}, x6647x);
	defparam lut_1846.LUT_SIZE = 4;
	defparam lut_1846.mask = 16'h0f04;

	lut_sub lut_1848 ({sk[557], i_9_, i_13_, i_1_, i_11_, i_2_, i_0_}, x6648x);
	defparam lut_1848.LUT_SIZE = 7;
	defparam lut_1848.mask = 128'h0f0fffffffffffff0010000000000000;

	lut_sub lut_1850 ({sk[558], n_n725, x303x, n_n837, x520x, x6647x, x6648x}, x519x);
	defparam lut_1850.LUT_SIZE = 7;
	defparam lut_1850.mask = 128'h0f0fffffffffffff005533770f5f3f7f;

	lut_sub lut_1854 ({sk[559], i_7_, i_8_, i_6_, i_3_, i_4_, i_1_}, x518x);
	defparam lut_1854.LUT_SIZE = 7;
	defparam lut_1854.mask = 128'h0f0fffffffffffff0000000040c00000;

	lut_sub lut_1857 ({sk[560], i_0_, n_n844, x303x, n_n729, x518x, x7988x}, x6651x);
	defparam lut_1857.LUT_SIZE = 7;
	defparam lut_1857.mask = 128'h0f0fffffffffffff00000a0a00330a3b;

	lut_sub lut_1860 ({sk[561], i_9_, i_10_, i_8_, i_3_, i_11_}, x392x);
	defparam lut_1860.LUT_SIZE = 6;
	defparam lut_1860.mask = 64'h5577ffff80000000;

	lut_sub lut_1862 ({sk[562], i_8_, i_5_, i_6_, i_3_, i_0_}, x522x);
	defparam lut_1862.LUT_SIZE = 6;
	defparam lut_1862.mask = 64'h5577ffff040c0000;

	lut_sub lut_1865 ({sk[563], i_5_, i_13_, i_12_, n_n346, x296x, x392x}, x1474x);
	defparam lut_1865.LUT_SIZE = 7;
	defparam lut_1865.mask = 128'h0f0fffffffffffff1111000011150000;

	lut_sub lut_1868 ({sk[564], i_7_, i_8_, i_6_, n_n755, x525x, x524x}, x1475x);
	defparam lut_1868.LUT_SIZE = 7;
	defparam lut_1868.mask = 128'h0f0fffffffffffff0000030500000000;

	lut_sub lut_1871 ({sk[565], i_0_, n_n853, x265x, x406x, x318x, x1510x}, x1504x);
	defparam lut_1871.LUT_SIZE = 7;
	defparam lut_1871.mask = 128'h0f0fffffffffffff00005f7f00005f5f;

	lut_sub lut_1875 ({sk[566], i_2_, x17x, x37x, x322x, x6743x, x7984x}, x6745x);
	defparam lut_1875.LUT_SIZE = 7;
	defparam lut_1875.mask = 128'h0f0fffffffffffffaabbafbfaabbaabb;

	lut_sub lut_1879 ({sk[567], n_n725, x14x, n_n735, x303x, x522x, x6753x}, x6757x);
	defparam lut_1879.LUT_SIZE = 7;
	defparam lut_1879.mask = 128'h0f0fffffffffffff0000030300550357;

	lut_sub lut_1882 ({sk[568], i_10_, i_8_, i_13_, i_4_, i_12_}, x49x);
	defparam lut_1882.LUT_SIZE = 6;
	defparam lut_1882.mask = 64'h5577ffff30b00000;

	lut_sub lut_1885 ({sk[569], i_7_, i_5_, i_6_, i_2_}, x350x);
	defparam lut_1885.LUT_SIZE = 5;
	defparam lut_1885.mask = 32'h0fff0080;

	lut_sub lut_1887 ({sk[570], i_10_, i_7_, i_5_, i_13_, i_11_}, x963x);
	defparam lut_1887.LUT_SIZE = 6;
	defparam lut_1887.mask = 64'h5577ffff80000000;

	lut_sub lut_1889 ({sk[571], i_10_, i_7_, i_8_, i_3_, n_n570, n_n729}, x7964x);
	defparam lut_1889.LUT_SIZE = 7;
	defparam lut_1889.mask = 128'h0f0fffffffffffffafcf8cccafffafff;

	lut_sub lut_1898 ({sk[572], i_5_, i_3_, i_4_, n_n842, x963x, x7964x}, x528x);
	defparam lut_1898.LUT_SIZE = 7;
	defparam lut_1898.mask = 128'h0f0fffffffffffffbbbfbbbb33333333;

	lut_sub lut_1902 ({sk[573], i_10_, i_7_, i_8_, i_6_, i_13_, i_12_}, x952x);
	defparam lut_1902.LUT_SIZE = 7;
	defparam lut_1902.mask = 128'h0f0fffffffffffff0080000000000000;

	lut_sub lut_1904 ({sk[574], i_10_, i_7_, i_8_}, n_n651);
	defparam lut_1904.LUT_SIZE = 4;
	defparam lut_1904.mask = 16'h0f01;

	lut_sub lut_1906 ({sk[575], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x542x);
	defparam lut_1906.LUT_SIZE = 7;
	defparam lut_1906.mask = 128'h0f0fffffffffffff4000000010010000;

	lut_sub lut_1910 ({sk[576], i_13_, i_1_, i_11_, i_2_, i_0_}, x6664x);
	defparam lut_1910.LUT_SIZE = 6;
	defparam lut_1910.mask = 64'h5577ffff08000000;

	lut_sub lut_1912 ({sk[577], i_9_, i_7_, i_5_, i_6_, i_3_, i_4_}, x1607x);
	defparam lut_1912.LUT_SIZE = 7;
	defparam lut_1912.mask = 128'h0f0fffffffffffff0000000800000000;

	lut_sub lut_1914 ({sk[578], i_5_, i_11_, n_n570, n_n699, x277x, x1607x}, x1604x);
	defparam lut_1914.LUT_SIZE = 7;
	defparam lut_1914.mask = 128'h0f0fffffffffffff0057000000550000;

	lut_sub lut_1917 ({sk[579], i_5_, i_3_, i_4_, n_n849, n_n746, x305x}, x6663x);
	defparam lut_1917.LUT_SIZE = 7;
	defparam lut_1917.mask = 128'h0f0fffffffffffff5503000055000000;

	lut_sub lut_1920 ({sk[580], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x544x);
	defparam lut_1920.LUT_SIZE = 7;
	defparam lut_1920.mask = 128'h0f0fffffffffffff0008000000040000;

	lut_sub lut_1923 ({sk[581], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x543x);
	defparam lut_1923.LUT_SIZE = 7;
	defparam lut_1923.mask = 128'h0f0fffffffffffff0010000000200000;

	lut_sub lut_1926 ({sk[582], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x573x);
	defparam lut_1926.LUT_SIZE = 7;
	defparam lut_1926.mask = 128'h0f0fffffffffffff0000020000000800;

	lut_sub lut_1929 ({sk[583], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x572x);
	defparam lut_1929.LUT_SIZE = 7;
	defparam lut_1929.mask = 128'h0f0fffffffffffff0000000000000440;

	lut_sub lut_1932 ({sk[584], i_5_, i_3_, i_4_, n_n849, x573x, x572x}, x1570x);
	defparam lut_1932.LUT_SIZE = 7;
	defparam lut_1932.mask = 128'h0f0fffffffffffff0005000000030000;

	lut_sub lut_1935 ({sk[585], i_10_, i_7_, i_6_, i_13_, i_12_, i_11_}, x6684x);
	defparam lut_1935.LUT_SIZE = 7;
	defparam lut_1935.mask = 128'h0f0fffffffffffff1000000000000000;

	lut_sub lut_1937 ({sk[586], i_6_, x17x, n_n822, x24x, n_n670, x6669x}, x6676x);
	defparam lut_1937.LUT_SIZE = 7;
	defparam lut_1937.mask = 128'h0f0fffffffffffff0003555700005555;

	lut_sub lut_1940 ({sk[587], i_13_, i_12_, x17x, n_n453, x399x, x480x}, x6677x);
	defparam lut_1940.LUT_SIZE = 7;
	defparam lut_1940.mask = 128'h0f0fffffffffffff0033003305370033;

	lut_sub lut_1943 ({sk[588], i_7_, i_5_, x313x, x17x, n_n685, x6679x}, x6681x);
	defparam lut_1943.LUT_SIZE = 7;
	defparam lut_1943.mask = 128'h0f0fffffffffffff0537050505050505;

	lut_sub lut_1946 ({sk[589], n_n822, x24x, n_n712, n_n752, x6680x, x570x}, x6682x);
	defparam lut_1946.LUT_SIZE = 7;
	defparam lut_1946.mask = 128'h0f0fffffffffffff0003000300035557;

	lut_sub lut_1949 ({sk[590], i_5_, i_6_, i_1_, i_2_, i_0_}, x551x);
	defparam lut_1949.LUT_SIZE = 6;
	defparam lut_1949.mask = 64'h5577ffff00400800;

	lut_sub lut_1952 ({sk[591], i_10_, i_7_, i_8_, i_5_, i_6_}, x6700x);
	defparam lut_1952.LUT_SIZE = 6;
	defparam lut_1952.mask = 64'h5577ffff00000200;

	lut_sub lut_1954 ({sk[592], i_3_, i_0_, x33x, n_n651, x551x, x6700x}, x1555x);
	defparam lut_1954.LUT_SIZE = 7;
	defparam lut_1954.mask = 128'h0f0fffffffffffff0357030300000000;

	lut_sub lut_1957 ({sk[593], i_5_, i_6_, i_3_, i_1_, i_0_}, x549x);
	defparam lut_1957.LUT_SIZE = 6;
	defparam lut_1957.mask = 64'h5577fffff0c0a080;

	lut_sub lut_1962 ({sk[594], i_7_, i_8_, i_5_, i_6_, i_3_}, x6696x);
	defparam lut_1962.LUT_SIZE = 6;
	defparam lut_1962.mask = 64'h5577ffff00000002;

	lut_sub lut_1964 ({sk[595], i_5_, i_6_, i_3_, i_1_, i_2_, i_0_}, x6697x);
	defparam lut_1964.LUT_SIZE = 7;
	defparam lut_1964.mask = 128'h0f0fffffffffffff0400000000000000;

	lut_sub lut_1966 ({sk[596], n_n835, n_n656, n_n651, x549x, x6696x, x6697x}, x6702x);
	defparam lut_1966.LUT_SIZE = 7;
	defparam lut_1966.mask = 128'h0f0fffffffffffff00550f5f33773f7f;

	lut_sub lut_1970 ({sk[597], i_10_, i_8_, i_12_, i_1_, i_11_}, x555x);
	defparam lut_1970.LUT_SIZE = 6;
	defparam lut_1970.mask = 64'h5577ffff0008000a;

	lut_sub lut_1973 ({sk[598], i_10_, i_7_, i_8_, i_4_, i_12_, i_1_}, x1226x);
	defparam lut_1973.LUT_SIZE = 7;
	defparam lut_1973.mask = 128'h0f0fffffffffffff0000000000000010;

	lut_sub lut_1975 ({sk[599], i_8_, i_1_, x14x, n_n318, x555x, x1226x}, x554x);
	defparam lut_1975.LUT_SIZE = 7;
	defparam lut_1975.mask = 128'h0f0fffffffffffff557755775577557f;

	lut_sub lut_1979 ({sk[600], i_9_, i_10_, i_7_, i_8_, i_6_, i_12_}, x552x);
	defparam lut_1979.LUT_SIZE = 7;
	defparam lut_1979.mask = 128'h0f0fffffffffffff0000000000010005;

	lut_sub lut_1982 ({sk[601], i_7_, i_2_}, x352x);
	defparam lut_1982.LUT_SIZE = 3;
	defparam lut_1982.mask = 8'h34;

	lut_sub lut_1984 ({sk[602], i_0_, x30x, n_n844, n_n311, x13x, x352x}, x557x);
	defparam lut_1984.LUT_SIZE = 7;
	defparam lut_1984.mask = 128'h0f0fffffffffffff010101ff000000ff;

	lut_sub lut_1987 ({sk[603], i_9_, i_10_, i_5_, i_12_, i_11_}, x46x);
	defparam lut_1987.LUT_SIZE = 6;
	defparam lut_1987.mask = 64'h5577ffff000000a8;

	lut_sub lut_1990 ({sk[604], i_9_, i_10_, i_5_, i_12_, i_1_, i_11_}, x192x);
	defparam lut_1990.LUT_SIZE = 7;
	defparam lut_1990.mask = 128'h0f0fffffffffffff0000000000002230;

	lut_sub lut_1994 ({sk[605], i_10_, i_5_, i_12_, i_0_}, x338x);
	defparam lut_1994.LUT_SIZE = 5;
	defparam lut_1994.mask = 32'h0fff0010;

	lut_sub lut_1996 ({sk[606], i_10_, i_5_, i_6_, i_1_, i_11_, i_0_}, x183x);
	defparam lut_1996.LUT_SIZE = 7;
	defparam lut_1996.mask = 128'h0f0fffffffffffff0000000008000a00;

	lut_sub lut_1999 ({sk[607], i_5_, i_6_, i_12_, i_1_, i_2_}, x559x);
	defparam lut_1999.LUT_SIZE = 6;
	defparam lut_1999.mask = 64'h5577ffff11150000;

	lut_sub lut_2002 ({sk[608], i_5_, i_12_, x285x, n_n840, n_n656, x183x}, x177x);
	defparam lut_2002.LUT_SIZE = 7;
	defparam lut_2002.mask = 128'h0f0fffffffffffff57570000575f0000;

	lut_sub lut_2006 ({sk[609], i_10_, i_5_, i_6_, i_1_, i_11_, i_0_}, x175x);
	defparam lut_2006.LUT_SIZE = 7;
	defparam lut_2006.mask = 128'h0f0fffffffffffff000000000d000000;

	lut_sub lut_2009 ({sk[610], i_2_, x269x, n_n656, x338x, x559x, x175x}, x7256x);
	defparam lut_2009.LUT_SIZE = 7;
	defparam lut_2009.mask = 128'h0f0fffffffffffff5577557755775f7f;

	lut_sub lut_2013 ({sk[611], i_9_, i_10_, i_5_, i_6_, i_12_, i_11_}, x168x);
	defparam lut_2013.LUT_SIZE = 7;
	defparam lut_2013.mask = 128'h0f0fffffffffffff0000000000000200;

	lut_sub lut_2015 ({sk[612], i_5_, i_6_, i_12_, i_11_, i_0_, x283x}, x162x);
	defparam lut_2015.LUT_SIZE = 7;
	defparam lut_2015.mask = 128'h0f0fffffffffffff0000404000005511;

	lut_sub lut_2020 ({sk[613], x8x, x264x, n_n421, x13x, n_n598, x332x}, x7260x);
	defparam lut_2020.LUT_SIZE = 7;
	defparam lut_2020.mask = 128'h0f0fffffffffffff003700370037ffff;

	lut_sub lut_2024 ({sk[614], i_9_, i_3_, i_2_, i_0_, n_n415, x7251x}, x7252x);
	defparam lut_2024.LUT_SIZE = 7;
	defparam lut_2024.mask = 128'h0f0fffffffffffff5555555555575757;

	lut_sub lut_2028 ({sk[615], i_10_, i_7_, i_3_, i_1_, i_0_}, x6679x);
	defparam lut_2028.LUT_SIZE = 6;
	defparam lut_2028.mask = 64'h5577ffff80000000;

	lut_sub lut_2030 ({sk[616], i_13_, i_12_, i_1_, i_2_, i_0_}, x6680x);
	defparam lut_2030.LUT_SIZE = 6;
	defparam lut_2030.mask = 64'h5577ffff00800000;

	lut_sub lut_2032 ({sk[617], i_7_, i_6_, i_3_, i_1_, i_0_}, x570x);
	defparam lut_2032.LUT_SIZE = 6;
	defparam lut_2032.mask = 64'h5577ffff50400000;

	lut_sub lut_2035 ({sk[618], i_10_, i_13_, n_n2368, n_n844, n_n843, n_n851}, x6773x);
	defparam lut_2035.LUT_SIZE = 7;
	defparam lut_2035.mask = 128'h0f0fffffffffffff01ff00ff00ff00ff;

	lut_sub lut_2038 ({sk[619], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x610x);
	defparam lut_2038.LUT_SIZE = 7;
	defparam lut_2038.mask = 128'h0f0fffffffffffff0220000008800000;

	lut_sub lut_2043 ({sk[620], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x609x);
	defparam lut_2043.LUT_SIZE = 7;
	defparam lut_2043.mask = 128'h0f0fffffffffffff0010000004400000;

	lut_sub lut_2047 ({sk[621], i_9_, i_5_, i_3_, i_4_, i_1_, i_0_}, x574x);
	defparam lut_2047.LUT_SIZE = 7;
	defparam lut_2047.mask = 128'h0f0fffffffffffff0003000100000000;

	lut_sub lut_2050 ({sk[622], i_5_, i_6_, i_2_}, n_n624);
	defparam lut_2050.LUT_SIZE = 4;
	defparam lut_2050.mask = 16'h0f02;

	lut_sub lut_2052 ({sk[623], i_3_, i_4_, i_12_, i_11_}, x6573x);
	defparam lut_2052.LUT_SIZE = 5;
	defparam lut_2052.mask = 32'h0fff0080;

	lut_sub lut_2054 ({sk[624], i_12_, n_n538, n_n541, n_n844, n_n843, n_n840}, x1420x);
	defparam lut_2054.LUT_SIZE = 7;
	defparam lut_2054.mask = 128'h0f0fffffffffffff0003111300030003;

	lut_sub lut_2057 ({sk[625], i_9_, i_7_, i_8_, i_6_, i_2_}, x6800x);
	defparam lut_2057.LUT_SIZE = 6;
	defparam lut_2057.mask = 64'h5577ffff20000000;

	lut_sub lut_2059 ({sk[626], n_n833, n_n538, n_n716, n_n550, n_n837, x6800x}, x6804x);
	defparam lut_2059.LUT_SIZE = 7;
	defparam lut_2059.mask = 128'h0f0fffffffffffff0000005500000357;

	lut_sub lut_2062 ({sk[627], i_5_, i_3_, i_13_, i_4_, i_12_}, x302x);
	defparam lut_2062.LUT_SIZE = 6;
	defparam lut_2062.mask = 64'h5577ffff00800000;

	lut_sub lut_2064 ({sk[628], i_5_, i_6_, i_13_, i_12_, n_n818, x272x}, x7981x);
	defparam lut_2064.LUT_SIZE = 7;
	defparam lut_2064.mask = 128'h0f0fffffffffffffffffffcfafafaf8f;

	lut_sub lut_2072 ({sk[629], i_6_, n_n637, x8x, n_n818, x384x, x7981x}, x1402x);
	defparam lut_2072.LUT_SIZE = 7;
	defparam lut_2072.mask = 128'h0f0fffffffffffff00aa00bf00aa00bb;

	lut_sub lut_2076 ({sk[630], i_5_, i_3_, i_13_, i_4_, i_12_, i_11_}, x390x);
	defparam lut_2076.LUT_SIZE = 7;
	defparam lut_2076.mask = 128'h0f0fffffffffffff0000000000002000;

	lut_sub lut_2078 ({sk[631], i_3_, i_13_, i_1_, i_2_, i_0_}, x1390x);
	defparam lut_2078.LUT_SIZE = 6;
	defparam lut_2078.mask = 64'h5577ffff00000001;

	lut_sub lut_2080 ({sk[632], i_5_, i_12_}, x276x);
	defparam lut_2080.LUT_SIZE = 3;
	defparam lut_2080.mask = 8'h32;

	lut_sub lut_2082 ({sk[633], i_9_, n_n538, n_n844, x360x, x272x, x276x}, x7213x);
	defparam lut_2082.LUT_SIZE = 7;
	defparam lut_2082.mask = 128'h0f0fffffffffffff03030303131313ff;

	lut_sub lut_2086 ({sk[634], i_7_, i_6_, i_3_, i_0_}, x123x);
	defparam lut_2086.LUT_SIZE = 5;
	defparam lut_2086.mask = 32'h0fff1000;

	lut_sub lut_2088 ({sk[635], i_3_, n_n818, x16x, n_n415, n_n318, x26x}, x596x);
	defparam lut_2088.LUT_SIZE = 7;
	defparam lut_2088.mask = 128'h0f0fffffffffffff00001111000f111f;

	lut_sub lut_2091 ({sk[636], i_9_, i_7_, i_11_}, n_n277);
	defparam lut_2091.LUT_SIZE = 4;
	defparam lut_2091.mask = 16'h0f80;

	lut_sub lut_2093 ({sk[637], i_9_, i_10_, i_3_, i_4_}, x6807x);
	defparam lut_2093.LUT_SIZE = 5;
	defparam lut_2093.mask = 32'h0fff0002;

	lut_sub lut_2095 ({sk[638], i_9_, i_10_, i_7_, i_6_, i_12_, i_11_}, x604x);
	defparam lut_2095.LUT_SIZE = 7;
	defparam lut_2095.mask = 128'h0f0fffffffffffff0000503005035533;

	lut_sub lut_2100 ({sk[639], i_9_, i_10_, i_13_, i_4_, i_11_}, x273x);
	defparam lut_2100.LUT_SIZE = 6;
	defparam lut_2100.mask = 64'h5577ffff10000000;

	lut_sub lut_2102 ({sk[640], i_9_, i_7_, i_6_, i_3_, i_0_}, x1467x);
	defparam lut_2102.LUT_SIZE = 6;
	defparam lut_2102.mask = 64'h5577ffff00010000;

	lut_sub lut_2104 ({sk[641], i_5_, i_6_, i_3_, i_2_, i_0_}, x605x);
	defparam lut_2104.LUT_SIZE = 6;
	defparam lut_2104.mask = 64'h5577ffff03000100;

	lut_sub lut_2107 ({sk[642], x37x, x15x, n_n827, x273x, x1467x, x605x}, x6766x);
	defparam lut_2107.LUT_SIZE = 7;
	defparam lut_2107.mask = 128'h0f0fffffffffffff05050505373737ff;

	lut_sub lut_2111 ({sk[643], i_3_, i_1_, i_2_, i_0_}, x292x);
	defparam lut_2111.LUT_SIZE = 5;
	defparam lut_2111.mask = 32'h0fff0001;

	lut_sub lut_2113 ({sk[644], i_9_, i_5_, i_3_, i_13_, i_4_}, x6774x);
	defparam lut_2113.LUT_SIZE = 6;
	defparam lut_2113.mask = 64'h5577ffff00040000;

	lut_sub lut_2115 ({sk[645], i_9_, i_5_, i_6_, i_3_, i_4_, i_2_}, x1448x);
	defparam lut_2115.LUT_SIZE = 7;
	defparam lut_2115.mask = 128'h0f0fffffffffffff0000000100000000;

	lut_sub lut_2117 ({sk[646], i_9_, i_10_, i_8_, i_4_, i_12_, i_2_}, x355x);
	defparam lut_2117.LUT_SIZE = 7;
	defparam lut_2117.mask = 128'h0f0fffffffffffff0000000000000010;

	lut_sub lut_2119 ({sk[647], i_10_, x27x, n_n665, x29x, x96x, x355x}, x6980x);
	defparam lut_2119.LUT_SIZE = 7;
	defparam lut_2119.mask = 128'h0f0fffffffffffff555f555f555fdddf;

	lut_sub lut_2123 ({sk[648], i_9_, i_7_, i_4_}, x351x);
	defparam lut_2123.LUT_SIZE = 4;
	defparam lut_2123.mask = 16'h0f10;

	lut_sub lut_2125 ({sk[649], i_9_, i_8_, i_3_, i_13_, i_4_, i_11_}, x618x);
	defparam lut_2125.LUT_SIZE = 7;
	defparam lut_2125.mask = 128'h0f0fffffffffffffb000300000000000;

	lut_sub lut_2128 ({sk[650], i_10_, i_7_, i_13_, i_11_, i_2_, n_n1574}, x6986x);
	defparam lut_2128.LUT_SIZE = 7;
	defparam lut_2128.mask = 128'h0f0fffffffffffff55d5555555f75555;

	lut_sub lut_2133 ({sk[651], i_10_, i_7_, i_8_, i_13_, i_12_, i_11_}, x625x);
	defparam lut_2133.LUT_SIZE = 7;
	defparam lut_2133.mask = 128'h0f0fffffffffffffa0c0000000000000;

	lut_sub lut_2137 ({sk[652], i_9_, i_8_, i_13_, i_4_}, x319x);
	defparam lut_2137.LUT_SIZE = 5;
	defparam lut_2137.mask = 32'h0fff0400;

	lut_sub lut_2139 ({sk[653], i_9_, i_8_, i_5_}, n_n768);
	defparam lut_2139.LUT_SIZE = 4;
	defparam lut_2139.mask = 16'h0f10;

	lut_sub lut_2141 ({sk[654], i_10_, i_7_, i_12_, i_11_}, x636x);
	defparam lut_2141.LUT_SIZE = 5;
	defparam lut_2141.mask = 32'h0fffa800;

	lut_sub lut_2144 ({sk[655], i_10_, i_7_, i_13_, i_12_, i_1_, i_2_}, x1193x);
	defparam lut_2144.LUT_SIZE = 7;
	defparam lut_2144.mask = 128'h0f0fffffffffffff0000200000000000;

	lut_sub lut_2146 ({sk[656], i_10_, i_7_, i_8_, i_11_, n_n570, x328x}, x7974x);
	defparam lut_2146.LUT_SIZE = 7;
	defparam lut_2146.mask = 128'h0f0fffffffffffffefeeffffffffffff;

	lut_sub lut_2160 ({sk[657], i_9_, i_5_, i_3_, i_13_, i_4_}, x877x);
	defparam lut_2160.LUT_SIZE = 6;
	defparam lut_2160.mask = 64'h5577ffff00400000;

	lut_sub lut_2162 ({sk[658], i_9_, i_8_, i_3_, x24x, n_n570, n_n719}, x7966x);
	defparam lut_2162.LUT_SIZE = 7;
	defparam lut_2162.mask = 128'h0f0fffffffffffffaaffc0f0aafff0f0;

	lut_sub lut_2170 ({sk[659], i_6_, i_3_, i_1_, i_0_}, x41x);
	defparam lut_2170.LUT_SIZE = 5;
	defparam lut_2170.mask = 32'h0fffa080;

	lut_sub lut_2173 ({sk[660], i_10_, i_7_, i_8_, i_11_}, x382x);
	defparam lut_2173.LUT_SIZE = 5;
	defparam lut_2173.mask = 32'h0fff8000;

	lut_sub lut_2175 ({sk[661], i_6_, i_0_}, x271x);
	defparam lut_2175.LUT_SIZE = 3;
	defparam lut_2175.mask = 8'h38;

	lut_sub lut_2177 ({sk[662], i_7_, i_8_, i_3_, i_1_, n_n835, x271x}, x7009x);
	defparam lut_2177.LUT_SIZE = 7;
	defparam lut_2177.mask = 128'h0f0fffffffffffff7373737373505050;

	lut_sub lut_2181 ({sk[663], i_9_, i_11_, n_n773, x289x, n_n671, x7009x}, x1076x);
	defparam lut_2181.LUT_SIZE = 7;
	defparam lut_2181.mask = 128'h0f0fffffffffffff5777000055770000;

	lut_sub lut_2185 ({sk[664], i_5_, i_3_, i_1_}, x324x);
	defparam lut_2185.LUT_SIZE = 4;
	defparam lut_2185.mask = 16'h0f80;

	lut_sub lut_2187 ({sk[665], i_9_, i_5_, i_6_, i_3_, i_1_, n_n275}, x47x);
	defparam lut_2187.LUT_SIZE = 7;
	defparam lut_2187.mask = 128'h0f0fffffffffffff0000cc4000004040;

	lut_sub lut_2190 ({sk[666], i_6_, i_3_, i_1_, i_0_, n_n275, x47x}, x7018x);
	defparam lut_2190.LUT_SIZE = 7;
	defparam lut_2190.mask = 128'h0f0fffffffffffff7555555575755555;

	lut_sub lut_2194 ({sk[667], i_5_, x265x, x31x, n_n242, n_n277, x382x}, x7020x);
	defparam lut_2194.LUT_SIZE = 7;
	defparam lut_2194.mask = 128'h0f0fffffffffffff00550f5f00003333;

	lut_sub lut_2198 ({sk[668], i_9_, i_10_, i_1_, n_n675, x11x, x357x}, x7997x);
	defparam lut_2198.LUT_SIZE = 7;
	defparam lut_2198.mask = 128'h0f0fffffffffffffc8fafafaccffffff;

	lut_sub lut_2208 ({sk[669], i_10_, i_5_, i_6_, i_11_}, x304x);
	defparam lut_2208.LUT_SIZE = 5;
	defparam lut_2208.mask = 32'h0fff0040;

	lut_sub lut_2210 ({sk[670], i_8_, i_12_, i_11_}, x356x);
	defparam lut_2210.LUT_SIZE = 4;
	defparam lut_2210.mask = 16'h0f02;

	lut_sub lut_2212 ({sk[671], i_9_, i_10_, i_5_, i_12_}, x10x);
	defparam lut_2212.LUT_SIZE = 5;
	defparam lut_2212.mask = 32'h0fff0405;

	lut_sub lut_2215 ({sk[672], i_8_, i_5_, n_n844, n_n316, n_n840, x10x}, x778x);
	defparam lut_2215.LUT_SIZE = 7;
	defparam lut_2215.mask = 128'h0f0fffffffffffff0000000003570055;

	lut_sub lut_2218 ({sk[673], i_10_, i_5_, n_n346, x296x, x270x, x356x}, x7187x);
	defparam lut_2218.LUT_SIZE = 7;
	defparam lut_2218.mask = 128'h0f0fffffffffffff0000030300550303;

	lut_sub lut_2221 ({sk[674], i_9_, i_10_, i_5_, i_12_, i_0_}, x656x);
	defparam lut_2221.LUT_SIZE = 6;
	defparam lut_2221.mask = 64'h5577ffff00100111;

	lut_sub lut_2224 ({sk[675], n_n638, n_n318, n_n316, x26x, n_n651, x36x}, x7185x);
	defparam lut_2224.LUT_SIZE = 7;
	defparam lut_2224.mask = 128'h0f0fffffffffffff0003000300035557;

	lut_sub lut_2227 ({sk[676], i_8_, i_5_, i_4_, i_1_, i_2_, i_0_}, x1089x);
	defparam lut_2227.LUT_SIZE = 7;
	defparam lut_2227.mask = 128'h0f0fffffffffffff00c0008000000000;

	lut_sub lut_2230 ({sk[677], i_7_, i_4_, i_12_, i_1_, x26x, n_n683}, x7972x);
	defparam lut_2230.LUT_SIZE = 7;
	defparam lut_2230.mask = 128'h0f0fffffffffffffcfff8aaacfffcfff;

	lut_sub lut_2240 ({sk[678], i_7_, i_8_, i_5_, i_6_, i_3_, i_11_}, x1814x);
	defparam lut_2240.LUT_SIZE = 7;
	defparam lut_2240.mask = 128'h0f0fffffffffffff5000100000000000;

	lut_sub lut_2243 ({sk[679], i_7_, i_2_, x343x, x348x, x304x, x1814x}, x6508x);
	defparam lut_2243.LUT_SIZE = 7;
	defparam lut_2243.mask = 128'h0f0fffffffffffff5fff7fff5fff5fff;

	lut_sub lut_2248 ({sk[680], i_9_, i_10_, i_6_, i_1_, i_0_}, x6505x);
	defparam lut_2248.LUT_SIZE = 6;
	defparam lut_2248.mask = 64'h5577ffff00000155;

	lut_sub lut_2251 ({sk[681], i_7_, i_3_, i_1_, i_0_}, x287x);
	defparam lut_2251.LUT_SIZE = 5;
	defparam lut_2251.mask = 32'h0fff0001;

	lut_sub lut_2253 ({sk[682], i_9_, i_10_, i_7_, i_8_, i_11_}, x662x);
	defparam lut_2253.LUT_SIZE = 6;
	defparam lut_2253.mask = 64'h5577ffff44544555;

	lut_sub lut_2257 ({sk[683], i_10_, i_7_, i_5_, i_6_, i_3_, i_4_}, x117x);
	defparam lut_2257.LUT_SIZE = 7;
	defparam lut_2257.mask = 128'h0f0fffffffffffff4000000000000000;

	lut_sub lut_2259 ({sk[684], i_5_, i_6_, i_1_, x9x, n_n849, x294x}, x7105x);
	defparam lut_2259.LUT_SIZE = 7;
	defparam lut_2259.mask = 128'h0f0fffffffffffff0000550003030303;

	lut_sub lut_2262 ({sk[685], i_13_, i_11_, x378x, x117x, x7105x}, x7107x);
	defparam lut_2262.LUT_SIZE = 6;
	defparam lut_2262.mask = 64'h5577ffff557f5555;

	lut_sub lut_2266 ({sk[686], i_9_, i_7_, i_5_, i_6_, i_3_, i_4_}, x401x);
	defparam lut_2266.LUT_SIZE = 7;
	defparam lut_2266.mask = 128'h0f0fffffffffffff0000000400000000;

	lut_sub lut_2268 ({sk[687], i_9_, i_7_, i_8_, i_5_, i_4_, i_1_}, x76x);
	defparam lut_2268.LUT_SIZE = 7;
	defparam lut_2268.mask = 128'h0f0fffffffffffff0000000200000000;

	lut_sub lut_2270 ({sk[688], i_9_, i_7_, i_5_, i_3_, i_4_, i_1_}, x403x);
	defparam lut_2270.LUT_SIZE = 7;
	defparam lut_2270.mask = 128'h0f0fffffffffffff0000002000000000;

	lut_sub lut_2272 ({sk[689], i_9_, i_8_, i_5_, i_6_, i_4_, i_2_}, x912x);
	defparam lut_2272.LUT_SIZE = 7;
	defparam lut_2272.mask = 128'h0f0fffffffffffff0000000200000000;

	lut_sub lut_2274 ({sk[690], i_5_, i_6_, i_3_, n_n716, n_n275, x47x}, x908x);
	defparam lut_2274.LUT_SIZE = 7;
	defparam lut_2274.mask = 128'h0f0fffffffffffff0505050505050705;

	lut_sub lut_2277 ({sk[691], i_9_, i_7_, i_6_, i_3_, i_4_, i_0_}, x398x);
	defparam lut_2277.LUT_SIZE = 7;
	defparam lut_2277.mask = 128'h0f0fffffffffffff0000002000000000;

	lut_sub lut_2279 ({sk[692], n_n769, n_n771, n_n835, x406x, x318x, x401x}, x7026x);
	defparam lut_2279.LUT_SIZE = 7;
	defparam lut_2279.mask = 128'h0f0fffffffffffff5f7f5f7f5f7fffff;

	lut_sub lut_2284 ({sk[693], i_5_, i_4_, i_2_, n_n769, x110x, x398x}, x7025x);
	defparam lut_2284.LUT_SIZE = 7;
	defparam lut_2284.mask = 128'h0f0fffffffffffff7777777777777f77;

	lut_sub lut_2288 ({sk[694], i_5_, i_6_, n_n764, n_n791, x346x, x7025x}, x7027x);
	defparam lut_2288.LUT_SIZE = 7;
	defparam lut_2288.mask = 128'h0f0fffffffffffff555f555f555f777f;

	lut_sub lut_2292 ({sk[695], i_9_, i_10_, i_4_, x394x, x117x, x111x}, x7031x);
	defparam lut_2292.LUT_SIZE = 7;
	defparam lut_2292.mask = 128'h0f0fffffffffffff7fff7f7f7f7f7f7f;

	lut_sub lut_2297 ({sk[696], i_5_, i_4_, i_2_, n_n773, n_n699, n_n678}, x7030x);
	defparam lut_2297.LUT_SIZE = 7;
	defparam lut_2297.mask = 128'h0f0fffffffffffff11111f1111111111;

	lut_sub lut_2300 ({sk[697], i_4_, n_n792, x11x, x399x, x271x, x7030x}, x7032x);
	defparam lut_2300.LUT_SIZE = 7;
	defparam lut_2300.mask = 128'h0f0fffffffffffff555555555f5f7fff;

	lut_sub lut_2305 ({sk[698], i_9_, i_7_, i_3_, i_4_, i_1_, i_0_}, x108x);
	defparam lut_2305.LUT_SIZE = 7;
	defparam lut_2305.mask = 128'h0f0fffffffffffff0000080000000000;

	lut_sub lut_2307 ({sk[699], i_10_, i_7_, i_8_, i_3_, i_2_}, x679x);
	defparam lut_2307.LUT_SIZE = 6;
	defparam lut_2307.mask = 64'h5577ffff0caa0000;

	lut_sub lut_2310 ({sk[700], i_9_, i_7_, i_6_, i_1_, i_2_, i_0_}, x7035x);
	defparam lut_2310.LUT_SIZE = 7;
	defparam lut_2310.mask = 128'h0f0fffffffffffff0000808800008080;

	lut_sub lut_2313 ({sk[701], n_n764, n_n683, n_n240, x271x, x679x, x7035x}, x678x);
	defparam lut_2313.LUT_SIZE = 7;
	defparam lut_2313.mask = 128'h0f0fffffffffffff575757ff5757ffff;

	lut_sub lut_2318 ({sk[702], i_12_, x7031x, x7032x, x678x}, x7040x);
	defparam lut_2318.LUT_SIZE = 5;
	defparam lut_2318.mask = 32'h0fff7f3f;

	lut_sub lut_2322 ({sk[703], i_9_, i_7_, i_6_, i_3_, i_1_, i_2_}, x6525x);
	defparam lut_2322.LUT_SIZE = 7;
	defparam lut_2322.mask = 128'h0f0fffffffffffff0101010101010155;

	lut_sub lut_2325 ({sk[704], i_11_, i_0_}, x380x);
	defparam lut_2325.LUT_SIZE = 3;
	defparam lut_2325.mask = 8'h38;

	lut_sub lut_2327 ({sk[705], i_9_, i_10_, i_8_, i_5_, i_6_, i_12_}, x686x);
	defparam lut_2327.LUT_SIZE = 7;
	defparam lut_2327.mask = 128'h0f0fffffffffffff0000000000010011;

	lut_sub lut_2330 ({sk[706], i_5_, i_3_, i_12_, i_1_, i_2_, i_0_}, x685x);
	defparam lut_2330.LUT_SIZE = 7;
	defparam lut_2330.mask = 128'h0f0fffffffffffff0000000000000301;

	lut_sub lut_2333 ({sk[707], i_9_, i_10_, i_5_, i_12_, i_11_, i_0_}, x689x);
	defparam lut_2333.LUT_SIZE = 7;
	defparam lut_2333.mask = 128'h0f0fffffffffffff0000000008000d00;

	lut_sub lut_2336 ({sk[708], i_9_, i_8_, i_5_, i_12_, i_11_}, x688x);
	defparam lut_2336.LUT_SIZE = 6;
	defparam lut_2336.mask = 64'h5577ffff000000a8;

	lut_sub lut_2339 ({sk[709], i_3_, i_0_, x33x, n_n752, x689x, x688x}, x373x);
	defparam lut_2339.LUT_SIZE = 7;
	defparam lut_2339.mask = 128'h0f0fffffffffffff0000000003570303;

	lut_sub lut_2342 ({sk[710], i_9_, i_3_, i_12_, i_2_, n_n176, x380x}, x7970x);
	defparam lut_2342.LUT_SIZE = 7;
	defparam lut_2342.mask = 128'h0f0ffffffffffffffffffffffffffffe;

	lut_sub lut_2357 ({sk[711], i_9_, i_8_, n_n818, x686x, x685x, x7970x}, x7192x);
	defparam lut_2357.LUT_SIZE = 7;
	defparam lut_2357.mask = 128'h0f0fffffffffffffaaafaaafaaafbbbf;

	lut_sub lut_2361 ({sk[712], i_9_, i_7_, i_5_, i_6_, i_2_}, x1031x);
	defparam lut_2361.LUT_SIZE = 6;
	defparam lut_2361.mask = 64'h5577ffff00020000;

	lut_sub lut_2363 ({sk[713], i_10_, i_5_, i_3_, i_2_, n_n769, x317x}, x7971x);
	defparam lut_2363.LUT_SIZE = 7;
	defparam lut_2363.mask = 128'h0f0fffffffffffffafaf8fafffffcfff;

	lut_sub lut_2371 ({sk[714], i_8_, n_n675, x274x, n_n768, x1031x, x7971x}, x692x);
	defparam lut_2371.LUT_SIZE = 7;
	defparam lut_2371.mask = 128'h0f0fffffffffffffbbbbbfbfbbffbfff;

	lut_sub lut_2376 ({sk[715], i_10_, x323x, x265x, x29x, n_n827, x350x}, x694x);
	defparam lut_2376.LUT_SIZE = 7;
	defparam lut_2376.mask = 128'h0f0fffffffffffff55775f7f00330033;

	lut_sub lut_2380 ({sk[716], i_8_, i_5_, i_3_, i_0_, x265x, x399x}, x7052x);
	defparam lut_2380.LUT_SIZE = 7;
	defparam lut_2380.mask = 128'h0f0fffffffffffff0000f0f07555f5f5;

	lut_sub lut_2384 ({sk[717], i_5_, n_n769, x31x, n_n671, n_n653, n_n240}, x7051x);
	defparam lut_2384.LUT_SIZE = 7;
	defparam lut_2384.mask = 128'h0f0fffffffffffff11551f5f11111f1f;

	lut_sub lut_2388 ({sk[718], i_6_, i_3_, i_1_, i_0_, n_n764, x7051x}, x7053x);
	defparam lut_2388.LUT_SIZE = 7;
	defparam lut_2388.mask = 128'h0f0fffffffffffff55555555f575f555;

	lut_sub lut_2392 ({sk[719], i_4_, x12x, n_n764, x31x, x276x, x263x}, x1023x);
	defparam lut_2392.LUT_SIZE = 7;
	defparam lut_2392.mask = 128'h0f0fffffffffffff00030003005700ff;

	lut_sub lut_2396 ({sk[720], i_5_, i_6_, i_3_, i_11_, n_n275, x412x}, x1011x);
	defparam lut_2396.LUT_SIZE = 7;
	defparam lut_2396.mask = 128'h0f0fffffffffffff0000000050507050;

	lut_sub lut_2399 ({sk[721], i_7_, i_8_, i_3_, i_2_, n_n741, x7047x}, x7048x);
	defparam lut_2399.LUT_SIZE = 7;
	defparam lut_2399.mask = 128'h0f0fffffffffffff7775757577555555;

	lut_sub lut_2403 ({sk[722], i_9_, i_5_, i_6_, i_11_}, x397x);
	defparam lut_2403.LUT_SIZE = 5;
	defparam lut_2403.mask = 32'h0fff0004;

	lut_sub lut_2405 ({sk[723], i_5_, i_3_, i_0_}, x366x);
	defparam lut_2405.LUT_SIZE = 4;
	defparam lut_2405.mask = 16'h0f01;

	lut_sub lut_2407 ({sk[724], i_11_, i_0_, x15x, n_n185, n_n432, n_n183}, x155x);
	defparam lut_2407.LUT_SIZE = 7;
	defparam lut_2407.mask = 128'h0f0fffffffffffff0005000300000003;

	lut_sub lut_2410 ({sk[725], i_11_, n_n826, x34x, x270x, x366x, x155x}, x7272x);
	defparam lut_2410.LUT_SIZE = 7;
	defparam lut_2410.mask = 128'h0f0fffffffffffff5555555f5757575f;

	lut_sub lut_2414 ({sk[726], i_7_, i_8_, i_5_, i_3_, i_1_, i_0_}, x146x);
	defparam lut_2414.LUT_SIZE = 7;
	defparam lut_2414.mask = 128'h0f0fffffffffffff0000000100000000;

	lut_sub lut_2416 ({sk[727], i_7_, i_5_, i_6_, n_n197, n_n598, x332x}, x7990x);
	defparam lut_2416.LUT_SIZE = 7;
	defparam lut_2416.mask = 128'h0f0ffffffffffffffffffffffffff8fc;

	lut_sub lut_2430 ({sk[728], i_9_, i_5_, i_13_, i_12_, i_0_, x7990x}, x7278x);
	defparam lut_2430.LUT_SIZE = 7;
	defparam lut_2430.mask = 128'h0f0fffffffffffffaaaaaaeaaaaaaafb;

	lut_sub lut_2434 ({sk[729], i_9_, i_8_, i_12_, i_0_, n_n637, x7999x}, x7277x);
	defparam lut_2434.LUT_SIZE = 7;
	defparam lut_2434.mask = 128'h0f0fffffffffffff300030003000baaa;

	lut_sub lut_2437 ({sk[730], i_9_, i_11_, n_n746, x146x, x366x, x7277x}, x7279x);
	defparam lut_2437.LUT_SIZE = 7;
	defparam lut_2437.mask = 128'h0f0fffffffffffff5555555555555f7f;

	lut_sub lut_2441 ({sk[731], i_5_, i_0_}, x280x);
	defparam lut_2441.LUT_SIZE = 3;
	defparam lut_2441.mask = 8'h38;

	lut_sub lut_2443 ({sk[732], i_7_, i_8_, i_6_, i_3_}, x7296x);
	defparam lut_2443.LUT_SIZE = 5;
	defparam lut_2443.mask = 32'h0fff4000;

	lut_sub lut_2445 ({sk[733], i_5_, i_12_, i_0_, x27x, x15x, x7296x}, x705x);
	defparam lut_2445.LUT_SIZE = 7;
	defparam lut_2445.mask = 128'h0f0fffffffffffff0055005557000000;

	lut_sub lut_2449 ({sk[734], i_10_, i_5_, i_13_, i_11_, i_0_}, x102x);
	defparam lut_2449.LUT_SIZE = 6;
	defparam lut_2449.mask = 64'h5577ffff08000c00;

	lut_sub lut_2452 ({sk[735], i_9_, i_10_, i_5_, i_13_, i_0_}, x7298x);
	defparam lut_2452.LUT_SIZE = 6;
	defparam lut_2452.mask = 64'h5577ffff00100011;

	lut_sub lut_2455 ({sk[736], i_9_, i_5_, n_n453, n_n665, x102x, x7298x}, x7300x);
	defparam lut_2455.LUT_SIZE = 7;
	defparam lut_2455.mask = 128'h0f0fffffffffffff77777777777f7f7f;

	lut_sub lut_2460 ({sk[737], i_9_, i_5_, i_3_, i_4_, i_1_, i_0_}, x708x);
	defparam lut_2460.LUT_SIZE = 7;
	defparam lut_2460.mask = 128'h0f0fffffffffffff0000002000000030;

	lut_sub lut_2463 ({sk[738], i_10_, i_5_, i_3_, i_4_, i_1_, i_0_}, x712x);
	defparam lut_2463.LUT_SIZE = 7;
	defparam lut_2463.mask = 128'h0f0fffffffffffff0020000000300000;

	lut_sub lut_2466 ({sk[739], i_7_, x12x, n_n183, n_n153, n_n316, x712x}, x785x);
	defparam lut_2466.LUT_SIZE = 7;
	defparam lut_2466.mask = 128'h0f0fffffffffffff000000001111111f;

	lut_sub lut_2469 ({sk[740], i_9_, i_10_, i_5_, i_12_, i_11_, i_0_}, x717x);
	defparam lut_2469.LUT_SIZE = 7;
	defparam lut_2469.mask = 128'h0f0fffffffffffff0000010000010101;

	lut_sub lut_2473 ({sk[741], i_0_, x12x, x14x, n_n176, x270x, x719x}, x256x);
	defparam lut_2473.LUT_SIZE = 7;
	defparam lut_2473.mask = 128'h0f0fffffffffffff0005000500050037;

	lut_sub lut_2476 ({sk[742], i_4_, x355x, x36x, x366x, x717x, x7193x}, x7196x);
	defparam lut_2476.LUT_SIZE = 7;
	defparam lut_2476.mask = 128'h0f0fffffffffffff373737ff050505ff;

	lut_sub lut_2480 ({sk[743], i_2_, i_0_, n_n792, n_n716, x31x, n_n699}, x865x);
	defparam lut_2480.LUT_SIZE = 7;
	defparam lut_2480.mask = 128'h0f0fffffffffffff0507000000030000;

	lut_sub lut_2483 ({sk[744], i_7_, i_8_, n_n849, x37x, n_n835, n_n791}, x7137x);
	defparam lut_2483.LUT_SIZE = 7;
	defparam lut_2483.mask = 128'h0f0fffffffffffff0357000003030000;

	lut_sub lut_2486 ({sk[745], i_7_, i_5_, i_6_, n_n849, n_n678, x862x}, x857x);
	defparam lut_2486.LUT_SIZE = 7;
	defparam lut_2486.mask = 128'h0f0fffffffffffff0000570000005500;

	lut_sub lut_2489 ({sk[746], i_8_, i_5_, i_3_, i_0_, x265x, n_n545}, x859x);
	defparam lut_2489.LUT_SIZE = 7;
	defparam lut_2489.mask = 128'h0f0fffffffffffff0000000010000000;

	lut_sub lut_2491 ({sk[747], i_7_, i_5_, x37x, n_n683, n_n710, x6664x}, x7139x);
	defparam lut_2491.LUT_SIZE = 7;
	defparam lut_2491.mask = 128'h0f0fffffffffffff1111111f11111111;

	lut_sub lut_2494 ({sk[748], i_5_, x865x, x7137x, x857x, x859x, x7139x}, n_n981);
	defparam lut_2494.LUT_SIZE = 7;
	defparam lut_2494.mask = 128'h0f0fffffffffffff7f7f7f7f7fffffff;

	lut_sub lut_2500 ({sk[749], i_5_, i_6_, i_3_, i_4_, i_2_, i_0_}, x849x);
	defparam lut_2500.LUT_SIZE = 7;
	defparam lut_2500.mask = 128'h0f0fffffffffffff0000080000000000;

	lut_sub lut_2502 ({sk[750], i_0_, n_n185, n_n176, x281x, x330x, x849x}, x7147x);
	defparam lut_2502.LUT_SIZE = 7;
	defparam lut_2502.mask = 128'h0f0fffffffffffff55775f7f55555555;

	lut_sub lut_2506 ({sk[751], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x7145x);
	defparam lut_2506.LUT_SIZE = 7;
	defparam lut_2506.mask = 128'h0f0fffffffffffff00008080000080aa;

	lut_sub lut_2509 ({sk[752], i_6_, i_0_}, x263x);
	defparam lut_2509.LUT_SIZE = 3;
	defparam lut_2509.mask = 8'h32;

	lut_sub lut_2511 ({sk[753], i_9_, i_7_, i_8_, i_5_, i_6_}, x7152x);
	defparam lut_2511.LUT_SIZE = 6;
	defparam lut_2511.mask = 64'h5577ffff00002000;

	lut_sub lut_2513 ({sk[754], n_n764, x17x, x6669x, x297x, x263x, x7152x}, x7155x);
	defparam lut_2513.LUT_SIZE = 7;
	defparam lut_2513.mask = 128'h0f0fffffffffffff050505ff050537ff;

	lut_sub lut_2517 ({sk[755], i_9_, i_8_, i_4_, i_1_, i_2_, i_0_}, x1509x);
	defparam lut_2517.LUT_SIZE = 7;
	defparam lut_2517.mask = 128'h0f0fffffffffffff0000008000000000;

	lut_sub lut_2519 ({sk[756], i_9_, i_8_, i_6_, i_4_, i_2_, i_0_}, x1510x);
	defparam lut_2519.LUT_SIZE = 7;
	defparam lut_2519.mask = 128'h0f0fffffffffffff0000000800000000;

	lut_sub lut_2521 ({sk[757], i_5_, i_4_, i_0_, n_n197, n_n843, x39x}, x837x);
	defparam lut_2521.LUT_SIZE = 7;
	defparam lut_2521.mask = 128'h0f0fffffffffffff1111000011130000;

	lut_sub lut_2524 ({sk[758], n_n853, x110x, x7155x, x1509x, x1510x, x837x}, n_n984);
	defparam lut_2524.LUT_SIZE = 7;
	defparam lut_2524.mask = 128'h0f0fffffffffffff55ff55ff7fffffff;

	lut_sub lut_2530 ({sk[759], i_8_, x267x, n_n853, x394x, n_n791, x108x}, x824x);
	defparam lut_2530.LUT_SIZE = 7;
	defparam lut_2530.mask = 128'h0f0fffffffffffff005f005f005f007f;

	lut_sub lut_2534 ({sk[760], i_10_, i_6_, i_0_, x27x, x17x, x6718x}, x7158x);
	defparam lut_2534.LUT_SIZE = 7;
	defparam lut_2534.mask = 128'h0f0fffffffffffff1311111111111111;

	lut_sub lut_2537 ({sk[761], i_10_, n_n853, x27x, x28x, n_n678, n_n791}, x7159x);
	defparam lut_2537.LUT_SIZE = 7;
	defparam lut_2537.mask = 128'h0f0fffffffffffff0000035700000000;

	lut_sub lut_2540 ({sk[762], x17x, x399x, x6679x, x824x, x7158x, x7159x}, n_n983);
	defparam lut_2540.LUT_SIZE = 7;
	defparam lut_2540.mask = 128'h0f0fffffffffffff7f7f7f7f7fffffff;

	lut_sub lut_2546 ({sk[763], i_8_, i_5_}, x357x);
	defparam lut_2546.LUT_SIZE = 3;
	defparam lut_2546.mask = 8'h34;

	lut_sub lut_2548 ({sk[764], i_9_, i_4_, i_11_}, x374x);
	defparam lut_2548.LUT_SIZE = 4;
	defparam lut_2548.mask = 16'h0f04;

	lut_sub lut_2550 ({sk[765], i_9_, i_5_, i_3_, i_4_, i_0_}, x730x);
	defparam lut_2550.LUT_SIZE = 6;
	defparam lut_2550.mask = 64'h5577ffff0008000c;

	lut_sub lut_2553 ({sk[766], i_9_, i_12_, i_11_}, x342x);
	defparam lut_2553.LUT_SIZE = 4;
	defparam lut_2553.mask = 16'h0f04;

	lut_sub lut_2555 ({sk[767], n_n197, n_n840, n_n346, x297x, x296x, x342x}, x729x);
	defparam lut_2555.LUT_SIZE = 7;
	defparam lut_2555.mask = 128'h0f0fffffffffffff00550f5f33773f7f;

	lut_sub lut_2559 ({sk[768], x288x, x28x, n_n213, n_n311, x296x, x730x}, x7205x);
	defparam lut_2559.LUT_SIZE = 7;
	defparam lut_2559.mask = 128'h0f0fffffffffffff0000050500330537;

	lut_sub lut_2562 ({sk[769], i_9_, i_3_, i_11_, n_n570, n_n819, n_n752}, x803x);
	defparam lut_2562.LUT_SIZE = 7;
	defparam lut_2562.mask = 128'h0f0fffffffffffff0705000003000000;

	lut_sub lut_2565 ({sk[770], i_9_, i_10_, i_5_, i_6_, i_12_, i_11_}, x737x);
	defparam lut_2565.LUT_SIZE = 7;
	defparam lut_2565.mask = 128'h0f0fffffffffffff0000030000530353;

	lut_sub lut_2570 ({sk[771], i_6_, i_12_, i_1_, i_11_, i_2_, i_0_}, x7220x);
	defparam lut_2570.LUT_SIZE = 7;
	defparam lut_2570.mask = 128'h0f0fffffffffffff0020002000202020;

	lut_sub lut_2573 ({sk[772], i_10_, i_1_, i_2_, i_0_, n_n541, x7220x}, x227x);
	defparam lut_2573.LUT_SIZE = 7;
	defparam lut_2573.mask = 128'h0f0fffffffffffff1111111111111113;

	lut_sub lut_2576 ({sk[773], i_10_, i_5_, i_6_, i_12_, i_11_, n_n412}, x7969x);
	defparam lut_2576.LUT_SIZE = 7;
	defparam lut_2576.mask = 128'h0f0ffffffffffffffffffffffffbffff;

	lut_sub lut_2592 ({sk[774], i_4_, n_n818, n_n844, x6807x, x737x, x7969x}, x7222x);
	defparam lut_2592.LUT_SIZE = 7;
	defparam lut_2592.mask = 128'h0f0fffffffffffffaaafbbbfaaafaaaf;

	lut_sub lut_2596 ({sk[775], i_9_, i_7_, i_8_, i_5_}, x741x);
	defparam lut_2596.LUT_SIZE = 5;
	defparam lut_2596.mask = 32'h0fff0203;

	lut_sub lut_2599 ({sk[776], i_10_, i_7_, i_8_, i_5_, i_0_}, x740x);
	defparam lut_2599.LUT_SIZE = 6;
	defparam lut_2599.mask = 64'h5577ffff0008000c;

	lut_sub lut_2602 ({sk[777], i_9_, i_7_, i_8_, i_5_, i_12_, i_0_}, x221x);
	defparam lut_2602.LUT_SIZE = 7;
	defparam lut_2602.mask = 128'h0f0fffffffffffff0000000000000001;

	lut_sub lut_2604 ({sk[778], i_0_, n_n318, n_n316, x741x, x740x, x221x}, x739x);
	defparam lut_2604.LUT_SIZE = 7;
	defparam lut_2604.mask = 128'h0f0fffffffffffff5577557755775f7f;

	lut_sub lut_2608 ({sk[779], i_4_, n_n818, n_n316, n_n752, x304x, x280x}, x214x);
	defparam lut_2608.LUT_SIZE = 7;
	defparam lut_2608.mask = 128'h0f0fffffffffffff0005333700000000;

	lut_sub lut_2611 ({sk[780], i_12_, i_1_, i_2_, i_0_, n_n538, x6573x}, x7211x);
	defparam lut_2611.LUT_SIZE = 7;
	defparam lut_2611.mask = 128'h0f0fffffffffffff0000007000000050;

	lut_sub lut_2614 ({sk[781], i_7_, i_6_, n_n541, x7208x, x236x}, x7212x);
	defparam lut_2614.LUT_SIZE = 6;
	defparam lut_2614.mask = 64'h5577ffff55555557;

	lut_sub lut_2617 ({sk[782], i_12_, i_11_, i_2_, n_n538, x271x, x213x}, x7230x);
	defparam lut_2617.LUT_SIZE = 7;
	defparam lut_2617.mask = 128'h0f0fffffffffffff5555555755555555;

	lut_sub lut_2620 ({sk[783], i_9_, i_7_, i_8_, i_5_, i_12_, i_11_}, x206x);
	defparam lut_2620.LUT_SIZE = 7;
	defparam lut_2620.mask = 128'h0f0fffffffffffff0000000004000000;

	lut_sub lut_2622 ({sk[784], i_5_, i_6_, i_3_, i_1_}, x751x);
	defparam lut_2622.LUT_SIZE = 5;
	defparam lut_2622.mask = 32'h0fff1300;

	lut_sub lut_2625 ({sk[785], i_0_, n_n213, n_n639, x96x, x11x, x332x}, x750x);
	defparam lut_2625.LUT_SIZE = 7;
	defparam lut_2625.mask = 128'h0f0fffffffffffff0000005500003030;

	lut_sub lut_2628 ({sk[786], i_3_, i_0_, x28x, n_n421, n_n358, n_n318}, x7289x);
	defparam lut_2628.LUT_SIZE = 7;
	defparam lut_2628.mask = 128'h0f0fffffffffffff000000000000111f;

	lut_sub lut_2631 ({sk[787], i_10_, i_8_, i_3_, n_n840, x276x, x128x}, x7290x);
	defparam lut_2631.LUT_SIZE = 7;
	defparam lut_2631.mask = 128'h0f0fffffffffffff5555555555575555;

	lut_sub lut_2634 ({sk[788], i_7_, i_12_, i_11_, x8x, n_n639, x7998x}, x7291x);
	defparam lut_2634.LUT_SIZE = 7;
	defparam lut_2634.mask = 128'h0f0fffffffffffff0003aa000000aa00;

	lut_sub lut_2637 ({sk[789], i_5_, x126x, n_n526, n_n844, n_n840, x7306x}, x7308x);
	defparam lut_2637.LUT_SIZE = 7;
	defparam lut_2637.mask = 128'h0f0fffffffffffff55555f7f55555577;

	lut_sub lut_2641 ({sk[790], i_8_, i_5_, n_n453, n_n814, n_n318, x287x}, x7307x);
	defparam lut_2641.LUT_SIZE = 7;
	defparam lut_2641.mask = 128'h0f0fffffffffffff111f000000000000;

	lut_sub lut_2644 ({sk[791], i_10_, i_5_, i_12_, i_11_, i_0_}, x754x);
	defparam lut_2644.LUT_SIZE = 6;
	defparam lut_2644.mask = 64'h5577ffff08000d00;

	lut_sub lut_2647 ({sk[792], i_7_, i_8_, i_3_, i_12_, i_2_}, x753x);
	defparam lut_2647.LUT_SIZE = 6;
	defparam lut_2647.mask = 64'h5577ffff00031113;

	lut_sub lut_2650 ({sk[793], i_5_, i_12_, i_1_, i_11_, i_2_, i_0_}, x752x);
	defparam lut_2650.LUT_SIZE = 7;
	defparam lut_2650.mask = 128'h0f0fffffffffffff0020002000330011;

	lut_sub lut_2655 ({sk[794], i_13_, i_12_, i_1_, i_11_, i_0_}, x862x);
	defparam lut_2655.LUT_SIZE = 6;
	defparam lut_2655.mask = 64'h5577ffff00800000;

	lut_sub lut_2657 ({sk[795], i_10_, i_5_, i_12_, i_11_, i_0_}, x39x);
	defparam lut_2657.LUT_SIZE = 6;
	defparam lut_2657.mask = 64'h5577ffff00201120;

	lut_sub lut_2660 ({sk[796], i_10_, i_7_, i_6_, i_11_}, x393x);
	defparam lut_2660.LUT_SIZE = 5;
	defparam lut_2660.mask = 32'h0fff0008;

	lut_sub lut_2662 ({sk[797], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x525x);
	defparam lut_2662.LUT_SIZE = 7;
	defparam lut_2662.mask = 128'h0f0fffffffffffff0000008000000040;

	lut_sub lut_2665 ({sk[798], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x524x);
	defparam lut_2665.LUT_SIZE = 7;
	defparam lut_2665.mask = 128'h0f0fffffffffffff0000000800000004;

	lut_sub lut_2668 ({sk[799], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x541x);
	defparam lut_2668.LUT_SIZE = 7;
	defparam lut_2668.mask = 128'h0f0fffffffffffff0400000008000000;

	lut_sub lut_2671 ({sk[800], i_9_, i_7_, i_8_, i_6_, i_13_, i_12_}, x569x);
	defparam lut_2671.LUT_SIZE = 7;
	defparam lut_2671.mask = 128'h0f0fffffffffffffc800000000000000;

	lut_sub lut_2674 ({sk[801], i_9_, i_5_, i_3_, i_4_, i_0_}, x613x);
	defparam lut_2674.LUT_SIZE = 6;
	defparam lut_2674.mask = 64'h5577ffff03010000;

	lut_sub lut_2677 ({sk[802], i_7_, i_5_, i_6_, i_1_, i_2_}, x675x);
	defparam lut_2677.LUT_SIZE = 6;
	defparam lut_2677.mask = 64'h5577ffff0000a800;

	lut_sub lut_2680 ({sk[803], i_9_, i_10_, i_7_, i_5_, i_12_, i_11_}, x710x);
	defparam lut_2680.LUT_SIZE = 7;
	defparam lut_2680.mask = 128'h0f0fffffffffffff0000500000035003;

	lut_sub lut_2683 ({sk[804], i_10_, i_12_, i_11_, i_0_}, x719x);
	defparam lut_2683.LUT_SIZE = 5;
	defparam lut_2683.mask = 32'h0fff080d;

	lut_sub lut_2687 ({sk[805], i_10_, i_7_, i_8_, i_5_, i_11_, n_n826}, x128x);
	defparam lut_2687.LUT_SIZE = 7;
	defparam lut_2687.mask = 128'h0f0fffffffffffff0000000010000000;

	lut_sub lut_2689 ({sk[806], i_7_, i_12_, i_2_, x20x, n_n358, n_n197}, x151x);
	defparam lut_2689.LUT_SIZE = 7;
	defparam lut_2689.mask = 128'h0f0fffffffffffff0000000300000007;

	lut_sub lut_2692 ({sk[807], i_9_, i_8_, i_4_, i_2_, i_0_}, x7236x);
	defparam lut_2692.LUT_SIZE = 6;
	defparam lut_2692.mask = 64'h5577ffff20003000;

	lut_sub lut_2695 ({sk[808], i_4_, i_2_, x288x, n_n581, n_n213, x290x}, x199x);
	defparam lut_2695.LUT_SIZE = 7;
	defparam lut_2695.mask = 128'h0f0fffffffffffff0101011100000000;

	lut_sub lut_2698 ({sk[809], x20x, x27x, n_n197, x22x, x206x, x39x}, x201x);
	defparam lut_2698.LUT_SIZE = 7;
	defparam lut_2698.mask = 128'h0f0fffffffffffff030307070303070f;

	lut_sub lut_2702 ({sk[810], i_5_, i_6_, i_3_, i_4_, i_2_, x342x}, x213x);
	defparam lut_2702.LUT_SIZE = 7;
	defparam lut_2702.mask = 128'h0f0fffffffffffff0000000000100000;

	lut_sub lut_2704 ({sk[811], i_10_, i_12_, i_11_, i_0_}, x7208x);
	defparam lut_2704.LUT_SIZE = 5;
	defparam lut_2704.mask = 32'h0fff080c;

	lut_sub lut_2707 ({sk[812], i_9_, i_7_, i_5_, i_6_, n_n318, n_n153}, x236x);
	defparam lut_2707.LUT_SIZE = 7;
	defparam lut_2707.mask = 128'h0f0fffffffffffff0000010000000101;

	lut_sub lut_2710 ({sk[813], i_7_, i_5_, i_3_, i_1_, i_0_, x374x}, x247x);
	defparam lut_2710.LUT_SIZE = 7;
	defparam lut_2710.mask = 128'h0f0fffffffffffff0000000100000000;

	lut_sub lut_2712 ({sk[814], i_9_, i_7_, i_8_, i_6_, i_12_}, x7193x);
	defparam lut_2712.LUT_SIZE = 6;
	defparam lut_2712.mask = 64'h5577ffff00000001;

	lut_sub lut_2714 ({sk[815], i_7_, i_4_, i_0_, x15x, x10x, x710x}, x784x);
	defparam lut_2714.LUT_SIZE = 7;
	defparam lut_2714.mask = 128'h0f0fffffffffffff0005000000070000;

	lut_sub lut_2717 ({sk[816], i_7_, i_5_, i_6_, i_3_, i_0_}, x7172x);
	defparam lut_2717.LUT_SIZE = 6;
	defparam lut_2717.mask = 64'h5577ffff00000004;

	lut_sub lut_2719 ({sk[817], i_7_, i_5_, i_3_, i_0_, x289x, n_n719}, x881x);
	defparam lut_2719.LUT_SIZE = 7;
	defparam lut_2719.mask = 128'h0f0fffffffffffff0000000000000100;

	lut_sub lut_2721 ({sk[818], i_9_, i_8_, i_5_, n_n675, n_n716, x412x}, x883x);
	defparam lut_2721.LUT_SIZE = 7;
	defparam lut_2721.mask = 128'h0f0fffffffffffff0013001100110011;

	lut_sub lut_2724 ({sk[819], i_5_, i_6_, i_4_, n_n675, n_n816, n_n672}, x894x);
	defparam lut_2724.LUT_SIZE = 7;
	defparam lut_2724.mask = 128'h0f0fffffffffffff1113000300000000;

	lut_sub lut_2727 ({sk[820], i_10_, i_8_, i_2_, n_n545, n_n653, x675x}, x896x);
	defparam lut_2727.LUT_SIZE = 7;
	defparam lut_2727.mask = 128'h0f0fffffffffffff0505070500000000;

	lut_sub lut_2730 ({sk[821], i_7_, i_8_, i_5_, n_n816, n_n779, n_n685}, x920x);
	defparam lut_2730.LUT_SIZE = 7;
	defparam lut_2730.mask = 128'h0f0fffffffffffff0700050003000000;

	lut_sub lut_2733 ({sk[822], i_5_, i_3_, i_0_}, x7083x);
	defparam lut_2733.LUT_SIZE = 4;
	defparam lut_2733.mask = 16'h0f40;

	lut_sub lut_2735 ({sk[823], i_8_, i_11_, i_0_, n_n575, n_n606, x413x}, x949x);
	defparam lut_2735.LUT_SIZE = 7;
	defparam lut_2735.mask = 128'h0f0fffffffffffff0003000005070505;

	lut_sub lut_2738 ({sk[824], i_5_, i_3_, i_11_, i_2_, n_n773}, x984x);
	defparam lut_2738.LUT_SIZE = 6;
	defparam lut_2738.mask = 64'h5577ffff40000000;

	lut_sub lut_2740 ({sk[825], i_9_, i_10_, i_3_, i_2_, n_n526, x11x}, x986x);
	defparam lut_2740.LUT_SIZE = 7;
	defparam lut_2740.mask = 128'h0f0fffffffffffff3330000010100000;

	lut_sub lut_2744 ({sk[826], i_10_, i_7_, i_8_, i_12_, i_11_, n_n653}, x987x);
	defparam lut_2744.LUT_SIZE = 7;
	defparam lut_2744.mask = 128'h0f0fffffffffffff4440000000000000;

	lut_sub lut_2747 ({sk[827], i_6_, i_2_, i_0_, n_n242, n_n277}, x1075x);
	defparam lut_2747.LUT_SIZE = 6;
	defparam lut_2747.mask = 64'h5577ffff30005000;

	lut_sub lut_2750 ({sk[828], i_7_, i_8_, i_3_, i_2_, x37x, n_n716}, x1095x);
	defparam lut_2750.LUT_SIZE = 7;
	defparam lut_2750.mask = 128'h0f0fffffffffffff0000000070300000;

	lut_sub lut_2753 ({sk[829], i_3_, i_13_, i_12_, i_11_, n_n275, x351x}, x1141x);
	defparam lut_2753.LUT_SIZE = 7;
	defparam lut_2753.mask = 128'h0f0fffffffffffff0075000000000000;

	lut_sub lut_2756 ({sk[830], i_7_, i_8_, i_3_, x294x, x273x}, x1142x);
	defparam lut_2756.LUT_SIZE = 6;
	defparam lut_2756.mask = 64'h5577ffff55750000;

	lut_sub lut_2759 ({sk[831], i_8_, i_3_, n_n741, x32x, x105x, x275x}, x1185x);
	defparam lut_2759.LUT_SIZE = 7;
	defparam lut_2759.mask = 128'h0f0fffffffffffff030f030703070307;

	lut_sub lut_2763 ({sk[832], i_6_, i_3_, i_4_, i_1_, i_11_, i_2_}, x1204x);
	defparam lut_2763.LUT_SIZE = 7;
	defparam lut_2763.mask = 128'h0f0fffffffffffff0000400000000000;

	lut_sub lut_2765 ({sk[833], i_9_, i_7_, i_6_, i_12_, i_1_, i_11_}, x1211x);
	defparam lut_2765.LUT_SIZE = 7;
	defparam lut_2765.mask = 128'h0f0fffffffffffff0040000000500000;

	lut_sub lut_2768 ({sk[834], i_4_, i_1_, n_n316, n_n35, n_n756, x393x}, x1220x);
	defparam lut_2768.LUT_SIZE = 7;
	defparam lut_2768.mask = 128'h0f0fffffffffffff0537050500000000;

	lut_sub lut_2771 ({sk[835], i_7_, i_6_, i_3_, i_12_}, x6913x);
	defparam lut_2771.LUT_SIZE = 5;
	defparam lut_2771.mask = 32'h0fff0010;

	lut_sub lut_2773 ({sk[836], i_9_, i_10_, i_6_, i_12_, i_11_, i_2_}, x1234x);
	defparam lut_2773.LUT_SIZE = 7;
	defparam lut_2773.mask = 128'h0f0fffffffffffff0000000000004450;

	lut_sub lut_2777 ({sk[837], i_10_, i_8_, i_6_, i_12_, i_11_, n_n534}, x1256x);
	defparam lut_2777.LUT_SIZE = 7;
	defparam lut_2777.mask = 128'h0f0fffffffffffff0000000040500000;

	lut_sub lut_2780 ({sk[838], i_9_, i_10_, i_7_, i_8_, i_6_, i_12_}, x1288x);
	defparam lut_2780.LUT_SIZE = 7;
	defparam lut_2780.mask = 128'h0f0fffffffffffff0000000000000004;

	lut_sub lut_2782 ({sk[839], i_10_, i_3_, i_13_, i_12_, i_11_}, x6862x);
	defparam lut_2782.LUT_SIZE = 6;
	defparam lut_2782.mask = 64'h5577ffff40000000;

	lut_sub lut_2784 ({sk[840], i_7_, i_8_, i_6_, n_n779, n_n849, n_n685}, x1364x);
	defparam lut_2784.LUT_SIZE = 7;
	defparam lut_2784.mask = 128'h0f0fffffffffffff0013001100030000;

	lut_sub lut_2787 ({sk[841], i_6_, i_4_, i_1_, n_n675, n_n792, n_n761}, x1365x);
	defparam lut_2787.LUT_SIZE = 7;
	defparam lut_2787.mask = 128'h0f0fffffffffffff0000000000001505;

	lut_sub lut_2790 ({sk[842], i_7_, i_5_, i_6_, i_3_, n_n814, n_n826}, x7994x);
	defparam lut_2790.LUT_SIZE = 7;
	defparam lut_2790.mask = 128'h0f0fffffffffffff8088aaaaccccffff;

	lut_sub lut_2796 ({sk[843], i_9_, i_10_, i_7_, i_6_, i_11_}, x6810x);
	defparam lut_2796.LUT_SIZE = 6;
	defparam lut_2796.mask = 64'h5577ffff00000004;

	lut_sub lut_2798 ({sk[844], i_10_, i_7_, i_8_, i_5_, i_6_, i_11_}, x6795x);
	defparam lut_2798.LUT_SIZE = 7;
	defparam lut_2798.mask = 128'h0f0fffffffffffff0000000080000000;

	lut_sub lut_2800 ({sk[845], i_13_, i_4_, i_1_, i_0_}, x6785x);
	defparam lut_2800.LUT_SIZE = 5;
	defparam lut_2800.mask = 32'h0fff0400;

	lut_sub lut_2802 ({sk[846], i_5_, i_6_, i_1_, i_2_, n_n822, x24x}, x7992x);
	defparam lut_2802.LUT_SIZE = 7;
	defparam lut_2802.mask = 128'h0f0ffffffffffffffffffffffefefffe;

	lut_sub lut_2816 ({sk[847], i_8_, n_n598, x273x, x385x, x42x, x7992x}, x1425x);
	defparam lut_2816.LUT_SIZE = 7;
	defparam lut_2816.mask = 128'h0f0fffffffffffffaabfaaff00000000;

	lut_sub lut_2821 ({sk[848], i_7_, i_1_}, x6775x);
	defparam lut_2821.LUT_SIZE = 3;
	defparam lut_2821.mask = 8'h34;

	lut_sub lut_2823 ({sk[849], i_7_, i_6_, n_n816, n_n822, x6774x, x613x}, x1438x);
	defparam lut_2823.LUT_SIZE = 7;
	defparam lut_2823.mask = 128'h0f0fffffffffffff0357000000000000;

	lut_sub lut_2826 ({sk[850], i_9_, i_6_, i_4_, n_n818, n_n849, x1448x}, x1439x);
	defparam lut_2826.LUT_SIZE = 7;
	defparam lut_2826.mask = 128'h0f0fffffffffffff1111111311111111;

	lut_sub lut_2829 ({sk[851], i_7_, i_6_, i_3_}, x6762x);
	defparam lut_2829.LUT_SIZE = 4;
	defparam lut_2829.mask = 16'h0f01;

	lut_sub lut_2831 ({sk[852], i_9_, i_5_, i_4_, i_2_, x15x, x287x}, x7983x);
	defparam lut_2831.LUT_SIZE = 7;
	defparam lut_2831.mask = 128'h0f0fffffffffffffffaaffa8ffffffff;

	lut_sub lut_2837 ({sk[853], i_10_, i_13_, i_12_, n_n819, n_n846, x7983x}, x1466x);
	defparam lut_2837.LUT_SIZE = 7;
	defparam lut_2837.mask = 128'h0f0fffffffffffff00ab000000000000;

	lut_sub lut_2840 ({sk[854], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x6753x);
	defparam lut_2840.LUT_SIZE = 7;
	defparam lut_2840.mask = 128'h0f0fffffffffffff0010000000000000;

	lut_sub lut_2842 ({sk[855], i_9_, i_7_, i_8_, i_1_, i_0_}, x6743x);
	defparam lut_2842.LUT_SIZE = 6;
	defparam lut_2842.mask = 64'h5577ffff00010000;

	lut_sub lut_2844 ({sk[856], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x6709x);
	defparam lut_2844.LUT_SIZE = 7;
	defparam lut_2844.mask = 128'h0f0fffffffffffff0000000000001000;

	lut_sub lut_2846 ({sk[857], i_10_, i_7_, i_8_, i_6_, i_11_}, x6710x);
	defparam lut_2846.LUT_SIZE = 6;
	defparam lut_2846.mask = 64'h5577ffff00001000;

	lut_sub lut_2848 ({sk[858], i_9_, i_10_, i_7_, i_6_, i_3_, i_0_}, x1540x);
	defparam lut_2848.LUT_SIZE = 7;
	defparam lut_2848.mask = 128'h0f0fffffffffffff0000000000000001;

	lut_sub lut_2850 ({sk[859], i_9_, i_10_, i_7_, i_5_, i_3_, i_1_}, x1541x);
	defparam lut_2850.LUT_SIZE = 7;
	defparam lut_2850.mask = 128'h0f0fffffffffffff0000000000000001;

	lut_sub lut_2852 ({sk[860], i_7_, i_8_, i_6_, i_3_, x35x, x6664x}, x1596x);
	defparam lut_2852.LUT_SIZE = 7;
	defparam lut_2852.mask = 128'h0f0fffffffffffff1000000000000000;

	lut_sub lut_2854 ({sk[861], i_5_, i_3_, i_4_, i_1_, i_2_, i_0_}, x6655x);
	defparam lut_2854.LUT_SIZE = 7;
	defparam lut_2854.mask = 128'h0f0fffffffffffff4000000000000000;

	lut_sub lut_2856 ({sk[862], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x6609x);
	defparam lut_2856.LUT_SIZE = 7;
	defparam lut_2856.mask = 128'h0f0fffffffffffff0000000000000001;

	lut_sub lut_2858 ({sk[863], i_8_, i_6_, i_3_, i_4_, i_2_, i_0_}, x6596x);
	defparam lut_2858.LUT_SIZE = 7;
	defparam lut_2858.mask = 128'h0f0fffffffffffff0000000010000000;

	lut_sub lut_2860 ({sk[864], i_9_, i_5_, i_3_, i_4_, i_11_}, x6568x);
	defparam lut_2860.LUT_SIZE = 6;
	defparam lut_2860.mask = 64'h5577ffff00000800;

	lut_sub lut_2862 ({sk[865], i_7_, i_8_, i_6_, i_1_, i_2_, i_0_}, x6540x);
	defparam lut_2862.LUT_SIZE = 7;
	defparam lut_2862.mask = 128'h0f0fffffffffffff0000004000000000;

	lut_sub lut_2864 ({sk[866], i_7_, i_8_, i_5_, i_6_, i_3_, i_4_}, x6542x);
	defparam lut_2864.LUT_SIZE = 7;
	defparam lut_2864.mask = 128'h0f0fffffffffffff0002000000000000;

	lut_sub lut_2866 ({sk[867], i_8_, i_1_, i_2_, i_0_, n_n538, x28x}, x7991x);
	defparam lut_2866.LUT_SIZE = 7;
	defparam lut_2866.mask = 128'h0f0fffffffffffffffffffffffffefff;

	lut_sub lut_2882 ({sk[868], i_9_, i_10_, i_8_, i_3_, i_13_, i_11_}, x6484x);
	defparam lut_2882.LUT_SIZE = 7;
	defparam lut_2882.mask = 128'h0f0fffffffffffff2000200020002303;

	lut_sub lut_2885 ({sk[869], i_9_, i_7_, i_8_, i_5_, i_6_, x277x}, x7988x);
	defparam lut_2885.LUT_SIZE = 7;
	defparam lut_2885.mask = 128'h0f0fffffffffffffbbffffffbfffffff;

	lut_sub lut_2891 ({sk[870], n_n849, n_n850, n_n748, n_n755, x544x, x543x}, x6665x);
	defparam lut_2891.LUT_SIZE = 7;
	defparam lut_2891.mask = 128'h0f0fffffffffffff0000030300550357;

	lut_sub lut_2894 ({sk[871], i_1_, n_n816, n_n795, x17x, x35x, x6718x}, x6726x);
	defparam lut_2894.LUT_SIZE = 7;
	defparam lut_2894.mask = 128'h0f0fffffffffffff0505050505050537;

	lut_sub lut_2897 ({sk[872], i_10_, i_8_, i_5_, n_n853, n_n779, x394x}, x6727x);
	defparam lut_2897.LUT_SIZE = 7;
	defparam lut_2897.mask = 128'h0f0fffffffffffff0705050505050505;

	lut_sub lut_2900 ({sk[873], i_6_, i_1_, i_2_, i_0_, n_n822, x24x}, x7993x);
	defparam lut_2900.LUT_SIZE = 7;
	defparam lut_2900.mask = 128'h0f0ffffffffffffffefffefffeffffff;

	lut_sub lut_2914 ({sk[874], i_8_, i_5_, i_2_, x17x, n_n773, x7993x}, x6728x);
	defparam lut_2914.LUT_SIZE = 7;
	defparam lut_2914.mask = 128'h0f0fffffffffffffabaaaaaa03000000;

	lut_sub lut_2917 ({sk[875], i_8_, i_1_, i_2_, n_n2368, x37x, x322x}, x6729x);
	defparam lut_2917.LUT_SIZE = 7;
	defparam lut_2917.mask = 128'h0f0fffffffffffff001100110011001f;

	lut_sub lut_2920 ({sk[876], i_9_, i_13_, n_n844, n_n752, n_n846}, x7984x);
	defparam lut_2920.LUT_SIZE = 6;
	defparam lut_2920.mask = 64'h5577fffffeffffff;

	lut_sub lut_2932 ({sk[877], i_2_, n_n2368, n_n822, x24x, n_n639, x6762x}, x6765x);
	defparam lut_2932.LUT_SIZE = 7;
	defparam lut_2932.mask = 128'h0f0fffffffffffff0000555500035557;

	lut_sub lut_2935 ({sk[878], i_5_, i_2_, x15x, x273x, x292x, x340x}, x6778x);
	defparam lut_2935.LUT_SIZE = 7;
	defparam lut_2935.mask = 128'h0f0fffffffffffff1111111f11111111;

	lut_sub lut_2938 ({sk[879], i_6_, n_n2368, n_n822, x96x, x6774x, x6775x}, x6779x);
	defparam lut_2938.LUT_SIZE = 7;
	defparam lut_2938.mask = 128'h0f0fffffffffffff001100110011f0f1;

	lut_sub lut_2941 ({sk[880], i_7_, n_n816, n_n795, n_n822, x574x, x6785x}, x6789x);
	defparam lut_2941.LUT_SIZE = 7;
	defparam lut_2941.mask = 128'h0f0fffffffffffff0005333700050005;

	lut_sub lut_2944 ({sk[881], i_9_, i_7_, i_6_, n_n761, n_n538, n_n453}, x7996x);
	defparam lut_2944.LUT_SIZE = 7;
	defparam lut_2944.mask = 128'h0f0ffffffffffffffffffffffffeffff;

	lut_sub lut_2959 ({sk[882], i_1_, i_2_, i_0_, x6807x, x7996x}, x6813x);
	defparam lut_2959.LUT_SIZE = 6;
	defparam lut_2959.mask = 64'h5577ffffa0000003;

	lut_sub lut_2962 ({sk[883], i_0_, x265x, x272x, x46x, x302x, x6810x}, x6814x);
	defparam lut_2962.LUT_SIZE = 7;
	defparam lut_2962.mask = 128'h0f0fffffffffffff000f111f000f000f;

	lut_sub lut_2965 ({sk[884], n_n675, x326x, n_n716, n_n545, x29x, x289x}, x6839x);
	defparam lut_2965.LUT_SIZE = 7;
	defparam lut_2965.mask = 128'h0f0fffffffffffff0000030300550357;

	lut_sub lut_2968 ({sk[885], i_7_, i_8_, i_6_, n_n761, x346x, x6862x}, x6866x);
	defparam lut_2968.LUT_SIZE = 7;
	defparam lut_2968.mask = 128'h0f0fffffffffffff0003550300030003;

	lut_sub lut_2971 ({sk[886], i_10_, i_7_, i_6_, i_1_, i_11_, i_2_}, x6888x);
	defparam lut_2971.LUT_SIZE = 7;
	defparam lut_2971.mask = 128'h0f0fffffffffffff0000000045000000;

	lut_sub lut_2974 ({sk[887], i_10_, i_7_, i_6_, i_1_, i_11_, x332x}, x7976x);
	defparam lut_2974.LUT_SIZE = 7;
	defparam lut_2974.mask = 128'h0f0fffffffffffffffffffffbfafffff;

	lut_sub lut_2988 ({sk[888], i_6_, i_4_, i_1_, i_2_, x270x, x552x}, x6926x);
	defparam lut_2988.LUT_SIZE = 7;
	defparam lut_2988.mask = 128'h0f0fffffffffffff0055000000570000;

	lut_sub lut_2991 ({sk[889], i_10_, i_12_, i_1_, i_11_, x268x, x1211x}, x7975x);
	defparam lut_2991.LUT_SIZE = 7;
	defparam lut_2991.mask = 128'h0f0fffffffffffffaaaa8aaaaaaa8a8a;

	lut_sub lut_2996 ({sk[890], i_5_, i_6_, i_2_, n_n242, n_n277}, x7047x);
	defparam lut_2996.LUT_SIZE = 6;
	defparam lut_2996.mask = 64'h5577ffff30000050;

	lut_sub lut_2999 ({sk[891], i_5_, i_12_, i_11_, i_0_, x986x}, x7060x);
	defparam lut_2999.LUT_SIZE = 6;
	defparam lut_2999.mask = 64'h5577ffffd5d5d555;

	lut_sub lut_3003 ({sk[892], i_9_, i_7_, n_n658, n_n526, x984x, x987x}, x7061x);
	defparam lut_3003.LUT_SIZE = 7;
	defparam lut_3003.mask = 128'h0f0fffffffffffff7777777f77777777;

	lut_sub lut_3007 ({sk[893], i_9_, i_10_, i_12_, i_11_, x323x, x325x}, x7071x);
	defparam lut_3007.LUT_SIZE = 7;
	defparam lut_3007.mask = 128'h0f0fffffffffffff7500000030000000;

	lut_sub lut_3010 ({sk[894], i_8_, n_n843, n_n729, x413x, x952x, x7083x}, x7088x);
	defparam lut_3010.LUT_SIZE = 7;
	defparam lut_3010.mask = 128'h0f0fffffffffffff111f115f11111155;

	lut_sub lut_3014 ({sk[895], n_n545, x370x, x6733x, n_n653, n_n240, x324x}, x7106x);
	defparam lut_3014.LUT_SIZE = 7;
	defparam lut_3014.mask = 128'h0f0fffffffffffff000000ff131313ff;

	lut_sub lut_3018 ({sk[896], i_5_, i_6_, i_1_, i_0_, n_n550, x881x}, x7124x);
	defparam lut_3018.LUT_SIZE = 7;
	defparam lut_3018.mask = 128'h0f0fffffffffffff5555555555555755;

	lut_sub lut_3021 ({sk[897], n_n819, n_n671, n_n176, x301x, x284x, x280x}, x7148x);
	defparam lut_3021.LUT_SIZE = 7;
	defparam lut_3021.mask = 128'h0f0fffffffffffff0000003305050537;

	lut_sub lut_3024 ({sk[898], i_7_, i_5_, i_0_, x265x, n_n545, x7148x}, x7149x);
	defparam lut_3024.LUT_SIZE = 7;
	defparam lut_3024.mask = 128'h0f0fffffffffffff5555555557555555;

	lut_sub lut_3027 ({sk[899], i_7_, n_n213, n_n153, x11x, x397x, x247x}, x7204x);
	defparam lut_3027.LUT_SIZE = 7;
	defparam lut_3027.mask = 128'h0f0fffffffffffff5577557f55555555;

	lut_sub lut_3031 ({sk[900], n_n311, x13x, n_n598, x357x, x374x, x7236x}, x7240x);
	defparam lut_3031.LUT_SIZE = 7;
	defparam lut_3031.mask = 128'h0f0fffffffffffff0003000300035557;

	lut_sub lut_3034 ({sk[901], i_7_, i_12_, i_11_, x708x, x357x, x729x}, x7968x);
	defparam lut_3034.LUT_SIZE = 7;
	defparam lut_3034.mask = 128'h0f0fffffffffffffeee0eeeeeeeeeeee;

	lut_sub lut_3043 ({sk[902], i_12_, x16x, x30x, n_n213, n_n598, x352x}, x7251x);
	defparam lut_3043.LUT_SIZE = 7;
	defparam lut_3043.mask = 128'h0f0fffffffffffff0003000300030507;

	lut_sub lut_3046 ({sk[903], i_9_, i_8_, i_2_, n_n311, n_n639, x151x}, x7270x);
	defparam lut_3046.LUT_SIZE = 7;
	defparam lut_3046.mask = 128'h0f0fffffffffffff5555555555555557;

	lut_sub lut_3049 ({sk[904], i_8_, i_5_, x8x, n_n818, x292x, x397x}, x7271x);
	defparam lut_3049.LUT_SIZE = 7;
	defparam lut_3049.mask = 128'h0f0fffffffffffff0000000005370505;

	lut_sub lut_3052 ({sk[905], i_7_, i_5_, i_6_, i_3_, i_1_, n_n311}, x7999x);
	defparam lut_3052.LUT_SIZE = 7;
	defparam lut_3052.mask = 128'h0f0ffffffffffffffffffafeffffffff;

	lut_sub lut_3066 ({sk[906], i_10_, i_8_, i_3_, i_2_, x26x, x314x}, x7998x);
	defparam lut_3066.LUT_SIZE = 7;
	defparam lut_3066.mask = 128'h0f0fffffffffffffffeeffeeffecffee;

	lut_sub lut_3080 ({sk[907], i_3_, n_n316, n_n837, n_n597, x338x, x751x}, x7306x);
	defparam lut_3080.LUT_SIZE = 7;
	defparam lut_3080.mask = 128'h0f0fffffffffffff0000050500330537;

	lut_sub lut_3083 ({sk[908], i_2_, i_0_, n_n421, n_n358, x754x, x753x}, x7316x);
	defparam lut_3083.LUT_SIZE = 7;
	defparam lut_3083.mask = 128'h0f0fffffffffffff0000005503030357;

	lut_sub lut_3086 ({sk[909], i_5_, i_6_, i_1_, i_0_, n_n2368, n_n729}, x7329x);
	defparam lut_3086.LUT_SIZE = 7;
	defparam lut_3086.mask = 128'h0f0fffffffffffff3733333333333333;

	lut_sub lut_3089 ({sk[910], x7082x, x947x, n_n838, x528x, x949x, x7088x}, x7332x);
	defparam lut_3089.LUT_SIZE = 7;
	defparam lut_3089.mask = 128'h0f0fffffffffffff777fffffffffffff;

	lut_sub lut_3095 ({sk[911], x7101x, x7102x, x884x, x883x, x7124x}, x7333x);
	defparam lut_3095.LUT_SIZE = 6;
	defparam lut_3095.mask = 64'h5577ffff7fffffff;


endmodule