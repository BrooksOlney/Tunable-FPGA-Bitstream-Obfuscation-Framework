module spla_qmap_map (sk, i_0_, i_1_, i_8_, i_6_, i_7_, i_9_, i_10_, i_11_, i_15_, i_12_, i_13_, i_14_, i_4_, i_3_, i_5_, i_2_, o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_, o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_, o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_, o_41_, o_42_, o_43_, o_44_, o_45_);

	input i_0_;
	input i_1_;
	input i_8_;
	input i_6_;
	input i_7_;
	input i_9_;
	input i_10_;
	input i_11_;
	input i_15_;
	input i_12_;
	input i_13_;
	input i_14_;
	input i_4_;
	input i_3_;
	input i_5_;
	input i_2_;
	output o_0_;
	output o_1_;
	output o_2_;
	output o_3_;
	output o_4_;
	output o_5_;
	output o_6_;
	output o_7_;
	output o_8_;
	output o_9_;
	output o_10_;
	output o_11_;
	output o_12_;
	output o_13_;
	output o_14_;
	output o_15_;
	output o_16_;
	output o_17_;
	output o_18_;
	output o_19_;
	output o_20_;
	output o_21_;
	output o_22_;
	output o_23_;
	output o_24_;
	output o_25_;
	output o_26_;
	output o_27_;
	output o_28_;
	output o_29_;
	output o_30_;
	output o_31_;
	output o_32_;
	output o_33_;
	output o_34_;
	output o_35_;
	output o_36_;
	output o_37_;
	output o_38_;
	output o_39_;
	output o_40_;
	output o_41_;
	output o_42_;
	output o_43_;
	output o_44_;
	output o_45_;



	wire g9, g11, g52, g456, g458, g621, g812, g845, g846, g923, g963, g989, g1003, g1456, g1018, g1057, g1454, g1077, g1125, g1128, g1129;
	wire g1253, g1346, g1393, g1417, g1422, g1424, g1426, g1437, g1449, g1451, g1, g2, g3, g4, g5, g6, g7, g8, g10, g12, g14;
	wire g15, g16, g17, g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29, g30, g31, g32, g33, g34, g35;
	wire g36, g37, g38, g39, g40, g41, g42, g43, g44, g45, g46, g47, g48, g49, g50, g51, g53, g54, g55, g56, g57;
	wire g58, g59, g60, g61, g62, g63, g64, g65, g66, g68, g69, g70, g71, g72, g73, g74, g75, g76, g77, g78, g79;
	wire g80, g81, g82, g83, g84, g85, g86, g87, g88, g89, g90, g91, g92, g93, g94, g95, g96, g97, g98, g99, g100;
	wire g101, g102, g103, g104, g105, g106, g107, g108, g109, g110, g111, g112, g113, g114, g115, g116, g117, g118, g119, g120, g121;
	wire g122, g123, g124, g125, g126, g127, g128, g129, g130, g131, g1639, g132, g133, g134, g135, g136, g137, g138, g139, g140, g141;
	wire g142, g143, g144, g145, g146, g147, g148, g149, g150, g151, g152, g153, g154, g155, g156, g157, g158, g159, g160, g161, g162;
	wire g163, g164, g165, g166, g167, g168, g169, g170, g171, g172, g173, g174, g175, g176, g177, g178, g179, g180, g181, g182, g183;
	wire g184, g185, g186, g187, g188, g189, g190, g191, g192, g193, g194, g195, g196, g197, g198, g199, g200, g201, g202, g203, g204;
	wire g205, g206, g207, g208, g209, g210, g211, g212, g213, g214, g215, g216, g217, g218, g219, g220, g221, g222, g223, g224, g225;
	wire g226, g227, g228, g229, g230, g231, g232, g233, g234, g235, g236, g237, g238, g239, g240, g241, g242, g243, g244, g245, g246;
	wire g247, g248, g249, g250, g251, g252, g253, g254, g255, g256, g257, g258, g259, g260, g261, g262, g263, g264, g265, g266, g267;
	wire g268, g269, g270, g271, g272, g273, g274, g275, g276, g277, g278, g279, g280, g281, g282, g283, g284, g285, g286, g287, g288;
	wire g289, g290, g291, g292, g293, g294, g295, g296, g297, g298, g299, g300, g301, g302, g303, g304, g305, g306, g307, g308, g309;
	wire g310, g311, g312, g313, g314, g315, g1632, g316, g317, g318, g319, g320, g1625, g321, g322, g323, g324, g325, g326, g327, g328;
	wire g329, g330, g1606, g331, g1613, g332, g333, g334, g335, g336, g337, g338, g339, g340, g341, g342, g343, g344, g345, g346, g347;
	wire g348, g349, g350, g351, g352, g353, g354, g355, g356, g357, g358, g359, g360, g361, g362, g363, g364, g365, g366, g367, g368;
	wire g369, g370, g371, g372, g373, g374, g375, g376, g377, g378, g379, g380, g381, g382, g383, g384, g385, g386, g387, g388, g389;
	wire g390, g391, g392, g393, g394, g395, g396, g397, g398, g399, g400, g401, g402, g403, g404, g405, g406, g407, g408, g409, g410;
	wire g411, g412, g413, g414, g415, g416, g417, g418, g419, g420, g421, g422, g423, g424, g425, g426, g427, g428, g429, g430, g431;
	wire g432, g433, g434, g435, g436, g437, g438, g439, g440, g441, g1593, g442, g443, g444, g445, g446, g447, g448, g449, g450, g451;
	wire g452, g453, g454, g1584, g455, g457, g459, g460, g461, g462, g463, g464, g465, g466, g467, g468, g469, g470, g471, g472, g473;
	wire g474, g475, g476, g477, g478, g479, g480, g481, g482, g483, g484, g485, g486, g487, g488, g489, g490, g491, g492, g493, g494;
	wire g495, g496, g497, g498, g499, g500, g501, g502, g503, g504, g505, g506, g507, g508, g509, g510, g511, g512, g513, g514, g515;
	wire g516, g517, g518, g1577, g519, g520, g521, g522, g523, g524, g1564, g525, g526, g527, g528, g529, g530, g531, g532, g533, g534;
	wire g535, g536, g1459, g537, g538, g539, g540, g541, g542, g543, g544, g545, g546, g547, g548, g549, g550, g551, g552, g553, g554;
	wire g555, g556, g557, g558, g559, g560, g561, g562, g563, g564, g565, g566, g567, g568, g569, g570, g571, g572, g573, g574, g575;
	wire g576, g577, g578, g579, g580, g1554, g1543, g581, g582, g583, g584, g585, g586, g587, g588, g589, g590, g591, g592, g593, g594;
	wire g595, g596, g597, g598, g599, g600, g601, g602, g603, g604, g605, g606, g607, g608, g609, g610, g611, g612, g613, g614, g615;
	wire g616, g617, g618, g1458, g619, g620, g623, g624, g625, g626, g627, g628, g629, g630, g631, g632, g633, g634, g635, g636, g637;
	wire g638, g639, g640, g641, g642, g643, g644, g645, g646, g647, g648, g649, g650, g651, g652, g653, g654, g655, g656, g657, g658;
	wire g659, g660, g661, g662, g663, g664, g665, g666, g667, g668, g669, g670, g671, g672, g673, g674, g675, g676, g677, g678, g679;
	wire g680, g681, g682, g683, g684, g685, g686, g687, g688, g689, g690, g1457, g691, g692, g693, g694, g695, g696, g697, g698, g699;
	wire g700, g701, g702, g703, g704, g705, g706, g1531, g707, g708, g709, g710, g711, g712, g713, g714, g715, g716, g717, g718, g719;
	wire g720, g721, g722, g723, g724, g725, g726, g727, g728, g729, g730, g731, g732, g733, g734, g735, g736, g737, g738, g739, g740;
	wire g741, g742, g743, g744, g745, g746, g747, g1518, g748, g749, g750, g751, g752, g753, g754, g755, g756, g757, g758, g759, g760;
	wire g761, g762, g763, g764, g765, g766, g767, g768, g769, g770, g771, g772, g773, g774, g775, g776, g777, g778, g779, g780, g781;
	wire g782, g783, g784, g785, g786, g787, g788, g789, g790, g791, g792, g793, g794, g795, g796, g797, g798, g799, g800, g801, g802;
	wire g803, g804, g805, g806, g807, g808, g809, g810, g811, g813, g814, g815, g816, g817, g818, g819, g820, g821, g822, g823, g824;
	wire g825, g826, g827, g828, g829, g830, g831, g832, g833, g834, g835, g836, g837, g838, g839, g840, g841, g842, g843, g1511, g844;
	wire g847, g848, g849, g850, g851, g852, g853, g854, g855, g856, g857, g858, g859, g860, g861, g862, g863, g864, g865, g866, g867;
	wire g868, g869, g870, g871, g872, g1501, g1488, g873, g874, g875, g876, g877, g878, g879, g880, g881, g882, g883, g884, g885, g886;
	wire g887, g888, g889, g890, g891, g892, g893, g894, g895, g896, g1478, g897, g898, g899, g900, g901, g902, g903, g904, g905, g906;
	wire g907, g908, g909, g910, g911, g912, g913, g914, g915, g916, g917, g918, g919, g920, g921, g922, g924, g925, g926, g927, g928;
	wire g929, g930, g931, g932, g933, g934, g935, g936, g937, g938, g939, g940, g941, g942, g943, g944, g945, g946, g947, g948, g949;
	wire g950, g1467, g951, g952, g953, g954, g955, g956, g957, g958, g959, g960, g961, g962, g964, g965, g966, g967, g968, g969, g970;
	wire g971, g972, g973, g974, g975, g976, g977, g978, g979, g980, g981, g982, g983, g984, g985, g986, g987, g988, g990, g991, g992;
	wire g993, g994, g995, g996, g997, g998, g999, g1000, g1001, g1002, g1004, g1005, g1006, g1007, g1008, g1009, g1010, g1011, g1012, g1013, g1455;
	wire g1014, g1015, g1016, g1017, g1019, g1020, g1021, g1022, g1023, g1024, g1025, g1026, g1027, g1028, g1029, g1030, g1031, g1032, g1033, g1034, g1035;
	wire g1036, g1037, g1038, g1039, g1040, g1041, g1042, g1043, g1044, g1045, g1046, g1047, g1048, g1049, g1050, g1051, g1052, g1053, g1054, g1055, g1056;
	wire g1058, g1060, g1062, g1063, g1064, g1065, g1067, g1068, g1069, g1070, g1071, g1072, g1073, g1074, g1075, g1076, g1080, g1081, g1082, g1084, g1085;
	wire g1086, g1087, g1088, g1090, g1091, g1094, g1095, g1096, g1097, g1098, g1099, g1100, g1101, g1102, g1103, g1104, g1105, g1106, g1107, g1108, g1109;
	wire g1110, g1111, g1112, g1460, g1113, g1114, g1115, g1116, g1117, g1118, g1119, g1122, g1123, g1124, g1126, g1127, g1130, g1131, g1132, g1133, g1134;
	wire g1135, g1136, g1137, g1138, g1139, g1140, g1141, g1142, g1143, g1144, g1145, g1146, g1147, g1148, g1149, g1150, g1151, g1152, g1153, g1154, g1155;
	wire g1156, g1157, g1158, g1159, g1160, g1161, g1162, g1163, g1164, g1165, g1166, g1167, g1168, g1169, g1170, g1171, g1172, g1173, g1174, g1175, g1176;
	wire g1177, g1178, g1179, g1180, g1181, g1182, g1453, g1183, g1184, g1185, g1186, g1452, g1187, g1188, g1189, g1190, g1191, g1192, g1193, g1194, g1195;
	wire g1196, g1197, g1198, g1199, g1200, g1201, g1202, g1203, g1204, g1205, g1206, g1207, g1208, g1209, g1210, g1211, g1212, g1213, g1214, g1215, g1216;
	wire g1217, g1218, g1219, g1220, g1221, g1222, g1223, g1224, g1225, g1226, g1227, g1228, g1229, g1230, g1231, g1232, g1233, g1234, g1235, g1236, g1237;
	wire g1238, g1239, g1240, g1241, g1242, g1243, g1244, g1245, g1246, g1247, g1248, g1249, g1250, g1251, g1252, g1254, g1255, g1256, g1257, g1258, g1259;
	wire g1260, g1261, g1262, g1263, g1264, g1265, g1266, g1267, g1268, g1269, g1270, g1271, g1272, g1273, g1274, g1275, g1276, g1277, g1278, g1279, g1280;
	wire g1281, g1282, g1283, g1284, g1285, g1286, g1287, g1288, g1289, g1290, g1291, g1292, g1293, g1294, g1295, g1296, g1297, g1298, g1299, g1300, g1301;
	wire g1302, g1303, g1304, g1305, g1306, g1307, g1308, g1309, g1310, g1311, g1312, g1313, g1314, g1315, g1316, g1317, g1318, g1319, g1320, g1321, g1322;
	wire g1323, g1324, g1325, g1326, g1327, g1328, g1329, g1330, g1331, g1332, g1333, g1334, g1335, g1336, g1337, g1338, g1339, g1340, g1341, g1342, g1343;
	wire g1344, g1345, g1347, g1348, g1349, g1350, g1351, g1352, g1353, g1354, g1355, g1356, g1357, g1358, g1359, g1360, g1361, g1362, g1363, g1364, g1365;
	wire g1366, g1367, g1368, g1369, g1370, g1371, g1372, g1373, g1374, g1375, g1376, g1377, g1378, g1379, g1380, g1381, g1382, g1383, g1384, g1385, g1386;
	wire g1387, g1388, g1389, g1390, g1391, g1392, g1394, g1395, g1396, g1397, g1398, g1399, g1400, g1401, g1402, g1403, g1404, g1405, g1406, g1407, g1408;
	wire g1409, g1410, g1411, g1412, g1413, g1414, g1415, g1416, g1418, g1419, g1420, g1421, g1423, g1427, g1428, g1429, g1430, g1431, g1432, g1433, g1434;
	wire g1435, g1436, g1438, g1439, g1440, g1441, g1442, g1443, g1444, g1445, g1446, g1447, g1448, g1450, g1461, g1462, g1463, g1464, g1465, g1466, g1468;
	wire g1469, g1470, g1472, g1471, g1475, g1473, g1474, g1476, g1477, g1479, g1480, g1481, g1482, g1485, g1483, g1484, g1486, g1487, g1489, g1490, g1491;
	wire g1494, g1492, g1493, g1497, g1498, g1495, g1496, g1499, g1500, g1502, g1503, g1504, g1505, g1508, g1506, g1507, g1509, g1510, g1512, g1513, g1514;
	wire g1515, g1516, g1517, g1519, g1520, g1521, g1524, g1522, g1523, g1527, g1528, g1525, g1526, g1529, g1530, g1532, g1533, g1534, g1537, g1535, g1536;
	wire g1540, g1538, g1539, g1541, g1542, g1544, g1545, g1546, g1549, g1547, g1548, g1550, g1551, g1552, g1553, g1555, g1556, g1557, g1558, g1561, g1559;
	wire g1560, g1562, g1563, g1565, g1566, g1567, g1570, g1568, g1569, g1573, g1574, g1571, g1572, g1575, g1576, g1578, g1579, g1580, g1581, g1582, g1583;
	wire g1585, g1586, g1587, g1589, g1588, g1591, g1590, g1592, g1594, g1595, g1596, g1599, g1597, g1598, g1602, g1603, g1600, g1601, g1604, g1605, g1607;
	wire g1608, g1609, g1610, g1611, g1612, g1614, g1615, g1616, g1619, g1617, g1618, g1622, g1623, g1620, g1621, g1624, g1626, g1627, g1628, g1629, g1630;
	wire g1631, g1633, g1634, g1635, g1636, g1637, g1638, g1640, g1641, g1642, g1643, g1646, g1644, g1645, g1647, g1648;

	lut_sub lut_5 ({g9}, o_0_);
	defparam lut_5.LUT_SIZE = 1;
	defparam lut_5.mask = 2'b10;

	lut_sub lut_9 ({g11}, o_1_);
	defparam lut_9.LUT_SIZE = 1;
	defparam lut_9.mask = 2'b10;

	lut_sub lut_13 ({g52}, o_3_);
	defparam lut_13.LUT_SIZE = 1;
	defparam lut_13.mask = 2'b10;

	lut_sub lut_17 ({g456}, o_5_);
	defparam lut_17.LUT_SIZE = 1;
	defparam lut_17.mask = 2'b10;

	lut_sub lut_21 ({g458}, o_6_);
	defparam lut_21.LUT_SIZE = 1;
	defparam lut_21.mask = 2'b10;

	lut_sub lut_25 ({g621}, o_7_);
	defparam lut_25.LUT_SIZE = 1;
	defparam lut_25.mask = 2'b10;

	lut_sub lut_29 ({g812}, o_9_);
	defparam lut_29.LUT_SIZE = 1;
	defparam lut_29.mask = 2'b10;

	lut_sub lut_33 ({g845}, o_10_);
	defparam lut_33.LUT_SIZE = 1;
	defparam lut_33.mask = 2'b10;

	lut_sub lut_37 ({g846}, o_11_);
	defparam lut_37.LUT_SIZE = 1;
	defparam lut_37.mask = 2'b10;

	lut_sub lut_41 ({g923}, o_12_);
	defparam lut_41.LUT_SIZE = 1;
	defparam lut_41.mask = 2'b10;

	lut_sub lut_45 ({g963}, o_13_);
	defparam lut_45.LUT_SIZE = 1;
	defparam lut_45.mask = 2'b10;

	lut_sub lut_49 ({g989}, o_14_);
	defparam lut_49.LUT_SIZE = 1;
	defparam lut_49.mask = 2'b10;

	lut_sub lut_53 ({g1003}, o_15_);
	defparam lut_53.LUT_SIZE = 1;
	defparam lut_53.mask = 2'b10;

	lut_sub lut_57 ({g1456}, o_16_);
	defparam lut_57.LUT_SIZE = 1;
	defparam lut_57.mask = 2'b10;

	lut_sub lut_61 ({g1018}, o_17_);
	defparam lut_61.LUT_SIZE = 1;
	defparam lut_61.mask = 2'b10;

	lut_sub lut_65 ({g1057}, o_18_);
	defparam lut_65.LUT_SIZE = 1;
	defparam lut_65.mask = 2'b10;

	lut_sub lut_69 ({g1454}, o_22_);
	defparam lut_69.LUT_SIZE = 1;
	defparam lut_69.mask = 2'b10;

	lut_sub lut_73 ({g1077}, o_23_);
	defparam lut_73.LUT_SIZE = 1;
	defparam lut_73.mask = 2'b10;

	lut_sub lut_77 ({g1125}, o_32_);
	defparam lut_77.LUT_SIZE = 1;
	defparam lut_77.mask = 2'b10;

	lut_sub lut_81 ({g1128}, o_33_);
	defparam lut_81.LUT_SIZE = 1;
	defparam lut_81.mask = 2'b10;

	lut_sub lut_85 ({g1129}, o_34_);
	defparam lut_85.LUT_SIZE = 1;
	defparam lut_85.mask = 2'b10;

	lut_sub lut_89 ({g1253}, o_35_);
	defparam lut_89.LUT_SIZE = 1;
	defparam lut_89.mask = 2'b10;

	lut_sub lut_93 ({g1346}, o_36_);
	defparam lut_93.LUT_SIZE = 1;
	defparam lut_93.mask = 2'b10;

	lut_sub lut_97 ({g1393}, o_37_);
	defparam lut_97.LUT_SIZE = 1;
	defparam lut_97.mask = 2'b10;

	lut_sub lut_101 ({g1417}, o_38_);
	defparam lut_101.LUT_SIZE = 1;
	defparam lut_101.mask = 2'b10;

	lut_sub lut_105 ({g1422}, o_39_);
	defparam lut_105.LUT_SIZE = 1;
	defparam lut_105.mask = 2'b10;

	lut_sub lut_109 ({g1424}, o_40_);
	defparam lut_109.LUT_SIZE = 1;
	defparam lut_109.mask = 2'b10;

	lut_sub lut_113 ({g1426}, o_42_);
	defparam lut_113.LUT_SIZE = 1;
	defparam lut_113.mask = 2'b10;

	lut_sub lut_117 ({g1437}, o_43_);
	defparam lut_117.LUT_SIZE = 1;
	defparam lut_117.mask = 2'b10;

	lut_sub lut_121 ({g1449}, o_44_);
	defparam lut_121.LUT_SIZE = 1;
	defparam lut_121.mask = 2'b10;

	lut_sub lut_125 ({g1451}, o_45_);
	defparam lut_125.LUT_SIZE = 1;
	defparam lut_125.mask = 2'b10;

	lut_sub lut_129 ({i_6_, i_7_}, g1);
	defparam lut_129.LUT_SIZE = 2;
	defparam lut_129.mask = 4'b1000;

	lut_sub lut_134 ({i_8_, g1}, g2);
	defparam lut_134.LUT_SIZE = 2;
	defparam lut_134.mask = 4'b0100;

	lut_sub lut_138 ({i_9_, i_10_, i_11_, i_15_}, g3);
	defparam lut_138.LUT_SIZE = 4;
	defparam lut_138.mask = 16'h8000;

	lut_sub lut_142 ({i_12_, i_13_, i_14_}, g4);
	defparam lut_142.LUT_SIZE = 3;
	defparam lut_142.mask = 8'h80;

	lut_sub lut_148 ({g3, g4}, g5);
	defparam lut_148.LUT_SIZE = 2;
	defparam lut_148.mask = 4'b0001;

	lut_sub lut_152 ({i_4_, i_3_, i_5_}, g6);
	defparam lut_152.LUT_SIZE = 3;
	defparam lut_152.mask = 8'h40;

	lut_sub lut_157 ({i_0_, i_1_, g6, i_2_}, g7);
	defparam lut_157.LUT_SIZE = 4;
	defparam lut_157.mask = 16'h0002;

	lut_sub lut_163 ({g5, g7}, g8);
	defparam lut_163.LUT_SIZE = 2;
	defparam lut_163.mask = 4'b0001;

	lut_sub lut_169 ({i_0_, i_1_, g2, g8}, g9);
	defparam lut_169.LUT_SIZE = 4;
	defparam lut_169.mask = 16'hee0e;

	lut_sub lut_181 ({i_6_, i_7_}, g10);
	defparam lut_181.LUT_SIZE = 2;
	defparam lut_181.mask = 4'b0100;

	lut_sub lut_187 ({i_0_, i_1_, i_8_, i_2_, g8, g10}, g11);
	defparam lut_187.LUT_SIZE = 6;
	defparam lut_187.mask = 64'he0f0e0f00e0feeff;

	lut_sub lut_226 ({i_0_, i_1_, g5, i_2_}, g12);
	defparam lut_226.LUT_SIZE = 4;
	defparam lut_226.mask = 16'h0002;

	lut_sub lut_232 ({i_8_, i_6_, g6, g12}, o_2_);
	defparam lut_232.LUT_SIZE = 4;
	defparam lut_232.mask = 16'h1000;

	lut_sub lut_236 ({i_0_, i_1_, i_2_}, g14);
	defparam lut_236.LUT_SIZE = 3;
	defparam lut_236.mask = 8'h20;

	lut_sub lut_240 ({i_4_, i_3_, i_5_}, g15);
	defparam lut_240.LUT_SIZE = 3;
	defparam lut_240.mask = 8'h80;

	lut_sub lut_246 ({g14, g15}, g16);
	defparam lut_246.LUT_SIZE = 2;
	defparam lut_246.mask = 4'b0001;

	lut_sub lut_250 ({i_9_, i_10_, i_11_, i_15_}, g17);
	defparam lut_250.LUT_SIZE = 4;
	defparam lut_250.mask = 16'h0040;

	lut_sub lut_256 ({g4, g17}, g18);
	defparam lut_256.LUT_SIZE = 2;
	defparam lut_256.mask = 4'b0001;

	lut_sub lut_260 ({i_12_, i_13_, i_14_}, g19);
	defparam lut_260.LUT_SIZE = 3;
	defparam lut_260.mask = 8'h20;

	lut_sub lut_264 ({i_9_, i_10_, i_11_, i_15_}, g20);
	defparam lut_264.LUT_SIZE = 4;
	defparam lut_264.mask = 16'h0800;

	lut_sub lut_270 ({g19, g20}, g21);
	defparam lut_270.LUT_SIZE = 2;
	defparam lut_270.mask = 4'b0001;

	lut_sub lut_274 ({i_9_, i_10_, i_11_, i_15_}, g22);
	defparam lut_274.LUT_SIZE = 4;
	defparam lut_274.mask = 16'hfbff;

	lut_sub lut_294 ({g4, g22}, g23);
	defparam lut_294.LUT_SIZE = 2;
	defparam lut_294.mask = 4'b1101;

	lut_sub lut_300 ({i_12_, i_13_, i_14_}, g24);
	defparam lut_300.LUT_SIZE = 3;
	defparam lut_300.mask = 8'hbf;

	lut_sub lut_312 ({g20, g24}, g25);
	defparam lut_312.LUT_SIZE = 2;
	defparam lut_312.mask = 4'b1101;

	lut_sub lut_322 ({g18, g21, g23, g25}, g26);
	defparam lut_322.LUT_SIZE = 4;
	defparam lut_322.mask = 16'h1000;

	lut_sub lut_326 ({i_9_, i_10_, i_11_, i_15_}, g27);
	defparam lut_326.LUT_SIZE = 4;
	defparam lut_326.mask = 16'h0080;

	lut_sub lut_332 ({g24, g27}, g28);
	defparam lut_332.LUT_SIZE = 2;
	defparam lut_332.mask = 4'b0100;

	lut_sub lut_340 ({g2, g10, g26, g28}, g29);
	defparam lut_340.LUT_SIZE = 4;
	defparam lut_340.mask = 16'hf020;

	lut_sub lut_349 ({i_8_, g1}, g30);
	defparam lut_349.LUT_SIZE = 2;
	defparam lut_349.mask = 4'b0001;

	lut_sub lut_356 ({g4, g20, g27}, g31);
	defparam lut_356.LUT_SIZE = 3;
	defparam lut_356.mask = 8'h07;

	lut_sub lut_367 ({g5, g16, g29, g30, g31}, g32);
	defparam lut_367.LUT_SIZE = 5;
	defparam lut_367.mask = 32'h00f100f3;

	lut_sub lut_383 ({g19, g27}, g33);
	defparam lut_383.LUT_SIZE = 2;
	defparam lut_383.mask = 4'b0001;

	lut_sub lut_387 ({i_9_, i_10_}, g34);
	defparam lut_387.LUT_SIZE = 2;
	defparam lut_387.mask = 4'b0001;

	lut_sub lut_392 ({i_11_, i_15_, g34}, g35);
	defparam lut_392.LUT_SIZE = 3;
	defparam lut_392.mask = 8'h40;

	lut_sub lut_396 ({i_9_, i_10_, i_11_, i_15_}, g36);
	defparam lut_396.LUT_SIZE = 4;
	defparam lut_396.mask = 16'h0004;

	lut_sub lut_402 ({g4, g36}, g37);
	defparam lut_402.LUT_SIZE = 2;
	defparam lut_402.mask = 4'b1110;

	lut_sub lut_412 ({g19, g24, g35, g37}, g38);
	defparam lut_412.LUT_SIZE = 4;
	defparam lut_412.mask = 16'h4544;

	lut_sub lut_424 ({g2, g16, g33, g38}, g39);
	defparam lut_424.LUT_SIZE = 4;
	defparam lut_424.mask = 16'h000b;

	lut_sub lut_430 ({i_0_, i_1_, i_3_}, g40);
	defparam lut_430.LUT_SIZE = 3;
	defparam lut_430.mask = 8'h08;

	lut_sub lut_436 ({i_4_, g39, g40}, g41);
	defparam lut_436.LUT_SIZE = 3;
	defparam lut_436.mask = 8'h8c;

	lut_sub lut_442 ({i_6_, i_7_}, g42);
	defparam lut_442.LUT_SIZE = 2;
	defparam lut_442.mask = 4'b0010;

	lut_sub lut_447 ({i_8_, g42}, g43);
	defparam lut_447.LUT_SIZE = 2;
	defparam lut_447.mask = 4'b0100;

	lut_sub lut_455 ({g16, g43, g33, g38}, g44);
	defparam lut_455.LUT_SIZE = 4;
	defparam lut_455.mask = 16'h000b;

	lut_sub lut_461 ({i_6_, i_7_}, g45);
	defparam lut_461.LUT_SIZE = 2;
	defparam lut_461.mask = 4'b0001;

	lut_sub lut_469 ({g16, g26, g43, g45}, g46);
	defparam lut_469.LUT_SIZE = 4;
	defparam lut_469.mask = 16'h0075;

	lut_sub lut_480 ({i_8_, g4, g16, g24}, g47);
	defparam lut_480.LUT_SIZE = 4;
	defparam lut_480.mask = 16'h2203;

	lut_sub lut_489 ({g4, g20}, g48);
	defparam lut_489.LUT_SIZE = 2;
	defparam lut_489.mask = 4'b0001;

	lut_sub lut_494 ({i_8_, g42}, g49);
	defparam lut_494.LUT_SIZE = 2;
	defparam lut_494.mask = 4'b0001;

	lut_sub lut_502 ({g5, g16, g48, g49}, g50);
	defparam lut_502.LUT_SIZE = 4;
	defparam lut_502.mask = 16'h0105;

	lut_sub lut_514 ({g27, g42, g44, g46, g47, g50}, g51);
	defparam lut_514.LUT_SIZE = 6;
	defparam lut_514.mask = 64'ha000a000a0008000;

	lut_sub lut_527 ({g32, g41, g51}, g52);
	defparam lut_527.LUT_SIZE = 3;
	defparam lut_527.mask = 8'h10;

	lut_sub lut_531 ({i_9_, i_10_}, g53);
	defparam lut_531.LUT_SIZE = 2;
	defparam lut_531.mask = 4'b0110;

	lut_sub lut_536 ({i_4_, i_3_, i_5_}, g54);
	defparam lut_536.LUT_SIZE = 3;
	defparam lut_536.mask = 8'h08;

	lut_sub lut_542 ({g14, g54}, g55);
	defparam lut_542.LUT_SIZE = 2;
	defparam lut_542.mask = 4'b0001;

	lut_sub lut_546 ({i_12_, i_13_, i_14_}, g56);
	defparam lut_546.LUT_SIZE = 3;
	defparam lut_546.mask = 8'h60;

	lut_sub lut_556 ({g2, g35, g37, g55, g56}, g57);
	defparam lut_556.LUT_SIZE = 5;
	defparam lut_556.mask = 32'h00003031;

	lut_sub lut_566 ({i_0_, i_1_, i_2_, g10, g54}, g58);
	defparam lut_566.LUT_SIZE = 5;
	defparam lut_566.mask = 32'h00105500;

	lut_sub lut_580 ({g2, g26, g28, g33, g55, g58}, g59);
	defparam lut_580.LUT_SIZE = 6;
	defparam lut_580.mask = 64'haaaaaaaa8888a888;

	lut_sub lut_609 ({i_11_, i_15_, g4}, g60);
	defparam lut_609.LUT_SIZE = 3;
	defparam lut_609.mask = 8'h40;

	lut_sub lut_619 ({g30, g53, g55, g57, g59, g60}, g61);
	defparam lut_619.LUT_SIZE = 6;
	defparam lut_619.mask = 64'h3030303030303020;

	lut_sub lut_637 ({i_4_, i_3_, i_5_}, g62);
	defparam lut_637.LUT_SIZE = 3;
	defparam lut_637.mask = 8'h04;

	lut_sub lut_642 ({i_0_, i_1_, g62}, g63);
	defparam lut_642.LUT_SIZE = 3;
	defparam lut_642.mask = 8'h04;

	lut_sub lut_651 ({g26, g28, g43, g33, g55}, g64);
	defparam lut_651.LUT_SIZE = 5;
	defparam lut_651.mask = 32'h05050105;

	lut_sub lut_664 ({i_6_, i_7_, g55, g63, g64}, g65);
	defparam lut_664.LUT_SIZE = 5;
	defparam lut_664.mask = 32'h88888880;

	lut_sub lut_679 ({i_8_, g31, g42, g38, g55, g65}, g66);
	defparam lut_679.LUT_SIZE = 6;
	defparam lut_679.mask = 64'h5545554555555544;

	lut_sub lut_712 ({g61, g66}, o_4_);
	defparam lut_712.LUT_SIZE = 2;
	defparam lut_712.mask = 4'b1110;

	lut_sub lut_718 ({i_12_, i_13_, i_14_}, g68);
	defparam lut_718.LUT_SIZE = 3;
	defparam lut_718.mask = 8'hf7;

	lut_sub lut_728 ({i_9_, i_10_, i_11_, i_15_}, g69);
	defparam lut_728.LUT_SIZE = 4;
	defparam lut_728.mask = 16'h4000;

	lut_sub lut_734 ({g68, g69}, g70);
	defparam lut_734.LUT_SIZE = 2;
	defparam lut_734.mask = 4'b0100;

	lut_sub lut_738 ({i_0_, i_1_, i_2_}, g71);
	defparam lut_738.LUT_SIZE = 3;
	defparam lut_738.mask = 8'h80;

	lut_sub lut_744 ({g62, g71}, g72);
	defparam lut_744.LUT_SIZE = 2;
	defparam lut_744.mask = 4'b0001;

	lut_sub lut_750 ({g10, g72}, g73);
	defparam lut_750.LUT_SIZE = 2;
	defparam lut_750.mask = 4'b0001;

	lut_sub lut_755 ({i_8_, g73}, g74);
	defparam lut_755.LUT_SIZE = 2;
	defparam lut_755.mask = 4'b0100;

	lut_sub lut_760 ({i_8_, g73}, g75);
	defparam lut_760.LUT_SIZE = 2;
	defparam lut_760.mask = 4'b1110;

	lut_sub lut_766 ({i_12_, i_13_, i_14_}, g76);
	defparam lut_766.LUT_SIZE = 3;
	defparam lut_766.mask = 8'hef;

	lut_sub lut_778 ({g3, g76}, g77);
	defparam lut_778.LUT_SIZE = 2;
	defparam lut_778.mask = 4'b0010;

	lut_sub lut_784 ({g22, g68}, g78);
	defparam lut_784.LUT_SIZE = 2;
	defparam lut_784.mask = 4'b0111;

	lut_sub lut_792 ({g20, g76}, g79);
	defparam lut_792.LUT_SIZE = 2;
	defparam lut_792.mask = 4'b1101;

	lut_sub lut_798 ({i_9_, i_10_}, g80);
	defparam lut_798.LUT_SIZE = 2;
	defparam lut_798.mask = 4'b1000;

	lut_sub lut_803 ({g80, i_11_, i_15_}, g81);
	defparam lut_803.LUT_SIZE = 3;
	defparam lut_803.mask = 8'h01;

	lut_sub lut_809 ({g68, g81}, g82);
	defparam lut_809.LUT_SIZE = 2;
	defparam lut_809.mask = 4'b0100;

	lut_sub lut_814 ({g80, i_11_, i_15_}, g83);
	defparam lut_814.LUT_SIZE = 3;
	defparam lut_814.mask = 8'h02;

	lut_sub lut_822 ({i_8_, g73, g76, g82, g83}, g84);
	defparam lut_822.LUT_SIZE = 5;
	defparam lut_822.mask = 32'h00000073;

	lut_sub lut_836 ({g75, g77, g70, g78, g79, g84}, g85);
	defparam lut_836.LUT_SIZE = 6;
	defparam lut_836.mask = 64'h02000000aaaaaaaa;

	lut_sub lut_856 ({i_9_, i_10_, i_11_, i_15_}, g86);
	defparam lut_856.LUT_SIZE = 4;
	defparam lut_856.mask = 16'h0020;

	lut_sub lut_862 ({g76, g86}, g87);
	defparam lut_862.LUT_SIZE = 2;
	defparam lut_862.mask = 4'b1011;

	lut_sub lut_868 ({i_9_, i_10_, i_11_, i_15_}, g88);
	defparam lut_868.LUT_SIZE = 4;
	defparam lut_868.mask = 16'h0010;

	lut_sub lut_874 ({g68, g88}, g89);
	defparam lut_874.LUT_SIZE = 2;
	defparam lut_874.mask = 4'b1011;

	lut_sub lut_882 ({g36, g68}, g90);
	defparam lut_882.LUT_SIZE = 2;
	defparam lut_882.mask = 4'b0010;

	lut_sub lut_886 ({i_9_, i_10_, i_11_, i_15_}, g91);
	defparam lut_886.LUT_SIZE = 4;
	defparam lut_886.mask = 16'hfffe;

	lut_sub lut_906 ({g68, g91}, g92);
	defparam lut_906.LUT_SIZE = 2;
	defparam lut_906.mask = 4'b1000;

	lut_sub lut_911 ({i_15_, g76}, g93);
	defparam lut_911.LUT_SIZE = 2;
	defparam lut_911.mask = 4'b1000;

	lut_sub lut_917 ({g80, g93}, g94);
	defparam lut_917.LUT_SIZE = 2;
	defparam lut_917.mask = 4'b0001;

	lut_sub lut_926 ({i_8_, g73, g90, g82, g92, g94}, g95);
	defparam lut_926.LUT_SIZE = 6;
	defparam lut_926.mask = 64'h00007fff000000ff;

	lut_sub lut_958 ({g87, g78, g74, g79, g89, g95}, g96);
	defparam lut_958.LUT_SIZE = 6;
	defparam lut_958.mask = 64'haa00aa00aa00aa02;

	lut_sub lut_980 ({g17, g68}, g97);
	defparam lut_980.LUT_SIZE = 2;
	defparam lut_980.mask = 4'b1101;

	lut_sub lut_988 ({g27, g76}, g98);
	defparam lut_988.LUT_SIZE = 2;
	defparam lut_988.mask = 4'b0010;

	lut_sub lut_995 ({g73, g97, g98}, g99);
	defparam lut_995.LUT_SIZE = 3;
	defparam lut_995.mask = 8'h0d;

	lut_sub lut_1006 ({g70, g74, g85, g96, g99}, g100);
	defparam lut_1006.LUT_SIZE = 5;
	defparam lut_1006.mask = 32'h02020200;

	lut_sub lut_1012 ({i_8_, i_6_, i_7_}, g101);
	defparam lut_1012.LUT_SIZE = 3;
	defparam lut_1012.mask = 8'h10;

	lut_sub lut_1018 ({g72, g101}, g102);
	defparam lut_1018.LUT_SIZE = 2;
	defparam lut_1018.mask = 4'b0001;

	lut_sub lut_1026 ({g76, g102, g82, g83}, g103);
	defparam lut_1026.LUT_SIZE = 4;
	defparam lut_1026.mask = 16'h0703;

	lut_sub lut_1037 ({g87, g102, g89}, g104);
	defparam lut_1037.LUT_SIZE = 3;
	defparam lut_1037.mask = 8'h32;

	lut_sub lut_1045 ({i_8_, g45, g72}, g105);
	defparam lut_1045.LUT_SIZE = 3;
	defparam lut_1045.mask = 8'hfe;

	lut_sub lut_1059 ({g76, g82, g83, g105}, g106);
	defparam lut_1059.LUT_SIZE = 4;
	defparam lut_1059.mask = 16'h2a0a;

	lut_sub lut_1068 ({i_11_, i_15_, g34}, g107);
	defparam lut_1068.LUT_SIZE = 3;
	defparam lut_1068.mask = 8'hfb;

	lut_sub lut_1080 ({g76, g107}, g108);
	defparam lut_1080.LUT_SIZE = 2;
	defparam lut_1080.mask = 4'b1000;

	lut_sub lut_1086 ({g35, g76}, g109);
	defparam lut_1086.LUT_SIZE = 2;
	defparam lut_1086.mask = 4'b0010;

	lut_sub lut_1096 ({g108, g109, g90, g98, g102, g78}, g110);
	defparam lut_1096.LUT_SIZE = 6;
	defparam lut_1096.mask = 64'h2333333333333333;

	lut_sub lut_1134 ({g103, g104, g106, g110}, g111);
	defparam lut_1134.LUT_SIZE = 4;
	defparam lut_1134.mask = 16'h8000;

	lut_sub lut_1138 ({i_9_, i_10_, i_11_}, g112);
	defparam lut_1138.LUT_SIZE = 3;
	defparam lut_1138.mask = 8'h10;

	lut_sub lut_1143 ({i_15_, g112}, g113);
	defparam lut_1143.LUT_SIZE = 2;
	defparam lut_1143.mask = 4'b1110;

	lut_sub lut_1151 ({g68, g113}, g114);
	defparam lut_1151.LUT_SIZE = 2;
	defparam lut_1151.mask = 4'b0111;

	lut_sub lut_1161 ({g109, g90, g77, g105}, g115);
	defparam lut_1161.LUT_SIZE = 4;
	defparam lut_1161.mask = 16'h2aaa;

	lut_sub lut_1176 ({g102, g92, g79, g114, g115}, g116);
	defparam lut_1176.LUT_SIZE = 5;
	defparam lut_1176.mask = 32'haaaa0200;

	lut_sub lut_1190 ({g111, g116}, g117);
	defparam lut_1190.LUT_SIZE = 2;
	defparam lut_1190.mask = 4'b0001;

	lut_sub lut_1196 ({g6, g71}, g118);
	defparam lut_1196.LUT_SIZE = 2;
	defparam lut_1196.mask = 4'b0001;

	lut_sub lut_1202 ({i_8_, g10, g118}, g119);
	defparam lut_1202.LUT_SIZE = 3;
	defparam lut_1202.mask = 8'h01;

	lut_sub lut_1208 ({g54, g71}, g120);
	defparam lut_1208.LUT_SIZE = 2;
	defparam lut_1208.mask = 4'b0001;

	lut_sub lut_1214 ({i_8_, g45, g120}, g121);
	defparam lut_1214.LUT_SIZE = 3;
	defparam lut_1214.mask = 8'h01;

	lut_sub lut_1220 ({g49, g118}, g122);
	defparam lut_1220.LUT_SIZE = 2;
	defparam lut_1220.mask = 4'b0001;

	lut_sub lut_1226 ({g30, g118}, g123);
	defparam lut_1226.LUT_SIZE = 2;
	defparam lut_1226.mask = 4'b1110;

	lut_sub lut_1236 ({g70, g122, g123, g114}, g124);
	defparam lut_1236.LUT_SIZE = 4;
	defparam lut_1236.mask = 16'h0ace;

	lut_sub lut_1248 ({g49, g120}, g125);
	defparam lut_1248.LUT_SIZE = 2;
	defparam lut_1248.mask = 4'b0001;

	lut_sub lut_1253 ({i_15_, g112}, g126);
	defparam lut_1253.LUT_SIZE = 2;
	defparam lut_1253.mask = 4'b1011;

	lut_sub lut_1261 ({g76, g126}, g127);
	defparam lut_1261.LUT_SIZE = 2;
	defparam lut_1261.mask = 4'b1000;

	lut_sub lut_1270 ({g125, g77, g127, g123, g119}, g128);
	defparam lut_1270.LUT_SIZE = 5;
	defparam lut_1270.mask = 32'hff22f020;

	lut_sub lut_1293 ({g70, g119, g121, g124, g128}, g129);
	defparam lut_1293.LUT_SIZE = 5;
	defparam lut_1293.mask = 32'h44444000;

	lut_sub lut_1303 ({g2, g118}, g130);
	defparam lut_1303.LUT_SIZE = 2;
	defparam lut_1303.mask = 4'b1110;

	lut_sub lut_1311 ({g43, g120}, g131);
	defparam lut_1311.LUT_SIZE = 2;
	defparam lut_1311.mask = 4'b1110;

	lut_sub lut_1321 ({i_8_, g73, g108, g92, g1639}, g132);
	defparam lut_1321.LUT_SIZE = 5;
	defparam lut_1321.mask = 32'h55505544;

	lut_sub lut_1339 ({g108, g92, g123}, g133);
	defparam lut_1339.LUT_SIZE = 3;
	defparam lut_1339.mask = 8'h2a;

	lut_sub lut_1348 ({g108, g92, g130}, g134);
	defparam lut_1348.LUT_SIZE = 3;
	defparam lut_1348.mask = 8'h2a;

	lut_sub lut_1356 ({g43, g118}, g135);
	defparam lut_1356.LUT_SIZE = 2;
	defparam lut_1356.mask = 4'b1110;

	lut_sub lut_1366 ({g76, g122, g82, g83}, g136);
	defparam lut_1366.LUT_SIZE = 4;
	defparam lut_1366.mask = 16'h0703;

	lut_sub lut_1378 ({g78, g135, g122, g89}, g137);
	defparam lut_1378.LUT_SIZE = 4;
	defparam lut_1378.mask = 16'hb3a0;

	lut_sub lut_1394 ({g97, g98, g135, g122, g136, g137}, g138);
	defparam lut_1394.LUT_SIZE = 6;
	defparam lut_1394.mask = 64'h0080008088880080;

	lut_sub lut_1408 ({g76, g82, g83, g130}, g139);
	defparam lut_1408.LUT_SIZE = 4;
	defparam lut_1408.mask = 16'h2a0a;

	lut_sub lut_1419 ({g109, g90, g130}, g140);
	defparam lut_1419.LUT_SIZE = 3;
	defparam lut_1419.mask = 8'h2a;

	lut_sub lut_1429 ({g87, g127, g79, g123}, g141);
	defparam lut_1429.LUT_SIZE = 4;
	defparam lut_1429.mask = 16'haa8a;

	lut_sub lut_1441 ({i_8_, g10, g118}, g142);
	defparam lut_1441.LUT_SIZE = 3;
	defparam lut_1441.mask = 8'hef;

	lut_sub lut_1454 ({g97, g82, g142}, g143);
	defparam lut_1454.LUT_SIZE = 3;
	defparam lut_1454.mask = 8'ha2;

	lut_sub lut_1462 ({g42, g120}, g144);
	defparam lut_1462.LUT_SIZE = 2;
	defparam lut_1462.mask = 4'b0001;

	lut_sub lut_1471 ({g87, g144, g122, g89, g105}, g145);
	defparam lut_1471.LUT_SIZE = 5;
	defparam lut_1471.mask = 32'h51117333;

	lut_sub lut_1493 ({g139, g140, g141, g143, g145}, g146);
	defparam lut_1493.LUT_SIZE = 5;
	defparam lut_1493.mask = 32'h40000000;

	lut_sub lut_1500 ({g109, g90, g123}, g147);
	defparam lut_1500.LUT_SIZE = 3;
	defparam lut_1500.mask = 8'h2a;

	lut_sub lut_1509 ({g97, g98, g105}, g148);
	defparam lut_1509.LUT_SIZE = 3;
	defparam lut_1509.mask = 8'ha2;

	lut_sub lut_1521 ({g127, g78, g135, g79, g114, g105}, g149);
	defparam lut_1521.LUT_SIZE = 6;
	defparam lut_1521.mask = 64'h1155135711551155;

	lut_sub lut_1556 ({g77, g97, g102, g147, g148, g149}, g150);
	defparam lut_1556.LUT_SIZE = 6;
	defparam lut_1556.mask = 64'h4000404040004000;

	lut_sub lut_1565 ({i_9_, i_10_, i_11_, g142}, g151);
	defparam lut_1565.LUT_SIZE = 4;
	defparam lut_1565.mask = 16'h2080;

	lut_sub lut_1575 ({g73, g127, g93, g114, g151}, g152);
	defparam lut_1575.LUT_SIZE = 5;
	defparam lut_1575.mask = 32'hfafa3200;

	lut_sub lut_1599 ({g133, g134, g138, g146, g150, g152}, g153);
	defparam lut_1599.LUT_SIZE = 6;
	defparam lut_1599.mask = 64'h0001000000000000;

	lut_sub lut_1605 ({i_8_, g10, g120}, g154);
	defparam lut_1605.LUT_SIZE = 3;
	defparam lut_1605.mask = 8'hfe;

	lut_sub lut_1618 ({g125, g154, g122}, g155);
	defparam lut_1618.LUT_SIZE = 3;
	defparam lut_1618.mask = 8'h20;

	lut_sub lut_1626 ({i_15_, g34, g108, g68, g155}, g156);
	defparam lut_1626.LUT_SIZE = 5;
	defparam lut_1626.mask = 32'h0a0a0a8a;

	lut_sub lut_1640 ({g43, g72}, g157);
	defparam lut_1640.LUT_SIZE = 2;
	defparam lut_1640.mask = 4'b0001;

	lut_sub lut_1648 ({g157, g90, g78, g135}, g158);
	defparam lut_1648.LUT_SIZE = 4;
	defparam lut_1648.mask = 16'h888f;

	lut_sub lut_1660 ({i_8_, g10, g120}, g159);
	defparam lut_1660.LUT_SIZE = 3;
	defparam lut_1660.mask = 8'hef;

	lut_sub lut_1674 ({g87, g98, g144, g159}, g160);
	defparam lut_1674.LUT_SIZE = 4;
	defparam lut_1674.mask = 16'hab03;

	lut_sub lut_1686 ({g49, g72}, g161);
	defparam lut_1686.LUT_SIZE = 2;
	defparam lut_1686.mask = 4'b0001;

	lut_sub lut_1695 ({i_8_, g73, g108, g109, g154, g122}, g162);
	defparam lut_1695.LUT_SIZE = 6;
	defparam lut_1695.mask = 64'hf2f2f0f0f2f2f000;

	lut_sub lut_1736 ({g109, g161, g87, g125, g78, g162}, g163);
	defparam lut_1736.LUT_SIZE = 6;
	defparam lut_1736.mask = 64'h5051505150500000;

	lut_sub lut_1755 ({g30, g120}, g164);
	defparam lut_1755.LUT_SIZE = 2;
	defparam lut_1755.mask = 4'b0001;

	lut_sub lut_1761 ({g42, g118}, g165);
	defparam lut_1761.LUT_SIZE = 2;
	defparam lut_1761.mask = 4'b0001;

	lut_sub lut_1766 ({i_4_, i_3_, i_5_, g71}, g166);
	defparam lut_1766.LUT_SIZE = 4;
	defparam lut_1766.mask = 16'h1040;

	lut_sub lut_1773 ({g101, g166}, g167);
	defparam lut_1773.LUT_SIZE = 2;
	defparam lut_1773.mask = 4'b0001;

	lut_sub lut_1779 ({g45, g72}, g168);
	defparam lut_1779.LUT_SIZE = 2;
	defparam lut_1779.mask = 4'b0001;

	lut_sub lut_1785 ({i_8_, i_6_, g120, g77}, g169);
	defparam lut_1785.LUT_SIZE = 4;
	defparam lut_1785.mask = 16'h0001;

	lut_sub lut_1795 ({g125, g167, g97, g70, g168, g169}, g170);
	defparam lut_1795.LUT_SIZE = 6;
	defparam lut_1795.mask = 64'ha8a800a8a0a000a0;

	lut_sub lut_1819 ({g87, g127, g164, g102, g165, g170}, g171);
	defparam lut_1819.LUT_SIZE = 6;
	defparam lut_1819.mask = 64'h4444400055555000;

	lut_sub lut_1842 ({g156, g158, g160, g163, g171}, g172);
	defparam lut_1842.LUT_SIZE = 5;
	defparam lut_1842.mask = 32'h10000000;

	lut_sub lut_1852 ({g100, g117, g129, g132, g153, g172}, g173);
	defparam lut_1852.LUT_SIZE = 6;
	defparam lut_1852.mask = 64'h0000000000000001;

	lut_sub lut_1856 ({i_12_, i_13_, i_14_}, g174);
	defparam lut_1856.LUT_SIZE = 3;
	defparam lut_1856.mask = 8'hfe;

	lut_sub lut_1868 ({g20, g174}, g175);
	defparam lut_1868.LUT_SIZE = 2;
	defparam lut_1868.mask = 4'b0010;

	lut_sub lut_1872 ({i_12_, i_13_, i_14_}, g176);
	defparam lut_1872.LUT_SIZE = 3;
	defparam lut_1872.mask = 8'hfb;

	lut_sub lut_1884 ({g22, g176}, g177);
	defparam lut_1884.LUT_SIZE = 2;
	defparam lut_1884.mask = 4'b1000;

	lut_sub lut_1891 ({g75, g175, g177}, g178);
	defparam lut_1891.LUT_SIZE = 3;
	defparam lut_1891.mask = 8'h70;

	lut_sub lut_1899 ({g17, g176}, g179);
	defparam lut_1899.LUT_SIZE = 2;
	defparam lut_1899.mask = 4'b0010;

	lut_sub lut_1905 ({g27, g174}, g180);
	defparam lut_1905.LUT_SIZE = 2;
	defparam lut_1905.mask = 4'b0010;

	lut_sub lut_1912 ({g75, g179, g180}, g181);
	defparam lut_1912.LUT_SIZE = 3;
	defparam lut_1912.mask = 8'h70;

	lut_sub lut_1920 ({g81, g176}, g182);
	defparam lut_1920.LUT_SIZE = 2;
	defparam lut_1920.mask = 4'b0010;

	lut_sub lut_1926 ({g83, g174}, g183);
	defparam lut_1926.LUT_SIZE = 2;
	defparam lut_1926.mask = 4'b0010;

	lut_sub lut_1933 ({g74, g182, g183}, g184);
	defparam lut_1933.LUT_SIZE = 3;
	defparam lut_1933.mask = 8'h07;

	lut_sub lut_1941 ({g91, g176}, g185);
	defparam lut_1941.LUT_SIZE = 2;
	defparam lut_1941.mask = 4'b1000;

	lut_sub lut_1947 ({g36, g176}, g186);
	defparam lut_1947.LUT_SIZE = 2;
	defparam lut_1947.mask = 4'b0010;

	lut_sub lut_1953 ({g88, g176}, g187);
	defparam lut_1953.LUT_SIZE = 2;
	defparam lut_1953.mask = 4'b0010;

	lut_sub lut_1959 ({g3, g174}, g188);
	defparam lut_1959.LUT_SIZE = 2;
	defparam lut_1959.mask = 4'b0010;

	lut_sub lut_1968 ({i_8_, g73, g179, g188, g175, g180}, g189);
	defparam lut_1968.LUT_SIZE = 6;
	defparam lut_1968.mask = 64'h00007fff00000000;

	lut_sub lut_1991 ({g75, g185, g186, g187, g189}, g190);
	defparam lut_1991.LUT_SIZE = 5;
	defparam lut_1991.mask = 32'h8000aaaa;

	lut_sub lut_2005 ({g86, g174}, g191);
	defparam lut_2005.LUT_SIZE = 2;
	defparam lut_2005.mask = 4'b0010;

	lut_sub lut_2011 ({g35, g174}, g192);
	defparam lut_2011.LUT_SIZE = 2;
	defparam lut_2011.mask = 4'b0010;

	lut_sub lut_2020 ({g74, g191, g186, g187, g192}, g193);
	defparam lut_2020.LUT_SIZE = 5;
	defparam lut_2020.mask = 32'h00007fff;

	lut_sub lut_2040 ({g69, g176}, g194);
	defparam lut_2040.LUT_SIZE = 2;
	defparam lut_2040.mask = 4'b0010;

	lut_sub lut_2049 ({g75, g194, g188, g182, g183}, g195);
	defparam lut_2049.LUT_SIZE = 5;
	defparam lut_2049.mask = 32'h7fff0000;

	lut_sub lut_2073 ({g178, g181, g184, g190, g193, g195}, g196);
	defparam lut_2073.LUT_SIZE = 6;
	defparam lut_2073.mask = 64'h0800000000000000;

	lut_sub lut_2079 ({g113, g176}, g197);
	defparam lut_2079.LUT_SIZE = 2;
	defparam lut_2079.mask = 4'b1000;

	lut_sub lut_2086 ({g123, g194, g188}, g198);
	defparam lut_2086.LUT_SIZE = 3;
	defparam lut_2086.mask = 8'h70;

	lut_sub lut_2095 ({g105, g119, g188}, g199);
	defparam lut_2095.LUT_SIZE = 3;
	defparam lut_2095.mask = 8'h51;

	lut_sub lut_2103 ({g126, g174}, g200);
	defparam lut_2103.LUT_SIZE = 2;
	defparam lut_2103.mask = 4'b1000;

	lut_sub lut_2112 ({g125, g122, g123, g197, g200}, g201);
	defparam lut_2112.LUT_SIZE = 5;
	defparam lut_2112.mask = 32'hcf888888;

	lut_sub lut_2132 ({g121, g194, g198, g199, g201}, g202);
	defparam lut_2132.LUT_SIZE = 5;
	defparam lut_2132.mask = 32'h40404000;

	lut_sub lut_2144 ({g75, g164, g122, g194, g197, g202}, g203);
	defparam lut_2144.LUT_SIZE = 6;
	defparam lut_2144.mask = 64'h4440444055504440;

	lut_sub lut_2167 ({g125, g131, g185, g186, g192}, g204);
	defparam lut_2167.LUT_SIZE = 5;
	defparam lut_2167.mask = 32'h88ff80f0;

	lut_sub lut_2188 ({g125, g194, g188}, g205);
	defparam lut_2188.LUT_SIZE = 3;
	defparam lut_2188.mask = 8'h07;

	lut_sub lut_2197 ({g131, g191, g187}, g206);
	defparam lut_2197.LUT_SIZE = 3;
	defparam lut_2197.mask = 8'h70;

	lut_sub lut_2206 ({g125, g175, g177}, g207);
	defparam lut_2206.LUT_SIZE = 3;
	defparam lut_2206.mask = 8'h07;

	lut_sub lut_2215 ({g131, g179, g177}, g208);
	defparam lut_2215.LUT_SIZE = 3;
	defparam lut_2215.mask = 8'h70;

	lut_sub lut_2226 ({g125, g179, g186, g187, g182}, g209);
	defparam lut_2226.LUT_SIZE = 5;
	defparam lut_2226.mask = 32'h00007fff;

	lut_sub lut_2249 ({g205, g206, g207, g208, g209}, g210);
	defparam lut_2249.LUT_SIZE = 5;
	defparam lut_2249.mask = 32'h80000000;

	lut_sub lut_2258 ({g131, g182, g183, g204, g210}, g211);
	defparam lut_2258.LUT_SIZE = 5;
	defparam lut_2258.mask = 32'h10001111;

	lut_sub lut_2268 ({g107, g174}, g212);
	defparam lut_2268.LUT_SIZE = 2;
	defparam lut_2268.mask = 4'b1000;

	lut_sub lut_2274 ({g45, g118}, g213);
	defparam lut_2274.LUT_SIZE = 2;
	defparam lut_2274.mask = 4'b0001;

	lut_sub lut_2281 ({g135, g159, g183}, g214);
	defparam lut_2281.LUT_SIZE = 3;
	defparam lut_2281.mask = 8'h54;

	lut_sub lut_2291 ({g75, g105, g191, g180}, g215);
	defparam lut_2291.LUT_SIZE = 4;
	defparam lut_2291.mask = 16'h7350;

	lut_sub lut_2307 ({g131, g194, g212, g213, g214, g215}, g216);
	defparam lut_2307.LUT_SIZE = 6;
	defparam lut_2307.mask = 64'h8800800088888080;

	lut_sub lut_2321 ({g10, g120}, g217);
	defparam lut_2321.LUT_SIZE = 2;
	defparam lut_2321.mask = 4'b0001;

	lut_sub lut_2326 ({i_8_, i_6_, g120}, g218);
	defparam lut_2326.LUT_SIZE = 3;
	defparam lut_2326.mask = 8'h04;

	lut_sub lut_2331 ({i_10_, i_11_, i_15_, g174}, g219);
	defparam lut_2331.LUT_SIZE = 4;
	defparam lut_2331.mask = 16'h0008;

	lut_sub lut_2341 ({g165, g217, g200, g212, g218, g219}, g220);
	defparam lut_2341.LUT_SIZE = 6;
	defparam lut_2341.mask = 64'h0011151515151515;

	lut_sub lut_2366 ({g165, g179}, g221);
	defparam lut_2366.LUT_SIZE = 2;
	defparam lut_2366.mask = 4'b0001;

	lut_sub lut_2373 ({g122, g175, g177}, g222);
	defparam lut_2373.LUT_SIZE = 3;
	defparam lut_2373.mask = 8'h07;

	lut_sub lut_2383 ({g135, g122, g180, g183}, g223);
	defparam lut_2383.LUT_SIZE = 4;
	defparam lut_2383.mask = 16'hc8f8;

	lut_sub lut_2400 ({g135, g122, g185, g191, g186, g187}, g224);
	defparam lut_2400.LUT_SIZE = 6;
	defparam lut_2400.mask = 64'h80808000ffffcc00;

	lut_sub lut_2428 ({g120, g101}, g225);
	defparam lut_2428.LUT_SIZE = 2;
	defparam lut_2428.mask = 4'b0001;

	lut_sub lut_2434 ({i_8_, g45, g118}, g226);
	defparam lut_2434.LUT_SIZE = 3;
	defparam lut_2434.mask = 8'hfe;

	lut_sub lut_2446 ({g101, g118}, g227);
	defparam lut_2446.LUT_SIZE = 2;
	defparam lut_2446.mask = 4'b0001;

	lut_sub lut_2454 ({g179, g225, g226, g227}, g228);
	defparam lut_2454.LUT_SIZE = 4;
	defparam lut_2454.mask = 16'h00df;

	lut_sub lut_2469 ({g221, g222, g223, g224, g228}, g229);
	defparam lut_2469.LUT_SIZE = 5;
	defparam lut_2469.mask = 32'h02000000;

	lut_sub lut_2477 ({g123, g192, g200, g212}, g230);
	defparam lut_2477.LUT_SIZE = 4;
	defparam lut_2477.mask = 16'h7f00;

	lut_sub lut_2490 ({g122, g123, g191}, g231);
	defparam lut_2490.LUT_SIZE = 3;
	defparam lut_2490.mask = 8'h45;

	lut_sub lut_2499 ({g161, g122, g187}, g232);
	defparam lut_2499.LUT_SIZE = 3;
	defparam lut_2499.mask = 8'h15;

	lut_sub lut_2509 ({g105, g191, g175, g200}, g233);
	defparam lut_2509.LUT_SIZE = 4;
	defparam lut_2509.mask = 16'h7f00;

	lut_sub lut_2524 ({g142, g130, g180, g182, g183}, g234);
	defparam lut_2524.LUT_SIZE = 5;
	defparam lut_2524.mask = 32'h80a088ff;

	lut_sub lut_2545 ({g230, g231, g232, g233, g234}, g235);
	defparam lut_2545.LUT_SIZE = 5;
	defparam lut_2545.mask = 32'h40000000;

	lut_sub lut_2551 ({g102, g212}, g236);
	defparam lut_2551.LUT_SIZE = 2;
	defparam lut_2551.mask = 4'b0001;

	lut_sub lut_2558 ({g102, g182, g183}, g237);
	defparam lut_2558.LUT_SIZE = 3;
	defparam lut_2558.mask = 8'h07;

	lut_sub lut_2567 ({g102, g175, g177}, g238);
	defparam lut_2567.LUT_SIZE = 3;
	defparam lut_2567.mask = 8'h07;

	lut_sub lut_2576 ({g130, g185, g212}, g239);
	defparam lut_2576.LUT_SIZE = 3;
	defparam lut_2576.mask = 8'h70;

	lut_sub lut_2586 ({g102, g105, g183, g192}, g240);
	defparam lut_2586.LUT_SIZE = 4;
	defparam lut_2586.mask = 16'h8f8a;

	lut_sub lut_2601 ({g102, g191, g180, g200}, g241);
	defparam lut_2601.LUT_SIZE = 4;
	defparam lut_2601.mask = 16'h007f;

	lut_sub lut_2617 ({g236, g237, g238, g239, g240, g241}, g242);
	defparam lut_2617.LUT_SIZE = 6;
	defparam lut_2617.mask = 64'h2000000000000000;

	lut_sub lut_2624 ({g130, g191, g187}, g243);
	defparam lut_2624.LUT_SIZE = 3;
	defparam lut_2624.mask = 8'h70;

	lut_sub lut_2633 ({g130, g186, g192}, g244);
	defparam lut_2633.LUT_SIZE = 3;
	defparam lut_2633.mask = 8'h70;

	lut_sub lut_2642 ({g123, g175, g177}, g245);
	defparam lut_2642.LUT_SIZE = 3;
	defparam lut_2642.mask = 8'h70;

	lut_sub lut_2651 ({i_8_, g73, g200, g212}, g246);
	defparam lut_2651.LUT_SIZE = 4;
	defparam lut_2651.mask = 16'h0703;

	lut_sub lut_2664 ({i_8_, g73, g135, g131, g185, g197}, g247);
	defparam lut_2664.LUT_SIZE = 6;
	defparam lut_2664.mask = 64'h8c8f8c8c8c8f8c8f;

	lut_sub lut_2702 ({g243, g244, g245, g246, g247}, g248);
	defparam lut_2702.LUT_SIZE = 5;
	defparam lut_2702.mask = 32'h40000000;

	lut_sub lut_2707 ({i_9_, i_11_, i_15_, g174}, g249);
	defparam lut_2707.LUT_SIZE = 4;
	defparam lut_2707.mask = 16'h8000;

	lut_sub lut_2717 ({g161, g157, g186, g187, g182, g192}, g250);
	defparam lut_2717.LUT_SIZE = 6;
	defparam lut_2717.mask = 64'hfffff0f088008000;

	lut_sub lut_2753 ({g102, g130, g188, g175, g249, g250}, g251);
	defparam lut_2753.LUT_SIZE = 6;
	defparam lut_2753.mask = 64'h5454555544445544;

	lut_sub lut_2786 ({g220, g229, g235, g242, g248, g251}, g252);
	defparam lut_2786.LUT_SIZE = 6;
	defparam lut_2786.mask = 64'h0000000100000000;

	lut_sub lut_2792 ({g2, g120}, g253);
	defparam lut_2792.LUT_SIZE = 2;
	defparam lut_2792.mask = 4'b1110;

	lut_sub lut_2800 ({g30, g166}, g254);
	defparam lut_2800.LUT_SIZE = 2;
	defparam lut_2800.mask = 4'b1110;

	lut_sub lut_2811 ({g157, g165, g182, g253, g254}, g255);
	defparam lut_2811.LUT_SIZE = 5;
	defparam lut_2811.mask = 32'h0e0f0f0f;

	lut_sub lut_2833 ({g80, i_11_, i_15_, g157, g121, g174}, g256);
	defparam lut_2833.LUT_SIZE = 6;
	defparam lut_2833.mask = 64'h0000000022000a00;

	lut_sub lut_2842 ({g2, g166}, g257);
	defparam lut_2842.LUT_SIZE = 2;
	defparam lut_2842.mask = 4'b0001;

	lut_sub lut_2849 ({i_8_, g73, g135, g257}, g258);
	defparam lut_2849.LUT_SIZE = 4;
	defparam lut_2849.mask = 16'h2022;

	lut_sub lut_2857 ({g164, g217}, g259);
	defparam lut_2857.LUT_SIZE = 2;
	defparam lut_2857.mask = 4'b1000;

	lut_sub lut_2862 ({i_9_, i_11_, i_15_, g176}, g260);
	defparam lut_2862.LUT_SIZE = 4;
	defparam lut_2862.mask = 16'h2000;

	lut_sub lut_2872 ({g74, g194, g258, g177, g259, g260}, g261);
	defparam lut_2872.LUT_SIZE = 6;
	defparam lut_2872.mask = 64'h4500454455005544;

	lut_sub lut_2894 ({i_8_, i_6_, i_7_, g120}, g262);
	defparam lut_2894.LUT_SIZE = 4;
	defparam lut_2894.mask = 16'h4010;

	lut_sub lut_2903 ({g159, g185, g262, g191}, g263);
	defparam lut_2903.LUT_SIZE = 4;
	defparam lut_2903.mask = 16'h5703;

	lut_sub lut_2917 ({g165, g154, g192, g263}, g264);
	defparam lut_2917.LUT_SIZE = 4;
	defparam lut_2917.mask = 16'h8a88;

	lut_sub lut_2928 ({g144, g130, g200}, g265);
	defparam lut_2928.LUT_SIZE = 3;
	defparam lut_2928.mask = 8'hb0;

	lut_sub lut_2936 ({i_9_, i_10_, i_11_, i_15_, g130, g174}, g266);
	defparam lut_2936.LUT_SIZE = 6;
	defparam lut_2936.mask = 64'h00000080a0000000;

	lut_sub lut_2947 ({g159, g197, g258, g265, g266}, g267);
	defparam lut_2947.LUT_SIZE = 5;
	defparam lut_2947.mask = 32'hbb00bb0b;

	lut_sub lut_2970 ({g255, g256, g261, g264, g267}, g268);
	defparam lut_2970.LUT_SIZE = 5;
	defparam lut_2970.mask = 32'h10000000;

	lut_sub lut_2980 ({g196, g203, g211, g216, g252, g268}, g269);
	defparam lut_2980.LUT_SIZE = 6;
	defparam lut_2980.mask = 64'h0000000000000001;

	lut_sub lut_2986 ({g3, g24}, g270);
	defparam lut_2986.LUT_SIZE = 2;
	defparam lut_2986.mask = 4'b0010;

	lut_sub lut_2992 ({i_9_, i_10_, i_11_, i_15_, g68, g74}, g271);
	defparam lut_2992.LUT_SIZE = 6;
	defparam lut_2992.mask = 64'h4040400000004040;

	lut_sub lut_3002 ({g24, g86}, g272);
	defparam lut_3002.LUT_SIZE = 2;
	defparam lut_3002.mask = 4'b0100;

	lut_sub lut_3008 ({g68, g86}, g273);
	defparam lut_3008.LUT_SIZE = 2;
	defparam lut_3008.mask = 4'b0100;

	lut_sub lut_3015 ({i_8_, g73, g272, g273}, g274);
	defparam lut_3015.LUT_SIZE = 4;
	defparam lut_3015.mask = 16'h0700;

	lut_sub lut_3023 ({g27, g68}, g275);
	defparam lut_3023.LUT_SIZE = 2;
	defparam lut_3023.mask = 4'b0010;

	lut_sub lut_3030 ({i_8_, g28, g73, g275}, g276);
	defparam lut_3030.LUT_SIZE = 4;
	defparam lut_3030.mask = 16'h0013;

	lut_sub lut_3039 ({i_8_, g28, g73, g275}, g277);
	defparam lut_3039.LUT_SIZE = 4;
	defparam lut_3039.mask = 16'h1300;

	lut_sub lut_3047 ({g20, g68}, g278);
	defparam lut_3047.LUT_SIZE = 2;
	defparam lut_3047.mask = 4'b0010;

	lut_sub lut_3054 ({i_8_, g25, g73, g278}, g279);
	defparam lut_3054.LUT_SIZE = 4;
	defparam lut_3054.mask = 16'h3031;

	lut_sub lut_3066 ({i_8_, g24, g73, g68, g83}, g280);
	defparam lut_3066.LUT_SIZE = 5;
	defparam lut_3066.mask = 32'h05000504;

	lut_sub lut_3076 ({g35, g68}, g281);
	defparam lut_3076.LUT_SIZE = 2;
	defparam lut_3076.mask = 4'b0010;

	lut_sub lut_3082 ({g3, g68}, g282);
	defparam lut_3082.LUT_SIZE = 2;
	defparam lut_3082.mask = 4'b0010;

	lut_sub lut_3091 ({i_8_, g73, g273, g281, g282, g270}, g283);
	defparam lut_3091.LUT_SIZE = 6;
	defparam lut_3091.mask = 64'h0000000000007fff;

	lut_sub lut_3115 ({g274, g276, g277, g279, g280, g283}, g284);
	defparam lut_3115.LUT_SIZE = 6;
	defparam lut_3115.mask = 64'h8000000000000000;

	lut_sub lut_3123 ({g74, g270, g271, g284}, g285);
	defparam lut_3123.LUT_SIZE = 4;
	defparam lut_3123.mask = 16'h4440;

	lut_sub lut_3131 ({g68, g126}, g286);
	defparam lut_3131.LUT_SIZE = 2;
	defparam lut_3131.mask = 4'b1000;

	lut_sub lut_3138 ({g121, g254, g282}, g287);
	defparam lut_3138.LUT_SIZE = 3;
	defparam lut_3138.mask = 8'h45;

	lut_sub lut_3149 ({g3, g24, g68, g125, g126}, g288);
	defparam lut_3149.LUT_SIZE = 5;
	defparam lut_3149.mask = 32'h22203230;

	lut_sub lut_3165 ({g123, g119, g226, g282, g270}, g289);
	defparam lut_3165.LUT_SIZE = 5;
	defparam lut_3165.mask = 32'h8a88cf88;

	lut_sub lut_3187 ({g75, g122, g286, g287, g288, g289}, g290);
	defparam lut_3187.LUT_SIZE = 6;
	defparam lut_3187.mask = 64'h4000400040404000;

	lut_sub lut_3198 ({i_8_, g73, g105, g272}, g291);
	defparam lut_3198.LUT_SIZE = 4;
	defparam lut_3198.mask = 16'h4445;

	lut_sub lut_3210 ({g142, g227, g275, g282}, g292);
	defparam lut_3210.LUT_SIZE = 4;
	defparam lut_3210.mask = 16'hc8f8;

	lut_sub lut_3225 ({i_8_, g24, g73, g126, g105}, g293);
	defparam lut_3225.LUT_SIZE = 5;
	defparam lut_3225.mask = 32'h88008c00;

	lut_sub lut_3236 ({g25, g28, g105}, g294);
	defparam lut_3236.LUT_SIZE = 3;
	defparam lut_3236.mask = 8'ha2;

	lut_sub lut_3244 ({g68, g83}, g295);
	defparam lut_3244.LUT_SIZE = 2;
	defparam lut_3244.mask = 4'b0100;

	lut_sub lut_3250 ({g107, g68}, g296);
	defparam lut_3250.LUT_SIZE = 2;
	defparam lut_3250.mask = 4'b1000;

	lut_sub lut_3259 ({g125, g142, g295, g296, g278}, g297);
	defparam lut_3259.LUT_SIZE = 5;
	defparam lut_3259.mask = 32'ha0ff80c0;

	lut_sub lut_3280 ({g291, g292, g293, g294, g297}, g298);
	defparam lut_3280.LUT_SIZE = 5;
	defparam lut_3280.mask = 32'h00400000;

	lut_sub lut_3288 ({g24, g68, g122, g83}, g299);
	defparam lut_3288.LUT_SIZE = 4;
	defparam lut_3288.mask = 16'h1110;

	lut_sub lut_3298 ({i_8_, g24, g73, g68, g126}, g300);
	defparam lut_3298.LUT_SIZE = 5;
	defparam lut_3298.mask = 32'h0a080000;

	lut_sub lut_3308 ({g28, g135, g122, g275}, g301);
	defparam lut_3308.LUT_SIZE = 4;
	defparam lut_3308.mask = 16'hae0c;

	lut_sub lut_3324 ({g135, g122, g273, g281, g296, g278}, g302);
	defparam lut_3324.LUT_SIZE = 6;
	defparam lut_3324.mask = 64'hc0008000ffffaa00;

	lut_sub lut_3355 ({g24, g35, g107, g123, g130}, g303);
	defparam lut_3355.LUT_SIZE = 5;
	defparam lut_3355.mask = 32'he0ee0000;

	lut_sub lut_3372 ({g299, g300, g301, g302, g303}, g304);
	defparam lut_3372.LUT_SIZE = 5;
	defparam lut_3372.mask = 32'h02000000;

	lut_sub lut_3379 ({g25, g102, g278}, g305);
	defparam lut_3379.LUT_SIZE = 3;
	defparam lut_3379.mask = 8'h31;

	lut_sub lut_3387 ({g225, g275}, g306);
	defparam lut_3387.LUT_SIZE = 2;
	defparam lut_3387.mask = 4'b0001;

	lut_sub lut_3396 ({g24, g35, g102, g83, g105}, g307);
	defparam lut_3396.LUT_SIZE = 5;
	defparam lut_3396.mask = 32'h22af0000;

	lut_sub lut_3412 ({g24, g27, g68, g102, g83}, g308);
	defparam lut_3412.LUT_SIZE = 5;
	defparam lut_3412.mask = 32'h11331010;

	lut_sub lut_3425 ({g24, g107}, g309);
	defparam lut_3425.LUT_SIZE = 2;
	defparam lut_3425.mask = 4'b1000;

	lut_sub lut_3432 ({g102, g272, g309}, g310);
	defparam lut_3432.LUT_SIZE = 3;
	defparam lut_3432.mask = 8'h07;

	lut_sub lut_3441 ({i_8_, g73, g309, g296}, g311);
	defparam lut_3441.LUT_SIZE = 4;
	defparam lut_3441.mask = 16'h0305;

	lut_sub lut_3454 ({g305, g306, g307, g308, g310, g311}, g312);
	defparam lut_3454.LUT_SIZE = 6;
	defparam lut_3454.mask = 64'h8000000000000000;

	lut_sub lut_3460 ({g43, g166}, g313);
	defparam lut_3460.LUT_SIZE = 2;
	defparam lut_3460.mask = 4'b0001;

	lut_sub lut_3467 ({g24, g83, g130}, g314);
	defparam lut_3467.LUT_SIZE = 3;
	defparam lut_3467.mask = 8'h20;

	lut_sub lut_3472 ({i_15_, g24}, g315);
	defparam lut_3472.LUT_SIZE = 2;
	defparam lut_3472.mask = 4'b1000;

	lut_sub lut_3482 ({g151, g313, g278, g314, g315, g1632}, g316);
	defparam lut_3482.LUT_SIZE = 6;
	defparam lut_3482.mask = 64'h5050500040404000;

	lut_sub lut_3497 ({g131, g272, g273}, g317);
	defparam lut_3497.LUT_SIZE = 3;
	defparam lut_3497.mask = 8'h70;

	lut_sub lut_3506 ({g25, g125, g278}, g318);
	defparam lut_3506.LUT_SIZE = 3;
	defparam lut_3506.mask = 8'h31;

	lut_sub lut_3516 ({g131, g295, g281, g296}, g319);
	defparam lut_3516.LUT_SIZE = 4;
	defparam lut_3516.mask = 16'h7f00;

	lut_sub lut_3530 ({g125, g275, g273, g281}, g320);
	defparam lut_3530.LUT_SIZE = 4;
	defparam lut_3530.mask = 16'h007f;

	lut_sub lut_3545 ({g317, g318, g1625, g319, g320}, g321);
	defparam lut_3545.LUT_SIZE = 5;
	defparam lut_3545.mask = 32'h08000000;

	lut_sub lut_3555 ({g290, g298, g304, g312, g316, g321}, g322);
	defparam lut_3555.LUT_SIZE = 6;
	defparam lut_3555.mask = 64'h0000000000000001;

	lut_sub lut_3560 ({i_10_, i_11_, i_15_, g24}, g323);
	defparam lut_3560.LUT_SIZE = 4;
	defparam lut_3560.mask = 16'hfff7;

	lut_sub lut_3578 ({i_8_, i_9_, i_10_, i_11_, i_15_}, g324);
	defparam lut_3578.LUT_SIZE = 5;
	defparam lut_3578.mask = 32'h20000008;

	lut_sub lut_3586 ({g68, g165, g324}, g325);
	defparam lut_3586.LUT_SIZE = 3;
	defparam lut_3586.mask = 8'h10;

	lut_sub lut_3591 ({i_9_, i_10_, i_11_, i_15_, g68}, g326);
	defparam lut_3591.LUT_SIZE = 5;
	defparam lut_3591.mask = 32'h00880800;

	lut_sub lut_3601 ({i_8_, g24, g35, g73, g107}, g327);
	defparam lut_3601.LUT_SIZE = 5;
	defparam lut_3601.mask = 32'h00002300;

	lut_sub lut_3612 ({g125, g105, g272, g326, g327}, g328);
	defparam lut_3612.LUT_SIZE = 5;
	defparam lut_3612.mask = 32'h88aa80a0;

	lut_sub lut_3630 ({g25, g102, g123, g275, g325, g328}, g329);
	defparam lut_3630.LUT_SIZE = 6;
	defparam lut_3630.mask = 64'h0044004044444040;

	lut_sub lut_3647 ({g24, g35, g157, g74, g155}, g330);
	defparam lut_3647.LUT_SIZE = 5;
	defparam lut_3647.mask = 32'h00bf0000;

	lut_sub lut_3663 ({g125, g168, g121, g270, g330, g1606}, g331);
	defparam lut_3663.LUT_SIZE = 6;
	defparam lut_3663.mask = 64'h4440404040404040;

	lut_sub lut_3680 ({g285, g322, g1613, g329, g331}, g332);
	defparam lut_3680.LUT_SIZE = 5;
	defparam lut_3680.mask = 32'h00000001;

	lut_sub lut_3685 ({i_12_, i_13_, i_14_, g20}, g333);
	defparam lut_3685.LUT_SIZE = 4;
	defparam lut_3685.mask = 16'h1101;

	lut_sub lut_3694 ({g28, g98, g180}, g334);
	defparam lut_3694.LUT_SIZE = 3;
	defparam lut_3694.mask = 8'h80;

	lut_sub lut_3699 ({i_12_, i_13_, i_14_, g83}, g335);
	defparam lut_3699.LUT_SIZE = 4;
	defparam lut_3699.mask = 16'h1101;

	lut_sub lut_3708 ({g87, g191, g272}, g336);
	defparam lut_3708.LUT_SIZE = 3;
	defparam lut_3708.mask = 8'h08;

	lut_sub lut_3714 ({g35, g176}, g337);
	defparam lut_3714.LUT_SIZE = 2;
	defparam lut_3714.mask = 4'b0010;

	lut_sub lut_3719 ({i_12_, i_13_, i_14_, g107}, g338);
	defparam lut_3719.LUT_SIZE = 4;
	defparam lut_3719.mask = 16'h2202;

	lut_sub lut_3726 ({i_12_, i_13_, i_14_, g35}, g339);
	defparam lut_3726.LUT_SIZE = 4;
	defparam lut_3726.mask = 16'h1101;

	lut_sub lut_3734 ({g83, g176}, g340);
	defparam lut_3734.LUT_SIZE = 2;
	defparam lut_3734.mask = 4'b1101;

	lut_sub lut_3743 ({g77, g188, g270}, g341);
	defparam lut_3743.LUT_SIZE = 3;
	defparam lut_3743.mask = 8'h80;

	lut_sub lut_3749 ({g86, g176}, g342);
	defparam lut_3749.LUT_SIZE = 2;
	defparam lut_3749.mask = 4'b0010;

	lut_sub lut_3755 ({g20, g176}, g343);
	defparam lut_3755.LUT_SIZE = 2;
	defparam lut_3755.mask = 4'b1101;

	lut_sub lut_3766 ({g164, g340, g341, g342, g343}, g344);
	defparam lut_3766.LUT_SIZE = 5;
	defparam lut_3766.mask = 32'h0000fffb;

	lut_sub lut_3790 ({g164, g253, g337, g338, g339, g344}, g345);
	defparam lut_3790.LUT_SIZE = 6;
	defparam lut_3790.mask = 64'h8800aaaa80008080;

	lut_sub lut_3812 ({g253, g333, g334, g335, g336, g345}, g346);
	defparam lut_3812.LUT_SIZE = 6;
	defparam lut_3812.mask = 64'h0010000055555555;

	lut_sub lut_3834 ({g154, g122}, g347);
	defparam lut_3834.LUT_SIZE = 2;
	defparam lut_3834.mask = 4'b0010;

	lut_sub lut_3840 ({i_8_, g73, g130}, g348);
	defparam lut_3840.LUT_SIZE = 3;
	defparam lut_3840.mask = 8'h45;

	lut_sub lut_3851 ({g144, g164, g347, g105, g348}, g349);
	defparam lut_3851.LUT_SIZE = 5;
	defparam lut_3851.mask = 32'h01000000;

	lut_sub lut_3858 ({i_8_, i_6_, i_7_, g120, g166, g118}, g350);
	defparam lut_3858.LUT_SIZE = 6;
	defparam lut_3858.mask = 64'h330f3300330f5f00;

	lut_sub lut_3889 ({i_7_, g72, g350}, g351);
	defparam lut_3889.LUT_SIZE = 3;
	defparam lut_3889.mask = 8'ha8;

	lut_sub lut_3899 ({g119, g121, g227, g351}, g352);
	defparam lut_3899.LUT_SIZE = 4;
	defparam lut_3899.mask = 16'h4000;

	lut_sub lut_3904 ({i_11_, i_15_, g53}, g353);
	defparam lut_3904.LUT_SIZE = 3;
	defparam lut_3904.mask = 8'h80;

	lut_sub lut_3914 ({g3, g35, g176, g349, g352, g353}, g354);
	defparam lut_3914.LUT_SIZE = 6;
	defparam lut_3914.mask = 64'h4000500044005400;

	lut_sub lut_3925 ({i_12_, i_14_}, g355);
	defparam lut_3925.LUT_SIZE = 2;
	defparam lut_3925.mask = 4'b0100;

	lut_sub lut_3931 ({g159, g313}, g356);
	defparam lut_3931.LUT_SIZE = 2;
	defparam lut_3931.mask = 4'b1101;

	lut_sub lut_3939 ({g27, g176}, g357);
	defparam lut_3939.LUT_SIZE = 2;
	defparam lut_3939.mask = 4'b0010;

	lut_sub lut_3945 ({g107, g176}, g358);
	defparam lut_3945.LUT_SIZE = 2;
	defparam lut_3945.mask = 4'b1000;

	lut_sub lut_3953 ({g27, g126, g102, g176}, g359);
	defparam lut_3953.LUT_SIZE = 4;
	defparam lut_3953.mask = 16'h2022;

	lut_sub lut_3963 ({g105, g342, g358, g359}, g360);
	defparam lut_3963.LUT_SIZE = 4;
	defparam lut_3963.mask = 16'h80aa;

	lut_sub lut_3977 ({g355, g83, g356, g357, g350, g360}, g361);
	defparam lut_3977.LUT_SIZE = 6;
	defparam lut_3977.mask = 64'h5454545454545400;

	lut_sub lut_4004 ({g154, g340, g335}, g362);
	defparam lut_4004.LUT_SIZE = 3;
	defparam lut_4004.mask = 8'hd0;

	lut_sub lut_4014 ({g159, g154, g333, g343}, g363);
	defparam lut_4014.LUT_SIZE = 4;
	defparam lut_4014.mask = 16'h4c4f;

	lut_sub lut_4030 ({g159, g154, g337, g334, g339}, g364);
	defparam lut_4030.LUT_SIZE = 5;
	defparam lut_4030.mask = 32'h202033ff;

	lut_sub lut_4053 ({g154, g342, g336, g362, g363, g364}, g365);
	defparam lut_4053.LUT_SIZE = 6;
	defparam lut_4053.mask = 64'h0010000010101010;

	lut_sub lut_4065 ({g102, g186, g296, g358}, g366);
	defparam lut_4065.LUT_SIZE = 4;
	defparam lut_4065.mask = 16'h007f;

	lut_sub lut_4079 ({g108, g105, g212, g309}, g367);
	defparam lut_4079.LUT_SIZE = 4;
	defparam lut_4079.mask = 16'h70f0;

	lut_sub lut_4093 ({g123, g185, g187, g337}, g368);
	defparam lut_4093.LUT_SIZE = 4;
	defparam lut_4093.mask = 16'h7f00;

	lut_sub lut_4104 ({i_12_, i_13_, i_14_, g126}, g369);
	defparam lut_4104.LUT_SIZE = 4;
	defparam lut_4104.mask = 16'h2202;

	lut_sub lut_4114 ({g253, g369, g338, g358}, g370);
	defparam lut_4114.LUT_SIZE = 4;
	defparam lut_4114.mask = 16'h7f00;

	lut_sub lut_4128 ({g135, g122, g131, g342}, g371);
	defparam lut_4128.LUT_SIZE = 4;
	defparam lut_4128.mask = 16'h5545;

	lut_sub lut_4142 ({g123, g130, g342, g358}, g372);
	defparam lut_4142.LUT_SIZE = 4;
	defparam lut_4142.mask = 16'h8c8f;

	lut_sub lut_4158 ({g367, g368, g370, g371, g372}, g373);
	defparam lut_4158.LUT_SIZE = 5;
	defparam lut_4158.mask = 32'h40000000;

	lut_sub lut_4166 ({g161, g157, g337, g343}, g374);
	defparam lut_4166.LUT_SIZE = 4;
	defparam lut_4166.mask = 16'hfc44;

	lut_sub lut_4180 ({i_8_, g73, g192, g212}, g375);
	defparam lut_4180.LUT_SIZE = 4;
	defparam lut_4180.mask = 16'h0007;

	lut_sub lut_4190 ({g125, g191, g192, g212}, g376);
	defparam lut_4190.LUT_SIZE = 4;
	defparam lut_4190.mask = 16'h007f;

	lut_sub lut_4203 ({i_8_, g73, g102, g337}, g377);
	defparam lut_4203.LUT_SIZE = 4;
	defparam lut_4203.mask = 16'h1115;

	lut_sub lut_4217 ({g102, g105, g186, g182, g295, g281}, g378);
	defparam lut_4217.LUT_SIZE = 6;
	defparam lut_4217.mask = 64'h8000ffff8000aaaa;

	lut_sub lut_4251 ({g374, g375, g376, g377, g378}, g379);
	defparam lut_4251.LUT_SIZE = 5;
	defparam lut_4251.mask = 32'h00004000;

	lut_sub lut_4259 ({g164, g123, g333, g335}, g380);
	defparam lut_4259.LUT_SIZE = 4;
	defparam lut_4259.mask = 16'haf88;

	lut_sub lut_4275 ({g226, g227, g275, g357, g334}, g381);
	defparam lut_4275.LUT_SIZE = 5;
	defparam lut_4275.mask = 32'h5040ff44;

	lut_sub lut_4297 ({g164, g225, g334, g336, g380, g381}, g382);
	defparam lut_4297.LUT_SIZE = 6;
	defparam lut_4297.mask = 64'h1111001100010001;

	lut_sub lut_4310 ({g125, g254}, g383);
	defparam lut_4310.LUT_SIZE = 2;
	defparam lut_4310.mask = 4'b0100;

	lut_sub lut_4319 ({g142, g257, g179, g254, g217}, g384);
	defparam lut_4319.LUT_SIZE = 5;
	defparam lut_4319.mask = 32'h0f0f0d0f;

	lut_sub lut_4340 ({i_8_, g73, g357, g358}, g385);
	defparam lut_4340.LUT_SIZE = 4;
	defparam lut_4340.mask = 16'h0507;

	lut_sub lut_4354 ({g347, g356, g383, g384, g358, g385}, g386);
	defparam lut_4354.LUT_SIZE = 6;
	defparam lut_4354.mask = 64'h8080808080a08080;

	lut_sub lut_4372 ({g365, g366, g373, g379, g382, g386}, g387);
	defparam lut_4372.LUT_SIZE = 6;
	defparam lut_4372.mask = 64'h0000000000010000;

	lut_sub lut_4379 ({i_12_, i_13_, i_14_, g20, g157, g130}, g388);
	defparam lut_4379.LUT_SIZE = 6;
	defparam lut_4379.mask = 64'h0000000a00030000;

	lut_sub lut_4390 ({g3, g176, g226, g341}, g389);
	defparam lut_4390.LUT_SIZE = 4;
	defparam lut_4390.mask = 16'h88c8;

	lut_sub lut_4404 ({g20, g126, g122, g123, g105, g176}, g390);
	defparam lut_4404.LUT_SIZE = 6;
	defparam lut_4404.mask = 64'ha8a80000a8aa88aa;

	lut_sub lut_4431 ({g125, g126, g176, g389, g390}, g391);
	defparam lut_4431.LUT_SIZE = 5;
	defparam lut_4431.mask = 32'h88880888;

	lut_sub lut_4443 ({g42, g72}, g392);
	defparam lut_4443.LUT_SIZE = 2;
	defparam lut_4443.mask = 4'b0001;

	lut_sub lut_4451 ({g102, g191, g273, g392}, g393);
	defparam lut_4451.LUT_SIZE = 4;
	defparam lut_4451.mask = 16'h0537;

	lut_sub lut_4463 ({g15, g71}, g394);
	defparam lut_4463.LUT_SIZE = 2;
	defparam lut_4463.mask = 4'b0001;

	lut_sub lut_4468 ({i_6_, i_7_, i_10_, i_11_, g394}, g395);
	defparam lut_4468.LUT_SIZE = 5;
	defparam lut_4468.mask = 32'h00040400;

	lut_sub lut_4476 ({g142, g333, g395}, g396);
	defparam lut_4476.LUT_SIZE = 3;
	defparam lut_4476.mask = 8'h8a;

	lut_sub lut_4484 ({g355, g126}, g397);
	defparam lut_4484.LUT_SIZE = 2;
	defparam lut_4484.mask = 4'b0010;

	lut_sub lut_4493 ({i_14_, g125, g154, g122, g83, g397}, g398);
	defparam lut_4493.LUT_SIZE = 6;
	defparam lut_4493.mask = 64'h5505550555057737;

	lut_sub lut_4531 ({g135, g123, g186, g227, g341, g337}, g399);
	defparam lut_4531.LUT_SIZE = 6;
	defparam lut_4531.mask = 64'ha200a2a2f300f3f3;

	lut_sub lut_4567 ({g356, g369, g393, g396, g398, g399}, g400);
	defparam lut_4567.LUT_SIZE = 6;
	defparam lut_4567.mask = 64'h0400040004000000;

	lut_sub lut_4577 ({g105, g257, g254, g217}, g401);
	defparam lut_4577.LUT_SIZE = 4;
	defparam lut_4577.mask = 16'h0020;

	lut_sub lut_4586 ({g159, g154, g122, g257, g313}, g402);
	defparam lut_4586.LUT_SIZE = 5;
	defparam lut_4586.mask = 32'h00000080;

	lut_sub lut_4590 ({i_9_, i_10_, i_11_}, g403);
	defparam lut_4590.LUT_SIZE = 3;
	defparam lut_4590.mask = 8'h42;

	lut_sub lut_4600 ({i_15_, g68, g257, g254, g217, g403}, g404);
	defparam lut_4600.LUT_SIZE = 6;
	defparam lut_4600.mask = 64'h5155000000000000;

	lut_sub lut_4615 ({g296, g282, g401, g402, g404}, g405);
	defparam lut_4615.LUT_SIZE = 5;
	defparam lut_4615.mask = 32'haa220a02;

	lut_sub lut_4632 ({g185, g197, g179, g187, g282}, g406);
	defparam lut_4632.LUT_SIZE = 5;
	defparam lut_4632.mask = 32'h80000000;

	lut_sub lut_4638 ({i_8_, i_6_, i_7_, g72, g120}, g407);
	defparam lut_4638.LUT_SIZE = 5;
	defparam lut_4638.mask = 32'h57030350;

	lut_sub lut_4654 ({g1, g118}, g408);
	defparam lut_4654.LUT_SIZE = 2;
	defparam lut_4654.mask = 4'b1110;

	lut_sub lut_4663 ({g272, g334, g408}, g409);
	defparam lut_4663.LUT_SIZE = 3;
	defparam lut_4663.mask = 8'h8a;

	lut_sub lut_4674 ({g168, g342, g406, g407, g409}, g410);
	defparam lut_4674.LUT_SIZE = 5;
	defparam lut_4674.mask = 32'haa880a08;

	lut_sub lut_4691 ({g388, g391, g400, g405, g410}, g411);
	defparam lut_4691.LUT_SIZE = 5;
	defparam lut_4691.mask = 32'h00010000;

	lut_sub lut_4700 ({g346, g354, g361, g387, g411}, g412);
	defparam lut_4700.LUT_SIZE = 5;
	defparam lut_4700.mask = 32'h00000100;

	lut_sub lut_4707 ({g102, g257, g313}, g413);
	defparam lut_4707.LUT_SIZE = 3;
	defparam lut_4707.mask = 8'h80;

	lut_sub lut_4714 ({g105, g119, g413}, g414);
	defparam lut_4714.LUT_SIZE = 3;
	defparam lut_4714.mask = 8'h04;

	lut_sub lut_4721 ({g78, g131, g333}, g415);
	defparam lut_4721.LUT_SIZE = 3;
	defparam lut_4721.mask = 8'hc4;

	lut_sub lut_4728 ({i_9_, i_10_, i_11_, i_15_, g176}, g416);
	defparam lut_4728.LUT_SIZE = 5;
	defparam lut_4728.mask = 32'h00000220;

	lut_sub lut_4737 ({i_6_, g120, g154, g197, g416}, g417);
	defparam lut_4737.LUT_SIZE = 5;
	defparam lut_4737.mask = 32'h30753030;

	lut_sub lut_4756 ({g355, g35, g107, g159, g313}, g418);
	defparam lut_4756.LUT_SIZE = 5;
	defparam lut_4756.mask = 32'h0000d0d5;

	lut_sub lut_4772 ({g20, g355, g135, g165, g174}, g419);
	defparam lut_4772.LUT_SIZE = 5;
	defparam lut_4772.mask = 32'h0000a0b3;

	lut_sub lut_4788 ({g194, g414, g415, g417, g418, g419}, g420);
	defparam lut_4788.LUT_SIZE = 6;
	defparam lut_4788.mask = 64'h8000800000008000;

	lut_sub lut_4796 ({g1, g120}, g421);
	defparam lut_4796.LUT_SIZE = 2;
	defparam lut_4796.mask = 4'b0001;

	lut_sub lut_4803 ({g159, g313, g421}, g422);
	defparam lut_4803.LUT_SIZE = 3;
	defparam lut_4803.mask = 8'hf7;

	lut_sub lut_4816 ({i_15_, g34, g68, g422}, g423);
	defparam lut_4816.LUT_SIZE = 4;
	defparam lut_4816.mask = 16'h0004;

	lut_sub lut_4823 ({g25, g130, g397}, g424);
	defparam lut_4823.LUT_SIZE = 3;
	defparam lut_4823.mask = 8'hc4;

	lut_sub lut_4832 ({g257, g254, g217}, g425);
	defparam lut_4832.LUT_SIZE = 3;
	defparam lut_4832.mask = 8'h20;

	lut_sub lut_4840 ({g92, g105, g275, g425}, g426);
	defparam lut_4840.LUT_SIZE = 4;
	defparam lut_4840.mask = 16'hcd0d;

	lut_sub lut_4856 ({g161, g183, g423, g424, g426}, g427);
	defparam lut_4856.LUT_SIZE = 5;
	defparam lut_4856.mask = 32'h40404000;

	lut_sub lut_4862 ({i_9_, i_10_, i_11_}, g428);
	defparam lut_4862.LUT_SIZE = 3;
	defparam lut_4862.mask = 8'hdf;

	lut_sub lut_4872 ({i_9_, i_10_, i_11_}, g429);
	defparam lut_4872.LUT_SIZE = 3;
	defparam lut_4872.mask = 8'h04;

	lut_sub lut_4879 ({i_15_, g428, g68, g429}, g430);
	defparam lut_4879.LUT_SIZE = 4;
	defparam lut_4879.mask = 16'hc444;

	lut_sub lut_4888 ({i_8_, i_6_, i_7_, g120}, g431);
	defparam lut_4888.LUT_SIZE = 4;
	defparam lut_4888.mask = 16'h1040;

	lut_sub lut_4897 ({g159, g185, g272, g431}, g432);
	defparam lut_4897.LUT_SIZE = 4;
	defparam lut_4897.mask = 16'h3705;

	lut_sub lut_4912 ({g425, g402, g341, g430, g432}, g433);
	defparam lut_4912.LUT_SIZE = 5;
	defparam lut_4912.mask = 32'h08880aaa;

	lut_sub lut_4927 ({i_8_, i_6_, i_7_, g72, g120, g118}, g434);
	defparam lut_4927.LUT_SIZE = 6;
	defparam lut_4927.mask = 64'h005f00330000005f;

	lut_sub lut_4950 ({g154, g253, g356, g383}, g435);
	defparam lut_4950.LUT_SIZE = 4;
	defparam lut_4950.mask = 16'h0004;

	lut_sub lut_4957 ({g164, g213, g402}, g436);
	defparam lut_4957.LUT_SIZE = 3;
	defparam lut_4957.mask = 8'hbf;

	lut_sub lut_4973 ({g70, g82, g357, g434, g435, g436}, g437);
	defparam lut_4973.LUT_SIZE = 6;
	defparam lut_4973.mask = 64'hfff03330aaa02220;

	lut_sub lut_5007 ({g102, g122, g257, g313}, g438);
	defparam lut_5007.LUT_SIZE = 4;
	defparam lut_5007.mask = 16'h8000;

	lut_sub lut_5015 ({g73, g159, g123, g142}, g439);
	defparam lut_5015.LUT_SIZE = 4;
	defparam lut_5015.mask = 16'h0100;

	lut_sub lut_5022 ({g105, g438, g439}, g440);
	defparam lut_5022.LUT_SIZE = 3;
	defparam lut_5022.mask = 8'h01;

	lut_sub lut_5031 ({g413, g217, g286, g340, g440}, g441);
	defparam lut_5031.LUT_SIZE = 5;
	defparam lut_5031.mask = 32'h70707770;

	lut_sub lut_5055 ({g420, g427, g433, g437, g441, g1593}, g442);
	defparam lut_5055.LUT_SIZE = 6;
	defparam lut_5055.mask = 64'h0000000000000001;

	lut_sub lut_5062 ({g73, g164, g402}, g443);
	defparam lut_5062.LUT_SIZE = 3;
	defparam lut_5062.mask = 8'h40;

	lut_sub lut_5069 ({g142, g105, g259}, g444);
	defparam lut_5069.LUT_SIZE = 3;
	defparam lut_5069.mask = 8'h01;

	lut_sub lut_5074 ({g80, i_11_}, g445);
	defparam lut_5074.LUT_SIZE = 2;
	defparam lut_5074.mask = 4'b0001;

	lut_sub lut_5081 ({g125, g413, g439}, g446);
	defparam lut_5081.LUT_SIZE = 3;
	defparam lut_5081.mask = 8'h10;

	lut_sub lut_5087 ({g142, g217}, g447);
	defparam lut_5087.LUT_SIZE = 2;
	defparam lut_5087.mask = 4'b0010;

	lut_sub lut_5096 ({i_15_, g428, g445, g176, g446, g447}, g448);
	defparam lut_5096.LUT_SIZE = 6;
	defparam lut_5096.mask = 64'hc0c0000000a000a0;

	lut_sub lut_5111 ({g78, g177, g278, g333}, g449);
	defparam lut_5111.LUT_SIZE = 4;
	defparam lut_5111.mask = 16'h0080;

	lut_sub lut_5120 ({g24, g35, g36, g161, g68}, g450);
	defparam lut_5120.LUT_SIZE = 5;
	defparam lut_5120.mask = 32'h0aff0a2a;

	lut_sub lut_5141 ({g20, g355, g78}, g451);
	defparam lut_5141.LUT_SIZE = 3;
	defparam lut_5141.mask = 8'h54;

	lut_sub lut_5152 ({g161, g175, g177, g278, g451}, g452);
	defparam lut_5152.LUT_SIZE = 5;
	defparam lut_5152.mask = 32'h0000bfff;

	lut_sub lut_5175 ({g109, g157, g186, g192, g452}, g453);
	defparam lut_5175.LUT_SIZE = 5;
	defparam lut_5175.mask = 32'haa80aa00;

	lut_sub lut_5191 ({i_8_, g392, g449, g450, g453}, g454);
	defparam lut_5191.LUT_SIZE = 5;
	defparam lut_5191.mask = 32'h55055544;

	lut_sub lut_5210 ({g66, g1584, g448, g454}, g455);
	defparam lut_5210.LUT_SIZE = 4;
	defparam lut_5210.mask = 16'h0004;

	lut_sub lut_5220 ({g173, g269, g332, g412, g442, g455}, g456);
	defparam lut_5220.LUT_SIZE = 6;
	defparam lut_5220.mask = 64'h0000000000000001;

	lut_sub lut_5225 ({i_0_, i_1_, g6}, g457);
	defparam lut_5225.LUT_SIZE = 3;
	defparam lut_5225.mask = 8'h04;

	lut_sub lut_5231 ({g457, g51}, g458);
	defparam lut_5231.LUT_SIZE = 2;
	defparam lut_5231.mask = 4'b0100;

	lut_sub lut_5239 ({g24, g74, g91, g257}, g459);
	defparam lut_5239.LUT_SIZE = 4;
	defparam lut_5239.mask = 16'h4c00;

	lut_sub lut_5245 ({i_12_, i_13_, i_14_}, g460);
	defparam lut_5245.LUT_SIZE = 3;
	defparam lut_5245.mask = 8'hfd;

	lut_sub lut_5257 ({g27, g460}, g461);
	defparam lut_5257.LUT_SIZE = 2;
	defparam lut_5257.mask = 4'b0010;

	lut_sub lut_5264 ({g75, g107, g460}, g462);
	defparam lut_5264.LUT_SIZE = 3;
	defparam lut_5264.mask = 8'h80;

	lut_sub lut_5272 ({i_8_, g27, g73, g86, g460}, g463);
	defparam lut_5272.LUT_SIZE = 5;
	defparam lut_5272.mask = 32'h020a000a;

	lut_sub lut_5284 ({i_8_, g3, g73, g83, g460}, g464);
	defparam lut_5284.LUT_SIZE = 5;
	defparam lut_5284.mask = 32'h0202020a;

	lut_sub lut_5296 ({i_8_, g20, g35, g73, g460}, g465);
	defparam lut_5296.LUT_SIZE = 5;
	defparam lut_5296.mask = 32'h00220222;

	lut_sub lut_5308 ({i_8_, g73, g107, g353, g460}, g466);
	defparam lut_5308.LUT_SIZE = 5;
	defparam lut_5308.mask = 32'h00a20000;

	lut_sub lut_5318 ({g463, g464, g465, g466}, g467);
	defparam lut_5318.LUT_SIZE = 4;
	defparam lut_5318.mask = 16'h8000;

	lut_sub lut_5324 ({g24, g69}, g468);
	defparam lut_5324.LUT_SIZE = 2;
	defparam lut_5324.mask = 4'b0100;

	lut_sub lut_5331 ({g3, g460, g468}, g469);
	defparam lut_5331.LUT_SIZE = 3;
	defparam lut_5331.mask = 8'ha2;

	lut_sub lut_5340 ({g121, g213, g469}, g470);
	defparam lut_5340.LUT_SIZE = 3;
	defparam lut_5340.mask = 8'h2a;

	lut_sub lut_5349 ({g161, g86, g460}, g471);
	defparam lut_5349.LUT_SIZE = 3;
	defparam lut_5349.mask = 8'h02;

	lut_sub lut_5357 ({g20, g27, g83, g460}, g472);
	defparam lut_5357.LUT_SIZE = 4;
	defparam lut_5357.mask = 16'h2aaa;

	lut_sub lut_5369 ({g24, g81}, g473);
	defparam lut_5369.LUT_SIZE = 2;
	defparam lut_5369.mask = 4'b0100;

	lut_sub lut_5377 ({g157, g86, g460, g473}, g474);
	defparam lut_5377.LUT_SIZE = 4;
	defparam lut_5377.mask = 16'h005d;

	lut_sub lut_5389 ({i_8_, g73, g86, g126, g460}, g475);
	defparam lut_5389.LUT_SIZE = 5;
	defparam lut_5389.mask = 32'h0088008a;

	lut_sub lut_5403 ({g142, g470, g471, g472, g474, g475}, g476);
	defparam lut_5403.LUT_SIZE = 6;
	defparam lut_5403.mask = 64'h8000000088000000;

	lut_sub lut_5411 ({g17, g24}, g477);
	defparam lut_5411.LUT_SIZE = 2;
	defparam lut_5411.mask = 4'b0010;

	lut_sub lut_5419 ({g80, i_11_, i_15_, g119, g392, g460}, g478);
	defparam lut_5419.LUT_SIZE = 6;
	defparam lut_5419.mask = 64'h000000000a002200;

	lut_sub lut_5430 ({g225, g213, g477, g478}, g479);
	defparam lut_5430.LUT_SIZE = 4;
	defparam lut_5430.mask = 16'ha888;

	lut_sub lut_5444 ({g167, g461, g462, g467, g476, g479}, g480);
	defparam lut_5444.LUT_SIZE = 6;
	defparam lut_5444.mask = 64'h0100010001000000;

	lut_sub lut_5454 ({g24, g154, g91, g175}, g481);
	defparam lut_5454.LUT_SIZE = 4;
	defparam lut_5454.mask = 16'hd050;

	lut_sub lut_5462 ({i_12_, i_13_, i_14_}, g482);
	defparam lut_5462.LUT_SIZE = 3;
	defparam lut_5462.mask = 8'h54;

	lut_sub lut_5470 ({g36, g482}, g483);
	defparam lut_5470.LUT_SIZE = 2;
	defparam lut_5470.mask = 4'b0001;

	lut_sub lut_5476 ({g91, g482}, g484);
	defparam lut_5476.LUT_SIZE = 2;
	defparam lut_5476.mask = 4'b0100;

	lut_sub lut_5484 ({g159, g154, g483, g484}, g485);
	defparam lut_5484.LUT_SIZE = 4;
	defparam lut_5484.mask = 16'h7530;

	lut_sub lut_5496 ({g91, g460}, g486);
	defparam lut_5496.LUT_SIZE = 2;
	defparam lut_5496.mask = 4'b1000;

	lut_sub lut_5502 ({g91, g174}, g487);
	defparam lut_5502.LUT_SIZE = 2;
	defparam lut_5502.mask = 4'b1000;

	lut_sub lut_5510 ({g102, g105, g486, g487}, g488);
	defparam lut_5510.LUT_SIZE = 4;
	defparam lut_5510.mask = 16'h3075;

	lut_sub lut_5522 ({g17, g482}, g489);
	defparam lut_5522.LUT_SIZE = 2;
	defparam lut_5522.mask = 4'b0001;

	lut_sub lut_5532 ({g105, g253, g200, g212, g356, g489}, g490);
	defparam lut_5532.LUT_SIZE = 6;
	defparam lut_5532.mask = 64'ha000a080ff00ffcc;

	lut_sub lut_5564 ({g481, g485, g488, g490}, g491);
	defparam lut_5564.LUT_SIZE = 4;
	defparam lut_5564.mask = 16'h4000;

	lut_sub lut_5572 ({g24, g36, g91, g88}, g492);
	defparam lut_5572.LUT_SIZE = 4;
	defparam lut_5572.mask = 16'hdf00;

	lut_sub lut_5588 ({g165, g131, g257, g383, g477, g492}, g493);
	defparam lut_5588.LUT_SIZE = 6;
	defparam lut_5588.mask = 64'h8888cfcc88888888;

	lut_sub lut_5615 ({i_9_, i_10_, i_11_, i_15_, g174, g460}, g494);
	defparam lut_5615.LUT_SIZE = 6;
	defparam lut_5615.mask = 64'ha0a0aaaea0aaaca0;

	lut_sub lut_5645 ({g22, g460}, g495);
	defparam lut_5645.LUT_SIZE = 2;
	defparam lut_5645.mask = 4'b1000;

	lut_sub lut_5651 ({g24, g88}, g496);
	defparam lut_5651.LUT_SIZE = 2;
	defparam lut_5651.mask = 4'b0100;

	lut_sub lut_5658 ({i_8_, i_6_, i_7_, g118, g495, g496}, g497);
	defparam lut_5658.LUT_SIZE = 6;
	defparam lut_5658.mask = 64'h0502000000000000;

	lut_sub lut_5669 ({g102, g350, g468, g494, g497}, g498);
	defparam lut_5669.LUT_SIZE = 5;
	defparam lut_5669.mask = 32'haa80a080;

	lut_sub lut_5685 ({g459, g480, g491, g493, g498}, g499);
	defparam lut_5685.LUT_SIZE = 5;
	defparam lut_5685.mask = 32'h00010000;

	lut_sub lut_5690 ({i_12_, i_13_, i_14_, g88}, g500);
	defparam lut_5690.LUT_SIZE = 4;
	defparam lut_5690.mask = 16'h1110;

	lut_sub lut_5698 ({g81, g460}, g501);
	defparam lut_5698.LUT_SIZE = 2;
	defparam lut_5698.mask = 4'b0010;

	lut_sub lut_5706 ({g161, g183, g501, g473}, g502);
	defparam lut_5706.LUT_SIZE = 4;
	defparam lut_5706.mask = 16'h007f;

	lut_sub lut_5722 ({g125, g164, g105, g487, g500, g502}, g503);
	defparam lut_5722.LUT_SIZE = 6;
	defparam lut_5722.mask = 64'h88aa888880a08080;

	lut_sub lut_5743 ({g355, g91, g212}, g504);
	defparam lut_5743.LUT_SIZE = 3;
	defparam lut_5743.mask = 8'ha2;

	lut_sub lut_5752 ({g157, g186, g192}, g505);
	defparam lut_5752.LUT_SIZE = 3;
	defparam lut_5752.mask = 8'h07;

	lut_sub lut_5763 ({g125, g253, g483, g504, g505}, g506);
	defparam lut_5763.LUT_SIZE = 5;
	defparam lut_5763.mask = 32'ha0aa2022;

	lut_sub lut_5775 ({i_12_, i_13_, i_14_}, g507);
	defparam lut_5775.LUT_SIZE = 3;
	defparam lut_5775.mask = 8'h14;

	lut_sub lut_5782 ({g69, g507}, g508);
	defparam lut_5782.LUT_SIZE = 2;
	defparam lut_5782.mask = 4'b0001;

	lut_sub lut_5790 ({g355, g125, g88, g191}, g509);
	defparam lut_5790.LUT_SIZE = 4;
	defparam lut_5790.mask = 16'h0507;

	lut_sub lut_5803 ({g122, g413, g473, g508, g509}, g510);
	defparam lut_5803.LUT_SIZE = 5;
	defparam lut_5803.mask = 32'h80aa80a0;

	lut_sub lut_5816 ({g69, g460}, g511);
	defparam lut_5816.LUT_SIZE = 2;
	defparam lut_5816.mask = 4'b0010;

	lut_sub lut_5824 ({g180, g225, g213, g425}, g512);
	defparam lut_5824.LUT_SIZE = 4;
	defparam lut_5824.mask = 16'h00bf;

	lut_sub lut_5836 ({g36, g76}, g513);
	defparam lut_5836.LUT_SIZE = 2;
	defparam lut_5836.mask = 4'b1101;

	lut_sub lut_5844 ({g24, g36}, g514);
	defparam lut_5844.LUT_SIZE = 2;
	defparam lut_5844.mask = 4'b0100;

	lut_sub lut_5852 ({g125, g192, g513, g514}, g515);
	defparam lut_5852.LUT_SIZE = 4;
	defparam lut_5852.mask = 16'h00df;

	lut_sub lut_5867 ({g188, g436, g511, g512, g515}, g516);
	defparam lut_5867.LUT_SIZE = 5;
	defparam lut_5867.mask = 32'h88808800;

	lut_sub lut_5879 ({g24, g113, g257, g356}, g517);
	defparam lut_5879.LUT_SIZE = 4;
	defparam lut_5879.mask = 16'h7000;

	lut_sub lut_5886 ({i_8_, i_6_, i_7_, g120}, g518);
	defparam lut_5886.LUT_SIZE = 4;
	defparam lut_5886.mask = 16'h4050;

	lut_sub lut_5896 ({g348, g514, g517, g1577}, g519);
	defparam lut_5896.LUT_SIZE = 4;
	defparam lut_5896.mask = 16'h4044;

	lut_sub lut_5904 ({i_9_, i_10_, i_11_, g225, g213}, g520);
	defparam lut_5904.LUT_SIZE = 5;
	defparam lut_5904.mask = 32'hffff8fff;

	lut_sub lut_5938 ({g22, g482}, g521);
	defparam lut_5938.LUT_SIZE = 2;
	defparam lut_5938.mask = 4'b0100;

	lut_sub lut_5944 ({g88, g174}, g522);
	defparam lut_5944.LUT_SIZE = 2;
	defparam lut_5944.mask = 4'b0010;

	lut_sub lut_5953 ({g164, g253, g483, g484, g500}, g523);
	defparam lut_5953.LUT_SIZE = 5;
	defparam lut_5953.mask = 32'haaff80c0;

	lut_sub lut_5975 ({g164, g521, g522, g523}, g524);
	defparam lut_5975.LUT_SIZE = 4;
	defparam lut_5975.mask = 16'h5540;

	lut_sub lut_5989 ({g503, g506, g510, g516, g519, g1564}, g525);
	defparam lut_5989.LUT_SIZE = 6;
	defparam lut_5989.mask = 64'h0000000000000001;

	lut_sub lut_5998 ({g22, g24, g125, g123, g438}, g526);
	defparam lut_5998.LUT_SIZE = 5;
	defparam lut_5998.mask = 32'hef000000;

	lut_sub lut_6012 ({g355, g75, g91, g212}, g527);
	defparam lut_6012.LUT_SIZE = 4;
	defparam lut_6012.mask = 16'h50d0;

	lut_sub lut_6024 ({g17, g22, g24, g81}, g528);
	defparam lut_6024.LUT_SIZE = 4;
	defparam lut_6024.mask = 16'hc4cc;

	lut_sub lut_6038 ({g73, g468, g487, g528}, g529);
	defparam lut_6038.LUT_SIZE = 4;
	defparam lut_6038.mask = 16'h007f;

	lut_sub lut_6054 ({g75, g192, g513, g514, g527, g529}, g530);
	defparam lut_6054.LUT_SIZE = 6;
	defparam lut_6054.mask = 64'h0080000088888888;

	lut_sub lut_6071 ({g69, g154, g113, g119, g482}, g531);
	defparam lut_6071.LUT_SIZE = 5;
	defparam lut_6071.mask = 32'h50005111;

	lut_sub lut_6087 ({g24, g122, g113, g105, g174, g531}, g532);
	defparam lut_6087.LUT_SIZE = 6;
	defparam lut_6087.mask = 64'h2aaa00aa2aaa2aaa;

	lut_sub lut_6117 ({i_9_, i_10_, i_11_, i_15_, g174, g460}, g533);
	defparam lut_6117.LUT_SIZE = 6;
	defparam lut_6117.mask = 64'ha0a0a0a0a0a0aca0;

	lut_sub lut_6140 ({g88, g460}, g534);
	defparam lut_6140.LUT_SIZE = 2;
	defparam lut_6140.mask = 4'b0010;

	lut_sub lut_6149 ({g157, g191, g534, g496, g522}, g535);
	defparam lut_6149.LUT_SIZE = 5;
	defparam lut_6149.mask = 32'h00007fff;

	lut_sub lut_6172 ({g168, g435, g501, g533, g535}, g536);
	defparam lut_6172.LUT_SIZE = 5;
	defparam lut_6172.mask = 32'ha0aa8088;

	lut_sub lut_6189 ({g526, g1459, g530, g532, g536}, g537);
	defparam lut_6189.LUT_SIZE = 5;
	defparam lut_6189.mask = 32'h01000000;

	lut_sub lut_6195 ({i_14_, g102, g113}, g538);
	defparam lut_6195.LUT_SIZE = 3;
	defparam lut_6195.mask = 8'h02;

	lut_sub lut_6203 ({g119, g121, g213, g351}, g539);
	defparam lut_6203.LUT_SIZE = 4;
	defparam lut_6203.mask = 16'h4000;

	lut_sub lut_6208 ({i_9_, i_10_, i_11_, i_15_, g174}, g540);
	defparam lut_6208.LUT_SIZE = 5;
	defparam lut_6208.mask = 32'h20000002;

	lut_sub lut_6219 ({g69, g254, g402, g487, g539, g540}, g541);
	defparam lut_6219.LUT_SIZE = 6;
	defparam lut_6219.mask = 64'h4545450045454544;

	lut_sub lut_6246 ({g105, g186, g513, g514}, g542);
	defparam lut_6246.LUT_SIZE = 4;
	defparam lut_6246.mask = 16'hdf00;

	lut_sub lut_6258 ({g76, g81}, g543);
	defparam lut_6258.LUT_SIZE = 2;
	defparam lut_6258.mask = 4'b0100;

	lut_sub lut_6266 ({g105, g182, g543, g473}, g544);
	defparam lut_6266.LUT_SIZE = 4;
	defparam lut_6266.mask = 16'h7f00;

	lut_sub lut_6281 ({g22, g69, g113, g105, g482}, g545);
	defparam lut_6281.LUT_SIZE = 5;
	defparam lut_6281.mask = 32'h44444044;

	lut_sub lut_6295 ({g105, g487, g484, g522}, g546);
	defparam lut_6295.LUT_SIZE = 4;
	defparam lut_6295.mask = 16'h7f00;

	lut_sub lut_6310 ({g102, g483, g489, g484, g500}, g547);
	defparam lut_6310.LUT_SIZE = 5;
	defparam lut_6310.mask = 32'h00007fff;

	lut_sub lut_6333 ({g542, g544, g545, g546, g547}, g548);
	defparam lut_6333.LUT_SIZE = 5;
	defparam lut_6333.mask = 32'h80000000;

	lut_sub lut_6340 ({g538, g541, g548}, g549);
	defparam lut_6340.LUT_SIZE = 3;
	defparam lut_6340.mask = 8'h40;

	lut_sub lut_6350 ({g17, g22, g81, g142, g174, g351}, g550);
	defparam lut_6350.LUT_SIZE = 6;
	defparam lut_6350.mask = 64'hc8c800c8c8c8c8c8;

	lut_sub lut_6376 ({g22, g76}, g551);
	defparam lut_6376.LUT_SIZE = 2;
	defparam lut_6376.mask = 4'b0111;

	lut_sub lut_6384 ({g76, g69}, g552);
	defparam lut_6384.LUT_SIZE = 2;
	defparam lut_6384.mask = 4'b1011;

	lut_sub lut_6395 ({g17, g76, g135, g88, g460}, g553);
	defparam lut_6395.LUT_SIZE = 5;
	defparam lut_6395.mask = 32'hcfff0f5f;

	lut_sub lut_6427 ({g17, g76, g122, g81, g460}, g554);
	defparam lut_6427.LUT_SIZE = 5;
	defparam lut_6427.mask = 32'hfcfdf0f5;

	lut_sub lut_6455 ({g36, g460}, g555);
	defparam lut_6455.LUT_SIZE = 2;
	defparam lut_6455.mask = 4'b0010;

	lut_sub lut_6465 ({g102, g105, g555, g501, g543, g534}, g556);
	defparam lut_6465.LUT_SIZE = 6;
	defparam lut_6465.mask = 64'hf000ffff80008000;

	lut_sub lut_6492 ({g76, g113}, g557);
	defparam lut_6492.LUT_SIZE = 2;
	defparam lut_6492.mask = 4'b1000;

	lut_sub lut_6502 ({g125, g122, g123, g552, g511, g557}, g558);
	defparam lut_6502.LUT_SIZE = 6;
	defparam lut_6502.mask = 64'h08ff08aa080a080a;

	lut_sub lut_6530 ({g119, g121, g552, g511, g558}, g559);
	defparam lut_6530.LUT_SIZE = 5;
	defparam lut_6530.mask = 32'h55044404;

	lut_sub lut_6546 ({g76, g161, g122, g91, g88}, g560);
	defparam lut_6546.LUT_SIZE = 5;
	defparam lut_6546.mask = 32'h0d5d0000;

	lut_sub lut_6562 ({g17, g88, g113, g105, g460}, g561);
	defparam lut_6562.LUT_SIZE = 5;
	defparam lut_6562.mask = 32'h80888888;

	lut_sub lut_6574 ({g76, g91}, g562);
	defparam lut_6574.LUT_SIZE = 2;
	defparam lut_6574.mask = 4'b1000;

	lut_sub lut_6581 ({i_8_, g73, g486, g562}, g563);
	defparam lut_6581.LUT_SIZE = 4;
	defparam lut_6581.mask = 16'h0700;

	lut_sub lut_6590 ({g123, g555, g486}, g564);
	defparam lut_6590.LUT_SIZE = 3;
	defparam lut_6590.mask = 8'h70;

	lut_sub lut_6601 ({g36, g76, g88, g130, g460}, g565);
	defparam lut_6601.LUT_SIZE = 5;
	defparam lut_6601.mask = 32'h0c00cc88;

	lut_sub lut_6617 ({g76, g81, g91, g130, g460}, g566);
	defparam lut_6617.LUT_SIZE = 5;
	defparam lut_6617.mask = 32'hc0cc8088;

	lut_sub lut_6635 ({g560, g561, g563, g564, g565, g566}, g567);
	defparam lut_6635.LUT_SIZE = 6;
	defparam lut_6635.mask = 64'h8000000000000000;

	lut_sub lut_6643 ({i_8_, g73, g76, g88, g460}, g568);
	defparam lut_6643.LUT_SIZE = 5;
	defparam lut_6643.mask = 32'h00000032;

	lut_sub lut_6654 ({g76, g161, g157, g81, g88}, g569);
	defparam lut_6654.LUT_SIZE = 5;
	defparam lut_6654.mask = 32'h05370000;

	lut_sub lut_6665 ({i_10_, i_11_, i_15_, g76}, g570);
	defparam lut_6665.LUT_SIZE = 4;
	defparam lut_6665.mask = 16'h2000;

	lut_sub lut_6673 ({g123, g213, g551, g570}, g571);
	defparam lut_6673.LUT_SIZE = 4;
	defparam lut_6673.mask = 16'hcd05;

	lut_sub lut_6688 ({g17, g76, g125, g81, g225}, g572);
	defparam lut_6688.LUT_SIZE = 5;
	defparam lut_6688.mask = 32'h03005f00;

	lut_sub lut_6703 ({g135, g131, g562, g557}, g573);
	defparam lut_6703.LUT_SIZE = 4;
	defparam lut_6703.mask = 16'h8c8f;

	lut_sub lut_6718 ({i_8_, g73, g76, g113, g460}, g574);
	defparam lut_6718.LUT_SIZE = 5;
	defparam lut_6718.mask = 32'h008800c8;

	lut_sub lut_6732 ({g568, g569, g571, g572, g573, g574}, g575);
	defparam lut_6732.LUT_SIZE = 6;
	defparam lut_6732.mask = 64'h2000000000000000;

	lut_sub lut_6741 ({g17, g36, g76, g88, g131}, g576);
	defparam lut_6741.LUT_SIZE = 5;
	defparam lut_6741.mask = 32'h20a0a0a0;

	lut_sub lut_6755 ({g125, g131, g551, g543}, g577);
	defparam lut_6755.LUT_SIZE = 4;
	defparam lut_6755.mask = 16'h2f23;

	lut_sub lut_6768 ({g17, g460}, g578);
	defparam lut_6768.LUT_SIZE = 2;
	defparam lut_6768.mask = 4'b0010;

	lut_sub lut_6776 ({g102, g105, g578, g495}, g579);
	defparam lut_6776.LUT_SIZE = 4;
	defparam lut_6776.mask = 16'h5073;

	lut_sub lut_6791 ({i_15_, g151, g460, g576, g577, g579}, g580);
	defparam lut_6791.LUT_SIZE = 6;
	defparam lut_6791.mask = 64'h2020202020200020;

	lut_sub lut_6807 ({g1554, g1543, g559, g567, g575, g580}, g581);
	defparam lut_6807.LUT_SIZE = 6;
	defparam lut_6807.mask = 64'h0000000000000001;

	lut_sub lut_6813 ({i_12_, i_13_, i_14_, g75, g81}, g582);
	defparam lut_6813.LUT_SIZE = 5;
	defparam lut_6813.mask = 32'h00040040;

	lut_sub lut_6821 ({i_8_, g73, g501, g543}, g583);
	defparam lut_6821.LUT_SIZE = 4;
	defparam lut_6821.mask = 16'h0700;

	lut_sub lut_6831 ({i_8_, g73, g76, g88, g460}, g584);
	defparam lut_6831.LUT_SIZE = 5;
	defparam lut_6831.mask = 32'h00320000;

	lut_sub lut_6840 ({i_8_, g73, g552, g511}, g585);
	defparam lut_6840.LUT_SIZE = 4;
	defparam lut_6840.mask = 16'h000d;

	lut_sub lut_6850 ({i_8_, g73, g551, g578, g495}, g586);
	defparam lut_6850.LUT_SIZE = 5;
	defparam lut_6850.mask = 32'h007700f7;

	lut_sub lut_6872 ({g74, g513, g583, g584, g585, g586}, g587);
	defparam lut_6872.LUT_SIZE = 6;
	defparam lut_6872.mask = 64'h8000800000008000;

	lut_sub lut_6882 ({i_8_, g17, g73, g76, g511}, g588);
	defparam lut_6882.LUT_SIZE = 5;
	defparam lut_6882.mask = 32'h050d000c;

	lut_sub lut_6895 ({g582, g587, g588}, g589);
	defparam lut_6895.LUT_SIZE = 3;
	defparam lut_6895.mask = 8'h20;

	lut_sub lut_6902 ({g74, g259, g552}, g590);
	defparam lut_6902.LUT_SIZE = 3;
	defparam lut_6902.mask = 8'h8a;

	lut_sub lut_6911 ({g125, g168, g511}, g591);
	defparam lut_6911.LUT_SIZE = 3;
	defparam lut_6911.mask = 8'h15;

	lut_sub lut_6922 ({i_8_, g73, g155, g555, g486, g591}, g592);
	defparam lut_6922.LUT_SIZE = 6;
	defparam lut_6922.mask = 64'h80aa80a080aa8080;

	lut_sub lut_6946 ({g157, g262, g258, g551, g562, g501}, g593);
	defparam lut_6946.LUT_SIZE = 6;
	defparam lut_6946.mask = 64'h0fff0ccc0aaa0888;

	lut_sub lut_6980 ({g157, g135, g253, g254}, g594);
	defparam lut_6980.LUT_SIZE = 4;
	defparam lut_6980.mask = 16'h0100;

	lut_sub lut_6989 ({g258, g431, g543, g557, g594}, g595);
	defparam lut_6989.LUT_SIZE = 5;
	defparam lut_6989.mask = 32'hc4c4f5c4;

	lut_sub lut_7013 ({g167, g578, g590, g592, g593, g595}, g596);
	defparam lut_7013.LUT_SIZE = 6;
	defparam lut_7013.mask = 64'h0100010001000000;

	lut_sub lut_7021 ({g81, g482}, g597);
	defparam lut_7021.LUT_SIZE = 2;
	defparam lut_7021.mask = 4'b0001;

	lut_sub lut_7030 ({g159, g521, g597, g483, g489}, g598);
	defparam lut_7030.LUT_SIZE = 5;
	defparam lut_7030.mask = 32'h7fff0000;

	lut_sub lut_7053 ({g159, g154, g500, g522, g598}, g599);
	defparam lut_7053.LUT_SIZE = 5;
	defparam lut_7053.mask = 32'h80a080aa;

	lut_sub lut_7069 ({g154, g521, g597, g489, g599}, g600);
	defparam lut_7069.LUT_SIZE = 5;
	defparam lut_7069.mask = 32'h40005555;

	lut_sub lut_7083 ({i_14_, g88, g123}, g601);
	defparam lut_7083.LUT_SIZE = 3;
	defparam lut_7083.mask = 8'h02;

	lut_sub lut_7091 ({g123, g186, g513, g514}, g602);
	defparam lut_7091.LUT_SIZE = 4;
	defparam lut_7091.mask = 16'hdf00;

	lut_sub lut_7103 ({i_12_, i_13_, i_14_, g91, g123}, g603);
	defparam lut_7103.LUT_SIZE = 5;
	defparam lut_7103.mask = 32'h08080800;

	lut_sub lut_7113 ({g142, g521, g597, g489}, g604);
	defparam lut_7113.LUT_SIZE = 4;
	defparam lut_7113.mask = 16'h7f00;

	lut_sub lut_7125 ({g36, g174}, g605);
	defparam lut_7125.LUT_SIZE = 2;
	defparam lut_7125.mask = 4'b0010;

	lut_sub lut_7133 ({g17, g421, g408, g507}, g606);
	defparam lut_7133.LUT_SIZE = 4;
	defparam lut_7133.mask = 16'h0045;

	lut_sub lut_7141 ({g226, g461}, g607);
	defparam lut_7141.LUT_SIZE = 2;
	defparam lut_7141.mask = 4'b0100;

	lut_sub lut_7147 ({g81, g174}, g608);
	defparam lut_7147.LUT_SIZE = 2;
	defparam lut_7147.mask = 4'b1101;

	lut_sub lut_7156 ({g177, g392, g608}, g609);
	defparam lut_7156.LUT_SIZE = 3;
	defparam lut_7156.mask = 8'h23;

	lut_sub lut_7163 ({i_9_, i_11_, i_15_, g24}, g610);
	defparam lut_7163.LUT_SIZE = 4;
	defparam lut_7163.mask = 16'h0200;

	lut_sub lut_7171 ({g24, g88, g113, g174}, g611);
	defparam lut_7171.LUT_SIZE = 4;
	defparam lut_7171.mask = 16'h3075;

	lut_sub lut_7185 ({g1, i_15_, g34, g120, g174}, g612);
	defparam lut_7185.LUT_SIZE = 5;
	defparam lut_7185.mask = 32'h00000200;

	lut_sub lut_7194 ({g73, g159, g192, g611, g612}, g613);
	defparam lut_7194.LUT_SIZE = 5;
	defparam lut_7194.mask = 32'ha0aa2022;

	lut_sub lut_7212 ({g183, g383, g607, g609, g610, g613}, g614);
	defparam lut_7212.LUT_SIZE = 6;
	defparam lut_7212.mask = 64'h4000500000005000;

	lut_sub lut_7225 ({g144, g257, g254, g217, g226}, g615);
	defparam lut_7225.LUT_SIZE = 5;
	defparam lut_7225.mask = 32'h04000000;

	lut_sub lut_7235 ({g175, g422, g615, g555, g486, g578}, g616);
	defparam lut_7235.LUT_SIZE = 6;
	defparam lut_7235.mask = 64'haaff80c0aaff0000;

	lut_sub lut_7270 ({g161, g191, g534, g496, g522}, g617);
	defparam lut_7270.LUT_SIZE = 5;
	defparam lut_7270.mask = 32'h00007fff;

	lut_sub lut_7293 ({g125, g159, g438, g522, g617}, g618);
	defparam lut_7293.LUT_SIZE = 5;
	defparam lut_7293.mask = 32'h888a8888;

	lut_sub lut_7310 ({g601, g1458, g614, g616, g618}, g619);
	defparam lut_7310.LUT_SIZE = 5;
	defparam lut_7310.mask = 32'h00010000;

	lut_sub lut_7320 ({g550, g581, g589, g596, g600, g619}, g620);
	defparam lut_7320.LUT_SIZE = 6;
	defparam lut_7320.mask = 64'h0000000100000000;

	lut_sub lut_7330 ({g269, g499, g525, g537, g549, g620}, g621);
	defparam lut_7330.LUT_SIZE = 6;
	defparam lut_7330.mask = 64'h0000000000000001;

	lut_sub lut_7334 ({i_0_, i_1_, i_3_}, o_8_);
	defparam lut_7334.LUT_SIZE = 3;
	defparam lut_7334.mask = 8'h40;

	lut_sub lut_7342 ({g117, g129, g132, g153}, g623);
	defparam lut_7342.LUT_SIZE = 4;
	defparam lut_7342.mask = 16'h0001;

	lut_sub lut_7349 ({g18, g97, g578}, g624);
	defparam lut_7349.LUT_SIZE = 3;
	defparam lut_7349.mask = 8'h20;

	lut_sub lut_7354 ({i_12_, i_13_, i_14_, g22}, g625);
	defparam lut_7354.LUT_SIZE = 4;
	defparam lut_7354.mask = 16'h8088;

	lut_sub lut_7362 ({g19, g22}, g626);
	defparam lut_7362.LUT_SIZE = 2;
	defparam lut_7362.mask = 4'b0010;

	lut_sub lut_7367 ({i_12_, i_13_, i_14_, g88}, g627);
	defparam lut_7367.LUT_SIZE = 4;
	defparam lut_7367.mask = 16'h4044;

	lut_sub lut_7375 ({g19, g81}, g628);
	defparam lut_7375.LUT_SIZE = 2;
	defparam lut_7375.mask = 4'b1110;

	lut_sub lut_7382 ({i_12_, i_13_, i_14_, g81}, g629);
	defparam lut_7382.LUT_SIZE = 4;
	defparam lut_7382.mask = 16'h4044;

	lut_sub lut_7390 ({g19, g88}, g630);
	defparam lut_7390.LUT_SIZE = 2;
	defparam lut_7390.mask = 4'b0001;

	lut_sub lut_7400 ({g154, g624, g627, g628, g629, g630}, g631);
	defparam lut_7400.LUT_SIZE = 6;
	defparam lut_7400.mask = 64'hfffff7ff00000000;

	lut_sub lut_7440 ({g159, g154, g624, g625, g626, g631}, g632);
	defparam lut_7440.LUT_SIZE = 6;
	defparam lut_7440.mask = 64'h008000a08080aaaa;

	lut_sub lut_7460 ({g75, g102, g513, g632}, g633);
	defparam lut_7460.LUT_SIZE = 4;
	defparam lut_7460.mask = 16'h1151;

	lut_sub lut_7470 ({g19, g35}, g634);
	defparam lut_7470.LUT_SIZE = 2;
	defparam lut_7470.mask = 4'b1110;

	lut_sub lut_7478 ({g19, g36}, g635);
	defparam lut_7478.LUT_SIZE = 2;
	defparam lut_7478.mask = 4'b0001;

	lut_sub lut_7484 ({i_8_, g45, g394}, g636);
	defparam lut_7484.LUT_SIZE = 3;
	defparam lut_7484.mask = 8'h01;

	lut_sub lut_7491 ({i_9_, i_10_, i_11_, g135, g630, g636}, g637);
	defparam lut_7491.LUT_SIZE = 6;
	defparam lut_7491.mask = 64'h3075757530303030;

	lut_sub lut_7525 ({g17, g19, g102, g91, g88, g105}, g638);
	defparam lut_7525.LUT_SIZE = 6;
	defparam lut_7525.mask = 64'h0000a2a20000a2ff;

	lut_sub lut_7551 ({g634, g105, g383, g635, g637, g638}, g639);
	defparam lut_7551.LUT_SIZE = 6;
	defparam lut_7551.mask = 64'h0000808880888088;

	lut_sub lut_7564 ({i_13_, i_14_, g91}, g640);
	defparam lut_7564.LUT_SIZE = 3;
	defparam lut_7564.mask = 8'h80;

	lut_sub lut_7569 ({i_12_, i_13_, i_14_, g36}, g641);
	defparam lut_7569.LUT_SIZE = 4;
	defparam lut_7569.mask = 16'h4044;

	lut_sub lut_7577 ({g19, g113}, g642);
	defparam lut_7577.LUT_SIZE = 2;
	defparam lut_7577.mask = 4'b0010;

	lut_sub lut_7585 ({g125, g642, g628, g629}, g643);
	defparam lut_7585.LUT_SIZE = 4;
	defparam lut_7585.mask = 16'h00df;

	lut_sub lut_7600 ({g356, g640, g641, g629, g643}, g644);
	defparam lut_7600.LUT_SIZE = 5;
	defparam lut_7600.mask = 32'haaaa8000;

	lut_sub lut_7615 ({g164, g625, g627}, g645);
	defparam lut_7615.LUT_SIZE = 3;
	defparam lut_7615.mask = 8'h07;

	lut_sub lut_7624 ({g122, g217, g635}, g646);
	defparam lut_7624.LUT_SIZE = 3;
	defparam lut_7624.mask = 8'h15;

	lut_sub lut_7632 ({i_12_, i_13_, i_14_, g91, g105}, g647);
	defparam lut_7632.LUT_SIZE = 5;
	defparam lut_7632.mask = 32'h80008080;

	lut_sub lut_7640 ({g19, g86}, g648);
	defparam lut_7640.LUT_SIZE = 2;
	defparam lut_7640.mask = 4'b0001;

	lut_sub lut_7648 ({g102, g642, g635, g648}, g649);
	defparam lut_7648.LUT_SIZE = 4;
	defparam lut_7648.mask = 16'h007f;

	lut_sub lut_7663 ({g36, g76, g91, g88, g123}, g650);
	defparam lut_7663.LUT_SIZE = 5;
	defparam lut_7663.mask = 32'ha200aa00;

	lut_sub lut_7675 ({g19, g107}, g651);
	defparam lut_7675.LUT_SIZE = 2;
	defparam lut_7675.mask = 4'b0010;

	lut_sub lut_7681 ({g19, g91}, g652);
	defparam lut_7681.LUT_SIZE = 2;
	defparam lut_7681.mask = 4'b0010;

	lut_sub lut_7689 ({g634, g102, g651, g652}, g653);
	defparam lut_7689.LUT_SIZE = 4;
	defparam lut_7689.mask = 16'h0f07;

	lut_sub lut_7701 ({g4, g69}, g654);
	defparam lut_7701.LUT_SIZE = 2;
	defparam lut_7701.mask = 4'b0001;

	lut_sub lut_7708 ({g70, g511, g654}, g655);
	defparam lut_7708.LUT_SIZE = 3;
	defparam lut_7708.mask = 8'h80;

	lut_sub lut_7715 ({i_8_, i_6_, i_7_, g118, g655, g630}, g656);
	defparam lut_7715.LUT_SIZE = 6;
	defparam lut_7715.mask = 64'h0500000c05000500;

	lut_sub lut_7731 ({g647, g649, g650, g653, g656}, g657);
	defparam lut_7731.LUT_SIZE = 5;
	defparam lut_7731.mask = 32'h80000000;

	lut_sub lut_7740 ({g17, g19, g27, g226, g227}, g658);
	defparam lut_7740.LUT_SIZE = 5;
	defparam lut_7740.mask = 32'h000c005d;

	lut_sub lut_7754 ({i_8_, g17, g19, g36, g73}, g659);
	defparam lut_7754.LUT_SIZE = 5;
	defparam lut_7754.mask = 32'h00000105;

	lut_sub lut_7764 ({g135, g130, g131, g635}, g660);
	defparam lut_7764.LUT_SIZE = 4;
	defparam lut_7764.mask = 16'h5554;

	lut_sub lut_7778 ({g105, g543, g513, g635}, g661);
	defparam lut_7778.LUT_SIZE = 4;
	defparam lut_7778.mask = 16'hdf00;

	lut_sub lut_7793 ({g36, g76, g125, g91, g88}, g662);
	defparam lut_7793.LUT_SIZE = 5;
	defparam lut_7793.mask = 32'h0d000f00;

	lut_sub lut_7808 ({g658, g659, g660, g661, g662}, g663);
	defparam lut_7808.LUT_SIZE = 5;
	defparam lut_7808.mask = 32'h80000000;

	lut_sub lut_7813 ({i_12_, i_13_, i_14_, g113}, g664);
	defparam lut_7813.LUT_SIZE = 4;
	defparam lut_7813.mask = 16'h8088;

	lut_sub lut_7820 ({i_12_, i_13_, i_14_, g91}, g665);
	defparam lut_7820.LUT_SIZE = 4;
	defparam lut_7820.mask = 16'h8088;

	lut_sub lut_7831 ({g164, g253, g624, g664, g665}, g666);
	defparam lut_7831.LUT_SIZE = 5;
	defparam lut_7831.mask = 32'h08ff080f;

	lut_sub lut_7853 ({g125, g226, g408, g624, g666}, g667);
	defparam lut_7853.LUT_SIZE = 5;
	defparam lut_7853.mask = 32'h11151111;

	lut_sub lut_7867 ({g3, g19}, g668);
	defparam lut_7867.LUT_SIZE = 2;
	defparam lut_7867.mask = 4'b0001;

	lut_sub lut_7874 ({i_11_, i_15_, g53, g76, g668}, g669);
	defparam lut_7874.LUT_SIZE = 5;
	defparam lut_7874.mask = 32'haaaaaaa2;

	lut_sub lut_7895 ({i_8_, g73, g635, g652}, g670);
	defparam lut_7895.LUT_SIZE = 4;
	defparam lut_7895.mask = 16'h0700;

	lut_sub lut_7907 ({g75, g168, g350, g652, g669, g670}, g671);
	defparam lut_7907.LUT_SIZE = 6;
	defparam lut_7907.mask = 64'ha0a02020aaa02220;

	lut_sub lut_7931 ({g645, g646, g657, g663, g667, g671}, g672);
	defparam lut_7931.LUT_SIZE = 6;
	defparam lut_7931.mask = 64'h0001000000000000;

	lut_sub lut_7938 ({g253, g641, g635}, g673);
	defparam lut_7938.LUT_SIZE = 3;
	defparam lut_7938.mask = 8'h70;

	lut_sub lut_7948 ({g30, g120, g626, g630}, g674);
	defparam lut_7948.LUT_SIZE = 4;
	defparam lut_7948.mask = 16'h0007;

	lut_sub lut_7960 ({g164, g641, g628, g655, g665, g674}, g675);
	defparam lut_7960.LUT_SIZE = 6;
	defparam lut_7960.mask = 64'haaaaaaaa00080000;

	lut_sub lut_7986 ({g253, g625, g627, g629, g673, g675}, g676);
	defparam lut_7986.LUT_SIZE = 6;
	defparam lut_7986.mask = 64'h4000000044444444;

	lut_sub lut_7999 ({i_12_, i_13_, g17}, g677);
	defparam lut_7999.LUT_SIZE = 3;
	defparam lut_7999.mask = 8'h10;

	lut_sub lut_8008 ({i_14_, g142, g254, g425, g402, g677}, g678);
	defparam lut_8008.LUT_SIZE = 6;
	defparam lut_8008.mask = 64'h5544554455555050;

	lut_sub lut_8038 ({i_11_, i_15_, g19, g53, g401}, g679);
	defparam lut_8038.LUT_SIZE = 5;
	defparam lut_8038.mask = 32'h00000800;

	lut_sub lut_8048 ({g3, g19, g35, g425, g402, g353}, g680);
	defparam lut_8048.LUT_SIZE = 6;
	defparam lut_8048.mask = 64'h0000405000004454;

	lut_sub lut_8061 ({g80, i_11_, g636}, g681);
	defparam lut_8061.LUT_SIZE = 3;
	defparam lut_8061.mask = 8'h04;

	lut_sub lut_8070 ({g122, g123, g105, g642, g626}, g682);
	defparam lut_8070.LUT_SIZE = 5;
	defparam lut_8070.mask = 32'h8c8f888a;

	lut_sub lut_8088 ({i_12_, i_14_, g88, g408}, g683);
	defparam lut_8088.LUT_SIZE = 4;
	defparam lut_8088.mask = 16'h0020;

	lut_sub lut_8094 ({g4, g113}, g684);
	defparam lut_8094.LUT_SIZE = 2;
	defparam lut_8094.mask = 4'b1101;

	lut_sub lut_8104 ({g135, g131, g664, g684}, g685);
	defparam lut_8104.LUT_SIZE = 4;
	defparam lut_8104.mask = 16'hba30;

	lut_sub lut_8117 ({i_12_, i_13_, i_14_, g22, g142, g408}, g686);
	defparam lut_8117.LUT_SIZE = 6;
	defparam lut_8117.mask = 64'hc0000000e000e000;

	lut_sub lut_8131 ({i_8_, g73, g102, g562}, g687);
	defparam lut_8131.LUT_SIZE = 4;
	defparam lut_8131.mask = 16'h1115;

	lut_sub lut_8140 ({i_12_, i_14_, g113}, g688);
	defparam lut_8140.LUT_SIZE = 3;
	defparam lut_8140.mask = 8'h08;

	lut_sub lut_8150 ({g125, g164, g254, g217, g629, g688}, g689);
	defparam lut_8150.LUT_SIZE = 6;
	defparam lut_8150.mask = 64'haafa88c8aaaa8888;

	lut_sub lut_8185 ({g683, g685, g686, g687, g689}, g690);
	defparam lut_8185.LUT_SIZE = 5;
	defparam lut_8185.mask = 32'h40000000;

	lut_sub lut_8195 ({g676, g678, g679, g680, g1457, g690}, g691);
	defparam lut_8195.LUT_SIZE = 6;
	defparam lut_8195.mask = 64'h0000000010000000;

	lut_sub lut_8205 ({g30, g42, g118, g113, g460, g629}, g692);
	defparam lut_8205.LUT_SIZE = 6;
	defparam lut_8205.mask = 64'h000000c0005500d5;

	lut_sub lut_8222 ({i_12_, i_13_, i_14_, g88, g392, g407}, g693);
	defparam lut_8222.LUT_SIZE = 6;
	defparam lut_8222.mask = 64'h0000050000000300;

	lut_sub lut_8233 ({g131, g624, g625, g630}, g694);
	defparam lut_8233.LUT_SIZE = 4;
	defparam lut_8233.mask = 16'hf700;

	lut_sub lut_8247 ({g17, g19, g125, g694}, g695);
	defparam lut_8247.LUT_SIZE = 4;
	defparam lut_8247.mask = 16'haaa8;

	lut_sub lut_8263 ({g19, g69, g352, g692, g693, g695}, g696);
	defparam lut_8263.LUT_SIZE = 6;
	defparam lut_8263.mask = 64'h4040404040400040;

	lut_sub lut_8279 ({g633, g639, g644, g672, g691, g696}, g697);
	defparam lut_8279.LUT_SIZE = 6;
	defparam lut_8279.mask = 64'h0000000000000001;

	lut_sub lut_8286 ({g355, g35, g555}, g698);
	defparam lut_8286.LUT_SIZE = 3;
	defparam lut_8286.mask = 8'ha8;

	lut_sub lut_8294 ({g4, g81}, g699);
	defparam lut_8294.LUT_SIZE = 2;
	defparam lut_8294.mask = 4'b1110;

	lut_sub lut_8302 ({g19, g83}, g700);
	defparam lut_8302.LUT_SIZE = 2;
	defparam lut_8302.mask = 4'b1110;

	lut_sub lut_8312 ({g4, g69, g91, g668}, g701);
	defparam lut_8312.LUT_SIZE = 4;
	defparam lut_8312.mask = 16'haa20;

	lut_sub lut_8325 ({g634, g37, g75, g654, g668}, g702);
	defparam lut_8325.LUT_SIZE = 5;
	defparam lut_8325.mask = 32'hf0f0f070;

	lut_sub lut_8345 ({g4, g88}, g703);
	defparam lut_8345.LUT_SIZE = 2;
	defparam lut_8345.mask = 4'b1110;

	lut_sub lut_8356 ({i_8_, g73, g651, g699, g648, g703}, g704);
	defparam lut_8356.LUT_SIZE = 6;
	defparam lut_8356.mask = 64'h0000fbff00003333;

	lut_sub lut_8385 ({g18, g33, g73}, g705);
	defparam lut_8385.LUT_SIZE = 3;
	defparam lut_8385.mask = 8'h15;

	lut_sub lut_8396 ({g21, g23, g74, g704, g705}, g706);
	defparam lut_8396.LUT_SIZE = 5;
	defparam lut_8396.mask = 32'h80888080;

	lut_sub lut_8410 ({g21, g23, g75, g1531, g702, g706}, g707);
	defparam lut_8410.LUT_SIZE = 6;
	defparam lut_8410.mask = 64'h0004040400040004;

	lut_sub lut_8421 ({i_8_, g73, g108, g309}, g708);
	defparam lut_8421.LUT_SIZE = 4;
	defparam lut_8421.mask = 16'h0007;

	lut_sub lut_8430 ({g75, g486, g708}, g709);
	defparam lut_8430.LUT_SIZE = 3;
	defparam lut_8430.mask = 8'h8a;

	lut_sub lut_8440 ({g355, g35, g75, g555}, g710);
	defparam lut_8440.LUT_SIZE = 4;
	defparam lut_8440.mask = 16'h444c;

	lut_sub lut_8454 ({g74, g698, g196, g707, g709, g710}, g711);
	defparam lut_8454.LUT_SIZE = 6;
	defparam lut_8454.mask = 64'h0002000200000002;

	lut_sub lut_8463 ({g119, g254, g668}, g712);
	defparam lut_8463.LUT_SIZE = 3;
	defparam lut_8463.mask = 8'h45;

	lut_sub lut_8472 ({g123, g119, g654}, g713);
	defparam lut_8472.LUT_SIZE = 3;
	defparam lut_8472.mask = 8'h51;

	lut_sub lut_8481 ({g105, g121, g654}, g714);
	defparam lut_8481.LUT_SIZE = 3;
	defparam lut_8481.mask = 8'h51;

	lut_sub lut_8491 ({g19, g126, g122, g684}, g715);
	defparam lut_8491.LUT_SIZE = 4;
	defparam lut_8491.mask = 16'h2232;

	lut_sub lut_8504 ({g3, g19, g125, g126, g121}, g716);
	defparam lut_8504.LUT_SIZE = 5;
	defparam lut_8504.mask = 32'h000c005f;

	lut_sub lut_8520 ({g19, g75, g126, g715, g716}, g717);
	defparam lut_8520.LUT_SIZE = 5;
	defparam lut_8520.mask = 32'h88880888;

	lut_sub lut_8534 ({g125, g226, g684, g668}, g718);
	defparam lut_8534.LUT_SIZE = 4;
	defparam lut_8534.mask = 16'h50dc;

	lut_sub lut_8547 ({g70, g270, g511}, g719);
	defparam lut_8547.LUT_SIZE = 3;
	defparam lut_8547.mask = 8'h80;

	lut_sub lut_8554 ({g77, g719, g654}, g720);
	defparam lut_8554.LUT_SIZE = 3;
	defparam lut_8554.mask = 8'h20;

	lut_sub lut_8561 ({i_8_, i_6_, i_7_, g120, g508, g720}, g721);
	defparam lut_8561.LUT_SIZE = 6;
	defparam lut_8561.mask = 64'h0000000003000800;

	lut_sub lut_8573 ({g712, g713, g714, g717, g718, g721}, g722);
	defparam lut_8573.LUT_SIZE = 6;
	defparam lut_8573.mask = 64'h0800000000000000;

	lut_sub lut_8579 ({g81, g507}, g723);
	defparam lut_8579.LUT_SIZE = 2;
	defparam lut_8579.mask = 4'b0001;

	lut_sub lut_8587 ({i_9_, i_10_, g123, g315, g408, g723}, g724);
	defparam lut_8587.LUT_SIZE = 6;
	defparam lut_8587.mask = 64'h55005d0c55005500;

	lut_sub lut_8612 ({g17, g19, g357}, g725);
	defparam lut_8612.LUT_SIZE = 3;
	defparam lut_8612.mask = 8'ha8;

	lut_sub lut_8622 ({g121, g434, g341, g725}, g726);
	defparam lut_8622.LUT_SIZE = 4;
	defparam lut_8622.mask = 16'h0ace;

	lut_sub lut_8638 ({g167, g144, g334, g624, g724, g726}, g727);
	defparam lut_8638.LUT_SIZE = 6;
	defparam lut_8638.mask = 64'h8888008808080008;

	lut_sub lut_8652 ({g355, g35}, g728);
	defparam lut_8652.LUT_SIZE = 2;
	defparam lut_8652.mask = 4'b0001;

	lut_sub lut_8659 ({g355, g107, g486}, g729);
	defparam lut_8659.LUT_SIZE = 3;
	defparam lut_8659.mask = 8'ha2;

	lut_sub lut_8667 ({i_13_, i_14_, g36, g625}, g730);
	defparam lut_8667.LUT_SIZE = 4;
	defparam lut_8667.mask = 16'h8aaa;

	lut_sub lut_8683 ({g125, g131, g728, g534, g729, g730}, g731);
	defparam lut_8683.LUT_SIZE = 6;
	defparam lut_8683.mask = 64'h3000ffff10005555;

	lut_sub lut_8717 ({g21, g313, g254, g333}, g732);
	defparam lut_8717.LUT_SIZE = 4;
	defparam lut_8717.mask = 16'h05cd;

	lut_sub lut_8732 ({g87, g125, g122, g272, g534}, g733);
	defparam lut_8732.LUT_SIZE = 5;
	defparam lut_8732.mask = 32'hf000f888;

	lut_sub lut_8750 ({g161, g451, g732, g733}, g734);
	defparam lut_8750.LUT_SIZE = 4;
	defparam lut_8750.mask = 16'h4404;

	lut_sub lut_8756 ({i_12_, i_13_, i_14_}, g735);
	defparam lut_8756.LUT_SIZE = 3;
	defparam lut_8756.mask = 8'h28;

	lut_sub lut_8762 ({i_9_, i_10_, i_15_, g19}, g736);
	defparam lut_8762.LUT_SIZE = 4;
	defparam lut_8762.mask = 16'h0400;

	lut_sub lut_8770 ({g68, g126, g508, g736}, g737);
	defparam lut_8770.LUT_SIZE = 4;
	defparam lut_8770.mask = 16'h0888;

	lut_sub lut_8778 ({g22, g507}, g738);
	defparam lut_8778.LUT_SIZE = 2;
	defparam lut_8778.mask = 4'b0100;

	lut_sub lut_8785 ({g562, g737, g738}, g739);
	defparam lut_8785.LUT_SIZE = 3;
	defparam lut_8785.mask = 8'h20;

	lut_sub lut_8793 ({i_15_, g19, g428, g68, g429}, g740);
	defparam lut_8793.LUT_SIZE = 5;
	defparam lut_8793.mask = 32'hc4d50000;

	lut_sub lut_8810 ({g27, g105, g425, g735, g739, g740}, g741);
	defparam lut_8810.LUT_SIZE = 6;
	defparam lut_8810.mask = 64'h2222aaff2022a0ff;

	lut_sub lut_8845 ({g126, g176, g642}, g742);
	defparam lut_8845.LUT_SIZE = 3;
	defparam lut_8845.mask = 8'h2a;

	lut_sub lut_8853 ({g3, i_12_, i_13_, i_14_, g69}, g743);
	defparam lut_8853.LUT_SIZE = 5;
	defparam lut_8853.mask = 32'h40447347;

	lut_sub lut_8873 ({g73, g164, g402, g742, g743}, g744);
	defparam lut_8873.LUT_SIZE = 5;
	defparam lut_8873.mask = 32'h2f232323;

	lut_sub lut_8894 ({g157, g78, g333, g723}, g745);
	defparam lut_8894.LUT_SIZE = 4;
	defparam lut_8894.mask = 16'h00f7;

	lut_sub lut_8909 ({g157, g90, g125, g728, g729}, g746);
	defparam lut_8909.LUT_SIZE = 5;
	defparam lut_8909.mask = 32'hf5f5c400;

	lut_sub lut_8932 ({g165, g217, g729, g745, g746}, g747);
	defparam lut_8932.LUT_SIZE = 5;
	defparam lut_8932.mask = 32'h44040404;

	lut_sub lut_8946 ({g727, g1518, g734, g741, g744, g747}, g748);
	defparam lut_8946.LUT_SIZE = 6;
	defparam lut_8946.mask = 64'h0000000000000001;

	lut_sub lut_8951 ({i_9_, i_10_, i_11_, i_15_, g507}, g749);
	defparam lut_8951.LUT_SIZE = 5;
	defparam lut_8951.mask = 32'h01100000;

	lut_sub lut_8960 ({i_6_, g120, g135, g113, g507}, g750);
	defparam lut_8960.LUT_SIZE = 5;
	defparam lut_8960.mask = 32'h40ff4040;

	lut_sub lut_8975 ({i_9_, i_10_, i_11_, i_15_, g76}, g751);
	defparam lut_8975.LUT_SIZE = 5;
	defparam lut_8975.mask = 32'h00000220;

	lut_sub lut_8984 ({g185, g416, g562, g751}, g752);
	defparam lut_8984.LUT_SIZE = 4;
	defparam lut_8984.mask = 16'h8000;

	lut_sub lut_8993 ({g113, g507, g749, g750, g752}, g753);
	defparam lut_8993.LUT_SIZE = 5;
	defparam lut_8993.mask = 32'h23332323;

	lut_sub lut_9010 ({i_15_, i_12_, i_13_, i_14_, g112}, g754);
	defparam lut_9010.LUT_SIZE = 5;
	defparam lut_9010.mask = 32'h01014044;

	lut_sub lut_9019 ({i_9_, i_10_, i_15_, g507}, g755);
	defparam lut_9019.LUT_SIZE = 4;
	defparam lut_9019.mask = 16'h0100;

	lut_sub lut_9027 ({i_8_, g73, g130, g754, g755}, g756);
	defparam lut_9027.LUT_SIZE = 5;
	defparam lut_9027.mask = 32'h70757070;

	lut_sub lut_9050 ({g161, g119, g175, g508, g505, g756}, g757);
	defparam lut_9050.LUT_SIZE = 6;
	defparam lut_9050.mask = 64'h8888808088008000;

	lut_sub lut_9067 ({g177, g183, g278, g392, g501}, g758);
	defparam lut_9067.LUT_SIZE = 5;
	defparam lut_9067.mask = 32'h13333333;

	lut_sub lut_9091 ({g161, g90, g125, g281, g728, g555}, g759);
	defparam lut_9091.LUT_SIZE = 6;
	defparam lut_9091.mask = 64'hff88ff88c0800000;

	lut_sub lut_9122 ({g159, g336, g627, g758, g759}, g760);
	defparam lut_9122.LUT_SIZE = 5;
	defparam lut_9122.mask = 32'h00404444;

	lut_sub lut_9132 ({g343, g626}, g761);
	defparam lut_9132.LUT_SIZE = 2;
	defparam lut_9132.mask = 4'b0010;

	lut_sub lut_9140 ({g27, g168, g735, g719}, g762);
	defparam lut_9140.LUT_SIZE = 4;
	defparam lut_9140.mask = 16'h0a0b;

	lut_sub lut_9153 ({g125, g413, g439, g761, g762}, g763);
	defparam lut_9153.LUT_SIZE = 5;
	defparam lut_9153.mask = 32'h222a2222;

	lut_sub lut_9171 ({g753, g582, g587, g757, g760, g763}, g764);
	defparam lut_9171.LUT_SIZE = 6;
	defparam lut_9171.mask = 64'h0001000000000000;

	lut_sub lut_9177 ({g75, g197}, g765);
	defparam lut_9177.LUT_SIZE = 2;
	defparam lut_9177.mask = 4'b0100;

	lut_sub lut_9184 ({g164, g102, g397}, g766);
	defparam lut_9184.LUT_SIZE = 3;
	defparam lut_9184.mask = 8'h15;

	lut_sub lut_9193 ({i_7_, g17, g72, g76}, g767);
	defparam lut_9193.LUT_SIZE = 4;
	defparam lut_9193.mask = 16'h0002;

	lut_sub lut_9203 ({g102, g257, g313, g217, g737, g684}, g768);
	defparam lut_9203.LUT_SIZE = 6;
	defparam lut_9203.mask = 64'hf131313131313131;

	lut_sub lut_9237 ({g142, g749, g766, g767, g768}, g769);
	defparam lut_9237.LUT_SIZE = 5;
	defparam lut_9237.mask = 32'h40004040;

	lut_sub lut_9246 ({i_15_, g19, g445, g176}, g770);
	defparam lut_9246.LUT_SIZE = 4;
	defparam lut_9246.mask = 16'h2203;

	lut_sub lut_9256 ({i_8_, g73, g508, g719}, g771);
	defparam lut_9256.LUT_SIZE = 4;
	defparam lut_9256.mask = 16'h0b00;

	lut_sub lut_9267 ({g105, g438, g439, g770, g771}, g772);
	defparam lut_9267.LUT_SIZE = 5;
	defparam lut_9267.mask = 32'h8888888a;

	lut_sub lut_9285 ({g765, g271, g284, g202, g769, g772}, g773);
	defparam lut_9285.LUT_SIZE = 6;
	defparam lut_9285.mask = 64'h0001000000000000;

	lut_sub lut_9294 ({i_8_, g165, g83, g182, g735, g723}, g774);
	defparam lut_9294.LUT_SIZE = 6;
	defparam lut_9294.mask = 64'h0000557700000f0f;

	lut_sub lut_9319 ({g87, g135, g272, g534}, g775);
	defparam lut_9319.LUT_SIZE = 4;
	defparam lut_9319.mask = 16'hf070;

	lut_sub lut_9333 ({g20, g355, g122, g495}, g776);
	defparam lut_9333.LUT_SIZE = 4;
	defparam lut_9333.mask = 16'h1113;

	lut_sub lut_9343 ({i_8_, i_12_, i_13_, i_14_, g22, g35}, g777);
	defparam lut_9343.LUT_SIZE = 6;
	defparam lut_9343.mask = 64'hc00cccc000505000;

	lut_sub lut_9363 ({g165, g339, g777}, g778);
	defparam lut_9363.LUT_SIZE = 3;
	defparam lut_9363.mask = 8'h07;

	lut_sub lut_9374 ({g122, g194, g775, g776, g778}, g779);
	defparam lut_9374.LUT_SIZE = 5;
	defparam lut_9374.mask = 32'h80808000;

	lut_sub lut_9385 ({g85, g96, g99, g774, g779}, g780);
	defparam lut_9385.LUT_SIZE = 5;
	defparam lut_9385.mask = 32'h00000040;

	lut_sub lut_9395 ({g722, g322, g748, g764, g773, g780}, g781);
	defparam lut_9395.LUT_SIZE = 6;
	defparam lut_9395.mask = 64'h0000000000000001;

	lut_sub lut_9405 ({g346, g354, g361, g387, g411, g581}, g782);
	defparam lut_9405.LUT_SIZE = 6;
	defparam lut_9405.mask = 64'h0000000000010000;

	lut_sub lut_9412 ({g21, g23, g122}, g783);
	defparam lut_9412.LUT_SIZE = 3;
	defparam lut_9412.mask = 8'h45;

	lut_sub lut_9421 ({g122, g699, g700}, g784);
	defparam lut_9421.LUT_SIZE = 3;
	defparam lut_9421.mask = 8'h0e;

	lut_sub lut_9432 ({g634, g135, g651, g648, g703}, g785);
	defparam lut_9432.LUT_SIZE = 5;
	defparam lut_9432.mask = 32'hff00bf00;

	lut_sub lut_9455 ({g18, g33, g135, g122, g785}, g786);
	defparam lut_9455.LUT_SIZE = 5;
	defparam lut_9455.mask = 32'haa080808;

	lut_sub lut_9470 ({g122, g648, g783, g784, g786}, g787);
	defparam lut_9470.LUT_SIZE = 5;
	defparam lut_9470.mask = 32'h40404000;

	lut_sub lut_9480 ({g23, g102, g684, g703}, g788);
	defparam lut_9480.LUT_SIZE = 4;
	defparam lut_9480.mask = 16'h0f0e;

	lut_sub lut_9495 ({g37, g102, g105, g699, g700}, g789);
	defparam lut_9495.LUT_SIZE = 5;
	defparam lut_9495.mask = 32'h0f003f11;

	lut_sub lut_9515 ({g4, g102, g91, g788, g789}, g790);
	defparam lut_9515.LUT_SIZE = 5;
	defparam lut_9515.mask = 32'h44444404;

	lut_sub lut_9529 ({g144, g164, g684, g703}, g791);
	defparam lut_9529.LUT_SIZE = 4;
	defparam lut_9529.mask = 16'h0cae;

	lut_sub lut_9544 ({g19, g126, g254, g790, g791}, g792);
	defparam lut_9544.LUT_SIZE = 5;
	defparam lut_9544.mask = 32'h22220222;

	lut_sub lut_9558 ({g19, g126, g74, g684}, g793);
	defparam lut_9558.LUT_SIZE = 4;
	defparam lut_9558.mask = 16'h2232;

	lut_sub lut_9570 ({g4, g75, g91, g651}, g794);
	defparam lut_9570.LUT_SIZE = 4;
	defparam lut_9570.mask = 16'h50d0;

	lut_sub lut_9583 ({g21, g49, g33, g120, g648}, g795);
	defparam lut_9583.LUT_SIZE = 5;
	defparam lut_9583.mask = 32'h00130033;

	lut_sub lut_9598 ({g634, g131, g648, g700, g795}, g796);
	defparam lut_9598.LUT_SIZE = 5;
	defparam lut_9598.mask = 32'h00aa20aa;

	lut_sub lut_9615 ({g634, g125, g131, g651, g796}, g797);
	defparam lut_9615.LUT_SIZE = 5;
	defparam lut_9615.mask = 32'h45004545;

	lut_sub lut_9631 ({g21, g142, g227, g668}, g798);
	defparam lut_9631.LUT_SIZE = 4;
	defparam lut_9631.mask = 16'h11f1;

	lut_sub lut_9645 ({g23, g123, g684, g703}, g799);
	defparam lut_9645.LUT_SIZE = 4;
	defparam lut_9645.mask = 16'hf0e0;

	lut_sub lut_9659 ({g18, g23, g105, g684}, g800);
	defparam lut_9659.LUT_SIZE = 4;
	defparam lut_9659.mask = 16'hc8cc;

	lut_sub lut_9673 ({g33, g131, g225, g227}, g801);
	defparam lut_9673.LUT_SIZE = 4;
	defparam lut_9673.mask = 16'h00f7;

	lut_sub lut_9686 ({i_8_, g73, g684, g703}, g802);
	defparam lut_9686.LUT_SIZE = 4;
	defparam lut_9686.mask = 16'h000e;

	lut_sub lut_9695 ({g18, g102, g654}, g803);
	defparam lut_9695.LUT_SIZE = 3;
	defparam lut_9695.mask = 8'h13;

	lut_sub lut_9705 ({g23, g130, g699, g703}, g804);
	defparam lut_9705.LUT_SIZE = 4;
	defparam lut_9705.mask = 16'hf0e0;

	lut_sub lut_9721 ({g799, g800, g801, g802, g803, g804}, g805);
	defparam lut_9721.LUT_SIZE = 6;
	defparam lut_9721.mask = 64'h8000000000000000;

	lut_sub lut_9728 ({g18, g33, g142}, g806);
	defparam lut_9728.LUT_SIZE = 3;
	defparam lut_9728.mask = 8'h2a;

	lut_sub lut_9739 ({g4, g36, g91, g123, g130}, g807);
	defparam lut_9739.LUT_SIZE = 5;
	defparam lut_9739.mask = 32'h0000e0ee;

	lut_sub lut_9757 ({g125, g122, g105, g651, g700, g703}, g808);
	defparam lut_9757.LUT_SIZE = 6;
	defparam lut_9757.mask = 64'h55ff505010301010;

	lut_sub lut_9787 ({g142, g699, g700, g806, g807, g808}, g809);
	defparam lut_9787.LUT_SIZE = 6;
	defparam lut_9787.mask = 64'h0000004040404040;

	lut_sub lut_9801 ({g793, g794, g797, g798, g805, g809}, g810);
	defparam lut_9801.LUT_SIZE = 6;
	defparam lut_9801.mask = 64'h0010000000000000;

	lut_sub lut_9811 ({g211, g216, g252, g787, g792, g810}, g811);
	defparam lut_9811.LUT_SIZE = 6;
	defparam lut_9811.mask = 64'h0000000000000001;

	lut_sub lut_9821 ({g623, g697, g711, g781, g782, g811}, g812);
	defparam lut_9821.LUT_SIZE = 6;
	defparam lut_9821.mask = 64'h0000000000000001;

	lut_sub lut_9828 ({g581, g589, g596}, g813);
	defparam lut_9828.LUT_SIZE = 3;
	defparam lut_9828.mask = 8'h01;

	lut_sub lut_9837 ({g712, g713, g714, g717, g718}, g814);
	defparam lut_9837.LUT_SIZE = 5;
	defparam lut_9837.mask = 32'h20000000;

	lut_sub lut_9844 ({i_11_, i_15_, g19, g53, g105}, g815);
	defparam lut_9844.LUT_SIZE = 5;
	defparam lut_9844.mask = 32'h00000200;

	lut_sub lut_9851 ({g112, g154, g130}, g816);
	defparam lut_9851.LUT_SIZE = 3;
	defparam lut_9851.mask = 8'h0e;

	lut_sub lut_9861 ({i_15_, g4, g34, g155, g816}, g817);
	defparam lut_9861.LUT_SIZE = 5;
	defparam lut_9861.mask = 32'h0000005d;

	lut_sub lut_9870 ({i_9_, i_11_, i_15_, g4}, g818);
	defparam lut_9870.LUT_SIZE = 4;
	defparam lut_9870.mask = 16'h1000;

	lut_sub lut_9878 ({g125, g159, g703, g818}, g819);
	defparam lut_9878.LUT_SIZE = 4;
	defparam lut_9878.mask = 16'hc0d5;

	lut_sub lut_9893 ({g19, g27, g102, g165, g324}, g820);
	defparam lut_9893.LUT_SIZE = 5;
	defparam lut_9893.mask = 32'h0000111f;

	lut_sub lut_9908 ({g21, g164, g105, g819, g820}, g821);
	defparam lut_9908.LUT_SIZE = 5;
	defparam lut_9908.mask = 32'h88880800;

	lut_sub lut_9921 ({g18, g167, g815, g817, g821}, g822);
	defparam lut_9921.LUT_SIZE = 5;
	defparam lut_9921.mask = 32'h40404000;

	lut_sub lut_9933 ({g814, g707, g787, g792, g810, g822}, g823);
	defparam lut_9933.LUT_SIZE = 6;
	defparam lut_9933.mask = 64'h0000000000000001;

	lut_sub lut_9941 ({g80, i_11_, i_15_, g76, g414, g447}, g824);
	defparam lut_9941.LUT_SIZE = 6;
	defparam lut_9941.mask = 64'h0000000000c000a0;

	lut_sub lut_9951 ({g164, g105, g562}, g825);
	defparam lut_9951.LUT_SIZE = 3;
	defparam lut_9951.mask = 8'h45;

	lut_sub lut_9961 ({g87, g154, g557, g518}, g826);
	defparam lut_9961.LUT_SIZE = 4;
	defparam lut_9961.mask = 16'h7530;

	lut_sub lut_9976 ({g17, g76, g107, g168, g105}, g827);
	defparam lut_9976.LUT_SIZE = 5;
	defparam lut_9976.mask = 32'ha000b300;

	lut_sub lut_9990 ({i_6_, g120, g159, g562, g751}, g828);
	defparam lut_9990.LUT_SIZE = 5;
	defparam lut_9990.mask = 32'h30753030;

	lut_sub lut_10010 ({g159, g89, g684, g826, g827, g828}, g829);
	defparam lut_10010.LUT_SIZE = 6;
	defparam lut_10010.mask = 64'h0000008080808080;

	lut_sub lut_10023 ({g125, g165, g495, g825, g829}, g830);
	defparam lut_10023.LUT_SIZE = 5;
	defparam lut_10023.mask = 32'h44404040;

	lut_sub lut_10037 ({g161, g90, g413, g217, g501, g736}, g831);
	defparam lut_10037.LUT_SIZE = 6;
	defparam lut_10037.mask = 64'haafaaafa88c80000;

	lut_sub lut_10071 ({g78, g356, g392, g486, g534, g831}, g832);
	defparam lut_10071.LUT_SIZE = 6;
	defparam lut_10071.mask = 64'h5500400055554040;

	lut_sub lut_10094 ({g127, g402, g443, g642, g655}, g833);
	defparam lut_10094.LUT_SIZE = 5;
	defparam lut_10094.mask = 32'h45cf00cf;

	lut_sub lut_10116 ({g440, g446, g626, g628}, g834);
	defparam lut_10116.LUT_SIZE = 4;
	defparam lut_10116.mask = 16'hba30;

	lut_sub lut_10132 ({g61, g824, g830, g832, g833, g834}, g835);
	defparam lut_10132.LUT_SIZE = 6;
	defparam lut_10132.mask = 64'h0000000000020000;

	lut_sub lut_10140 ({g98, g225, g213, g425}, g836);
	defparam lut_10140.LUT_SIZE = 4;
	defparam lut_10140.mask = 16'h00bf;

	lut_sub lut_10155 ({g164, g79, g142, g402, g392}, g837);
	defparam lut_10155.LUT_SIZE = 5;
	defparam lut_10155.mask = 32'hfd00ff00;

	lut_sub lut_10178 ({g49, g33, g166, g401, g534}, g838);
	defparam lut_10178.LUT_SIZE = 5;
	defparam lut_10178.mask = 32'h00cc05cd;

	lut_sub lut_10197 ({g130, g425, g648, g688, g838}, g839);
	defparam lut_10197.LUT_SIZE = 5;
	defparam lut_10197.mask = 32'h8088a0aa;

	lut_sub lut_10214 ({g22, g76, g83, g435, g444}, g840);
	defparam lut_10214.LUT_SIZE = 5;
	defparam lut_10214.mask = 32'hae000c00;

	lut_sub lut_10227 ({i_8_, i_6_, i_7_, g21, g23, g118}, g841);
	defparam lut_10227.LUT_SIZE = 6;
	defparam lut_10227.mask = 64'h0000440005000000;

	lut_sub lut_10238 ({g17, g19, g434, g841}, g842);
	defparam lut_10238.LUT_SIZE = 4;
	defparam lut_10238.mask = 16'haaa8;

	lut_sub lut_10252 ({g109, g157, g422, g842}, g843);
	defparam lut_10252.LUT_SIZE = 4;
	defparam lut_10252.mask = 16'h5540;

	lut_sub lut_10266 ({g836, g837, g1511, g839, g840, g843}, g844);
	defparam lut_10266.LUT_SIZE = 6;
	defparam lut_10266.mask = 64'h0004000000000000;

	lut_sub lut_10276 ({g173, g813, g697, g823, g835, g844}, g845);
	defparam lut_10276.LUT_SIZE = 6;
	defparam lut_10276.mask = 64'h0000000000000001;

	lut_sub lut_10283 ({i_0_, i_1_, g15, g32, g39}, g846);
	defparam lut_10283.LUT_SIZE = 5;
	defparam lut_10283.mask = 32'h88888088;

	lut_sub lut_10295 ({g4, g86}, g847);
	defparam lut_10295.LUT_SIZE = 2;
	defparam lut_10295.mask = 4'b1110;

	lut_sub lut_10302 ({i_12_, i_13_, i_14_, g86}, g848);
	defparam lut_10302.LUT_SIZE = 4;
	defparam lut_10302.mask = 16'hfbbb;

	lut_sub lut_10319 ({i_12_, i_13_, i_14_, g35}, g849);
	defparam lut_10319.LUT_SIZE = 4;
	defparam lut_10319.mask = 16'h0444;

	lut_sub lut_10326 ({i_12_, i_13_, i_14_, g83}, g850);
	defparam lut_10326.LUT_SIZE = 4;
	defparam lut_10326.mask = 16'h0444;

	lut_sub lut_10334 ({g4, g35}, g851);
	defparam lut_10334.LUT_SIZE = 2;
	defparam lut_10334.mask = 4'b1110;

	lut_sub lut_10342 ({g4, g107}, g852);
	defparam lut_10342.LUT_SIZE = 2;
	defparam lut_10342.mask = 4'b0010;

	lut_sub lut_10347 ({i_12_, i_13_, i_14_, g107}, g853);
	defparam lut_10347.LUT_SIZE = 4;
	defparam lut_10347.mask = 16'h0888;

	lut_sub lut_10358 ({g253, g849, g852, g848, g853}, g854);
	defparam lut_10358.LUT_SIZE = 5;
	defparam lut_10358.mask = 32'hdfff0000;

	lut_sub lut_10382 ({g164, g849, g847, g850, g851, g854}, g855);
	defparam lut_10382.LUT_SIZE = 6;
	defparam lut_10382.mask = 64'haaaaaaaa00200000;

	lut_sub lut_10407 ({g125, g164, g847, g848, g855}, g856);
	defparam lut_10407.LUT_SIZE = 5;
	defparam lut_10407.mask = 32'h55110501;

	lut_sub lut_10421 ({g4, g126}, g857);
	defparam lut_10421.LUT_SIZE = 2;
	defparam lut_10421.mask = 4'b0010;

	lut_sub lut_10429 ({i_8_, g73, g102, g851, g857}, g858);
	defparam lut_10429.LUT_SIZE = 5;
	defparam lut_10429.mask = 32'h0cdd0c5d;

	lut_sub lut_10452 ({g21, g73, g413, g847, g858}, g859);
	defparam lut_10452.LUT_SIZE = 5;
	defparam lut_10452.mask = 32'h2a220a02;

	lut_sub lut_10464 ({i_9_, i_10_, i_11_, i_15_, g460}, g860);
	defparam lut_10464.LUT_SIZE = 5;
	defparam lut_10464.mask = 32'h00000880;

	lut_sub lut_10473 ({i_9_, g101, g165, g394, g860}, g861);
	defparam lut_10473.LUT_SIZE = 5;
	defparam lut_10473.mask = 32'h05050537;

	lut_sub lut_10491 ({g122, g847, g851, g861}, g862);
	defparam lut_10491.LUT_SIZE = 4;
	defparam lut_10491.mask = 16'haa02;

	lut_sub lut_10503 ({g130, g278, g421, g392}, g863);
	defparam lut_10503.LUT_SIZE = 4;
	defparam lut_10503.mask = 16'h0f07;

	lut_sub lut_10518 ({g25, g164, g402, g392, g863}, g864);
	defparam lut_10518.LUT_SIZE = 5;
	defparam lut_10518.mask = 32'h0800aaaa;

	lut_sub lut_10531 ({i_12_, i_13_, i_14_, g20}, g865);
	defparam lut_10531.LUT_SIZE = 4;
	defparam lut_10531.mask = 16'h0444;

	lut_sub lut_10541 ({g123, g130, g849, g853}, g866);
	defparam lut_10541.LUT_SIZE = 4;
	defparam lut_10541.mask = 16'h8c8f;

	lut_sub lut_10557 ({g4, g126, g91, g105, g309}, g867);
	defparam lut_10557.LUT_SIZE = 5;
	defparam lut_10557.mask = 32'h4444ccc4;

	lut_sub lut_10576 ({g123, g850, g865, g866, g867}, g868);
	defparam lut_10576.LUT_SIZE = 5;
	defparam lut_10576.mask = 32'h20002222;

	lut_sub lut_10585 ({i_9_, i_10_, i_11_, i_15_, g735}, g869);
	defparam lut_10585.LUT_SIZE = 5;
	defparam lut_10585.mask = 32'h04004000;

	lut_sub lut_10593 ({g24, g113, g492}, g870);
	defparam lut_10593.LUT_SIZE = 3;
	defparam lut_10593.mask = 8'h2a;

	lut_sub lut_10603 ({g24, g35, g161, g68}, g871);
	defparam lut_10603.LUT_SIZE = 4;
	defparam lut_10603.mask = 16'h0302;

	lut_sub lut_10614 ({g257, g351, g869, g870, g871}, g872);
	defparam lut_10614.LUT_SIZE = 5;
	defparam lut_10614.mask = 32'h22aa20a0;

	lut_sub lut_10631 ({g856, g859, g1501, g864, g1488}, g873);
	defparam lut_10631.LUT_SIZE = 5;
	defparam lut_10631.mask = 32'h00000001;

	lut_sub lut_10639 ({g159, g847, g850, g865}, g874);
	defparam lut_10639.LUT_SIZE = 4;
	defparam lut_10639.mask = 16'hf700;

	lut_sub lut_10650 ({i_12_, i_13_, i_14_, g27}, g875);
	defparam lut_10650.LUT_SIZE = 4;
	defparam lut_10650.mask = 16'h0444;

	lut_sub lut_10660 ({g159, g852, g853, g875}, g876);
	defparam lut_10660.LUT_SIZE = 4;
	defparam lut_10660.mask = 16'h7f00;

	lut_sub lut_10671 ({g3, i_12_, i_13_, i_14_}, g877);
	defparam lut_10671.LUT_SIZE = 4;
	defparam lut_10671.mask = 16'h002a;

	lut_sub lut_10680 ({g154, g849, g851}, g878);
	defparam lut_10680.LUT_SIZE = 3;
	defparam lut_10680.mask = 8'hb0;

	lut_sub lut_10691 ({g154, g877, g850, g865, g878}, g879);
	defparam lut_10691.LUT_SIZE = 5;
	defparam lut_10691.mask = 32'h8000aaaa;

	lut_sub lut_10709 ({g154, g847, g848, g874, g876, g879}, g880);
	defparam lut_10709.LUT_SIZE = 6;
	defparam lut_10709.mask = 64'h0000004040404040;

	lut_sub lut_10718 ({i_12_, i_13_, i_14_, g126}, g881);
	defparam lut_10718.LUT_SIZE = 4;
	defparam lut_10718.mask = 16'h0888;

	lut_sub lut_10725 ({i_9_, i_10_, i_11_, i_15_, g460}, g882);
	defparam lut_10725.LUT_SIZE = 5;
	defparam lut_10725.mask = 32'h00000888;

	lut_sub lut_10736 ({g24, g144, g126, g402, g882}, g883);
	defparam lut_10736.LUT_SIZE = 5;
	defparam lut_10736.mask = 32'hc0d50055;

	lut_sub lut_10754 ({g257, g356, g881, g883}, g884);
	defparam lut_10754.LUT_SIZE = 4;
	defparam lut_10754.mask = 16'ha888;

	lut_sub lut_10767 ({g125, g159, g438, g472, g877}, g885);
	defparam lut_10767.LUT_SIZE = 5;
	defparam lut_10767.mask = 32'h8a8f888c;

	lut_sub lut_10787 ({g480, g880, g884, g885}, g886);
	defparam lut_10787.LUT_SIZE = 4;
	defparam lut_10787.mask = 16'h0001;

	lut_sub lut_10793 ({g102, g881}, g887);
	defparam lut_10793.LUT_SIZE = 2;
	defparam lut_10793.mask = 4'b0001;

	lut_sub lut_10799 ({i_12_, i_13_, i_14_, g35, g102}, g888);
	defparam lut_10799.LUT_SIZE = 5;
	defparam lut_10799.mask = 32'h00101010;

	lut_sub lut_10807 ({i_12_, i_13_, i_14_, g86, g102}, g889);
	defparam lut_10807.LUT_SIZE = 5;
	defparam lut_10807.mask = 32'h00101010;

	lut_sub lut_10815 ({i_12_, i_13_, i_14_, g107, g102}, g890);
	defparam lut_10815.LUT_SIZE = 5;
	defparam lut_10815.mask = 32'h00404040;

	lut_sub lut_10824 ({g3, i_12_, i_13_, i_14_, g35, g105}, g891);
	defparam lut_10824.LUT_SIZE = 6;
	defparam lut_10824.mask = 64'h0020202000a0a0a0;

	lut_sub lut_10838 ({g83, g460}, g892);
	defparam lut_10838.LUT_SIZE = 2;
	defparam lut_10838.mask = 4'b0010;

	lut_sub lut_10848 ({g105, g295, g892, g700, g847, g852}, g893);
	defparam lut_10848.LUT_SIZE = 6;
	defparam lut_10848.mask = 64'hfdffffff00000000;

	lut_sub lut_10887 ({g888, g889, g890, g891, g893}, g894);
	defparam lut_10887.LUT_SIZE = 5;
	defparam lut_10887.mask = 32'h80000000;

	lut_sub lut_10895 ({g20, g164, g105, g460}, g895);
	defparam lut_10895.LUT_SIZE = 4;
	defparam lut_10895.mask = 16'h008a;

	lut_sub lut_10905 ({g159, g154, g849, g881}, g896);
	defparam lut_10905.LUT_SIZE = 4;
	defparam lut_10905.mask = 16'h8caf;

	lut_sub lut_10922 ({g3, g383, g460, g895, g1478}, g897);
	defparam lut_10922.LUT_SIZE = 5;
	defparam lut_10922.mask = 32'h44440444;

	lut_sub lut_10934 ({g4, g83}, g898);
	defparam lut_10934.LUT_SIZE = 2;
	defparam lut_10934.mask = 4'b1110;

	lut_sub lut_10943 ({g31, g528, g898}, g899);
	defparam lut_10943.LUT_SIZE = 3;
	defparam lut_10943.mask = 8'h40;

	lut_sub lut_10950 ({g107, g165, g460}, g900);
	defparam lut_10950.LUT_SIZE = 3;
	defparam lut_10950.mask = 8'h20;

	lut_sub lut_10960 ({g142, g392, g351, g496, g899, g900}, g901);
	defparam lut_10960.LUT_SIZE = 6;
	defparam lut_10960.mask = 64'h2222202022aa20a0;

	lut_sub lut_10983 ({g73, g144, g102, g165, g130}, g902);
	defparam lut_10983.LUT_SIZE = 5;
	defparam lut_10983.mask = 32'h40000000;

	lut_sub lut_10989 ({i_9_, i_10_, i_11_, i_15_, g4, g24}, g903);
	defparam lut_10989.LUT_SIZE = 6;
	defparam lut_10989.mask = 64'h000003000000a3a3;

	lut_sub lut_11005 ({g45, g86, g460}, g904);
	defparam lut_11005.LUT_SIZE = 3;
	defparam lut_11005.mask = 8'h02;

	lut_sub lut_11013 ({i_8_, g42, g72, g473, g904}, g905);
	defparam lut_11013.LUT_SIZE = 5;
	defparam lut_11013.mask = 32'h00000407;

	lut_sub lut_11025 ({g422, g852, g902, g903, g905}, g906);
	defparam lut_11025.LUT_SIZE = 5;
	defparam lut_11025.mask = 32'haa0a8808;

	lut_sub lut_11042 ({g119, g272, g425, g351, g468}, g907);
	defparam lut_11042.LUT_SIZE = 5;
	defparam lut_11042.mask = 32'hbb0baa0a;

	lut_sub lut_11066 ({g887, g894, g897, g901, g906, g907}, g908);
	defparam lut_11066.LUT_SIZE = 6;
	defparam lut_11066.mask = 64'h0000000100000000;

	lut_sub lut_11071 ({i_9_, i_10_, i_11_, i_15_, g4}, g909);
	defparam lut_11071.LUT_SIZE = 5;
	defparam lut_11071.mask = 32'h00041000;

	lut_sub lut_11080 ({i_15_, g102, g615, g350, g909}, g910);
	defparam lut_11080.LUT_SIZE = 5;
	defparam lut_11080.mask = 32'h11555050;

	lut_sub lut_11097 ({i_11_, i_15_, g4, g34, g125, g218}, g911);
	defparam lut_11097.LUT_SIZE = 6;
	defparam lut_11097.mask = 64'h0003000000050000;

	lut_sub lut_11106 ({i_14_, g27, g226}, g912);
	defparam lut_11106.LUT_SIZE = 3;
	defparam lut_11106.mask = 8'h20;

	lut_sub lut_11115 ({g123, g105, g852, g853, g875}, g913);
	defparam lut_11115.LUT_SIZE = 5;
	defparam lut_11115.mask = 32'h808088ff;

	lut_sub lut_11135 ({g164, g154, g853, g875, g913}, g914);
	defparam lut_11135.LUT_SIZE = 5;
	defparam lut_11135.mask = 32'h40554040;

	lut_sub lut_11150 ({g105, g851, g911, g912, g914}, g915);
	defparam lut_11150.LUT_SIZE = 5;
	defparam lut_11150.mask = 32'h00404040;

	lut_sub lut_11161 ({g126, g122, g105, g383, g460}, g916);
	defparam lut_11161.LUT_SIZE = 5;
	defparam lut_11161.mask = 32'ha8aa0000;

	lut_sub lut_11174 ({g24, g83, g699}, g917);
	defparam lut_11174.LUT_SIZE = 3;
	defparam lut_11174.mask = 8'h45;

	lut_sub lut_11185 ({g164, g213, g270, g402, g654}, g918);
	defparam lut_11185.LUT_SIZE = 5;
	defparam lut_11185.mask = 32'hb3a0a0a0;

	lut_sub lut_11201 ({i_12_, i_13_, i_14_, g27, g167}, g919);
	defparam lut_11201.LUT_SIZE = 5;
	defparam lut_11201.mask = 32'h13000000;

	lut_sub lut_11211 ({i_14_, g225, g213, g425, g919}, g920);
	defparam lut_11211.LUT_SIZE = 5;
	defparam lut_11211.mask = 32'h55554555;

	lut_sub lut_11234 ({g435, g916, g917, g918, g920}, g921);
	defparam lut_11234.LUT_SIZE = 5;
	defparam lut_11234.mask = 32'h02002200;

	lut_sub lut_11245 ({g5, g539, g910, g915, g921}, g922);
	defparam lut_11245.LUT_SIZE = 5;
	defparam lut_11245.mask = 32'h10100010;

	lut_sub lut_11257 ({g332, g823, g873, g886, g908, g922}, g923);
	defparam lut_11257.LUT_SIZE = 6;
	defparam lut_11257.mask = 64'h0000000000000001;

	lut_sub lut_11262 ({i_11_, g34}, g924);
	defparam lut_11262.LUT_SIZE = 2;
	defparam lut_11262.mask = 4'b0100;

	lut_sub lut_11271 ({g102, g337, g605, g635, g851}, g925);
	defparam lut_11271.LUT_SIZE = 5;
	defparam lut_11271.mask = 32'h0000bfff;

	lut_sub lut_11293 ({g43, g924, g394, g925}, g926);
	defparam lut_11293.LUT_SIZE = 4;
	defparam lut_11293.mask = 16'haaa8;

	lut_sub lut_11305 ({g3, i_12_, i_13_, i_14_, g69}, g927);
	defparam lut_11305.LUT_SIZE = 5;
	defparam lut_11305.mask = 32'h0401c431;

	lut_sub lut_11320 ({g17, g81, g174, g927}, g928);
	defparam lut_11320.LUT_SIZE = 4;
	defparam lut_11320.mask = 16'ha222;

	lut_sub lut_11331 ({g4, g27, g928}, g929);
	defparam lut_11331.LUT_SIZE = 3;
	defparam lut_11331.mask = 8'h54;

	lut_sub lut_11339 ({g892, g473}, g930);
	defparam lut_11339.LUT_SIZE = 2;
	defparam lut_11339.mask = 4'b1000;

	lut_sub lut_11346 ({i_15_, g428, g24, g460}, g931);
	defparam lut_11346.LUT_SIZE = 4;
	defparam lut_11346.mask = 16'ha0c0;

	lut_sub lut_11357 ({g468, g743, g770, g877}, g932);
	defparam lut_11357.LUT_SIZE = 4;
	defparam lut_11357.mask = 16'h8000;

	lut_sub lut_11365 ({g929, g930, g931, g932}, g933);
	defparam lut_11365.LUT_SIZE = 4;
	defparam lut_11365.mask = 16'h0004;

	lut_sub lut_11372 ({g342, g522, g630}, g934);
	defparam lut_11372.LUT_SIZE = 3;
	defparam lut_11372.mask = 8'h80;

	lut_sub lut_11380 ({g21, g397, g508, g934}, g935);
	defparam lut_11380.LUT_SIZE = 4;
	defparam lut_11380.mask = 16'h4000;

	lut_sub lut_11389 ({i_8_, g168, g898, g928, g933, g935}, g936);
	defparam lut_11389.LUT_SIZE = 6;
	defparam lut_11389.mask = 64'h0000ffee0000f0f0;

	lut_sub lut_11419 ({g102, g358, g487, g652, g852}, g937);
	defparam lut_11419.LUT_SIZE = 5;
	defparam lut_11419.mask = 32'h00007fff;

	lut_sub lut_11442 ({g19, g102, g113, g105, g174}, g938);
	defparam lut_11442.LUT_SIZE = 5;
	defparam lut_11442.mask = 32'h8080c0f0;

	lut_sub lut_11458 ({g4, g126, g102, g105, g176}, g939);
	defparam lut_11458.LUT_SIZE = 5;
	defparam lut_11458.mask = 32'h8800cf00;

	lut_sub lut_11474 ({g105, g853, g937, g938, g939}, g940);
	defparam lut_11474.LUT_SIZE = 5;
	defparam lut_11474.mask = 32'h80008080;

	lut_sub lut_11484 ({g102, g105, g654, g847}, g941);
	defparam lut_11484.LUT_SIZE = 4;
	defparam lut_11484.mask = 16'h30ba;

	lut_sub lut_11499 ({g305, g307, g308, g310, g941}, g942);
	defparam lut_11499.LUT_SIZE = 5;
	defparam lut_11499.mask = 32'h80000000;

	lut_sub lut_11505 ({i_15_, i_12_, i_13_, i_14_, g112, g105}, g943);
	defparam lut_11505.LUT_SIZE = 6;
	defparam lut_11505.mask = 64'h0222202220002020;

	lut_sub lut_11520 ({g105, g719, g943}, g944);
	defparam lut_11520.LUT_SIZE = 3;
	defparam lut_11520.mask = 8'h2a;

	lut_sub lut_11529 ({g22, g48, g174}, g945);
	defparam lut_11529.LUT_SIZE = 3;
	defparam lut_11529.mask = 8'h4c;

	lut_sub lut_11538 ({g105, g188, g875}, g946);
	defparam lut_11538.LUT_SIZE = 3;
	defparam lut_11538.mask = 8'h70;

	lut_sub lut_11550 ({g236, g237, g238, g240, g241, g946}, g947);
	defparam lut_11550.LUT_SIZE = 6;
	defparam lut_11550.mask = 64'h0800000000000000;

	lut_sub lut_11557 ({g337, g605, g635}, g948);
	defparam lut_11557.LUT_SIZE = 3;
	defparam lut_11557.mask = 8'h80;

	lut_sub lut_11563 ({g770, g898}, g949);
	defparam lut_11563.LUT_SIZE = 2;
	defparam lut_11563.mask = 4'b0100;

	lut_sub lut_11571 ({g105, g948, g949, g638}, g950);
	defparam lut_11571.LUT_SIZE = 4;
	defparam lut_11571.mask = 16'h02aa;

	lut_sub lut_11585 ({g944, g360, g1543, g1467, g947, g950}, g951);
	defparam lut_11585.LUT_SIZE = 6;
	defparam lut_11585.mask = 64'h0000000000000001;

	lut_sub lut_11591 ({i_15_, i_12_, i_13_, i_14_, g429, g105}, g952);
	defparam lut_11591.LUT_SIZE = 6;
	defparam lut_11591.mask = 64'h0222202220002020;

	lut_sub lut_11605 ({i_15_, i_12_, i_13_, i_14_, g428, g105}, g953);
	defparam lut_11605.LUT_SIZE = 6;
	defparam lut_11605.mask = 64'h0888808880008080;

	lut_sub lut_11622 ({g18, g97, g102, g578, g875}, g954);
	defparam lut_11622.LUT_SIZE = 5;
	defparam lut_11622.mask = 32'h0f070f0f;

	lut_sub lut_11643 ({g105, g500, g954}, g955);
	defparam lut_11643.LUT_SIZE = 3;
	defparam lut_11643.mask = 8'h8a;

	lut_sub lut_11655 ({g887, g790, g894, g952, g953, g955}, g956);
	defparam lut_11655.LUT_SIZE = 6;
	defparam lut_11655.mask = 64'h0000004000000000;

	lut_sub lut_11662 ({i_12_, i_13_, i_14_, g107, g91, g105}, g957);
	defparam lut_11662.LUT_SIZE = 6;
	defparam lut_11662.mask = 64'h88a000a0880088a0;

	lut_sub lut_11680 ({i_12_, i_13_, i_14_, g17, g27, g105}, g958);
	defparam lut_11680.LUT_SIZE = 6;
	defparam lut_11680.mask = 64'h2a2a0a2a0a2a0a22;

	lut_sub lut_11705 ({g957, g958}, g959);
	defparam lut_11705.LUT_SIZE = 2;
	defparam lut_11705.mask = 4'b1000;

	lut_sub lut_11714 ({g538, g111, g116, g548, g959}, g960);
	defparam lut_11714.LUT_SIZE = 5;
	defparam lut_11714.mask = 32'h00010000;

	lut_sub lut_11724 ({g936, g940, g942, g951, g956, g960}, g961);
	defparam lut_11724.LUT_SIZE = 6;
	defparam lut_11724.mask = 64'h0000000100000000;

	lut_sub lut_11730 ({i_8_, i_9_, i_10_, i_11_, g42, g394}, g962);
	defparam lut_11730.LUT_SIZE = 6;
	defparam lut_11730.mask = 64'h0110010001100110;

	lut_sub lut_11743 ({g926, g961, g962}, g963);
	defparam lut_11743.LUT_SIZE = 3;
	defparam lut_11743.mask = 8'h02;

	lut_sub lut_11751 ({g107, g176, g487, g652}, g964);
	defparam lut_11751.LUT_SIZE = 4;
	defparam lut_11751.mask = 16'h0888;

	lut_sub lut_11761 ({g83, g735, g738, g933}, g965);
	defparam lut_11761.LUT_SIZE = 4;
	defparam lut_11761.mask = 16'h4440;

	lut_sub lut_11770 ({g605, g761, g934}, g966);
	defparam lut_11770.LUT_SIZE = 3;
	defparam lut_11770.mask = 8'h10;

	lut_sub lut_11778 ({g489, g723, g851, g964}, g967);
	defparam lut_11778.LUT_SIZE = 4;
	defparam lut_11778.mask = 16'h1000;

	lut_sub lut_11787 ({g20, g735, g847, g966, g967}, g968);
	defparam lut_11787.LUT_SIZE = 5;
	defparam lut_11787.mask = 32'h01010100;

	lut_sub lut_11797 ({i_8_, g421, g964, g965, g968}, g969);
	defparam lut_11797.LUT_SIZE = 5;
	defparam lut_11797.mask = 32'h00ee00e0;

	lut_sub lut_11814 ({g164, g253, g468, g483, g855}, g970);
	defparam lut_11814.LUT_SIZE = 5;
	defparam lut_11814.mask = 32'h44554050;

	lut_sub lut_11828 ({g898, g945}, g971);
	defparam lut_11828.LUT_SIZE = 2;
	defparam lut_11828.mask = 4'b0001;

	lut_sub lut_11836 ({g421, g508, g725, g971}, g972);
	defparam lut_11836.LUT_SIZE = 4;
	defparam lut_11836.mask = 16'h00ef;

	lut_sub lut_11850 ({g253, g338, g484, g665}, g973);
	defparam lut_11850.LUT_SIZE = 4;
	defparam lut_11850.mask = 16'h7f00;

	lut_sub lut_11861 ({i_15_, i_12_, i_13_, i_14_, g112}, g974);
	defparam lut_11861.LUT_SIZE = 5;
	defparam lut_11861.mask = 32'h15454044;

	lut_sub lut_11876 ({g336, g627, g848}, g975);
	defparam lut_11876.LUT_SIZE = 3;
	defparam lut_11876.mask = 8'h04;

	lut_sub lut_11884 ({g164, g335, g597, g629}, g976);
	defparam lut_11884.LUT_SIZE = 4;
	defparam lut_11884.mask = 16'h007f;

	lut_sub lut_11898 ({g164, g974, g975, g976}, g977);
	defparam lut_11898.LUT_SIZE = 4;
	defparam lut_11898.mask = 16'haa20;

	lut_sub lut_11909 ({g333, g625, g865}, g978);
	defparam lut_11909.LUT_SIZE = 3;
	defparam lut_11909.mask = 8'h80;

	lut_sub lut_11919 ({g164, g334, g489, g624, g877, g875}, g979);
	defparam lut_11919.LUT_SIZE = 6;
	defparam lut_11919.mask = 64'h00000000fffff7ff;

	lut_sub lut_11958 ({g164, g948, g929, g978, g979}, g980);
	defparam lut_11958.LUT_SIZE = 5;
	defparam lut_11958.mask = 32'haaaa0002;

	lut_sub lut_11975 ({g972, g973, g676, g977, g980}, g981);
	defparam lut_11975.LUT_SIZE = 5;
	defparam lut_11975.mask = 32'h01000000;

	lut_sub lut_11984 ({g164, g253, g500, g624, g875}, g982);
	defparam lut_11984.LUT_SIZE = 5;
	defparam lut_11984.mask = 32'h22ff20f0;

	lut_sub lut_12003 ({i_15_, i_12_, i_13_, i_14_, g112}, g983);
	defparam lut_12003.LUT_SIZE = 5;
	defparam lut_12003.mask = 32'h40100401;

	lut_sub lut_12012 ({g113, g482}, g984);
	defparam lut_12012.LUT_SIZE = 2;
	defparam lut_12012.mask = 4'b0100;

	lut_sub lut_12021 ({g164, g253, g369, g664, g853}, g985);
	defparam lut_12021.LUT_SIZE = 5;
	defparam lut_12021.mask = 32'hc0ff80aa;

	lut_sub lut_12045 ({g164, g253, g984, g881, g852, g985}, g986);
	defparam lut_12045.LUT_SIZE = 6;
	defparam lut_12045.mask = 64'h5000555540004400;

	lut_sub lut_12064 ({g421, g983, g986}, g987);
	defparam lut_12064.LUT_SIZE = 3;
	defparam lut_12064.mask = 8'h54;

	lut_sub lut_12074 ({g346, g524, g982, g987}, g988);
	defparam lut_12074.LUT_SIZE = 4;
	defparam lut_12074.mask = 16'h0001;

	lut_sub lut_12082 ({g969, g970, g981, g988}, g989);
	defparam lut_12082.LUT_SIZE = 4;
	defparam lut_12082.mask = 16'h0100;

	lut_sub lut_12087 ({i_9_, i_10_, i_11_, g225}, g990);
	defparam lut_12087.LUT_SIZE = 4;
	defparam lut_12087.mask = 16'h0040;

	lut_sub lut_12093 ({g3, i_12_, i_13_, i_14_, g69}, g991);
	defparam lut_12093.LUT_SIZE = 5;
	defparam lut_12093.mask = 32'hbfba0c88;

	lut_sub lut_12116 ({g3, g227, g735, g927}, g992);
	defparam lut_12116.LUT_SIZE = 4;
	defparam lut_12116.mask = 16'h0507;

	lut_sub lut_12126 ({g17, g174}, g993);
	defparam lut_12126.LUT_SIZE = 2;
	defparam lut_12126.mask = 4'b0010;

	lut_sub lut_12133 ({g17, g27, g227}, g994);
	defparam lut_12133.LUT_SIZE = 3;
	defparam lut_12133.mask = 8'h15;

	lut_sub lut_12143 ({g226, g993, g725, g994}, g995);
	defparam lut_12143.LUT_SIZE = 4;
	defparam lut_12143.mask = 16'h20aa;

	lut_sub lut_12156 ({g3, g19, g68, g69, g226}, g996);
	defparam lut_12156.LUT_SIZE = 5;
	defparam lut_12156.mask = 32'h0022a0aa;

	lut_sub lut_12171 ({g227, g341, g655, g996}, g997);
	defparam lut_12171.LUT_SIZE = 4;
	defparam lut_12171.mask = 16'haa02;

	lut_sub lut_12183 ({g194, g213, g912, g997}, g998);
	defparam lut_12183.LUT_SIZE = 4;
	defparam lut_12183.mask = 16'h4440;

	lut_sub lut_12192 ({i_12_, i_13_, i_14_, g17, g27, g226}, g999);
	defparam lut_12192.LUT_SIZE = 6;
	defparam lut_12192.mask = 64'h0a2a002a0a0a0a22;

	lut_sub lut_12215 ({g213, g552, g469, g999}, g1000);
	defparam lut_12215.LUT_SIZE = 4;
	defparam lut_12215.mask = 16'haa02;

	lut_sub lut_12229 ({g226, g991, g992, g995, g998, g1000}, g1001);
	defparam lut_12229.LUT_SIZE = 6;
	defparam lut_12229.mask = 64'h0000010001000100;

	lut_sub lut_12235 ({i_9_, i_10_, i_11_, i_15_, i_13_, i_14_}, g1002);
	defparam lut_12235.LUT_SIZE = 6;
	defparam lut_12235.mask = 64'hf700000000000000;

	lut_sub lut_12251 ({g70, g121, g654, g990, g1001, g1002}, g1003);
	defparam lut_12251.LUT_SIZE = 6;
	defparam lut_12251.mask = 64'h3030200030300000;

	lut_sub lut_12265 ({g445, g142}, g1004);
	defparam lut_12265.LUT_SIZE = 2;
	defparam lut_12265.mask = 4'b0010;

	lut_sub lut_12272 ({g17, g27, g142}, g1005);
	defparam lut_12272.LUT_SIZE = 3;
	defparam lut_12272.mask = 8'h2a;

	lut_sub lut_12280 ({g428, g142}, g1006);
	defparam lut_12280.LUT_SIZE = 2;
	defparam lut_12280.mask = 4'b1000;

	lut_sub lut_12286 ({i_12_, i_13_, i_14_, g107, g91}, g1007);
	defparam lut_12286.LUT_SIZE = 5;
	defparam lut_12286.mask = 32'h51f15553;

	lut_sub lut_12310 ({g154, g984, g852, g853, g1007}, g1008);
	defparam lut_12310.LUT_SIZE = 5;
	defparam lut_12310.mask = 32'hbfff0000;

	lut_sub lut_12334 ({g159, g217, g984, g974, g983, g1008}, g1009);
	defparam lut_12334.LUT_SIZE = 6;
	defparam lut_12334.mask = 64'ha0008000aaaa8888;

	lut_sub lut_12357 ({g159, g154, g641, g849, g964}, g1010);
	defparam lut_12357.LUT_SIZE = 5;
	defparam lut_12357.mask = 32'h40c055ff;

	lut_sub lut_12380 ({g159, g975, g964, g1010, g1007}, g1011);
	defparam lut_12380.LUT_SIZE = 5;
	defparam lut_12380.mask = 32'h00013333;

	lut_sub lut_12396 ({g69, g154, g482, g743}, g1012);
	defparam lut_12396.LUT_SIZE = 4;
	defparam lut_12396.mask = 16'h5070;

	lut_sub lut_12408 ({g725, g929, g971, g1012}, g1013);
	defparam lut_12408.LUT_SIZE = 4;
	defparam lut_12408.mask = 16'h0002;

	lut_sub lut_12417 ({g154, g217, g974, g1013, g1455}, g1014);
	defparam lut_12417.LUT_SIZE = 5;
	defparam lut_12417.mask = 32'ha020aa22;

	lut_sub lut_12433 ({g335, g508, g629, g851}, g1015);
	defparam lut_12433.LUT_SIZE = 4;
	defparam lut_12433.mask = 16'h4000;

	lut_sub lut_12442 ({g159, g635, g932, g966, g1015}, g1016);
	defparam lut_12442.LUT_SIZE = 5;
	defparam lut_12442.mask = 32'hfeff0000;

	lut_sub lut_12466 ({g154, g875, g1016, g365, g632, g880}, g1017);
	defparam lut_12466.LUT_SIZE = 6;
	defparam lut_12466.mask = 64'h0100000001000100;

	lut_sub lut_12477 ({g600, g1009, g1011, g1014, g1017}, g1018);
	defparam lut_12477.LUT_SIZE = 5;
	defparam lut_12477.mask = 32'h00000001;

	lut_sub lut_12484 ({g357, g857, g948}, g1019);
	defparam lut_12484.LUT_SIZE = 3;
	defparam lut_12484.mask = 8'h40;

	lut_sub lut_12493 ({g125, g469, g720, g929, g1019}, g1020);
	defparam lut_12493.LUT_SIZE = 5;
	defparam lut_12493.mask = 32'h0000fffe;

	lut_sub lut_12512 ({i_15_, i_12_, i_13_, i_14_, g112}, g1021);
	defparam lut_12512.LUT_SIZE = 5;
	defparam lut_12512.mask = 32'h55550400;

	lut_sub lut_12526 ({i_12_, i_13_, i_14_, g144, g113}, g1022);
	defparam lut_12526.LUT_SIZE = 5;
	defparam lut_12526.mask = 32'h02000002;

	lut_sub lut_12535 ({g131, g197, g557, g664}, g1023);
	defparam lut_12535.LUT_SIZE = 4;
	defparam lut_12535.mask = 16'h7f00;

	lut_sub lut_12547 ({i_15_, i_12_, i_13_, i_14_, g125, g112}, g1024);
	defparam lut_12547.LUT_SIZE = 6;
	defparam lut_12547.mask = 64'h0111010000010100;

	lut_sub lut_12561 ({g131, g1021, g1022, g1023, g1024}, g1025);
	defparam lut_12561.LUT_SIZE = 5;
	defparam lut_12561.mask = 32'h80008080;

	lut_sub lut_12568 ({i_15_, i_12_, i_13_, i_14_, g112}, g1026);
	defparam lut_12568.LUT_SIZE = 5;
	defparam lut_12568.mask = 32'h00454044;

	lut_sub lut_12580 ({i_12_, i_13_, i_14_, g107, g91, g131}, g1027);
	defparam lut_12580.LUT_SIZE = 6;
	defparam lut_12580.mask = 64'h00a800a8008888a0;

	lut_sub lut_12598 ({g107, g460, g640}, g1028);
	defparam lut_12598.LUT_SIZE = 3;
	defparam lut_12598.mask = 8'h2a;

	lut_sub lut_12608 ({g4, g107, g176, g652}, g1029);
	defparam lut_12608.LUT_SIZE = 4;
	defparam lut_12608.mask = 16'h2a0a;

	lut_sub lut_12621 ({g125, g296, g651, g1028, g1029}, g1030);
	defparam lut_12621.LUT_SIZE = 5;
	defparam lut_12621.mask = 32'h0000efff;

	lut_sub lut_12643 ({g125, g1026, g1027, g1030}, g1031);
	defparam lut_12643.LUT_SIZE = 4;
	defparam lut_12643.mask = 16'h8880;

	lut_sub lut_12654 ({g20, g496, g522, g735, g847}, g1032);
	defparam lut_12654.LUT_SIZE = 5;
	defparam lut_12654.mask = 32'h50004000;

	lut_sub lut_12663 ({g508, g514, g852}, g1033);
	defparam lut_12663.LUT_SIZE = 3;
	defparam lut_12663.mask = 8'h80;

	lut_sub lut_12669 ({i_12_, i_14_, g88, g477}, g1034);
	defparam lut_12669.LUT_SIZE = 4;
	defparam lut_12669.mask = 16'haa8a;

	lut_sub lut_12682 ({i_12_, i_13_, i_14_, g20, g27, g91}, g1035);
	defparam lut_12682.LUT_SIZE = 6;
	defparam lut_12682.mask = 64'h0033bb3f330033bf;

	lut_sub lut_12721 ({g725, g1032, g1033, g1034, g1035}, g1036);
	defparam lut_12721.LUT_SIZE = 5;
	defparam lut_12721.mask = 32'h00000002;

	lut_sub lut_12727 ({i_12_, i_13_, i_14_, g86, g83}, g1037);
	defparam lut_12727.LUT_SIZE = 5;
	defparam lut_12727.mask = 32'h55050030;

	lut_sub lut_12742 ({g629, g703, g851, g1037}, g1038);
	defparam lut_12742.LUT_SIZE = 4;
	defparam lut_12742.mask = 16'h0200;

	lut_sub lut_12750 ({g25, g358, g933, g1038}, g1039);
	defparam lut_12750.LUT_SIZE = 4;
	defparam lut_12750.mask = 16'h0010;

	lut_sub lut_12758 ({i_8_, g144, g898, g1036, g1039}, g1040);
	defparam lut_12758.LUT_SIZE = 5;
	defparam lut_12758.mask = 32'h00ee00e0;

	lut_sub lut_12772 ({g761, g945}, g1041);
	defparam lut_12772.LUT_SIZE = 2;
	defparam lut_12772.mask = 4'b0001;

	lut_sub lut_12780 ({g125, g144, g851, g1041}, g1042);
	defparam lut_12780.LUT_SIZE = 4;
	defparam lut_12780.mask = 16'h0ace;

	lut_sub lut_12794 ({g317, g318, g319, g320}, g1043);
	defparam lut_12794.LUT_SIZE = 4;
	defparam lut_12794.mask = 16'h8000;

	lut_sub lut_12802 ({g355, g35, g460, g641}, g1044);
	defparam lut_12802.LUT_SIZE = 4;
	defparam lut_12802.mask = 16'ha2a0;

	lut_sub lut_12815 ({g125, g131, g487, g948, g1044}, g1045);
	defparam lut_12815.LUT_SIZE = 5;
	defparam lut_12815.mask = 32'h11ff10f0;

	lut_sub lut_12836 ({i_12_, i_13_, i_14_, g17, g27, g125}, g1046);
	defparam lut_12836.LUT_SIZE = 6;
	defparam lut_12836.mask = 64'h0515001505001511;

	lut_sub lut_12858 ({g125, g79, g625, g931}, g1047);
	defparam lut_12858.LUT_SIZE = 4;
	defparam lut_12858.mask = 16'h00f7;

	lut_sub lut_12871 ({i_12_, i_13_, i_14_, g35, g36, g125}, g1048);
	defparam lut_12871.LUT_SIZE = 6;
	defparam lut_12871.mask = 64'h1111001111000505;

	lut_sub lut_12888 ({i_15_, i_12_, i_13_, i_14_, g429, g125}, g1049);
	defparam lut_12888.LUT_SIZE = 6;
	defparam lut_12888.mask = 64'h1101011111111011;

	lut_sub lut_12909 ({g125, g282, g552, g668, g698}, g1050);
	defparam lut_12909.LUT_SIZE = 5;
	defparam lut_12909.mask = 32'h0000fbff;

	lut_sub lut_12932 ({g87, g131, g342, g1028, g1050}, g1051);
	defparam lut_12932.LUT_SIZE = 5;
	defparam lut_12932.mask = 32'h00aa20aa;

	lut_sub lut_12949 ({g1046, g1047, g1048, g1049, g1051}, g1052);
	defparam lut_12949.LUT_SIZE = 5;
	defparam lut_12949.mask = 32'h40000000;

	lut_sub lut_12959 ({g1042, g1043, g576, g577, g1045, g1052}, g1053);
	defparam lut_12959.LUT_SIZE = 6;
	defparam lut_12959.mask = 64'h0000010000000000;

	lut_sub lut_12965 ({i_15_, i_12_, i_13_, i_14_, g125, g445}, g1054);
	defparam lut_12965.LUT_SIZE = 6;
	defparam lut_12965.mask = 64'h0111111101010000;

	lut_sub lut_12982 ({g125, g504, g729, g643, g1054}, g1055);
	defparam lut_12982.LUT_SIZE = 5;
	defparam lut_12982.mask = 32'h88880008;

	lut_sub lut_12994 ({g211, g695, g797, g1055}, g1056);
	defparam lut_12994.LUT_SIZE = 4;
	defparam lut_12994.mask = 16'h0001;

	lut_sub lut_13004 ({g1020, g1025, g1031, g1040, g1053, g1056}, g1057);
	defparam lut_13004.LUT_SIZE = 6;
	defparam lut_13004.mask = 64'h0000001000000000;

	lut_sub lut_13010 ({g2, g12}, g1058);
	defparam lut_13010.LUT_SIZE = 2;
	defparam lut_13010.mask = 4'b0001;

	lut_sub lut_13015 ({i_4_, i_3_, i_5_, g1058}, o_19_);
	defparam lut_13015.LUT_SIZE = 4;
	defparam lut_13015.mask = 16'h0100;

	lut_sub lut_13019 ({i_4_, i_3_, i_5_}, g1060);
	defparam lut_13019.LUT_SIZE = 3;
	defparam lut_13019.mask = 8'h02;

	lut_sub lut_13025 ({g1058, g1060}, o_20_);
	defparam lut_13025.LUT_SIZE = 2;
	defparam lut_13025.mask = 4'b0001;

	lut_sub lut_13032 ({g6, g14, g101}, g1062);
	defparam lut_13032.LUT_SIZE = 3;
	defparam lut_13032.mask = 8'h01;

	lut_sub lut_13040 ({g18, g23, g28, g33}, g1063);
	defparam lut_13040.LUT_SIZE = 4;
	defparam lut_13040.mask = 16'h0800;

	lut_sub lut_13048 ({g20, g56, g1062, g1063}, g1064);
	defparam lut_13048.LUT_SIZE = 4;
	defparam lut_13048.mask = 16'h2223;

	lut_sub lut_13057 ({i_8_, i_7_, g48}, g1065);
	defparam lut_13057.LUT_SIZE = 3;
	defparam lut_13057.mask = 8'h04;

	lut_sub lut_13064 ({g55, g1064, g1065}, o_21_);
	defparam lut_13064.LUT_SIZE = 3;
	defparam lut_13064.mask = 8'h37;

	lut_sub lut_13075 ({g26, g28, g33}, g1067);
	defparam lut_13075.LUT_SIZE = 3;
	defparam lut_13075.mask = 8'h08;

	lut_sub lut_13082 ({g14, g62, g101}, g1068);
	defparam lut_13082.LUT_SIZE = 3;
	defparam lut_13082.mask = 8'h01;

	lut_sub lut_13088 ({i_8_, i_7_, g14, g62}, g1069);
	defparam lut_13088.LUT_SIZE = 4;
	defparam lut_13088.mask = 16'h1000;

	lut_sub lut_13096 ({g6, g14, g43, g1069}, g1070);
	defparam lut_13096.LUT_SIZE = 4;
	defparam lut_13096.mask = 16'haaa8;

	lut_sub lut_13110 ({g2, g16, g43, g1070}, g1071);
	defparam lut_13110.LUT_SIZE = 4;
	defparam lut_13110.mask = 16'h5450;

	lut_sub lut_13120 ({g1068, g1071}, g1072);
	defparam lut_13120.LUT_SIZE = 2;
	defparam lut_13120.mask = 4'b0100;

	lut_sub lut_13128 ({g26, g28, g1068, g1070}, g1073);
	defparam lut_13128.LUT_SIZE = 4;
	defparam lut_13128.mask = 16'h44f4;

	lut_sub lut_13140 ({g59, g65}, g1074);
	defparam lut_13140.LUT_SIZE = 2;
	defparam lut_13140.mask = 4'b0001;

	lut_sub lut_13146 ({i_0_, i_1_, g6, g15}, g1075);
	defparam lut_13146.LUT_SIZE = 4;
	defparam lut_13146.mask = 16'h0070;

	lut_sub lut_13158 ({g16, g28, g29, g43, g46, g1064}, g1076);
	defparam lut_13158.LUT_SIZE = 6;
	defparam lut_13158.mask = 64'h8888888800880080;

	lut_sub lut_13178 ({g33, g1072, g1073, g1074, g1075, g1076}, g1077);
	defparam lut_13178.LUT_SIZE = 6;
	defparam lut_13178.mask = 64'h0004000400000004;

	lut_sub lut_13186 ({i_4_, i_3_, g14, g42}, o_24_);
	defparam lut_13186.LUT_SIZE = 4;
	defparam lut_13186.mask = 16'h0001;

	lut_sub lut_13192 ({i_4_, i_3_, g10, g14}, o_25_);
	defparam lut_13192.LUT_SIZE = 4;
	defparam lut_13192.mask = 16'h0001;

	lut_sub lut_13199 ({g2, g43, g55}, g1080);
	defparam lut_13199.LUT_SIZE = 3;
	defparam lut_13199.mask = 8'h15;

	lut_sub lut_13208 ({g1062, g1072, g1080}, g1081);
	defparam lut_13208.LUT_SIZE = 3;
	defparam lut_13208.mask = 8'h20;

	lut_sub lut_13215 ({i_6_, i_7_, g14, g40, g1060}, g1082);
	defparam lut_13215.LUT_SIZE = 5;
	defparam lut_13215.mask = 32'h33053705;

	lut_sub lut_13236 ({g21, g23, g25, g1081, g1082}, o_26_);
	defparam lut_13236.LUT_SIZE = 5;
	defparam lut_13236.mask = 32'hddd5dddd;

	lut_sub lut_13264 ({g1, i_4_, i_3_, i_5_, g14}, g1084);
	defparam lut_13264.LUT_SIZE = 5;
	defparam lut_13264.mask = 32'h00010000;

	lut_sub lut_13273 ({g10, g18, g40, g457, g1081}, g1085);
	defparam lut_13273.LUT_SIZE = 5;
	defparam lut_13273.mask = 32'h00aa0fbf;

	lut_sub lut_13295 ({g33, g1062, g1072, g1080}, g1086);
	defparam lut_13295.LUT_SIZE = 4;
	defparam lut_13295.mask = 16'h00df;

	lut_sub lut_13307 ({i_4_, g40, g1075}, g1087);
	defparam lut_13307.LUT_SIZE = 3;
	defparam lut_13307.mask = 8'ha8;

	lut_sub lut_13319 ({g28, g45, g1062, g1072, g1080, g1087}, g1088);
	defparam lut_13319.LUT_SIZE = 6;
	defparam lut_13319.mask = 64'hffff55550c000400;

	lut_sub lut_13353 ({g1084, g1085, g1086, g1088}, o_27_);
	defparam lut_13353.LUT_SIZE = 4;
	defparam lut_13353.mask = 16'hbfff;

	lut_sub lut_13373 ({g1071, g1080}, g1090);
	defparam lut_13373.LUT_SIZE = 2;
	defparam lut_13373.mask = 4'b0010;

	lut_sub lut_13379 ({g1, g40}, g1091);
	defparam lut_13379.LUT_SIZE = 2;
	defparam lut_13379.mask = 4'b0001;

	lut_sub lut_13389 ({g23, g37, g1081, g1085, g1090, g1091}, o_28_);
	defparam lut_13389.LUT_SIZE = 6;
	defparam lut_13389.mask = 64'hffdfff5fdfdf5f5f;

	lut_sub lut_13452 ({g21, g634, g1081, g1086, g1090}, o_29_);
	defparam lut_13452.LUT_SIZE = 5;
	defparam lut_13452.mask = 32'hbb33fbf3;

	lut_sub lut_13481 ({g127, g74, g114}, g1094);
	defparam lut_13481.LUT_SIZE = 3;
	defparam lut_13481.mask = 8'h23;

	lut_sub lut_13490 ({i_12_, i_13_, i_14_, g107, g74, g91}, g1095);
	defparam lut_13490.LUT_SIZE = 6;
	defparam lut_13490.mask = 64'h0032003200222230;

	lut_sub lut_13508 ({i_12_, i_13_, i_14_, g75, g107, g91}, g1096);
	defparam lut_13508.LUT_SIZE = 6;
	defparam lut_13508.mask = 64'ha000c000e000c000;

	lut_sub lut_13522 ({i_15_, i_12_, i_13_, i_14_, g75, g112}, g1097);
	defparam lut_13522.LUT_SIZE = 6;
	defparam lut_13522.mask = 64'h0444404444044440;

	lut_sub lut_13539 ({i_15_, i_12_, i_13_, i_14_, g112, g74}, g1098);
	defparam lut_13539.LUT_SIZE = 6;
	defparam lut_13539.mask = 64'h0100101101010110;

	lut_sub lut_13556 ({g1094, g793, g1095, g1096, g1097, g1098}, g1099);
	defparam lut_13556.LUT_SIZE = 6;
	defparam lut_13556.mask = 64'h8000000000000000;

	lut_sub lut_13562 ({i_8_, g73, g358}, g1100);
	defparam lut_13562.LUT_SIZE = 3;
	defparam lut_13562.mask = 8'h10;

	lut_sub lut_13572 ({g1100, g670, g463, g464, g465, g466}, g1101);
	defparam lut_13572.LUT_SIZE = 6;
	defparam lut_13572.mask = 64'h8000000000000000;

	lut_sub lut_13577 ({i_15_, i_12_, i_13_, i_14_, g112}, g1102);
	defparam lut_13577.LUT_SIZE = 5;
	defparam lut_13577.mask = 32'h00100401;

	lut_sub lut_13586 ({g22, g174, g761}, g1103);
	defparam lut_13586.LUT_SIZE = 3;
	defparam lut_13586.mask = 8'h15;

	lut_sub lut_13595 ({i_8_, g73, g605, g635}, g1104);
	defparam lut_13595.LUT_SIZE = 4;
	defparam lut_13595.mask = 16'h0007;

	lut_sub lut_13604 ({i_8_, g73, g337, g851}, g1105);
	defparam lut_13604.LUT_SIZE = 4;
	defparam lut_13604.mask = 16'h000b;

	lut_sub lut_13616 ({g75, g949, g1102, g1103, g1104, g1105}, g1106);
	defparam lut_13616.LUT_SIZE = 6;
	defparam lut_13616.mask = 64'h0000080088888888;

	lut_sub lut_13631 ({g4, g27, g725}, g1107);
	defparam lut_13631.LUT_SIZE = 3;
	defparam lut_13631.mask = 8'h54;

	lut_sub lut_13640 ({i_8_, g4, g27, g73}, g1108);
	defparam lut_13640.LUT_SIZE = 4;
	defparam lut_13640.mask = 16'h0001;

	lut_sub lut_13650 ({g74, g847, g934, g1107, g1041, g1108}, g1109);
	defparam lut_13650.LUT_SIZE = 6;
	defparam lut_13650.mask = 64'haaaaaaaa00000002;

	lut_sub lut_13675 ({g102, g337, g605, g635, g858}, g1110);
	defparam lut_13675.LUT_SIZE = 5;
	defparam lut_13675.mask = 32'haaaa8000;

	lut_sub lut_13691 ({i_8_, g48, g73, g337, g605}, g1111);
	defparam lut_13691.LUT_SIZE = 5;
	defparam lut_13691.mask = 32'h0707000f;

	lut_sub lut_13708 ({g75, g725, g1029, g1111}, g1112);
	defparam lut_13708.LUT_SIZE = 4;
	defparam lut_13708.mask = 16'h02aa;

	lut_sub lut_13722 ({g1460, g1101, g1106, g1109, g1110, g1112}, g1113);
	defparam lut_13722.LUT_SIZE = 6;
	defparam lut_13722.mask = 64'h0000000000000001;

	lut_sub lut_13730 ({g496, g738, g1102, g1033}, g1114);
	defparam lut_13730.LUT_SIZE = 4;
	defparam lut_13730.mask = 16'h4000;

	lut_sub lut_13736 ({i_15_, i_12_, i_13_, i_14_, g75, g429}, g1115);
	defparam lut_13736.LUT_SIZE = 6;
	defparam lut_13736.mask = 64'h0404044444444044;

	lut_sub lut_13756 ({i_8_, g73, g993, g927, g1114, g1115}, g1116);
	defparam lut_13756.LUT_SIZE = 6;
	defparam lut_13756.mask = 64'haaaa2000aaaaa000;

	lut_sub lut_13784 ({g285, g589, g530, g1099, g1113, g1116}, g1117);
	defparam lut_13784.LUT_SIZE = 6;
	defparam lut_13784.mask = 64'h0000000000000001;

	lut_sub lut_13791 ({g24, g35, g1090}, g1118);
	defparam lut_13791.LUT_SIZE = 3;
	defparam lut_13791.mask = 8'h20;

	lut_sub lut_13801 ({g25, g42, g40, g1081, g1118, g1088}, g1119);
	defparam lut_13801.LUT_SIZE = 6;
	defparam lut_13801.mask = 64'h0404040044444400;

	lut_sub lut_13818 ({g100, g711, g961, g1117, g1119}, o_30_);
	defparam lut_13818.LUT_SIZE = 5;
	defparam lut_13818.mask = 32'hfffffffe;

	lut_sub lut_13853 ({i_6_, i_7_, i_4_, i_3_, i_5_, g14}, o_31_);
	defparam lut_13853.LUT_SIZE = 6;
	defparam lut_13853.mask = 64'h0001404000004045;

	lut_sub lut_13865 ({g1, i_4_, i_3_, i_5_, g14}, g1122);
	defparam lut_13865.LUT_SIZE = 5;
	defparam lut_13865.mask = 32'h00000001;

	lut_sub lut_13874 ({g43, g38, g55, g57, g1122}, g1123);
	defparam lut_13874.LUT_SIZE = 5;
	defparam lut_13874.mask = 32'h88888088;

	lut_sub lut_13889 ({g38, g1067, g1068, g1069, g1074}, g1124);
	defparam lut_13889.LUT_SIZE = 5;
	defparam lut_13889.mask = 32'h40444055;

	lut_sub lut_13906 ({g100, g711, g961, g1117, g1123, g1124}, g1125);
	defparam lut_13906.LUT_SIZE = 6;
	defparam lut_13906.mask = 64'h0000000000000001;

	lut_sub lut_13912 ({g38, g1067}, g1126);
	defparam lut_13912.LUT_SIZE = 2;
	defparam lut_13912.mask = 4'b0001;

	lut_sub lut_13920 ({g6, g14, g43, g1126}, g1127);
	defparam lut_13920.LUT_SIZE = 4;
	defparam lut_13920.mask = 16'h0002;

	lut_sub lut_13928 ({g44, g41, g1127, g1076}, g1128);
	defparam lut_13928.LUT_SIZE = 4;
	defparam lut_13928.mask = 16'h0400;

	lut_sub lut_13936 ({g100, g711, g961, g1117}, g1129);
	defparam lut_13936.LUT_SIZE = 4;
	defparam lut_13936.mask = 16'h0001;

	lut_sub lut_13944 ({i_8_, g73, g112, g636, g857}, g1130);
	defparam lut_13944.LUT_SIZE = 5;
	defparam lut_13944.mask = 32'h03030357;

	lut_sub lut_13962 ({g164, g154, g974, g1130}, g1131);
	defparam lut_13962.LUT_SIZE = 4;
	defparam lut_13962.mask = 16'h8a88;

	lut_sub lut_13974 ({g154, g106, g784, g964}, g1132);
	defparam lut_13974.LUT_SIZE = 4;
	defparam lut_13974.mask = 16'h40c0;

	lut_sub lut_13984 ({g123, g770, g629, g1132}, g1133);
	defparam lut_13984.LUT_SIZE = 4;
	defparam lut_13984.mask = 16'h4055;

	lut_sub lut_13996 ({g164, g123, g597, g628}, g1134);
	defparam lut_13996.LUT_SIZE = 4;
	defparam lut_13996.mask = 16'h30ba;

	lut_sub lut_14012 ({g75, g182, g183, g582, g976, g1134}, g1135);
	defparam lut_14012.LUT_SIZE = 6;
	defparam lut_14012.mask = 64'h8000000080808080;

	lut_sub lut_14024 ({g24, g75, g68, g83}, g1136);
	defparam lut_14024.LUT_SIZE = 4;
	defparam lut_14024.mask = 16'h5040;

	lut_sub lut_14032 ({i_8_, i_6_, i_7_, g445, g394}, g1137);
	defparam lut_14032.LUT_SIZE = 5;
	defparam lut_14032.mask = 32'h00000111;

	lut_sub lut_14042 ({g154, g597, g628, g629}, g1138);
	defparam lut_14042.LUT_SIZE = 4;
	defparam lut_14042.mask = 16'hdf00;

	lut_sub lut_14054 ({i_12_, i_13_, i_14_, g122, g83}, g1139);
	defparam lut_14054.LUT_SIZE = 5;
	defparam lut_14054.mask = 32'h01001001;

	lut_sub lut_14063 ({g123, g335, g850}, g1140);
	defparam lut_14063.LUT_SIZE = 3;
	defparam lut_14063.mask = 8'h70;

	lut_sub lut_14071 ({i_15_, i_12_, i_13_, i_14_, g445, g105}, g1141);
	defparam lut_14071.LUT_SIZE = 6;
	defparam lut_14071.mask = 64'h0220202222020222;

	lut_sub lut_14090 ({g1137, g1138, g1139, g1140, g1141}, g1142);
	defparam lut_14090.LUT_SIZE = 5;
	defparam lut_14090.mask = 32'h80000000;

	lut_sub lut_14098 ({g161, g125, g185, g182}, g1143);
	defparam lut_14098.LUT_SIZE = 4;
	defparam lut_14098.mask = 16'hf8a8;

	lut_sub lut_14113 ({g164, g154, g340, g850}, g1144);
	defparam lut_14113.LUT_SIZE = 4;
	defparam lut_14113.mask = 16'haf22;

	lut_sub lut_14128 ({g161, g122, g501, g543}, g1145);
	defparam lut_14128.LUT_SIZE = 4;
	defparam lut_14128.mask = 16'hf8a8;

	lut_sub lut_14143 ({g362, g1143, g1144, g1145}, g1146);
	defparam lut_14143.LUT_SIZE = 4;
	defparam lut_14143.mask = 16'h0100;

	lut_sub lut_14151 ({g75, g84, g699, g700}, g1147);
	defparam lut_14151.LUT_SIZE = 4;
	defparam lut_14151.mask = 16'h10f0;

	lut_sub lut_14164 ({g136, g1136, g1142, g1146, g1147}, g1148);
	defparam lut_14164.LUT_SIZE = 5;
	defparam lut_14164.mask = 32'h01000000;

	lut_sub lut_14170 ({g892, g608}, g1149);
	defparam lut_14170.LUT_SIZE = 2;
	defparam lut_14170.mask = 4'b0100;

	lut_sub lut_14179 ({g75, g105, g892, g473, g949}, g1150);
	defparam lut_14179.LUT_SIZE = 5;
	defparam lut_14179.mask = 32'h404055ff;

	lut_sub lut_14201 ({g161, g1149, g503, g1055, g1150}, g1151);
	defparam lut_14201.LUT_SIZE = 5;
	defparam lut_14201.mask = 32'h01010001;

	lut_sub lut_14212 ({g1131, g1133, g1135, g1148, g1151}, g1152);
	defparam lut_14212.LUT_SIZE = 5;
	defparam lut_14212.mask = 32'h00000001;

	lut_sub lut_14218 ({g1104, g1105}, g1153);
	defparam lut_14218.LUT_SIZE = 2;
	defparam lut_14218.mask = 4'b1000;

	lut_sub lut_14225 ({i_12_, i_13_, i_14_, g35, g36, g123}, g1154);
	defparam lut_14225.LUT_SIZE = 6;
	defparam lut_14225.mask = 64'h2a2a2a2a2a2a2a0a;

	lut_sub lut_14255 ({g125, g122, g186, g513}, g1155);
	defparam lut_14255.LUT_SIZE = 4;
	defparam lut_14255.mask = 16'hf4c4;

	lut_sub lut_14268 ({i_8_, i_6_, i_7_, g924, g394}, g1156);
	defparam lut_14268.LUT_SIZE = 5;
	defparam lut_14268.mask = 32'h00000110;

	lut_sub lut_14275 ({i_12_, i_13_, i_14_, g35, g105}, g1157);
	defparam lut_14275.LUT_SIZE = 5;
	defparam lut_14275.mask = 32'h02202022;

	lut_sub lut_14288 ({g164, g483, g641, g1156, g1157}, g1158);
	defparam lut_14288.LUT_SIZE = 5;
	defparam lut_14288.mask = 32'h88888000;

	lut_sub lut_14302 ({g161, g186, g192, g878, g1155, g1158}, g1159);
	defparam lut_14302.LUT_SIZE = 6;
	defparam lut_14302.mask = 64'h1010101010000000;

	lut_sub lut_14313 ({i_12_, i_13_, i_14_, g35, g36, g105}, g1160);
	defparam lut_14313.LUT_SIZE = 6;
	defparam lut_14313.mask = 64'h2222002a22222200;

	lut_sub lut_14334 ({g161, g122, g337, g851, g1160}, g1161);
	defparam lut_14334.LUT_SIZE = 5;
	defparam lut_14334.mask = 32'haa22a020;

	lut_sub lut_14351 ({g75, g192, g513, g514, g1161}, g1162);
	defparam lut_14351.LUT_SIZE = 5;
	defparam lut_14351.mask = 32'h04005555;

	lut_sub lut_14368 ({g634, g37, g75, g759, g710}, g1163);
	defparam lut_14368.LUT_SIZE = 5;
	defparam lut_14368.mask = 32'h02020222;

	lut_sub lut_14380 ({g164, g339, g849, g851}, g1164);
	defparam lut_14380.LUT_SIZE = 4;
	defparam lut_14380.mask = 16'h00bf;

	lut_sub lut_14394 ({i_8_, g35, g73, g68, g460}, g1165);
	defparam lut_14394.LUT_SIZE = 5;
	defparam lut_14394.mask = 32'h0000000e;

	lut_sub lut_14405 ({g30, g49, g118, g605, g514}, g1166);
	defparam lut_14405.LUT_SIZE = 5;
	defparam lut_14405.mask = 32'h0105030f;

	lut_sub lut_14418 ({i_8_, i_7_, i_12_, i_13_, i_14_, g36}, g1167);
	defparam lut_14418.LUT_SIZE = 6;
	defparam lut_14418.mask = 64'h0000000010010000;

	lut_sub lut_14428 ({i_8_, g73, g90, g186, g1166, g1167}, g1168);
	defparam lut_14428.LUT_SIZE = 6;
	defparam lut_14428.mask = 64'h1111111111111fff;

	lut_sub lut_14461 ({g634, g125, g281, g1165, g1168}, g1169);
	defparam lut_14461.LUT_SIZE = 5;
	defparam lut_14461.mask = 32'h88008880;

	lut_sub lut_14474 ({g125, g164, g122, g105, g948}, g1170);
	defparam lut_14474.LUT_SIZE = 5;
	defparam lut_14474.mask = 32'h8aaaaaaa;

	lut_sub lut_14497 ({g1455, g1048, g1164, g1169, g1170}, g1171);
	defparam lut_14497.LUT_SIZE = 5;
	defparam lut_14497.mask = 32'h20000000;

	lut_sub lut_14507 ({g1153, g1154, g1159, g1162, g1163, g1171}, g1172);
	defparam lut_14507.LUT_SIZE = 6;
	defparam lut_14507.mask = 64'h0000000000010000;

	lut_sub lut_14515 ({g125, g122, g648, g847}, g1173);
	defparam lut_14515.LUT_SIZE = 4;
	defparam lut_14515.mask = 16'hf4c4;

	lut_sub lut_14528 ({i_8_, i_6_, i_7_, g429, g394}, g1174);
	defparam lut_14528.LUT_SIZE = 5;
	defparam lut_14528.mask = 32'h00000110;

	lut_sub lut_14538 ({g68, g86, g125, g122, g460}, g1175);
	defparam lut_14538.LUT_SIZE = 5;
	defparam lut_14538.mask = 32'h003f0022;

	lut_sub lut_14554 ({g75, g273, g648, g1174, g1175}, g1176);
	defparam lut_14554.LUT_SIZE = 5;
	defparam lut_14554.mask = 32'h80008888;

	lut_sub lut_14567 ({g75, g125, g187, g1173, g1176}, g1177);
	defparam lut_14567.LUT_SIZE = 5;
	defparam lut_14567.mask = 32'h10101110;

	lut_sub lut_14577 ({i_15_, i_14_, g429, g122}, g1178);
	defparam lut_14577.LUT_SIZE = 4;
	defparam lut_14577.mask = 16'h0111;

	lut_sub lut_14585 ({i_15_, i_12_, i_13_, i_14_, g161, g429}, g1179);
	defparam lut_14585.LUT_SIZE = 6;
	defparam lut_14585.mask = 64'h0000001101010111;

	lut_sub lut_14601 ({g164, g105, g342, g522, g630, g847}, g1180);
	defparam lut_14601.LUT_SIZE = 6;
	defparam lut_14601.mask = 64'h4000ffff40004000;

	lut_sub lut_14625 ({g429, g123}, g1181);
	defparam lut_14625.LUT_SIZE = 2;
	defparam lut_14625.mask = 4'b0010;

	lut_sub lut_14633 ({g164, g975, g952, g1181}, g1182);
	defparam lut_14633.LUT_SIZE = 4;
	defparam lut_14633.mask = 16'h8808;

	lut_sub lut_14644 ({g1049, g1115, g1177, g1453, g1182}, g1183);
	defparam lut_14644.LUT_SIZE = 5;
	defparam lut_14644.mask = 32'h01000000;

	lut_sub lut_14651 ({g122, g487, g1029}, g1184);
	defparam lut_14651.LUT_SIZE = 3;
	defparam lut_14651.mask = 8'h0b;

	lut_sub lut_14660 ({i_14_, g107, g91, g123}, g1185);
	defparam lut_14660.LUT_SIZE = 4;
	defparam lut_14660.mask = 16'h88a8;

	lut_sub lut_14672 ({g105, g487, g484, g652}, g1186);
	defparam lut_14672.LUT_SIZE = 4;
	defparam lut_14672.mask = 16'h7f00;

	lut_sub lut_14687 ({g105, g358, g852, g1186, g1452}, g1187);
	defparam lut_14687.LUT_SIZE = 5;
	defparam lut_14687.mask = 32'h80008888;

	lut_sub lut_14701 ({g75, g122, g185, g486, g487, g708}, g1188);
	defparam lut_14701.LUT_SIZE = 6;
	defparam lut_14701.mask = 64'h80008000aaaaaa00;

	lut_sub lut_14723 ({g1184, g527, g1185, g1187, g1188}, g1189);
	defparam lut_14723.LUT_SIZE = 5;
	defparam lut_14723.mask = 32'h10000000;

	lut_sub lut_14731 ({g154, g334, g489, g624}, g1190);
	defparam lut_14731.LUT_SIZE = 4;
	defparam lut_14731.mask = 16'hfb00;

	lut_sub lut_14747 ({g18, g33, g97, g98, g122, g1190}, g1191);
	defparam lut_14747.LUT_SIZE = 6;
	defparam lut_14747.mask = 64'h88a8888888888888;

	lut_sub lut_14770 ({g105, g993, g1191}, g1192);
	defparam lut_14770.LUT_SIZE = 3;
	defparam lut_14770.mask = 8'h45;

	lut_sub lut_14779 ({i_8_, g73, g578, g461}, g1193);
	defparam lut_14779.LUT_SIZE = 4;
	defparam lut_14779.mask = 16'h0007;

	lut_sub lut_14790 ({g17, g76, g122, g91, g460}, g1194);
	defparam lut_14790.LUT_SIZE = 5;
	defparam lut_14790.mask = 32'h0c000f0a;

	lut_sub lut_14805 ({g28, g122, g180, g275}, g1195);
	defparam lut_14805.LUT_SIZE = 4;
	defparam lut_14805.mask = 16'h070f;

	lut_sub lut_14818 ({i_12_, i_13_, i_14_, g17, g27, g125}, g1196);
	defparam lut_14818.LUT_SIZE = 6;
	defparam lut_14818.mask = 64'h1100150011150000;

	lut_sub lut_14836 ({g276, g1193, g1194, g1195, g1196}, g1197);
	defparam lut_14836.LUT_SIZE = 5;
	defparam lut_14836.mask = 32'h80000000;

	lut_sub lut_14846 ({g164, g123, g334, g489, g624, g1107}, g1198);
	defparam lut_14846.LUT_SIZE = 6;
	defparam lut_14846.mask = 64'h0010ffff00100010;

	lut_sub lut_14871 ({i_12_, i_13_, i_14_, g17, g27, g86}, g1199);
	defparam lut_14871.LUT_SIZE = 6;
	defparam lut_14871.mask = 64'h770f000f0000000f;

	lut_sub lut_14898 ({g75, g97, g98, g725, g1029, g1199}, g1200);
	defparam lut_14898.LUT_SIZE = 6;
	defparam lut_14898.mask = 64'hfffffdff00000000;

	lut_sub lut_14937 ({g18, g33, g75, g1030, g1046}, g1201);
	defparam lut_14937.LUT_SIZE = 5;
	defparam lut_14937.mask = 32'h88080808;

	lut_sub lut_14951 ({g181, g1096, g1197, g1198, g1200, g1201}, g1202);
	defparam lut_14951.LUT_SIZE = 6;
	defparam lut_14951.mask = 64'h0004000000000000;

	lut_sub lut_14957 ({g461, g477}, g1203);
	defparam lut_14957.LUT_SIZE = 2;
	defparam lut_14957.mask = 4'b1000;

	lut_sub lut_14962 ({i_11_, i_15_, i_12_, i_13_, i_14_, g34}, g1204);
	defparam lut_14962.LUT_SIZE = 6;
	defparam lut_14962.mask = 64'h1545404411015044;

	lut_sub lut_14985 ({g179, g853, g1203, g1204}, g1205);
	defparam lut_14985.LUT_SIZE = 4;
	defparam lut_14985.mask = 16'h2000;

	lut_sub lut_14994 ({g154, g122, g1007, g1205, g999}, g1206);
	defparam lut_14994.LUT_SIZE = 5;
	defparam lut_14994.mask = 32'h0a02aa22;

	lut_sub lut_15012 ({g915, g959, g1189, g1192, g1202, g1206}, g1207);
	defparam lut_15012.LUT_SIZE = 6;
	defparam lut_15012.mask = 64'h0000000000000001;

	lut_sub lut_15018 ({g722, g203}, g1208);
	defparam lut_15018.LUT_SIZE = 2;
	defparam lut_15018.mask = 4'b0001;

	lut_sub lut_15025 ({i_8_, g73, g551, g495}, g1209);
	defparam lut_15025.LUT_SIZE = 4;
	defparam lut_15025.mask = 16'h000d;

	lut_sub lut_15035 ({g78, g122, g278, g551}, g1210);
	defparam lut_15035.LUT_SIZE = 4;
	defparam lut_15035.mask = 16'h0f0b;

	lut_sub lut_15049 ({g164, g154, g333, g343}, g1211);
	defparam lut_15049.LUT_SIZE = 4;
	defparam lut_15049.mask = 16'h4f45;

	lut_sub lut_15064 ({g21, g25, g125, g278}, g1212);
	defparam lut_15064.LUT_SIZE = 4;
	defparam lut_15064.mask = 16'h3133;

	lut_sub lut_15079 ({g154, g105, g521, g625, g626}, g1213);
	defparam lut_15079.LUT_SIZE = 5;
	defparam lut_15079.mask = 32'h8080f0ff;

	lut_sub lut_15101 ({g1209, g1210, g1211, g1212, g1213}, g1214);
	defparam lut_15101.LUT_SIZE = 5;
	defparam lut_15101.mask = 32'h04000000;

	lut_sub lut_15107 ({i_8_, i_6_, i_7_, g428, g394}, g1215);
	defparam lut_15107.LUT_SIZE = 5;
	defparam lut_15107.mask = 32'h00000444;

	lut_sub lut_15117 ({i_8_, g25, g73, g278, g1215}, g1216);
	defparam lut_15117.LUT_SIZE = 5;
	defparam lut_15117.mask = 32'haaaaa0a8;

	lut_sub lut_15138 ({g222, g207, g776, g783, g1216}, g1217);
	defparam lut_15138.LUT_SIZE = 5;
	defparam lut_15138.mask = 32'h40000000;

	lut_sub lut_15144 ({i_15_, i_12_, i_13_, i_14_, g428, g75}, g1218);
	defparam lut_15144.LUT_SIZE = 6;
	defparam lut_15144.mask = 64'h0088088888808808;

	lut_sub lut_15162 ({g125, g164, g551, g626}, g1219);
	defparam lut_15162.LUT_SIZE = 4;
	defparam lut_15162.mask = 16'h05cd;

	lut_sub lut_15178 ({g161, g164, g343, g452, g521, g1219}, g1220);
	defparam lut_15178.LUT_SIZE = 6;
	defparam lut_15178.mask = 64'ha0a0808000a00080;

	lut_sub lut_15195 ({g164, g154, g865, g978, g1047}, g1221);
	defparam lut_15195.LUT_SIZE = 5;
	defparam lut_15195.mask = 32'ha0aa2022;

	lut_sub lut_15209 ({i_15_, i_12_, i_13_, i_14_, g428, g123}, g1222);
	defparam lut_15209.LUT_SIZE = 6;
	defparam lut_15209.mask = 64'h0088808888080800;

	lut_sub lut_15223 ({g953, g1222}, g1223);
	defparam lut_15223.LUT_SIZE = 2;
	defparam lut_15223.mask = 4'b1000;

	lut_sub lut_15233 ({g1214, g1217, g1218, g1220, g1221, g1223}, g1224);
	defparam lut_15233.LUT_SIZE = 6;
	defparam lut_15233.mask = 64'h0000000000000100;

	lut_sub lut_15241 ({g3, g48, g119, g460}, g1225);
	defparam lut_15241.LUT_SIZE = 4;
	defparam lut_15241.mask = 16'hf0d0;

	lut_sub lut_15253 ({i_8_, i_3_, i_5_, g10, g71}, g1226);
	defparam lut_15253.LUT_SIZE = 5;
	defparam lut_15253.mask = 32'h00000100;

	lut_sub lut_15262 ({g3, g75, g460, g927, g1226}, g1227);
	defparam lut_15262.LUT_SIZE = 5;
	defparam lut_15262.mask = 32'h55115551;

	lut_sub lut_15283 ({g468, g608, g927, g1225, g1227}, g1228);
	defparam lut_15283.LUT_SIZE = 5;
	defparam lut_15283.mask = 32'h55455555;

	lut_sub lut_15305 ({g69, g113, g105, g482}, g1229);
	defparam lut_15305.LUT_SIZE = 4;
	defparam lut_15305.mask = 16'h4044;

	lut_sub lut_15317 ({g355, g126, g122, g182, g460, g552}, g1230);
	defparam lut_15317.LUT_SIZE = 6;
	defparam lut_15317.mask = 64'h00ef00af00ff00af;

	lut_sub lut_15352 ({g75, g282, g270, g585, g1230}, g1231);
	defparam lut_15352.LUT_SIZE = 5;
	defparam lut_15352.mask = 32'h80008888;

	lut_sub lut_15365 ({g105, g1229, g877, g857, g1231}, g1232);
	defparam lut_15365.LUT_SIZE = 5;
	defparam lut_15365.mask = 32'h40005500;

	lut_sub lut_15375 ({i_15_, i_12_, i_13_, i_14_, g75, g112}, g1233);
	defparam lut_15375.LUT_SIZE = 6;
	defparam lut_15375.mask = 64'h0404044444444044;

	lut_sub lut_15396 ({g125, g154, g688, g877, g929, g1012}, g1234);
	defparam lut_15396.LUT_SIZE = 6;
	defparam lut_15396.mask = 64'h2020aaaa2000aa00;

	lut_sub lut_15418 ({g5, g17, g69, g174}, g1235);
	defparam lut_15418.LUT_SIZE = 4;
	defparam lut_15418.mask = 16'hd500;

	lut_sub lut_15431 ({g226, g469, g508, g725, g1235}, g1236);
	defparam lut_15431.LUT_SIZE = 5;
	defparam lut_15431.mask = 32'hffef0000;

	lut_sub lut_15454 ({g164, g341, g742, g655, g1236}, g1237);
	defparam lut_15454.LUT_SIZE = 5;
	defparam lut_15454.mask = 32'haaaa0002;

	lut_sub lut_15469 ({g341, g469, g927}, g1238);
	defparam lut_15469.LUT_SIZE = 3;
	defparam lut_15469.mask = 8'h02;

	lut_sub lut_15479 ({g347, g121, g725, g945, g983, g1238}, g1239);
	defparam lut_15479.LUT_SIZE = 6;
	defparam lut_15479.mask = 64'h000c0004ffff5555;

	lut_sub lut_15514 ({g290, g1233, g1234, g1237, g1239}, g1240);
	defparam lut_15514.LUT_SIZE = 5;
	defparam lut_15514.mask = 32'h00000100;

	lut_sub lut_15522 ({g24, g113, g174, g857}, g1241);
	defparam lut_15522.LUT_SIZE = 4;
	defparam lut_15522.mask = 16'h0a2a;

	lut_sub lut_15535 ({g383, g469, g928, g971, g1241}, g1242);
	defparam lut_15535.LUT_SIZE = 5;
	defparam lut_15535.mask = 32'hfffe0000;

	lut_sub lut_15557 ({g77, g105, g927, g945}, g1243);
	defparam lut_15557.LUT_SIZE = 4;
	defparam lut_15557.mask = 16'hb0f0;

	lut_sub lut_15571 ({g125, g205, g761, g1243}, g1244);
	defparam lut_15571.LUT_SIZE = 4;
	defparam lut_15571.mask = 16'ha020;

	lut_sub lut_15580 ({g3, i_12_, i_13_, i_14_, g75, g69}, g1245);
	defparam lut_15580.LUT_SIZE = 6;
	defparam lut_15580.mask = 64'h4000440040cc44cc;

	lut_sub lut_15603 ({g944, g1242, g129, g391, g1244, g1245}, g1246);
	defparam lut_15603.LUT_SIZE = 6;
	defparam lut_15603.mask = 64'h0000000000020000;

	lut_sub lut_15611 ({i_15_, g125, g112, g122, g460}, g1247);
	defparam lut_15611.LUT_SIZE = 5;
	defparam lut_15611.mask = 32'h000a0202;

	lut_sub lut_15619 ({i_15_, i_12_, i_13_, i_14_, g428}, g1248);
	defparam lut_15619.LUT_SIZE = 5;
	defparam lut_15619.mask = 32'h20200888;

	lut_sub lut_15630 ({g123, g1248, g974}, g1249);
	defparam lut_15630.LUT_SIZE = 3;
	defparam lut_15630.mask = 8'h70;

	lut_sub lut_15642 ({g164, g347, g557, g898, g1247, g1249}, g1250);
	defparam lut_15642.LUT_SIZE = 6;
	defparam lut_15642.mask = 64'h0808888808008800;

	lut_sub lut_15660 ({g122, g933, g559, g532, g1457, g1250}, g1251);
	defparam lut_15660.LUT_SIZE = 6;
	defparam lut_15660.mask = 64'h0001000100000001;

	lut_sub lut_15672 ({g1224, g1228, g1232, g1240, g1246, g1251}, g1252);
	defparam lut_15672.LUT_SIZE = 6;
	defparam lut_15672.mask = 64'h0000000000010000;

	lut_sub lut_15682 ({g1152, g1172, g1183, g1207, g1208, g1252}, g1253);
	defparam lut_15682.LUT_SIZE = 6;
	defparam lut_15682.mask = 64'h0000000000000001;

	lut_sub lut_15689 ({i_12_, i_13_, i_14_, g107, g91, g130}, g1254);
	defparam lut_15689.LUT_SIZE = 6;
	defparam lut_15689.mask = 64'h88a8a0a8a8a8a8a0;

	lut_sub lut_15715 ({i_12_, i_13_, i_14_, g107, g102}, g1255);
	defparam lut_15715.LUT_SIZE = 5;
	defparam lut_15715.mask = 32'h04444040;

	lut_sub lut_15727 ({i_8_, g73, g107, g176, g460}, g1256);
	defparam lut_15727.LUT_SIZE = 5;
	defparam lut_15727.mask = 32'h00e00000;

	lut_sub lut_15735 ({i_12_, i_13_, i_14_, g102, g91}, g1257);
	defparam lut_15735.LUT_SIZE = 5;
	defparam lut_15735.mask = 32'h20002020;

	lut_sub lut_15746 ({g159, g253, g852, g853, g964}, g1258);
	defparam lut_15746.LUT_SIZE = 5;
	defparam lut_15746.mask = 32'h40c040ff;

	lut_sub lut_15765 ({g1255, g1256, g1257, g1258}, g1259);
	defparam lut_15765.LUT_SIZE = 4;
	defparam lut_15765.mask = 16'h4000;

	lut_sub lut_15771 ({g130, g652}, g1260);
	defparam lut_15771.LUT_SIZE = 2;
	defparam lut_15771.mask = 4'b0100;

	lut_sub lut_15778 ({i_8_, g4, g73, g91}, g1261);
	defparam lut_15778.LUT_SIZE = 4;
	defparam lut_15778.mask = 16'h0200;

	lut_sub lut_15786 ({g135, g131, g296, g651}, g1262);
	defparam lut_15786.LUT_SIZE = 4;
	defparam lut_15786.mask = 16'h888f;

	lut_sub lut_15801 ({i_8_, g19, g73, g107, g68, g91}, g1263);
	defparam lut_15801.LUT_SIZE = 6;
	defparam lut_15801.mask = 64'h00c800fa00000000;

	lut_sub lut_15819 ({g131, g1028, g1260, g1261, g1262, g1263}, g1264);
	defparam lut_15819.LUT_SIZE = 6;
	defparam lut_15819.mask = 64'h0000200020002000;

	lut_sub lut_15828 ({i_11_, g34, g101, g394}, g1265);
	defparam lut_15828.LUT_SIZE = 4;
	defparam lut_15828.mask = 16'h0001;

	lut_sub lut_15838 ({g131, g348, g487, g852, g964, g1265}, g1266);
	defparam lut_15838.LUT_SIZE = 6;
	defparam lut_15838.mask = 64'h20002020a000aaaa;

	lut_sub lut_15856 ({i_12_, i_13_, i_14_, g107, g91}, g1267);
	defparam lut_15856.LUT_SIZE = 5;
	defparam lut_15856.mask = 32'hae0ca0ec;

	lut_sub lut_15877 ({g135, g562, g1029, g1267}, g1268);
	defparam lut_15877.LUT_SIZE = 4;
	defparam lut_15877.mask = 16'hdf00;

	lut_sub lut_15891 ({g159, g964, g1007, g1268}, g1269);
	defparam lut_15891.LUT_SIZE = 4;
	defparam lut_15891.mask = 16'h02aa;

	lut_sub lut_15905 ({g973, g1254, g1259, g1264, g1266, g1269}, g1270);
	defparam lut_15905.LUT_SIZE = 6;
	defparam lut_15905.mask = 64'h0001000000000000;

	lut_sub lut_15911 ({i_4_, i_3_, i_5_, g43, g71}, g1271);
	defparam lut_15911.LUT_SIZE = 5;
	defparam lut_15911.mask = 32'h01001100;

	lut_sub lut_15921 ({i_15_, g429, g74, g460, g1271}, g1272);
	defparam lut_15921.LUT_SIZE = 5;
	defparam lut_15921.mask = 32'h004c0000;

	lut_sub lut_15929 ({i_12_, i_14_, g88, g130}, g1273);
	defparam lut_15929.LUT_SIZE = 4;
	defparam lut_15929.mask = 16'h0020;

	lut_sub lut_15937 ({g135, g648, g703, g775}, g1274);
	defparam lut_15937.LUT_SIZE = 4;
	defparam lut_15937.mask = 16'h20aa;

	lut_sub lut_15950 ({g74, g104, g847, g1273, g1274}, g1275);
	defparam lut_15950.LUT_SIZE = 5;
	defparam lut_15950.mask = 32'h44000400;

	lut_sub lut_15960 ({g313, g348, g496, g535}, g1276);
	defparam lut_15960.LUT_SIZE = 4;
	defparam lut_15960.mask = 16'h8a88;

	lut_sub lut_15972 ({g413, g522, g847, g1276}, g1277);
	defparam lut_15972.LUT_SIZE = 4;
	defparam lut_15972.mask = 16'h1055;

	lut_sub lut_15983 ({g135, g191, g187}, g1278);
	defparam lut_15983.LUT_SIZE = 3;
	defparam lut_15983.mask = 8'h70;

	lut_sub lut_15993 ({g102, g534, g500, g703}, g1279);
	defparam lut_15993.LUT_SIZE = 4;
	defparam lut_15993.mask = 16'h00bf;

	lut_sub lut_16006 ({g135, g89, g630}, g1280);
	defparam lut_16006.LUT_SIZE = 3;
	defparam lut_16006.mask = 8'hd0;

	lut_sub lut_16014 ({i_12_, i_13_, i_14_, g86, g102}, g1281);
	defparam lut_16014.LUT_SIZE = 5;
	defparam lut_16014.mask = 32'h01101011;

	lut_sub lut_16024 ({i_15_, i_12_, i_13_, i_14_, g429, g131}, g1282);
	defparam lut_16024.LUT_SIZE = 6;
	defparam lut_16024.mask = 64'h0222200020222020;

	lut_sub lut_16041 ({g1278, g1279, g1280, g1281, g1282}, g1283);
	defparam lut_16041.LUT_SIZE = 5;
	defparam lut_16041.mask = 32'h80000000;

	lut_sub lut_16049 ({g135, g131, g273, g342}, g1284);
	defparam lut_16049.LUT_SIZE = 4;
	defparam lut_16049.mask = 16'h88af;

	lut_sub lut_16066 ({g159, g253, g336, g500, g627, g848}, g1285);
	defparam lut_16066.LUT_SIZE = 6;
	defparam lut_16066.mask = 64'h0040f0f00040ffff;

	lut_sub lut_16099 ({g274, g584, g1284, g1285}, g1286);
	defparam lut_16099.LUT_SIZE = 4;
	defparam lut_16099.mask = 16'h1000;

	lut_sub lut_16105 ({i_15_, i_12_, i_13_, i_14_, g429, g130}, g1287);
	defparam lut_16105.LUT_SIZE = 6;
	defparam lut_16105.mask = 64'h0222222220220200;

	lut_sub lut_16124 ({g76, g157, g135, g88, g176}, g1288);
	defparam lut_16124.LUT_SIZE = 5;
	defparam lut_16124.mask = 32'h30330022;

	lut_sub lut_16137 ({i_8_, i_6_, i_7_, g429, g394}, g1289);
	defparam lut_16137.LUT_SIZE = 5;
	defparam lut_16137.mask = 32'h01110000;

	lut_sub lut_16147 ({g206, g1287, g1288, g1289}, g1290);
	defparam lut_16147.LUT_SIZE = 4;
	defparam lut_16147.mask = 16'h8000;

	lut_sub lut_16153 ({i_15_, i_12_, i_13_, i_14_, g429, g74}, g1291);
	defparam lut_16153.LUT_SIZE = 6;
	defparam lut_16153.mask = 64'h0011010110101101;

	lut_sub lut_16169 ({g102, g253, g342, g630}, g1292);
	defparam lut_16169.LUT_SIZE = 4;
	defparam lut_16169.mask = 16'h8f88;

	lut_sub lut_16184 ({g159, g847, g934, g975, g1292}, g1293);
	defparam lut_16184.LUT_SIZE = 5;
	defparam lut_16184.mask = 32'h00015555;

	lut_sub lut_16201 ({g1283, g1286, g1290, g1291, g1293}, g1294);
	defparam lut_16201.LUT_SIZE = 5;
	defparam lut_16201.mask = 32'h00000004;

	lut_sub lut_16210 ({g1270, g1272, g1275, g1277, g1294}, g1295);
	defparam lut_16210.LUT_SIZE = 5;
	defparam lut_16210.mask = 32'h00000100;

	lut_sub lut_16217 ({i_12_, i_13_, i_14_, g35, g36, g130}, g1296);
	defparam lut_16217.LUT_SIZE = 6;
	defparam lut_16217.mask = 64'h220a0a2a2a222a0a;

	lut_sub lut_16245 ({g135, g130, g337, g635, g851, g1296}, g1297);
	defparam lut_16245.LUT_SIZE = 6;
	defparam lut_16245.mask = 64'h2000a0002000aaaa;

	lut_sub lut_16264 ({g157, g135, g186, g337}, g1298);
	defparam lut_16264.LUT_SIZE = 4;
	defparam lut_16264.mask = 16'h3075;

	lut_sub lut_16277 ({g109, g90, g102}, g1299);
	defparam lut_16277.LUT_SIZE = 3;
	defparam lut_16277.mask = 8'h15;

	lut_sub lut_16286 ({g35, g157, g460}, g1300);
	defparam lut_16286.LUT_SIZE = 3;
	defparam lut_16286.mask = 8'hc4;

	lut_sub lut_16294 ({i_12_, i_14_, g35, g72}, g1301);
	defparam lut_16294.LUT_SIZE = 4;
	defparam lut_16294.mask = 16'h0010;

	lut_sub lut_16299 ({i_8_, i_6_, i_7_, g1301}, g1302);
	defparam lut_16299.LUT_SIZE = 4;
	defparam lut_16299.mask = 16'h1400;

	lut_sub lut_16309 ({g74, g1299, g281, g1300, g1302}, g1303);
	defparam lut_16309.LUT_SIZE = 5;
	defparam lut_16309.mask = 32'hfb00bb00;

	lut_sub lut_16331 ({g74, g313, g253, g851, g1298, g1303}, g1304);
	defparam lut_16331.LUT_SIZE = 6;
	defparam lut_16331.mask = 64'h0444040404040404;

	lut_sub lut_16347 ({g253, g337, g339, g849}, g1305);
	defparam lut_16347.LUT_SIZE = 4;
	defparam lut_16347.mask = 16'h7f00;

	lut_sub lut_16361 ({g37, g102, g555, g483}, g1306);
	defparam lut_16361.LUT_SIZE = 4;
	defparam lut_16361.mask = 16'h0f07;

	lut_sub lut_16373 ({i_12_, i_13_, i_14_, g35, g102}, g1307);
	defparam lut_16373.LUT_SIZE = 5;
	defparam lut_16373.mask = 32'h01101011;

	lut_sub lut_16386 ({g634, g135, g131, g281, g513}, g1308);
	defparam lut_16386.LUT_SIZE = 5;
	defparam lut_16386.mask = 32'h000f444f;

	lut_sub lut_16404 ({g1305, g1306, g1307, g1308}, g1309);
	defparam lut_16404.LUT_SIZE = 4;
	defparam lut_16404.mask = 16'h4000;

	lut_sub lut_16411 ({i_12_, i_13_, i_14_, g35, g36, g159}, g1310);
	defparam lut_16411.LUT_SIZE = 6;
	defparam lut_16411.mask = 64'h0a2a222a002a002a;

	lut_sub lut_16436 ({g90, g74, g281, g513, g635, g1310}, g1311);
	defparam lut_16436.LUT_SIZE = 6;
	defparam lut_16436.mask = 64'haaaa0800aaaa0000;

	lut_sub lut_16461 ({g673, g926, g1045, g1309, g1311}, g1312);
	defparam lut_16461.LUT_SIZE = 5;
	defparam lut_16461.mask = 32'h00010000;

	lut_sub lut_16468 ({i_12_, i_13_, i_14_, g35, g36, g74}, g1313);
	defparam lut_16468.LUT_SIZE = 6;
	defparam lut_16468.mask = 64'h1105050500111105;

	lut_sub lut_16489 ({g35, g339, g460, g641}, g1314);
	defparam lut_16489.LUT_SIZE = 4;
	defparam lut_16489.mask = 16'ha020;

	lut_sub lut_16497 ({i_8_, i_7_, g924, g394}, g1315);
	defparam lut_16497.LUT_SIZE = 4;
	defparam lut_16497.mask = 16'h0100;

	lut_sub lut_16505 ({g135, g1314, g1315, g204}, g1316);
	defparam lut_16505.LUT_SIZE = 4;
	defparam lut_16505.mask = 16'h0444;

	lut_sub lut_16515 ({g313, g348, g514, g746}, g1317);
	defparam lut_16515.LUT_SIZE = 4;
	defparam lut_16515.mask = 16'h4544;

	lut_sub lut_16528 ({g257, g605, g1313, g1316, g1317}, g1318);
	defparam lut_16528.LUT_SIZE = 5;
	defparam lut_16528.mask = 32'h10101000;

	lut_sub lut_16540 ({g1010, g506, g1297, g1304, g1312, g1318}, g1319);
	defparam lut_16540.LUT_SIZE = 6;
	defparam lut_16540.mask = 64'h0000000000000001;

	lut_sub lut_16546 ({i_14_, g27, g102}, g1320);
	defparam lut_16546.LUT_SIZE = 3;
	defparam lut_16546.mask = 8'h01;

	lut_sub lut_16554 ({g17, g76, g135, g460}, g1321);
	defparam lut_16554.LUT_SIZE = 4;
	defparam lut_16554.mask = 16'h00c8;

	lut_sub lut_16564 ({g159, g253, g334, g875}, g1322);
	defparam lut_16564.LUT_SIZE = 4;
	defparam lut_16564.mask = 16'h223f;

	lut_sub lut_16580 ({g135, g185, g180, g1321, g1322}, g1323);
	defparam lut_16580.LUT_SIZE = 5;
	defparam lut_16580.mask = 32'h40004444;

	lut_sub lut_16593 ({g74, g180, g461, g1320, g1323}, g1324);
	defparam lut_16593.LUT_SIZE = 5;
	defparam lut_16593.mask = 32'h44444000;

	lut_sub lut_16604 ({g28, g135, g275}, g1325);
	defparam lut_16604.LUT_SIZE = 3;
	defparam lut_16604.mask = 8'h4c;

	lut_sub lut_16612 ({i_12_, i_13_, i_14_, g17, g102}, g1326);
	defparam lut_16612.LUT_SIZE = 5;
	defparam lut_16612.mask = 32'h01110101;

	lut_sub lut_16623 ({i_8_, g73, g578, g993}, g1327);
	defparam lut_16623.LUT_SIZE = 4;
	defparam lut_16623.mask = 16'h0700;

	lut_sub lut_16632 ({i_12_, i_13_, i_14_, g17, g159, g131}, g1328);
	defparam lut_16632.LUT_SIZE = 6;
	defparam lut_16632.mask = 64'h0e0c000e0e0e0e00;

	lut_sub lut_16657 ({g1325, g277, g1326, g1327, g1328}, g1329);
	defparam lut_16657.LUT_SIZE = 5;
	defparam lut_16657.mask = 32'h80000000;

	lut_sub lut_16667 ({g74, g402, g337, g605, g993, g1107}, g1330);
	defparam lut_16667.LUT_SIZE = 6;
	defparam lut_16667.mask = 64'h4444ffff40005000;

	lut_sub lut_16697 ({g130, g131, g334, g875}, g1331);
	defparam lut_16697.LUT_SIZE = 4;
	defparam lut_16697.mask = 16'h222f;

	lut_sub lut_16712 ({g18, g33, g74, g1331, g937}, g1332);
	defparam lut_16712.LUT_SIZE = 5;
	defparam lut_16712.mask = 32'h22202020;

	lut_sub lut_16725 ({g1095, g1005, g1329, g1330, g1332}, g1333);
	defparam lut_16725.LUT_SIZE = 5;
	defparam lut_16725.mask = 32'h01000000;

	lut_sub lut_16732 ({g97, g98, g135}, g1334);
	defparam lut_16732.LUT_SIZE = 3;
	defparam lut_16732.mask = 8'ha2;

	lut_sub lut_16741 ({g102, g212, g484}, g1335);
	defparam lut_16741.LUT_SIZE = 3;
	defparam lut_16741.mask = 8'h07;

	lut_sub lut_16749 ({i_4_, i_3_, i_5_, g71, g101}, g1336);
	defparam lut_16749.LUT_SIZE = 5;
	defparam lut_16749.mask = 32'h10000100;

	lut_sub lut_16755 ({i_9_, i_10_, i_11_, g1336}, g1337);
	defparam lut_16755.LUT_SIZE = 4;
	defparam lut_16755.mask = 16'h0040;

	lut_sub lut_16763 ({g4, g27, g394, g1337}, g1338);
	defparam lut_16763.LUT_SIZE = 4;
	defparam lut_16763.mask = 16'h1115;

	lut_sub lut_16776 ({g18, g33, g135, g130, g624}, g1339);
	defparam lut_16776.LUT_SIZE = 5;
	defparam lut_16776.mask = 32'h77070707;

	lut_sub lut_16800 ({g1334, g383, g993, g1335, g1338, g1339}, g1340);
	defparam lut_16800.LUT_SIZE = 6;
	defparam lut_16800.mask = 64'h4000404000000000;

	lut_sub lut_16810 ({g179, g461, g605, g487}, g1341);
	defparam lut_16810.LUT_SIZE = 4;
	defparam lut_16810.mask = 16'h8000;

	lut_sub lut_16819 ({g135, g313, g477, g1341, g990}, g1342);
	defparam lut_16819.LUT_SIZE = 5;
	defparam lut_16819.mask = 32'h2220aaa0;

	lut_sub lut_16836 ({g97, g98, g74, g257, g489}, g1343);
	defparam lut_16836.LUT_SIZE = 5;
	defparam lut_16836.mask = 32'he0e0eae0;

	lut_sub lut_16858 ({g1027, g995, g1340, g1342, g1343}, g1344);
	defparam lut_16858.LUT_SIZE = 5;
	defparam lut_16858.mask = 32'h00010000;

	lut_sub lut_16867 ({g955, g982, g1324, g1333, g1344}, g1345);
	defparam lut_16867.LUT_SIZE = 5;
	defparam lut_16867.mask = 32'h00000001;

	lut_sub lut_16877 ({g1172, g1183, g1207, g1295, g1319, g1345}, g1346);
	defparam lut_16877.LUT_SIZE = 6;
	defparam lut_16877.mask = 64'h0000000000000001;

	lut_sub lut_16884 ({g123, g852, g853}, g1347);
	defparam lut_16884.LUT_SIZE = 3;
	defparam lut_16884.mask = 8'h70;

	lut_sub lut_16894 ({g113, g174, g408, g857}, g1348);
	defparam lut_16894.LUT_SIZE = 4;
	defparam lut_16894.mask = 16'hc444;

	lut_sub lut_16904 ({i_15_, i_12_, i_13_, i_14_, g112, g123}, g1349);
	defparam lut_16904.LUT_SIZE = 6;
	defparam lut_16904.mask = 64'h0000020000220200;

	lut_sub lut_16916 ({g130, g742, g1347, g1348, g1349}, g1350);
	defparam lut_16916.LUT_SIZE = 5;
	defparam lut_16916.mask = 32'h00808080;

	lut_sub lut_16927 ({g123, g113, g130, g507, g974}, g1351);
	defparam lut_16927.LUT_SIZE = 5;
	defparam lut_16927.mask = 32'h75557050;

	lut_sub lut_16949 ({g24, g113, g408, g1350, g1351}, g1352);
	defparam lut_16949.LUT_SIZE = 5;
	defparam lut_16949.mask = 32'h02222222;

	lut_sub lut_16961 ({i_15_, i_12_, i_13_, i_14_, g73, g112}, g1353);
	defparam lut_16961.LUT_SIZE = 6;
	defparam lut_16961.mask = 64'h0505050005155555;

	lut_sub lut_16987 ({g10, g72, g101, g1102}, g1354);
	defparam lut_16987.LUT_SIZE = 4;
	defparam lut_16987.mask = 16'h0307;

	lut_sub lut_16999 ({i_8_, g73, g125, g857, g1029}, g1355);
	defparam lut_16999.LUT_SIZE = 5;
	defparam lut_16999.mask = 32'h033303ab;

	lut_sub lut_17021 ({g102, g200, g212, g484, g684, g881}, g1356);
	defparam lut_17021.LUT_SIZE = 6;
	defparam lut_17021.mask = 64'h00000000dfffffff;

	lut_sub lut_17060 ({g105, g984, g943, g957, g1356}, g1357);
	defparam lut_17060.LUT_SIZE = 5;
	defparam lut_17060.mask = 32'h80008080;

	lut_sub lut_17071 ({g940, g1353, g1354, g1355, g1357}, g1358);
	defparam lut_17071.LUT_SIZE = 5;
	defparam lut_17071.mask = 32'h00004440;

	lut_sub lut_17078 ({i_15_, i_12_, i_13_, i_14_, g112}, g1359);
	defparam lut_17078.LUT_SIZE = 5;
	defparam lut_17078.mask = 32'h15455154;

	lut_sub lut_17094 ({i_15_, i_12_, i_13_, i_14_, g112}, g1360);
	defparam lut_17094.LUT_SIZE = 5;
	defparam lut_17094.mask = 32'h11041004;

	lut_sub lut_17106 ({i_8_, g107, g735, g1267, g1360}, g1361);
	defparam lut_17106.LUT_SIZE = 5;
	defparam lut_17106.mask = 32'h00008088;

	lut_sub lut_17116 ({i_8_, g165, g487, g1359, g1361}, g1362);
	defparam lut_17116.LUT_SIZE = 5;
	defparam lut_17116.mask = 32'h002a00aa;

	lut_sub lut_17130 ({g135, g122, g185, g562}, g1363);
	defparam lut_17130.LUT_SIZE = 4;
	defparam lut_17130.mask = 16'h3705;

	lut_sub lut_17146 ({g165, g122, g114, g286, g557, g983}, g1364);
	defparam lut_17146.LUT_SIZE = 6;
	defparam lut_17146.mask = 64'hffff00c0aaaa0080;

	lut_sub lut_17182 ({g122, g197, g200, g715, g1363, g1364}, g1365);
	defparam lut_17182.LUT_SIZE = 6;
	defparam lut_17182.mask = 64'h4040404040000000;

	lut_sub lut_17194 ({g1025, g1031, g1362, g1365}, g1366);
	defparam lut_17194.LUT_SIZE = 4;
	defparam lut_17194.mask = 16'h0004;

	lut_sub lut_17204 ({g1184, g527, g1009, g1185, g1187, g1188}, g1367);
	defparam lut_17204.LUT_SIZE = 6;
	defparam lut_17204.mask = 64'h0010000000000000;

	lut_sub lut_17214 ({g987, g1099, g1352, g1358, g1366, g1367}, g1368);
	defparam lut_17214.LUT_SIZE = 6;
	defparam lut_17214.mask = 64'h0000000000000001;

	lut_sub lut_17223 ({g165, g122, g343, g626, g945}, g1369);
	defparam lut_17223.LUT_SIZE = 5;
	defparam lut_17223.mask = 32'hff0c5504;

	lut_sub lut_17245 ({g135, g605, g761, g1369}, g1370);
	defparam lut_17245.LUT_SIZE = 4;
	defparam lut_17245.mask = 16'h1055;

	lut_sub lut_17257 ({g159, g253, g333, g865}, g1371);
	defparam lut_17257.LUT_SIZE = 4;
	defparam lut_17257.mask = 16'h88cf;

	lut_sub lut_17272 ({g20, g24, g74, g460}, g1372);
	defparam lut_17272.LUT_SIZE = 4;
	defparam lut_17272.mask = 16'h0032;

	lut_sub lut_17280 ({i_12_, i_13_, i_14_, g22, g102}, g1373);
	defparam lut_17280.LUT_SIZE = 5;
	defparam lut_17280.mask = 32'h40044040;

	lut_sub lut_17291 ({g257, g313, g278, g333}, g1374);
	defparam lut_17291.LUT_SIZE = 4;
	defparam lut_17291.mask = 16'hf8c8;

	lut_sub lut_17308 ({g122, g1314, g1371, g1372, g1373, g1374}, g1375);
	defparam lut_17308.LUT_SIZE = 6;
	defparam lut_17308.mask = 64'h0040004000000040;

	lut_sub lut_17318 ({g125, g159, g521, g642}, g1376);
	defparam lut_17318.LUT_SIZE = 4;
	defparam lut_17318.mask = 16'h3075;

	lut_sub lut_17334 ({g23, g157, g130, g175, g449, g1376}, g1377);
	defparam lut_17334.LUT_SIZE = 6;
	defparam lut_17334.mask = 64'h00aa0022a0aa2022;

	lut_sub lut_17357 ({g165, g257, g738, g777, g1377}, g1378);
	defparam lut_17357.LUT_SIZE = 5;
	defparam lut_17357.mask = 32'h55504440;

	lut_sub lut_17374 ({g425, g408, g945, g1248, g1111}, g1379);
	defparam lut_17374.LUT_SIZE = 5;
	defparam lut_17374.mask = 32'h080a88aa;

	lut_sub lut_17390 ({g74, g521, g1041, g388}, g1380);
	defparam lut_17390.LUT_SIZE = 4;
	defparam lut_17390.mask = 16'haa20;

	lut_sub lut_17403 ({g1370, g1375, g1378, g1379, g1380}, g1381);
	defparam lut_17403.LUT_SIZE = 5;
	defparam lut_17403.mask = 32'h00000001;

	lut_sub lut_17409 ({i_8_, i_6_, g120, g761}, g1382);
	defparam lut_17409.LUT_SIZE = 4;
	defparam lut_17409.mask = 16'h2000;

	lut_sub lut_17418 ({g21, g23, g74, g495, g1382}, g1383);
	defparam lut_17418.LUT_SIZE = 5;
	defparam lut_17418.mask = 32'ha0a8a0a0;

	lut_sub lut_17433 ({g78, g74, g79}, g1384);
	defparam lut_17433.LUT_SIZE = 3;
	defparam lut_17433.mask = 8'h32;

	lut_sub lut_17442 ({g74, g175, g278}, g1385);
	defparam lut_17442.LUT_SIZE = 3;
	defparam lut_17442.mask = 8'h07;

	lut_sub lut_17452 ({g159, g131, g253, g625}, g1386);
	defparam lut_17452.LUT_SIZE = 4;
	defparam lut_17452.mask = 16'h5554;

	lut_sub lut_17464 ({i_8_, i_6_, i_7_, g428, g394}, g1387);
	defparam lut_17464.LUT_SIZE = 5;
	defparam lut_17464.mask = 32'h04400000;

	lut_sub lut_17474 ({g25, g102, g79, g278, g1387}, g1388);
	defparam lut_17474.LUT_SIZE = 5;
	defparam lut_17474.mask = 32'haa00aa08;

	lut_sub lut_17491 ({g131, g177, g551, g1386, g1388}, g1389);
	defparam lut_17491.LUT_SIZE = 5;
	defparam lut_17491.mask = 32'h04004444;

	lut_sub lut_17503 ({g21, g122, g413, g931}, g1390);
	defparam lut_17503.LUT_SIZE = 4;
	defparam lut_17503.mask = 16'hba32;

	lut_sub lut_17520 ({g1384, g238, g1131, g1385, g1389, g1390}, g1391);
	defparam lut_17520.LUT_SIZE = 6;
	defparam lut_17520.mask = 64'h0010000000000000;

	lut_sub lut_17530 ({g1042, g1467, g1006, g1270, g1383, g1391}, g1392);
	defparam lut_17530.LUT_SIZE = 6;
	defparam lut_17530.mask = 64'h0000010000000000;

	lut_sub lut_17540 ({g1172, g1224, g1319, g1368, g1381, g1392}, g1393);
	defparam lut_17540.LUT_SIZE = 6;
	defparam lut_17540.mask = 64'h0000000000000001;

	lut_sub lut_17548 ({g74, g182, g183, g699}, g1394);
	defparam lut_17548.LUT_SIZE = 4;
	defparam lut_17548.mask = 16'h00bf;

	lut_sub lut_17563 ({g355, g83, g356, g629, g1394}, g1395);
	defparam lut_17563.LUT_SIZE = 5;
	defparam lut_17563.mask = 32'ha8a8a8a0;

	lut_sub lut_17580 ({g102, g699, g700}, g1396);
	defparam lut_17580.LUT_SIZE = 3;
	defparam lut_17580.mask = 8'h0e;

	lut_sub lut_17589 ({g24, g74, g445}, g1397);
	defparam lut_17589.LUT_SIZE = 3;
	defparam lut_17589.mask = 8'h10;

	lut_sub lut_17597 ({g24, g68, g102, g83}, g1398);
	defparam lut_17597.LUT_SIZE = 4;
	defparam lut_17597.mask = 16'h1110;

	lut_sub lut_17606 ({g102, g501, g543}, g1399);
	defparam lut_17606.LUT_SIZE = 3;
	defparam lut_17606.mask = 8'h07;

	lut_sub lut_17616 ({i_8_, g19, g73, g76, g83}, g1400);
	defparam lut_17616.LUT_SIZE = 5;
	defparam lut_17616.mask = 32'h04050000;

	lut_sub lut_17624 ({i_8_, i_6_, i_7_, g445, g394}, g1401);
	defparam lut_17624.LUT_SIZE = 5;
	defparam lut_17624.mask = 32'h01100000;

	lut_sub lut_17633 ({i_8_, g73, g82, g295, g1401}, g1402);
	defparam lut_17633.LUT_SIZE = 5;
	defparam lut_17633.mask = 32'haa80aaaa;

	lut_sub lut_17654 ({g1398, g1399, g583, g1400, g1402}, g1403);
	defparam lut_17654.LUT_SIZE = 5;
	defparam lut_17654.mask = 32'h40000000;

	lut_sub lut_17663 ({g131, g182, g183, g295, g700}, g1404);
	defparam lut_17663.LUT_SIZE = 5;
	defparam lut_17663.mask = 32'hbfff0000;

	lut_sub lut_17687 ({g157, g74, g183, g892, g608, g1404}, g1405);
	defparam lut_17687.LUT_SIZE = 6;
	defparam lut_17687.mask = 64'haaaaa0a020002000;

	lut_sub lut_17709 ({g159, g214, g438, g770, g930}, g1406);
	defparam lut_17709.LUT_SIZE = 5;
	defparam lut_17709.mask = 32'h4c004f00;

	lut_sub lut_17725 ({g1396, g1397, g1403, g1405, g1406}, g1407);
	defparam lut_17725.LUT_SIZE = 5;
	defparam lut_17725.mask = 32'h01000000;

	lut_sub lut_17731 ({i_15_, i_12_, i_13_, i_14_, g445, g130}, g1408);
	defparam lut_17731.LUT_SIZE = 6;
	defparam lut_17731.mask = 64'h0202000220022220;

	lut_sub lut_17746 ({g157, g131, g501, g543}, g1409);
	defparam lut_17746.LUT_SIZE = 4;
	defparam lut_17746.mask = 16'h5073;

	lut_sub lut_17762 ({g157, g159, g253, g335, g597, g850}, g1410);
	defparam lut_17762.LUT_SIZE = 6;
	defparam lut_17762.mask = 64'h8088f0ff8088c0cc;

	lut_sub lut_17794 ({g103, g253, g237, g629, g1410}, g1411);
	defparam lut_17794.LUT_SIZE = 5;
	defparam lut_17794.mask = 32'h40500000;

	lut_sub lut_17802 ({i_4_, i_3_, i_5_, g83, g735}, g1412);
	defparam lut_17802.LUT_SIZE = 5;
	defparam lut_17802.mask = 32'h01001000;

	lut_sub lut_17812 ({g2, g54, g71, g723, g1412}, g1413);
	defparam lut_17812.LUT_SIZE = 5;
	defparam lut_17812.mask = 32'h00000407;

	lut_sub lut_17824 ({g102, g350, g608, g898, g1413}, g1414);
	defparam lut_17824.LUT_SIZE = 5;
	defparam lut_17824.mask = 32'haa020202;

	lut_sub lut_17839 ({g774, g1408, g1409, g1411, g1414}, g1415);
	defparam lut_17839.LUT_SIZE = 5;
	defparam lut_17839.mask = 32'h10000000;

	lut_sub lut_17848 ({g1460, g1004, g1395, g1407, g1415}, g1416);
	defparam lut_17848.LUT_SIZE = 5;
	defparam lut_17848.mask = 32'h00000100;

	lut_sub lut_17857 ({g1152, g1183, g1295, g1368, g1416}, g1417);
	defparam lut_17857.LUT_SIZE = 5;
	defparam lut_17857.mask = 32'h00000001;

	lut_sub lut_17867 ({g109, g161, g392, g569, g1149, g374}, g1418);
	defparam lut_17867.LUT_SIZE = 6;
	defparam lut_17867.mask = 64'h5010501050100000;

	lut_sub lut_17881 ({i_15_, i_12_, i_13_, i_14_, g429, g445}, g1419);
	defparam lut_17881.LUT_SIZE = 6;
	defparam lut_17881.mask = 64'h0000003707050573;

	lut_sub lut_17905 ({g24, g35, g36, g68}, g1420);
	defparam lut_17905.LUT_SIZE = 4;
	defparam lut_17905.mask = 16'hd0d5;

	lut_sub lut_17921 ({g157, g343, g502, g1419, g1420}, g1421);
	defparam lut_17921.LUT_SIZE = 5;
	defparam lut_17921.mask = 32'hf0f00040;

	lut_sub lut_17938 ({g250, g454, g1179, g1418, g1421}, g1422);
	defparam lut_17938.LUT_SIZE = 5;
	defparam lut_17938.mask = 32'h00000010;

	lut_sub lut_17946 ({g5, g16, g30, g49}, g1423);
	defparam lut_17946.LUT_SIZE = 4;
	defparam lut_17946.mask = 16'h0007;

	lut_sub lut_17957 ({g2, g14, g62, g1126, g1423}, g1424);
	defparam lut_17957.LUT_SIZE = 5;
	defparam lut_17957.mask = 32'haaaaaaa2;

	lut_sub lut_17978 ({g80, i_11_, g7, g101}, o_41_);
	defparam lut_17978.LUT_SIZE = 4;
	defparam lut_17978.mask = 16'h0010;

	lut_sub lut_17984 ({g395, g1459}, g1426);
	defparam lut_17984.LUT_SIZE = 2;
	defparam lut_17984.mask = 4'b1000;

	lut_sub lut_17990 ({g774, g779}, g1427);
	defparam lut_17990.LUT_SIZE = 2;
	defparam lut_17990.mask = 4'b0100;

	lut_sub lut_18000 ({g135, g299, g342, g681, g301, g302}, g1428);
	defparam lut_18000.LUT_SIZE = 6;
	defparam lut_18000.mask = 64'h1000000010100000;

	lut_sub lut_18010 ({g122, g948, g1184, g1268}, g1429);
	defparam lut_18010.LUT_SIZE = 4;
	defparam lut_18010.mask = 16'h8808;

	lut_sub lut_18018 ({g122, g898}, g1430);
	defparam lut_18018.LUT_SIZE = 2;
	defparam lut_18018.mask = 4'b0010;

	lut_sub lut_18028 ({g221, g222, g1430, g223, g224, g1178}, g1431);
	defparam lut_18028.LUT_SIZE = 6;
	defparam lut_18028.mask = 64'h0200000000000000;

	lut_sub lut_18038 ({g637, g138, g1554, g862, g1429, g1431}, g1432);
	defparam lut_18038.LUT_SIZE = 6;
	defparam lut_18038.mask = 64'h0000000100000000;

	lut_sub lut_18046 ({i_8_, g333, g898, g1015, g1032}, g1433);
	defparam lut_18046.LUT_SIZE = 5;
	defparam lut_18046.mask = 32'hfeff0000;

	lut_sub lut_18068 ({g514, g725, g641, g1203}, g1434);
	defparam lut_18068.LUT_SIZE = 4;
	defparam lut_18068.mask = 16'h0400;

	lut_sub lut_18078 ({g165, g933, g1433, g1434, g1362, g1365}, g1435);
	defparam lut_18078.LUT_SIZE = 6;
	defparam lut_18078.mask = 64'h4444444400000400;

	lut_sub lut_18096 ({g1427, g787, g1370, g1428, g1432, g1435}, g1436);
	defparam lut_18096.LUT_SIZE = 6;
	defparam lut_18096.mask = 64'h0000000000000001;

	lut_sub lut_18105 ({g135, g337, g635, g1001, g1436}, g1437);
	defparam lut_18105.LUT_SIZE = 5;
	defparam lut_18105.mask = 32'h10001111;

	lut_sub lut_18118 ({g17, g23, g507, g624, g1036}, g1438);
	defparam lut_18118.LUT_SIZE = 5;
	defparam lut_18118.mask = 32'h00110010;

	lut_sub lut_18129 ({g408, g605, g971, g1248, g1181}, g1439);
	defparam lut_18129.LUT_SIZE = 5;
	defparam lut_18129.mask = 32'h0800aaaa;

	lut_sub lut_18146 ({g130, g965, g1438, g1185, g1439}, g1440);
	defparam lut_18146.LUT_SIZE = 5;
	defparam lut_18146.mask = 32'h00044444;

	lut_sub lut_18157 ({g123, g850, g1154}, g1441);
	defparam lut_18157.LUT_SIZE = 3;
	defparam lut_18157.mask = 8'h8a;

	lut_sub lut_18167 ({g597, g489, g624, g629}, g1442);
	defparam lut_18167.LUT_SIZE = 4;
	defparam lut_18167.mask = 16'h2000;

	lut_sub lut_18176 ({g70, g335, g468, g770, g877}, g1443);
	defparam lut_18176.LUT_SIZE = 5;
	defparam lut_18176.mask = 32'h80000000;

	lut_sub lut_18185 ({g334, g875, g928, g1442, g1443}, g1444);
	defparam lut_18185.LUT_SIZE = 5;
	defparam lut_18185.mask = 32'h00000100;

	lut_sub lut_18193 ({g123, g552, g511, g654}, g1445);
	defparam lut_18193.LUT_SIZE = 4;
	defparam lut_18193.mask = 16'hf700;

	lut_sub lut_18208 ({g77, g123, g270, g1287, g1445}, g1446);
	defparam lut_18208.LUT_SIZE = 5;
	defparam lut_18208.mask = 32'h80880088;

	lut_sub lut_18222 ({g123, g198, g1107, g1444, g1222, g1446}, g1447);
	defparam lut_18222.LUT_SIZE = 6;
	defparam lut_18222.mask = 64'h0004000044440000;

	lut_sub lut_18235 ({g1254, g1352, g1408, g1441, g1447}, g1448);
	defparam lut_18235.LUT_SIZE = 5;
	defparam lut_18235.mask = 32'h00100000;

	lut_sub lut_18244 ({g1456, g1297, g1436, g1440, g1448}, g1449);
	defparam lut_18244.LUT_SIZE = 5;
	defparam lut_18244.mask = 32'h00000001;

	lut_sub lut_18253 ({g2, g16, g43, g38, g1070}, g1450);
	defparam lut_18253.LUT_SIZE = 5;
	defparam lut_18253.mask = 32'h888c88cc;

	lut_sub lut_18273 ({g100, g711, g961, g1117, g1123, g1450}, g1451);
	defparam lut_18273.LUT_SIZE = 6;
	defparam lut_18273.mask = 64'h0000000000000002;

	lut_sub lut_18280 ({g91, g107, i_14_, g164}, g1452);
	defparam lut_18280.LUT_SIZE = 4;
	defparam lut_18280.mask = 16'h5510;

	lut_sub lut_18294 ({g88, g154, g86, g1180, g1179, g1178}, g1453);
	defparam lut_18294.LUT_SIZE = 6;
	defparam lut_18294.mask = 64'h0800080800000808;

	lut_sub lut_18306 ({g48, i_7_, i_8_, g1068, g1067, g16}, g1454);
	defparam lut_18306.LUT_SIZE = 6;
	defparam lut_18306.mask = 64'hf3f3f3f3f3a2f3f3;

	lut_sub lut_18357 ({g36, g35, i_14_, g154}, g1455);
	defparam lut_18357.LUT_SIZE = 4;
	defparam lut_18357.mask = 16'h02aa;

	lut_sub lut_18367 ({i_10_, i_9_, g118, g10, i_8_, i_11_}, g1456);
	defparam lut_18367.LUT_SIZE = 6;
	defparam lut_18367.mask = 64'hfff9fff7fff7ffff;

	lut_sub lut_18434 ({i_14_, g682, g681, g226, g69}, g1457);
	defparam lut_18434.LUT_SIZE = 5;
	defparam lut_18434.mask = 32'h00b000f0;

	lut_sub lut_18450 ({g605, g73, g606, g604, g603, g602}, g1458);
	defparam lut_18450.LUT_SIZE = 6;
	defparam lut_18450.mask = 64'h8000800080000000;

	lut_sub lut_18458 ({g71, g15, i_7_, i_6_, i_11_, i_10_}, g1459);
	defparam lut_18458.LUT_SIZE = 6;
	defparam lut_18458.mask = 64'h0000000000000220;

	lut_sub lut_18465 ({g73, g1461}, g1460);
	defparam lut_18465.LUT_SIZE = 2;
	defparam lut_18465.mask = 4'b0010;

	lut_sub lut_18471 ({g73, g1462}, g1461);
	defparam lut_18471.LUT_SIZE = 2;
	defparam lut_18471.mask = 4'b0001;

	lut_sub lut_18477 ({g1463, g1464}, g1462);
	defparam lut_18477.LUT_SIZE = 2;
	defparam lut_18477.mask = 4'b1000;

	lut_sub lut_18482 ({i_8_, g1465}, g1463);
	defparam lut_18482.LUT_SIZE = 2;
	defparam lut_18482.mask = 4'b0100;

	lut_sub lut_18487 ({i_8_, g1466}, g1464);
	defparam lut_18487.LUT_SIZE = 2;
	defparam lut_18487.mask = 4'b0001;

	lut_sub lut_18495 ({g628, g608, g898, g340}, g1465);
	defparam lut_18495.LUT_SIZE = 4;
	defparam lut_18495.mask = 16'h0001;

	lut_sub lut_18501 ({g608, g847}, g1466);
	defparam lut_18501.LUT_SIZE = 2;
	defparam lut_18501.mask = 4'b0001;

	lut_sub lut_18507 ({g1468, g1469}, g1467);
	defparam lut_18507.LUT_SIZE = 2;
	defparam lut_18507.mask = 4'b1000;

	lut_sub lut_18513 ({g168, g1470}, g1468);
	defparam lut_18513.LUT_SIZE = 2;
	defparam lut_18513.mask = 4'b0100;

	lut_sub lut_18519 ({g168, g1472}, g1469);
	defparam lut_18519.LUT_SIZE = 2;
	defparam lut_18519.mask = 4'b0001;

	lut_sub lut_18525 ({g105, g1471}, g1470);
	defparam lut_18525.LUT_SIZE = 2;
	defparam lut_18525.mask = 4'b1000;

	lut_sub lut_18531 ({g105, g1475}, g1471);
	defparam lut_18531.LUT_SIZE = 2;
	defparam lut_18531.mask = 4'b0100;

	lut_sub lut_18537 ({g1473, g1474}, g1472);
	defparam lut_18537.LUT_SIZE = 2;
	defparam lut_18537.mask = 4'b1000;

	lut_sub lut_18543 ({g105, g1476}, g1473);
	defparam lut_18543.LUT_SIZE = 2;
	defparam lut_18543.mask = 4'b0100;

	lut_sub lut_18549 ({g105, g1477}, g1474);
	defparam lut_18549.LUT_SIZE = 2;
	defparam lut_18549.mask = 4'b0001;

	lut_sub lut_18556 ({g626, g343, g851}, g1475);
	defparam lut_18556.LUT_SIZE = 3;
	defparam lut_18556.mask = 8'h10;

	lut_sub lut_18564 ({g626, g343, g851, g945}, g1476);
	defparam lut_18564.LUT_SIZE = 4;
	defparam lut_18564.mask = 16'h0100;

	lut_sub lut_18572 ({g626, g343, g102, g945}, g1477);
	defparam lut_18572.LUT_SIZE = 4;
	defparam lut_18572.mask = 16'h4544;

	lut_sub lut_18582 ({g1479, g1480}, g1478);
	defparam lut_18582.LUT_SIZE = 2;
	defparam lut_18582.mask = 4'b1000;

	lut_sub lut_18588 ({g23, g1481}, g1479);
	defparam lut_18588.LUT_SIZE = 2;
	defparam lut_18588.mask = 4'b0100;

	lut_sub lut_18594 ({g23, g1482}, g1480);
	defparam lut_18594.LUT_SIZE = 2;
	defparam lut_18594.mask = 4'b0001;

	lut_sub lut_18600 ({g142, g1485}, g1481);
	defparam lut_18600.LUT_SIZE = 2;
	defparam lut_18600.mask = 4'b0001;

	lut_sub lut_18606 ({g1483, g1484}, g1482);
	defparam lut_18606.LUT_SIZE = 2;
	defparam lut_18606.mask = 4'b1000;

	lut_sub lut_18612 ({g142, g1486}, g1483);
	defparam lut_18612.LUT_SIZE = 2;
	defparam lut_18612.mask = 4'b0100;

	lut_sub lut_18618 ({g142, g1487}, g1484);
	defparam lut_18618.LUT_SIZE = 2;
	defparam lut_18618.mask = 4'b0001;

	lut_sub lut_18626 ({g703, g518, g154, g896}, g1485);
	defparam lut_18626.LUT_SIZE = 4;
	defparam lut_18626.mask = 16'h1011;

	lut_sub lut_18636 ({g703, g518, g25, g896}, g1486);
	defparam lut_18636.LUT_SIZE = 4;
	defparam lut_18636.mask = 16'h1011;

	lut_sub lut_18645 ({g703, g518, g896}, g1487);
	defparam lut_18645.LUT_SIZE = 3;
	defparam lut_18645.mask = 8'h45;

	lut_sub lut_18653 ({g1489, g1490}, g1488);
	defparam lut_18653.LUT_SIZE = 2;
	defparam lut_18653.mask = 4'b1000;

	lut_sub lut_18659 ({g130, g1491}, g1489);
	defparam lut_18659.LUT_SIZE = 2;
	defparam lut_18659.mask = 4'b0100;

	lut_sub lut_18665 ({g130, g1494}, g1490);
	defparam lut_18665.LUT_SIZE = 2;
	defparam lut_18665.mask = 4'b0001;

	lut_sub lut_18671 ({g1492, g1493}, g1491);
	defparam lut_18671.LUT_SIZE = 2;
	defparam lut_18671.mask = 4'b1000;

	lut_sub lut_18677 ({g123, g1497}, g1492);
	defparam lut_18677.LUT_SIZE = 2;
	defparam lut_18677.mask = 4'b0100;

	lut_sub lut_18683 ({g123, g1498}, g1493);
	defparam lut_18683.LUT_SIZE = 2;
	defparam lut_18683.mask = 4'b0001;

	lut_sub lut_18689 ({g1495, g1496}, g1494);
	defparam lut_18689.LUT_SIZE = 2;
	defparam lut_18689.mask = 4'b1000;

	lut_sub lut_18695 ({g123, g1499}, g1495);
	defparam lut_18695.LUT_SIZE = 2;
	defparam lut_18695.mask = 4'b0100;

	lut_sub lut_18701 ({g123, g1500}, g1496);
	defparam lut_18701.LUT_SIZE = 2;
	defparam lut_18701.mask = 4'b0001;

	lut_sub lut_18709 ({g872, g868, g847, g848}, g1497);
	defparam lut_18709.LUT_SIZE = 4;
	defparam lut_18709.mask = 16'h0001;

	lut_sub lut_18716 ({g872, g868, g848}, g1498);
	defparam lut_18716.LUT_SIZE = 3;
	defparam lut_18716.mask = 8'h01;

	lut_sub lut_18724 ({g872, g868, g847, g848}, g1499);
	defparam lut_18724.LUT_SIZE = 4;
	defparam lut_18724.mask = 16'h0001;

	lut_sub lut_18732 ({g872, g868, g159, g848}, g1500);
	defparam lut_18732.LUT_SIZE = 4;
	defparam lut_18732.mask = 16'h0007;

	lut_sub lut_18740 ({g1502, g1503}, g1501);
	defparam lut_18740.LUT_SIZE = 2;
	defparam lut_18740.mask = 4'b1000;

	lut_sub lut_18746 ({g253, g1504}, g1502);
	defparam lut_18746.LUT_SIZE = 2;
	defparam lut_18746.mask = 4'b0100;

	lut_sub lut_18752 ({g253, g1505}, g1503);
	defparam lut_18752.LUT_SIZE = 2;
	defparam lut_18752.mask = 4'b0001;

	lut_sub lut_18758 ({g851, g1508}, g1504);
	defparam lut_18758.LUT_SIZE = 2;
	defparam lut_18758.mask = 4'b0001;

	lut_sub lut_18764 ({g1506, g1507}, g1505);
	defparam lut_18764.LUT_SIZE = 2;
	defparam lut_18764.mask = 4'b1000;

	lut_sub lut_18770 ({g851, g1509}, g1506);
	defparam lut_18770.LUT_SIZE = 2;
	defparam lut_18770.mask = 4'b0100;

	lut_sub lut_18776 ({g851, g1510}, g1507);
	defparam lut_18776.LUT_SIZE = 2;
	defparam lut_18776.mask = 4'b0001;

	lut_sub lut_18782 ({g862, g684}, g1508);
	defparam lut_18782.LUT_SIZE = 2;
	defparam lut_18782.mask = 4'b0001;

	lut_sub lut_18790 ({g75, g862, g408, g356}, g1509);
	defparam lut_18790.LUT_SIZE = 4;
	defparam lut_18790.mask = 16'h0002;

	lut_sub lut_18797 ({g862, g684, g356}, g1510);
	defparam lut_18797.LUT_SIZE = 3;
	defparam lut_18797.mask = 8'h0b;

	lut_sub lut_18805 ({g76, g1512}, g1511);
	defparam lut_18805.LUT_SIZE = 2;
	defparam lut_18805.mask = 4'b1000;

	lut_sub lut_18811 ({g76, g1513}, g1512);
	defparam lut_18811.LUT_SIZE = 2;
	defparam lut_18811.mask = 4'b0100;

	lut_sub lut_18817 ({g1514, g1515}, g1513);
	defparam lut_18817.LUT_SIZE = 2;
	defparam lut_18817.mask = 4'b1000;

	lut_sub lut_18822 ({i_11_, g1516}, g1514);
	defparam lut_18822.LUT_SIZE = 2;
	defparam lut_18822.mask = 4'b0100;

	lut_sub lut_18827 ({i_11_, g1517}, g1515);
	defparam lut_18827.LUT_SIZE = 2;
	defparam lut_18827.mask = 4'b0001;

	lut_sub lut_18832 ({i_15_, i_10_, g436, i_9_}, g1516);
	defparam lut_18832.LUT_SIZE = 4;
	defparam lut_18832.mask = 16'hdfff;

	lut_sub lut_18851 ({i_15_, i_10_, g422, i_9_}, g1517);
	defparam lut_18851.LUT_SIZE = 4;
	defparam lut_18851.mask = 16'hfeff;

	lut_sub lut_18871 ({g1519, g1520}, g1518);
	defparam lut_18871.LUT_SIZE = 2;
	defparam lut_18871.mask = 4'b1000;

	lut_sub lut_18877 ({g125, g1521}, g1519);
	defparam lut_18877.LUT_SIZE = 2;
	defparam lut_18877.mask = 4'b0100;

	lut_sub lut_18883 ({g125, g1524}, g1520);
	defparam lut_18883.LUT_SIZE = 2;
	defparam lut_18883.mask = 4'b0001;

	lut_sub lut_18889 ({g1522, g1523}, g1521);
	defparam lut_18889.LUT_SIZE = 2;
	defparam lut_18889.mask = 4'b1000;

	lut_sub lut_18895 ({g154, g1527}, g1522);
	defparam lut_18895.LUT_SIZE = 2;
	defparam lut_18895.mask = 4'b0100;

	lut_sub lut_18901 ({g154, g1528}, g1523);
	defparam lut_18901.LUT_SIZE = 2;
	defparam lut_18901.mask = 4'b0001;

	lut_sub lut_18907 ({g1525, g1526}, g1524);
	defparam lut_18907.LUT_SIZE = 2;
	defparam lut_18907.mask = 4'b1000;

	lut_sub lut_18913 ({g154, g1529}, g1525);
	defparam lut_18913.LUT_SIZE = 2;
	defparam lut_18913.mask = 4'b0100;

	lut_sub lut_18919 ({g154, g1530}, g1526);
	defparam lut_18919.LUT_SIZE = 2;
	defparam lut_18919.mask = 4'b0001;

	lut_sub lut_18927 ({g731, g641, g339, g640}, g1527);
	defparam lut_18927.LUT_SIZE = 4;
	defparam lut_18927.mask = 16'h0080;

	lut_sub lut_18935 ({g731, g641, g122, g640}, g1528);
	defparam lut_18935.LUT_SIZE = 4;
	defparam lut_18935.mask = 16'h00ec;

	lut_sub lut_18947 ({g731, g641, g339, g640}, g1529);
	defparam lut_18947.LUT_SIZE = 4;
	defparam lut_18947.mask = 16'h0080;

	lut_sub lut_18955 ({g731, g641, g122, g640}, g1530);
	defparam lut_18955.LUT_SIZE = 4;
	defparam lut_18955.mask = 16'h00a8;

	lut_sub lut_18963 ({g1532, g1533}, g1531);
	defparam lut_18963.LUT_SIZE = 2;
	defparam lut_18963.mask = 4'b1000;

	lut_sub lut_18969 ({g634, g1534}, g1532);
	defparam lut_18969.LUT_SIZE = 2;
	defparam lut_18969.mask = 4'b0100;

	lut_sub lut_18975 ({g634, g1537}, g1533);
	defparam lut_18975.LUT_SIZE = 2;
	defparam lut_18975.mask = 4'b0001;

	lut_sub lut_18981 ({g1535, g1536}, g1534);
	defparam lut_18981.LUT_SIZE = 2;
	defparam lut_18981.mask = 4'b1000;

	lut_sub lut_18986 ({i_8_, g73}, g1535);
	defparam lut_18986.LUT_SIZE = 2;
	defparam lut_18986.mask = 4'b1000;

	lut_sub lut_18991 ({i_8_, g1540}, g1536);
	defparam lut_18991.LUT_SIZE = 2;
	defparam lut_18991.mask = 4'b0001;

	lut_sub lut_18997 ({g1538, g1539}, g1537);
	defparam lut_18997.LUT_SIZE = 2;
	defparam lut_18997.mask = 4'b1000;

	lut_sub lut_19002 ({i_8_, g1541}, g1538);
	defparam lut_19002.LUT_SIZE = 2;
	defparam lut_19002.mask = 4'b0100;

	lut_sub lut_19007 ({i_8_, g1542}, g1539);
	defparam lut_19007.LUT_SIZE = 2;
	defparam lut_19007.mask = 4'b0001;

	lut_sub lut_19014 ({g700, g699, g73}, g1540);
	defparam lut_19014.LUT_SIZE = 3;
	defparam lut_19014.mask = 8'hab;

	lut_sub lut_19026 ({g701, g700, g37, g73}, g1541);
	defparam lut_19026.LUT_SIZE = 4;
	defparam lut_19026.mask = 16'haaab;

	lut_sub lut_19041 ({g700, g699, g73}, g1542);
	defparam lut_19041.LUT_SIZE = 3;
	defparam lut_19041.mask = 8'hab;

	lut_sub lut_19051 ({g1544, g1545}, g1543);
	defparam lut_19051.LUT_SIZE = 2;
	defparam lut_19051.mask = 4'b1000;

	lut_sub lut_19057 ({g102, g1546}, g1544);
	defparam lut_19057.LUT_SIZE = 2;
	defparam lut_19057.mask = 4'b0100;

	lut_sub lut_19063 ({g102, g1549}, g1545);
	defparam lut_19063.LUT_SIZE = 2;
	defparam lut_19063.mask = 4'b0001;

	lut_sub lut_19069 ({g1547, g1548}, g1546);
	defparam lut_19069.LUT_SIZE = 2;
	defparam lut_19069.mask = 4'b1000;

	lut_sub lut_19075 ({g22, g556}, g1547);
	defparam lut_19075.LUT_SIZE = 2;
	defparam lut_19075.mask = 4'b0100;

	lut_sub lut_19081 ({g22, g556}, g1548);
	defparam lut_19081.LUT_SIZE = 2;
	defparam lut_19081.mask = 4'b0001;

	lut_sub lut_19087 ({g1550, g1551}, g1549);
	defparam lut_19087.LUT_SIZE = 2;
	defparam lut_19087.mask = 4'b1000;

	lut_sub lut_19093 ({g22, g1552}, g1550);
	defparam lut_19093.LUT_SIZE = 2;
	defparam lut_19093.mask = 4'b0100;

	lut_sub lut_19099 ({g22, g1553}, g1551);
	defparam lut_19099.LUT_SIZE = 2;
	defparam lut_19099.mask = 4'b0001;

	lut_sub lut_19106 ({g460, g76, g556}, g1552);
	defparam lut_19106.LUT_SIZE = 3;
	defparam lut_19106.mask = 8'h01;

	lut_sub lut_19114 ({g460, g91, g113, g556}, g1553);
	defparam lut_19114.LUT_SIZE = 4;
	defparam lut_19114.mask = 16'h0155;

	lut_sub lut_19124 ({g1555, g1556}, g1554);
	defparam lut_19124.LUT_SIZE = 2;
	defparam lut_19124.mask = 4'b1000;

	lut_sub lut_19130 ({g513, g1557}, g1555);
	defparam lut_19130.LUT_SIZE = 2;
	defparam lut_19130.mask = 4'b0100;

	lut_sub lut_19136 ({g513, g1558}, g1556);
	defparam lut_19136.LUT_SIZE = 2;
	defparam lut_19136.mask = 4'b0001;

	lut_sub lut_19142 ({g122, g1561}, g1557);
	defparam lut_19142.LUT_SIZE = 2;
	defparam lut_19142.mask = 4'b0100;

	lut_sub lut_19148 ({g1559, g1560}, g1558);
	defparam lut_19148.LUT_SIZE = 2;
	defparam lut_19148.mask = 4'b1000;

	lut_sub lut_19154 ({g122, g1562}, g1559);
	defparam lut_19154.LUT_SIZE = 2;
	defparam lut_19154.mask = 4'b0100;

	lut_sub lut_19160 ({g122, g1563}, g1560);
	defparam lut_19160.LUT_SIZE = 2;
	defparam lut_19160.mask = 4'b0001;

	lut_sub lut_19167 ({g554, g135, g553}, g1561);
	defparam lut_19167.LUT_SIZE = 3;
	defparam lut_19167.mask = 8'h01;

	lut_sub lut_19173 ({g554, g553}, g1562);
	defparam lut_19173.LUT_SIZE = 2;
	defparam lut_19173.mask = 4'b0001;

	lut_sub lut_19181 ({g552, g554, g551, g553}, g1563);
	defparam lut_19181.LUT_SIZE = 4;
	defparam lut_19181.mask = 16'h0001;

	lut_sub lut_19187 ({g1565, g1566}, g1564);
	defparam lut_19187.LUT_SIZE = 2;
	defparam lut_19187.mask = 4'b1000;

	lut_sub lut_19193 ({g392, g1567}, g1565);
	defparam lut_19193.LUT_SIZE = 2;
	defparam lut_19193.mask = 4'b0100;

	lut_sub lut_19199 ({g392, g1570}, g1566);
	defparam lut_19199.LUT_SIZE = 2;
	defparam lut_19199.mask = 4'b0001;

	lut_sub lut_19205 ({g1568, g1569}, g1567);
	defparam lut_19205.LUT_SIZE = 2;
	defparam lut_19205.mask = 4'b1000;

	lut_sub lut_19210 ({i_15_, g1573}, g1568);
	defparam lut_19210.LUT_SIZE = 2;
	defparam lut_19210.mask = 4'b0100;

	lut_sub lut_19215 ({i_15_, g1574}, g1569);
	defparam lut_19215.LUT_SIZE = 2;
	defparam lut_19215.mask = 4'b0001;

	lut_sub lut_19221 ({g1571, g1572}, g1570);
	defparam lut_19221.LUT_SIZE = 2;
	defparam lut_19221.mask = 4'b1000;

	lut_sub lut_19226 ({i_15_, g1575}, g1571);
	defparam lut_19226.LUT_SIZE = 2;
	defparam lut_19226.mask = 4'b0100;

	lut_sub lut_19231 ({i_15_, g1576}, g1572);
	defparam lut_19231.LUT_SIZE = 2;
	defparam lut_19231.mask = 4'b0001;

	lut_sub lut_19239 ({g174, g428, g142, g524}, g1573);
	defparam lut_19239.LUT_SIZE = 4;
	defparam lut_19239.mask = 16'h1555;

	lut_sub lut_19252 ({g174, g520, g524}, g1574);
	defparam lut_19252.LUT_SIZE = 3;
	defparam lut_19252.mask = 8'h15;

	lut_sub lut_19261 ({g174, g428, g524}, g1575);
	defparam lut_19261.LUT_SIZE = 3;
	defparam lut_19261.mask = 8'h15;

	lut_sub lut_19270 ({g174, g520, g524}, g1576);
	defparam lut_19270.LUT_SIZE = 3;
	defparam lut_19270.mask = 8'h15;

	lut_sub lut_19278 ({g174, g1578}, g1577);
	defparam lut_19278.LUT_SIZE = 2;
	defparam lut_19278.mask = 4'b1000;

	lut_sub lut_19284 ({g174, g1579}, g1578);
	defparam lut_19284.LUT_SIZE = 2;
	defparam lut_19284.mask = 4'b0100;

	lut_sub lut_19290 ({g1580, g1581}, g1579);
	defparam lut_19290.LUT_SIZE = 2;
	defparam lut_19290.mask = 4'b1000;

	lut_sub lut_19295 ({i_9_, g1582}, g1580);
	defparam lut_19295.LUT_SIZE = 2;
	defparam lut_19295.mask = 4'b0100;

	lut_sub lut_19300 ({i_9_, g1583}, g1581);
	defparam lut_19300.LUT_SIZE = 2;
	defparam lut_19300.mask = 4'b0001;

	lut_sub lut_19305 ({i_15_, i_11_, g262, i_10_}, g1582);
	defparam lut_19305.LUT_SIZE = 4;
	defparam lut_19305.mask = 16'hfdff;

	lut_sub lut_19324 ({i_15_, i_11_, g518, i_10_}, g1583);
	defparam lut_19324.LUT_SIZE = 4;
	defparam lut_19324.mask = 16'hfdff;

	lut_sub lut_19344 ({g1585, g1586}, g1584);
	defparam lut_19344.LUT_SIZE = 2;
	defparam lut_19344.mask = 4'b1000;

	lut_sub lut_19349 ({i_15_, g1587}, g1585);
	defparam lut_19349.LUT_SIZE = 2;
	defparam lut_19349.mask = 4'b0100;

	lut_sub lut_19354 ({i_15_, g1589}, g1586);
	defparam lut_19354.LUT_SIZE = 2;
	defparam lut_19354.mask = 4'b0001;

	lut_sub lut_19359 ({i_11_, g1588}, g1587);
	defparam lut_19359.LUT_SIZE = 2;
	defparam lut_19359.mask = 4'b0010;

	lut_sub lut_19364 ({i_11_, g1591}, g1588);
	defparam lut_19364.LUT_SIZE = 2;
	defparam lut_19364.mask = 4'b0001;

	lut_sub lut_19369 ({i_11_, g1590}, g1589);
	defparam lut_19369.LUT_SIZE = 2;
	defparam lut_19369.mask = 4'b1000;

	lut_sub lut_19374 ({i_11_, g1592}, g1590);
	defparam lut_19374.LUT_SIZE = 2;
	defparam lut_19374.mask = 4'b0100;

	lut_sub lut_19380 ({g176, i_10_, g443, i_9_}, g1591);
	defparam lut_19380.LUT_SIZE = 4;
	defparam lut_19380.mask = 16'hf7ff;

	lut_sub lut_19400 ({g176, i_10_, g444, i_9_}, g1592);
	defparam lut_19400.LUT_SIZE = 4;
	defparam lut_19400.mask = 16'hf7ff;

	lut_sub lut_19420 ({g1594, g1595}, g1593);
	defparam lut_19420.LUT_SIZE = 2;
	defparam lut_19420.mask = 4'b1000;

	lut_sub lut_19426 ({g78, g1596}, g1594);
	defparam lut_19426.LUT_SIZE = 2;
	defparam lut_19426.mask = 4'b0100;

	lut_sub lut_19432 ({g78, g1599}, g1595);
	defparam lut_19432.LUT_SIZE = 2;
	defparam lut_19432.mask = 4'b0001;

	lut_sub lut_19438 ({g1597, g1598}, g1596);
	defparam lut_19438.LUT_SIZE = 2;
	defparam lut_19438.mask = 4'b1000;

	lut_sub lut_19444 ({g97, g1602}, g1597);
	defparam lut_19444.LUT_SIZE = 2;
	defparam lut_19444.mask = 4'b0100;

	lut_sub lut_19450 ({g97, g1603}, g1598);
	defparam lut_19450.LUT_SIZE = 2;
	defparam lut_19450.mask = 4'b0001;

	lut_sub lut_19456 ({g1600, g1601}, g1599);
	defparam lut_19456.LUT_SIZE = 2;
	defparam lut_19456.mask = 4'b1000;

	lut_sub lut_19462 ({g97, g1604}, g1600);
	defparam lut_19462.LUT_SIZE = 2;
	defparam lut_19462.mask = 4'b0100;

	lut_sub lut_19468 ({g97, g1605}, g1601);
	defparam lut_19468.LUT_SIZE = 2;
	defparam lut_19468.mask = 4'b0001;

	lut_sub lut_19476 ({g144, g425, g226, g142}, g1602);
	defparam lut_19476.LUT_SIZE = 4;
	defparam lut_19476.mask = 16'h0100;

	lut_sub lut_19484 ({g144, g425, g114, g142}, g1603);
	defparam lut_19484.LUT_SIZE = 4;
	defparam lut_19484.mask = 16'h0501;

	lut_sub lut_19493 ({g144, g425, g226}, g1604);
	defparam lut_19493.LUT_SIZE = 3;
	defparam lut_19493.mask = 8'h10;

	lut_sub lut_19500 ({g144, g425, g114}, g1605);
	defparam lut_19500.LUT_SIZE = 3;
	defparam lut_19500.mask = 8'h75;

	lut_sub lut_19510 ({g24, g1607}, g1606);
	defparam lut_19510.LUT_SIZE = 2;
	defparam lut_19510.mask = 4'b1000;

	lut_sub lut_19516 ({g24, g1608}, g1607);
	defparam lut_19516.LUT_SIZE = 2;
	defparam lut_19516.mask = 4'b0100;

	lut_sub lut_19522 ({g1609, g1610}, g1608);
	defparam lut_19522.LUT_SIZE = 2;
	defparam lut_19522.mask = 4'b1000;

	lut_sub lut_19527 ({i_11_, g1611}, g1609);
	defparam lut_19527.LUT_SIZE = 2;
	defparam lut_19527.mask = 4'b0100;

	lut_sub lut_19532 ({i_11_, g1612}, g1610);
	defparam lut_19532.LUT_SIZE = 2;
	defparam lut_19532.mask = 4'b0001;

	lut_sub lut_19537 ({i_15_, i_10_, g144, i_9_}, g1611);
	defparam lut_19537.LUT_SIZE = 4;
	defparam lut_19537.mask = 16'hefff;

	lut_sub lut_19556 ({i_15_, i_10_, g165, i_9_}, g1612);
	defparam lut_19556.LUT_SIZE = 4;
	defparam lut_19556.mask = 16'hefff;

	lut_sub lut_19576 ({g1614, g1615}, g1613);
	defparam lut_19576.LUT_SIZE = 2;
	defparam lut_19576.mask = 4'b1000;

	lut_sub lut_19582 ({g102, g1616}, g1614);
	defparam lut_19582.LUT_SIZE = 2;
	defparam lut_19582.mask = 4'b0100;

	lut_sub lut_19588 ({g102, g1619}, g1615);
	defparam lut_19588.LUT_SIZE = 2;
	defparam lut_19588.mask = 4'b0001;

	lut_sub lut_19594 ({g1617, g1618}, g1616);
	defparam lut_19594.LUT_SIZE = 2;
	defparam lut_19594.mask = 4'b1000;

	lut_sub lut_19600 ({g155, g1622}, g1617);
	defparam lut_19600.LUT_SIZE = 2;
	defparam lut_19600.mask = 4'b0100;

	lut_sub lut_19606 ({g155, g1623}, g1618);
	defparam lut_19606.LUT_SIZE = 2;
	defparam lut_19606.mask = 4'b0001;

	lut_sub lut_19612 ({g1620, g1621}, g1619);
	defparam lut_19612.LUT_SIZE = 2;
	defparam lut_19612.mask = 4'b1000;

	lut_sub lut_19618 ({g155, g323}, g1620);
	defparam lut_19618.LUT_SIZE = 2;
	defparam lut_19618.mask = 4'b0100;

	lut_sub lut_19624 ({g155, g1624}, g1621);
	defparam lut_19624.LUT_SIZE = 2;
	defparam lut_19624.mask = 4'b0001;

	lut_sub lut_19632 ({g24, g323, g107, g254}, g1622);
	defparam lut_19632.LUT_SIZE = 4;
	defparam lut_19632.mask = 16'h1f5f;

	lut_sub lut_19650 ({g24, g323, g126, g254}, g1623);
	defparam lut_19650.LUT_SIZE = 4;
	defparam lut_19650.mask = 16'h7fff;

	lut_sub lut_19671 ({g24, g323, g126}, g1624);
	defparam lut_19671.LUT_SIZE = 3;
	defparam lut_19671.mask = 8'h7f;

	lut_sub lut_19683 ({g68, g1626}, g1625);
	defparam lut_19683.LUT_SIZE = 2;
	defparam lut_19683.mask = 4'b1000;

	lut_sub lut_19689 ({g68, g1627}, g1626);
	defparam lut_19689.LUT_SIZE = 2;
	defparam lut_19689.mask = 4'b0100;

	lut_sub lut_19695 ({g1628, g1629}, g1627);
	defparam lut_19695.LUT_SIZE = 2;
	defparam lut_19695.mask = 4'b1000;

	lut_sub lut_19700 ({i_11_, g1630}, g1628);
	defparam lut_19700.LUT_SIZE = 2;
	defparam lut_19700.mask = 4'b0100;

	lut_sub lut_19705 ({i_11_, g1631}, g1629);
	defparam lut_19705.LUT_SIZE = 2;
	defparam lut_19705.mask = 4'b0001;

	lut_sub lut_19710 ({i_15_, i_10_, g157, i_9_}, g1630);
	defparam lut_19710.LUT_SIZE = 4;
	defparam lut_19710.mask = 16'hfeff;

	lut_sub lut_19729 ({i_15_, i_10_, g254, i_9_}, g1631);
	defparam lut_19729.LUT_SIZE = 4;
	defparam lut_19729.mask = 16'hf7ff;

	lut_sub lut_19749 ({g68, g1633}, g1632);
	defparam lut_19749.LUT_SIZE = 2;
	defparam lut_19749.mask = 4'b1000;

	lut_sub lut_19755 ({g68, g1634}, g1633);
	defparam lut_19755.LUT_SIZE = 2;
	defparam lut_19755.mask = 4'b0100;

	lut_sub lut_19761 ({g1635, g1636}, g1634);
	defparam lut_19761.LUT_SIZE = 2;
	defparam lut_19761.mask = 4'b1000;

	lut_sub lut_19766 ({i_11_, g1637}, g1635);
	defparam lut_19766.LUT_SIZE = 2;
	defparam lut_19766.mask = 4'b0100;

	lut_sub lut_19771 ({i_11_, g1638}, g1636);
	defparam lut_19771.LUT_SIZE = 2;
	defparam lut_19771.mask = 4'b0001;

	lut_sub lut_19776 ({i_15_, i_10_, g131, i_9_}, g1637);
	defparam lut_19776.LUT_SIZE = 4;
	defparam lut_19776.mask = 16'hbfff;

	lut_sub lut_19795 ({i_15_, i_10_, g122, i_9_}, g1638);
	defparam lut_19795.LUT_SIZE = 4;
	defparam lut_19795.mask = 16'hfeff;

	lut_sub lut_19815 ({g1640, g1641}, g1639);
	defparam lut_19815.LUT_SIZE = 2;
	defparam lut_19815.mask = 4'b1000;

	lut_sub lut_19821 ({g75, g1642}, g1640);
	defparam lut_19821.LUT_SIZE = 2;
	defparam lut_19821.mask = 4'b0100;

	lut_sub lut_19827 ({g75, g1643}, g1641);
	defparam lut_19827.LUT_SIZE = 2;
	defparam lut_19827.mask = 4'b0001;

	lut_sub lut_19833 ({g87, g1646}, g1642);
	defparam lut_19833.LUT_SIZE = 2;
	defparam lut_19833.mask = 4'b0001;

	lut_sub lut_19839 ({g1644, g1645}, g1643);
	defparam lut_19839.LUT_SIZE = 2;
	defparam lut_19839.mask = 4'b1000;

	lut_sub lut_19845 ({g87, g1647}, g1644);
	defparam lut_19845.LUT_SIZE = 2;
	defparam lut_19845.mask = 4'b0100;

	lut_sub lut_19851 ({g87, g1648}, g1645);
	defparam lut_19851.LUT_SIZE = 2;
	defparam lut_19851.mask = 4'b0001;

	lut_sub lut_19858 ({g79, g89, g125}, g1646);
	defparam lut_19858.LUT_SIZE = 3;
	defparam lut_19858.mask = 8'h23;

	lut_sub lut_19868 ({g131, g79, g130, g125}, g1647);
	defparam lut_19868.LUT_SIZE = 4;
	defparam lut_19868.mask = 16'h0023;

	lut_sub lut_19876 ({g79, g125}, g1648);
	defparam lut_19876.LUT_SIZE = 2;
	defparam lut_19876.mask = 4'b1011;


endmodule