module diffeq (
	PCLK, PRESET, Pdxport_0_0_, Pdxport_1_1_, Pdxport_2_2_, Pdxport_3_3_, Pdxport_4_4_, Pdxport_5_5_, 
	Pdxport_6_6_, Pdxport_7_7_, Pdxport_8_8_, Pdxport_9_9_, Pdxport_10_10_, Pdxport_11_11_, Paport_0_0_, Paport_1_1_, Paport_2_2_, Paport_3_3_, 
	Paport_4_4_, Paport_5_5_, Paport_6_6_, Paport_7_7_, Paport_8_8_, Paport_9_9_, Paport_10_10_, Paport_11_11_, Preset_0_0_, Pready_0_0_, 
	PDN, Pnext_0_0_, Pover_0_0_);

input PCLK, PRESET, Pdxport_0_0_, Pdxport_1_1_, Pdxport_2_2_, Pdxport_3_3_, Pdxport_4_4_, Pdxport_5_5_, Pdxport_6_6_, Pdxport_7_7_, Pdxport_8_8_, Pdxport_9_9_, Pdxport_10_10_, Pdxport_11_11_, Paport_0_0_, Paport_1_1_, Paport_2_2_, Paport_3_3_, Paport_4_4_, Paport_5_5_, Paport_6_6_, Paport_7_7_, Paport_8_8_, Paport_9_9_, Paport_10_10_, Paport_11_11_, Preset_0_0_, Pready_0_0_;

output PDN, Pnext_0_0_, Pover_0_0_;

wire n3, n2, N_N4254, n4, N_N4238, n5, N_N4231, n6, N_N4229, n7, N_N4217, n8, N_N4174, n9, N_N4166, n11, N_N4139, n12, N_N4113, n13, N_N4110, n14, N_N4105, n15, N_N4098, n16, N_N4094, n17, N_N4089, n18, N_N4085, n19, N_N4074, n22, N_N4055, n23, N_N4053, n24, N_N4046, n25, N_N4044, n26, N_N4041, n27, N_N4038, n28, N_N4032, n29, N_N4029, n30, N_N4028, n31, N_N4023, n32, N_N4020, n34, N_N4007, n35, N_N3987, n36, N_N3980, n38, N_N3969, n39, N_N3967, n40, N_N3963, n41, N_N3958, n42, N_N3956, n43, N_N3946, n44, N_N3941, n46, N_N3915, n47, N_N3914, n48, N_N3913, n49, N_N3909, N_N3904, n51, N_N3895, n56, N_N3847, n57, N_N3828, n58, N_N3825, n59, N_N3823, n60, N_N3817, n61, N_N3814, n62, N_N3804, n63, N_N3801, n64, N_N3798, n65, N_N3795, n66, N_N3787, n67, N_N3785, n68, N_N3772, n72, N_N3752, n73, N_N3744, n74, N_N3740, N_N3739, n78, N_N3723, n80, N_N3720, n81, N_N3717, n82, N_N3712, n83, N_N3710, N_N3707, n84, N_N3705, n86, N_N3695, N_N3690, n89, N_N3683, n90, N_N3671, n91, N_N3668, n92, N_N3666, n93, N_N3664, n94, N_N3662, n95, N_N3661, n96, N_N3658, n97, N_N3653, n98, N_N3652, n102, N_N3640, N_N3638, n104, N_N3633, n108, n106, N_N3811, N_N3620, n111, N_N3618, n112, N_N3616, n113, N_N3615, n114, N_N3614, n115, N_N3611, n118, N_N3602, n119, N_N3599, n120, N_N3596, n121, N_N3595, n122, N_N3592, n123, N_N3589, n124, N_N3586, n125, N_N3584, n126, N_N3579, n127, N_N3570, n130, N_N3559, n131, N_N3558, N_N3530, n135, N_N3524, n136, N_N3523, n137, N_N3511, n138, N_N3506, n139, N_N3503, n140, N_N3499, n143, N_N3488, n144, N_N3487, n145, N_N3486, n146, N_N3483, n147, N_N3481, n148, N_N3479, n149, N_N3476, n150, N_N3474, n151, N_N3472, N_N3465, n152, N_N3458, n153, N_N3456, n154, N_N3454, n156, N_N3449, n158, N_N3437, n159, N_N3435, N_N3432, n160, N_N3431, N_N3425, n162, N_N3423, n163, N_N3416, n164, N_N3413, n165, N_N3409, n166, N_N3406, n167, N_N3401, n168, N_N3400, n169, N_N3399, N_N3390, N_N3389, N_N3374, n172, N_N3372, n173, N_N3366, n175, N_N3352, n176, N_N3349, N_N3348, n178, N_N3339, N_N3338, n179, N_N3335, n180, N_N3334, n181, N_N3332, n183, N_N3325, n184, N_N3322, n185, N_N3321, n186, N_N3320, n187, N_N3318, n188, N_N3316, n189, N_N3315, N_N3314, n190, N_N3310, N_N3305, N_N3287, n193, N_N3284, n194, N_N3277, n195, N_N3276, n196, N_N3273, n197, N_N3266, n198, N_N3263, n199, N_N3259, n200, N_N3249, n201, N_N3247, n203, N_N3244, n204, N_N3241, n205, N_N3240, n206, N_N3231, n207, N_N3227, n208, N_N3222, n209, N_N3216, n210, N_N3215, n211, N_N3213, n212, N_N3211, n213, N_N3210, n214, N_N3209, N_N3206, n215, N_N3204, n216, N_N3202, n217, N_N3201, n218, N_N3200, n220, N_N3194, n221, N_N3193, n222, N_N3192, n223, N_N3191, n224, N_N3190, n225, N_N3189, n228, N_N3178, n229, N_N3177, n230, N_N3174, n231, N_N3173, n232, N_N3172, n234, N_N3165, n235, N_N3163, n236, N_N3162, N_N3160, N_N3156, N_N3155, n239, N_N3153, n240, N_N3152, n242, N_N3147, n243, N_N3146, n244, N_N3145, n245, N_N3144, n247, N_N3136, n248, N_N3133, n249, N_N3132, n250, N_N3130, n251, N_N3129, n253, N_N3123, N_N3119, n255, N_N3117, n256, N_N3115, n257, N_N3113, n258, N_N3106, n259, N_N3104, n260, N_N3103, n261, N_N3102, n262, N_N3101, n263, N_N3093, n264, N_N3091, n265, N_N3087, n266, N_N3086, N_N3078, n267, N_N3075, n269, N_N3070, n270, N_N3068, N_N3063, n275, N_N3058, n276, N_N3057, n277, N_N3053, n278, N_N3052, n279, N_N3051, n280, N_N3050, n281, N_N3049, n282, N_N3048, N_N3041, n286, N_N3040, N_N3038, n287, N_N3037, n288, N_N3034, n291, N_N3028, n292, N_N3027, N_N3016, n296, N_N3015, n297, N_N3014, n299, N_N3010, n300, N_N3009, n301, N_N3008, n302, N_N3007, n303, N_N3004, n304, N_N3003, n307, N_N2998, n308, N_N2997, N_N2996, n310, N_N2992, n312, N_N2988, n313, N_N2987, n315, N_N2984, n316, N_N2983, n318, N_N2980, n319, N_N2979, n320, N_N2978, n321, N_N2977, n322, N_N2976, n323, N_N2975, n324, N_N2974, n325, N_N2973, n326, N_N2972, n328, N_N2969, N_N2966, N_N2965, n330, N_N2964, n331, N_N2963, n332, N_N2962, n333, N_N2961, N_N2958, N_N2957, n335, N_N2956, n336, N_N2955, n337, N_N2953, n338, N_N2952, n339, N_N46, n340, N_N45, n341, N_N44, n342, N_N43, n343, N_N42, n344, N_N41, n345, N_N40, n346, N_N39, n347, N_N38, n348, N_N37, n349, N_N36, n351, n352, n350, n355, n353, n357, n356, n361, n362, n360, n358, n365, n366, n363, n369, n370, n367, n374, n375, n372, n371, n378, n379, n376, n382, n383, n380, n387, n388, n385, n384, n392, n393, n390, n389, n396, n397, n394, n400, n401, n398, n404, n405, n402, n408, n409, n406, n411, n412, n410, n414, n413, n417, n416, N_N47, n421, n418, n424, n422, n428, n425, n432, n429, n436, n433, n440, n437, n444, n441, n448, n445, n452, n449, n461, n460, n458, n463, n464, n466, n475, n476, n473, n478, n481, n484, n487, n490, n493, n496, n499, n502, n505, n508, n511, n514, n518, n517, n519, n522, n525, n528, n534, n533, n536, n537, n540, n542, n543, n544, n546, n550, n549, n551, n553, n554, n557, n559, n560, n564, n563, n565, n567, n568, n571, n573, n575, n574, n576, n577, n580, n581, n583, n585, n584, n586, n591, n596, n594, n597, n599, n602, n600, n604, n607, n609, n610, n616, n613, n619, n618, n623, n621, n624, n625, n626, n635, n636, n637, n638, n639, n640, n641, n642, n645, n648, n650, n653, n656, n659, n662, n665, n668, n671, n676, n678, n679, n680, n681, n682, n684, n687, n688, n689, n691, n694, n695, n696, n698, n701, n702, n703, n706, n709, n710, n711, n712, n713, n716, n719, n720, n722, n724, n725, n726, n727, n729, n730, n731, n735, n736, n739, n741, n742, n744, n746, n748, n750, n752, n754, n756, n759, n760, n761, n764, n765, n767, n769, n771, n773, n775, n776, n778, n781, n783, n784, n793, n802, n803, n800, n806, n807, n804, n810, n811, n808, n814, n815, n812, n818, n819, n816, n822, n823, n820, n826, n827, n824, n830, n831, n828, n834, n835, n832, n838, n839, n836, n842, n843, n840, n846, n847, n844, n849, n848, n850, n852, n854, n855, n857, n858, n860, n861, n863, n864, n866, n867, n869, n870, n872, n873, n875, n876, n878, n882, n880, n881, n879, n885, n886, n887, n888, n889, n892, n897, n895, n899, n900, n909, n914, n916, n918, n926, n929, n927, n931, n930, n932, n934, n935, n939, n944, n946, n947, n950, n951, n955, n954, n956, n958, n957, n961, n960, n963, n962, n965, n964, n966, n971, n969, n980, n979, n983, n981, n987, n985, n991, n994, n997, n999, n1001, n1003, n1005, n1006, n1007, n1014, n1012, n1016, n1015, n1018, n1017, n1031, n1030, n1034, n1033, n1032, n1041, n1042, n1047, n1048, n1049, n1050, n1052, n1051, n1058, n1059, n1061, n1063, n1062, n1064, n1066, n1067, n1072, n1073, n1082, n1081, n1086, n1091, n1090, n1100, n1102, n1105, n1104, n1108, n1115, n1116, n1118, n1117, n1129, n1128, n1127, n1138, n1141, n1162, n1172, n1173, n1178, n1179, n1180, N_N3542, n1181, N_N3061, n1182, N_N3042, N_N3005, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1192, n1191, n1195, n1196, n1194, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1216, n1217, n1221, n1226, n1227, n1228, n1230, n1233, n1235, n1237, n1238, n1242, n1245, n1247, n1250, n1252, n1254, n1271, n1273, n1275, n1276, N_N3859, n1277, n1283, N_N3538, N_N3029, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1299;

reg N_N4054, N_N3745, N_N4119, N_N3826, N_N3818, N_N3345, N_N3924, N_N3815, N_N3691, N_N3157, N_N3872, N_N3788, N_N3375, N_N3143, N_N4197, N_N3843, N_N3426, N_N4118, N_N3580, N_N3175, N_N3071, N_N3808, N_N3923, N_N3250, N_N4221, N_N3069, N_N3464, N_N3535, N_N3871, N_N3248, N_N4180, N_N3311, N_N3442, N_N3981, N_N3842, N_N3105, N_N4133, N_N4117, N_N3420, N_N3761, N_N3062, N_N4071, N_N4227, N_N3807, N_N4145, N_N3922, N_N3516, N_N3489, N_N4030, N_N3540, N_N3513, N_N4083, N_N3841, N_N4018, N_N3971, N_N4232, N_N4246, N_N3806, N_N3992, N_N4086, N_N4230, N_N4212, Pnext_0_0_, N_N3626, N_N3965, N_N3890, NDN3_11, NDN5_10, N_N3786, N_N4171, NDN5_16, N_N3799, N_N3844, N_N3196, N_N4126, N_N3681, N_N3679, N_N3340, N_N4116, N_N3810, N_N3235, N_N3283, N_N3716, N_N3701, N_N3921, N_N3625, N_N3751, N_N3736, N_N3870, N_N4024, N_N3876, N_N3840, N_N4021, N_N3932, NLC1_2, N_N3805, N_N3700, N_N3735, NLak3_2, NLak3_9, N_N3906, N_N3388, N_N4057, N_N3011, N_N3346, N_N3677, N_N4165, N_N4080, N_N3373, N_N3709, N_N4206, N_N3324, N_N3575, N_N4159, NAK5_2, N_N3916, N_N3743, N_N4242, N_N3312, N_N3733, N_N3774, N_N4214, N_N3294, N_N3796, N_N3574, N_N3791, N_N3480, N_N4243, N_N3940, N_N3509, N_N4015, N_N2989, N_N3919, N_N3578, N_N3529, N_N4222, N_N3910, N_N3868, N_N3947, N_N4181, N_N3793, N_N3822, N_N3813, N_N4114, N_N4134, N_N3866, N_N4218, N_N3939, N_N3776, N_N3387, N_N4194, N_N3821, N_N3882, N_N4167, N_N3800, N_N4237, N_N3417, N_N3918, N_N4158, N_N3630, N_N3344, N_N4072, N_N3274, N_N3473, N_N4205, N_N4111, N_N3680, N_N3838, N_N3262, N_N4099, N_N3607, N_N3323, N_N3612, N_N4079, PDN, N_N3457, N_N3445, N_N3794, N_N3663, N_N3715, N_N4039, N_N3280, N_N4239, N_N3988, N_N3433, N_N4075, N_N3468, N_N4045, N_N3482, N_N3832, N_N3304, N_N3750, N_N3634, N_N3293, N_N3659, N_N4252, N_N3912, N_N3862, N_N3221, N_N3875, N_N3949, N_N3908, N_N3711, N_N3931, N_N3469, N_N3436, N_N3974, N_N3905, N_N3741, N_N3369, N_N3164, N_N3500, N_N3996, N_N3356, N_N4093, Pover_0_0_, N_N4224, N_N4027, NDN1_4, N_N3384, N_N4036, N_N3968, N_N4183, NGFDN_3, N_N4090, N_N4004, N_N3205, N_N4136, N_N3303, N_N3533, N_N3336, N_N3961, N_N3331, N_N3203, N_N4236, N_N3884, N_N3367, N_N4140, NDN2_2, N_N4106, N_N3100, N_N4193, N_N3470, N_N3424, N_N3959, N_N3393, N_N4042, N_N3188, N_N4095, N_N3957, N_N3517, N_N4047, N_N3081, N_N3541, N_N4177, NDN3_3, N_N4176, N_N3585, NDN3_8, N_N4209, N_N3824, N_N4208, N_N4120, N_N3708, N_N4220, N_N3999, N_N4223, N_N3179, N_N4179, N_N3475, N_N4132, N_N4182, N_N3797, N_N3214, N_N4070, N_N4135, NLD3_9, NDN5_2, NDN5_3, N_N3778, NDN5_4, N_N3212, NDN5_5, NDN5_6, NDN5_7, NDN5_8, N_N4073, NDN5_9, NEN5_9, N_N3684, N_N4056, N_N3713, N_N3829, N_N4060, NSr3_2, NSr5_2, NSr5_3, N_N3462, N_N3460, NSr5_4, NSr3_9, NSr5_5, NSr5_7, NSr5_8, N_N3998;

always  @(posedge PCLK)
	N_N4054<=N_N4053;

 always  @(posedge PCLK)
	N_N3745<=N_N3744;

 always  @(posedge PCLK)
	N_N4119<=N_N3406;

 always  @(posedge PCLK)
	N_N3826<=N_N3825;

 always  @(posedge PCLK)
	N_N3818<=N_N3817;

 always  @(posedge PCLK)
	N_N3345<=N_N3078;

 always  @(posedge PCLK)
	N_N3924<=N_N3409;

 always  @(posedge PCLK)
	N_N3815<=N_N3814;

 always  @(posedge PCLK)
	N_N3691<=N_N3690;

 always  @(posedge PCLK)
	N_N3157<=N_N2972;

 always  @(posedge PCLK)
	N_N3872<=N_N3123;

 always  @(posedge PCLK)
	N_N3788<=N_N3787;

 always  @(posedge PCLK)
	N_N3375<=N_N3374;

 always  @(posedge PCLK)
	N_N3143<=N_N3136;

 always  @(posedge PCLK)
	N_N4197<=N_N3847;

 always  @(posedge PCLK)
	N_N3843<=N_N3668;

 always  @(posedge PCLK)
	N_N3426<=N_N3425;

 always  @(posedge PCLK)
	N_N4118<=N_N3506;

 always  @(posedge PCLK)
	N_N3580<=N_N3579;

 always  @(posedge PCLK)
	N_N3175<=N_N3174;

 always  @(posedge PCLK)
	N_N3071<=N_N3070;

 always  @(posedge PCLK)
	N_N3808<=N_N3349;

 always  @(posedge PCLK)
	N_N3923<=N_N3227;

 always  @(posedge PCLK)
	N_N3250<=N_N3249;

 always  @(posedge PCLK)
	N_N4221<=N_N3486;

 always  @(posedge PCLK)
	N_N3069<=N_N3068;

 always  @(posedge PCLK)
	N_N3464<=N_N3216;

 always  @(posedge PCLK)
	N_N3535<=N_N3454;

 always  @(posedge PCLK)
	N_N3871<=N_N2952;

 always  @(posedge PCLK)
	N_N3248<=N_N3247;

 always  @(posedge PCLK)
	N_N4180<=N_N3334;

 always  @(posedge PCLK)
	N_N3311<=N_N3310;

 always  @(posedge PCLK)
	N_N3442<=N_N3215;

 always  @(posedge PCLK)
	N_N3981<=N_N3980;

 always  @(posedge PCLK)
	N_N3842<=N_N3413;

 always  @(posedge PCLK)
	N_N3105<=N_N3104;

 always  @(posedge PCLK)
	N_N4133<=N_N2997;

 always  @(posedge PCLK)
	N_N4117<=N_N3661;

 always  @(posedge PCLK)
	N_N3420<=N_N2973;

 always  @(posedge PCLK)
	N_N3761<=N_N3640;

 always  @(posedge PCLK)
	N_N3062<=N_N3009;

 always  @(posedge PCLK)
	N_N4071<=N_N3615;

 always  @(posedge PCLK)
	N_N4227<=N_N3859;

 always  @(posedge PCLK)
	N_N3807<=N_N3129;

 always  @(posedge PCLK)
	N_N4145<=N_N3222;

 always  @(posedge PCLK)
	N_N3922<=N_N3652;

 always  @(posedge PCLK)
	N_N3516<=N_N2992;

 always  @(posedge PCLK)
	N_N3489<=N_N3488;

 always  @(posedge PCLK)
	N_N4030<=N_N4029;

 always  @(posedge PCLK)
	N_N3540<=N_N3050;

 always  @(posedge PCLK)
	N_N3513<=N_N3487;

 always  @(posedge PCLK)
	N_N4083<=N_N2963;

 always  @(posedge PCLK)
	N_N3841<=N_N3431;

 always  @(posedge PCLK)
	N_N4018<=N_N3717;

 always  @(posedge PCLK)
	N_N3971<=N_N3801;

 always  @(posedge PCLK)
	N_N4232<=N_N4231;

 always  @(posedge PCLK)
	N_N4246<=N_N3276;

 always  @(posedge PCLK)
	N_N3806<=N_N3173;

 always  @(posedge PCLK)
	N_N3992<=N_N3723;

 always  @(posedge PCLK)
	N_N4086<=N_N4085;

 always  @(posedge PCLK)
	N_N4230<=N_N4229;

 always  @(posedge PCLK)
	N_N4212<=N_N3599;

 always  @(posedge PCLK)
	Pnext_0_0_<=N_N3005;

 always  @(posedge PCLK)
	N_N3626<=N_N3162;

 always  @(posedge PCLK)
	N_N3965<=N_N3106;

 always  @(posedge PCLK)
	N_N3890<=N_N3570;

 always  @(posedge PCLK)
	NDN3_11<=N_N3287;

 always  @(posedge PCLK)
	NDN5_10<=N_N3231;

 always  @(posedge PCLK)
	N_N3786<=N_N3785;

 always  @(posedge PCLK)
	N_N4171<=N_N3596;

 always  @(posedge PCLK)
	NDN5_16<=N_N3063;

 always  @(posedge PCLK)
	N_N3799<=N_N3798;

 always  @(posedge PCLK)
	N_N3844<=N_N3315;

 always  @(posedge PCLK)
	N_N3196<=N_N3152;

 always  @(posedge PCLK)
	N_N4126<=N_N3277;

 always  @(posedge PCLK)
	N_N3681<=N_N3400;

 always  @(posedge PCLK)
	N_N3679<=N_N3049;

 always  @(posedge PCLK)
	N_N3340<=N_N3339;

 always  @(posedge PCLK)
	N_N4116<=N_N3969;

 always  @(posedge PCLK)
	N_N3810<=N_N3316;

 always  @(posedge PCLK)
	N_N3235<=N_N2974;

 always  @(posedge PCLK)
	N_N3283<=N_N3053;

 always  @(posedge PCLK)
	N_N3716<=N_N3399;

 always  @(posedge PCLK)
	N_N3701<=N_N3048;

 always  @(posedge PCLK)
	N_N3921<=N_N3524;

 always  @(posedge PCLK)
	N_N3625<=N_N3558;

 always  @(posedge PCLK)
	N_N3751<=N_N3115;

 always  @(posedge PCLK)
	N_N3736<=N_N3456;

 always  @(posedge PCLK)
	N_N3870<=N_N3772;

 always  @(posedge PCLK)
	N_N4024<=N_N4023;

 always  @(posedge PCLK)
	N_N3876<=N_N3804;

 always  @(posedge PCLK)
	N_N3840<=N_N3133;

 always  @(posedge PCLK)
	N_N4021<=N_N4020;

 always  @(posedge PCLK)
	N_N3932<=N_N3189;

 always  @(posedge PCLK)
	NLC1_2<=N_N3811;

 always  @(posedge PCLK)
	N_N3805<=N_N3132;

 always  @(posedge PCLK)
	N_N3700<=N_N3259;

 always  @(posedge PCLK)
	N_N3735<=N_N3015;

 always  @(posedge PCLK)
	NLak3_2<=N_N2987;

 always  @(posedge PCLK)
	NLak3_9<=N_N3465;

 always  @(posedge PCLK)
	N_N3906<=N_N3003;

 always  @(posedge PCLK)
	N_N3388<=N_N2953;

 always  @(posedge PCLK)
	N_N4057<=N_N4007;

 always  @(posedge PCLK)
	N_N3011<=N_N2969;

 always  @(posedge PCLK)
	N_N3346<=N_N3037;

 always  @(posedge PCLK)
	N_N3677<=N_N2998;

 always  @(posedge PCLK)
	N_N4165<=N_N3146;

 always  @(posedge PCLK)
	N_N4080<=N_N3010;

 always  @(posedge PCLK)
	N_N3373<=N_N3372;

 always  @(posedge PCLK)
	N_N3709<=N_N3616;

 always  @(posedge PCLK)
	N_N4206<=N_N3483;

 always  @(posedge PCLK)
	N_N3324<=N_N3119;

 always  @(posedge PCLK)
	N_N3575<=N_N3325;

 always  @(posedge PCLK)
	N_N4159<=N_N3058;

 always  @(posedge PCLK)
	NAK5_2<=N_N3638;

 always  @(posedge PCLK)
	N_N3916<=N_N3915;

 always  @(posedge PCLK)
	N_N3743<=N_N3666;

 always  @(posedge PCLK)
	N_N4242<=N_N3052;

 always  @(posedge PCLK)
	N_N3312<=N_N2966;

 always  @(posedge PCLK)
	N_N3733<=N_N3595;

 always  @(posedge PCLK)
	N_N3774<=N_N3664;

 always  @(posedge PCLK)
	N_N4214<=N_N3332;

 always  @(posedge PCLK)
	N_N3294<=N_N2965;

 always  @(posedge PCLK)
	N_N3796<=N_N3795;

 always  @(posedge PCLK)
	N_N3574<=N_N3523;

 always  @(posedge PCLK)
	N_N3791<=N_N3653;

 always  @(posedge PCLK)
	N_N3480<=N_N3266;

 always  @(posedge PCLK)
	N_N4243<=N_N3914;

 always  @(posedge PCLK)
	N_N3940<=N_N3263;

 always  @(posedge PCLK)
	N_N3509<=N_N3241;

 always  @(posedge PCLK)
	N_N4015<=N_N3913;

 always  @(posedge PCLK)
	N_N2989<=N_N2988;

 always  @(posedge PCLK)
	N_N3919<=N_N2955;

 always  @(posedge PCLK)
	N_N3578<=N_N3389;

 always  @(posedge PCLK)
	N_N3529<=N_N3240;

 always  @(posedge PCLK)
	N_N4222<=N_N4174;

 always  @(posedge PCLK)
	N_N3910<=N_N3909;

 always  @(posedge PCLK)
	N_N3868<=N_N2956;

 always  @(posedge PCLK)
	N_N3947<=N_N3946;

 always  @(posedge PCLK)
	N_N4181<=N_N3390;

 always  @(posedge PCLK)
	N_N3793<=N_N3695;

 always  @(posedge PCLK)
	N_N3822<=N_N3004;

 always  @(posedge PCLK)
	N_N3813<=N_N3153;

 always  @(posedge PCLK)
	N_N4114<=N_N4113;

 always  @(posedge PCLK)
	N_N4134<=N_N3156;

 always  @(posedge PCLK)
	N_N3866<=N_N2961;

 always  @(posedge PCLK)
	N_N4218<=N_N4217;

 always  @(posedge PCLK)
	N_N3939<=N_N3589;

 always  @(posedge PCLK)
	N_N3776<=N_N3614;

 always  @(posedge PCLK)
	N_N3387<=N_N3145;

 always  @(posedge PCLK)
	N_N4194<=N_N3051;

 always  @(posedge PCLK)
	N_N3821<=N_N3014;

 always  @(posedge PCLK)
	N_N3882<=N_N3705;

 always  @(posedge PCLK)
	N_N4167<=N_N4166;

 always  @(posedge PCLK)
	N_N3800<=N_N3201;

 always  @(posedge PCLK)
	N_N4237<=N_N3192;

 always  @(posedge PCLK)
	N_N3417<=N_N3416;

 always  @(posedge PCLK)
	N_N3918<=N_N3592;

 always  @(posedge PCLK)
	N_N4158<=N_N3437;

 always  @(posedge PCLK)
	N_N3630<=N_N2976;

 always  @(posedge PCLK)
	N_N3344<=N_N3103;

 always  @(posedge PCLK)
	N_N4072<=N_N3206;

 always  @(posedge PCLK)
	N_N3274<=N_N3273;

 always  @(posedge PCLK)
	N_N3473<=N_N3472;

 always  @(posedge PCLK)
	N_N4205<=N_N3511;

 always  @(posedge PCLK)
	N_N4111<=N_N4110;

 always  @(posedge PCLK)
	N_N3680<=N_N3008;

 always  @(posedge PCLK)
	N_N3838<=N_N3432;

 always  @(posedge PCLK)
	N_N3262<=N_N2984;

 always  @(posedge PCLK)
	N_N4099<=N_N4098;

 always  @(posedge PCLK)
	N_N3607<=N_N2975;

 always  @(posedge PCLK)
	N_N3323<=N_N3320;

 always  @(posedge PCLK)
	N_N3612<=N_N3611;

 always  @(posedge PCLK)
	N_N4079<=N_N4032;

 always  @(posedge PCLK)
	PDN<=N_N3620;

 always  @(posedge PCLK)
	N_N3457<=N_N3102;

 always  @(posedge PCLK)
	N_N3445<=N_N3155;

 always  @(posedge PCLK)
	N_N3794<=N_N3559;

 always  @(posedge PCLK)
	N_N3663<=N_N3662;

 always  @(posedge PCLK)
	N_N3715<=N_N3007;

 always  @(posedge PCLK)
	N_N4039<=N_N4038;

 always  @(posedge PCLK)
	N_N3280<=N_N2983;

 always  @(posedge PCLK)
	N_N4239<=N_N4238;

 always  @(posedge PCLK)
	N_N3988<=N_N3987;

 always  @(posedge PCLK)
	N_N3433<=N_N3172;

 always  @(posedge PCLK)
	N_N4075<=N_N4074;

 always  @(posedge PCLK)
	N_N3468<=N_N3038;

 always  @(posedge PCLK)
	N_N4045<=N_N4044;

 always  @(posedge PCLK)
	N_N3482<=N_N3481;

 always  @(posedge PCLK)
	N_N3832<=N_N3086;

 always  @(posedge PCLK)
	N_N3304<=N_N3210;

 always  @(posedge PCLK)
	N_N3750<=N_N3040;

 always  @(posedge PCLK)
	N_N3634<=N_N3633;

 always  @(posedge PCLK)
	N_N3293<=N_N3177;

 always  @(posedge PCLK)
	N_N3659<=N_N3658;

 always  @(posedge PCLK)
	N_N4252<=N_N3671;

 always  @(posedge PCLK)
	N_N3912<=N_N3449;

 always  @(posedge PCLK)
	N_N3862<=N_N3117;

 always  @(posedge PCLK)
	N_N3221<=N_N3209;

 always  @(posedge PCLK)
	N_N3875<=N_N3113;

 always  @(posedge PCLK)
	N_N3949<=N_N3602;

 always  @(posedge PCLK)
	N_N3908<=N_N3322;

 always  @(posedge PCLK)
	N_N3711<=N_N3710;

 always  @(posedge PCLK)
	N_N3931<=N_N3244;

 always  @(posedge PCLK)
	N_N3469<=N_N2996;

 always  @(posedge PCLK)
	N_N3436<=N_N3435;

 always  @(posedge PCLK)
	N_N3974<=N_N3027;

 always  @(posedge PCLK)
	N_N3905<=N_N3904;

 always  @(posedge PCLK)
	N_N3741<=N_N3740;

 always  @(posedge PCLK)
	N_N3369<=N_N3165;

 always  @(posedge PCLK)
	N_N3164<=N_N3144;

 always  @(posedge PCLK)
	N_N3500<=N_N3499;

 always  @(posedge PCLK)
	N_N3996<=N_N3200;

 always  @(posedge PCLK)
	N_N3356<=N_N2979;

 always  @(posedge PCLK)
	N_N4093<=N_N3147;

 always  @(posedge PCLK)
	Pover_0_0_<=N_N3061;

 always  @(posedge PCLK)
	N_N4224<=N_N3586;

 always  @(posedge PCLK)
	N_N4027<=N_N2980;

 always  @(posedge PCLK)
	NDN1_4<=N_N3305;

 always  @(posedge PCLK)
	N_N3384<=N_N2978;

 always  @(posedge PCLK)
	N_N4036<=N_N3093;

 always  @(posedge PCLK)
	N_N3968<=N_N3967;

 always  @(posedge PCLK)
	N_N4183<=N_N3190;

 always  @(posedge PCLK)
	NGFDN_3<=N_N3542;

 always  @(posedge PCLK)
	N_N4090<=N_N4089;

 always  @(posedge PCLK)
	N_N4004<=N_N3091;

 always  @(posedge PCLK)
	N_N3205<=N_N3204;

 always  @(posedge PCLK)
	N_N4136<=N_N3191;

 always  @(posedge PCLK)
	N_N3303<=N_N3101;

 always  @(posedge PCLK)
	N_N3533<=N_N3352;

 always  @(posedge PCLK)
	N_N3336<=N_N3335;

 always  @(posedge PCLK)
	N_N3961<=N_N2964;

 always  @(posedge PCLK)
	N_N3331<=N_N3057;

 always  @(posedge PCLK)
	N_N3203<=N_N3202;

 always  @(posedge PCLK)
	N_N4236<=N_N4028;

 always  @(posedge PCLK)
	N_N3884<=N_N3321;

 always  @(posedge PCLK)
	N_N3367<=N_N3366;

 always  @(posedge PCLK)
	N_N4140<=N_N4139;

 always  @(posedge PCLK)
	NDN2_2<=N_N3476;

 always  @(posedge PCLK)
	N_N4106<=N_N4105;

 always  @(posedge PCLK)
	N_N3100<=N_N3028;

 always  @(posedge PCLK)
	N_N4193<=N_N3720;

 always  @(posedge PCLK)
	N_N3470<=N_N3034;

 always  @(posedge PCLK)
	N_N3424<=N_N3423;

 always  @(posedge PCLK)
	N_N3959<=N_N3958;

 always  @(posedge PCLK)
	N_N3393<=N_N3318;

 always  @(posedge PCLK)
	N_N4042<=N_N4041;

 always  @(posedge PCLK)
	N_N3188<=N_N3075;

 always  @(posedge PCLK)
	N_N4095<=N_N4094;

 always  @(posedge PCLK)
	N_N3957<=N_N3956;

 always  @(posedge PCLK)
	N_N3517<=N_N3401;

 always  @(posedge PCLK)
	N_N4047<=N_N4046;

 always  @(posedge PCLK)
	N_N3081<=N_N2977;

 always  @(posedge PCLK)
	N_N3541<=N_N2962;

 always  @(posedge PCLK)
	N_N4177<=N_N3087;

 always  @(posedge PCLK)
	NDN3_3<=N_N3530;

 always  @(posedge PCLK)
	N_N4176<=N_N3479;

 always  @(posedge PCLK)
	N_N3585<=N_N3584;

 always  @(posedge PCLK)
	NDN3_8<=N_N3752;

 always  @(posedge PCLK)
	N_N4209<=N_N3503;

 always  @(posedge PCLK)
	N_N3824<=N_N3823;

 always  @(posedge PCLK)
	N_N4208<=N_N3130;

 always  @(posedge PCLK)
	N_N4120<=N_N3895;

 always  @(posedge PCLK)
	N_N3708<=N_N3707;

 always  @(posedge PCLK)
	N_N4220<=N_N3941;

 always  @(posedge PCLK)
	N_N3999<=N_N4254;

 always  @(posedge PCLK)
	N_N4223<=N_N3314;

 always  @(posedge PCLK)
	N_N3179<=N_N3178;

 always  @(posedge PCLK)
	N_N4179<=N_N3963;

 always  @(posedge PCLK)
	N_N3475<=N_N3474;

 always  @(posedge PCLK)
	N_N4132<=N_N3194;

 always  @(posedge PCLK)
	N_N4182<=N_N2958;

 always  @(posedge PCLK)
	N_N3797<=N_N3163;

 always  @(posedge PCLK)
	N_N3214<=N_N3213;

 always  @(posedge PCLK)
	N_N4070<=N_N3193;

 always  @(posedge PCLK)
	N_N4135<=N_N2957;

 always  @(posedge PCLK)
	NLD3_9<=N_N3042;

 always  @(posedge PCLK)
	NDN5_2<=N_N3160;

 always  @(posedge PCLK)
	NDN5_3<=N_N3041;

 always  @(posedge PCLK)
	N_N3778<=N_N3284;

 always  @(posedge PCLK)
	NDN5_4<=N_N3739;

 always  @(posedge PCLK)
	N_N3212<=N_N3211;

 always  @(posedge PCLK)
	NDN5_5<=N_N3348;

 always  @(posedge PCLK)
	NDN5_6<=N_N3016;

 always  @(posedge PCLK)
	NDN5_7<=N_N3538;

 always  @(posedge PCLK)
	NDN5_8<=N_N3029;

 always  @(posedge PCLK)
	N_N4073<=N_N3338;

 always  @(posedge PCLK)
	NDN5_9<=N_N3458;

 always  @(posedge PCLK)
	NEN5_9<=N_N3618;

 always  @(posedge PCLK)
	N_N3684<=N_N3683;

 always  @(posedge PCLK)
	N_N4056<=N_N4055;

 always  @(posedge PCLK)
	N_N3713<=N_N3712;

 always  @(posedge PCLK)
	N_N3829<=N_N3828;

 always  @(posedge PCLK)
	N_N4060<=N_N47;

 always  @(posedge PCLK)
	NSr3_2<=N_N46;

 always  @(posedge PCLK)
	NSr5_2<=N_N45;

 always  @(posedge PCLK)
	NSr5_3<=N_N44;

 always  @(posedge PCLK)
	N_N3462<=N_N43;

 always  @(posedge PCLK)
	N_N3460<=N_N42;

 always  @(posedge PCLK)
	NSr5_4<=N_N41;

 always  @(posedge PCLK)
	NSr3_9<=N_N40;

 always  @(posedge PCLK)
	NSr5_5<=N_N39;

 always  @(posedge PCLK)
	NSr5_7<=N_N38;

 always  @(posedge PCLK)
	NSr5_8<=N_N37;

 always  @(posedge PCLK)
	N_N3998<=N_N36;

 assign n3 = ( (~ PRESET)  &  n410 ) ;
 assign n2 = ( N_N3460  &  (~ n411)  &  n412 ) ;
 assign N_N4254 = ( n3  &  n2 ) | ( n3  &  N_N3999 ) ;
 assign n4 = ( PRESET  &  n463 ) | ( n458  &  n463 ) | ( PRESET  &  (~ N_N4239) ) | ( n458  &  (~ N_N4239) ) ;
 assign N_N4238 = ( (~ n4) ) ;
 assign n5 = ( n464 ) | ( (~ N_N4232) ) ;
 assign N_N4231 = ( (~ n5) ) ;
 assign n6 = ( n464 ) | ( (~ N_N4230) ) ;
 assign N_N4229 = ( (~ n6) ) ;
 assign n7 = ( n464 ) | ( (~ N_N4218) ) ;
 assign N_N4217 = ( (~ n7) ) ;
 assign n8 = ( (~ PRESET)  &  n1235 ) ;
 assign N_N4174 = ( N_N4222  &  n8 ) ;
 assign n9 = ( n591  &  (~ n1237) ) | ( (~ n1194)  &  (~ n1237) ) | ( n591  &  (~ N_N4167) ) | ( (~ n1194)  &  (~ N_N4167) ) ;
 assign N_N4166 = ( (~ n9) ) ;
 assign n11 = ( PRESET  &  n463 ) | ( n463  &  n594 ) | ( PRESET  &  (~ N_N4140) ) | ( n594  &  (~ N_N4140) ) ;
 assign N_N4139 = ( (~ n11) ) ;
 assign n12 = ( n597  &  n599 ) | ( n597  &  (~ n1194) ) | ( n599  &  (~ N_N4114) ) | ( (~ n1194)  &  (~ N_N4114) ) ;
 assign N_N4113 = ( (~ n12) ) ;
 assign n13 = ( n607  &  n609 ) | ( n607  &  n610 ) | ( n609  &  (~ N_N4111) ) | ( n610  &  (~ N_N4111) ) ;
 assign N_N4110 = ( (~ n13) ) ;
 assign n14 = ( n464 ) | ( (~ N_N4106) ) ;
 assign N_N4105 = ( (~ n14) ) ;
 assign n15 = ( PRESET  &  n463 ) | ( n463  &  n613 ) | ( PRESET  &  (~ N_N4099) ) | ( n613  &  (~ N_N4099) ) ;
 assign N_N4098 = ( (~ n15) ) ;
 assign n16 = ( PRESET  &  n463 ) | ( n463  &  n618 ) | ( PRESET  &  (~ N_N4095) ) | ( n618  &  (~ N_N4095) ) ;
 assign N_N4094 = ( (~ n16) ) ;
 assign n17 = ( n464 ) | ( (~ N_N4090) ) ;
 assign N_N4089 = ( (~ n17) ) ;
 assign n18 = ( PRESET  &  n463 ) | ( n463  &  n621 ) | ( PRESET  &  (~ N_N4086) ) | ( n621  &  (~ N_N4086) ) ;
 assign N_N4085 = ( (~ n18) ) ;
 assign n19 = ( n624  &  n625 ) | ( n624  &  n626 ) | ( n625  &  (~ N_N4075) ) | ( n626  &  (~ N_N4075) ) ;
 assign N_N4074 = ( (~ n19) ) ;
 assign n22 = ( (~ Paport_5_5_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Paport_5_5_)  &  (~ N_N4056) ) | ( n466  &  (~ N_N4056) ) ;
 assign N_N4055 = ( (~ n22) ) ;
 assign n23 = ( (~ Paport_7_7_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Paport_7_7_)  &  (~ N_N4054) ) | ( n466  &  (~ N_N4054) ) ;
 assign N_N4053 = ( (~ n23) ) ;
 assign n24 = ( n635  &  n636 ) | ( n635  &  n637 ) | ( n636  &  (~ N_N4047) ) | ( n637  &  (~ N_N4047) ) ;
 assign N_N4046 = ( (~ n24) ) ;
 assign n25 = ( n626  &  n635 ) | ( n635  &  n636 ) | ( n626  &  (~ N_N4045) ) | ( n636  &  (~ N_N4045) ) ;
 assign N_N4044 = ( (~ n25) ) ;
 assign n26 = ( n638  &  n639 ) | ( n638  &  n640 ) | ( n639  &  (~ N_N4042) ) | ( n640  &  (~ N_N4042) ) ;
 assign N_N4041 = ( (~ n26) ) ;
 assign n27 = ( n638  &  n639 ) | ( n638  &  n641 ) | ( n639  &  (~ N_N4039) ) | ( n641  &  (~ N_N4039) ) ;
 assign N_N4038 = ( (~ n27) ) ;
 assign n28 = ( n597  &  n599 ) | ( n597  &  n722 ) | ( n599  &  (~ N_N4079) ) | ( n722  &  (~ N_N4079) ) ;
 assign N_N4032 = ( (~ n28) ) ;
 assign n29 = ( n724  &  n725 ) | ( n724  &  n726 ) | ( n725  &  (~ N_N4030) ) | ( n726  &  (~ N_N4030) ) ;
 assign N_N4029 = ( (~ n29) ) ;
 assign n30 = ( n641  &  n727 ) | ( n727  &  n729 ) | ( n641  &  (~ N_N4236) ) | ( n729  &  (~ N_N4236) ) ;
 assign N_N4028 = ( (~ n30) ) ;
 assign n31 = ( n624  &  n625 ) | ( n624  &  n730 ) | ( n625  &  (~ N_N4024) ) | ( n730  &  (~ N_N4024) ) ;
 assign N_N4023 = ( (~ n31) ) ;
 assign n32 = ( n624  &  n625 ) | ( n624  &  n731 ) | ( n625  &  (~ N_N4021) ) | ( n731  &  (~ N_N4021) ) ;
 assign N_N4020 = ( (~ n32) ) ;
 assign n34 = ( (~ Pdxport_2_2_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Pdxport_2_2_)  &  (~ N_N4057) ) | ( n466  &  (~ N_N4057) ) ;
 assign N_N4007 = ( (~ n34) ) ;
 assign n35 = ( n773  &  n775 ) | ( n773  &  n776 ) | ( n775  &  (~ N_N3988) ) | ( n776  &  (~ N_N3988) ) ;
 assign N_N3987 = ( (~ n35) ) ;
 assign n36 = ( n607  &  n610 ) | ( n610  &  (~ N_N3981) ) | ( n607  &  n778 ) | ( (~ N_N3981)  &  n778 ) ;
 assign N_N3980 = ( (~ n36) ) ;
 assign n38 = ( n635  &  n636 ) | ( n635  &  n781 ) | ( n636  &  (~ N_N4116) ) | ( n781  &  (~ N_N4116) ) ;
 assign N_N3969 = ( (~ n38) ) ;
 assign n39 = ( n638  &  n639 ) | ( n638  &  n781 ) | ( n639  &  (~ N_N3968) ) | ( n781  &  (~ N_N3968) ) ;
 assign N_N3967 = ( (~ n39) ) ;
 assign n40 = ( (~ Pdxport_5_5_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Pdxport_5_5_)  &  (~ N_N4179) ) | ( n466  &  (~ N_N4179) ) ;
 assign N_N3963 = ( (~ n40) ) ;
 assign n41 = ( n624  &  n625 ) | ( n624  &  n781 ) | ( n625  &  (~ N_N3959) ) | ( n781  &  (~ N_N3959) ) ;
 assign N_N3958 = ( (~ n41) ) ;
 assign n42 = ( n624  &  n625 ) | ( n624  &  n783 ) | ( n625  &  (~ N_N3957) ) | ( n783  &  (~ N_N3957) ) ;
 assign N_N3956 = ( (~ n42) ) ;
 assign n43 = ( n591  &  (~ n1237) ) | ( n784  &  (~ n1237) ) | ( n591  &  (~ N_N3947) ) | ( n784  &  (~ N_N3947) ) ;
 assign N_N3946 = ( (~ n43) ) ;
 assign n44 = ( (~ Pdxport_3_3_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Pdxport_3_3_)  &  (~ N_N4220) ) | ( n466  &  (~ N_N4220) ) ;
 assign N_N3941 = ( (~ n44) ) ;
 assign n46 = ( (~ Paport_0_0_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Paport_0_0_)  &  (~ N_N3916) ) | ( n466  &  (~ N_N3916) ) ;
 assign N_N3915 = ( (~ n46) ) ;
 assign n47 = ( (~ Paport_6_6_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Paport_6_6_)  &  (~ N_N4243) ) | ( n466  &  (~ N_N4243) ) ;
 assign N_N3914 = ( (~ n47) ) ;
 assign n48 = ( (~ Paport_8_8_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Paport_8_8_)  &  (~ N_N4015) ) | ( n466  &  (~ N_N4015) ) ;
 assign N_N3913 = ( (~ n48) ) ;
 assign n49 = ( n727  &  n729 ) | ( n727  &  n793 ) | ( n729  &  (~ N_N3910) ) | ( n793  &  (~ N_N3910) ) ;
 assign N_N3909 = ( (~ n49) ) ;
 assign N_N3904 = ( N_N3905  &  n8 ) ;
 assign n51 = ( (~ Pdxport_1_1_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Pdxport_1_1_)  &  (~ N_N4120) ) | ( n466  &  (~ N_N4120) ) ;
 assign N_N3895 = ( (~ n51) ) ;
 assign n56 = ( n885  &  n887 ) | ( n886  &  n887 ) | ( n885  &  (~ N_N4197) ) | ( n886  &  (~ N_N4197) ) ;
 assign N_N3847 = ( (~ n56) ) ;
 assign n57 = ( n591  &  (~ n1237) ) | ( n888  &  (~ n1237) ) | ( n591  &  (~ N_N3829) ) | ( n888  &  (~ N_N3829) ) ;
 assign N_N3828 = ( (~ n57) ) ;
 assign n58 = ( n591  &  (~ n1237) ) | ( n889  &  (~ n1237) ) | ( n591  &  (~ N_N3826) ) | ( n889  &  (~ N_N3826) ) ;
 assign N_N3825 = ( (~ n58) ) ;
 assign n59 = ( n624  &  n625 ) | ( n624  &  n640 ) | ( n625  &  (~ N_N3824) ) | ( n640  &  (~ N_N3824) ) ;
 assign N_N3823 = ( (~ n59) ) ;
 assign n60 = ( (~ Paport_9_9_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Paport_9_9_)  &  (~ N_N3818) ) | ( n466  &  (~ N_N3818) ) ;
 assign N_N3817 = ( (~ n60) ) ;
 assign n61 = ( n591  &  (~ n1237) ) | ( n892  &  (~ n1237) ) | ( n591  &  (~ N_N3815) ) | ( n892  &  (~ N_N3815) ) ;
 assign N_N3814 = ( (~ n61) ) ;
 assign n62 = ( n464 ) | ( (~ N_N3876) ) ;
 assign N_N3804 = ( (~ n62) ) ;
 assign n63 = ( PRESET  &  n463 ) | ( n463  &  n895 ) | ( PRESET  &  (~ N_N3971) ) | ( n895  &  (~ N_N3971) ) ;
 assign N_N3801 = ( (~ n63) ) ;
 assign n64 = ( n638  &  n639 ) | ( n638  &  n730 ) | ( n639  &  (~ N_N3799) ) | ( n730  &  (~ N_N3799) ) ;
 assign N_N3798 = ( (~ n64) ) ;
 assign n65 = ( n591  &  (~ n1237) ) | ( n899  &  (~ n1237) ) | ( n591  &  (~ N_N3796) ) | ( n899  &  (~ N_N3796) ) ;
 assign N_N3795 = ( (~ n65) ) ;
 assign n66 = ( n591  &  (~ n1237) ) | ( n900  &  (~ n1237) ) | ( n591  &  (~ N_N3788) ) | ( n900  &  (~ N_N3788) ) ;
 assign N_N3787 = ( (~ n66) ) ;
 assign n67 = ( n464 ) | ( (~ N_N3786) ) ;
 assign N_N3785 = ( (~ n67) ) ;
 assign n68 = ( n635  &  n636 ) | ( n635  &  n726 ) | ( n636  &  (~ N_N3870) ) | ( n726  &  (~ N_N3870) ) ;
 assign N_N3772 = ( (~ n68) ) ;
 assign n72 = ( (~ PRESET)  &  (~ NGFDN_3) ) ;
 assign N_N3752 = ( n72  &  NDN3_8 ) | ( n72  &  NDN3_3 ) ;
 assign n73 = ( PRESET  &  n909 ) | ( n909  &  (~ N_N3745) ) ;
 assign N_N3744 = ( (~ n73) ) ;
 assign n74 = ( n464 ) | ( (~ N_N3741) ) ;
 assign N_N3740 = ( (~ n74) ) ;
 assign N_N3739 = ( (~ PRESET)  &  (~ NSr5_4) ) ;
 assign n78 = ( n886  &  n887 ) | ( n887  &  n914 ) | ( n886  &  (~ N_N3992) ) | ( n914  &  (~ N_N3992) ) ;
 assign N_N3723 = ( (~ n78) ) ;
 assign n80 = ( n626  &  n727 ) | ( n727  &  n729 ) | ( n626  &  (~ N_N4193) ) | ( n729  &  (~ N_N4193) ) ;
 assign N_N3720 = ( (~ n80) ) ;
 assign n81 = ( n886  &  n887 ) | ( n887  &  n916 ) | ( n886  &  (~ N_N4018) ) | ( n916  &  (~ N_N4018) ) ;
 assign N_N3717 = ( (~ n81) ) ;
 assign n82 = ( n597  &  n599 ) | ( n597  &  n918 ) | ( n599  &  (~ N_N3713) ) | ( n918  &  (~ N_N3713) ) ;
 assign N_N3712 = ( (~ n82) ) ;
 assign n83 = ( n724  &  n725 ) | ( n724  &  n731 ) | ( n725  &  (~ N_N3711) ) | ( n731  &  (~ N_N3711) ) ;
 assign N_N3710 = ( (~ n83) ) ;
 assign N_N3707 = ( N_N3708  &  n8 ) ;
 assign n84 = ( (~ Paport_10_10_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Paport_10_10_)  &  (~ N_N3882) ) | ( n466  &  (~ N_N3882) ) ;
 assign N_N3705 = ( (~ n84) ) ;
 assign n86 = ( n727  &  n729 ) | ( n727  &  n730 ) | ( n729  &  (~ N_N3793) ) | ( n730  &  (~ N_N3793) ) ;
 assign N_N3695 = ( (~ n86) ) ;
 assign N_N3690 = ( N_N3691  &  n8 ) ;
 assign n89 = ( n591  &  (~ n1237) ) | ( n926  &  (~ n1237) ) | ( n591  &  (~ N_N3684) ) | ( n926  &  (~ N_N3684) ) ;
 assign N_N3683 = ( (~ n89) ) ;
 assign n90 = ( PRESET  &  n463 ) | ( n463  &  n927 ) | ( PRESET  &  (~ N_N4252) ) | ( n927  &  (~ N_N4252) ) ;
 assign N_N3671 = ( (~ n90) ) ;
 assign n91 = ( PRESET  &  n463 ) | ( n463  &  n930 ) | ( PRESET  &  (~ N_N3843) ) | ( n930  &  (~ N_N3843) ) ;
 assign N_N3668 = ( (~ n91) ) ;
 assign n92 = ( n597  &  n599 ) | ( n597  &  n932 ) | ( n599  &  (~ N_N3743) ) | ( n932  &  (~ N_N3743) ) ;
 assign N_N3666 = ( (~ n92) ) ;
 assign n93 = ( n597  &  n599 ) | ( n597  &  n934 ) | ( n599  &  (~ N_N3774) ) | ( n934  &  (~ N_N3774) ) ;
 assign N_N3664 = ( (~ n93) ) ;
 assign n94 = ( n641  &  n773 ) | ( n773  &  n775 ) | ( n641  &  (~ N_N3663) ) | ( n775  &  (~ N_N3663) ) ;
 assign N_N3662 = ( (~ n94) ) ;
 assign n95 = ( n724  &  n725 ) | ( n724  &  n781 ) | ( n725  &  (~ N_N4117) ) | ( n781  &  (~ N_N4117) ) ;
 assign N_N3661 = ( (~ n95) ) ;
 assign n96 = ( n635  &  n636 ) | ( n635  &  n641 ) | ( n636  &  (~ N_N3659) ) | ( n641  &  (~ N_N3659) ) ;
 assign N_N3658 = ( (~ n96) ) ;
 assign n97 = ( n597  &  n599 ) | ( n597  &  n935 ) | ( n599  &  (~ N_N3791) ) | ( n935  &  (~ N_N3791) ) ;
 assign N_N3653 = ( (~ n97) ) ;
 assign n98 = ( n724  &  n725 ) | ( n724  &  n783 ) | ( n725  &  (~ N_N3922) ) | ( n783  &  (~ N_N3922) ) ;
 assign N_N3652 = ( (~ n98) ) ;
 assign n102 = ( n607  &  n610 ) | ( n607  &  n939 ) | ( n610  &  (~ N_N3761) ) | ( n939  &  (~ N_N3761) ) ;
 assign N_N3640 = ( (~ n102) ) ;
 assign N_N3638 = ( (~ PRESET)  &  (~ n410) ) ;
 assign n104 = ( n464 ) | ( (~ N_N3634) ) ;
 assign N_N3633 = ( (~ n104) ) ;
 assign n108 = ( N_N3336  &  n769 ) | ( N_N3336  &  n771 ) | ( n769  &  (~ N_N4205) ) | ( n771  &  (~ N_N4205) ) ;
 assign n106 = ( NLD3_9  &  n108 ) | ( NLD3_9  &  N_N3336  &  (~ N_N4205) ) ;
 assign N_N3811 = ( (~ PRESET)  &  (~ PDN) ) ;
 assign N_N3620 = ( N_N3811  &  NGFDN_3 ) | ( N_N3811  &  (~ n149) ) ;
 assign n111 = ( NLD3_9  &  n944 ) | ( n944  &  n946 ) | ( NLD3_9  &  (~ NEN5_9) ) | ( n946  &  (~ NEN5_9) ) ;
 assign N_N3618 = ( (~ n111) ) ;
 assign n112 = ( n597  &  n599 ) | ( n597  &  n947 ) | ( n599  &  (~ N_N3709) ) | ( n947  &  (~ N_N3709) ) ;
 assign N_N3616 = ( (~ n112) ) ;
 assign n113 = ( n640  &  n773 ) | ( n773  &  n775 ) | ( n640  &  (~ N_N4071) ) | ( n775  &  (~ N_N4071) ) ;
 assign N_N3615 = ( (~ n113) ) ;
 assign n114 = ( n727  &  n729 ) | ( n727  &  n731 ) | ( n729  &  (~ N_N3776) ) | ( n731  &  (~ N_N3776) ) ;
 assign N_N3614 = ( (~ n114) ) ;
 assign n115 = ( n624  &  n625 ) | ( n624  &  n641 ) | ( n625  &  (~ N_N3612) ) | ( n641  &  (~ N_N3612) ) ;
 assign N_N3611 = ( (~ n115) ) ;
 assign n118 = ( n886  &  n887 ) | ( n887  &  n950 ) | ( n886  &  (~ N_N3949) ) | ( n950  &  (~ N_N3949) ) ;
 assign N_N3602 = ( (~ n118) ) ;
 assign n119 = ( PRESET  &  n956 ) | ( n954  &  n956 ) | ( PRESET  &  (~ N_N4212) ) | ( n954  &  (~ N_N4212) ) ;
 assign N_N3599 = ( (~ n119) ) ;
 assign n120 = ( PRESET  &  n956 ) | ( n956  &  n957 ) | ( PRESET  &  (~ N_N4171) ) | ( n957  &  (~ N_N4171) ) ;
 assign N_N3596 = ( (~ n120) ) ;
 assign n121 = ( (~ Paport_2_2_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Paport_2_2_)  &  (~ N_N3733) ) | ( n466  &  (~ N_N3733) ) ;
 assign N_N3595 = ( (~ n121) ) ;
 assign n122 = ( PRESET  &  n463 ) | ( n463  &  n960 ) | ( PRESET  &  (~ N_N3918) ) | ( n960  &  (~ N_N3918) ) ;
 assign N_N3592 = ( (~ n122) ) ;
 assign n123 = ( PRESET  &  n463 ) | ( n463  &  n962 ) | ( PRESET  &  (~ N_N3939) ) | ( n962  &  (~ N_N3939) ) ;
 assign N_N3589 = ( (~ n123) ) ;
 assign n124 = ( PRESET  &  n463 ) | ( n463  &  n964 ) | ( PRESET  &  (~ N_N4224) ) | ( n964  &  (~ N_N4224) ) ;
 assign N_N3586 = ( (~ n124) ) ;
 assign n125 = ( n624  &  n625 ) | ( n624  &  n966 ) | ( n625  &  (~ N_N3585) ) | ( n966  &  (~ N_N3585) ) ;
 assign N_N3584 = ( (~ n125) ) ;
 assign n126 = ( n464 ) | ( (~ N_N3580) ) ;
 assign N_N3579 = ( (~ n126) ) ;
 assign n127 = ( n971  &  n969 ) | ( n971  &  (~ N_N3751) ) ;
 assign N_N3570 = ( (~ n127) ) ;
 assign n130 = ( n607  &  n610 ) | ( n610  &  (~ N_N3794) ) | ( n607  &  n947 ) | ( (~ N_N3794)  &  n947 ) ;
 assign N_N3559 = ( (~ n130) ) ;
 assign n131 = ( n624  &  n625 ) | ( n624  &  n793 ) | ( n625  &  (~ N_N3625) ) | ( n793  &  (~ N_N3625) ) ;
 assign N_N3558 = ( (~ n131) ) ;
 assign N_N3530 = ( n72  &  NDN3_3 ) | ( n72  &  (~ NSr3_2) ) ;
 assign n135 = ( n635  &  n636 ) | ( n635  &  n783 ) | ( n636  &  (~ N_N3921) ) | ( n783  &  (~ N_N3921) ) ;
 assign N_N3524 = ( (~ n135) ) ;
 assign n136 = ( (~ Paport_4_4_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Paport_4_4_)  &  (~ N_N3574) ) | ( n466  &  (~ N_N3574) ) ;
 assign N_N3523 = ( (~ n136) ) ;
 assign n137 = ( (~ Paport_11_11_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Paport_11_11_)  &  (~ N_N4205) ) | ( n466  &  (~ N_N4205) ) ;
 assign N_N3511 = ( (~ n137) ) ;
 assign n138 = ( PRESET  &  n463 ) | ( n463  &  n979 ) | ( PRESET  &  (~ N_N4118) ) | ( n979  &  (~ N_N4118) ) ;
 assign N_N3506 = ( (~ n138) ) ;
 assign n139 = ( PRESET  &  n463 ) | ( n463  &  n981 ) | ( PRESET  &  (~ N_N4209) ) | ( n981  &  (~ N_N4209) ) ;
 assign N_N3503 = ( (~ n139) ) ;
 assign n140 = ( PRESET  &  n463 ) | ( n463  &  n985 ) | ( PRESET  &  (~ N_N3500) ) | ( n985  &  (~ N_N3500) ) ;
 assign N_N3499 = ( (~ n140) ) ;
 assign n143 = ( n607  &  n610 ) | ( n610  &  (~ N_N3489) ) | ( n607  &  n991 ) | ( (~ N_N3489)  &  n991 ) ;
 assign N_N3488 = ( (~ n143) ) ;
 assign n144 = ( n607  &  n610 ) | ( n607  &  n918 ) | ( n610  &  (~ N_N3513) ) | ( n918  &  (~ N_N3513) ) ;
 assign N_N3487 = ( (~ n144) ) ;
 assign n145 = ( n773  &  n775 ) | ( n773  &  n783 ) | ( n775  &  (~ N_N4221) ) | ( n783  &  (~ N_N4221) ) ;
 assign N_N3486 = ( (~ n145) ) ;
 assign n146 = ( (~ Pdxport_6_6_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Pdxport_6_6_)  &  (~ N_N4206) ) | ( n466  &  (~ N_N4206) ) ;
 assign N_N3483 = ( (~ n146) ) ;
 assign n147 = ( n626  &  n638 ) | ( n638  &  n639 ) | ( n626  &  (~ N_N3482) ) | ( n639  &  (~ N_N3482) ) ;
 assign N_N3481 = ( (~ n147) ) ;
 assign n148 = ( n969  &  n994 ) | ( n994  &  (~ N_N4080) ) ;
 assign N_N3479 = ( (~ n148) ) ;
 assign n149 = ( (~ Preset_0_0_) ) | ( PDN ) | ( NLC1_2 ) ;
 assign N_N3476 = ( (~ PRESET)  &  n149  &  NDN2_2 ) ;
 assign n150 = ( n597  &  n599 ) | ( n597  &  n778 ) | ( n599  &  (~ N_N3475) ) | ( n778  &  (~ N_N3475) ) ;
 assign N_N3474 = ( (~ n150) ) ;
 assign n151 = ( n626  &  n773 ) | ( n773  &  n775 ) | ( n626  &  (~ N_N3473) ) | ( n775  &  (~ N_N3473) ) ;
 assign N_N3472 = ( (~ n151) ) ;
 assign N_N3465 = ( (~ PRESET)  &  n106 ) ;
 assign n152 = ( n944  &  (~ N_N3042) ) | ( (~ N_N3042)  &  (~ NEN5_9) ) ;
 assign N_N3458 = ( (~ n152) ) ;
 assign n153 = ( n637  &  n638 ) | ( n638  &  n639 ) | ( n637  &  (~ N_N3736) ) | ( n639  &  (~ N_N3736) ) ;
 assign N_N3456 = ( (~ n153) ) ;
 assign n154 = ( n607  &  n610 ) | ( n610  &  (~ N_N3535) ) | ( n607  &  n997 ) | ( (~ N_N3535)  &  n997 ) ;
 assign N_N3454 = ( (~ n154) ) ;
 assign n156 = ( n886  &  n887 ) | ( n887  &  n999 ) | ( n886  &  (~ N_N3912) ) | ( n999  &  (~ N_N3912) ) ;
 assign N_N3449 = ( (~ n156) ) ;
 assign n158 = ( n597  &  n599 ) | ( n597  &  n1007 ) | ( n599  &  (~ N_N4158) ) | ( n1007  &  (~ N_N4158) ) ;
 assign N_N3437 = ( (~ n158) ) ;
 assign n159 = ( n724  &  n725 ) | ( n724  &  n776 ) | ( n725  &  (~ N_N3436) ) | ( n776  &  (~ N_N3436) ) ;
 assign N_N3435 = ( (~ n159) ) ;
 assign N_N3432 = ( (~ PRESET)  &  n2 ) | ( (~ PRESET)  &  N_N3838 ) ;
 assign n160 = ( n724  &  n725 ) | ( n724  &  n966 ) | ( n725  &  (~ N_N3841) ) | ( n966  &  (~ N_N3841) ) ;
 assign N_N3431 = ( (~ n160) ) ;
 assign N_N3425 = ( N_N3426  &  n8 ) ;
 assign n162 = ( n635  &  n636 ) | ( n635  &  n731 ) | ( n636  &  (~ N_N3424) ) | ( n731  &  (~ N_N3424) ) ;
 assign N_N3423 = ( (~ n162) ) ;
 assign n163 = ( n464 ) | ( (~ N_N3417) ) ;
 assign N_N3416 = ( (~ n163) ) ;
 assign n164 = ( PRESET  &  n463 ) | ( n463  &  n1012 ) | ( PRESET  &  (~ N_N3842) ) | ( n1012  &  (~ N_N3842) ) ;
 assign N_N3413 = ( (~ n164) ) ;
 assign n165 = ( PRESET  &  n463 ) | ( n463  &  n1015 ) | ( PRESET  &  (~ N_N3924) ) | ( n1015  &  (~ N_N3924) ) ;
 assign N_N3409 = ( (~ n165) ) ;
 assign n166 = ( PRESET  &  n463 ) | ( n463  &  n1017 ) | ( PRESET  &  (~ N_N4119) ) | ( n1017  &  (~ N_N4119) ) ;
 assign N_N3406 = ( (~ n166) ) ;
 assign n167 = ( n464 ) | ( (~ N_N3517) ) ;
 assign N_N3401 = ( (~ n167) ) ;
 assign n168 = ( n464 ) | ( (~ N_N3681) ) ;
 assign N_N3400 = ( (~ n168) ) ;
 assign n169 = ( n464 ) | ( (~ N_N3716) ) ;
 assign N_N3399 = ( (~ n169) ) ;
 assign N_N3390 = ( N_N4181  &  n8 ) ;
 assign N_N3389 = ( N_N3578  &  n3 ) ;
 assign N_N3374 = ( N_N3375  &  n8 ) ;
 assign n172 = ( n464 ) | ( (~ N_N3373) ) ;
 assign N_N3372 = ( (~ n172) ) ;
 assign n173 = ( n635  &  n636 ) | ( n635  &  n730 ) | ( n636  &  (~ N_N3367) ) | ( n730  &  (~ N_N3367) ) ;
 assign N_N3366 = ( (~ n173) ) ;
 assign n175 = ( n464 ) | ( (~ N_N3533) ) ;
 assign N_N3352 = ( (~ n175) ) ;
 assign n176 = ( PRESET  &  n463 ) | ( n463  &  n1030 ) | ( PRESET  &  (~ N_N3808) ) | ( n1030  &  (~ N_N3808) ) ;
 assign N_N3349 = ( (~ n176) ) ;
 assign N_N3348 = ( (~ PRESET)  &  (~ NSr5_5) ) ;
 assign n178 = ( PRESET  &  n956 ) | ( n956  &  n1032 ) | ( PRESET  &  (~ N_N3340) ) | ( n1032  &  (~ N_N3340) ) ;
 assign N_N3339 = ( (~ n178) ) ;
 assign N_N3338 = ( N_N4073  &  n8 ) ;
 assign n179 = ( (~ N_N3336)  &  n610 ) | ( n607  &  n610 ) | ( (~ N_N3336)  &  n1007 ) | ( n607  &  n1007 ) ;
 assign N_N3335 = ( (~ n179) ) ;
 assign n180 = ( n726  &  n773 ) | ( n773  &  n775 ) | ( n726  &  (~ N_N4180) ) | ( n775  &  (~ N_N4180) ) ;
 assign N_N3334 = ( (~ n180) ) ;
 assign n181 = ( (~ PRESET)  &  n1221 ) | ( (~ PRESET)  &  (~ n183)  &  N_N4214 ) ;
 assign N_N3332 = ( n181  &  N_N3462 ) ;
 assign n183 = ( (~ N_N4060)  &  n441  &  n445  &  n449  &  (~ n880)  &  n1033  &  n1128  &  n1226 ) ;
 assign N_N3325 = ( (~ PRESET)  &  n183 ) ;
 assign n184 = ( n607  &  n610 ) | ( n607  &  n935 ) | ( n610  &  (~ N_N3908) ) | ( n935  &  (~ N_N3908) ) ;
 assign N_N3322 = ( (~ n184) ) ;
 assign n185 = ( n607  &  n610 ) | ( n607  &  n722 ) | ( n610  &  (~ N_N3884) ) | ( n722  &  (~ N_N3884) ) ;
 assign N_N3321 = ( (~ n185) ) ;
 assign n186 = ( n731  &  n773 ) | ( n773  &  n775 ) | ( n731  &  (~ N_N3323) ) | ( n775  &  (~ N_N3323) ) ;
 assign N_N3320 = ( (~ n186) ) ;
 assign n187 = ( n464 ) | ( (~ N_N3393) ) ;
 assign N_N3318 = ( (~ n187) ) ;
 assign n188 = ( n969  &  n1041 ) | ( n1041  &  (~ N_N3932) ) ;
 assign N_N3316 = ( (~ n188) ) ;
 assign n189 = ( n969  &  n1042 ) | ( n1042  &  (~ N_N3876) ) ;
 assign N_N3315 = ( (~ n189) ) ;
 assign N_N3314 = ( N_N4223  &  n8 ) ;
 assign n190 = ( n640  &  n727 ) | ( n727  &  n729 ) | ( n640  &  (~ N_N3311) ) | ( n729  &  (~ N_N3311) ) ;
 assign N_N3310 = ( (~ n190) ) ;
 assign N_N3305 = ( NDN1_4  &  N_N3811 ) ;
 assign N_N3287 = ( NDN3_11  &  n72 ) ;
 assign n193 = ( (~ Paport_3_3_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Paport_3_3_)  &  (~ N_N3778) ) | ( n466  &  (~ N_N3778) ) ;
 assign N_N3284 = ( (~ n193) ) ;
 assign n194 = ( n1047  &  n441 ) | ( n1047  &  n886 ) ;
 assign N_N3277 = ( (~ n194) ) ;
 assign n195 = ( n1048  &  n433 ) | ( n1048  &  n886 ) ;
 assign N_N3276 = ( (~ n195) ) ;
 assign n196 = ( n591  &  (~ n1237) ) | ( n1049  &  (~ n1237) ) | ( n591  &  (~ N_N3274) ) | ( n1049  &  (~ N_N3274) ) ;
 assign N_N3273 = ( (~ n196) ) ;
 assign n197 = ( n591  &  (~ n1237) ) | ( n1050  &  (~ n1237) ) | ( n591  &  (~ N_N3480) ) | ( n1050  &  (~ N_N3480) ) ;
 assign N_N3266 = ( (~ n197) ) ;
 assign n198 = ( PRESET  &  n463 ) | ( n463  &  n1051 ) | ( PRESET  &  (~ N_N3940) ) | ( n1051  &  (~ N_N3940) ) ;
 assign N_N3263 = ( (~ n198) ) ;
 assign n199 = ( n624  &  n625 ) | ( n624  &  n776 ) | ( n625  &  (~ N_N3700) ) | ( n776  &  (~ N_N3700) ) ;
 assign N_N3259 = ( (~ n199) ) ;
 assign n200 = ( n464 ) | ( (~ N_N3250) ) ;
 assign N_N3249 = ( (~ n200) ) ;
 assign n201 = ( n464 ) | ( (~ N_N3248) ) ;
 assign N_N3247 = ( (~ n201) ) ;
 assign n203 = ( n597  &  n599 ) | ( n597  &  n784 ) | ( n599  &  (~ N_N3931) ) | ( n784  &  (~ N_N3931) ) ;
 assign N_N3244 = ( (~ n203) ) ;
 assign n204 = ( n591  &  (~ n1237) ) | ( n1058  &  (~ n1237) ) | ( n591  &  (~ N_N3509) ) | ( n1058  &  (~ N_N3509) ) ;
 assign N_N3241 = ( (~ n204) ) ;
 assign n205 = ( n591  &  (~ n1237) ) | ( n1059  &  (~ n1237) ) | ( n591  &  (~ N_N3529) ) | ( n1059  &  (~ N_N3529) ) ;
 assign N_N3240 = ( (~ n205) ) ;
 assign n206 = ( NLD3_9  &  n944 ) | ( n944  &  n1061 ) | ( NLD3_9  &  (~ NDN5_10) ) | ( n1061  &  (~ NDN5_10) ) ;
 assign N_N3231 = ( (~ n206) ) ;
 assign n207 = ( PRESET  &  n463 ) | ( n463  &  n1062 ) | ( PRESET  &  (~ N_N3923) ) | ( n1062  &  (~ N_N3923) ) ;
 assign N_N3227 = ( (~ n207) ) ;
 assign n208 = ( n886  &  n887 ) | ( n887  &  n1064 ) | ( n886  &  (~ N_N4145) ) | ( n1064  &  (~ N_N4145) ) ;
 assign N_N3222 = ( (~ n208) ) ;
 assign n209 = ( n597  &  n599 ) | ( n597  &  n926 ) | ( n599  &  (~ N_N3464) ) | ( n926  &  (~ N_N3464) ) ;
 assign N_N3216 = ( (~ n209) ) ;
 assign n210 = ( n597  &  n599 ) | ( n597  &  n888 ) | ( n599  &  (~ N_N3442) ) | ( n888  &  (~ N_N3442) ) ;
 assign N_N3215 = ( (~ n210) ) ;
 assign n211 = ( n597  &  n599 ) | ( n597  &  n939 ) | ( n599  &  (~ N_N3214) ) | ( n939  &  (~ N_N3214) ) ;
 assign N_N3213 = ( (~ n211) ) ;
 assign n212 = ( n597  &  n599 ) | ( n597  &  n991 ) | ( n599  &  (~ N_N3212) ) | ( n991  &  (~ N_N3212) ) ;
 assign N_N3211 = ( (~ n212) ) ;
 assign n213 = ( n724  &  n725 ) | ( n724  &  n793 ) | ( n725  &  (~ N_N3304) ) | ( n793  &  (~ N_N3304) ) ;
 assign N_N3210 = ( (~ n213) ) ;
 assign n214 = ( n724  &  n725 ) | ( n724  &  n730 ) | ( n725  &  (~ N_N3221) ) | ( n730  &  (~ N_N3221) ) ;
 assign N_N3209 = ( (~ n214) ) ;
 assign N_N3206 = ( N_N4072  &  n8 ) ;
 assign n215 = ( n638  &  n639 ) | ( n638  &  n783 ) | ( n639  &  (~ N_N3205) ) | ( n783  &  (~ N_N3205) ) ;
 assign N_N3204 = ( (~ n215) ) ;
 assign n216 = ( n638  &  n639 ) | ( n638  &  n726 ) | ( n639  &  (~ N_N3203) ) | ( n726  &  (~ N_N3203) ) ;
 assign N_N3202 = ( (~ n216) ) ;
 assign n217 = ( n969  &  n1066 ) | ( n1066  &  (~ N_N3634) ) ;
 assign N_N3201 = ( (~ n217) ) ;
 assign n218 = ( n886  &  n887 ) | ( n887  &  n1067 ) | ( n886  &  (~ N_N3996) ) | ( n1067  &  (~ N_N3996) ) ;
 assign N_N3200 = ( (~ n218) ) ;
 assign n220 = ( (~ Pdxport_7_7_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Pdxport_7_7_)  &  (~ N_N4132) ) | ( n466  &  (~ N_N4132) ) ;
 assign N_N3194 = ( (~ n220) ) ;
 assign n221 = ( (~ Pdxport_9_9_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Pdxport_9_9_)  &  (~ N_N4070) ) | ( n466  &  (~ N_N4070) ) ;
 assign N_N3193 = ( (~ n221) ) ;
 assign n222 = ( (~ Pdxport_11_11_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Pdxport_11_11_)  &  (~ N_N4237) ) | ( n466  &  (~ N_N4237) ) ;
 assign N_N3192 = ( (~ n222) ) ;
 assign n223 = ( n969  &  n1072 ) | ( n1072  &  (~ N_N3517) ) ;
 assign N_N3191 = ( (~ n223) ) ;
 assign n224 = ( n969  &  n1073 ) | ( n1073  &  (~ N_N3393) ) ;
 assign N_N3190 = ( (~ n224) ) ;
 assign n225 = ( n464 ) | ( (~ N_N3932) ) ;
 assign N_N3189 = ( (~ n225) ) ;
 assign n228 = ( n597  &  n599 ) | ( n597  &  n997 ) | ( n599  &  (~ N_N3179) ) | ( n997  &  (~ N_N3179) ) ;
 assign N_N3178 = ( (~ n228) ) ;
 assign n229 = ( n637  &  n773 ) | ( n773  &  n775 ) | ( n637  &  (~ N_N3293) ) | ( n775  &  (~ N_N3293) ) ;
 assign N_N3177 = ( (~ n229) ) ;
 assign n230 = ( n773  &  n775 ) | ( n773  &  n781 ) | ( n775  &  (~ N_N3175) ) | ( n781  &  (~ N_N3175) ) ;
 assign N_N3174 = ( (~ n230) ) ;
 assign n231 = ( n640  &  n724 ) | ( n724  &  n725 ) | ( n640  &  (~ N_N3806) ) | ( n725  &  (~ N_N3806) ) ;
 assign N_N3173 = ( (~ n231) ) ;
 assign n232 = ( n641  &  n724 ) | ( n724  &  n725 ) | ( n641  &  (~ N_N3433) ) | ( n725  &  (~ N_N3433) ) ;
 assign N_N3172 = ( (~ n232) ) ;
 assign n234 = ( PRESET  &  n956 ) | ( n956  &  n1081 ) | ( PRESET  &  (~ N_N3369) ) | ( n1081  &  (~ N_N3369) ) ;
 assign N_N3165 = ( (~ n234) ) ;
 assign n235 = ( (~ Paport_1_1_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Paport_1_1_)  &  (~ N_N3797) ) | ( n466  &  (~ N_N3797) ) ;
 assign N_N3163 = ( (~ n235) ) ;
 assign n236 = ( n638  &  n639 ) | ( n638  &  n793 ) | ( n639  &  (~ N_N3626) ) | ( n793  &  (~ N_N3626) ) ;
 assign N_N3162 = ( (~ n236) ) ;
 assign N_N3160 = ( (~ PRESET)  &  (~ NSr5_2) ) ;
 assign N_N3156 = ( N_N4134  &  n8 ) ;
 assign N_N3155 = ( N_N3445  &  n8 ) ;
 assign n239 = ( n969  &  n1086 ) | ( n1086  &  (~ N_N3280) ) ;
 assign N_N3153 = ( (~ n239) ) ;
 assign n240 = ( n464 ) | ( (~ N_N3196) ) ;
 assign N_N3152 = ( (~ n240) ) ;
 assign n242 = ( PRESET  &  n956 ) | ( n956  &  n1090 ) | ( PRESET  &  (~ N_N4093) ) | ( n1090  &  (~ N_N4093) ) ;
 assign N_N3147 = ( (~ n242) ) ;
 assign n243 = ( (~ Pdxport_4_4_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Pdxport_4_4_)  &  (~ N_N4165) ) | ( n466  &  (~ N_N4165) ) ;
 assign N_N3146 = ( (~ n243) ) ;
 assign n244 = ( n773  &  n775 ) | ( n773  &  n793 ) | ( n775  &  (~ N_N3387) ) | ( n793  &  (~ N_N3387) ) ;
 assign N_N3145 = ( (~ n244) ) ;
 assign n245 = ( n637  &  n724 ) | ( n724  &  n725 ) | ( n637  &  (~ N_N3164) ) | ( n725  &  (~ N_N3164) ) ;
 assign N_N3144 = ( (~ n245) ) ;
 assign n247 = ( n727  &  n729 ) | ( n727  &  n783 ) | ( n729  &  (~ N_N3143) ) | ( n783  &  (~ N_N3143) ) ;
 assign N_N3136 = ( (~ n247) ) ;
 assign n248 = ( n635  &  n636 ) | ( n635  &  n966 ) | ( n636  &  (~ N_N3840) ) | ( n966  &  (~ N_N3840) ) ;
 assign N_N3133 = ( (~ n248) ) ;
 assign n249 = ( n635  &  n636 ) | ( n635  &  n640 ) | ( n636  &  (~ N_N3805) ) | ( n640  &  (~ N_N3805) ) ;
 assign N_N3132 = ( (~ n249) ) ;
 assign n250 = ( n969  &  n1100 ) | ( n1100  &  (~ N_N4159) ) ;
 assign N_N3130 = ( (~ n250) ) ;
 assign n251 = ( n969  &  n1102 ) | ( n1102  &  (~ N_N3235) ) ;
 assign N_N3129 = ( (~ n251) ) ;
 assign n253 = ( PRESET  &  n463 ) | ( n463  &  n1104 ) | ( PRESET  &  (~ N_N3872) ) | ( n1104  &  (~ N_N3872) ) ;
 assign N_N3123 = ( (~ n253) ) ;
 assign N_N3119 = ( N_N3324  &  n8 ) ;
 assign n255 = ( n607  &  n610 ) | ( n610  &  (~ N_N3862) ) | ( n607  &  n934 ) | ( (~ N_N3862)  &  n934 ) ;
 assign N_N3117 = ( (~ n255) ) ;
 assign n256 = ( n464 ) | ( (~ N_N3751) ) ;
 assign N_N3115 = ( (~ n256) ) ;
 assign n257 = ( n597  &  n599 ) | ( n597  &  n1059 ) | ( n599  &  (~ N_N3875) ) | ( n1059  &  (~ N_N3875) ) ;
 assign N_N3113 = ( (~ n257) ) ;
 assign n258 = ( n886  &  n887 ) | ( n887  &  n1108 ) | ( n886  &  (~ N_N3965) ) | ( n1108  &  (~ N_N3965) ) ;
 assign N_N3106 = ( (~ n258) ) ;
 assign n259 = ( n464 ) | ( (~ N_N3105) ) ;
 assign N_N3104 = ( (~ n259) ) ;
 assign n260 = ( n730  &  n773 ) | ( n773  &  n775 ) | ( n730  &  (~ N_N3344) ) | ( n775  &  (~ N_N3344) ) ;
 assign N_N3103 = ( (~ n260) ) ;
 assign n261 = ( n626  &  n724 ) | ( n724  &  n725 ) | ( n626  &  (~ N_N3457) ) | ( n725  &  (~ N_N3457) ) ;
 assign N_N3102 = ( (~ n261) ) ;
 assign n262 = ( n635  &  n636 ) | ( n635  &  n793 ) | ( n636  &  (~ N_N3303) ) | ( n793  &  (~ N_N3303) ) ;
 assign N_N3101 = ( (~ n262) ) ;
 assign n263 = ( n1115  &  n445 ) | ( n1115  &  n886 ) ;
 assign N_N3093 = ( (~ n263) ) ;
 assign n264 = ( n1116  &  n449 ) | ( n1116  &  n886 ) ;
 assign N_N3091 = ( (~ n264) ) ;
 assign n265 = ( PRESET  &  n463 ) | ( n463  &  n1117 ) | ( PRESET  &  (~ N_N4177) ) | ( n1117  &  (~ N_N4177) ) ;
 assign N_N3087 = ( (~ n265) ) ;
 assign n266 = ( n607  &  n610 ) | ( n607  &  n932 ) | ( n610  &  (~ N_N3832) ) | ( n932  &  (~ N_N3832) ) ;
 assign N_N3086 = ( (~ n266) ) ;
 assign N_N3078 = ( N_N3345  &  n8 ) ;
 assign n267 = ( n635  &  n636 ) | ( n635  &  n776 ) | ( n636  &  (~ N_N3188) ) | ( n776  &  (~ N_N3188) ) ;
 assign N_N3075 = ( (~ n267) ) ;
 assign n269 = ( n726  &  n727 ) | ( n727  &  n729 ) | ( n726  &  (~ N_N3071) ) | ( n729  &  (~ N_N3071) ) ;
 assign N_N3070 = ( (~ n269) ) ;
 assign n270 = ( n727  &  n729 ) | ( n727  &  n966 ) | ( n729  &  (~ N_N3069) ) | ( n966  &  (~ N_N3069) ) ;
 assign N_N3068 = ( (~ n270) ) ;
 assign N_N3063 = ( NDN5_16  &  (~ n944) ) ;
 assign n275 = ( n464 ) | ( (~ N_N4159) ) ;
 assign N_N3058 = ( (~ n275) ) ;
 assign n276 = ( n464 ) | ( (~ N_N3331) ) ;
 assign N_N3057 = ( (~ n276) ) ;
 assign n277 = ( PRESET  &  n956 ) | ( n956  &  n1127 ) | ( PRESET  &  (~ N_N3283) ) | ( n1127  &  (~ N_N3283) ) ;
 assign N_N3053 = ( (~ n277) ) ;
 assign n278 = ( (~ Pdxport_8_8_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Pdxport_8_8_)  &  (~ N_N4242) ) | ( n466  &  (~ N_N4242) ) ;
 assign N_N3052 = ( (~ n278) ) ;
 assign n279 = ( (~ Pdxport_10_10_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Pdxport_10_10_)  &  (~ N_N4194) ) | ( n466  &  (~ N_N4194) ) ;
 assign N_N3051 = ( (~ n279) ) ;
 assign n280 = ( n597  &  n599 ) | ( n597  &  n900 ) | ( n599  &  (~ N_N3540) ) | ( n900  &  (~ N_N3540) ) ;
 assign N_N3050 = ( (~ n280) ) ;
 assign n281 = ( n638  &  n639 ) | ( n638  &  n731 ) | ( n639  &  (~ N_N3679) ) | ( n731  &  (~ N_N3679) ) ;
 assign N_N3049 = ( (~ n281) ) ;
 assign n282 = ( n638  &  n639 ) | ( n638  &  n776 ) | ( n639  &  (~ N_N3701) ) | ( n776  &  (~ N_N3701) ) ;
 assign N_N3048 = ( (~ n282) ) ;
 assign N_N3041 = ( (~ PRESET)  &  (~ NSr5_3) ) ;
 assign n286 = ( n597  &  n599 ) | ( n597  &  n1058 ) | ( n599  &  (~ N_N3750) ) | ( n1058  &  (~ N_N3750) ) ;
 assign N_N3040 = ( (~ n286) ) ;
 assign N_N3038 = ( N_N3468  &  n8 ) ;
 assign n287 = ( PRESET  &  n909 ) | ( n909  &  (~ N_N3346) ) ;
 assign N_N3037 = ( (~ n287) ) ;
 assign n288 = ( n969  &  n1138 ) | ( n1138  &  (~ N_N3822) ) ;
 assign N_N3034 = ( (~ n288) ) ;
 assign n291 = ( n638  &  n639 ) | ( n638  &  n966 ) | ( n639  &  (~ N_N3100) ) | ( n966  &  (~ N_N3100) ) ;
 assign N_N3028 = ( (~ n291) ) ;
 assign n292 = ( n886  &  n887 ) | ( n887  &  n1141 ) | ( n886  &  (~ N_N3974) ) | ( n1141  &  (~ N_N3974) ) ;
 assign N_N3027 = ( (~ n292) ) ;
 assign N_N3016 = ( NDN5_6  &  (~ n944) ) | ( (~ n357)  &  (~ n944) ) ;
 assign n296 = ( n624  &  n625 ) | ( n624  &  n637 ) | ( n625  &  (~ N_N3735) ) | ( n637  &  (~ N_N3735) ) ;
 assign N_N3015 = ( (~ n296) ) ;
 assign n297 = ( n597  &  n599 ) | ( n597  &  n1049 ) | ( n599  &  (~ N_N3821) ) | ( n1049  &  (~ N_N3821) ) ;
 assign N_N3014 = ( (~ n297) ) ;
 assign n299 = ( n464 ) | ( (~ N_N4080) ) ;
 assign N_N3010 = ( (~ n299) ) ;
 assign n300 = ( n464 ) | ( (~ N_N3062) ) ;
 assign N_N3009 = ( (~ n300) ) ;
 assign n301 = ( n597  &  n599 ) | ( n597  &  n899 ) | ( n599  &  (~ N_N3680) ) | ( n899  &  (~ N_N3680) ) ;
 assign N_N3008 = ( (~ n301) ) ;
 assign n302 = ( n597  &  n599 ) | ( n597  &  n1050 ) | ( n599  &  (~ N_N3715) ) | ( n1050  &  (~ N_N3715) ) ;
 assign N_N3007 = ( (~ n302) ) ;
 assign n303 = ( n464 ) | ( (~ N_N3822) ) ;
 assign N_N3004 = ( (~ n303) ) ;
 assign n304 = ( (~ Pdxport_0_0_)  &  n464 ) | ( n464  &  n466 ) | ( (~ Pdxport_0_0_)  &  (~ N_N3906) ) | ( n466  &  (~ N_N3906) ) ;
 assign N_N3003 = ( (~ n304) ) ;
 assign n307 = ( n597  &  n599 ) | ( n597  &  n609 ) | ( n599  &  (~ N_N3677) ) | ( n609  &  (~ N_N3677) ) ;
 assign N_N2998 = ( (~ n307) ) ;
 assign n308 = ( n773  &  n775 ) | ( n773  &  n966 ) | ( n775  &  (~ N_N4133) ) | ( n966  &  (~ N_N4133) ) ;
 assign N_N2997 = ( (~ n308) ) ;
 assign N_N2996 = ( N_N3469  &  n8 ) ;
 assign n310 = ( n597  &  n599 ) | ( n597  &  n892 ) | ( n599  &  (~ N_N3516) ) | ( n892  &  (~ N_N3516) ) ;
 assign N_N2992 = ( (~ n310) ) ;
 assign n312 = ( PRESET  &  n909 ) | ( n909  &  (~ N_N2989) ) ;
 assign N_N2988 = ( (~ n312) ) ;
 assign n313 = ( Pready_0_0_  &  (~ PDN)  &  n1230  &  (~ NLak3_2) ) ;
 assign N_N2987 = ( (~ PRESET)  &  NSr3_2  &  n313 ) ;
 assign n315 = ( n464 ) | ( (~ N_N3262) ) ;
 assign N_N2984 = ( (~ n315) ) ;
 assign n316 = ( n464 ) | ( (~ N_N3280) ) ;
 assign N_N2983 = ( (~ n316) ) ;
 assign n318 = ( n886  &  n887 ) | ( n887  &  n1162 ) | ( n886  &  (~ N_N4027) ) | ( n1162  &  (~ N_N4027) ) ;
 assign N_N2980 = ( (~ n318) ) ;
 assign n319 = ( n464 ) | ( (~ N_N3356) ) ;
 assign N_N2979 = ( (~ n319) ) ;
 assign n320 = ( n464 ) | ( (~ N_N3384) ) ;
 assign N_N2978 = ( (~ n320) ) ;
 assign n321 = ( n624  &  n625 ) | ( n624  &  n726 ) | ( n625  &  (~ N_N3081) ) | ( n726  &  (~ N_N3081) ) ;
 assign N_N2977 = ( (~ n321) ) ;
 assign n322 = ( n727  &  n729 ) | ( n727  &  n776 ) | ( n729  &  (~ N_N3630) ) | ( n776  &  (~ N_N3630) ) ;
 assign N_N2976 = ( (~ n322) ) ;
 assign n323 = ( n637  &  n727 ) | ( n727  &  n729 ) | ( n637  &  (~ N_N3607) ) | ( n729  &  (~ N_N3607) ) ;
 assign N_N2975 = ( (~ n323) ) ;
 assign n324 = ( n464 ) | ( (~ N_N3235) ) ;
 assign N_N2974 = ( (~ n324) ) ;
 assign n325 = ( n597  &  n599 ) | ( n597  &  n889 ) | ( n599  &  (~ N_N3420) ) | ( n889  &  (~ N_N3420) ) ;
 assign N_N2973 = ( (~ n325) ) ;
 assign n326 = ( n727  &  n729 ) | ( n727  &  n781 ) | ( n729  &  (~ N_N3157) ) | ( n781  &  (~ N_N3157) ) ;
 assign N_N2972 = ( (~ n326) ) ;
 assign n328 = ( n464 ) | ( (~ N_N3011) ) ;
 assign N_N2969 = ( (~ n328) ) ;
 assign N_N2966 = ( N_N3312  &  n8 ) ;
 assign N_N2965 = ( N_N3294  &  n8 ) ;
 assign n330 = ( n1172  &  n422 ) | ( n1172  &  n886 ) ;
 assign N_N2964 = ( (~ n330) ) ;
 assign n331 = ( n886  &  n887 ) | ( n887  &  n1173 ) | ( n886  &  (~ N_N4083) ) | ( n1173  &  (~ N_N4083) ) ;
 assign N_N2963 = ( (~ n331) ) ;
 assign n332 = ( n464 ) | ( (~ N_N3541) ) ;
 assign N_N2962 = ( (~ n332) ) ;
 assign n333 = ( n464 ) | ( (~ N_N3866) ) ;
 assign N_N2961 = ( (~ n333) ) ;
 assign N_N2958 = ( N_N4182  &  n8 ) ;
 assign N_N2957 = ( N_N4135  &  n8 ) ;
 assign n335 = ( n969  &  n1178 ) | ( n1178  &  (~ N_N3262) ) ;
 assign N_N2956 = ( (~ n335) ) ;
 assign n336 = ( n969  &  n1179 ) | ( n1179  &  (~ N_N3417) ) ;
 assign N_N2955 = ( (~ n336) ) ;
 assign n337 = ( PRESET  &  n909 ) | ( n909  &  (~ N_N3388) ) ;
 assign N_N2953 = ( (~ n337) ) ;
 assign n338 = ( n969  &  n1180 ) | ( n1180  &  (~ N_N3786) ) ;
 assign N_N2952 = ( (~ n338) ) ;
 assign n339 = ( N_N3811  &  (~ NSr3_2) ) | ( N_N3811  &  n313 ) ;
 assign N_N46 = ( (~ n339) ) ;
 assign n340 = ( (~ n944)  &  (~ NSr5_2) ) | ( (~ n357)  &  NAK5_2  &  (~ n944) ) ;
 assign N_N45 = ( (~ n340) ) ;
 assign n341 = ( (~ n944)  &  (~ NSr5_3) ) | ( NAK5_2  &  (~ n944)  &  (~ NSr5_2) ) ;
 assign N_N44 = ( (~ n341) ) ;
 assign n342 = ( n3  &  (~ N_N3462) ) | ( n3  &  n183 ) ;
 assign N_N43 = ( (~ n342) ) ;
 assign n343 = ( n3  &  (~ N_N3462)  &  (~ n411) ) | ( n3  &  n183  &  (~ n411) ) ;
 assign N_N42 = ( (~ n343) ) ;
 assign n344 = ( (~ NSr5_4)  &  (~ n944) ) | ( NAK5_2  &  (~ n944)  &  (~ NSr5_3) ) ;
 assign N_N41 = ( (~ n344) ) ;
 assign n345 = ( N_N3811  &  (~ NSr3_9) ) | ( NDN3_8  &  n106  &  N_N3811 ) ;
 assign N_N40 = ( (~ n345) ) ;
 assign n346 = ( (~ n944)  &  (~ NSr5_5) ) | ( (~ NSr5_4)  &  NAK5_2  &  (~ n944) ) ;
 assign N_N39 = ( (~ n346) ) ;
 assign n347 = ( (~ n944)  &  (~ NSr5_7) ) | ( NAK5_2  &  (~ n944)  &  (~ NSr5_5) ) ;
 assign N_N38 = ( (~ n347) ) ;
 assign n348 = ( (~ n944)  &  (~ NSr5_8) ) | ( NAK5_2  &  (~ n944)  &  (~ NSr5_7) ) ;
 assign N_N37 = ( (~ n348) ) ;
 assign n349 = ( (~ PRESET)  &  n951  &  (~ n1299) ) | ( (~ PRESET)  &  (~ N_N3998)  &  (~ n1299) ) ;
 assign N_N36 = ( (~ n349) ) ;
 assign n351 = ( (~ n1228)  &  n1230 ) ;
 assign n352 = ( (~ NLD3_9)  &  n460  &  n1228 ) ;
 assign n350 = ( (~ PRESET)  &  n351 ) | ( (~ PRESET)  &  n352 ) ;
 assign n355 = ( n414  &  (~ n882) ) ;
 assign n353 = ( (~ PRESET)  &  n355 ) | ( (~ PRESET)  &  (~ n1271) ) ;
 assign n357 = ( (~ NDN3_8) ) | ( (~ NSr3_9) ) | ( NLak3_9 ) ;
 assign n356 = ( NSr5_4  &  n357 ) | ( n357  &  (~ NSr5_5) ) | ( NSr5_4  &  (~ NSr5_2) ) | ( (~ NSr5_5)  &  (~ NSr5_2) ) ;
 assign n361 = ( n356  &  n372 ) | ( n372  &  (~ N_N3906) ) | ( n356  &  (~ N_N3303) ) | ( (~ N_N3906)  &  (~ N_N3303) ) ;
 assign n362 = ( n385  &  n390 ) | ( n390  &  (~ N_N3939) ) | ( n385  &  (~ N_N3940) ) | ( (~ N_N3939)  &  (~ N_N3940) ) ;
 assign n360 = ( (~ NSr5_7) ) | ( NSr5_5 ) ;
 assign n358 = ( n361  &  n362  &  n360 ) | ( n361  &  n362  &  (~ N_N3304) ) ;
 assign n365 = ( n356  &  n372 ) | ( n372  &  (~ N_N4206) ) | ( n356  &  (~ N_N3188) ) | ( (~ N_N4206)  &  (~ N_N3188) ) ;
 assign n366 = ( n385  &  n390 ) | ( n385  &  (~ N_N3813) ) | ( n390  &  (~ N_N4239) ) | ( (~ N_N3813)  &  (~ N_N4239) ) ;
 assign n363 = ( n360  &  n365  &  n366 ) | ( n365  &  n366  &  (~ N_N3436) ) ;
 assign n369 = ( n356  &  n372 ) | ( n372  &  (~ N_N4165) ) | ( n356  &  (~ N_N3424) ) | ( (~ N_N4165)  &  (~ N_N3424) ) ;
 assign n370 = ( n385  &  n390 ) | ( n385  &  (~ N_N3868) ) | ( n390  &  (~ N_N4099) ) | ( (~ N_N3868)  &  (~ N_N4099) ) ;
 assign n367 = ( n360  &  n369  &  n370 ) | ( n369  &  n370  &  (~ N_N3711) ) ;
 assign n374 = ( n356  &  n360 ) | ( n360  &  (~ N_N4057) ) | ( n356  &  (~ N_N3221) ) | ( (~ N_N4057)  &  (~ N_N3221) ) ;
 assign n375 = ( n385  &  n390 ) | ( n390  &  (~ N_N3918) ) | ( n385  &  (~ N_N3919) ) | ( (~ N_N3918)  &  (~ N_N3919) ) ;
 assign n372 = ( NSr5_7 ) | ( (~ NSr5_8) ) ;
 assign n371 = ( n374  &  n375  &  n372 ) | ( n374  &  n375  &  (~ N_N3367) ) ;
 assign n378 = ( n356  &  n372 ) | ( n372  &  (~ N_N4120) ) | ( n356  &  (~ N_N4116) ) | ( (~ N_N4120)  &  (~ N_N4116) ) ;
 assign n379 = ( n385  &  n390 ) | ( n390  &  (~ N_N4118) ) | ( n385  &  (~ N_N4119) ) | ( (~ N_N4118)  &  (~ N_N4119) ) ;
 assign n376 = ( n360  &  n378  &  n379 ) | ( n378  &  n379  &  (~ N_N4117) ) ;
 assign n382 = ( n356  &  n372 ) | ( n372  &  (~ N_N4220) ) | ( n356  &  (~ N_N3921) ) | ( (~ N_N4220)  &  (~ N_N3921) ) ;
 assign n383 = ( n385  &  n390 ) | ( n390  &  (~ N_N3923) ) | ( n385  &  (~ N_N3924) ) | ( (~ N_N3923)  &  (~ N_N3924) ) ;
 assign n380 = ( n360  &  n382  &  n383 ) | ( n382  &  n383  &  (~ N_N3922) ) ;
 assign n387 = ( n356  &  n372 ) | ( n372  &  (~ N_N4179) ) | ( n356  &  (~ N_N3870) ) | ( (~ N_N4179)  &  (~ N_N3870) ) ;
 assign n388 = ( n360  &  n390 ) | ( n360  &  (~ N_N3872) ) | ( n390  &  (~ N_N4030) ) | ( (~ N_N3872)  &  (~ N_N4030) ) ;
 assign n385 = ( (~ NSr5_4) ) | ( NSr5_3 ) ;
 assign n384 = ( n387  &  n388  &  n385 ) | ( n387  &  n388  &  (~ N_N3871) ) ;
 assign n392 = ( n356  &  n360 ) | ( n360  &  (~ N_N4242) ) | ( n356  &  (~ N_N3164) ) | ( (~ N_N4242)  &  (~ N_N3164) ) ;
 assign n393 = ( n372  &  n385 ) | ( n385  &  (~ N_N4047) ) | ( n372  &  (~ N_N4252) ) | ( (~ N_N4047)  &  (~ N_N4252) ) ;
 assign n390 = ( (~ NSr5_3) ) | ( NSr5_2 ) ;
 assign n389 = ( n392  &  n393  &  n390 ) | ( n392  &  n393  &  (~ N_N3800) ) ;
 assign n396 = ( n356  &  n372 ) | ( n372  &  (~ N_N4070) ) | ( n356  &  (~ N_N3805) ) | ( (~ N_N4070)  &  (~ N_N3805) ) ;
 assign n397 = ( n385  &  n390 ) | ( n390  &  (~ N_N3807) ) | ( n385  &  (~ N_N3808) ) | ( (~ N_N3807)  &  (~ N_N3808) ) ;
 assign n394 = ( n360  &  n396  &  n397 ) | ( n396  &  n397  &  (~ N_N3806) ) ;
 assign n400 = ( n356  &  n372 ) | ( n372  &  (~ N_N4132) ) | ( n356  &  (~ N_N3840) ) | ( (~ N_N4132)  &  (~ N_N3840) ) ;
 assign n401 = ( n385  &  n390 ) | ( n390  &  (~ N_N3842) ) | ( n385  &  (~ N_N3843) ) | ( (~ N_N3842)  &  (~ N_N3843) ) ;
 assign n398 = ( n360  &  n400  &  n401 ) | ( n400  &  n401  &  (~ N_N3841) ) ;
 assign n404 = ( n356  &  n360 ) | ( n360  &  (~ N_N4237) ) | ( n356  &  (~ N_N3433) ) | ( (~ N_N4237)  &  (~ N_N3433) ) ;
 assign n405 = ( n385  &  n390 ) | ( n390  &  (~ N_N4208) ) | ( n385  &  (~ N_N4209) ) | ( (~ N_N4208)  &  (~ N_N4209) ) ;
 assign n402 = ( n372  &  n404  &  n405 ) | ( n404  &  n405  &  (~ N_N3659) ) ;
 assign n408 = ( n356  &  n360 ) | ( n360  &  (~ N_N4194) ) | ( n356  &  (~ N_N3457) ) | ( (~ N_N4194)  &  (~ N_N3457) ) ;
 assign n409 = ( n385  &  n390 ) | ( n390  &  (~ N_N4176) ) | ( n385  &  (~ N_N4177) ) | ( (~ N_N4176)  &  (~ N_N4177) ) ;
 assign n406 = ( n372  &  n408  &  n409 ) | ( n408  &  n409  &  (~ N_N4045) ) ;
 assign n411 = ( n390  &  n385  &  n360  &  n372  &  n356 ) ;
 assign n412 = ( (~ N_N3999)  &  (~ n1297) ) | ( N_N3838  &  (~ n1297) ) ;
 assign n410 = ( N_N3460  &  n411 ) | ( N_N3460  &  n412 ) ;
 assign n414 = ( N_N3578 ) | ( n410 ) ;
 assign n413 = ( n412  &  (~ n1221) ) | ( n414  &  (~ n1221) ) ;
 assign n417 = ( (~ n353)  &  (~ N_N4060) ) | ( (~ n353)  &  n886 ) | ( N_N4060  &  n886 ) ;
 assign n416 = ( PRESET ) | ( n413 ) ;
 assign N_N47 = ( n417  &  n358 ) | ( n417  &  n416 ) ;
 assign n421 = ( N_N3369 ) | ( n436 ) ;
 assign n418 = ( n421  &  (~ n436) ) | ( n421  &  (~ N_N3369) ) ;
 assign n424 = ( (~ N_N4060) ) | ( N_N3961 ) ;
 assign n422 = ( n424  &  N_N4060 ) | ( n424  &  (~ N_N3961) ) ;
 assign n428 = ( N_N4093 ) | ( n432 ) ;
 assign n425 = ( n428  &  (~ n432) ) | ( n428  &  (~ N_N4093) ) ;
 assign n432 = ( N_N4212 ) | ( n448 ) ;
 assign n429 = ( n432  &  (~ n448) ) | ( n432  &  (~ N_N4212) ) ;
 assign n436 = ( N_N4246 ) | ( n428 ) ;
 assign n433 = ( (~ n428)  &  n436 ) | ( n436  &  (~ N_N4246) ) ;
 assign n440 = ( N_N4171 ) | ( n452 ) ;
 assign n437 = ( n440  &  (~ n452) ) | ( n440  &  (~ N_N4171) ) ;
 assign n444 = ( N_N4126 ) | ( n424 ) ;
 assign n441 = ( (~ n424)  &  n444 ) | ( n444  &  (~ N_N4126) ) ;
 assign n448 = ( N_N4036 ) | ( n440 ) ;
 assign n445 = ( (~ n440)  &  n448 ) | ( n448  &  (~ N_N4036) ) ;
 assign n452 = ( N_N4004 ) | ( n444 ) ;
 assign n449 = ( (~ n444)  &  n452 ) | ( n452  &  (~ N_N4004) ) ;
 assign n461 = ( (~ NLD3_9)  &  (~ n351) ) | ( (~ NLD3_9)  &  (~ N_N4239) ) | ( (~ n351)  &  (~ N_N3774) ) | ( (~ N_N4239)  &  (~ N_N3774) ) ;
 assign n460 = ( NDN3_8 ) | ( (~ NDN3_3) ) ;
 assign n458 = ( n461  &  n460 ) | ( n461  &  (~ N_N4090) ) ;
 assign n463 = ( PRESET ) | ( (~ n352) ) ;
 assign n464 = ( n1233 ) | ( PRESET ) ;
 assign n466 = ( PRESET ) | ( (~ n1233) ) ;
 assign n475 = ( NDN5_9 ) | ( (~ NEN5_9) ) ;
 assign n476 = ( NDN5_10 ) | ( NSr5_7 ) ;
 assign n473 = ( n475  &  n476 ) | ( n476  &  (~ N_N3612) ) | ( n475  &  (~ N_N4039) ) | ( (~ N_N3612)  &  (~ N_N4039) ) ;
 assign n478 = ( n475  &  n476 ) | ( n475  &  (~ N_N3482) ) | ( n476  &  (~ N_N4075) ) | ( (~ N_N3482)  &  (~ N_N4075) ) ;
 assign n481 = ( n475  &  n476 ) | ( n476  &  (~ N_N3735) ) | ( n475  &  (~ N_N3736) ) | ( (~ N_N3735)  &  (~ N_N3736) ) ;
 assign n484 = ( n475  &  n476 ) | ( n476  &  (~ N_N3700) ) | ( n475  &  (~ N_N3701) ) | ( (~ N_N3700)  &  (~ N_N3701) ) ;
 assign n487 = ( n475  &  n476 ) | ( n475  &  (~ N_N3679) ) | ( n476  &  (~ N_N4021) ) | ( (~ N_N3679)  &  (~ N_N4021) ) ;
 assign n490 = ( n475  &  n476 ) | ( n476  &  (~ N_N3625) ) | ( n475  &  (~ N_N3626) ) | ( (~ N_N3625)  &  (~ N_N3626) ) ;
 assign n493 = ( n475  &  n476 ) | ( n475  &  (~ N_N3799) ) | ( n476  &  (~ N_N4024) ) | ( (~ N_N3799)  &  (~ N_N4024) ) ;
 assign n496 = ( n475  &  n476 ) | ( n476  &  (~ N_N3959) ) | ( n475  &  (~ N_N3968) ) | ( (~ N_N3959)  &  (~ N_N3968) ) ;
 assign n499 = ( n475  &  n476 ) | ( n475  &  (~ N_N3205) ) | ( n476  &  (~ N_N3957) ) | ( (~ N_N3205)  &  (~ N_N3957) ) ;
 assign n502 = ( n475  &  n476 ) | ( n476  &  (~ N_N3081) ) | ( n475  &  (~ N_N3203) ) | ( (~ N_N3081)  &  (~ N_N3203) ) ;
 assign n505 = ( n475  &  n476 ) | ( n475  &  (~ N_N3100) ) | ( n476  &  (~ N_N3585) ) | ( (~ N_N3100)  &  (~ N_N3585) ) ;
 assign n508 = ( n475  &  n476 ) | ( n476  &  (~ N_N3824) ) | ( n475  &  (~ N_N4042) ) | ( (~ N_N3824)  &  (~ N_N4042) ) ;
 assign n511 = ( n475  &  n476 ) | ( n476  &  (~ N_N3274) ) | ( n475  &  (~ N_N3470) ) | ( (~ N_N3274)  &  (~ N_N3470) ) ;
 assign n514 = ( n475  &  n476 ) | ( n475  &  (~ N_N3810) ) | ( n476  &  (~ N_N3947) ) | ( (~ N_N3810)  &  (~ N_N3947) ) ;
 assign n518 = ( n502  &  n484  &  n564 ) ;
 assign n517 = ( n518  &  n505 ) ;
 assign n519 = ( n475  &  n476 ) | ( n476  &  (~ N_N3829) ) | ( n475  &  (~ N_N4224) ) | ( (~ N_N3829)  &  (~ N_N4224) ) ;
 assign n522 = ( n475  &  n476 ) | ( n476  &  (~ N_N3796) ) | ( n475  &  (~ N_N3971) ) | ( (~ N_N3796)  &  (~ N_N3971) ) ;
 assign n525 = ( n475  &  n476 ) | ( n475  &  (~ N_N3500) ) | ( n476  &  (~ N_N3684) ) | ( (~ N_N3500)  &  (~ N_N3684) ) ;
 assign n528 = ( (~ n490)  &  (~ n522)  &  (~ n525) ) | ( (~ n490)  &  (~ n522)  &  (~ n534) ) ;
 assign n534 = ( n490  &  n496 ) | ( (~ n490)  &  (~ n496) ) ;
 assign n533 = ( n525  &  (~ n528) ) | ( (~ n528)  &  n534 ) ;
 assign n536 = ( n490  &  n496 ) ;
 assign n537 = ( n475  &  n476 ) | ( n476  &  (~ N_N3480) ) | ( n475  &  (~ N_N4086) ) | ( (~ N_N3480)  &  (~ N_N4086) ) ;
 assign n540 = ( n537  &  (~ n1184) ) ;
 assign n542 = ( n533  &  n537 ) | ( n537  &  n540 ) | ( n533  &  (~ n1184) ) | ( n540  &  (~ n1184) ) ;
 assign n543 = ( n519  &  n542 ) ;
 assign n544 = ( n519  &  n543 ) | ( n542  &  n543 ) | ( n519  &  (~ n1185) ) | ( n542  &  (~ n1185) ) ;
 assign n546 = ( n475  &  n476 ) | ( n476  &  (~ N_N3509) ) | ( n475  &  (~ N_N3890) ) | ( (~ N_N3509)  &  (~ N_N3890) ) ;
 assign n550 = ( n496  &  n493  &  n490 ) ;
 assign n549 = ( n550  &  n499 ) ;
 assign n551 = ( n546  &  (~ n1186) ) ;
 assign n553 = ( n544  &  n546 ) | ( n546  &  n551 ) | ( n544  &  (~ n1186) ) | ( n551  &  (~ n1186) ) ;
 assign n554 = ( n475  &  n476 ) | ( n476  &  (~ N_N3826) ) | ( n475  &  (~ N_N4183) ) | ( (~ N_N3826)  &  (~ N_N4183) ) ;
 assign n557 = ( n554  &  (~ n1187) ) ;
 assign n559 = ( n553  &  n554 ) | ( n554  &  n557 ) | ( n553  &  (~ n1187) ) | ( n557  &  (~ n1187) ) ;
 assign n560 = ( n475  &  n476 ) | ( n476  &  (~ N_N3529) ) | ( n475  &  (~ N_N3844) ) | ( (~ N_N3529)  &  (~ N_N3844) ) ;
 assign n564 = ( n499  &  n487  &  n550 ) ;
 assign n563 = ( n564  &  n502 ) ;
 assign n565 = ( n560  &  (~ n1188) ) ;
 assign n567 = ( n559  &  n560 ) | ( n560  &  n565 ) | ( n559  &  (~ n1188) ) | ( n565  &  (~ n1188) ) ;
 assign n568 = ( n475  &  n476 ) | ( n476  &  (~ N_N3815) ) | ( n475  &  (~ N_N4136) ) | ( (~ N_N3815)  &  (~ N_N4136) ) ;
 assign n571 = ( n568  &  (~ n1189) ) ;
 assign n573 = ( n567  &  n568 ) | ( n568  &  n571 ) | ( n567  &  (~ n1189) ) | ( n571  &  (~ n1189) ) ;
 assign n575 = ( n481  &  n517 ) | ( (~ n481)  &  (~ n517) ) ;
 assign n574 = ( n573  &  n575 ) ;
 assign n576 = ( n514  &  n573 ) | ( n574  &  n573 ) | ( n514  &  n575 ) | ( n574  &  n575 ) ;
 assign n577 = ( n475  &  n476 ) | ( n476  &  (~ N_N3788) ) | ( n475  &  (~ N_N4140) ) | ( (~ N_N3788)  &  (~ N_N4140) ) ;
 assign n580 = ( n576  &  n577 ) ;
 assign n581 = ( n576  &  n580 ) | ( n577  &  n580 ) | ( n576  &  (~ n1191) ) | ( n577  &  (~ n1191) ) ;
 assign n583 = ( n511  &  n581 ) ;
 assign n585 = ( n478  &  n1238 ) | ( (~ n478)  &  (~ n1238) ) ;
 assign n584 = ( n583  &  n511 ) | ( n585  &  n511 ) | ( n583  &  n581 ) | ( n585  &  n581 ) ;
 assign n586 = ( n475  &  n476 ) | ( n476  &  (~ N_N4167) ) | ( n475  &  (~ N_N4095) ) | ( (~ N_N4167)  &  (~ N_N4095) ) ;
 assign n591 = ( PRESET ) | ( n476 ) ;
 assign n596 = ( (~ NLD3_9)  &  (~ n351) ) | ( (~ NLD3_9)  &  (~ N_N4140) ) | ( (~ n351)  &  (~ N_N3540) ) | ( (~ N_N4140)  &  (~ N_N3540) ) ;
 assign n594 = ( n460  &  n596 ) | ( n596  &  (~ N_N3541) ) ;
 assign n597 = ( PRESET ) | ( (~ n475) ) ;
 assign n599 = ( PRESET ) | ( n475 ) ;
 assign n602 = ( NDN5_6 ) | ( n357 ) ;
 assign n600 = ( n475  &  n602 ) | ( n475  &  (~ N_N3906) ) | ( n602  &  (~ N_N3910) ) | ( (~ N_N3906)  &  (~ N_N3910) ) ;
 assign n604 = ( n475  &  n602 ) | ( n602  &  (~ N_N3939) ) | ( n475  &  (~ N_N3940) ) | ( (~ N_N3939)  &  (~ N_N3940) ) ;
 assign n607 = ( PRESET ) | ( (~ n602) ) ;
 assign n609 = ( n600  &  n604 ) | ( (~ n600)  &  (~ n604) ) ;
 assign n610 = ( PRESET ) | ( n602 ) ;
 assign n616 = ( (~ n351)  &  n460 ) | ( n460  &  (~ N_N4099) ) | ( (~ n351)  &  (~ N_N3384) ) | ( (~ N_N4099)  &  (~ N_N3384) ) ;
 assign n613 = ( (~ NLD3_9)  &  n616 ) | ( n616  &  (~ N_N3743) ) ;
 assign n619 = ( (~ n351)  &  n460 ) | ( n460  &  (~ N_N4095) ) | ( (~ n351)  &  (~ N_N3866) ) | ( (~ N_N4095)  &  (~ N_N3866) ) ;
 assign n618 = ( (~ NLD3_9)  &  n619 ) | ( n619  &  (~ N_N4114) ) ;
 assign n623 = ( (~ NLD3_9)  &  (~ n351) ) | ( (~ NLD3_9)  &  (~ N_N4086) ) | ( (~ n351)  &  (~ N_N3715) ) | ( (~ N_N4086)  &  (~ N_N3715) ) ;
 assign n621 = ( n460  &  n623 ) | ( n623  &  (~ N_N3716) ) ;
 assign n624 = ( PRESET ) | ( (~ n1242) ) ;
 assign n625 = ( PRESET ) | ( n1242 ) ;
 assign n626 = ( (~ n412) ) | ( (~ N_N4197) ) ;
 assign n635 = ( PRESET ) | ( (~ n1245) ) ;
 assign n636 = ( PRESET ) | ( n1245 ) ;
 assign n637 = ( (~ n412) ) | ( (~ N_N4145) ) ;
 assign n638 = ( PRESET ) | ( (~ n1247) ) ;
 assign n639 = ( PRESET ) | ( n1247 ) ;
 assign n640 = ( (~ n412) ) | ( (~ N_N3912) ) ;
 assign n641 = ( (~ n412) ) | ( (~ N_N4227) ) ;
 assign n642 = ( n475  &  n602 ) | ( n475  &  (~ N_N4194) ) | ( n602  &  (~ N_N4193) ) | ( (~ N_N4194)  &  (~ N_N4193) ) ;
 assign n645 = ( n475  &  n602 ) | ( n602  &  (~ N_N4176) ) | ( n475  &  (~ N_N4177) ) | ( (~ N_N4176)  &  (~ N_N4177) ) ;
 assign n648 = ( n475  &  n602 ) | ( n475  &  (~ N_N3800) ) | ( n602  &  (~ N_N4252) ) | ( (~ N_N3800)  &  (~ N_N4252) ) ;
 assign n650 = ( n475  &  n602 ) | ( n475  &  (~ N_N4242) ) | ( n602  &  (~ N_N3607) ) | ( (~ N_N4242)  &  (~ N_N3607) ) ;
 assign n653 = ( n475  &  n602 ) | ( n475  &  (~ N_N4220) ) | ( n602  &  (~ N_N3143) ) | ( (~ N_N4220)  &  (~ N_N3143) ) ;
 assign n656 = ( n475  &  n602 ) | ( n602  &  (~ N_N3923) ) | ( n475  &  (~ N_N3924) ) | ( (~ N_N3923)  &  (~ N_N3924) ) ;
 assign n659 = ( n475  &  n602 ) | ( n602  &  (~ N_N3918) ) | ( n475  &  (~ N_N3919) ) | ( (~ N_N3918)  &  (~ N_N3919) ) ;
 assign n662 = ( n475  &  n602 ) | ( n475  &  (~ N_N4057) ) | ( n602  &  (~ N_N3793) ) | ( (~ N_N4057)  &  (~ N_N3793) ) ;
 assign n665 = ( n475  &  n602 ) | ( n602  &  (~ N_N4118) ) | ( n475  &  (~ N_N4119) ) | ( (~ N_N4118)  &  (~ N_N4119) ) ;
 assign n668 = ( n475  &  n602 ) | ( n475  &  (~ N_N4120) ) | ( n602  &  (~ N_N3157) ) | ( (~ N_N4120)  &  (~ N_N3157) ) ;
 assign n671 = ( (~ n600)  &  (~ n604)  &  (~ n665) ) | ( (~ n600)  &  (~ n604)  &  (~ n668) ) ;
 assign n676 = ( n665  &  (~ n671) ) | ( n668  &  (~ n671) ) ;
 assign n678 = ( n662  &  n676 ) ;
 assign n679 = ( n659  &  n662 ) | ( n678  &  n662 ) | ( n659  &  n676 ) | ( n678  &  n676 ) ;
 assign n680 = ( n656  &  n679 ) ;
 assign n681 = ( n653  &  n656 ) | ( n680  &  n656 ) | ( n653  &  n679 ) | ( n680  &  n679 ) ;
 assign n682 = ( n475  &  n602 ) | ( n475  &  (~ N_N3868) ) | ( n602  &  (~ N_N4099) ) | ( (~ N_N3868)  &  (~ N_N4099) ) ;
 assign n684 = ( n475  &  n602 ) | ( n475  &  (~ N_N4165) ) | ( n602  &  (~ N_N3776) ) | ( (~ N_N4165)  &  (~ N_N3776) ) ;
 assign n687 = ( n682  &  n684 ) ;
 assign n688 = ( n681  &  n682 ) | ( n687  &  n682 ) | ( n681  &  n684 ) | ( n687  &  n684 ) ;
 assign n689 = ( n475  &  n602 ) | ( n602  &  (~ N_N3871) ) | ( n475  &  (~ N_N3872) ) | ( (~ N_N3871)  &  (~ N_N3872) ) ;
 assign n691 = ( n475  &  n602 ) | ( n475  &  (~ N_N4179) ) | ( n602  &  (~ N_N3071) ) | ( (~ N_N4179)  &  (~ N_N3071) ) ;
 assign n694 = ( n689  &  n691 ) ;
 assign n695 = ( n688  &  n689 ) | ( n694  &  n689 ) | ( n688  &  n691 ) | ( n694  &  n691 ) ;
 assign n696 = ( n475  &  n602 ) | ( n475  &  (~ N_N3813) ) | ( n602  &  (~ N_N4239) ) | ( (~ N_N3813)  &  (~ N_N4239) ) ;
 assign n698 = ( n475  &  n602 ) | ( n475  &  (~ N_N4206) ) | ( n602  &  (~ N_N3630) ) | ( (~ N_N4206)  &  (~ N_N3630) ) ;
 assign n701 = ( n696  &  n698 ) ;
 assign n702 = ( n695  &  n696 ) | ( n701  &  n696 ) | ( n695  &  n698 ) | ( n701  &  n698 ) ;
 assign n703 = ( n475  &  n602 ) | ( n602  &  (~ N_N3842) ) | ( n475  &  (~ N_N3843) ) | ( (~ N_N3842)  &  (~ N_N3843) ) ;
 assign n706 = ( n475  &  n602 ) | ( n475  &  (~ N_N4132) ) | ( n602  &  (~ N_N3069) ) | ( (~ N_N4132)  &  (~ N_N3069) ) ;
 assign n709 = ( n703  &  n706 ) ;
 assign n710 = ( n702  &  n703 ) | ( n709  &  n703 ) | ( n702  &  n706 ) | ( n709  &  n706 ) ;
 assign n711 = ( n650  &  n710 ) ;
 assign n712 = ( n648  &  n650 ) | ( n711  &  n650 ) | ( n648  &  n710 ) | ( n711  &  n710 ) ;
 assign n713 = ( n475  &  n602 ) | ( n602  &  (~ N_N3807) ) | ( n475  &  (~ N_N3808) ) | ( (~ N_N3807)  &  (~ N_N3808) ) ;
 assign n716 = ( n475  &  n602 ) | ( n475  &  (~ N_N4070) ) | ( n602  &  (~ N_N3311) ) | ( (~ N_N4070)  &  (~ N_N3311) ) ;
 assign n719 = ( n713  &  n716 ) ;
 assign n720 = ( n712  &  n713 ) | ( n719  &  n713 ) | ( n712  &  n716 ) | ( n719  &  n716 ) ;
 assign n722 = ( (~ n720)  &  n1286 ) | ( n720  &  (~ n1286) ) ;
 assign n724 = ( PRESET ) | ( (~ n1250) ) ;
 assign n725 = ( PRESET ) | ( n1250 ) ;
 assign n726 = ( (~ n412) ) | ( (~ N_N3974) ) ;
 assign n727 = ( PRESET ) | ( (~ n1252) ) ;
 assign n729 = ( PRESET ) | ( n1252 ) ;
 assign n730 = ( (~ n412) ) | ( (~ N_N3992) ) ;
 assign n731 = ( (~ n412) ) | ( (~ N_N4018) ) ;
 assign n735 = ( N_N3916  &  N_N3797  &  (~ N_N4111) ) | ( N_N3916  &  (~ N_N3535)  &  (~ N_N4111) ) ;
 assign n736 = ( (~ N_N3797)  &  (~ n735) ) | ( (~ n735)  &  N_N3535 ) ;
 assign n739 = ( n736  &  (~ N_N3733) ) ;
 assign n741 = ( n736  &  n739 ) | ( n736  &  N_N3794 ) | ( n739  &  (~ N_N3733) ) | ( N_N3794  &  (~ N_N3733) ) ;
 assign n742 = ( n741  &  (~ N_N3778) ) ;
 assign n744 = ( n741  &  n742 ) | ( n741  &  N_N3981 ) | ( n742  &  (~ N_N3778) ) | ( N_N3981  &  (~ N_N3778) ) ;
 assign n746 = ( (~ n744)  &  N_N3574 ) ;
 assign n748 = ( (~ n744)  &  n746 ) | ( N_N3574  &  n746 ) | ( (~ n744)  &  (~ N_N3832) ) | ( N_N3574  &  (~ N_N3832) ) ;
 assign n750 = ( n748  &  (~ N_N3761) ) ;
 assign n752 = ( n748  &  n750 ) | ( n748  &  N_N4056 ) | ( n750  &  (~ N_N3761) ) | ( N_N4056  &  (~ N_N3761) ) ;
 assign n754 = ( (~ n752)  &  N_N3862 ) ;
 assign n756 = ( (~ n752)  &  n754 ) | ( N_N3862  &  n754 ) | ( (~ n752)  &  (~ N_N4243) ) | ( N_N3862  &  (~ N_N4243) ) ;
 assign n759 = ( n756  &  N_N3489 ) ;
 assign n760 = ( n756  &  n759 ) | ( N_N3489  &  n759 ) | ( n756  &  (~ N_N4054) ) | ( N_N3489  &  (~ N_N4054) ) ;
 assign n761 = ( (~ n760)  &  (~ N_N3908) ) ;
 assign n764 = ( (~ n760)  &  n761 ) | ( (~ n760)  &  N_N4015 ) | ( n761  &  (~ N_N3908) ) | ( N_N4015  &  (~ N_N3908) ) ;
 assign n765 = ( n764  &  (~ N_N3513) ) ;
 assign n767 = ( n764  &  n765 ) | ( n764  &  N_N3818 ) | ( n765  &  (~ N_N3513) ) | ( N_N3818  &  (~ N_N3513) ) ;
 assign n769 = ( (~ n767)  &  N_N3884 ) | ( (~ N_N3882)  &  N_N3884 ) ;
 assign n771 = ( (~ n767)  &  (~ N_N3882) ) ;
 assign n773 = ( PRESET ) | ( (~ n1254) ) ;
 assign n775 = ( PRESET ) | ( n1254 ) ;
 assign n776 = ( (~ n412) ) | ( (~ N_N4083) ) ;
 assign n778 = ( (~ n679)  &  n1287 ) | ( n679  &  (~ n1287) ) ;
 assign n781 = ( (~ n412) ) | ( (~ N_N4027) ) ;
 assign n783 = ( (~ n412) ) | ( (~ N_N3996) ) ;
 assign n784 = ( (~ n575)  &  n1197 ) | ( n575  &  (~ n1197) ) ;
 assign n793 = ( (~ n412) ) | ( (~ N_N3965) ) ;
 assign n802 = ( (~ N_N3445)  &  n356 ) | ( n356  &  n385 ) | ( (~ N_N3445)  &  (~ N_N4095) ) | ( n385  &  (~ N_N4095) ) ;
 assign n803 = ( (~ N_N3905)  &  n372 ) | ( n372  &  n390 ) | ( (~ N_N3905)  &  (~ N_N4237) ) | ( n390  &  (~ N_N4237) ) ;
 assign n800 = ( n360  &  n802  &  n803 ) | ( n802  &  n803  &  (~ N_N3663) ) ;
 assign n806 = ( (~ N_N3468)  &  n356 ) | ( n356  &  n385 ) | ( (~ N_N3468)  &  (~ N_N3470) ) | ( n385  &  (~ N_N3470) ) ;
 assign n807 = ( n360  &  n372 ) | ( n360  &  (~ N_N4194) ) | ( n372  &  (~ N_N3473) ) | ( (~ N_N4194)  &  (~ N_N3473) ) ;
 assign n804 = ( (~ N_N3469)  &  n806  &  n807 ) | ( n390  &  n806  &  n807 ) ;
 assign n810 = ( n356  &  n372 ) | ( n356  &  (~ N_N4070) ) | ( n372  &  (~ N_N4140) ) | ( (~ N_N4070)  &  (~ N_N4140) ) ;
 assign n811 = ( (~ N_N4073)  &  (~ N_N4072) ) | ( (~ N_N4073)  &  n385 ) | ( (~ N_N4072)  &  n390 ) | ( n385  &  n390 ) ;
 assign n808 = ( n360  &  n810  &  n811 ) | ( n810  &  n811  &  (~ N_N4071) ) ;
 assign n814 = ( n356  &  n360 ) | ( n360  &  (~ N_N3810) ) | ( n356  &  (~ N_N3293) ) | ( (~ N_N3810)  &  (~ N_N3293) ) ;
 assign n815 = ( (~ N_N3426)  &  n372 ) | ( n372  &  n385 ) | ( (~ N_N3426)  &  (~ N_N4242) ) | ( n385  &  (~ N_N4242) ) ;
 assign n812 = ( (~ N_N3294)  &  n814  &  n815 ) | ( n390  &  n814  &  n815 ) ;
 assign n818 = ( n356  &  n372 ) | ( n356  &  (~ N_N4132) ) | ( n372  &  (~ N_N4136) ) | ( (~ N_N4132)  &  (~ N_N4136) ) ;
 assign n819 = ( (~ N_N4134)  &  (~ N_N4135) ) | ( (~ N_N4135)  &  n385 ) | ( (~ N_N4134)  &  n390 ) | ( n385  &  n390 ) ;
 assign n816 = ( n360  &  n818  &  n819 ) | ( n818  &  n819  &  (~ N_N4133) ) ;
 assign n822 = ( (~ N_N3312)  &  n356 ) | ( n356  &  n390 ) | ( (~ N_N3312)  &  (~ N_N3844) ) | ( n390  &  (~ N_N3844) ) ;
 assign n823 = ( n360  &  n372 ) | ( n360  &  (~ N_N4206) ) | ( n372  &  (~ N_N3988) ) | ( (~ N_N4206)  &  (~ N_N3988) ) ;
 assign n820 = ( (~ N_N3375)  &  n822  &  n823 ) | ( n385  &  n822  &  n823 ) ;
 assign n826 = ( n356  &  n372 ) | ( n356  &  (~ N_N4179) ) | ( n372  &  (~ N_N4183) ) | ( (~ N_N4179)  &  (~ N_N4183) ) ;
 assign n827 = ( (~ N_N4181)  &  (~ N_N4182) ) | ( (~ N_N4182)  &  n385 ) | ( (~ N_N4181)  &  n390 ) | ( n385  &  n390 ) ;
 assign n824 = ( n360  &  n826  &  n827 ) | ( n826  &  n827  &  (~ N_N4180) ) ;
 assign n830 = ( n356  &  n360 ) | ( n360  &  (~ N_N3890) ) | ( n356  &  (~ N_N3323) ) | ( (~ N_N3890)  &  (~ N_N3323) ) ;
 assign n831 = ( (~ N_N3691)  &  n372 ) | ( n372  &  n385 ) | ( (~ N_N3691)  &  (~ N_N4165) ) | ( n385  &  (~ N_N4165) ) ;
 assign n828 = ( (~ N_N3324)  &  n830  &  n831 ) | ( n390  &  n830  &  n831 ) ;
 assign n834 = ( n356  &  n372 ) | ( n356  &  (~ N_N4220) ) | ( n372  &  (~ N_N4224) ) | ( (~ N_N4220)  &  (~ N_N4224) ) ;
 assign n835 = ( (~ N_N4222)  &  (~ N_N4223) ) | ( (~ N_N4223)  &  n385 ) | ( (~ N_N4222)  &  n390 ) | ( n385  &  n390 ) ;
 assign n832 = ( n360  &  n834  &  n835 ) | ( n834  &  n835  &  (~ N_N4221) ) ;
 assign n838 = ( n356  &  n360 ) | ( n360  &  (~ N_N4086) ) | ( n356  &  (~ N_N3344) ) | ( (~ N_N4086)  &  (~ N_N3344) ) ;
 assign n839 = ( n372  &  n390 ) | ( n390  &  (~ N_N4057) ) | ( n372  &  (~ N_N3346) ) | ( (~ N_N4057)  &  (~ N_N3346) ) ;
 assign n836 = ( (~ N_N3345)  &  n838  &  n839 ) | ( n385  &  n838  &  n839 ) ;
 assign n842 = ( n356  &  n385 ) | ( n385  &  (~ N_N3500) ) | ( n356  &  (~ N_N2989) ) | ( (~ N_N3500)  &  (~ N_N2989) ) ;
 assign n843 = ( (~ N_N3708)  &  n372 ) | ( n372  &  n390 ) | ( (~ N_N3708)  &  (~ N_N4120) ) | ( n390  &  (~ N_N4120) ) ;
 assign n840 = ( n360  &  n842  &  n843 ) | ( n842  &  n843  &  (~ N_N3175) ) ;
 assign n846 = ( n356  &  n360 ) | ( n360  &  (~ N_N3971) ) | ( n356  &  (~ N_N3387) ) | ( (~ N_N3971)  &  (~ N_N3387) ) ;
 assign n847 = ( n372  &  n385 ) | ( n385  &  (~ N_N3906) ) | ( n372  &  (~ N_N3745) ) | ( (~ N_N3906)  &  (~ N_N3745) ) ;
 assign n844 = ( n390  &  n846  &  n847 ) | ( n846  &  n847  &  (~ N_N3388) ) ;
 assign n849 = ( n844 ) | ( (~ N_N3965) ) ;
 assign n848 = ( n840  &  n849 ) ;
 assign n850 = ( n840  &  n848 ) | ( n849  &  n848 ) | ( n840  &  (~ N_N4027) ) | ( n849  &  (~ N_N4027) ) ;
 assign n852 = ( n850  &  (~ N_N3992) ) ;
 assign n854 = ( n836  &  n850 ) | ( n850  &  n852 ) | ( n836  &  (~ N_N3992) ) | ( n852  &  (~ N_N3992) ) ;
 assign n855 = ( n854  &  (~ N_N3996) ) ;
 assign n857 = ( n832  &  n854 ) | ( n854  &  n855 ) | ( n832  &  (~ N_N3996) ) | ( n855  &  (~ N_N3996) ) ;
 assign n858 = ( n857  &  (~ N_N4018) ) ;
 assign n860 = ( n828  &  n857 ) | ( n857  &  n858 ) | ( n828  &  (~ N_N4018) ) | ( n858  &  (~ N_N4018) ) ;
 assign n861 = ( n860  &  (~ N_N3974) ) ;
 assign n863 = ( n824  &  n860 ) | ( n860  &  n861 ) | ( n824  &  (~ N_N3974) ) | ( n861  &  (~ N_N3974) ) ;
 assign n864 = ( n863  &  (~ N_N4083) ) ;
 assign n866 = ( n820  &  n863 ) | ( n863  &  n864 ) | ( n820  &  (~ N_N4083) ) | ( n864  &  (~ N_N4083) ) ;
 assign n867 = ( n866  &  (~ N_N3949) ) ;
 assign n869 = ( n816  &  n866 ) | ( n866  &  n867 ) | ( n816  &  (~ N_N3949) ) | ( n867  &  (~ N_N3949) ) ;
 assign n870 = ( n869  &  (~ N_N4145) ) ;
 assign n872 = ( n812  &  n869 ) | ( n869  &  n870 ) | ( n812  &  (~ N_N4145) ) | ( n870  &  (~ N_N4145) ) ;
 assign n873 = ( n872  &  (~ N_N3912) ) ;
 assign n875 = ( n808  &  n872 ) | ( n872  &  n873 ) | ( n808  &  (~ N_N3912) ) | ( n873  &  (~ N_N3912) ) ;
 assign n876 = ( n875  &  (~ N_N4197) ) ;
 assign n878 = ( n804  &  n875 ) | ( n875  &  n876 ) | ( n804  &  (~ N_N4197) ) | ( n876  &  (~ N_N4197) ) ;
 assign n882 = ( (~ n880) ) | ( n1221 ) ;
 assign n880 = ( (~ N_N3462) ) | ( N_N3575 ) | ( (~ N_N4214) ) ;
 assign n881 = ( (~ n878)  &  n800 ) | ( n878  &  (~ n800) ) ;
 assign n879 = ( n882  &  n880 ) | ( n882  &  n881 ) ;
 assign n885 = ( (~ n875)  &  n1198 ) | ( n875  &  (~ n1198) ) ;
 assign n886 = ( PRESET ) | ( n880 ) ;
 assign n887 = ( PRESET ) | ( n882 ) ;
 assign n888 = ( n1185  &  n1199 ) | ( (~ n1185)  &  (~ n1199) ) ;
 assign n889 = ( n1187  &  n1200 ) | ( (~ n1187)  &  (~ n1200) ) ;
 assign n892 = ( n1189  &  n1201 ) | ( (~ n1189)  &  (~ n1201) ) ;
 assign n897 = ( (~ NLD3_9)  &  (~ n351) ) | ( (~ NLD3_9)  &  (~ N_N3971) ) | ( (~ n351)  &  (~ N_N3680) ) | ( (~ N_N3971)  &  (~ N_N3680) ) ;
 assign n895 = ( n460  &  n897 ) | ( n897  &  (~ N_N3681) ) ;
 assign n899 = ( n490  &  n522 ) | ( (~ n490)  &  (~ n522) ) ;
 assign n900 = ( n1191  &  n1202 ) | ( (~ n1191)  &  (~ n1202) ) ;
 assign n909 = ( PRESET ) | ( n1235 ) ;
 assign n914 = ( (~ n850)  &  n1203 ) | ( n850  &  (~ n1203) ) ;
 assign n916 = ( (~ n857)  &  n1204 ) | ( n857  &  (~ n1204) ) ;
 assign n918 = ( (~ n716)  &  n1288 ) | ( n716  &  (~ n1288) ) ;
 assign n926 = ( (~ n534)  &  n1289 ) | ( n534  &  (~ n1289) ) ;
 assign n929 = ( (~ n351)  &  n460 ) | ( n460  &  (~ N_N4252) ) | ( (~ n351)  &  (~ N_N3533) ) | ( (~ N_N4252)  &  (~ N_N3533) ) ;
 assign n927 = ( (~ NLD3_9)  &  n929 ) | ( n929  &  (~ N_N3791) ) ;
 assign n931 = ( (~ n351)  &  n460 ) | ( n460  &  (~ N_N3843) ) | ( (~ n351)  &  (~ N_N3105) ) | ( (~ N_N3843)  &  (~ N_N3105) ) ;
 assign n930 = ( (~ NLD3_9)  &  n931 ) | ( (~ N_N3489)  &  n931 ) ;
 assign n932 = ( (~ n684)  &  n1290 ) | ( n684  &  (~ n1290) ) ;
 assign n934 = ( (~ n698)  &  n1291 ) | ( n698  &  (~ n1291) ) ;
 assign n935 = ( (~ n710)  &  n1292 ) | ( n710  &  (~ n1292) ) ;
 assign n939 = ( (~ n691)  &  n1293 ) | ( n691  &  (~ n1293) ) ;
 assign n944 = ( PRESET ) | ( NLD3_9 ) ;
 assign n946 = ( NSr5_8 ) | ( PRESET ) ;
 assign n947 = ( (~ n676)  &  n1294 ) | ( n676  &  (~ n1294) ) ;
 assign n950 = ( (~ n866)  &  n1205 ) | ( n866  &  (~ n1205) ) ;
 assign n951 = ( (~ PDN)  &  (~ NLC1_2) ) ;
 assign n955 = ( n363  &  (~ N_N4212) ) | ( n413  &  (~ N_N4212) ) | ( n363  &  n1271 ) | ( n413  &  n1271 ) ;
 assign n954 = ( n955  &  n429 ) | ( n955  &  n880 ) ;
 assign n956 = ( PRESET ) | ( (~ n355) ) ;
 assign n958 = ( n367  &  (~ N_N4171) ) | ( n413  &  (~ N_N4171) ) | ( n367  &  n1271 ) | ( n413  &  n1271 ) ;
 assign n957 = ( n958  &  n437 ) | ( n958  &  n880 ) ;
 assign n961 = ( (~ n351)  &  n460 ) | ( n460  &  (~ N_N3918) ) | ( (~ n351)  &  (~ N_N3356) ) | ( (~ N_N3918)  &  (~ N_N3356) ) ;
 assign n960 = ( (~ NLD3_9)  &  n961 ) | ( n961  &  (~ N_N3709) ) ;
 assign n963 = ( (~ NLD3_9)  &  (~ n351) ) | ( (~ NLD3_9)  &  (~ N_N3939) ) | ( (~ n351)  &  (~ N_N3677) ) | ( (~ N_N3939)  &  (~ N_N3677) ) ;
 assign n962 = ( n460  &  n963 ) | ( n963  &  (~ N_N3741) ) ;
 assign n965 = ( (~ NLD3_9)  &  (~ n351) ) | ( (~ NLD3_9)  &  (~ N_N4224) ) | ( (~ n351)  &  (~ N_N3442) ) | ( (~ N_N4224)  &  (~ N_N3442) ) ;
 assign n964 = ( n460  &  n965 ) | ( n965  &  (~ N_N4106) ) ;
 assign n966 = ( (~ n412) ) | ( (~ N_N3949) ) ;
 assign n971 = ( (~ n350)  &  n1273 ) | ( (~ N_N3890)  &  n1273 ) | ( (~ n350)  &  (~ N_N3750) ) | ( (~ N_N3890)  &  (~ N_N3750) ) ;
 assign n969 = ( PRESET ) | ( n460 ) ;
 assign n980 = ( (~ NLD3_9)  &  (~ n351) ) | ( (~ NLD3_9)  &  (~ N_N4118) ) | ( (~ n351)  &  (~ N_N3179) ) | ( (~ N_N4118)  &  (~ N_N3179) ) ;
 assign n979 = ( n460  &  n980 ) | ( n980  &  (~ N_N4232) ) ;
 assign n983 = ( (~ NLD3_9)  &  (~ n351) ) | ( (~ N_N3336)  &  (~ n351) ) | ( (~ NLD3_9)  &  (~ N_N4209) ) | ( (~ N_N3336)  &  (~ N_N4209) ) ;
 assign n981 = ( n460  &  n983 ) | ( n983  &  (~ N_N3373) ) ;
 assign n987 = ( (~ n351)  &  n460 ) | ( n460  &  (~ N_N3500) ) | ( (~ n351)  &  (~ N_N3331) ) | ( (~ N_N3500)  &  (~ N_N3331) ) ;
 assign n985 = ( (~ NLD3_9)  &  n987 ) | ( n987  &  (~ N_N3464) ) ;
 assign n991 = ( (~ n706)  &  n1295 ) | ( n706  &  (~ n1295) ) ;
 assign n994 = ( (~ n350)  &  (~ N_N4079) ) | ( (~ N_N4176)  &  (~ N_N4079) ) | ( (~ n350)  &  n1273 ) | ( (~ N_N4176)  &  n1273 ) ;
 assign n997 = ( (~ n1206)  &  n1207 ) | ( n1206  &  (~ n1207) ) ;
 assign n999 = ( (~ n872)  &  n1208 ) | ( n872  &  (~ n1208) ) ;
 assign n1001 = ( n475  &  n602 ) | ( n475  &  (~ N_N4237) ) | ( n602  &  (~ N_N4236) ) | ( (~ N_N4237)  &  (~ N_N4236) ) ;
 assign n1003 = ( n475  &  n602 ) | ( n602  &  (~ N_N4208) ) | ( n475  &  (~ N_N4209) ) | ( (~ N_N4208)  &  (~ N_N4209) ) ;
 assign n1005 = ( n720  &  n645 ) ;
 assign n1006 = ( n642  &  n645 ) | ( n1005  &  n645 ) | ( n642  &  n720 ) | ( n1005  &  n720 ) ;
 assign n1007 = ( (~ n1006)  &  n1296 ) | ( n1006  &  (~ n1296) ) ;
 assign n1014 = ( (~ n351)  &  n460 ) | ( n460  &  (~ N_N3842) ) | ( (~ n351)  &  (~ N_N3196) ) | ( (~ N_N3842)  &  (~ N_N3196) ) ;
 assign n1012 = ( (~ NLD3_9)  &  n1014 ) | ( n1014  &  (~ N_N3212) ) ;
 assign n1016 = ( (~ n351)  &  n460 ) | ( n460  &  (~ N_N3924) ) | ( (~ n351)  &  (~ N_N3250) ) | ( (~ N_N3924)  &  (~ N_N3250) ) ;
 assign n1015 = ( (~ NLD3_9)  &  n1016 ) | ( (~ N_N3981)  &  n1016 ) ;
 assign n1018 = ( (~ NLD3_9)  &  (~ n351) ) | ( (~ n351)  &  (~ N_N3535) ) | ( (~ NLD3_9)  &  (~ N_N4119) ) | ( (~ N_N3535)  &  (~ N_N4119) ) ;
 assign n1017 = ( n460  &  n1018 ) | ( n1018  &  (~ N_N3580) ) ;
 assign n1031 = ( (~ n351)  &  n460 ) | ( n460  &  (~ N_N3808) ) | ( (~ n351)  &  (~ N_N3062) ) | ( (~ N_N3808)  &  (~ N_N3062) ) ;
 assign n1030 = ( (~ NLD3_9)  &  n1031 ) | ( n1031  &  (~ N_N3513) ) ;
 assign n1034 = ( n402  &  (~ N_N3340) ) | ( n413  &  (~ N_N3340) ) | ( n402  &  n1271 ) | ( n413  &  n1271 ) ;
 assign n1033 = ( (~ N_N3340)  &  n1183 ) | ( N_N3340  &  (~ n1183) ) ;
 assign n1032 = ( n1034  &  n1033 ) | ( n1034  &  n880 ) ;
 assign n1041 = ( (~ n350)  &  (~ N_N3931) ) | ( (~ N_N3810)  &  (~ N_N3931) ) | ( (~ n350)  &  n1273 ) | ( (~ N_N3810)  &  n1273 ) ;
 assign n1042 = ( (~ n350)  &  (~ N_N3875) ) | ( (~ N_N3844)  &  (~ N_N3875) ) | ( (~ n350)  &  n1273 ) | ( (~ N_N3844)  &  n1273 ) ;
 assign n1047 = ( (~ n353)  &  n371 ) | ( (~ n353)  &  n416 ) | ( n371  &  (~ N_N4126) ) | ( n416  &  (~ N_N4126) ) ;
 assign n1048 = ( (~ n353)  &  n389 ) | ( (~ n353)  &  n416 ) | ( n389  &  (~ N_N4246) ) | ( n416  &  (~ N_N4246) ) ;
 assign n1049 = ( (~ n585)  &  n1209 ) | ( n585  &  (~ n1209) ) ;
 assign n1050 = ( n1184  &  n1210 ) | ( (~ n1184)  &  (~ n1210) ) ;
 assign n1052 = ( (~ NLD3_9)  &  (~ n351) ) | ( (~ NLD3_9)  &  (~ N_N3940) ) | ( (~ n351)  &  (~ N_N4111) ) | ( (~ N_N3940)  &  (~ N_N4111) ) ;
 assign n1051 = ( n460  &  n1052 ) | ( n1052  &  (~ N_N4218) ) ;
 assign n1058 = ( n1186  &  n1211 ) | ( (~ n1186)  &  (~ n1211) ) ;
 assign n1059 = ( n1188  &  n1212 ) | ( (~ n1188)  &  (~ n1212) ) ;
 assign n1061 = ( NSr5_7 ) | ( PRESET ) ;
 assign n1063 = ( (~ NLD3_9)  &  (~ n351) ) | ( (~ NLD3_9)  &  (~ N_N3923) ) | ( (~ n351)  &  (~ N_N3475) ) | ( (~ N_N3923)  &  (~ N_N3475) ) ;
 assign n1062 = ( n460  &  n1063 ) | ( n1063  &  (~ N_N4230) ) ;
 assign n1064 = ( (~ n869)  &  n1213 ) | ( n869  &  (~ n1213) ) ;
 assign n1066 = ( (~ n350)  &  (~ N_N3908) ) | ( (~ N_N3800)  &  (~ N_N3908) ) | ( (~ n350)  &  n1273 ) | ( (~ N_N3800)  &  n1273 ) ;
 assign n1067 = ( (~ n854)  &  n1214 ) | ( n854  &  (~ n1214) ) ;
 assign n1072 = ( (~ n350)  &  n1273 ) | ( (~ N_N4136)  &  n1273 ) | ( (~ n350)  &  (~ N_N3516) ) | ( (~ N_N4136)  &  (~ N_N3516) ) ;
 assign n1073 = ( (~ n350)  &  n1273 ) | ( (~ N_N4183)  &  n1273 ) | ( (~ n350)  &  (~ N_N3420) ) | ( (~ N_N4183)  &  (~ N_N3420) ) ;
 assign n1082 = ( n394  &  (~ N_N3369) ) | ( n413  &  (~ N_N3369) ) | ( n394  &  n1271 ) | ( n413  &  n1271 ) ;
 assign n1081 = ( n1082  &  n418 ) | ( n1082  &  n880 ) ;
 assign n1086 = ( (~ n350)  &  (~ N_N3862) ) | ( (~ N_N3862)  &  (~ N_N3813) ) | ( (~ n350)  &  n1273 ) | ( (~ N_N3813)  &  n1273 ) ;
 assign n1091 = ( n398  &  (~ N_N4093) ) | ( n413  &  (~ N_N4093) ) | ( n398  &  n1271 ) | ( n413  &  n1271 ) ;
 assign n1090 = ( n1091  &  n425 ) | ( n1091  &  n880 ) ;
 assign n1100 = ( (~ n350)  &  (~ N_N4158) ) | ( (~ N_N4208)  &  (~ N_N4158) ) | ( (~ n350)  &  n1273 ) | ( (~ N_N4208)  &  n1273 ) ;
 assign n1102 = ( (~ n350)  &  (~ N_N3713) ) | ( (~ N_N3807)  &  (~ N_N3713) ) | ( (~ n350)  &  n1273 ) | ( (~ N_N3807)  &  n1273 ) ;
 assign n1105 = ( (~ n351)  &  n460 ) | ( n460  &  (~ N_N3872) ) | ( (~ n351)  &  (~ N_N3248) ) | ( (~ N_N3872)  &  (~ N_N3248) ) ;
 assign n1104 = ( (~ NLD3_9)  &  n1105 ) | ( n1105  &  (~ N_N3761) ) ;
 assign n1108 = ( (~ N_N3965)  &  n844 ) | ( N_N3965  &  (~ n844) ) ;
 assign n1115 = ( (~ n353)  &  n384 ) | ( (~ n353)  &  n416 ) | ( n384  &  (~ N_N4036) ) | ( n416  &  (~ N_N4036) ) ;
 assign n1116 = ( (~ n353)  &  n380 ) | ( (~ n353)  &  n416 ) | ( n380  &  (~ N_N4004) ) | ( n416  &  (~ N_N4004) ) ;
 assign n1118 = ( (~ n351)  &  n460 ) | ( n460  &  (~ N_N4177) ) | ( (~ n351)  &  (~ N_N3011) ) | ( (~ N_N4177)  &  (~ N_N3011) ) ;
 assign n1117 = ( (~ NLD3_9)  &  n1118 ) | ( (~ N_N3884)  &  n1118 ) ;
 assign n1129 = ( n406  &  (~ N_N3283) ) | ( n413  &  (~ N_N3283) ) | ( n406  &  n1271 ) | ( n413  &  n1271 ) ;
 assign n1128 = ( (~ N_N3283)  &  n421 ) | ( N_N3283  &  (~ n421) ) ;
 assign n1127 = ( n1129  &  n1128 ) | ( n1129  &  n880 ) ;
 assign n1138 = ( (~ n350)  &  (~ N_N3821) ) | ( (~ N_N3470)  &  (~ N_N3821) ) | ( (~ n350)  &  n1273 ) | ( (~ N_N3470)  &  n1273 ) ;
 assign n1141 = ( (~ n860)  &  n1216 ) | ( n860  &  (~ n1216) ) ;
 assign n1162 = ( (~ n840)  &  n1275 ) | ( n840  &  (~ n1275) ) ;
 assign n1172 = ( (~ n353)  &  n376 ) | ( (~ n353)  &  n416 ) | ( n376  &  (~ N_N3961) ) | ( n416  &  (~ N_N3961) ) ;
 assign n1173 = ( (~ n863)  &  n1217 ) | ( n863  &  (~ n1217) ) ;
 assign n1178 = ( (~ n350)  &  (~ N_N3832) ) | ( (~ N_N3868)  &  (~ N_N3832) ) | ( (~ n350)  &  n1273 ) | ( (~ N_N3868)  &  n1273 ) ;
 assign n1179 = ( (~ n350)  &  (~ N_N3794) ) | ( (~ N_N3794)  &  (~ N_N3919) ) | ( (~ n350)  &  n1273 ) | ( (~ N_N3919)  &  n1273 ) ;
 assign n1180 = ( (~ n350)  &  (~ N_N3214) ) | ( (~ N_N3871)  &  (~ N_N3214) ) | ( (~ n350)  &  n1273 ) | ( (~ N_N3871)  &  n1273 ) ;
 assign N_N3542 = ( n72  &  (~ NSr3_9) ) ;
 assign n1181 = ( (~ PRESET)  &  Pover_0_0_  &  (~ NGFDN_3) ) | ( (~ PRESET)  &  Pover_0_0_  &  NDN3_11 ) ;
 assign N_N3061 = ( N_N3542 ) | ( n1181 ) ;
 assign n1182 = ( (~ PRESET)  &  Pnext_0_0_  &  (~ NLD3_9) ) | ( (~ PRESET)  &  Pnext_0_0_  &  NDN5_16 ) ;
 assign N_N3042 = ( (~ PRESET)  &  n1227 ) ;
 assign N_N3005 = ( n1182 ) | ( N_N3042 ) ;
 assign n1183 = ( N_N3283 ) | ( n421 ) ;
 assign n1184 = ( (~ n536)  &  n493 ) | ( n536  &  (~ n493) ) ;
 assign n1185 = ( (~ n550)  &  n499 ) | ( n550  &  (~ n499) ) ;
 assign n1186 = ( (~ n549)  &  n487 ) | ( n549  &  (~ n487) ) ;
 assign n1187 = ( (~ n564)  &  n502 ) | ( n564  &  (~ n502) ) ;
 assign n1188 = ( (~ n563)  &  n484 ) | ( n563  &  (~ n484) ) ;
 assign n1189 = ( (~ n518)  &  n505 ) | ( n518  &  (~ n505) ) ;
 assign n1192 = ( n505  &  n481  &  n518 ) ;
 assign n1191 = ( (~ n1192)  &  n508 ) | ( n1192  &  (~ n508) ) ;
 assign n1195 = ( (~ n584)  &  n586 ) | ( n584  &  (~ n586) ) ;
 assign n1196 = ( (~ n473)  &  n1284 ) | ( n473  &  (~ n1284) ) ;
 assign n1194 = ( (~ n1195)  &  n1196 ) | ( n1195  &  (~ n1196) ) ;
 assign n1197 = ( (~ n573)  &  n514 ) | ( n573  &  (~ n514) ) ;
 assign n1198 = ( n804  &  N_N4197 ) | ( (~ n804)  &  (~ N_N4197) ) ;
 assign n1199 = ( (~ n542)  &  n519 ) | ( n542  &  (~ n519) ) ;
 assign n1200 = ( (~ n553)  &  n554 ) | ( n553  &  (~ n554) ) ;
 assign n1201 = ( (~ n567)  &  n568 ) | ( n567  &  (~ n568) ) ;
 assign n1202 = ( (~ n576)  &  n577 ) | ( n576  &  (~ n577) ) ;
 assign n1203 = ( n836  &  N_N3992 ) | ( (~ n836)  &  (~ N_N3992) ) ;
 assign n1204 = ( n828  &  N_N4018 ) | ( (~ n828)  &  (~ N_N4018) ) ;
 assign n1205 = ( n816  &  N_N3949 ) | ( (~ n816)  &  (~ N_N3949) ) ;
 assign n1206 = ( (~ n665)  &  n668 ) | ( n665  &  (~ n668) ) ;
 assign n1207 = ( n604 ) | ( n600 ) ;
 assign n1208 = ( n808  &  N_N3912 ) | ( (~ n808)  &  (~ N_N3912) ) ;
 assign n1209 = ( (~ n581)  &  n511 ) | ( n581  &  (~ n511) ) ;
 assign n1210 = ( (~ n533)  &  n537 ) | ( n533  &  (~ n537) ) ;
 assign n1211 = ( (~ n544)  &  n546 ) | ( n544  &  (~ n546) ) ;
 assign n1212 = ( (~ n559)  &  n560 ) | ( n559  &  (~ n560) ) ;
 assign n1213 = ( n812  &  N_N4145 ) | ( (~ n812)  &  (~ N_N4145) ) ;
 assign n1214 = ( n832  &  N_N3996 ) | ( (~ n832)  &  (~ N_N3996) ) ;
 assign n1216 = ( n824  &  N_N3974 ) | ( (~ n824)  &  (~ N_N3974) ) ;
 assign n1217 = ( n820  &  N_N4083 ) | ( (~ n820)  &  (~ N_N4083) ) ;
 assign n1221 = ( n2  &  (~ N_N4214) ) ;
 assign n1226 = ( n425  &  n422  &  n418  &  n437  &  n433  &  n429 ) ;
 assign n1227 = ( (~ NLD3_9)  &  NDN5_9 ) ;
 assign n1228 = ( (~ PDN) ) | ( NDN1_4 ) ;
 assign n1230 = ( (~ Preset_0_0_)  &  (~ NLC1_2) ) | ( (~ Preset_0_0_)  &  N_N3998 ) | ( NLC1_2  &  N_N3998 ) ;
 assign n1233 = ( (~ NDN3_3)  &  (~ NSr3_2) ) ;
 assign n1235 = ( NDN2_2 ) | ( n149 ) ;
 assign n1237 = ( (~ PRESET)  &  n476 ) ;
 assign n1238 = ( n508  &  n1192 ) ;
 assign n1242 = ( NSr5_8 ) | ( NDN5_8 ) ;
 assign n1245 = ( NSr5_4 ) | ( NDN5_4 ) ;
 assign n1247 = ( NSr5_7 ) | ( NDN5_7 ) ;
 assign n1250 = ( NSr5_3 ) | ( NDN5_3 ) ;
 assign n1252 = ( NSr5_5 ) | ( NDN5_5 ) ;
 assign n1254 = ( NSr5_2 ) | ( NDN5_2 ) ;
 assign n1271 = ( (~ n412) ) | ( n414 ) ;
 assign n1273 = ( PRESET ) | ( (~ NLD3_9) ) ;
 assign n1275 = ( n849  &  N_N4027 ) | ( (~ n849)  &  (~ N_N4027) ) ;
 assign n1276 = ( PRESET  &  n1283 ) | ( n879  &  n1283 ) | ( (~ N_N4227)  &  n1283 ) ;
 assign N_N3859 = ( (~ n1276) ) ;
 assign n1277 = ( n371  &  n367  &  n363  &  n384  &  n380  &  n376 ) ;
 assign n1283 = ( (~ n881) ) | ( n886 ) | ( N_N4227 ) ;
 assign N_N3538 = ( (~ n1061) ) ;
 assign N_N3029 = ( (~ n946) ) ;
 assign n1284 = ( n1238  &  n478 ) ;
 assign n1285 = ( n490 ) | ( n522 ) ;
 assign n1286 = ( (~ n642)  &  n645 ) | ( n642  &  (~ n645) ) ;
 assign n1287 = ( (~ n653)  &  n656 ) | ( n653  &  (~ n656) ) ;
 assign n1288 = ( (~ n712)  &  n713 ) | ( n712  &  (~ n713) ) ;
 assign n1289 = ( (~ n525)  &  n1285 ) | ( n525  &  (~ n1285) ) ;
 assign n1290 = ( (~ n681)  &  n682 ) | ( n681  &  (~ n682) ) ;
 assign n1291 = ( (~ n695)  &  n696 ) | ( n695  &  (~ n696) ) ;
 assign n1292 = ( (~ n648)  &  n650 ) | ( n648  &  (~ n650) ) ;
 assign n1293 = ( (~ n688)  &  n689 ) | ( n688  &  (~ n689) ) ;
 assign n1294 = ( (~ n659)  &  n662 ) | ( n659  &  (~ n662) ) ;
 assign n1295 = ( (~ n702)  &  n703 ) | ( n702  &  (~ n703) ) ;
 assign n1296 = ( (~ n1001)  &  n1003 ) | ( n1001  &  (~ n1003) ) ;
 assign n1297 = ( (~ N_N3999)  &  n358  &  n389  &  n394  &  n398  &  n402  &  n406  &  n1277 ) ;
 assign n1299 = ( (~ Preset_0_0_)  &  n951 ) ;


endmodule

