module ks_bar_qmap_map (sk, shiftx6x, shiftx4x, shiftx5x, shiftx2x, shiftx3x, ax16x, ax15x, ax14x, ax13x, shiftx0x, shiftx1x, ax12x, ax11x, ax10x, ax9x, ax4x, ax3x, ax2x, ax1x, ax8x, ax7x, ax6x, ax5x, ax32x, ax31x, ax30x, ax29x, ax28x, ax27x, ax26x, ax25x, ax20x, ax19x, ax18x, ax17x, ax24x, ax23x, ax22x, ax21x, ax64x, ax63x, ax62x, ax61x, ax60x, ax59x, ax58x, ax57x, ax52x, ax51x, ax50x, ax49x, ax56x, ax55x, ax54x, ax53x, ax48x, ax47x, ax46x, ax45x, ax44x, ax43x, ax42x, ax41x, ax36x, ax35x, ax34x, ax33x, ax40x, ax38x, ax39x, ax37x, ax80x, ax79x, ax78x, ax77x, ax76x, ax75x, ax74x, ax73x, ax68x, ax67x, ax66x, ax65x, ax72x, ax71x, ax70x, ax69x, ax96x, ax95x, ax94x, ax93x, ax92x, ax91x, ax90x, ax89x, ax84x, ax83x, ax82x, ax81x, ax88x, ax87x, ax86x, ax85x, ax0x, ax127x, ax126x, ax125x, ax124x, ax123x, ax122x, ax121x, ax116x, ax115x, ax114x, ax113x, ax120x, ax119x, ax118x, ax117x, ax112x, ax111x, ax110x, ax109x, ax108x, ax107x, ax106x, ax105x, ax100x, ax99x, ax98x, ax97x, ax104x, ax103x, ax102x, ax101x, resultx0x, resultx1x, resultx2x, resultx3x, resultx4x, resultx5x, resultx6x, resultx7x, resultx8x, resultx9x, resultx10x, resultx11x, resultx12x, resultx13x, resultx14x, resultx15x, resultx16x, resultx17x, resultx18x, resultx19x, resultx20x, resultx21x, resultx22x, resultx23x, resultx24x, resultx25x, resultx26x, resultx27x, resultx28x, resultx29x, resultx30x, resultx31x, resultx32x, resultx33x, resultx34x, resultx35x, resultx36x, resultx37x, resultx38x, resultx39x, resultx40x, resultx41x, resultx42x, resultx43x, resultx44x, resultx45x, resultx46x, resultx47x, resultx48x, resultx49x, resultx50x, resultx51x, resultx52x, resultx53x, resultx54x, resultx55x, resultx56x, resultx57x, resultx58x, resultx59x, resultx60x, resultx61x, resultx62x, resultx63x, resultx64x, resultx65x, resultx66x, resultx67x, resultx68x, resultx69x, resultx70x, resultx71x, resultx72x, resultx73x, resultx74x, resultx75x, resultx76x, resultx77x, resultx78x, resultx79x, resultx80x, resultx81x, resultx82x, resultx83x, resultx84x, resultx85x, resultx86x, resultx87x, resultx88x, resultx89x, resultx90x, resultx91x, resultx92x, resultx93x, resultx94x, resultx95x, resultx96x, resultx97x, resultx98x, resultx99x, resultx100x, resultx101x, resultx102x, resultx103x, resultx104x, resultx105x, resultx106x, resultx107x, resultx108x, resultx109x, resultx110x, resultx111x, resultx112x, resultx113x, resultx114x, resultx115x, resultx116x, resultx117x, resultx118x, resultx119x, resultx120x, resultx121x, resultx122x, resultx123x, resultx124x, resultx125x, resultx126x, resultx127x);

	input shiftx6x;
	input shiftx4x;
	input shiftx5x;
	input shiftx2x;
	input shiftx3x;
	input ax16x;
	input ax15x;
	input ax14x;
	input ax13x;
	input shiftx0x;
	input shiftx1x;
	input ax12x;
	input ax11x;
	input ax10x;
	input ax9x;
	input ax4x;
	input ax3x;
	input ax2x;
	input ax1x;
	input ax8x;
	input ax7x;
	input ax6x;
	input ax5x;
	input ax32x;
	input ax31x;
	input ax30x;
	input ax29x;
	input ax28x;
	input ax27x;
	input ax26x;
	input ax25x;
	input ax20x;
	input ax19x;
	input ax18x;
	input ax17x;
	input ax24x;
	input ax23x;
	input ax22x;
	input ax21x;
	input ax64x;
	input ax63x;
	input ax62x;
	input ax61x;
	input ax60x;
	input ax59x;
	input ax58x;
	input ax57x;
	input ax52x;
	input ax51x;
	input ax50x;
	input ax49x;
	input ax56x;
	input ax55x;
	input ax54x;
	input ax53x;
	input ax48x;
	input ax47x;
	input ax46x;
	input ax45x;
	input ax44x;
	input ax43x;
	input ax42x;
	input ax41x;
	input ax36x;
	input ax35x;
	input ax34x;
	input ax33x;
	input ax40x;
	input ax38x;
	input ax39x;
	input ax37x;
	input ax80x;
	input ax79x;
	input ax78x;
	input ax77x;
	input ax76x;
	input ax75x;
	input ax74x;
	input ax73x;
	input ax68x;
	input ax67x;
	input ax66x;
	input ax65x;
	input ax72x;
	input ax71x;
	input ax70x;
	input ax69x;
	input ax96x;
	input ax95x;
	input ax94x;
	input ax93x;
	input ax92x;
	input ax91x;
	input ax90x;
	input ax89x;
	input ax84x;
	input ax83x;
	input ax82x;
	input ax81x;
	input ax88x;
	input ax87x;
	input ax86x;
	input ax85x;
	input ax0x;
	input ax127x;
	input ax126x;
	input ax125x;
	input ax124x;
	input ax123x;
	input ax122x;
	input ax121x;
	input ax116x;
	input ax115x;
	input ax114x;
	input ax113x;
	input ax120x;
	input ax119x;
	input ax118x;
	input ax117x;
	input ax112x;
	input ax111x;
	input ax110x;
	input ax109x;
	input ax108x;
	input ax107x;
	input ax106x;
	input ax105x;
	input ax100x;
	input ax99x;
	input ax98x;
	input ax97x;
	input ax104x;
	input ax103x;
	input ax102x;
	input ax101x;
	output resultx0x;
	output resultx1x;
	output resultx2x;
	output resultx3x;
	output resultx4x;
	output resultx5x;
	output resultx6x;
	output resultx7x;
	output resultx8x;
	output resultx9x;
	output resultx10x;
	output resultx11x;
	output resultx12x;
	output resultx13x;
	output resultx14x;
	output resultx15x;
	output resultx16x;
	output resultx17x;
	output resultx18x;
	output resultx19x;
	output resultx20x;
	output resultx21x;
	output resultx22x;
	output resultx23x;
	output resultx24x;
	output resultx25x;
	output resultx26x;
	output resultx27x;
	output resultx28x;
	output resultx29x;
	output resultx30x;
	output resultx31x;
	output resultx32x;
	output resultx33x;
	output resultx34x;
	output resultx35x;
	output resultx36x;
	output resultx37x;
	output resultx38x;
	output resultx39x;
	output resultx40x;
	output resultx41x;
	output resultx42x;
	output resultx43x;
	output resultx44x;
	output resultx45x;
	output resultx46x;
	output resultx47x;
	output resultx48x;
	output resultx49x;
	output resultx50x;
	output resultx51x;
	output resultx52x;
	output resultx53x;
	output resultx54x;
	output resultx55x;
	output resultx56x;
	output resultx57x;
	output resultx58x;
	output resultx59x;
	output resultx60x;
	output resultx61x;
	output resultx62x;
	output resultx63x;
	output resultx64x;
	output resultx65x;
	output resultx66x;
	output resultx67x;
	output resultx68x;
	output resultx69x;
	output resultx70x;
	output resultx71x;
	output resultx72x;
	output resultx73x;
	output resultx74x;
	output resultx75x;
	output resultx76x;
	output resultx77x;
	output resultx78x;
	output resultx79x;
	output resultx80x;
	output resultx81x;
	output resultx82x;
	output resultx83x;
	output resultx84x;
	output resultx85x;
	output resultx86x;
	output resultx87x;
	output resultx88x;
	output resultx89x;
	output resultx90x;
	output resultx91x;
	output resultx92x;
	output resultx93x;
	output resultx94x;
	output resultx95x;
	output resultx96x;
	output resultx97x;
	output resultx98x;
	output resultx99x;
	output resultx100x;
	output resultx101x;
	output resultx102x;
	output resultx103x;
	output resultx104x;
	output resultx105x;
	output resultx106x;
	output resultx107x;
	output resultx108x;
	output resultx109x;
	output resultx110x;
	output resultx111x;
	output resultx112x;
	output resultx113x;
	output resultx114x;
	output resultx115x;
	output resultx116x;
	output resultx117x;
	output resultx118x;
	output resultx119x;
	output resultx120x;
	output resultx121x;
	output resultx122x;
	output resultx123x;
	output resultx124x;
	output resultx125x;
	output resultx126x;
	output resultx127x;

	input [127 : 0] sk /* synthesis noprune */;


	wire g1, g2, g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g20, g21;
	wire g22, g23, g24, g25, g26, g27, g28, g29, g30, g31, g32, g33, g34, g35, g36, g37, g38, g39, g40, g41, g42;
	wire g44, g45, g46, g47, g48, g49, g50, g51, g52, g53, g54, g55, g56, g57, g58, g59, g60, g61, g62, g63, g64;
	wire g65, g66, g67, g68, g69, g70, g71, g72, g73, g74, g75, g76, g77, g78, g79, g80, g81, g82, g83, g84, g85;
	wire g87, g88, g89, g90, g91, g92, g93, g94, g95, g96, g97, g98, g99, g100, g101, g102, g103, g104, g105, g106, g107;
	wire g108, g109, g110, g111, g112, g113, g114, g115, g116, g117, g118, g119, g120, g121, g122, g123, g124, g125, g126, g127, g128;
	wire g130, g131, g132, g133, g134, g135, g136, g137, g138, g139, g140, g141, g142, g143, g144, g145, g146, g147, g148, g149, g150;
	wire g151, g152, g153, g154, g155, g156, g157, g158, g159, g160, g161, g162, g163, g164, g165, g166, g167, g168, g169, g170, g171;
	wire g173, g174, g175, g176, g177, g178, g179, g180, g181, g182, g184, g185, g186, g187, g188, g189, g190, g191, g192, g193, g195;
	wire g196, g197, g198, g199, g200, g201, g202, g203, g204, g206, g207, g208, g209, g210, g211, g212, g213, g214, g215, g217, g218;
	wire g219, g220, g221, g222, g223, g224, g225, g226, g228, g229, g230, g231, g232, g233, g234, g235, g236, g237, g239, g240, g241;
	wire g242, g243, g244, g245, g246, g247, g248, g250, g251, g252, g253, g254, g255, g256, g257, g258, g259, g261, g262, g263, g264;
	wire g265, g266, g267, g268, g269, g270, g272, g273, g274, g275, g276, g277, g278, g279, g280, g281, g283, g284, g285, g286, g287;
	wire g288, g289, g290, g291, g292, g294, g295, g296, g297, g298, g299, g300, g301, g302, g303, g305, g306, g308, g309, g311, g312;
	wire g314, g315, g317, g318, g320, g321, g323, g324, g326, g327, g329, g330, g332, g333, g335, g336, g338, g339, g341, g342, g344;
	wire g345, g347, g348, g350, g351, g353, g354, g356, g357, g359, g360, g362, g363, g365, g366, g368, g369, g371, g372, g374, g375;
	wire g377, g378, g380, g381, g383, g384, g386, g387, g389, g390, g392, g393, g395, g396, g398, g399, g401, g402, g404, g405, g407;
	wire g408, g410, g411, g413, g414, g416, g417, g419, g420, g422, g423, g425, g426, g428, g429, g431, g432, g434, g435, g437, g438;
	wire g440, g441, g443, g444, g446, g447;

	assign g1 = (((!ax16x) & (!ax15x) & (!ax14x) & (ax13x) & (shiftx0x) & (shiftx1x)) + ((!ax16x) & (!ax15x) & (ax14x) & (!ax13x) & (!shiftx0x) & (shiftx1x)) + ((!ax16x) & (!ax15x) & (ax14x) & (ax13x) & (!shiftx0x) & (shiftx1x)) + ((!ax16x) & (!ax15x) & (ax14x) & (ax13x) & (shiftx0x) & (shiftx1x)) + ((!ax16x) & (ax15x) & (!ax14x) & (!ax13x) & (shiftx0x) & (!shiftx1x)) + ((!ax16x) & (ax15x) & (!ax14x) & (ax13x) & (shiftx0x) & (!shiftx1x)) + ((!ax16x) & (ax15x) & (!ax14x) & (ax13x) & (shiftx0x) & (shiftx1x)) + ((!ax16x) & (ax15x) & (ax14x) & (!ax13x) & (!shiftx0x) & (shiftx1x)) + ((!ax16x) & (ax15x) & (ax14x) & (!ax13x) & (shiftx0x) & (!shiftx1x)) + ((!ax16x) & (ax15x) & (ax14x) & (ax13x) & (!shiftx0x) & (shiftx1x)) + ((!ax16x) & (ax15x) & (ax14x) & (ax13x) & (shiftx0x) & (!shiftx1x)) + ((!ax16x) & (ax15x) & (ax14x) & (ax13x) & (shiftx0x) & (shiftx1x)) + ((ax16x) & (!ax15x) & (!ax14x) & (!ax13x) & (!shiftx0x) & (!shiftx1x)) + ((ax16x) & (!ax15x) & (!ax14x) & (ax13x) & (!shiftx0x) & (!shiftx1x)) + ((ax16x) & (!ax15x) & (!ax14x) & (ax13x) & (shiftx0x) & (shiftx1x)) + ((ax16x) & (!ax15x) & (ax14x) & (!ax13x) & (!shiftx0x) & (!shiftx1x)) + ((ax16x) & (!ax15x) & (ax14x) & (!ax13x) & (!shiftx0x) & (shiftx1x)) + ((ax16x) & (!ax15x) & (ax14x) & (ax13x) & (!shiftx0x) & (!shiftx1x)) + ((ax16x) & (!ax15x) & (ax14x) & (ax13x) & (!shiftx0x) & (shiftx1x)) + ((ax16x) & (!ax15x) & (ax14x) & (ax13x) & (shiftx0x) & (shiftx1x)) + ((ax16x) & (ax15x) & (!ax14x) & (!ax13x) & (!shiftx0x) & (!shiftx1x)) + ((ax16x) & (ax15x) & (!ax14x) & (!ax13x) & (shiftx0x) & (!shiftx1x)) + ((ax16x) & (ax15x) & (!ax14x) & (ax13x) & (!shiftx0x) & (!shiftx1x)) + ((ax16x) & (ax15x) & (!ax14x) & (ax13x) & (shiftx0x) & (!shiftx1x)) + ((ax16x) & (ax15x) & (!ax14x) & (ax13x) & (shiftx0x) & (shiftx1x)) + ((ax16x) & (ax15x) & (ax14x) & (!ax13x) & (!shiftx0x) & (!shiftx1x)) + ((ax16x) & (ax15x) & (ax14x) & (!ax13x) & (!shiftx0x) & (shiftx1x)) + ((ax16x) & (ax15x) & (ax14x) & (!ax13x) & (shiftx0x) & (!shiftx1x)) + ((ax16x) & (ax15x) & (ax14x) & (ax13x) & (!shiftx0x) & (!shiftx1x)) + ((ax16x) & (ax15x) & (ax14x) & (ax13x) & (!shiftx0x) & (shiftx1x)) + ((ax16x) & (ax15x) & (ax14x) & (ax13x) & (shiftx0x) & (!shiftx1x)) + ((ax16x) & (ax15x) & (ax14x) & (ax13x) & (shiftx0x) & (shiftx1x)));
	assign g2 = (((!ax12x) & (!ax11x) & (!ax10x) & (ax9x) & (shiftx0x) & (shiftx1x)) + ((!ax12x) & (!ax11x) & (ax10x) & (!ax9x) & (!shiftx0x) & (shiftx1x)) + ((!ax12x) & (!ax11x) & (ax10x) & (ax9x) & (!shiftx0x) & (shiftx1x)) + ((!ax12x) & (!ax11x) & (ax10x) & (ax9x) & (shiftx0x) & (shiftx1x)) + ((!ax12x) & (ax11x) & (!ax10x) & (!ax9x) & (shiftx0x) & (!shiftx1x)) + ((!ax12x) & (ax11x) & (!ax10x) & (ax9x) & (shiftx0x) & (!shiftx1x)) + ((!ax12x) & (ax11x) & (!ax10x) & (ax9x) & (shiftx0x) & (shiftx1x)) + ((!ax12x) & (ax11x) & (ax10x) & (!ax9x) & (!shiftx0x) & (shiftx1x)) + ((!ax12x) & (ax11x) & (ax10x) & (!ax9x) & (shiftx0x) & (!shiftx1x)) + ((!ax12x) & (ax11x) & (ax10x) & (ax9x) & (!shiftx0x) & (shiftx1x)) + ((!ax12x) & (ax11x) & (ax10x) & (ax9x) & (shiftx0x) & (!shiftx1x)) + ((!ax12x) & (ax11x) & (ax10x) & (ax9x) & (shiftx0x) & (shiftx1x)) + ((ax12x) & (!ax11x) & (!ax10x) & (!ax9x) & (!shiftx0x) & (!shiftx1x)) + ((ax12x) & (!ax11x) & (!ax10x) & (ax9x) & (!shiftx0x) & (!shiftx1x)) + ((ax12x) & (!ax11x) & (!ax10x) & (ax9x) & (shiftx0x) & (shiftx1x)) + ((ax12x) & (!ax11x) & (ax10x) & (!ax9x) & (!shiftx0x) & (!shiftx1x)) + ((ax12x) & (!ax11x) & (ax10x) & (!ax9x) & (!shiftx0x) & (shiftx1x)) + ((ax12x) & (!ax11x) & (ax10x) & (ax9x) & (!shiftx0x) & (!shiftx1x)) + ((ax12x) & (!ax11x) & (ax10x) & (ax9x) & (!shiftx0x) & (shiftx1x)) + ((ax12x) & (!ax11x) & (ax10x) & (ax9x) & (shiftx0x) & (shiftx1x)) + ((ax12x) & (ax11x) & (!ax10x) & (!ax9x) & (!shiftx0x) & (!shiftx1x)) + ((ax12x) & (ax11x) & (!ax10x) & (!ax9x) & (shiftx0x) & (!shiftx1x)) + ((ax12x) & (ax11x) & (!ax10x) & (ax9x) & (!shiftx0x) & (!shiftx1x)) + ((ax12x) & (ax11x) & (!ax10x) & (ax9x) & (shiftx0x) & (!shiftx1x)) + ((ax12x) & (ax11x) & (!ax10x) & (ax9x) & (shiftx0x) & (shiftx1x)) + ((ax12x) & (ax11x) & (ax10x) & (!ax9x) & (!shiftx0x) & (!shiftx1x)) + ((ax12x) & (ax11x) & (ax10x) & (!ax9x) & (!shiftx0x) & (shiftx1x)) + ((ax12x) & (ax11x) & (ax10x) & (!ax9x) & (shiftx0x) & (!shiftx1x)) + ((ax12x) & (ax11x) & (ax10x) & (ax9x) & (!shiftx0x) & (!shiftx1x)) + ((ax12x) & (ax11x) & (ax10x) & (ax9x) & (!shiftx0x) & (shiftx1x)) + ((ax12x) & (ax11x) & (ax10x) & (ax9x) & (shiftx0x) & (!shiftx1x)) + ((ax12x) & (ax11x) & (ax10x) & (ax9x) & (shiftx0x) & (shiftx1x)));
	assign g3 = (((!ax4x) & (!ax3x) & (!ax2x) & (ax1x) & (shiftx0x) & (shiftx1x)) + ((!ax4x) & (!ax3x) & (ax2x) & (!ax1x) & (!shiftx0x) & (shiftx1x)) + ((!ax4x) & (!ax3x) & (ax2x) & (ax1x) & (!shiftx0x) & (shiftx1x)) + ((!ax4x) & (!ax3x) & (ax2x) & (ax1x) & (shiftx0x) & (shiftx1x)) + ((!ax4x) & (ax3x) & (!ax2x) & (!ax1x) & (shiftx0x) & (!shiftx1x)) + ((!ax4x) & (ax3x) & (!ax2x) & (ax1x) & (shiftx0x) & (!shiftx1x)) + ((!ax4x) & (ax3x) & (!ax2x) & (ax1x) & (shiftx0x) & (shiftx1x)) + ((!ax4x) & (ax3x) & (ax2x) & (!ax1x) & (!shiftx0x) & (shiftx1x)) + ((!ax4x) & (ax3x) & (ax2x) & (!ax1x) & (shiftx0x) & (!shiftx1x)) + ((!ax4x) & (ax3x) & (ax2x) & (ax1x) & (!shiftx0x) & (shiftx1x)) + ((!ax4x) & (ax3x) & (ax2x) & (ax1x) & (shiftx0x) & (!shiftx1x)) + ((!ax4x) & (ax3x) & (ax2x) & (ax1x) & (shiftx0x) & (shiftx1x)) + ((ax4x) & (!ax3x) & (!ax2x) & (!ax1x) & (!shiftx0x) & (!shiftx1x)) + ((ax4x) & (!ax3x) & (!ax2x) & (ax1x) & (!shiftx0x) & (!shiftx1x)) + ((ax4x) & (!ax3x) & (!ax2x) & (ax1x) & (shiftx0x) & (shiftx1x)) + ((ax4x) & (!ax3x) & (ax2x) & (!ax1x) & (!shiftx0x) & (!shiftx1x)) + ((ax4x) & (!ax3x) & (ax2x) & (!ax1x) & (!shiftx0x) & (shiftx1x)) + ((ax4x) & (!ax3x) & (ax2x) & (ax1x) & (!shiftx0x) & (!shiftx1x)) + ((ax4x) & (!ax3x) & (ax2x) & (ax1x) & (!shiftx0x) & (shiftx1x)) + ((ax4x) & (!ax3x) & (ax2x) & (ax1x) & (shiftx0x) & (shiftx1x)) + ((ax4x) & (ax3x) & (!ax2x) & (!ax1x) & (!shiftx0x) & (!shiftx1x)) + ((ax4x) & (ax3x) & (!ax2x) & (!ax1x) & (shiftx0x) & (!shiftx1x)) + ((ax4x) & (ax3x) & (!ax2x) & (ax1x) & (!shiftx0x) & (!shiftx1x)) + ((ax4x) & (ax3x) & (!ax2x) & (ax1x) & (shiftx0x) & (!shiftx1x)) + ((ax4x) & (ax3x) & (!ax2x) & (ax1x) & (shiftx0x) & (shiftx1x)) + ((ax4x) & (ax3x) & (ax2x) & (!ax1x) & (!shiftx0x) & (!shiftx1x)) + ((ax4x) & (ax3x) & (ax2x) & (!ax1x) & (!shiftx0x) & (shiftx1x)) + ((ax4x) & (ax3x) & (ax2x) & (!ax1x) & (shiftx0x) & (!shiftx1x)) + ((ax4x) & (ax3x) & (ax2x) & (ax1x) & (!shiftx0x) & (!shiftx1x)) + ((ax4x) & (ax3x) & (ax2x) & (ax1x) & (!shiftx0x) & (shiftx1x)) + ((ax4x) & (ax3x) & (ax2x) & (ax1x) & (shiftx0x) & (!shiftx1x)) + ((ax4x) & (ax3x) & (ax2x) & (ax1x) & (shiftx0x) & (shiftx1x)));
	assign g4 = (((!ax8x) & (!ax7x) & (!ax6x) & (ax5x) & (shiftx0x) & (shiftx1x)) + ((!ax8x) & (!ax7x) & (ax6x) & (!ax5x) & (!shiftx0x) & (shiftx1x)) + ((!ax8x) & (!ax7x) & (ax6x) & (ax5x) & (!shiftx0x) & (shiftx1x)) + ((!ax8x) & (!ax7x) & (ax6x) & (ax5x) & (shiftx0x) & (shiftx1x)) + ((!ax8x) & (ax7x) & (!ax6x) & (!ax5x) & (shiftx0x) & (!shiftx1x)) + ((!ax8x) & (ax7x) & (!ax6x) & (ax5x) & (shiftx0x) & (!shiftx1x)) + ((!ax8x) & (ax7x) & (!ax6x) & (ax5x) & (shiftx0x) & (shiftx1x)) + ((!ax8x) & (ax7x) & (ax6x) & (!ax5x) & (!shiftx0x) & (shiftx1x)) + ((!ax8x) & (ax7x) & (ax6x) & (!ax5x) & (shiftx0x) & (!shiftx1x)) + ((!ax8x) & (ax7x) & (ax6x) & (ax5x) & (!shiftx0x) & (shiftx1x)) + ((!ax8x) & (ax7x) & (ax6x) & (ax5x) & (shiftx0x) & (!shiftx1x)) + ((!ax8x) & (ax7x) & (ax6x) & (ax5x) & (shiftx0x) & (shiftx1x)) + ((ax8x) & (!ax7x) & (!ax6x) & (!ax5x) & (!shiftx0x) & (!shiftx1x)) + ((ax8x) & (!ax7x) & (!ax6x) & (ax5x) & (!shiftx0x) & (!shiftx1x)) + ((ax8x) & (!ax7x) & (!ax6x) & (ax5x) & (shiftx0x) & (shiftx1x)) + ((ax8x) & (!ax7x) & (ax6x) & (!ax5x) & (!shiftx0x) & (!shiftx1x)) + ((ax8x) & (!ax7x) & (ax6x) & (!ax5x) & (!shiftx0x) & (shiftx1x)) + ((ax8x) & (!ax7x) & (ax6x) & (ax5x) & (!shiftx0x) & (!shiftx1x)) + ((ax8x) & (!ax7x) & (ax6x) & (ax5x) & (!shiftx0x) & (shiftx1x)) + ((ax8x) & (!ax7x) & (ax6x) & (ax5x) & (shiftx0x) & (shiftx1x)) + ((ax8x) & (ax7x) & (!ax6x) & (!ax5x) & (!shiftx0x) & (!shiftx1x)) + ((ax8x) & (ax7x) & (!ax6x) & (!ax5x) & (shiftx0x) & (!shiftx1x)) + ((ax8x) & (ax7x) & (!ax6x) & (ax5x) & (!shiftx0x) & (!shiftx1x)) + ((ax8x) & (ax7x) & (!ax6x) & (ax5x) & (shiftx0x) & (!shiftx1x)) + ((ax8x) & (ax7x) & (!ax6x) & (ax5x) & (shiftx0x) & (shiftx1x)) + ((ax8x) & (ax7x) & (ax6x) & (!ax5x) & (!shiftx0x) & (!shiftx1x)) + ((ax8x) & (ax7x) & (ax6x) & (!ax5x) & (!shiftx0x) & (shiftx1x)) + ((ax8x) & (ax7x) & (ax6x) & (!ax5x) & (shiftx0x) & (!shiftx1x)) + ((ax8x) & (ax7x) & (ax6x) & (ax5x) & (!shiftx0x) & (!shiftx1x)) + ((ax8x) & (ax7x) & (ax6x) & (ax5x) & (!shiftx0x) & (shiftx1x)) + ((ax8x) & (ax7x) & (ax6x) & (ax5x) & (shiftx0x) & (!shiftx1x)) + ((ax8x) & (ax7x) & (ax6x) & (ax5x) & (shiftx0x) & (shiftx1x)));
	assign g5 = (((!shiftx2x) & (!shiftx3x) & (g1) & (!g2) & (!g3) & (!g4)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (!g2) & (!g3) & (g4)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (!g2) & (g3) & (!g4)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (!g2) & (g3) & (g4)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (g2) & (!g3) & (!g4)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (g2) & (!g3) & (g4)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (g2) & (g3) & (!g4)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (g2) & (g3) & (g4)) + ((!shiftx2x) & (shiftx3x) & (!g1) & (!g2) & (!g3) & (g4)) + ((!shiftx2x) & (shiftx3x) & (!g1) & (!g2) & (g3) & (g4)) + ((!shiftx2x) & (shiftx3x) & (!g1) & (g2) & (!g3) & (g4)) + ((!shiftx2x) & (shiftx3x) & (!g1) & (g2) & (g3) & (g4)) + ((!shiftx2x) & (shiftx3x) & (g1) & (!g2) & (!g3) & (g4)) + ((!shiftx2x) & (shiftx3x) & (g1) & (!g2) & (g3) & (g4)) + ((!shiftx2x) & (shiftx3x) & (g1) & (g2) & (!g3) & (g4)) + ((!shiftx2x) & (shiftx3x) & (g1) & (g2) & (g3) & (g4)) + ((shiftx2x) & (!shiftx3x) & (!g1) & (g2) & (!g3) & (!g4)) + ((shiftx2x) & (!shiftx3x) & (!g1) & (g2) & (!g3) & (g4)) + ((shiftx2x) & (!shiftx3x) & (!g1) & (g2) & (g3) & (!g4)) + ((shiftx2x) & (!shiftx3x) & (!g1) & (g2) & (g3) & (g4)) + ((shiftx2x) & (!shiftx3x) & (g1) & (g2) & (!g3) & (!g4)) + ((shiftx2x) & (!shiftx3x) & (g1) & (g2) & (!g3) & (g4)) + ((shiftx2x) & (!shiftx3x) & (g1) & (g2) & (g3) & (!g4)) + ((shiftx2x) & (!shiftx3x) & (g1) & (g2) & (g3) & (g4)) + ((shiftx2x) & (shiftx3x) & (!g1) & (!g2) & (g3) & (!g4)) + ((shiftx2x) & (shiftx3x) & (!g1) & (!g2) & (g3) & (g4)) + ((shiftx2x) & (shiftx3x) & (!g1) & (g2) & (g3) & (!g4)) + ((shiftx2x) & (shiftx3x) & (!g1) & (g2) & (g3) & (g4)) + ((shiftx2x) & (shiftx3x) & (g1) & (!g2) & (g3) & (!g4)) + ((shiftx2x) & (shiftx3x) & (g1) & (!g2) & (g3) & (g4)) + ((shiftx2x) & (shiftx3x) & (g1) & (g2) & (g3) & (!g4)) + ((shiftx2x) & (shiftx3x) & (g1) & (g2) & (g3) & (g4)));
	assign g6 = (((!ax32x) & (!ax31x) & (!ax30x) & (ax29x) & (shiftx0x) & (shiftx1x)) + ((!ax32x) & (!ax31x) & (ax30x) & (!ax29x) & (!shiftx0x) & (shiftx1x)) + ((!ax32x) & (!ax31x) & (ax30x) & (ax29x) & (!shiftx0x) & (shiftx1x)) + ((!ax32x) & (!ax31x) & (ax30x) & (ax29x) & (shiftx0x) & (shiftx1x)) + ((!ax32x) & (ax31x) & (!ax30x) & (!ax29x) & (shiftx0x) & (!shiftx1x)) + ((!ax32x) & (ax31x) & (!ax30x) & (ax29x) & (shiftx0x) & (!shiftx1x)) + ((!ax32x) & (ax31x) & (!ax30x) & (ax29x) & (shiftx0x) & (shiftx1x)) + ((!ax32x) & (ax31x) & (ax30x) & (!ax29x) & (!shiftx0x) & (shiftx1x)) + ((!ax32x) & (ax31x) & (ax30x) & (!ax29x) & (shiftx0x) & (!shiftx1x)) + ((!ax32x) & (ax31x) & (ax30x) & (ax29x) & (!shiftx0x) & (shiftx1x)) + ((!ax32x) & (ax31x) & (ax30x) & (ax29x) & (shiftx0x) & (!shiftx1x)) + ((!ax32x) & (ax31x) & (ax30x) & (ax29x) & (shiftx0x) & (shiftx1x)) + ((ax32x) & (!ax31x) & (!ax30x) & (!ax29x) & (!shiftx0x) & (!shiftx1x)) + ((ax32x) & (!ax31x) & (!ax30x) & (ax29x) & (!shiftx0x) & (!shiftx1x)) + ((ax32x) & (!ax31x) & (!ax30x) & (ax29x) & (shiftx0x) & (shiftx1x)) + ((ax32x) & (!ax31x) & (ax30x) & (!ax29x) & (!shiftx0x) & (!shiftx1x)) + ((ax32x) & (!ax31x) & (ax30x) & (!ax29x) & (!shiftx0x) & (shiftx1x)) + ((ax32x) & (!ax31x) & (ax30x) & (ax29x) & (!shiftx0x) & (!shiftx1x)) + ((ax32x) & (!ax31x) & (ax30x) & (ax29x) & (!shiftx0x) & (shiftx1x)) + ((ax32x) & (!ax31x) & (ax30x) & (ax29x) & (shiftx0x) & (shiftx1x)) + ((ax32x) & (ax31x) & (!ax30x) & (!ax29x) & (!shiftx0x) & (!shiftx1x)) + ((ax32x) & (ax31x) & (!ax30x) & (!ax29x) & (shiftx0x) & (!shiftx1x)) + ((ax32x) & (ax31x) & (!ax30x) & (ax29x) & (!shiftx0x) & (!shiftx1x)) + ((ax32x) & (ax31x) & (!ax30x) & (ax29x) & (shiftx0x) & (!shiftx1x)) + ((ax32x) & (ax31x) & (!ax30x) & (ax29x) & (shiftx0x) & (shiftx1x)) + ((ax32x) & (ax31x) & (ax30x) & (!ax29x) & (!shiftx0x) & (!shiftx1x)) + ((ax32x) & (ax31x) & (ax30x) & (!ax29x) & (!shiftx0x) & (shiftx1x)) + ((ax32x) & (ax31x) & (ax30x) & (!ax29x) & (shiftx0x) & (!shiftx1x)) + ((ax32x) & (ax31x) & (ax30x) & (ax29x) & (!shiftx0x) & (!shiftx1x)) + ((ax32x) & (ax31x) & (ax30x) & (ax29x) & (!shiftx0x) & (shiftx1x)) + ((ax32x) & (ax31x) & (ax30x) & (ax29x) & (shiftx0x) & (!shiftx1x)) + ((ax32x) & (ax31x) & (ax30x) & (ax29x) & (shiftx0x) & (shiftx1x)));
	assign g7 = (((!ax28x) & (!ax27x) & (!ax26x) & (ax25x) & (shiftx0x) & (shiftx1x)) + ((!ax28x) & (!ax27x) & (ax26x) & (!ax25x) & (!shiftx0x) & (shiftx1x)) + ((!ax28x) & (!ax27x) & (ax26x) & (ax25x) & (!shiftx0x) & (shiftx1x)) + ((!ax28x) & (!ax27x) & (ax26x) & (ax25x) & (shiftx0x) & (shiftx1x)) + ((!ax28x) & (ax27x) & (!ax26x) & (!ax25x) & (shiftx0x) & (!shiftx1x)) + ((!ax28x) & (ax27x) & (!ax26x) & (ax25x) & (shiftx0x) & (!shiftx1x)) + ((!ax28x) & (ax27x) & (!ax26x) & (ax25x) & (shiftx0x) & (shiftx1x)) + ((!ax28x) & (ax27x) & (ax26x) & (!ax25x) & (!shiftx0x) & (shiftx1x)) + ((!ax28x) & (ax27x) & (ax26x) & (!ax25x) & (shiftx0x) & (!shiftx1x)) + ((!ax28x) & (ax27x) & (ax26x) & (ax25x) & (!shiftx0x) & (shiftx1x)) + ((!ax28x) & (ax27x) & (ax26x) & (ax25x) & (shiftx0x) & (!shiftx1x)) + ((!ax28x) & (ax27x) & (ax26x) & (ax25x) & (shiftx0x) & (shiftx1x)) + ((ax28x) & (!ax27x) & (!ax26x) & (!ax25x) & (!shiftx0x) & (!shiftx1x)) + ((ax28x) & (!ax27x) & (!ax26x) & (ax25x) & (!shiftx0x) & (!shiftx1x)) + ((ax28x) & (!ax27x) & (!ax26x) & (ax25x) & (shiftx0x) & (shiftx1x)) + ((ax28x) & (!ax27x) & (ax26x) & (!ax25x) & (!shiftx0x) & (!shiftx1x)) + ((ax28x) & (!ax27x) & (ax26x) & (!ax25x) & (!shiftx0x) & (shiftx1x)) + ((ax28x) & (!ax27x) & (ax26x) & (ax25x) & (!shiftx0x) & (!shiftx1x)) + ((ax28x) & (!ax27x) & (ax26x) & (ax25x) & (!shiftx0x) & (shiftx1x)) + ((ax28x) & (!ax27x) & (ax26x) & (ax25x) & (shiftx0x) & (shiftx1x)) + ((ax28x) & (ax27x) & (!ax26x) & (!ax25x) & (!shiftx0x) & (!shiftx1x)) + ((ax28x) & (ax27x) & (!ax26x) & (!ax25x) & (shiftx0x) & (!shiftx1x)) + ((ax28x) & (ax27x) & (!ax26x) & (ax25x) & (!shiftx0x) & (!shiftx1x)) + ((ax28x) & (ax27x) & (!ax26x) & (ax25x) & (shiftx0x) & (!shiftx1x)) + ((ax28x) & (ax27x) & (!ax26x) & (ax25x) & (shiftx0x) & (shiftx1x)) + ((ax28x) & (ax27x) & (ax26x) & (!ax25x) & (!shiftx0x) & (!shiftx1x)) + ((ax28x) & (ax27x) & (ax26x) & (!ax25x) & (!shiftx0x) & (shiftx1x)) + ((ax28x) & (ax27x) & (ax26x) & (!ax25x) & (shiftx0x) & (!shiftx1x)) + ((ax28x) & (ax27x) & (ax26x) & (ax25x) & (!shiftx0x) & (!shiftx1x)) + ((ax28x) & (ax27x) & (ax26x) & (ax25x) & (!shiftx0x) & (shiftx1x)) + ((ax28x) & (ax27x) & (ax26x) & (ax25x) & (shiftx0x) & (!shiftx1x)) + ((ax28x) & (ax27x) & (ax26x) & (ax25x) & (shiftx0x) & (shiftx1x)));
	assign g8 = (((!ax20x) & (!ax19x) & (!ax18x) & (ax17x) & (shiftx0x) & (shiftx1x)) + ((!ax20x) & (!ax19x) & (ax18x) & (!ax17x) & (!shiftx0x) & (shiftx1x)) + ((!ax20x) & (!ax19x) & (ax18x) & (ax17x) & (!shiftx0x) & (shiftx1x)) + ((!ax20x) & (!ax19x) & (ax18x) & (ax17x) & (shiftx0x) & (shiftx1x)) + ((!ax20x) & (ax19x) & (!ax18x) & (!ax17x) & (shiftx0x) & (!shiftx1x)) + ((!ax20x) & (ax19x) & (!ax18x) & (ax17x) & (shiftx0x) & (!shiftx1x)) + ((!ax20x) & (ax19x) & (!ax18x) & (ax17x) & (shiftx0x) & (shiftx1x)) + ((!ax20x) & (ax19x) & (ax18x) & (!ax17x) & (!shiftx0x) & (shiftx1x)) + ((!ax20x) & (ax19x) & (ax18x) & (!ax17x) & (shiftx0x) & (!shiftx1x)) + ((!ax20x) & (ax19x) & (ax18x) & (ax17x) & (!shiftx0x) & (shiftx1x)) + ((!ax20x) & (ax19x) & (ax18x) & (ax17x) & (shiftx0x) & (!shiftx1x)) + ((!ax20x) & (ax19x) & (ax18x) & (ax17x) & (shiftx0x) & (shiftx1x)) + ((ax20x) & (!ax19x) & (!ax18x) & (!ax17x) & (!shiftx0x) & (!shiftx1x)) + ((ax20x) & (!ax19x) & (!ax18x) & (ax17x) & (!shiftx0x) & (!shiftx1x)) + ((ax20x) & (!ax19x) & (!ax18x) & (ax17x) & (shiftx0x) & (shiftx1x)) + ((ax20x) & (!ax19x) & (ax18x) & (!ax17x) & (!shiftx0x) & (!shiftx1x)) + ((ax20x) & (!ax19x) & (ax18x) & (!ax17x) & (!shiftx0x) & (shiftx1x)) + ((ax20x) & (!ax19x) & (ax18x) & (ax17x) & (!shiftx0x) & (!shiftx1x)) + ((ax20x) & (!ax19x) & (ax18x) & (ax17x) & (!shiftx0x) & (shiftx1x)) + ((ax20x) & (!ax19x) & (ax18x) & (ax17x) & (shiftx0x) & (shiftx1x)) + ((ax20x) & (ax19x) & (!ax18x) & (!ax17x) & (!shiftx0x) & (!shiftx1x)) + ((ax20x) & (ax19x) & (!ax18x) & (!ax17x) & (shiftx0x) & (!shiftx1x)) + ((ax20x) & (ax19x) & (!ax18x) & (ax17x) & (!shiftx0x) & (!shiftx1x)) + ((ax20x) & (ax19x) & (!ax18x) & (ax17x) & (shiftx0x) & (!shiftx1x)) + ((ax20x) & (ax19x) & (!ax18x) & (ax17x) & (shiftx0x) & (shiftx1x)) + ((ax20x) & (ax19x) & (ax18x) & (!ax17x) & (!shiftx0x) & (!shiftx1x)) + ((ax20x) & (ax19x) & (ax18x) & (!ax17x) & (!shiftx0x) & (shiftx1x)) + ((ax20x) & (ax19x) & (ax18x) & (!ax17x) & (shiftx0x) & (!shiftx1x)) + ((ax20x) & (ax19x) & (ax18x) & (ax17x) & (!shiftx0x) & (!shiftx1x)) + ((ax20x) & (ax19x) & (ax18x) & (ax17x) & (!shiftx0x) & (shiftx1x)) + ((ax20x) & (ax19x) & (ax18x) & (ax17x) & (shiftx0x) & (!shiftx1x)) + ((ax20x) & (ax19x) & (ax18x) & (ax17x) & (shiftx0x) & (shiftx1x)));
	assign g9 = (((!ax24x) & (!ax23x) & (!ax22x) & (ax21x) & (shiftx0x) & (shiftx1x)) + ((!ax24x) & (!ax23x) & (ax22x) & (!ax21x) & (!shiftx0x) & (shiftx1x)) + ((!ax24x) & (!ax23x) & (ax22x) & (ax21x) & (!shiftx0x) & (shiftx1x)) + ((!ax24x) & (!ax23x) & (ax22x) & (ax21x) & (shiftx0x) & (shiftx1x)) + ((!ax24x) & (ax23x) & (!ax22x) & (!ax21x) & (shiftx0x) & (!shiftx1x)) + ((!ax24x) & (ax23x) & (!ax22x) & (ax21x) & (shiftx0x) & (!shiftx1x)) + ((!ax24x) & (ax23x) & (!ax22x) & (ax21x) & (shiftx0x) & (shiftx1x)) + ((!ax24x) & (ax23x) & (ax22x) & (!ax21x) & (!shiftx0x) & (shiftx1x)) + ((!ax24x) & (ax23x) & (ax22x) & (!ax21x) & (shiftx0x) & (!shiftx1x)) + ((!ax24x) & (ax23x) & (ax22x) & (ax21x) & (!shiftx0x) & (shiftx1x)) + ((!ax24x) & (ax23x) & (ax22x) & (ax21x) & (shiftx0x) & (!shiftx1x)) + ((!ax24x) & (ax23x) & (ax22x) & (ax21x) & (shiftx0x) & (shiftx1x)) + ((ax24x) & (!ax23x) & (!ax22x) & (!ax21x) & (!shiftx0x) & (!shiftx1x)) + ((ax24x) & (!ax23x) & (!ax22x) & (ax21x) & (!shiftx0x) & (!shiftx1x)) + ((ax24x) & (!ax23x) & (!ax22x) & (ax21x) & (shiftx0x) & (shiftx1x)) + ((ax24x) & (!ax23x) & (ax22x) & (!ax21x) & (!shiftx0x) & (!shiftx1x)) + ((ax24x) & (!ax23x) & (ax22x) & (!ax21x) & (!shiftx0x) & (shiftx1x)) + ((ax24x) & (!ax23x) & (ax22x) & (ax21x) & (!shiftx0x) & (!shiftx1x)) + ((ax24x) & (!ax23x) & (ax22x) & (ax21x) & (!shiftx0x) & (shiftx1x)) + ((ax24x) & (!ax23x) & (ax22x) & (ax21x) & (shiftx0x) & (shiftx1x)) + ((ax24x) & (ax23x) & (!ax22x) & (!ax21x) & (!shiftx0x) & (!shiftx1x)) + ((ax24x) & (ax23x) & (!ax22x) & (!ax21x) & (shiftx0x) & (!shiftx1x)) + ((ax24x) & (ax23x) & (!ax22x) & (ax21x) & (!shiftx0x) & (!shiftx1x)) + ((ax24x) & (ax23x) & (!ax22x) & (ax21x) & (shiftx0x) & (!shiftx1x)) + ((ax24x) & (ax23x) & (!ax22x) & (ax21x) & (shiftx0x) & (shiftx1x)) + ((ax24x) & (ax23x) & (ax22x) & (!ax21x) & (!shiftx0x) & (!shiftx1x)) + ((ax24x) & (ax23x) & (ax22x) & (!ax21x) & (!shiftx0x) & (shiftx1x)) + ((ax24x) & (ax23x) & (ax22x) & (!ax21x) & (shiftx0x) & (!shiftx1x)) + ((ax24x) & (ax23x) & (ax22x) & (ax21x) & (!shiftx0x) & (!shiftx1x)) + ((ax24x) & (ax23x) & (ax22x) & (ax21x) & (!shiftx0x) & (shiftx1x)) + ((ax24x) & (ax23x) & (ax22x) & (ax21x) & (shiftx0x) & (!shiftx1x)) + ((ax24x) & (ax23x) & (ax22x) & (ax21x) & (shiftx0x) & (shiftx1x)));
	assign g10 = (((!shiftx2x) & (!shiftx3x) & (g6) & (!g7) & (!g8) & (!g9)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (!g7) & (!g8) & (g9)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (!g7) & (g8) & (!g9)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (!g7) & (g8) & (g9)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (g7) & (!g8) & (!g9)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (g7) & (!g8) & (g9)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (g7) & (g8) & (!g9)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (g7) & (g8) & (g9)) + ((!shiftx2x) & (shiftx3x) & (!g6) & (!g7) & (!g8) & (g9)) + ((!shiftx2x) & (shiftx3x) & (!g6) & (!g7) & (g8) & (g9)) + ((!shiftx2x) & (shiftx3x) & (!g6) & (g7) & (!g8) & (g9)) + ((!shiftx2x) & (shiftx3x) & (!g6) & (g7) & (g8) & (g9)) + ((!shiftx2x) & (shiftx3x) & (g6) & (!g7) & (!g8) & (g9)) + ((!shiftx2x) & (shiftx3x) & (g6) & (!g7) & (g8) & (g9)) + ((!shiftx2x) & (shiftx3x) & (g6) & (g7) & (!g8) & (g9)) + ((!shiftx2x) & (shiftx3x) & (g6) & (g7) & (g8) & (g9)) + ((shiftx2x) & (!shiftx3x) & (!g6) & (g7) & (!g8) & (!g9)) + ((shiftx2x) & (!shiftx3x) & (!g6) & (g7) & (!g8) & (g9)) + ((shiftx2x) & (!shiftx3x) & (!g6) & (g7) & (g8) & (!g9)) + ((shiftx2x) & (!shiftx3x) & (!g6) & (g7) & (g8) & (g9)) + ((shiftx2x) & (!shiftx3x) & (g6) & (g7) & (!g8) & (!g9)) + ((shiftx2x) & (!shiftx3x) & (g6) & (g7) & (!g8) & (g9)) + ((shiftx2x) & (!shiftx3x) & (g6) & (g7) & (g8) & (!g9)) + ((shiftx2x) & (!shiftx3x) & (g6) & (g7) & (g8) & (g9)) + ((shiftx2x) & (shiftx3x) & (!g6) & (!g7) & (g8) & (!g9)) + ((shiftx2x) & (shiftx3x) & (!g6) & (!g7) & (g8) & (g9)) + ((shiftx2x) & (shiftx3x) & (!g6) & (g7) & (g8) & (!g9)) + ((shiftx2x) & (shiftx3x) & (!g6) & (g7) & (g8) & (g9)) + ((shiftx2x) & (shiftx3x) & (g6) & (!g7) & (g8) & (!g9)) + ((shiftx2x) & (shiftx3x) & (g6) & (!g7) & (g8) & (g9)) + ((shiftx2x) & (shiftx3x) & (g6) & (g7) & (g8) & (!g9)) + ((shiftx2x) & (shiftx3x) & (g6) & (g7) & (g8) & (g9)));
	assign g11 = (((!ax64x) & (!ax63x) & (!ax62x) & (ax61x) & (shiftx0x) & (shiftx1x)) + ((!ax64x) & (!ax63x) & (ax62x) & (!ax61x) & (!shiftx0x) & (shiftx1x)) + ((!ax64x) & (!ax63x) & (ax62x) & (ax61x) & (!shiftx0x) & (shiftx1x)) + ((!ax64x) & (!ax63x) & (ax62x) & (ax61x) & (shiftx0x) & (shiftx1x)) + ((!ax64x) & (ax63x) & (!ax62x) & (!ax61x) & (shiftx0x) & (!shiftx1x)) + ((!ax64x) & (ax63x) & (!ax62x) & (ax61x) & (shiftx0x) & (!shiftx1x)) + ((!ax64x) & (ax63x) & (!ax62x) & (ax61x) & (shiftx0x) & (shiftx1x)) + ((!ax64x) & (ax63x) & (ax62x) & (!ax61x) & (!shiftx0x) & (shiftx1x)) + ((!ax64x) & (ax63x) & (ax62x) & (!ax61x) & (shiftx0x) & (!shiftx1x)) + ((!ax64x) & (ax63x) & (ax62x) & (ax61x) & (!shiftx0x) & (shiftx1x)) + ((!ax64x) & (ax63x) & (ax62x) & (ax61x) & (shiftx0x) & (!shiftx1x)) + ((!ax64x) & (ax63x) & (ax62x) & (ax61x) & (shiftx0x) & (shiftx1x)) + ((ax64x) & (!ax63x) & (!ax62x) & (!ax61x) & (!shiftx0x) & (!shiftx1x)) + ((ax64x) & (!ax63x) & (!ax62x) & (ax61x) & (!shiftx0x) & (!shiftx1x)) + ((ax64x) & (!ax63x) & (!ax62x) & (ax61x) & (shiftx0x) & (shiftx1x)) + ((ax64x) & (!ax63x) & (ax62x) & (!ax61x) & (!shiftx0x) & (!shiftx1x)) + ((ax64x) & (!ax63x) & (ax62x) & (!ax61x) & (!shiftx0x) & (shiftx1x)) + ((ax64x) & (!ax63x) & (ax62x) & (ax61x) & (!shiftx0x) & (!shiftx1x)) + ((ax64x) & (!ax63x) & (ax62x) & (ax61x) & (!shiftx0x) & (shiftx1x)) + ((ax64x) & (!ax63x) & (ax62x) & (ax61x) & (shiftx0x) & (shiftx1x)) + ((ax64x) & (ax63x) & (!ax62x) & (!ax61x) & (!shiftx0x) & (!shiftx1x)) + ((ax64x) & (ax63x) & (!ax62x) & (!ax61x) & (shiftx0x) & (!shiftx1x)) + ((ax64x) & (ax63x) & (!ax62x) & (ax61x) & (!shiftx0x) & (!shiftx1x)) + ((ax64x) & (ax63x) & (!ax62x) & (ax61x) & (shiftx0x) & (!shiftx1x)) + ((ax64x) & (ax63x) & (!ax62x) & (ax61x) & (shiftx0x) & (shiftx1x)) + ((ax64x) & (ax63x) & (ax62x) & (!ax61x) & (!shiftx0x) & (!shiftx1x)) + ((ax64x) & (ax63x) & (ax62x) & (!ax61x) & (!shiftx0x) & (shiftx1x)) + ((ax64x) & (ax63x) & (ax62x) & (!ax61x) & (shiftx0x) & (!shiftx1x)) + ((ax64x) & (ax63x) & (ax62x) & (ax61x) & (!shiftx0x) & (!shiftx1x)) + ((ax64x) & (ax63x) & (ax62x) & (ax61x) & (!shiftx0x) & (shiftx1x)) + ((ax64x) & (ax63x) & (ax62x) & (ax61x) & (shiftx0x) & (!shiftx1x)) + ((ax64x) & (ax63x) & (ax62x) & (ax61x) & (shiftx0x) & (shiftx1x)));
	assign g12 = (((!ax60x) & (!ax59x) & (!ax58x) & (ax57x) & (shiftx0x) & (shiftx1x)) + ((!ax60x) & (!ax59x) & (ax58x) & (!ax57x) & (!shiftx0x) & (shiftx1x)) + ((!ax60x) & (!ax59x) & (ax58x) & (ax57x) & (!shiftx0x) & (shiftx1x)) + ((!ax60x) & (!ax59x) & (ax58x) & (ax57x) & (shiftx0x) & (shiftx1x)) + ((!ax60x) & (ax59x) & (!ax58x) & (!ax57x) & (shiftx0x) & (!shiftx1x)) + ((!ax60x) & (ax59x) & (!ax58x) & (ax57x) & (shiftx0x) & (!shiftx1x)) + ((!ax60x) & (ax59x) & (!ax58x) & (ax57x) & (shiftx0x) & (shiftx1x)) + ((!ax60x) & (ax59x) & (ax58x) & (!ax57x) & (!shiftx0x) & (shiftx1x)) + ((!ax60x) & (ax59x) & (ax58x) & (!ax57x) & (shiftx0x) & (!shiftx1x)) + ((!ax60x) & (ax59x) & (ax58x) & (ax57x) & (!shiftx0x) & (shiftx1x)) + ((!ax60x) & (ax59x) & (ax58x) & (ax57x) & (shiftx0x) & (!shiftx1x)) + ((!ax60x) & (ax59x) & (ax58x) & (ax57x) & (shiftx0x) & (shiftx1x)) + ((ax60x) & (!ax59x) & (!ax58x) & (!ax57x) & (!shiftx0x) & (!shiftx1x)) + ((ax60x) & (!ax59x) & (!ax58x) & (ax57x) & (!shiftx0x) & (!shiftx1x)) + ((ax60x) & (!ax59x) & (!ax58x) & (ax57x) & (shiftx0x) & (shiftx1x)) + ((ax60x) & (!ax59x) & (ax58x) & (!ax57x) & (!shiftx0x) & (!shiftx1x)) + ((ax60x) & (!ax59x) & (ax58x) & (!ax57x) & (!shiftx0x) & (shiftx1x)) + ((ax60x) & (!ax59x) & (ax58x) & (ax57x) & (!shiftx0x) & (!shiftx1x)) + ((ax60x) & (!ax59x) & (ax58x) & (ax57x) & (!shiftx0x) & (shiftx1x)) + ((ax60x) & (!ax59x) & (ax58x) & (ax57x) & (shiftx0x) & (shiftx1x)) + ((ax60x) & (ax59x) & (!ax58x) & (!ax57x) & (!shiftx0x) & (!shiftx1x)) + ((ax60x) & (ax59x) & (!ax58x) & (!ax57x) & (shiftx0x) & (!shiftx1x)) + ((ax60x) & (ax59x) & (!ax58x) & (ax57x) & (!shiftx0x) & (!shiftx1x)) + ((ax60x) & (ax59x) & (!ax58x) & (ax57x) & (shiftx0x) & (!shiftx1x)) + ((ax60x) & (ax59x) & (!ax58x) & (ax57x) & (shiftx0x) & (shiftx1x)) + ((ax60x) & (ax59x) & (ax58x) & (!ax57x) & (!shiftx0x) & (!shiftx1x)) + ((ax60x) & (ax59x) & (ax58x) & (!ax57x) & (!shiftx0x) & (shiftx1x)) + ((ax60x) & (ax59x) & (ax58x) & (!ax57x) & (shiftx0x) & (!shiftx1x)) + ((ax60x) & (ax59x) & (ax58x) & (ax57x) & (!shiftx0x) & (!shiftx1x)) + ((ax60x) & (ax59x) & (ax58x) & (ax57x) & (!shiftx0x) & (shiftx1x)) + ((ax60x) & (ax59x) & (ax58x) & (ax57x) & (shiftx0x) & (!shiftx1x)) + ((ax60x) & (ax59x) & (ax58x) & (ax57x) & (shiftx0x) & (shiftx1x)));
	assign g13 = (((!ax52x) & (!ax51x) & (!ax50x) & (ax49x) & (shiftx0x) & (shiftx1x)) + ((!ax52x) & (!ax51x) & (ax50x) & (!ax49x) & (!shiftx0x) & (shiftx1x)) + ((!ax52x) & (!ax51x) & (ax50x) & (ax49x) & (!shiftx0x) & (shiftx1x)) + ((!ax52x) & (!ax51x) & (ax50x) & (ax49x) & (shiftx0x) & (shiftx1x)) + ((!ax52x) & (ax51x) & (!ax50x) & (!ax49x) & (shiftx0x) & (!shiftx1x)) + ((!ax52x) & (ax51x) & (!ax50x) & (ax49x) & (shiftx0x) & (!shiftx1x)) + ((!ax52x) & (ax51x) & (!ax50x) & (ax49x) & (shiftx0x) & (shiftx1x)) + ((!ax52x) & (ax51x) & (ax50x) & (!ax49x) & (!shiftx0x) & (shiftx1x)) + ((!ax52x) & (ax51x) & (ax50x) & (!ax49x) & (shiftx0x) & (!shiftx1x)) + ((!ax52x) & (ax51x) & (ax50x) & (ax49x) & (!shiftx0x) & (shiftx1x)) + ((!ax52x) & (ax51x) & (ax50x) & (ax49x) & (shiftx0x) & (!shiftx1x)) + ((!ax52x) & (ax51x) & (ax50x) & (ax49x) & (shiftx0x) & (shiftx1x)) + ((ax52x) & (!ax51x) & (!ax50x) & (!ax49x) & (!shiftx0x) & (!shiftx1x)) + ((ax52x) & (!ax51x) & (!ax50x) & (ax49x) & (!shiftx0x) & (!shiftx1x)) + ((ax52x) & (!ax51x) & (!ax50x) & (ax49x) & (shiftx0x) & (shiftx1x)) + ((ax52x) & (!ax51x) & (ax50x) & (!ax49x) & (!shiftx0x) & (!shiftx1x)) + ((ax52x) & (!ax51x) & (ax50x) & (!ax49x) & (!shiftx0x) & (shiftx1x)) + ((ax52x) & (!ax51x) & (ax50x) & (ax49x) & (!shiftx0x) & (!shiftx1x)) + ((ax52x) & (!ax51x) & (ax50x) & (ax49x) & (!shiftx0x) & (shiftx1x)) + ((ax52x) & (!ax51x) & (ax50x) & (ax49x) & (shiftx0x) & (shiftx1x)) + ((ax52x) & (ax51x) & (!ax50x) & (!ax49x) & (!shiftx0x) & (!shiftx1x)) + ((ax52x) & (ax51x) & (!ax50x) & (!ax49x) & (shiftx0x) & (!shiftx1x)) + ((ax52x) & (ax51x) & (!ax50x) & (ax49x) & (!shiftx0x) & (!shiftx1x)) + ((ax52x) & (ax51x) & (!ax50x) & (ax49x) & (shiftx0x) & (!shiftx1x)) + ((ax52x) & (ax51x) & (!ax50x) & (ax49x) & (shiftx0x) & (shiftx1x)) + ((ax52x) & (ax51x) & (ax50x) & (!ax49x) & (!shiftx0x) & (!shiftx1x)) + ((ax52x) & (ax51x) & (ax50x) & (!ax49x) & (!shiftx0x) & (shiftx1x)) + ((ax52x) & (ax51x) & (ax50x) & (!ax49x) & (shiftx0x) & (!shiftx1x)) + ((ax52x) & (ax51x) & (ax50x) & (ax49x) & (!shiftx0x) & (!shiftx1x)) + ((ax52x) & (ax51x) & (ax50x) & (ax49x) & (!shiftx0x) & (shiftx1x)) + ((ax52x) & (ax51x) & (ax50x) & (ax49x) & (shiftx0x) & (!shiftx1x)) + ((ax52x) & (ax51x) & (ax50x) & (ax49x) & (shiftx0x) & (shiftx1x)));
	assign g14 = (((!ax56x) & (!ax55x) & (!ax54x) & (ax53x) & (shiftx0x) & (shiftx1x)) + ((!ax56x) & (!ax55x) & (ax54x) & (!ax53x) & (!shiftx0x) & (shiftx1x)) + ((!ax56x) & (!ax55x) & (ax54x) & (ax53x) & (!shiftx0x) & (shiftx1x)) + ((!ax56x) & (!ax55x) & (ax54x) & (ax53x) & (shiftx0x) & (shiftx1x)) + ((!ax56x) & (ax55x) & (!ax54x) & (!ax53x) & (shiftx0x) & (!shiftx1x)) + ((!ax56x) & (ax55x) & (!ax54x) & (ax53x) & (shiftx0x) & (!shiftx1x)) + ((!ax56x) & (ax55x) & (!ax54x) & (ax53x) & (shiftx0x) & (shiftx1x)) + ((!ax56x) & (ax55x) & (ax54x) & (!ax53x) & (!shiftx0x) & (shiftx1x)) + ((!ax56x) & (ax55x) & (ax54x) & (!ax53x) & (shiftx0x) & (!shiftx1x)) + ((!ax56x) & (ax55x) & (ax54x) & (ax53x) & (!shiftx0x) & (shiftx1x)) + ((!ax56x) & (ax55x) & (ax54x) & (ax53x) & (shiftx0x) & (!shiftx1x)) + ((!ax56x) & (ax55x) & (ax54x) & (ax53x) & (shiftx0x) & (shiftx1x)) + ((ax56x) & (!ax55x) & (!ax54x) & (!ax53x) & (!shiftx0x) & (!shiftx1x)) + ((ax56x) & (!ax55x) & (!ax54x) & (ax53x) & (!shiftx0x) & (!shiftx1x)) + ((ax56x) & (!ax55x) & (!ax54x) & (ax53x) & (shiftx0x) & (shiftx1x)) + ((ax56x) & (!ax55x) & (ax54x) & (!ax53x) & (!shiftx0x) & (!shiftx1x)) + ((ax56x) & (!ax55x) & (ax54x) & (!ax53x) & (!shiftx0x) & (shiftx1x)) + ((ax56x) & (!ax55x) & (ax54x) & (ax53x) & (!shiftx0x) & (!shiftx1x)) + ((ax56x) & (!ax55x) & (ax54x) & (ax53x) & (!shiftx0x) & (shiftx1x)) + ((ax56x) & (!ax55x) & (ax54x) & (ax53x) & (shiftx0x) & (shiftx1x)) + ((ax56x) & (ax55x) & (!ax54x) & (!ax53x) & (!shiftx0x) & (!shiftx1x)) + ((ax56x) & (ax55x) & (!ax54x) & (!ax53x) & (shiftx0x) & (!shiftx1x)) + ((ax56x) & (ax55x) & (!ax54x) & (ax53x) & (!shiftx0x) & (!shiftx1x)) + ((ax56x) & (ax55x) & (!ax54x) & (ax53x) & (shiftx0x) & (!shiftx1x)) + ((ax56x) & (ax55x) & (!ax54x) & (ax53x) & (shiftx0x) & (shiftx1x)) + ((ax56x) & (ax55x) & (ax54x) & (!ax53x) & (!shiftx0x) & (!shiftx1x)) + ((ax56x) & (ax55x) & (ax54x) & (!ax53x) & (!shiftx0x) & (shiftx1x)) + ((ax56x) & (ax55x) & (ax54x) & (!ax53x) & (shiftx0x) & (!shiftx1x)) + ((ax56x) & (ax55x) & (ax54x) & (ax53x) & (!shiftx0x) & (!shiftx1x)) + ((ax56x) & (ax55x) & (ax54x) & (ax53x) & (!shiftx0x) & (shiftx1x)) + ((ax56x) & (ax55x) & (ax54x) & (ax53x) & (shiftx0x) & (!shiftx1x)) + ((ax56x) & (ax55x) & (ax54x) & (ax53x) & (shiftx0x) & (shiftx1x)));
	assign g15 = (((!shiftx2x) & (!shiftx3x) & (g11) & (!g12) & (!g13) & (!g14)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (!g12) & (!g13) & (g14)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (!g12) & (g13) & (!g14)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (!g12) & (g13) & (g14)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (g12) & (!g13) & (!g14)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (g12) & (!g13) & (g14)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (g12) & (g13) & (!g14)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (g12) & (g13) & (g14)) + ((!shiftx2x) & (shiftx3x) & (!g11) & (!g12) & (!g13) & (g14)) + ((!shiftx2x) & (shiftx3x) & (!g11) & (!g12) & (g13) & (g14)) + ((!shiftx2x) & (shiftx3x) & (!g11) & (g12) & (!g13) & (g14)) + ((!shiftx2x) & (shiftx3x) & (!g11) & (g12) & (g13) & (g14)) + ((!shiftx2x) & (shiftx3x) & (g11) & (!g12) & (!g13) & (g14)) + ((!shiftx2x) & (shiftx3x) & (g11) & (!g12) & (g13) & (g14)) + ((!shiftx2x) & (shiftx3x) & (g11) & (g12) & (!g13) & (g14)) + ((!shiftx2x) & (shiftx3x) & (g11) & (g12) & (g13) & (g14)) + ((shiftx2x) & (!shiftx3x) & (!g11) & (g12) & (!g13) & (!g14)) + ((shiftx2x) & (!shiftx3x) & (!g11) & (g12) & (!g13) & (g14)) + ((shiftx2x) & (!shiftx3x) & (!g11) & (g12) & (g13) & (!g14)) + ((shiftx2x) & (!shiftx3x) & (!g11) & (g12) & (g13) & (g14)) + ((shiftx2x) & (!shiftx3x) & (g11) & (g12) & (!g13) & (!g14)) + ((shiftx2x) & (!shiftx3x) & (g11) & (g12) & (!g13) & (g14)) + ((shiftx2x) & (!shiftx3x) & (g11) & (g12) & (g13) & (!g14)) + ((shiftx2x) & (!shiftx3x) & (g11) & (g12) & (g13) & (g14)) + ((shiftx2x) & (shiftx3x) & (!g11) & (!g12) & (g13) & (!g14)) + ((shiftx2x) & (shiftx3x) & (!g11) & (!g12) & (g13) & (g14)) + ((shiftx2x) & (shiftx3x) & (!g11) & (g12) & (g13) & (!g14)) + ((shiftx2x) & (shiftx3x) & (!g11) & (g12) & (g13) & (g14)) + ((shiftx2x) & (shiftx3x) & (g11) & (!g12) & (g13) & (!g14)) + ((shiftx2x) & (shiftx3x) & (g11) & (!g12) & (g13) & (g14)) + ((shiftx2x) & (shiftx3x) & (g11) & (g12) & (g13) & (!g14)) + ((shiftx2x) & (shiftx3x) & (g11) & (g12) & (g13) & (g14)));
	assign g16 = (((!ax48x) & (!ax47x) & (!ax46x) & (ax45x) & (shiftx0x) & (shiftx1x)) + ((!ax48x) & (!ax47x) & (ax46x) & (!ax45x) & (!shiftx0x) & (shiftx1x)) + ((!ax48x) & (!ax47x) & (ax46x) & (ax45x) & (!shiftx0x) & (shiftx1x)) + ((!ax48x) & (!ax47x) & (ax46x) & (ax45x) & (shiftx0x) & (shiftx1x)) + ((!ax48x) & (ax47x) & (!ax46x) & (!ax45x) & (shiftx0x) & (!shiftx1x)) + ((!ax48x) & (ax47x) & (!ax46x) & (ax45x) & (shiftx0x) & (!shiftx1x)) + ((!ax48x) & (ax47x) & (!ax46x) & (ax45x) & (shiftx0x) & (shiftx1x)) + ((!ax48x) & (ax47x) & (ax46x) & (!ax45x) & (!shiftx0x) & (shiftx1x)) + ((!ax48x) & (ax47x) & (ax46x) & (!ax45x) & (shiftx0x) & (!shiftx1x)) + ((!ax48x) & (ax47x) & (ax46x) & (ax45x) & (!shiftx0x) & (shiftx1x)) + ((!ax48x) & (ax47x) & (ax46x) & (ax45x) & (shiftx0x) & (!shiftx1x)) + ((!ax48x) & (ax47x) & (ax46x) & (ax45x) & (shiftx0x) & (shiftx1x)) + ((ax48x) & (!ax47x) & (!ax46x) & (!ax45x) & (!shiftx0x) & (!shiftx1x)) + ((ax48x) & (!ax47x) & (!ax46x) & (ax45x) & (!shiftx0x) & (!shiftx1x)) + ((ax48x) & (!ax47x) & (!ax46x) & (ax45x) & (shiftx0x) & (shiftx1x)) + ((ax48x) & (!ax47x) & (ax46x) & (!ax45x) & (!shiftx0x) & (!shiftx1x)) + ((ax48x) & (!ax47x) & (ax46x) & (!ax45x) & (!shiftx0x) & (shiftx1x)) + ((ax48x) & (!ax47x) & (ax46x) & (ax45x) & (!shiftx0x) & (!shiftx1x)) + ((ax48x) & (!ax47x) & (ax46x) & (ax45x) & (!shiftx0x) & (shiftx1x)) + ((ax48x) & (!ax47x) & (ax46x) & (ax45x) & (shiftx0x) & (shiftx1x)) + ((ax48x) & (ax47x) & (!ax46x) & (!ax45x) & (!shiftx0x) & (!shiftx1x)) + ((ax48x) & (ax47x) & (!ax46x) & (!ax45x) & (shiftx0x) & (!shiftx1x)) + ((ax48x) & (ax47x) & (!ax46x) & (ax45x) & (!shiftx0x) & (!shiftx1x)) + ((ax48x) & (ax47x) & (!ax46x) & (ax45x) & (shiftx0x) & (!shiftx1x)) + ((ax48x) & (ax47x) & (!ax46x) & (ax45x) & (shiftx0x) & (shiftx1x)) + ((ax48x) & (ax47x) & (ax46x) & (!ax45x) & (!shiftx0x) & (!shiftx1x)) + ((ax48x) & (ax47x) & (ax46x) & (!ax45x) & (!shiftx0x) & (shiftx1x)) + ((ax48x) & (ax47x) & (ax46x) & (!ax45x) & (shiftx0x) & (!shiftx1x)) + ((ax48x) & (ax47x) & (ax46x) & (ax45x) & (!shiftx0x) & (!shiftx1x)) + ((ax48x) & (ax47x) & (ax46x) & (ax45x) & (!shiftx0x) & (shiftx1x)) + ((ax48x) & (ax47x) & (ax46x) & (ax45x) & (shiftx0x) & (!shiftx1x)) + ((ax48x) & (ax47x) & (ax46x) & (ax45x) & (shiftx0x) & (shiftx1x)));
	assign g17 = (((!ax44x) & (!ax43x) & (!ax42x) & (ax41x) & (shiftx0x) & (shiftx1x)) + ((!ax44x) & (!ax43x) & (ax42x) & (!ax41x) & (!shiftx0x) & (shiftx1x)) + ((!ax44x) & (!ax43x) & (ax42x) & (ax41x) & (!shiftx0x) & (shiftx1x)) + ((!ax44x) & (!ax43x) & (ax42x) & (ax41x) & (shiftx0x) & (shiftx1x)) + ((!ax44x) & (ax43x) & (!ax42x) & (!ax41x) & (shiftx0x) & (!shiftx1x)) + ((!ax44x) & (ax43x) & (!ax42x) & (ax41x) & (shiftx0x) & (!shiftx1x)) + ((!ax44x) & (ax43x) & (!ax42x) & (ax41x) & (shiftx0x) & (shiftx1x)) + ((!ax44x) & (ax43x) & (ax42x) & (!ax41x) & (!shiftx0x) & (shiftx1x)) + ((!ax44x) & (ax43x) & (ax42x) & (!ax41x) & (shiftx0x) & (!shiftx1x)) + ((!ax44x) & (ax43x) & (ax42x) & (ax41x) & (!shiftx0x) & (shiftx1x)) + ((!ax44x) & (ax43x) & (ax42x) & (ax41x) & (shiftx0x) & (!shiftx1x)) + ((!ax44x) & (ax43x) & (ax42x) & (ax41x) & (shiftx0x) & (shiftx1x)) + ((ax44x) & (!ax43x) & (!ax42x) & (!ax41x) & (!shiftx0x) & (!shiftx1x)) + ((ax44x) & (!ax43x) & (!ax42x) & (ax41x) & (!shiftx0x) & (!shiftx1x)) + ((ax44x) & (!ax43x) & (!ax42x) & (ax41x) & (shiftx0x) & (shiftx1x)) + ((ax44x) & (!ax43x) & (ax42x) & (!ax41x) & (!shiftx0x) & (!shiftx1x)) + ((ax44x) & (!ax43x) & (ax42x) & (!ax41x) & (!shiftx0x) & (shiftx1x)) + ((ax44x) & (!ax43x) & (ax42x) & (ax41x) & (!shiftx0x) & (!shiftx1x)) + ((ax44x) & (!ax43x) & (ax42x) & (ax41x) & (!shiftx0x) & (shiftx1x)) + ((ax44x) & (!ax43x) & (ax42x) & (ax41x) & (shiftx0x) & (shiftx1x)) + ((ax44x) & (ax43x) & (!ax42x) & (!ax41x) & (!shiftx0x) & (!shiftx1x)) + ((ax44x) & (ax43x) & (!ax42x) & (!ax41x) & (shiftx0x) & (!shiftx1x)) + ((ax44x) & (ax43x) & (!ax42x) & (ax41x) & (!shiftx0x) & (!shiftx1x)) + ((ax44x) & (ax43x) & (!ax42x) & (ax41x) & (shiftx0x) & (!shiftx1x)) + ((ax44x) & (ax43x) & (!ax42x) & (ax41x) & (shiftx0x) & (shiftx1x)) + ((ax44x) & (ax43x) & (ax42x) & (!ax41x) & (!shiftx0x) & (!shiftx1x)) + ((ax44x) & (ax43x) & (ax42x) & (!ax41x) & (!shiftx0x) & (shiftx1x)) + ((ax44x) & (ax43x) & (ax42x) & (!ax41x) & (shiftx0x) & (!shiftx1x)) + ((ax44x) & (ax43x) & (ax42x) & (ax41x) & (!shiftx0x) & (!shiftx1x)) + ((ax44x) & (ax43x) & (ax42x) & (ax41x) & (!shiftx0x) & (shiftx1x)) + ((ax44x) & (ax43x) & (ax42x) & (ax41x) & (shiftx0x) & (!shiftx1x)) + ((ax44x) & (ax43x) & (ax42x) & (ax41x) & (shiftx0x) & (shiftx1x)));
	assign g18 = (((!ax36x) & (!ax35x) & (!ax34x) & (ax33x) & (shiftx0x) & (shiftx1x)) + ((!ax36x) & (!ax35x) & (ax34x) & (!ax33x) & (!shiftx0x) & (shiftx1x)) + ((!ax36x) & (!ax35x) & (ax34x) & (ax33x) & (!shiftx0x) & (shiftx1x)) + ((!ax36x) & (!ax35x) & (ax34x) & (ax33x) & (shiftx0x) & (shiftx1x)) + ((!ax36x) & (ax35x) & (!ax34x) & (!ax33x) & (shiftx0x) & (!shiftx1x)) + ((!ax36x) & (ax35x) & (!ax34x) & (ax33x) & (shiftx0x) & (!shiftx1x)) + ((!ax36x) & (ax35x) & (!ax34x) & (ax33x) & (shiftx0x) & (shiftx1x)) + ((!ax36x) & (ax35x) & (ax34x) & (!ax33x) & (!shiftx0x) & (shiftx1x)) + ((!ax36x) & (ax35x) & (ax34x) & (!ax33x) & (shiftx0x) & (!shiftx1x)) + ((!ax36x) & (ax35x) & (ax34x) & (ax33x) & (!shiftx0x) & (shiftx1x)) + ((!ax36x) & (ax35x) & (ax34x) & (ax33x) & (shiftx0x) & (!shiftx1x)) + ((!ax36x) & (ax35x) & (ax34x) & (ax33x) & (shiftx0x) & (shiftx1x)) + ((ax36x) & (!ax35x) & (!ax34x) & (!ax33x) & (!shiftx0x) & (!shiftx1x)) + ((ax36x) & (!ax35x) & (!ax34x) & (ax33x) & (!shiftx0x) & (!shiftx1x)) + ((ax36x) & (!ax35x) & (!ax34x) & (ax33x) & (shiftx0x) & (shiftx1x)) + ((ax36x) & (!ax35x) & (ax34x) & (!ax33x) & (!shiftx0x) & (!shiftx1x)) + ((ax36x) & (!ax35x) & (ax34x) & (!ax33x) & (!shiftx0x) & (shiftx1x)) + ((ax36x) & (!ax35x) & (ax34x) & (ax33x) & (!shiftx0x) & (!shiftx1x)) + ((ax36x) & (!ax35x) & (ax34x) & (ax33x) & (!shiftx0x) & (shiftx1x)) + ((ax36x) & (!ax35x) & (ax34x) & (ax33x) & (shiftx0x) & (shiftx1x)) + ((ax36x) & (ax35x) & (!ax34x) & (!ax33x) & (!shiftx0x) & (!shiftx1x)) + ((ax36x) & (ax35x) & (!ax34x) & (!ax33x) & (shiftx0x) & (!shiftx1x)) + ((ax36x) & (ax35x) & (!ax34x) & (ax33x) & (!shiftx0x) & (!shiftx1x)) + ((ax36x) & (ax35x) & (!ax34x) & (ax33x) & (shiftx0x) & (!shiftx1x)) + ((ax36x) & (ax35x) & (!ax34x) & (ax33x) & (shiftx0x) & (shiftx1x)) + ((ax36x) & (ax35x) & (ax34x) & (!ax33x) & (!shiftx0x) & (!shiftx1x)) + ((ax36x) & (ax35x) & (ax34x) & (!ax33x) & (!shiftx0x) & (shiftx1x)) + ((ax36x) & (ax35x) & (ax34x) & (!ax33x) & (shiftx0x) & (!shiftx1x)) + ((ax36x) & (ax35x) & (ax34x) & (ax33x) & (!shiftx0x) & (!shiftx1x)) + ((ax36x) & (ax35x) & (ax34x) & (ax33x) & (!shiftx0x) & (shiftx1x)) + ((ax36x) & (ax35x) & (ax34x) & (ax33x) & (shiftx0x) & (!shiftx1x)) + ((ax36x) & (ax35x) & (ax34x) & (ax33x) & (shiftx0x) & (shiftx1x)));
	assign g19 = (((!ax40x) & (!ax38x) & (!ax39x) & (ax37x) & (shiftx1x) & (shiftx0x)) + ((!ax40x) & (!ax38x) & (ax39x) & (!ax37x) & (!shiftx1x) & (shiftx0x)) + ((!ax40x) & (!ax38x) & (ax39x) & (ax37x) & (!shiftx1x) & (shiftx0x)) + ((!ax40x) & (!ax38x) & (ax39x) & (ax37x) & (shiftx1x) & (shiftx0x)) + ((!ax40x) & (ax38x) & (!ax39x) & (!ax37x) & (shiftx1x) & (!shiftx0x)) + ((!ax40x) & (ax38x) & (!ax39x) & (ax37x) & (shiftx1x) & (!shiftx0x)) + ((!ax40x) & (ax38x) & (!ax39x) & (ax37x) & (shiftx1x) & (shiftx0x)) + ((!ax40x) & (ax38x) & (ax39x) & (!ax37x) & (!shiftx1x) & (shiftx0x)) + ((!ax40x) & (ax38x) & (ax39x) & (!ax37x) & (shiftx1x) & (!shiftx0x)) + ((!ax40x) & (ax38x) & (ax39x) & (ax37x) & (!shiftx1x) & (shiftx0x)) + ((!ax40x) & (ax38x) & (ax39x) & (ax37x) & (shiftx1x) & (!shiftx0x)) + ((!ax40x) & (ax38x) & (ax39x) & (ax37x) & (shiftx1x) & (shiftx0x)) + ((ax40x) & (!ax38x) & (!ax39x) & (!ax37x) & (!shiftx1x) & (!shiftx0x)) + ((ax40x) & (!ax38x) & (!ax39x) & (ax37x) & (!shiftx1x) & (!shiftx0x)) + ((ax40x) & (!ax38x) & (!ax39x) & (ax37x) & (shiftx1x) & (shiftx0x)) + ((ax40x) & (!ax38x) & (ax39x) & (!ax37x) & (!shiftx1x) & (!shiftx0x)) + ((ax40x) & (!ax38x) & (ax39x) & (!ax37x) & (!shiftx1x) & (shiftx0x)) + ((ax40x) & (!ax38x) & (ax39x) & (ax37x) & (!shiftx1x) & (!shiftx0x)) + ((ax40x) & (!ax38x) & (ax39x) & (ax37x) & (!shiftx1x) & (shiftx0x)) + ((ax40x) & (!ax38x) & (ax39x) & (ax37x) & (shiftx1x) & (shiftx0x)) + ((ax40x) & (ax38x) & (!ax39x) & (!ax37x) & (!shiftx1x) & (!shiftx0x)) + ((ax40x) & (ax38x) & (!ax39x) & (!ax37x) & (shiftx1x) & (!shiftx0x)) + ((ax40x) & (ax38x) & (!ax39x) & (ax37x) & (!shiftx1x) & (!shiftx0x)) + ((ax40x) & (ax38x) & (!ax39x) & (ax37x) & (shiftx1x) & (!shiftx0x)) + ((ax40x) & (ax38x) & (!ax39x) & (ax37x) & (shiftx1x) & (shiftx0x)) + ((ax40x) & (ax38x) & (ax39x) & (!ax37x) & (!shiftx1x) & (!shiftx0x)) + ((ax40x) & (ax38x) & (ax39x) & (!ax37x) & (!shiftx1x) & (shiftx0x)) + ((ax40x) & (ax38x) & (ax39x) & (!ax37x) & (shiftx1x) & (!shiftx0x)) + ((ax40x) & (ax38x) & (ax39x) & (ax37x) & (!shiftx1x) & (!shiftx0x)) + ((ax40x) & (ax38x) & (ax39x) & (ax37x) & (!shiftx1x) & (shiftx0x)) + ((ax40x) & (ax38x) & (ax39x) & (ax37x) & (shiftx1x) & (!shiftx0x)) + ((ax40x) & (ax38x) & (ax39x) & (ax37x) & (shiftx1x) & (shiftx0x)));
	assign g20 = (((!shiftx2x) & (!shiftx3x) & (g16) & (!g17) & (!g18) & (!g19)) + ((!shiftx2x) & (!shiftx3x) & (g16) & (!g17) & (!g18) & (g19)) + ((!shiftx2x) & (!shiftx3x) & (g16) & (!g17) & (g18) & (!g19)) + ((!shiftx2x) & (!shiftx3x) & (g16) & (!g17) & (g18) & (g19)) + ((!shiftx2x) & (!shiftx3x) & (g16) & (g17) & (!g18) & (!g19)) + ((!shiftx2x) & (!shiftx3x) & (g16) & (g17) & (!g18) & (g19)) + ((!shiftx2x) & (!shiftx3x) & (g16) & (g17) & (g18) & (!g19)) + ((!shiftx2x) & (!shiftx3x) & (g16) & (g17) & (g18) & (g19)) + ((!shiftx2x) & (shiftx3x) & (!g16) & (!g17) & (!g18) & (g19)) + ((!shiftx2x) & (shiftx3x) & (!g16) & (!g17) & (g18) & (g19)) + ((!shiftx2x) & (shiftx3x) & (!g16) & (g17) & (!g18) & (g19)) + ((!shiftx2x) & (shiftx3x) & (!g16) & (g17) & (g18) & (g19)) + ((!shiftx2x) & (shiftx3x) & (g16) & (!g17) & (!g18) & (g19)) + ((!shiftx2x) & (shiftx3x) & (g16) & (!g17) & (g18) & (g19)) + ((!shiftx2x) & (shiftx3x) & (g16) & (g17) & (!g18) & (g19)) + ((!shiftx2x) & (shiftx3x) & (g16) & (g17) & (g18) & (g19)) + ((shiftx2x) & (!shiftx3x) & (!g16) & (g17) & (!g18) & (!g19)) + ((shiftx2x) & (!shiftx3x) & (!g16) & (g17) & (!g18) & (g19)) + ((shiftx2x) & (!shiftx3x) & (!g16) & (g17) & (g18) & (!g19)) + ((shiftx2x) & (!shiftx3x) & (!g16) & (g17) & (g18) & (g19)) + ((shiftx2x) & (!shiftx3x) & (g16) & (g17) & (!g18) & (!g19)) + ((shiftx2x) & (!shiftx3x) & (g16) & (g17) & (!g18) & (g19)) + ((shiftx2x) & (!shiftx3x) & (g16) & (g17) & (g18) & (!g19)) + ((shiftx2x) & (!shiftx3x) & (g16) & (g17) & (g18) & (g19)) + ((shiftx2x) & (shiftx3x) & (!g16) & (!g17) & (g18) & (!g19)) + ((shiftx2x) & (shiftx3x) & (!g16) & (!g17) & (g18) & (g19)) + ((shiftx2x) & (shiftx3x) & (!g16) & (g17) & (g18) & (!g19)) + ((shiftx2x) & (shiftx3x) & (!g16) & (g17) & (g18) & (g19)) + ((shiftx2x) & (shiftx3x) & (g16) & (!g17) & (g18) & (!g19)) + ((shiftx2x) & (shiftx3x) & (g16) & (!g17) & (g18) & (g19)) + ((shiftx2x) & (shiftx3x) & (g16) & (g17) & (g18) & (!g19)) + ((shiftx2x) & (shiftx3x) & (g16) & (g17) & (g18) & (g19)));
	assign g21 = (((!shiftx4x) & (!shiftx5x) & (!g5) & (!g10) & (g15) & (!g20)) + ((!shiftx4x) & (!shiftx5x) & (!g5) & (!g10) & (g15) & (g20)) + ((!shiftx4x) & (!shiftx5x) & (!g5) & (g10) & (g15) & (!g20)) + ((!shiftx4x) & (!shiftx5x) & (!g5) & (g10) & (g15) & (g20)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (!g10) & (g15) & (!g20)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (!g10) & (g15) & (g20)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (g10) & (g15) & (!g20)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (g10) & (g15) & (g20)) + ((!shiftx4x) & (shiftx5x) & (!g5) & (g10) & (!g15) & (!g20)) + ((!shiftx4x) & (shiftx5x) & (!g5) & (g10) & (!g15) & (g20)) + ((!shiftx4x) & (shiftx5x) & (!g5) & (g10) & (g15) & (!g20)) + ((!shiftx4x) & (shiftx5x) & (!g5) & (g10) & (g15) & (g20)) + ((!shiftx4x) & (shiftx5x) & (g5) & (g10) & (!g15) & (!g20)) + ((!shiftx4x) & (shiftx5x) & (g5) & (g10) & (!g15) & (g20)) + ((!shiftx4x) & (shiftx5x) & (g5) & (g10) & (g15) & (!g20)) + ((!shiftx4x) & (shiftx5x) & (g5) & (g10) & (g15) & (g20)) + ((shiftx4x) & (!shiftx5x) & (!g5) & (!g10) & (!g15) & (g20)) + ((shiftx4x) & (!shiftx5x) & (!g5) & (!g10) & (g15) & (g20)) + ((shiftx4x) & (!shiftx5x) & (!g5) & (g10) & (!g15) & (g20)) + ((shiftx4x) & (!shiftx5x) & (!g5) & (g10) & (g15) & (g20)) + ((shiftx4x) & (!shiftx5x) & (g5) & (!g10) & (!g15) & (g20)) + ((shiftx4x) & (!shiftx5x) & (g5) & (!g10) & (g15) & (g20)) + ((shiftx4x) & (!shiftx5x) & (g5) & (g10) & (!g15) & (g20)) + ((shiftx4x) & (!shiftx5x) & (g5) & (g10) & (g15) & (g20)) + ((shiftx4x) & (shiftx5x) & (g5) & (!g10) & (!g15) & (!g20)) + ((shiftx4x) & (shiftx5x) & (g5) & (!g10) & (!g15) & (g20)) + ((shiftx4x) & (shiftx5x) & (g5) & (!g10) & (g15) & (!g20)) + ((shiftx4x) & (shiftx5x) & (g5) & (!g10) & (g15) & (g20)) + ((shiftx4x) & (shiftx5x) & (g5) & (g10) & (!g15) & (!g20)) + ((shiftx4x) & (shiftx5x) & (g5) & (g10) & (!g15) & (g20)) + ((shiftx4x) & (shiftx5x) & (g5) & (g10) & (g15) & (!g20)) + ((shiftx4x) & (shiftx5x) & (g5) & (g10) & (g15) & (g20)));
	assign g22 = (((!ax80x) & (!ax79x) & (!ax78x) & (ax77x) & (shiftx0x) & (shiftx1x)) + ((!ax80x) & (!ax79x) & (ax78x) & (!ax77x) & (!shiftx0x) & (shiftx1x)) + ((!ax80x) & (!ax79x) & (ax78x) & (ax77x) & (!shiftx0x) & (shiftx1x)) + ((!ax80x) & (!ax79x) & (ax78x) & (ax77x) & (shiftx0x) & (shiftx1x)) + ((!ax80x) & (ax79x) & (!ax78x) & (!ax77x) & (shiftx0x) & (!shiftx1x)) + ((!ax80x) & (ax79x) & (!ax78x) & (ax77x) & (shiftx0x) & (!shiftx1x)) + ((!ax80x) & (ax79x) & (!ax78x) & (ax77x) & (shiftx0x) & (shiftx1x)) + ((!ax80x) & (ax79x) & (ax78x) & (!ax77x) & (!shiftx0x) & (shiftx1x)) + ((!ax80x) & (ax79x) & (ax78x) & (!ax77x) & (shiftx0x) & (!shiftx1x)) + ((!ax80x) & (ax79x) & (ax78x) & (ax77x) & (!shiftx0x) & (shiftx1x)) + ((!ax80x) & (ax79x) & (ax78x) & (ax77x) & (shiftx0x) & (!shiftx1x)) + ((!ax80x) & (ax79x) & (ax78x) & (ax77x) & (shiftx0x) & (shiftx1x)) + ((ax80x) & (!ax79x) & (!ax78x) & (!ax77x) & (!shiftx0x) & (!shiftx1x)) + ((ax80x) & (!ax79x) & (!ax78x) & (ax77x) & (!shiftx0x) & (!shiftx1x)) + ((ax80x) & (!ax79x) & (!ax78x) & (ax77x) & (shiftx0x) & (shiftx1x)) + ((ax80x) & (!ax79x) & (ax78x) & (!ax77x) & (!shiftx0x) & (!shiftx1x)) + ((ax80x) & (!ax79x) & (ax78x) & (!ax77x) & (!shiftx0x) & (shiftx1x)) + ((ax80x) & (!ax79x) & (ax78x) & (ax77x) & (!shiftx0x) & (!shiftx1x)) + ((ax80x) & (!ax79x) & (ax78x) & (ax77x) & (!shiftx0x) & (shiftx1x)) + ((ax80x) & (!ax79x) & (ax78x) & (ax77x) & (shiftx0x) & (shiftx1x)) + ((ax80x) & (ax79x) & (!ax78x) & (!ax77x) & (!shiftx0x) & (!shiftx1x)) + ((ax80x) & (ax79x) & (!ax78x) & (!ax77x) & (shiftx0x) & (!shiftx1x)) + ((ax80x) & (ax79x) & (!ax78x) & (ax77x) & (!shiftx0x) & (!shiftx1x)) + ((ax80x) & (ax79x) & (!ax78x) & (ax77x) & (shiftx0x) & (!shiftx1x)) + ((ax80x) & (ax79x) & (!ax78x) & (ax77x) & (shiftx0x) & (shiftx1x)) + ((ax80x) & (ax79x) & (ax78x) & (!ax77x) & (!shiftx0x) & (!shiftx1x)) + ((ax80x) & (ax79x) & (ax78x) & (!ax77x) & (!shiftx0x) & (shiftx1x)) + ((ax80x) & (ax79x) & (ax78x) & (!ax77x) & (shiftx0x) & (!shiftx1x)) + ((ax80x) & (ax79x) & (ax78x) & (ax77x) & (!shiftx0x) & (!shiftx1x)) + ((ax80x) & (ax79x) & (ax78x) & (ax77x) & (!shiftx0x) & (shiftx1x)) + ((ax80x) & (ax79x) & (ax78x) & (ax77x) & (shiftx0x) & (!shiftx1x)) + ((ax80x) & (ax79x) & (ax78x) & (ax77x) & (shiftx0x) & (shiftx1x)));
	assign g23 = (((!ax76x) & (!ax75x) & (!ax74x) & (ax73x) & (shiftx0x) & (shiftx1x)) + ((!ax76x) & (!ax75x) & (ax74x) & (!ax73x) & (!shiftx0x) & (shiftx1x)) + ((!ax76x) & (!ax75x) & (ax74x) & (ax73x) & (!shiftx0x) & (shiftx1x)) + ((!ax76x) & (!ax75x) & (ax74x) & (ax73x) & (shiftx0x) & (shiftx1x)) + ((!ax76x) & (ax75x) & (!ax74x) & (!ax73x) & (shiftx0x) & (!shiftx1x)) + ((!ax76x) & (ax75x) & (!ax74x) & (ax73x) & (shiftx0x) & (!shiftx1x)) + ((!ax76x) & (ax75x) & (!ax74x) & (ax73x) & (shiftx0x) & (shiftx1x)) + ((!ax76x) & (ax75x) & (ax74x) & (!ax73x) & (!shiftx0x) & (shiftx1x)) + ((!ax76x) & (ax75x) & (ax74x) & (!ax73x) & (shiftx0x) & (!shiftx1x)) + ((!ax76x) & (ax75x) & (ax74x) & (ax73x) & (!shiftx0x) & (shiftx1x)) + ((!ax76x) & (ax75x) & (ax74x) & (ax73x) & (shiftx0x) & (!shiftx1x)) + ((!ax76x) & (ax75x) & (ax74x) & (ax73x) & (shiftx0x) & (shiftx1x)) + ((ax76x) & (!ax75x) & (!ax74x) & (!ax73x) & (!shiftx0x) & (!shiftx1x)) + ((ax76x) & (!ax75x) & (!ax74x) & (ax73x) & (!shiftx0x) & (!shiftx1x)) + ((ax76x) & (!ax75x) & (!ax74x) & (ax73x) & (shiftx0x) & (shiftx1x)) + ((ax76x) & (!ax75x) & (ax74x) & (!ax73x) & (!shiftx0x) & (!shiftx1x)) + ((ax76x) & (!ax75x) & (ax74x) & (!ax73x) & (!shiftx0x) & (shiftx1x)) + ((ax76x) & (!ax75x) & (ax74x) & (ax73x) & (!shiftx0x) & (!shiftx1x)) + ((ax76x) & (!ax75x) & (ax74x) & (ax73x) & (!shiftx0x) & (shiftx1x)) + ((ax76x) & (!ax75x) & (ax74x) & (ax73x) & (shiftx0x) & (shiftx1x)) + ((ax76x) & (ax75x) & (!ax74x) & (!ax73x) & (!shiftx0x) & (!shiftx1x)) + ((ax76x) & (ax75x) & (!ax74x) & (!ax73x) & (shiftx0x) & (!shiftx1x)) + ((ax76x) & (ax75x) & (!ax74x) & (ax73x) & (!shiftx0x) & (!shiftx1x)) + ((ax76x) & (ax75x) & (!ax74x) & (ax73x) & (shiftx0x) & (!shiftx1x)) + ((ax76x) & (ax75x) & (!ax74x) & (ax73x) & (shiftx0x) & (shiftx1x)) + ((ax76x) & (ax75x) & (ax74x) & (!ax73x) & (!shiftx0x) & (!shiftx1x)) + ((ax76x) & (ax75x) & (ax74x) & (!ax73x) & (!shiftx0x) & (shiftx1x)) + ((ax76x) & (ax75x) & (ax74x) & (!ax73x) & (shiftx0x) & (!shiftx1x)) + ((ax76x) & (ax75x) & (ax74x) & (ax73x) & (!shiftx0x) & (!shiftx1x)) + ((ax76x) & (ax75x) & (ax74x) & (ax73x) & (!shiftx0x) & (shiftx1x)) + ((ax76x) & (ax75x) & (ax74x) & (ax73x) & (shiftx0x) & (!shiftx1x)) + ((ax76x) & (ax75x) & (ax74x) & (ax73x) & (shiftx0x) & (shiftx1x)));
	assign g24 = (((!ax68x) & (!ax67x) & (!ax66x) & (ax65x) & (shiftx0x) & (shiftx1x)) + ((!ax68x) & (!ax67x) & (ax66x) & (!ax65x) & (!shiftx0x) & (shiftx1x)) + ((!ax68x) & (!ax67x) & (ax66x) & (ax65x) & (!shiftx0x) & (shiftx1x)) + ((!ax68x) & (!ax67x) & (ax66x) & (ax65x) & (shiftx0x) & (shiftx1x)) + ((!ax68x) & (ax67x) & (!ax66x) & (!ax65x) & (shiftx0x) & (!shiftx1x)) + ((!ax68x) & (ax67x) & (!ax66x) & (ax65x) & (shiftx0x) & (!shiftx1x)) + ((!ax68x) & (ax67x) & (!ax66x) & (ax65x) & (shiftx0x) & (shiftx1x)) + ((!ax68x) & (ax67x) & (ax66x) & (!ax65x) & (!shiftx0x) & (shiftx1x)) + ((!ax68x) & (ax67x) & (ax66x) & (!ax65x) & (shiftx0x) & (!shiftx1x)) + ((!ax68x) & (ax67x) & (ax66x) & (ax65x) & (!shiftx0x) & (shiftx1x)) + ((!ax68x) & (ax67x) & (ax66x) & (ax65x) & (shiftx0x) & (!shiftx1x)) + ((!ax68x) & (ax67x) & (ax66x) & (ax65x) & (shiftx0x) & (shiftx1x)) + ((ax68x) & (!ax67x) & (!ax66x) & (!ax65x) & (!shiftx0x) & (!shiftx1x)) + ((ax68x) & (!ax67x) & (!ax66x) & (ax65x) & (!shiftx0x) & (!shiftx1x)) + ((ax68x) & (!ax67x) & (!ax66x) & (ax65x) & (shiftx0x) & (shiftx1x)) + ((ax68x) & (!ax67x) & (ax66x) & (!ax65x) & (!shiftx0x) & (!shiftx1x)) + ((ax68x) & (!ax67x) & (ax66x) & (!ax65x) & (!shiftx0x) & (shiftx1x)) + ((ax68x) & (!ax67x) & (ax66x) & (ax65x) & (!shiftx0x) & (!shiftx1x)) + ((ax68x) & (!ax67x) & (ax66x) & (ax65x) & (!shiftx0x) & (shiftx1x)) + ((ax68x) & (!ax67x) & (ax66x) & (ax65x) & (shiftx0x) & (shiftx1x)) + ((ax68x) & (ax67x) & (!ax66x) & (!ax65x) & (!shiftx0x) & (!shiftx1x)) + ((ax68x) & (ax67x) & (!ax66x) & (!ax65x) & (shiftx0x) & (!shiftx1x)) + ((ax68x) & (ax67x) & (!ax66x) & (ax65x) & (!shiftx0x) & (!shiftx1x)) + ((ax68x) & (ax67x) & (!ax66x) & (ax65x) & (shiftx0x) & (!shiftx1x)) + ((ax68x) & (ax67x) & (!ax66x) & (ax65x) & (shiftx0x) & (shiftx1x)) + ((ax68x) & (ax67x) & (ax66x) & (!ax65x) & (!shiftx0x) & (!shiftx1x)) + ((ax68x) & (ax67x) & (ax66x) & (!ax65x) & (!shiftx0x) & (shiftx1x)) + ((ax68x) & (ax67x) & (ax66x) & (!ax65x) & (shiftx0x) & (!shiftx1x)) + ((ax68x) & (ax67x) & (ax66x) & (ax65x) & (!shiftx0x) & (!shiftx1x)) + ((ax68x) & (ax67x) & (ax66x) & (ax65x) & (!shiftx0x) & (shiftx1x)) + ((ax68x) & (ax67x) & (ax66x) & (ax65x) & (shiftx0x) & (!shiftx1x)) + ((ax68x) & (ax67x) & (ax66x) & (ax65x) & (shiftx0x) & (shiftx1x)));
	assign g25 = (((!ax72x) & (!ax71x) & (!ax70x) & (ax69x) & (shiftx0x) & (shiftx1x)) + ((!ax72x) & (!ax71x) & (ax70x) & (!ax69x) & (!shiftx0x) & (shiftx1x)) + ((!ax72x) & (!ax71x) & (ax70x) & (ax69x) & (!shiftx0x) & (shiftx1x)) + ((!ax72x) & (!ax71x) & (ax70x) & (ax69x) & (shiftx0x) & (shiftx1x)) + ((!ax72x) & (ax71x) & (!ax70x) & (!ax69x) & (shiftx0x) & (!shiftx1x)) + ((!ax72x) & (ax71x) & (!ax70x) & (ax69x) & (shiftx0x) & (!shiftx1x)) + ((!ax72x) & (ax71x) & (!ax70x) & (ax69x) & (shiftx0x) & (shiftx1x)) + ((!ax72x) & (ax71x) & (ax70x) & (!ax69x) & (!shiftx0x) & (shiftx1x)) + ((!ax72x) & (ax71x) & (ax70x) & (!ax69x) & (shiftx0x) & (!shiftx1x)) + ((!ax72x) & (ax71x) & (ax70x) & (ax69x) & (!shiftx0x) & (shiftx1x)) + ((!ax72x) & (ax71x) & (ax70x) & (ax69x) & (shiftx0x) & (!shiftx1x)) + ((!ax72x) & (ax71x) & (ax70x) & (ax69x) & (shiftx0x) & (shiftx1x)) + ((ax72x) & (!ax71x) & (!ax70x) & (!ax69x) & (!shiftx0x) & (!shiftx1x)) + ((ax72x) & (!ax71x) & (!ax70x) & (ax69x) & (!shiftx0x) & (!shiftx1x)) + ((ax72x) & (!ax71x) & (!ax70x) & (ax69x) & (shiftx0x) & (shiftx1x)) + ((ax72x) & (!ax71x) & (ax70x) & (!ax69x) & (!shiftx0x) & (!shiftx1x)) + ((ax72x) & (!ax71x) & (ax70x) & (!ax69x) & (!shiftx0x) & (shiftx1x)) + ((ax72x) & (!ax71x) & (ax70x) & (ax69x) & (!shiftx0x) & (!shiftx1x)) + ((ax72x) & (!ax71x) & (ax70x) & (ax69x) & (!shiftx0x) & (shiftx1x)) + ((ax72x) & (!ax71x) & (ax70x) & (ax69x) & (shiftx0x) & (shiftx1x)) + ((ax72x) & (ax71x) & (!ax70x) & (!ax69x) & (!shiftx0x) & (!shiftx1x)) + ((ax72x) & (ax71x) & (!ax70x) & (!ax69x) & (shiftx0x) & (!shiftx1x)) + ((ax72x) & (ax71x) & (!ax70x) & (ax69x) & (!shiftx0x) & (!shiftx1x)) + ((ax72x) & (ax71x) & (!ax70x) & (ax69x) & (shiftx0x) & (!shiftx1x)) + ((ax72x) & (ax71x) & (!ax70x) & (ax69x) & (shiftx0x) & (shiftx1x)) + ((ax72x) & (ax71x) & (ax70x) & (!ax69x) & (!shiftx0x) & (!shiftx1x)) + ((ax72x) & (ax71x) & (ax70x) & (!ax69x) & (!shiftx0x) & (shiftx1x)) + ((ax72x) & (ax71x) & (ax70x) & (!ax69x) & (shiftx0x) & (!shiftx1x)) + ((ax72x) & (ax71x) & (ax70x) & (ax69x) & (!shiftx0x) & (!shiftx1x)) + ((ax72x) & (ax71x) & (ax70x) & (ax69x) & (!shiftx0x) & (shiftx1x)) + ((ax72x) & (ax71x) & (ax70x) & (ax69x) & (shiftx0x) & (!shiftx1x)) + ((ax72x) & (ax71x) & (ax70x) & (ax69x) & (shiftx0x) & (shiftx1x)));
	assign g26 = (((!shiftx2x) & (!shiftx3x) & (g22) & (!g23) & (!g24) & (!g25)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (!g23) & (!g24) & (g25)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (!g23) & (g24) & (!g25)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (!g23) & (g24) & (g25)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (g23) & (!g24) & (!g25)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (g23) & (!g24) & (g25)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (g23) & (g24) & (!g25)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (g23) & (g24) & (g25)) + ((!shiftx2x) & (shiftx3x) & (!g22) & (!g23) & (!g24) & (g25)) + ((!shiftx2x) & (shiftx3x) & (!g22) & (!g23) & (g24) & (g25)) + ((!shiftx2x) & (shiftx3x) & (!g22) & (g23) & (!g24) & (g25)) + ((!shiftx2x) & (shiftx3x) & (!g22) & (g23) & (g24) & (g25)) + ((!shiftx2x) & (shiftx3x) & (g22) & (!g23) & (!g24) & (g25)) + ((!shiftx2x) & (shiftx3x) & (g22) & (!g23) & (g24) & (g25)) + ((!shiftx2x) & (shiftx3x) & (g22) & (g23) & (!g24) & (g25)) + ((!shiftx2x) & (shiftx3x) & (g22) & (g23) & (g24) & (g25)) + ((shiftx2x) & (!shiftx3x) & (!g22) & (g23) & (!g24) & (!g25)) + ((shiftx2x) & (!shiftx3x) & (!g22) & (g23) & (!g24) & (g25)) + ((shiftx2x) & (!shiftx3x) & (!g22) & (g23) & (g24) & (!g25)) + ((shiftx2x) & (!shiftx3x) & (!g22) & (g23) & (g24) & (g25)) + ((shiftx2x) & (!shiftx3x) & (g22) & (g23) & (!g24) & (!g25)) + ((shiftx2x) & (!shiftx3x) & (g22) & (g23) & (!g24) & (g25)) + ((shiftx2x) & (!shiftx3x) & (g22) & (g23) & (g24) & (!g25)) + ((shiftx2x) & (!shiftx3x) & (g22) & (g23) & (g24) & (g25)) + ((shiftx2x) & (shiftx3x) & (!g22) & (!g23) & (g24) & (!g25)) + ((shiftx2x) & (shiftx3x) & (!g22) & (!g23) & (g24) & (g25)) + ((shiftx2x) & (shiftx3x) & (!g22) & (g23) & (g24) & (!g25)) + ((shiftx2x) & (shiftx3x) & (!g22) & (g23) & (g24) & (g25)) + ((shiftx2x) & (shiftx3x) & (g22) & (!g23) & (g24) & (!g25)) + ((shiftx2x) & (shiftx3x) & (g22) & (!g23) & (g24) & (g25)) + ((shiftx2x) & (shiftx3x) & (g22) & (g23) & (g24) & (!g25)) + ((shiftx2x) & (shiftx3x) & (g22) & (g23) & (g24) & (g25)));
	assign g27 = (((!ax96x) & (!ax95x) & (!ax94x) & (ax93x) & (shiftx0x) & (shiftx1x)) + ((!ax96x) & (!ax95x) & (ax94x) & (!ax93x) & (!shiftx0x) & (shiftx1x)) + ((!ax96x) & (!ax95x) & (ax94x) & (ax93x) & (!shiftx0x) & (shiftx1x)) + ((!ax96x) & (!ax95x) & (ax94x) & (ax93x) & (shiftx0x) & (shiftx1x)) + ((!ax96x) & (ax95x) & (!ax94x) & (!ax93x) & (shiftx0x) & (!shiftx1x)) + ((!ax96x) & (ax95x) & (!ax94x) & (ax93x) & (shiftx0x) & (!shiftx1x)) + ((!ax96x) & (ax95x) & (!ax94x) & (ax93x) & (shiftx0x) & (shiftx1x)) + ((!ax96x) & (ax95x) & (ax94x) & (!ax93x) & (!shiftx0x) & (shiftx1x)) + ((!ax96x) & (ax95x) & (ax94x) & (!ax93x) & (shiftx0x) & (!shiftx1x)) + ((!ax96x) & (ax95x) & (ax94x) & (ax93x) & (!shiftx0x) & (shiftx1x)) + ((!ax96x) & (ax95x) & (ax94x) & (ax93x) & (shiftx0x) & (!shiftx1x)) + ((!ax96x) & (ax95x) & (ax94x) & (ax93x) & (shiftx0x) & (shiftx1x)) + ((ax96x) & (!ax95x) & (!ax94x) & (!ax93x) & (!shiftx0x) & (!shiftx1x)) + ((ax96x) & (!ax95x) & (!ax94x) & (ax93x) & (!shiftx0x) & (!shiftx1x)) + ((ax96x) & (!ax95x) & (!ax94x) & (ax93x) & (shiftx0x) & (shiftx1x)) + ((ax96x) & (!ax95x) & (ax94x) & (!ax93x) & (!shiftx0x) & (!shiftx1x)) + ((ax96x) & (!ax95x) & (ax94x) & (!ax93x) & (!shiftx0x) & (shiftx1x)) + ((ax96x) & (!ax95x) & (ax94x) & (ax93x) & (!shiftx0x) & (!shiftx1x)) + ((ax96x) & (!ax95x) & (ax94x) & (ax93x) & (!shiftx0x) & (shiftx1x)) + ((ax96x) & (!ax95x) & (ax94x) & (ax93x) & (shiftx0x) & (shiftx1x)) + ((ax96x) & (ax95x) & (!ax94x) & (!ax93x) & (!shiftx0x) & (!shiftx1x)) + ((ax96x) & (ax95x) & (!ax94x) & (!ax93x) & (shiftx0x) & (!shiftx1x)) + ((ax96x) & (ax95x) & (!ax94x) & (ax93x) & (!shiftx0x) & (!shiftx1x)) + ((ax96x) & (ax95x) & (!ax94x) & (ax93x) & (shiftx0x) & (!shiftx1x)) + ((ax96x) & (ax95x) & (!ax94x) & (ax93x) & (shiftx0x) & (shiftx1x)) + ((ax96x) & (ax95x) & (ax94x) & (!ax93x) & (!shiftx0x) & (!shiftx1x)) + ((ax96x) & (ax95x) & (ax94x) & (!ax93x) & (!shiftx0x) & (shiftx1x)) + ((ax96x) & (ax95x) & (ax94x) & (!ax93x) & (shiftx0x) & (!shiftx1x)) + ((ax96x) & (ax95x) & (ax94x) & (ax93x) & (!shiftx0x) & (!shiftx1x)) + ((ax96x) & (ax95x) & (ax94x) & (ax93x) & (!shiftx0x) & (shiftx1x)) + ((ax96x) & (ax95x) & (ax94x) & (ax93x) & (shiftx0x) & (!shiftx1x)) + ((ax96x) & (ax95x) & (ax94x) & (ax93x) & (shiftx0x) & (shiftx1x)));
	assign g28 = (((!ax92x) & (!ax91x) & (!ax90x) & (ax89x) & (shiftx0x) & (shiftx1x)) + ((!ax92x) & (!ax91x) & (ax90x) & (!ax89x) & (!shiftx0x) & (shiftx1x)) + ((!ax92x) & (!ax91x) & (ax90x) & (ax89x) & (!shiftx0x) & (shiftx1x)) + ((!ax92x) & (!ax91x) & (ax90x) & (ax89x) & (shiftx0x) & (shiftx1x)) + ((!ax92x) & (ax91x) & (!ax90x) & (!ax89x) & (shiftx0x) & (!shiftx1x)) + ((!ax92x) & (ax91x) & (!ax90x) & (ax89x) & (shiftx0x) & (!shiftx1x)) + ((!ax92x) & (ax91x) & (!ax90x) & (ax89x) & (shiftx0x) & (shiftx1x)) + ((!ax92x) & (ax91x) & (ax90x) & (!ax89x) & (!shiftx0x) & (shiftx1x)) + ((!ax92x) & (ax91x) & (ax90x) & (!ax89x) & (shiftx0x) & (!shiftx1x)) + ((!ax92x) & (ax91x) & (ax90x) & (ax89x) & (!shiftx0x) & (shiftx1x)) + ((!ax92x) & (ax91x) & (ax90x) & (ax89x) & (shiftx0x) & (!shiftx1x)) + ((!ax92x) & (ax91x) & (ax90x) & (ax89x) & (shiftx0x) & (shiftx1x)) + ((ax92x) & (!ax91x) & (!ax90x) & (!ax89x) & (!shiftx0x) & (!shiftx1x)) + ((ax92x) & (!ax91x) & (!ax90x) & (ax89x) & (!shiftx0x) & (!shiftx1x)) + ((ax92x) & (!ax91x) & (!ax90x) & (ax89x) & (shiftx0x) & (shiftx1x)) + ((ax92x) & (!ax91x) & (ax90x) & (!ax89x) & (!shiftx0x) & (!shiftx1x)) + ((ax92x) & (!ax91x) & (ax90x) & (!ax89x) & (!shiftx0x) & (shiftx1x)) + ((ax92x) & (!ax91x) & (ax90x) & (ax89x) & (!shiftx0x) & (!shiftx1x)) + ((ax92x) & (!ax91x) & (ax90x) & (ax89x) & (!shiftx0x) & (shiftx1x)) + ((ax92x) & (!ax91x) & (ax90x) & (ax89x) & (shiftx0x) & (shiftx1x)) + ((ax92x) & (ax91x) & (!ax90x) & (!ax89x) & (!shiftx0x) & (!shiftx1x)) + ((ax92x) & (ax91x) & (!ax90x) & (!ax89x) & (shiftx0x) & (!shiftx1x)) + ((ax92x) & (ax91x) & (!ax90x) & (ax89x) & (!shiftx0x) & (!shiftx1x)) + ((ax92x) & (ax91x) & (!ax90x) & (ax89x) & (shiftx0x) & (!shiftx1x)) + ((ax92x) & (ax91x) & (!ax90x) & (ax89x) & (shiftx0x) & (shiftx1x)) + ((ax92x) & (ax91x) & (ax90x) & (!ax89x) & (!shiftx0x) & (!shiftx1x)) + ((ax92x) & (ax91x) & (ax90x) & (!ax89x) & (!shiftx0x) & (shiftx1x)) + ((ax92x) & (ax91x) & (ax90x) & (!ax89x) & (shiftx0x) & (!shiftx1x)) + ((ax92x) & (ax91x) & (ax90x) & (ax89x) & (!shiftx0x) & (!shiftx1x)) + ((ax92x) & (ax91x) & (ax90x) & (ax89x) & (!shiftx0x) & (shiftx1x)) + ((ax92x) & (ax91x) & (ax90x) & (ax89x) & (shiftx0x) & (!shiftx1x)) + ((ax92x) & (ax91x) & (ax90x) & (ax89x) & (shiftx0x) & (shiftx1x)));
	assign g29 = (((!ax84x) & (!ax83x) & (!ax82x) & (ax81x) & (shiftx0x) & (shiftx1x)) + ((!ax84x) & (!ax83x) & (ax82x) & (!ax81x) & (!shiftx0x) & (shiftx1x)) + ((!ax84x) & (!ax83x) & (ax82x) & (ax81x) & (!shiftx0x) & (shiftx1x)) + ((!ax84x) & (!ax83x) & (ax82x) & (ax81x) & (shiftx0x) & (shiftx1x)) + ((!ax84x) & (ax83x) & (!ax82x) & (!ax81x) & (shiftx0x) & (!shiftx1x)) + ((!ax84x) & (ax83x) & (!ax82x) & (ax81x) & (shiftx0x) & (!shiftx1x)) + ((!ax84x) & (ax83x) & (!ax82x) & (ax81x) & (shiftx0x) & (shiftx1x)) + ((!ax84x) & (ax83x) & (ax82x) & (!ax81x) & (!shiftx0x) & (shiftx1x)) + ((!ax84x) & (ax83x) & (ax82x) & (!ax81x) & (shiftx0x) & (!shiftx1x)) + ((!ax84x) & (ax83x) & (ax82x) & (ax81x) & (!shiftx0x) & (shiftx1x)) + ((!ax84x) & (ax83x) & (ax82x) & (ax81x) & (shiftx0x) & (!shiftx1x)) + ((!ax84x) & (ax83x) & (ax82x) & (ax81x) & (shiftx0x) & (shiftx1x)) + ((ax84x) & (!ax83x) & (!ax82x) & (!ax81x) & (!shiftx0x) & (!shiftx1x)) + ((ax84x) & (!ax83x) & (!ax82x) & (ax81x) & (!shiftx0x) & (!shiftx1x)) + ((ax84x) & (!ax83x) & (!ax82x) & (ax81x) & (shiftx0x) & (shiftx1x)) + ((ax84x) & (!ax83x) & (ax82x) & (!ax81x) & (!shiftx0x) & (!shiftx1x)) + ((ax84x) & (!ax83x) & (ax82x) & (!ax81x) & (!shiftx0x) & (shiftx1x)) + ((ax84x) & (!ax83x) & (ax82x) & (ax81x) & (!shiftx0x) & (!shiftx1x)) + ((ax84x) & (!ax83x) & (ax82x) & (ax81x) & (!shiftx0x) & (shiftx1x)) + ((ax84x) & (!ax83x) & (ax82x) & (ax81x) & (shiftx0x) & (shiftx1x)) + ((ax84x) & (ax83x) & (!ax82x) & (!ax81x) & (!shiftx0x) & (!shiftx1x)) + ((ax84x) & (ax83x) & (!ax82x) & (!ax81x) & (shiftx0x) & (!shiftx1x)) + ((ax84x) & (ax83x) & (!ax82x) & (ax81x) & (!shiftx0x) & (!shiftx1x)) + ((ax84x) & (ax83x) & (!ax82x) & (ax81x) & (shiftx0x) & (!shiftx1x)) + ((ax84x) & (ax83x) & (!ax82x) & (ax81x) & (shiftx0x) & (shiftx1x)) + ((ax84x) & (ax83x) & (ax82x) & (!ax81x) & (!shiftx0x) & (!shiftx1x)) + ((ax84x) & (ax83x) & (ax82x) & (!ax81x) & (!shiftx0x) & (shiftx1x)) + ((ax84x) & (ax83x) & (ax82x) & (!ax81x) & (shiftx0x) & (!shiftx1x)) + ((ax84x) & (ax83x) & (ax82x) & (ax81x) & (!shiftx0x) & (!shiftx1x)) + ((ax84x) & (ax83x) & (ax82x) & (ax81x) & (!shiftx0x) & (shiftx1x)) + ((ax84x) & (ax83x) & (ax82x) & (ax81x) & (shiftx0x) & (!shiftx1x)) + ((ax84x) & (ax83x) & (ax82x) & (ax81x) & (shiftx0x) & (shiftx1x)));
	assign g30 = (((!ax88x) & (!ax87x) & (!ax86x) & (ax85x) & (shiftx0x) & (shiftx1x)) + ((!ax88x) & (!ax87x) & (ax86x) & (!ax85x) & (!shiftx0x) & (shiftx1x)) + ((!ax88x) & (!ax87x) & (ax86x) & (ax85x) & (!shiftx0x) & (shiftx1x)) + ((!ax88x) & (!ax87x) & (ax86x) & (ax85x) & (shiftx0x) & (shiftx1x)) + ((!ax88x) & (ax87x) & (!ax86x) & (!ax85x) & (shiftx0x) & (!shiftx1x)) + ((!ax88x) & (ax87x) & (!ax86x) & (ax85x) & (shiftx0x) & (!shiftx1x)) + ((!ax88x) & (ax87x) & (!ax86x) & (ax85x) & (shiftx0x) & (shiftx1x)) + ((!ax88x) & (ax87x) & (ax86x) & (!ax85x) & (!shiftx0x) & (shiftx1x)) + ((!ax88x) & (ax87x) & (ax86x) & (!ax85x) & (shiftx0x) & (!shiftx1x)) + ((!ax88x) & (ax87x) & (ax86x) & (ax85x) & (!shiftx0x) & (shiftx1x)) + ((!ax88x) & (ax87x) & (ax86x) & (ax85x) & (shiftx0x) & (!shiftx1x)) + ((!ax88x) & (ax87x) & (ax86x) & (ax85x) & (shiftx0x) & (shiftx1x)) + ((ax88x) & (!ax87x) & (!ax86x) & (!ax85x) & (!shiftx0x) & (!shiftx1x)) + ((ax88x) & (!ax87x) & (!ax86x) & (ax85x) & (!shiftx0x) & (!shiftx1x)) + ((ax88x) & (!ax87x) & (!ax86x) & (ax85x) & (shiftx0x) & (shiftx1x)) + ((ax88x) & (!ax87x) & (ax86x) & (!ax85x) & (!shiftx0x) & (!shiftx1x)) + ((ax88x) & (!ax87x) & (ax86x) & (!ax85x) & (!shiftx0x) & (shiftx1x)) + ((ax88x) & (!ax87x) & (ax86x) & (ax85x) & (!shiftx0x) & (!shiftx1x)) + ((ax88x) & (!ax87x) & (ax86x) & (ax85x) & (!shiftx0x) & (shiftx1x)) + ((ax88x) & (!ax87x) & (ax86x) & (ax85x) & (shiftx0x) & (shiftx1x)) + ((ax88x) & (ax87x) & (!ax86x) & (!ax85x) & (!shiftx0x) & (!shiftx1x)) + ((ax88x) & (ax87x) & (!ax86x) & (!ax85x) & (shiftx0x) & (!shiftx1x)) + ((ax88x) & (ax87x) & (!ax86x) & (ax85x) & (!shiftx0x) & (!shiftx1x)) + ((ax88x) & (ax87x) & (!ax86x) & (ax85x) & (shiftx0x) & (!shiftx1x)) + ((ax88x) & (ax87x) & (!ax86x) & (ax85x) & (shiftx0x) & (shiftx1x)) + ((ax88x) & (ax87x) & (ax86x) & (!ax85x) & (!shiftx0x) & (!shiftx1x)) + ((ax88x) & (ax87x) & (ax86x) & (!ax85x) & (!shiftx0x) & (shiftx1x)) + ((ax88x) & (ax87x) & (ax86x) & (!ax85x) & (shiftx0x) & (!shiftx1x)) + ((ax88x) & (ax87x) & (ax86x) & (ax85x) & (!shiftx0x) & (!shiftx1x)) + ((ax88x) & (ax87x) & (ax86x) & (ax85x) & (!shiftx0x) & (shiftx1x)) + ((ax88x) & (ax87x) & (ax86x) & (ax85x) & (shiftx0x) & (!shiftx1x)) + ((ax88x) & (ax87x) & (ax86x) & (ax85x) & (shiftx0x) & (shiftx1x)));
	assign g31 = (((!shiftx2x) & (!shiftx3x) & (g27) & (!g28) & (!g29) & (!g30)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (!g28) & (!g29) & (g30)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (!g28) & (g29) & (!g30)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (!g28) & (g29) & (g30)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (g28) & (!g29) & (!g30)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (g28) & (!g29) & (g30)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (g28) & (g29) & (!g30)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (g28) & (g29) & (g30)) + ((!shiftx2x) & (shiftx3x) & (!g27) & (!g28) & (!g29) & (g30)) + ((!shiftx2x) & (shiftx3x) & (!g27) & (!g28) & (g29) & (g30)) + ((!shiftx2x) & (shiftx3x) & (!g27) & (g28) & (!g29) & (g30)) + ((!shiftx2x) & (shiftx3x) & (!g27) & (g28) & (g29) & (g30)) + ((!shiftx2x) & (shiftx3x) & (g27) & (!g28) & (!g29) & (g30)) + ((!shiftx2x) & (shiftx3x) & (g27) & (!g28) & (g29) & (g30)) + ((!shiftx2x) & (shiftx3x) & (g27) & (g28) & (!g29) & (g30)) + ((!shiftx2x) & (shiftx3x) & (g27) & (g28) & (g29) & (g30)) + ((shiftx2x) & (!shiftx3x) & (!g27) & (g28) & (!g29) & (!g30)) + ((shiftx2x) & (!shiftx3x) & (!g27) & (g28) & (!g29) & (g30)) + ((shiftx2x) & (!shiftx3x) & (!g27) & (g28) & (g29) & (!g30)) + ((shiftx2x) & (!shiftx3x) & (!g27) & (g28) & (g29) & (g30)) + ((shiftx2x) & (!shiftx3x) & (g27) & (g28) & (!g29) & (!g30)) + ((shiftx2x) & (!shiftx3x) & (g27) & (g28) & (!g29) & (g30)) + ((shiftx2x) & (!shiftx3x) & (g27) & (g28) & (g29) & (!g30)) + ((shiftx2x) & (!shiftx3x) & (g27) & (g28) & (g29) & (g30)) + ((shiftx2x) & (shiftx3x) & (!g27) & (!g28) & (g29) & (!g30)) + ((shiftx2x) & (shiftx3x) & (!g27) & (!g28) & (g29) & (g30)) + ((shiftx2x) & (shiftx3x) & (!g27) & (g28) & (g29) & (!g30)) + ((shiftx2x) & (shiftx3x) & (!g27) & (g28) & (g29) & (g30)) + ((shiftx2x) & (shiftx3x) & (g27) & (!g28) & (g29) & (!g30)) + ((shiftx2x) & (shiftx3x) & (g27) & (!g28) & (g29) & (g30)) + ((shiftx2x) & (shiftx3x) & (g27) & (g28) & (g29) & (!g30)) + ((shiftx2x) & (shiftx3x) & (g27) & (g28) & (g29) & (g30)));
	assign g32 = (((!ax0x) & (!ax127x) & (!ax126x) & (ax125x) & (shiftx0x) & (shiftx1x)) + ((!ax0x) & (!ax127x) & (ax126x) & (!ax125x) & (!shiftx0x) & (shiftx1x)) + ((!ax0x) & (!ax127x) & (ax126x) & (ax125x) & (!shiftx0x) & (shiftx1x)) + ((!ax0x) & (!ax127x) & (ax126x) & (ax125x) & (shiftx0x) & (shiftx1x)) + ((!ax0x) & (ax127x) & (!ax126x) & (!ax125x) & (shiftx0x) & (!shiftx1x)) + ((!ax0x) & (ax127x) & (!ax126x) & (ax125x) & (shiftx0x) & (!shiftx1x)) + ((!ax0x) & (ax127x) & (!ax126x) & (ax125x) & (shiftx0x) & (shiftx1x)) + ((!ax0x) & (ax127x) & (ax126x) & (!ax125x) & (!shiftx0x) & (shiftx1x)) + ((!ax0x) & (ax127x) & (ax126x) & (!ax125x) & (shiftx0x) & (!shiftx1x)) + ((!ax0x) & (ax127x) & (ax126x) & (ax125x) & (!shiftx0x) & (shiftx1x)) + ((!ax0x) & (ax127x) & (ax126x) & (ax125x) & (shiftx0x) & (!shiftx1x)) + ((!ax0x) & (ax127x) & (ax126x) & (ax125x) & (shiftx0x) & (shiftx1x)) + ((ax0x) & (!ax127x) & (!ax126x) & (!ax125x) & (!shiftx0x) & (!shiftx1x)) + ((ax0x) & (!ax127x) & (!ax126x) & (ax125x) & (!shiftx0x) & (!shiftx1x)) + ((ax0x) & (!ax127x) & (!ax126x) & (ax125x) & (shiftx0x) & (shiftx1x)) + ((ax0x) & (!ax127x) & (ax126x) & (!ax125x) & (!shiftx0x) & (!shiftx1x)) + ((ax0x) & (!ax127x) & (ax126x) & (!ax125x) & (!shiftx0x) & (shiftx1x)) + ((ax0x) & (!ax127x) & (ax126x) & (ax125x) & (!shiftx0x) & (!shiftx1x)) + ((ax0x) & (!ax127x) & (ax126x) & (ax125x) & (!shiftx0x) & (shiftx1x)) + ((ax0x) & (!ax127x) & (ax126x) & (ax125x) & (shiftx0x) & (shiftx1x)) + ((ax0x) & (ax127x) & (!ax126x) & (!ax125x) & (!shiftx0x) & (!shiftx1x)) + ((ax0x) & (ax127x) & (!ax126x) & (!ax125x) & (shiftx0x) & (!shiftx1x)) + ((ax0x) & (ax127x) & (!ax126x) & (ax125x) & (!shiftx0x) & (!shiftx1x)) + ((ax0x) & (ax127x) & (!ax126x) & (ax125x) & (shiftx0x) & (!shiftx1x)) + ((ax0x) & (ax127x) & (!ax126x) & (ax125x) & (shiftx0x) & (shiftx1x)) + ((ax0x) & (ax127x) & (ax126x) & (!ax125x) & (!shiftx0x) & (!shiftx1x)) + ((ax0x) & (ax127x) & (ax126x) & (!ax125x) & (!shiftx0x) & (shiftx1x)) + ((ax0x) & (ax127x) & (ax126x) & (!ax125x) & (shiftx0x) & (!shiftx1x)) + ((ax0x) & (ax127x) & (ax126x) & (ax125x) & (!shiftx0x) & (!shiftx1x)) + ((ax0x) & (ax127x) & (ax126x) & (ax125x) & (!shiftx0x) & (shiftx1x)) + ((ax0x) & (ax127x) & (ax126x) & (ax125x) & (shiftx0x) & (!shiftx1x)) + ((ax0x) & (ax127x) & (ax126x) & (ax125x) & (shiftx0x) & (shiftx1x)));
	assign g33 = (((!ax124x) & (!ax123x) & (!ax122x) & (ax121x) & (shiftx0x) & (shiftx1x)) + ((!ax124x) & (!ax123x) & (ax122x) & (!ax121x) & (!shiftx0x) & (shiftx1x)) + ((!ax124x) & (!ax123x) & (ax122x) & (ax121x) & (!shiftx0x) & (shiftx1x)) + ((!ax124x) & (!ax123x) & (ax122x) & (ax121x) & (shiftx0x) & (shiftx1x)) + ((!ax124x) & (ax123x) & (!ax122x) & (!ax121x) & (shiftx0x) & (!shiftx1x)) + ((!ax124x) & (ax123x) & (!ax122x) & (ax121x) & (shiftx0x) & (!shiftx1x)) + ((!ax124x) & (ax123x) & (!ax122x) & (ax121x) & (shiftx0x) & (shiftx1x)) + ((!ax124x) & (ax123x) & (ax122x) & (!ax121x) & (!shiftx0x) & (shiftx1x)) + ((!ax124x) & (ax123x) & (ax122x) & (!ax121x) & (shiftx0x) & (!shiftx1x)) + ((!ax124x) & (ax123x) & (ax122x) & (ax121x) & (!shiftx0x) & (shiftx1x)) + ((!ax124x) & (ax123x) & (ax122x) & (ax121x) & (shiftx0x) & (!shiftx1x)) + ((!ax124x) & (ax123x) & (ax122x) & (ax121x) & (shiftx0x) & (shiftx1x)) + ((ax124x) & (!ax123x) & (!ax122x) & (!ax121x) & (!shiftx0x) & (!shiftx1x)) + ((ax124x) & (!ax123x) & (!ax122x) & (ax121x) & (!shiftx0x) & (!shiftx1x)) + ((ax124x) & (!ax123x) & (!ax122x) & (ax121x) & (shiftx0x) & (shiftx1x)) + ((ax124x) & (!ax123x) & (ax122x) & (!ax121x) & (!shiftx0x) & (!shiftx1x)) + ((ax124x) & (!ax123x) & (ax122x) & (!ax121x) & (!shiftx0x) & (shiftx1x)) + ((ax124x) & (!ax123x) & (ax122x) & (ax121x) & (!shiftx0x) & (!shiftx1x)) + ((ax124x) & (!ax123x) & (ax122x) & (ax121x) & (!shiftx0x) & (shiftx1x)) + ((ax124x) & (!ax123x) & (ax122x) & (ax121x) & (shiftx0x) & (shiftx1x)) + ((ax124x) & (ax123x) & (!ax122x) & (!ax121x) & (!shiftx0x) & (!shiftx1x)) + ((ax124x) & (ax123x) & (!ax122x) & (!ax121x) & (shiftx0x) & (!shiftx1x)) + ((ax124x) & (ax123x) & (!ax122x) & (ax121x) & (!shiftx0x) & (!shiftx1x)) + ((ax124x) & (ax123x) & (!ax122x) & (ax121x) & (shiftx0x) & (!shiftx1x)) + ((ax124x) & (ax123x) & (!ax122x) & (ax121x) & (shiftx0x) & (shiftx1x)) + ((ax124x) & (ax123x) & (ax122x) & (!ax121x) & (!shiftx0x) & (!shiftx1x)) + ((ax124x) & (ax123x) & (ax122x) & (!ax121x) & (!shiftx0x) & (shiftx1x)) + ((ax124x) & (ax123x) & (ax122x) & (!ax121x) & (shiftx0x) & (!shiftx1x)) + ((ax124x) & (ax123x) & (ax122x) & (ax121x) & (!shiftx0x) & (!shiftx1x)) + ((ax124x) & (ax123x) & (ax122x) & (ax121x) & (!shiftx0x) & (shiftx1x)) + ((ax124x) & (ax123x) & (ax122x) & (ax121x) & (shiftx0x) & (!shiftx1x)) + ((ax124x) & (ax123x) & (ax122x) & (ax121x) & (shiftx0x) & (shiftx1x)));
	assign g34 = (((!ax116x) & (!ax115x) & (!ax114x) & (ax113x) & (shiftx0x) & (shiftx1x)) + ((!ax116x) & (!ax115x) & (ax114x) & (!ax113x) & (!shiftx0x) & (shiftx1x)) + ((!ax116x) & (!ax115x) & (ax114x) & (ax113x) & (!shiftx0x) & (shiftx1x)) + ((!ax116x) & (!ax115x) & (ax114x) & (ax113x) & (shiftx0x) & (shiftx1x)) + ((!ax116x) & (ax115x) & (!ax114x) & (!ax113x) & (shiftx0x) & (!shiftx1x)) + ((!ax116x) & (ax115x) & (!ax114x) & (ax113x) & (shiftx0x) & (!shiftx1x)) + ((!ax116x) & (ax115x) & (!ax114x) & (ax113x) & (shiftx0x) & (shiftx1x)) + ((!ax116x) & (ax115x) & (ax114x) & (!ax113x) & (!shiftx0x) & (shiftx1x)) + ((!ax116x) & (ax115x) & (ax114x) & (!ax113x) & (shiftx0x) & (!shiftx1x)) + ((!ax116x) & (ax115x) & (ax114x) & (ax113x) & (!shiftx0x) & (shiftx1x)) + ((!ax116x) & (ax115x) & (ax114x) & (ax113x) & (shiftx0x) & (!shiftx1x)) + ((!ax116x) & (ax115x) & (ax114x) & (ax113x) & (shiftx0x) & (shiftx1x)) + ((ax116x) & (!ax115x) & (!ax114x) & (!ax113x) & (!shiftx0x) & (!shiftx1x)) + ((ax116x) & (!ax115x) & (!ax114x) & (ax113x) & (!shiftx0x) & (!shiftx1x)) + ((ax116x) & (!ax115x) & (!ax114x) & (ax113x) & (shiftx0x) & (shiftx1x)) + ((ax116x) & (!ax115x) & (ax114x) & (!ax113x) & (!shiftx0x) & (!shiftx1x)) + ((ax116x) & (!ax115x) & (ax114x) & (!ax113x) & (!shiftx0x) & (shiftx1x)) + ((ax116x) & (!ax115x) & (ax114x) & (ax113x) & (!shiftx0x) & (!shiftx1x)) + ((ax116x) & (!ax115x) & (ax114x) & (ax113x) & (!shiftx0x) & (shiftx1x)) + ((ax116x) & (!ax115x) & (ax114x) & (ax113x) & (shiftx0x) & (shiftx1x)) + ((ax116x) & (ax115x) & (!ax114x) & (!ax113x) & (!shiftx0x) & (!shiftx1x)) + ((ax116x) & (ax115x) & (!ax114x) & (!ax113x) & (shiftx0x) & (!shiftx1x)) + ((ax116x) & (ax115x) & (!ax114x) & (ax113x) & (!shiftx0x) & (!shiftx1x)) + ((ax116x) & (ax115x) & (!ax114x) & (ax113x) & (shiftx0x) & (!shiftx1x)) + ((ax116x) & (ax115x) & (!ax114x) & (ax113x) & (shiftx0x) & (shiftx1x)) + ((ax116x) & (ax115x) & (ax114x) & (!ax113x) & (!shiftx0x) & (!shiftx1x)) + ((ax116x) & (ax115x) & (ax114x) & (!ax113x) & (!shiftx0x) & (shiftx1x)) + ((ax116x) & (ax115x) & (ax114x) & (!ax113x) & (shiftx0x) & (!shiftx1x)) + ((ax116x) & (ax115x) & (ax114x) & (ax113x) & (!shiftx0x) & (!shiftx1x)) + ((ax116x) & (ax115x) & (ax114x) & (ax113x) & (!shiftx0x) & (shiftx1x)) + ((ax116x) & (ax115x) & (ax114x) & (ax113x) & (shiftx0x) & (!shiftx1x)) + ((ax116x) & (ax115x) & (ax114x) & (ax113x) & (shiftx0x) & (shiftx1x)));
	assign g35 = (((!ax120x) & (!ax119x) & (!ax118x) & (ax117x) & (shiftx0x) & (shiftx1x)) + ((!ax120x) & (!ax119x) & (ax118x) & (!ax117x) & (!shiftx0x) & (shiftx1x)) + ((!ax120x) & (!ax119x) & (ax118x) & (ax117x) & (!shiftx0x) & (shiftx1x)) + ((!ax120x) & (!ax119x) & (ax118x) & (ax117x) & (shiftx0x) & (shiftx1x)) + ((!ax120x) & (ax119x) & (!ax118x) & (!ax117x) & (shiftx0x) & (!shiftx1x)) + ((!ax120x) & (ax119x) & (!ax118x) & (ax117x) & (shiftx0x) & (!shiftx1x)) + ((!ax120x) & (ax119x) & (!ax118x) & (ax117x) & (shiftx0x) & (shiftx1x)) + ((!ax120x) & (ax119x) & (ax118x) & (!ax117x) & (!shiftx0x) & (shiftx1x)) + ((!ax120x) & (ax119x) & (ax118x) & (!ax117x) & (shiftx0x) & (!shiftx1x)) + ((!ax120x) & (ax119x) & (ax118x) & (ax117x) & (!shiftx0x) & (shiftx1x)) + ((!ax120x) & (ax119x) & (ax118x) & (ax117x) & (shiftx0x) & (!shiftx1x)) + ((!ax120x) & (ax119x) & (ax118x) & (ax117x) & (shiftx0x) & (shiftx1x)) + ((ax120x) & (!ax119x) & (!ax118x) & (!ax117x) & (!shiftx0x) & (!shiftx1x)) + ((ax120x) & (!ax119x) & (!ax118x) & (ax117x) & (!shiftx0x) & (!shiftx1x)) + ((ax120x) & (!ax119x) & (!ax118x) & (ax117x) & (shiftx0x) & (shiftx1x)) + ((ax120x) & (!ax119x) & (ax118x) & (!ax117x) & (!shiftx0x) & (!shiftx1x)) + ((ax120x) & (!ax119x) & (ax118x) & (!ax117x) & (!shiftx0x) & (shiftx1x)) + ((ax120x) & (!ax119x) & (ax118x) & (ax117x) & (!shiftx0x) & (!shiftx1x)) + ((ax120x) & (!ax119x) & (ax118x) & (ax117x) & (!shiftx0x) & (shiftx1x)) + ((ax120x) & (!ax119x) & (ax118x) & (ax117x) & (shiftx0x) & (shiftx1x)) + ((ax120x) & (ax119x) & (!ax118x) & (!ax117x) & (!shiftx0x) & (!shiftx1x)) + ((ax120x) & (ax119x) & (!ax118x) & (!ax117x) & (shiftx0x) & (!shiftx1x)) + ((ax120x) & (ax119x) & (!ax118x) & (ax117x) & (!shiftx0x) & (!shiftx1x)) + ((ax120x) & (ax119x) & (!ax118x) & (ax117x) & (shiftx0x) & (!shiftx1x)) + ((ax120x) & (ax119x) & (!ax118x) & (ax117x) & (shiftx0x) & (shiftx1x)) + ((ax120x) & (ax119x) & (ax118x) & (!ax117x) & (!shiftx0x) & (!shiftx1x)) + ((ax120x) & (ax119x) & (ax118x) & (!ax117x) & (!shiftx0x) & (shiftx1x)) + ((ax120x) & (ax119x) & (ax118x) & (!ax117x) & (shiftx0x) & (!shiftx1x)) + ((ax120x) & (ax119x) & (ax118x) & (ax117x) & (!shiftx0x) & (!shiftx1x)) + ((ax120x) & (ax119x) & (ax118x) & (ax117x) & (!shiftx0x) & (shiftx1x)) + ((ax120x) & (ax119x) & (ax118x) & (ax117x) & (shiftx0x) & (!shiftx1x)) + ((ax120x) & (ax119x) & (ax118x) & (ax117x) & (shiftx0x) & (shiftx1x)));
	assign g36 = (((!shiftx2x) & (!shiftx3x) & (g32) & (!g33) & (!g34) & (!g35)) + ((!shiftx2x) & (!shiftx3x) & (g32) & (!g33) & (!g34) & (g35)) + ((!shiftx2x) & (!shiftx3x) & (g32) & (!g33) & (g34) & (!g35)) + ((!shiftx2x) & (!shiftx3x) & (g32) & (!g33) & (g34) & (g35)) + ((!shiftx2x) & (!shiftx3x) & (g32) & (g33) & (!g34) & (!g35)) + ((!shiftx2x) & (!shiftx3x) & (g32) & (g33) & (!g34) & (g35)) + ((!shiftx2x) & (!shiftx3x) & (g32) & (g33) & (g34) & (!g35)) + ((!shiftx2x) & (!shiftx3x) & (g32) & (g33) & (g34) & (g35)) + ((!shiftx2x) & (shiftx3x) & (!g32) & (!g33) & (!g34) & (g35)) + ((!shiftx2x) & (shiftx3x) & (!g32) & (!g33) & (g34) & (g35)) + ((!shiftx2x) & (shiftx3x) & (!g32) & (g33) & (!g34) & (g35)) + ((!shiftx2x) & (shiftx3x) & (!g32) & (g33) & (g34) & (g35)) + ((!shiftx2x) & (shiftx3x) & (g32) & (!g33) & (!g34) & (g35)) + ((!shiftx2x) & (shiftx3x) & (g32) & (!g33) & (g34) & (g35)) + ((!shiftx2x) & (shiftx3x) & (g32) & (g33) & (!g34) & (g35)) + ((!shiftx2x) & (shiftx3x) & (g32) & (g33) & (g34) & (g35)) + ((shiftx2x) & (!shiftx3x) & (!g32) & (g33) & (!g34) & (!g35)) + ((shiftx2x) & (!shiftx3x) & (!g32) & (g33) & (!g34) & (g35)) + ((shiftx2x) & (!shiftx3x) & (!g32) & (g33) & (g34) & (!g35)) + ((shiftx2x) & (!shiftx3x) & (!g32) & (g33) & (g34) & (g35)) + ((shiftx2x) & (!shiftx3x) & (g32) & (g33) & (!g34) & (!g35)) + ((shiftx2x) & (!shiftx3x) & (g32) & (g33) & (!g34) & (g35)) + ((shiftx2x) & (!shiftx3x) & (g32) & (g33) & (g34) & (!g35)) + ((shiftx2x) & (!shiftx3x) & (g32) & (g33) & (g34) & (g35)) + ((shiftx2x) & (shiftx3x) & (!g32) & (!g33) & (g34) & (!g35)) + ((shiftx2x) & (shiftx3x) & (!g32) & (!g33) & (g34) & (g35)) + ((shiftx2x) & (shiftx3x) & (!g32) & (g33) & (g34) & (!g35)) + ((shiftx2x) & (shiftx3x) & (!g32) & (g33) & (g34) & (g35)) + ((shiftx2x) & (shiftx3x) & (g32) & (!g33) & (g34) & (!g35)) + ((shiftx2x) & (shiftx3x) & (g32) & (!g33) & (g34) & (g35)) + ((shiftx2x) & (shiftx3x) & (g32) & (g33) & (g34) & (!g35)) + ((shiftx2x) & (shiftx3x) & (g32) & (g33) & (g34) & (g35)));
	assign g37 = (((!ax112x) & (!ax111x) & (!ax110x) & (ax109x) & (shiftx0x) & (shiftx1x)) + ((!ax112x) & (!ax111x) & (ax110x) & (!ax109x) & (!shiftx0x) & (shiftx1x)) + ((!ax112x) & (!ax111x) & (ax110x) & (ax109x) & (!shiftx0x) & (shiftx1x)) + ((!ax112x) & (!ax111x) & (ax110x) & (ax109x) & (shiftx0x) & (shiftx1x)) + ((!ax112x) & (ax111x) & (!ax110x) & (!ax109x) & (shiftx0x) & (!shiftx1x)) + ((!ax112x) & (ax111x) & (!ax110x) & (ax109x) & (shiftx0x) & (!shiftx1x)) + ((!ax112x) & (ax111x) & (!ax110x) & (ax109x) & (shiftx0x) & (shiftx1x)) + ((!ax112x) & (ax111x) & (ax110x) & (!ax109x) & (!shiftx0x) & (shiftx1x)) + ((!ax112x) & (ax111x) & (ax110x) & (!ax109x) & (shiftx0x) & (!shiftx1x)) + ((!ax112x) & (ax111x) & (ax110x) & (ax109x) & (!shiftx0x) & (shiftx1x)) + ((!ax112x) & (ax111x) & (ax110x) & (ax109x) & (shiftx0x) & (!shiftx1x)) + ((!ax112x) & (ax111x) & (ax110x) & (ax109x) & (shiftx0x) & (shiftx1x)) + ((ax112x) & (!ax111x) & (!ax110x) & (!ax109x) & (!shiftx0x) & (!shiftx1x)) + ((ax112x) & (!ax111x) & (!ax110x) & (ax109x) & (!shiftx0x) & (!shiftx1x)) + ((ax112x) & (!ax111x) & (!ax110x) & (ax109x) & (shiftx0x) & (shiftx1x)) + ((ax112x) & (!ax111x) & (ax110x) & (!ax109x) & (!shiftx0x) & (!shiftx1x)) + ((ax112x) & (!ax111x) & (ax110x) & (!ax109x) & (!shiftx0x) & (shiftx1x)) + ((ax112x) & (!ax111x) & (ax110x) & (ax109x) & (!shiftx0x) & (!shiftx1x)) + ((ax112x) & (!ax111x) & (ax110x) & (ax109x) & (!shiftx0x) & (shiftx1x)) + ((ax112x) & (!ax111x) & (ax110x) & (ax109x) & (shiftx0x) & (shiftx1x)) + ((ax112x) & (ax111x) & (!ax110x) & (!ax109x) & (!shiftx0x) & (!shiftx1x)) + ((ax112x) & (ax111x) & (!ax110x) & (!ax109x) & (shiftx0x) & (!shiftx1x)) + ((ax112x) & (ax111x) & (!ax110x) & (ax109x) & (!shiftx0x) & (!shiftx1x)) + ((ax112x) & (ax111x) & (!ax110x) & (ax109x) & (shiftx0x) & (!shiftx1x)) + ((ax112x) & (ax111x) & (!ax110x) & (ax109x) & (shiftx0x) & (shiftx1x)) + ((ax112x) & (ax111x) & (ax110x) & (!ax109x) & (!shiftx0x) & (!shiftx1x)) + ((ax112x) & (ax111x) & (ax110x) & (!ax109x) & (!shiftx0x) & (shiftx1x)) + ((ax112x) & (ax111x) & (ax110x) & (!ax109x) & (shiftx0x) & (!shiftx1x)) + ((ax112x) & (ax111x) & (ax110x) & (ax109x) & (!shiftx0x) & (!shiftx1x)) + ((ax112x) & (ax111x) & (ax110x) & (ax109x) & (!shiftx0x) & (shiftx1x)) + ((ax112x) & (ax111x) & (ax110x) & (ax109x) & (shiftx0x) & (!shiftx1x)) + ((ax112x) & (ax111x) & (ax110x) & (ax109x) & (shiftx0x) & (shiftx1x)));
	assign g38 = (((!ax108x) & (!ax107x) & (!ax106x) & (ax105x) & (shiftx0x) & (shiftx1x)) + ((!ax108x) & (!ax107x) & (ax106x) & (!ax105x) & (!shiftx0x) & (shiftx1x)) + ((!ax108x) & (!ax107x) & (ax106x) & (ax105x) & (!shiftx0x) & (shiftx1x)) + ((!ax108x) & (!ax107x) & (ax106x) & (ax105x) & (shiftx0x) & (shiftx1x)) + ((!ax108x) & (ax107x) & (!ax106x) & (!ax105x) & (shiftx0x) & (!shiftx1x)) + ((!ax108x) & (ax107x) & (!ax106x) & (ax105x) & (shiftx0x) & (!shiftx1x)) + ((!ax108x) & (ax107x) & (!ax106x) & (ax105x) & (shiftx0x) & (shiftx1x)) + ((!ax108x) & (ax107x) & (ax106x) & (!ax105x) & (!shiftx0x) & (shiftx1x)) + ((!ax108x) & (ax107x) & (ax106x) & (!ax105x) & (shiftx0x) & (!shiftx1x)) + ((!ax108x) & (ax107x) & (ax106x) & (ax105x) & (!shiftx0x) & (shiftx1x)) + ((!ax108x) & (ax107x) & (ax106x) & (ax105x) & (shiftx0x) & (!shiftx1x)) + ((!ax108x) & (ax107x) & (ax106x) & (ax105x) & (shiftx0x) & (shiftx1x)) + ((ax108x) & (!ax107x) & (!ax106x) & (!ax105x) & (!shiftx0x) & (!shiftx1x)) + ((ax108x) & (!ax107x) & (!ax106x) & (ax105x) & (!shiftx0x) & (!shiftx1x)) + ((ax108x) & (!ax107x) & (!ax106x) & (ax105x) & (shiftx0x) & (shiftx1x)) + ((ax108x) & (!ax107x) & (ax106x) & (!ax105x) & (!shiftx0x) & (!shiftx1x)) + ((ax108x) & (!ax107x) & (ax106x) & (!ax105x) & (!shiftx0x) & (shiftx1x)) + ((ax108x) & (!ax107x) & (ax106x) & (ax105x) & (!shiftx0x) & (!shiftx1x)) + ((ax108x) & (!ax107x) & (ax106x) & (ax105x) & (!shiftx0x) & (shiftx1x)) + ((ax108x) & (!ax107x) & (ax106x) & (ax105x) & (shiftx0x) & (shiftx1x)) + ((ax108x) & (ax107x) & (!ax106x) & (!ax105x) & (!shiftx0x) & (!shiftx1x)) + ((ax108x) & (ax107x) & (!ax106x) & (!ax105x) & (shiftx0x) & (!shiftx1x)) + ((ax108x) & (ax107x) & (!ax106x) & (ax105x) & (!shiftx0x) & (!shiftx1x)) + ((ax108x) & (ax107x) & (!ax106x) & (ax105x) & (shiftx0x) & (!shiftx1x)) + ((ax108x) & (ax107x) & (!ax106x) & (ax105x) & (shiftx0x) & (shiftx1x)) + ((ax108x) & (ax107x) & (ax106x) & (!ax105x) & (!shiftx0x) & (!shiftx1x)) + ((ax108x) & (ax107x) & (ax106x) & (!ax105x) & (!shiftx0x) & (shiftx1x)) + ((ax108x) & (ax107x) & (ax106x) & (!ax105x) & (shiftx0x) & (!shiftx1x)) + ((ax108x) & (ax107x) & (ax106x) & (ax105x) & (!shiftx0x) & (!shiftx1x)) + ((ax108x) & (ax107x) & (ax106x) & (ax105x) & (!shiftx0x) & (shiftx1x)) + ((ax108x) & (ax107x) & (ax106x) & (ax105x) & (shiftx0x) & (!shiftx1x)) + ((ax108x) & (ax107x) & (ax106x) & (ax105x) & (shiftx0x) & (shiftx1x)));
	assign g39 = (((!ax100x) & (!ax99x) & (!ax98x) & (ax97x) & (shiftx0x) & (shiftx1x)) + ((!ax100x) & (!ax99x) & (ax98x) & (!ax97x) & (!shiftx0x) & (shiftx1x)) + ((!ax100x) & (!ax99x) & (ax98x) & (ax97x) & (!shiftx0x) & (shiftx1x)) + ((!ax100x) & (!ax99x) & (ax98x) & (ax97x) & (shiftx0x) & (shiftx1x)) + ((!ax100x) & (ax99x) & (!ax98x) & (!ax97x) & (shiftx0x) & (!shiftx1x)) + ((!ax100x) & (ax99x) & (!ax98x) & (ax97x) & (shiftx0x) & (!shiftx1x)) + ((!ax100x) & (ax99x) & (!ax98x) & (ax97x) & (shiftx0x) & (shiftx1x)) + ((!ax100x) & (ax99x) & (ax98x) & (!ax97x) & (!shiftx0x) & (shiftx1x)) + ((!ax100x) & (ax99x) & (ax98x) & (!ax97x) & (shiftx0x) & (!shiftx1x)) + ((!ax100x) & (ax99x) & (ax98x) & (ax97x) & (!shiftx0x) & (shiftx1x)) + ((!ax100x) & (ax99x) & (ax98x) & (ax97x) & (shiftx0x) & (!shiftx1x)) + ((!ax100x) & (ax99x) & (ax98x) & (ax97x) & (shiftx0x) & (shiftx1x)) + ((ax100x) & (!ax99x) & (!ax98x) & (!ax97x) & (!shiftx0x) & (!shiftx1x)) + ((ax100x) & (!ax99x) & (!ax98x) & (ax97x) & (!shiftx0x) & (!shiftx1x)) + ((ax100x) & (!ax99x) & (!ax98x) & (ax97x) & (shiftx0x) & (shiftx1x)) + ((ax100x) & (!ax99x) & (ax98x) & (!ax97x) & (!shiftx0x) & (!shiftx1x)) + ((ax100x) & (!ax99x) & (ax98x) & (!ax97x) & (!shiftx0x) & (shiftx1x)) + ((ax100x) & (!ax99x) & (ax98x) & (ax97x) & (!shiftx0x) & (!shiftx1x)) + ((ax100x) & (!ax99x) & (ax98x) & (ax97x) & (!shiftx0x) & (shiftx1x)) + ((ax100x) & (!ax99x) & (ax98x) & (ax97x) & (shiftx0x) & (shiftx1x)) + ((ax100x) & (ax99x) & (!ax98x) & (!ax97x) & (!shiftx0x) & (!shiftx1x)) + ((ax100x) & (ax99x) & (!ax98x) & (!ax97x) & (shiftx0x) & (!shiftx1x)) + ((ax100x) & (ax99x) & (!ax98x) & (ax97x) & (!shiftx0x) & (!shiftx1x)) + ((ax100x) & (ax99x) & (!ax98x) & (ax97x) & (shiftx0x) & (!shiftx1x)) + ((ax100x) & (ax99x) & (!ax98x) & (ax97x) & (shiftx0x) & (shiftx1x)) + ((ax100x) & (ax99x) & (ax98x) & (!ax97x) & (!shiftx0x) & (!shiftx1x)) + ((ax100x) & (ax99x) & (ax98x) & (!ax97x) & (!shiftx0x) & (shiftx1x)) + ((ax100x) & (ax99x) & (ax98x) & (!ax97x) & (shiftx0x) & (!shiftx1x)) + ((ax100x) & (ax99x) & (ax98x) & (ax97x) & (!shiftx0x) & (!shiftx1x)) + ((ax100x) & (ax99x) & (ax98x) & (ax97x) & (!shiftx0x) & (shiftx1x)) + ((ax100x) & (ax99x) & (ax98x) & (ax97x) & (shiftx0x) & (!shiftx1x)) + ((ax100x) & (ax99x) & (ax98x) & (ax97x) & (shiftx0x) & (shiftx1x)));
	assign g40 = (((!ax104x) & (!ax103x) & (!ax102x) & (ax101x) & (shiftx0x) & (shiftx1x)) + ((!ax104x) & (!ax103x) & (ax102x) & (!ax101x) & (!shiftx0x) & (shiftx1x)) + ((!ax104x) & (!ax103x) & (ax102x) & (ax101x) & (!shiftx0x) & (shiftx1x)) + ((!ax104x) & (!ax103x) & (ax102x) & (ax101x) & (shiftx0x) & (shiftx1x)) + ((!ax104x) & (ax103x) & (!ax102x) & (!ax101x) & (shiftx0x) & (!shiftx1x)) + ((!ax104x) & (ax103x) & (!ax102x) & (ax101x) & (shiftx0x) & (!shiftx1x)) + ((!ax104x) & (ax103x) & (!ax102x) & (ax101x) & (shiftx0x) & (shiftx1x)) + ((!ax104x) & (ax103x) & (ax102x) & (!ax101x) & (!shiftx0x) & (shiftx1x)) + ((!ax104x) & (ax103x) & (ax102x) & (!ax101x) & (shiftx0x) & (!shiftx1x)) + ((!ax104x) & (ax103x) & (ax102x) & (ax101x) & (!shiftx0x) & (shiftx1x)) + ((!ax104x) & (ax103x) & (ax102x) & (ax101x) & (shiftx0x) & (!shiftx1x)) + ((!ax104x) & (ax103x) & (ax102x) & (ax101x) & (shiftx0x) & (shiftx1x)) + ((ax104x) & (!ax103x) & (!ax102x) & (!ax101x) & (!shiftx0x) & (!shiftx1x)) + ((ax104x) & (!ax103x) & (!ax102x) & (ax101x) & (!shiftx0x) & (!shiftx1x)) + ((ax104x) & (!ax103x) & (!ax102x) & (ax101x) & (shiftx0x) & (shiftx1x)) + ((ax104x) & (!ax103x) & (ax102x) & (!ax101x) & (!shiftx0x) & (!shiftx1x)) + ((ax104x) & (!ax103x) & (ax102x) & (!ax101x) & (!shiftx0x) & (shiftx1x)) + ((ax104x) & (!ax103x) & (ax102x) & (ax101x) & (!shiftx0x) & (!shiftx1x)) + ((ax104x) & (!ax103x) & (ax102x) & (ax101x) & (!shiftx0x) & (shiftx1x)) + ((ax104x) & (!ax103x) & (ax102x) & (ax101x) & (shiftx0x) & (shiftx1x)) + ((ax104x) & (ax103x) & (!ax102x) & (!ax101x) & (!shiftx0x) & (!shiftx1x)) + ((ax104x) & (ax103x) & (!ax102x) & (!ax101x) & (shiftx0x) & (!shiftx1x)) + ((ax104x) & (ax103x) & (!ax102x) & (ax101x) & (!shiftx0x) & (!shiftx1x)) + ((ax104x) & (ax103x) & (!ax102x) & (ax101x) & (shiftx0x) & (!shiftx1x)) + ((ax104x) & (ax103x) & (!ax102x) & (ax101x) & (shiftx0x) & (shiftx1x)) + ((ax104x) & (ax103x) & (ax102x) & (!ax101x) & (!shiftx0x) & (!shiftx1x)) + ((ax104x) & (ax103x) & (ax102x) & (!ax101x) & (!shiftx0x) & (shiftx1x)) + ((ax104x) & (ax103x) & (ax102x) & (!ax101x) & (shiftx0x) & (!shiftx1x)) + ((ax104x) & (ax103x) & (ax102x) & (ax101x) & (!shiftx0x) & (!shiftx1x)) + ((ax104x) & (ax103x) & (ax102x) & (ax101x) & (!shiftx0x) & (shiftx1x)) + ((ax104x) & (ax103x) & (ax102x) & (ax101x) & (shiftx0x) & (!shiftx1x)) + ((ax104x) & (ax103x) & (ax102x) & (ax101x) & (shiftx0x) & (shiftx1x)));
	assign g41 = (((!shiftx2x) & (!shiftx3x) & (g37) & (!g38) & (!g39) & (!g40)) + ((!shiftx2x) & (!shiftx3x) & (g37) & (!g38) & (!g39) & (g40)) + ((!shiftx2x) & (!shiftx3x) & (g37) & (!g38) & (g39) & (!g40)) + ((!shiftx2x) & (!shiftx3x) & (g37) & (!g38) & (g39) & (g40)) + ((!shiftx2x) & (!shiftx3x) & (g37) & (g38) & (!g39) & (!g40)) + ((!shiftx2x) & (!shiftx3x) & (g37) & (g38) & (!g39) & (g40)) + ((!shiftx2x) & (!shiftx3x) & (g37) & (g38) & (g39) & (!g40)) + ((!shiftx2x) & (!shiftx3x) & (g37) & (g38) & (g39) & (g40)) + ((!shiftx2x) & (shiftx3x) & (!g37) & (!g38) & (!g39) & (g40)) + ((!shiftx2x) & (shiftx3x) & (!g37) & (!g38) & (g39) & (g40)) + ((!shiftx2x) & (shiftx3x) & (!g37) & (g38) & (!g39) & (g40)) + ((!shiftx2x) & (shiftx3x) & (!g37) & (g38) & (g39) & (g40)) + ((!shiftx2x) & (shiftx3x) & (g37) & (!g38) & (!g39) & (g40)) + ((!shiftx2x) & (shiftx3x) & (g37) & (!g38) & (g39) & (g40)) + ((!shiftx2x) & (shiftx3x) & (g37) & (g38) & (!g39) & (g40)) + ((!shiftx2x) & (shiftx3x) & (g37) & (g38) & (g39) & (g40)) + ((shiftx2x) & (!shiftx3x) & (!g37) & (g38) & (!g39) & (!g40)) + ((shiftx2x) & (!shiftx3x) & (!g37) & (g38) & (!g39) & (g40)) + ((shiftx2x) & (!shiftx3x) & (!g37) & (g38) & (g39) & (!g40)) + ((shiftx2x) & (!shiftx3x) & (!g37) & (g38) & (g39) & (g40)) + ((shiftx2x) & (!shiftx3x) & (g37) & (g38) & (!g39) & (!g40)) + ((shiftx2x) & (!shiftx3x) & (g37) & (g38) & (!g39) & (g40)) + ((shiftx2x) & (!shiftx3x) & (g37) & (g38) & (g39) & (!g40)) + ((shiftx2x) & (!shiftx3x) & (g37) & (g38) & (g39) & (g40)) + ((shiftx2x) & (shiftx3x) & (!g37) & (!g38) & (g39) & (!g40)) + ((shiftx2x) & (shiftx3x) & (!g37) & (!g38) & (g39) & (g40)) + ((shiftx2x) & (shiftx3x) & (!g37) & (g38) & (g39) & (!g40)) + ((shiftx2x) & (shiftx3x) & (!g37) & (g38) & (g39) & (g40)) + ((shiftx2x) & (shiftx3x) & (g37) & (!g38) & (g39) & (!g40)) + ((shiftx2x) & (shiftx3x) & (g37) & (!g38) & (g39) & (g40)) + ((shiftx2x) & (shiftx3x) & (g37) & (g38) & (g39) & (!g40)) + ((shiftx2x) & (shiftx3x) & (g37) & (g38) & (g39) & (g40)));
	assign g42 = (((!shiftx4x) & (!shiftx5x) & (!g26) & (!g31) & (g36) & (!g41)) + ((!shiftx4x) & (!shiftx5x) & (!g26) & (!g31) & (g36) & (g41)) + ((!shiftx4x) & (!shiftx5x) & (!g26) & (g31) & (g36) & (!g41)) + ((!shiftx4x) & (!shiftx5x) & (!g26) & (g31) & (g36) & (g41)) + ((!shiftx4x) & (!shiftx5x) & (g26) & (!g31) & (g36) & (!g41)) + ((!shiftx4x) & (!shiftx5x) & (g26) & (!g31) & (g36) & (g41)) + ((!shiftx4x) & (!shiftx5x) & (g26) & (g31) & (g36) & (!g41)) + ((!shiftx4x) & (!shiftx5x) & (g26) & (g31) & (g36) & (g41)) + ((!shiftx4x) & (shiftx5x) & (!g26) & (g31) & (!g36) & (!g41)) + ((!shiftx4x) & (shiftx5x) & (!g26) & (g31) & (!g36) & (g41)) + ((!shiftx4x) & (shiftx5x) & (!g26) & (g31) & (g36) & (!g41)) + ((!shiftx4x) & (shiftx5x) & (!g26) & (g31) & (g36) & (g41)) + ((!shiftx4x) & (shiftx5x) & (g26) & (g31) & (!g36) & (!g41)) + ((!shiftx4x) & (shiftx5x) & (g26) & (g31) & (!g36) & (g41)) + ((!shiftx4x) & (shiftx5x) & (g26) & (g31) & (g36) & (!g41)) + ((!shiftx4x) & (shiftx5x) & (g26) & (g31) & (g36) & (g41)) + ((shiftx4x) & (!shiftx5x) & (!g26) & (!g31) & (!g36) & (g41)) + ((shiftx4x) & (!shiftx5x) & (!g26) & (!g31) & (g36) & (g41)) + ((shiftx4x) & (!shiftx5x) & (!g26) & (g31) & (!g36) & (g41)) + ((shiftx4x) & (!shiftx5x) & (!g26) & (g31) & (g36) & (g41)) + ((shiftx4x) & (!shiftx5x) & (g26) & (!g31) & (!g36) & (g41)) + ((shiftx4x) & (!shiftx5x) & (g26) & (!g31) & (g36) & (g41)) + ((shiftx4x) & (!shiftx5x) & (g26) & (g31) & (!g36) & (g41)) + ((shiftx4x) & (!shiftx5x) & (g26) & (g31) & (g36) & (g41)) + ((shiftx4x) & (shiftx5x) & (g26) & (!g31) & (!g36) & (!g41)) + ((shiftx4x) & (shiftx5x) & (g26) & (!g31) & (!g36) & (g41)) + ((shiftx4x) & (shiftx5x) & (g26) & (!g31) & (g36) & (!g41)) + ((shiftx4x) & (shiftx5x) & (g26) & (!g31) & (g36) & (g41)) + ((shiftx4x) & (shiftx5x) & (g26) & (g31) & (!g36) & (!g41)) + ((shiftx4x) & (shiftx5x) & (g26) & (g31) & (!g36) & (g41)) + ((shiftx4x) & (shiftx5x) & (g26) & (g31) & (g36) & (!g41)) + ((shiftx4x) & (shiftx5x) & (g26) & (g31) & (g36) & (g41)));
	assign resultx0x = (((!sk[42]) & (shiftx6x) & (!g21) & (!g42)) + ((!sk[42]) & (shiftx6x) & (!g21) & (g42)) + ((!sk[42]) & (shiftx6x) & (g21) & (!g42)) + ((!sk[42]) & (shiftx6x) & (g21) & (g42)) + ((sk[42]) & (!shiftx6x) & (!g21) & (g42)) + ((sk[42]) & (!shiftx6x) & (g21) & (g42)) + ((sk[42]) & (shiftx6x) & (g21) & (!g42)) + ((sk[42]) & (shiftx6x) & (g21) & (g42)));
	assign g44 = (((!shiftx0x) & (!shiftx1x) & (!ax64x) & (!ax63x) & (!ax62x) & (ax65x)) + ((!shiftx0x) & (!shiftx1x) & (!ax64x) & (!ax63x) & (ax62x) & (ax65x)) + ((!shiftx0x) & (!shiftx1x) & (!ax64x) & (ax63x) & (!ax62x) & (ax65x)) + ((!shiftx0x) & (!shiftx1x) & (!ax64x) & (ax63x) & (ax62x) & (ax65x)) + ((!shiftx0x) & (!shiftx1x) & (ax64x) & (!ax63x) & (!ax62x) & (ax65x)) + ((!shiftx0x) & (!shiftx1x) & (ax64x) & (!ax63x) & (ax62x) & (ax65x)) + ((!shiftx0x) & (!shiftx1x) & (ax64x) & (ax63x) & (!ax62x) & (ax65x)) + ((!shiftx0x) & (!shiftx1x) & (ax64x) & (ax63x) & (ax62x) & (ax65x)) + ((!shiftx0x) & (shiftx1x) & (!ax64x) & (ax63x) & (!ax62x) & (!ax65x)) + ((!shiftx0x) & (shiftx1x) & (!ax64x) & (ax63x) & (!ax62x) & (ax65x)) + ((!shiftx0x) & (shiftx1x) & (!ax64x) & (ax63x) & (ax62x) & (!ax65x)) + ((!shiftx0x) & (shiftx1x) & (!ax64x) & (ax63x) & (ax62x) & (ax65x)) + ((!shiftx0x) & (shiftx1x) & (ax64x) & (ax63x) & (!ax62x) & (!ax65x)) + ((!shiftx0x) & (shiftx1x) & (ax64x) & (ax63x) & (!ax62x) & (ax65x)) + ((!shiftx0x) & (shiftx1x) & (ax64x) & (ax63x) & (ax62x) & (!ax65x)) + ((!shiftx0x) & (shiftx1x) & (ax64x) & (ax63x) & (ax62x) & (ax65x)) + ((shiftx0x) & (!shiftx1x) & (ax64x) & (!ax63x) & (!ax62x) & (!ax65x)) + ((shiftx0x) & (!shiftx1x) & (ax64x) & (!ax63x) & (!ax62x) & (ax65x)) + ((shiftx0x) & (!shiftx1x) & (ax64x) & (!ax63x) & (ax62x) & (!ax65x)) + ((shiftx0x) & (!shiftx1x) & (ax64x) & (!ax63x) & (ax62x) & (ax65x)) + ((shiftx0x) & (!shiftx1x) & (ax64x) & (ax63x) & (!ax62x) & (!ax65x)) + ((shiftx0x) & (!shiftx1x) & (ax64x) & (ax63x) & (!ax62x) & (ax65x)) + ((shiftx0x) & (!shiftx1x) & (ax64x) & (ax63x) & (ax62x) & (!ax65x)) + ((shiftx0x) & (!shiftx1x) & (ax64x) & (ax63x) & (ax62x) & (ax65x)) + ((shiftx0x) & (shiftx1x) & (!ax64x) & (!ax63x) & (ax62x) & (!ax65x)) + ((shiftx0x) & (shiftx1x) & (!ax64x) & (!ax63x) & (ax62x) & (ax65x)) + ((shiftx0x) & (shiftx1x) & (!ax64x) & (ax63x) & (ax62x) & (!ax65x)) + ((shiftx0x) & (shiftx1x) & (!ax64x) & (ax63x) & (ax62x) & (ax65x)) + ((shiftx0x) & (shiftx1x) & (ax64x) & (!ax63x) & (ax62x) & (!ax65x)) + ((shiftx0x) & (shiftx1x) & (ax64x) & (!ax63x) & (ax62x) & (ax65x)) + ((shiftx0x) & (shiftx1x) & (ax64x) & (ax63x) & (ax62x) & (!ax65x)) + ((shiftx0x) & (shiftx1x) & (ax64x) & (ax63x) & (ax62x) & (ax65x)));
	assign g45 = (((!shiftx0x) & (!shiftx1x) & (ax61x) & (!ax60x) & (!ax59x) & (!ax58x)) + ((!shiftx0x) & (!shiftx1x) & (ax61x) & (!ax60x) & (!ax59x) & (ax58x)) + ((!shiftx0x) & (!shiftx1x) & (ax61x) & (!ax60x) & (ax59x) & (!ax58x)) + ((!shiftx0x) & (!shiftx1x) & (ax61x) & (!ax60x) & (ax59x) & (ax58x)) + ((!shiftx0x) & (!shiftx1x) & (ax61x) & (ax60x) & (!ax59x) & (!ax58x)) + ((!shiftx0x) & (!shiftx1x) & (ax61x) & (ax60x) & (!ax59x) & (ax58x)) + ((!shiftx0x) & (!shiftx1x) & (ax61x) & (ax60x) & (ax59x) & (!ax58x)) + ((!shiftx0x) & (!shiftx1x) & (ax61x) & (ax60x) & (ax59x) & (ax58x)) + ((!shiftx0x) & (shiftx1x) & (!ax61x) & (!ax60x) & (ax59x) & (!ax58x)) + ((!shiftx0x) & (shiftx1x) & (!ax61x) & (!ax60x) & (ax59x) & (ax58x)) + ((!shiftx0x) & (shiftx1x) & (!ax61x) & (ax60x) & (ax59x) & (!ax58x)) + ((!shiftx0x) & (shiftx1x) & (!ax61x) & (ax60x) & (ax59x) & (ax58x)) + ((!shiftx0x) & (shiftx1x) & (ax61x) & (!ax60x) & (ax59x) & (!ax58x)) + ((!shiftx0x) & (shiftx1x) & (ax61x) & (!ax60x) & (ax59x) & (ax58x)) + ((!shiftx0x) & (shiftx1x) & (ax61x) & (ax60x) & (ax59x) & (!ax58x)) + ((!shiftx0x) & (shiftx1x) & (ax61x) & (ax60x) & (ax59x) & (ax58x)) + ((shiftx0x) & (!shiftx1x) & (!ax61x) & (ax60x) & (!ax59x) & (!ax58x)) + ((shiftx0x) & (!shiftx1x) & (!ax61x) & (ax60x) & (!ax59x) & (ax58x)) + ((shiftx0x) & (!shiftx1x) & (!ax61x) & (ax60x) & (ax59x) & (!ax58x)) + ((shiftx0x) & (!shiftx1x) & (!ax61x) & (ax60x) & (ax59x) & (ax58x)) + ((shiftx0x) & (!shiftx1x) & (ax61x) & (ax60x) & (!ax59x) & (!ax58x)) + ((shiftx0x) & (!shiftx1x) & (ax61x) & (ax60x) & (!ax59x) & (ax58x)) + ((shiftx0x) & (!shiftx1x) & (ax61x) & (ax60x) & (ax59x) & (!ax58x)) + ((shiftx0x) & (!shiftx1x) & (ax61x) & (ax60x) & (ax59x) & (ax58x)) + ((shiftx0x) & (shiftx1x) & (!ax61x) & (!ax60x) & (!ax59x) & (ax58x)) + ((shiftx0x) & (shiftx1x) & (!ax61x) & (!ax60x) & (ax59x) & (ax58x)) + ((shiftx0x) & (shiftx1x) & (!ax61x) & (ax60x) & (!ax59x) & (ax58x)) + ((shiftx0x) & (shiftx1x) & (!ax61x) & (ax60x) & (ax59x) & (ax58x)) + ((shiftx0x) & (shiftx1x) & (ax61x) & (!ax60x) & (!ax59x) & (ax58x)) + ((shiftx0x) & (shiftx1x) & (ax61x) & (!ax60x) & (ax59x) & (ax58x)) + ((shiftx0x) & (shiftx1x) & (ax61x) & (ax60x) & (!ax59x) & (ax58x)) + ((shiftx0x) & (shiftx1x) & (ax61x) & (ax60x) & (ax59x) & (ax58x)));
	assign g46 = (((!shiftx0x) & (!shiftx1x) & (!ax52x) & (!ax51x) & (!ax50x) & (ax53x)) + ((!shiftx0x) & (!shiftx1x) & (!ax52x) & (!ax51x) & (ax50x) & (ax53x)) + ((!shiftx0x) & (!shiftx1x) & (!ax52x) & (ax51x) & (!ax50x) & (ax53x)) + ((!shiftx0x) & (!shiftx1x) & (!ax52x) & (ax51x) & (ax50x) & (ax53x)) + ((!shiftx0x) & (!shiftx1x) & (ax52x) & (!ax51x) & (!ax50x) & (ax53x)) + ((!shiftx0x) & (!shiftx1x) & (ax52x) & (!ax51x) & (ax50x) & (ax53x)) + ((!shiftx0x) & (!shiftx1x) & (ax52x) & (ax51x) & (!ax50x) & (ax53x)) + ((!shiftx0x) & (!shiftx1x) & (ax52x) & (ax51x) & (ax50x) & (ax53x)) + ((!shiftx0x) & (shiftx1x) & (!ax52x) & (ax51x) & (!ax50x) & (!ax53x)) + ((!shiftx0x) & (shiftx1x) & (!ax52x) & (ax51x) & (!ax50x) & (ax53x)) + ((!shiftx0x) & (shiftx1x) & (!ax52x) & (ax51x) & (ax50x) & (!ax53x)) + ((!shiftx0x) & (shiftx1x) & (!ax52x) & (ax51x) & (ax50x) & (ax53x)) + ((!shiftx0x) & (shiftx1x) & (ax52x) & (ax51x) & (!ax50x) & (!ax53x)) + ((!shiftx0x) & (shiftx1x) & (ax52x) & (ax51x) & (!ax50x) & (ax53x)) + ((!shiftx0x) & (shiftx1x) & (ax52x) & (ax51x) & (ax50x) & (!ax53x)) + ((!shiftx0x) & (shiftx1x) & (ax52x) & (ax51x) & (ax50x) & (ax53x)) + ((shiftx0x) & (!shiftx1x) & (ax52x) & (!ax51x) & (!ax50x) & (!ax53x)) + ((shiftx0x) & (!shiftx1x) & (ax52x) & (!ax51x) & (!ax50x) & (ax53x)) + ((shiftx0x) & (!shiftx1x) & (ax52x) & (!ax51x) & (ax50x) & (!ax53x)) + ((shiftx0x) & (!shiftx1x) & (ax52x) & (!ax51x) & (ax50x) & (ax53x)) + ((shiftx0x) & (!shiftx1x) & (ax52x) & (ax51x) & (!ax50x) & (!ax53x)) + ((shiftx0x) & (!shiftx1x) & (ax52x) & (ax51x) & (!ax50x) & (ax53x)) + ((shiftx0x) & (!shiftx1x) & (ax52x) & (ax51x) & (ax50x) & (!ax53x)) + ((shiftx0x) & (!shiftx1x) & (ax52x) & (ax51x) & (ax50x) & (ax53x)) + ((shiftx0x) & (shiftx1x) & (!ax52x) & (!ax51x) & (ax50x) & (!ax53x)) + ((shiftx0x) & (shiftx1x) & (!ax52x) & (!ax51x) & (ax50x) & (ax53x)) + ((shiftx0x) & (shiftx1x) & (!ax52x) & (ax51x) & (ax50x) & (!ax53x)) + ((shiftx0x) & (shiftx1x) & (!ax52x) & (ax51x) & (ax50x) & (ax53x)) + ((shiftx0x) & (shiftx1x) & (ax52x) & (!ax51x) & (ax50x) & (!ax53x)) + ((shiftx0x) & (shiftx1x) & (ax52x) & (!ax51x) & (ax50x) & (ax53x)) + ((shiftx0x) & (shiftx1x) & (ax52x) & (ax51x) & (ax50x) & (!ax53x)) + ((shiftx0x) & (shiftx1x) & (ax52x) & (ax51x) & (ax50x) & (ax53x)));
	assign g47 = (((!shiftx0x) & (!shiftx1x) & (ax57x) & (!ax56x) & (!ax55x) & (!ax54x)) + ((!shiftx0x) & (!shiftx1x) & (ax57x) & (!ax56x) & (!ax55x) & (ax54x)) + ((!shiftx0x) & (!shiftx1x) & (ax57x) & (!ax56x) & (ax55x) & (!ax54x)) + ((!shiftx0x) & (!shiftx1x) & (ax57x) & (!ax56x) & (ax55x) & (ax54x)) + ((!shiftx0x) & (!shiftx1x) & (ax57x) & (ax56x) & (!ax55x) & (!ax54x)) + ((!shiftx0x) & (!shiftx1x) & (ax57x) & (ax56x) & (!ax55x) & (ax54x)) + ((!shiftx0x) & (!shiftx1x) & (ax57x) & (ax56x) & (ax55x) & (!ax54x)) + ((!shiftx0x) & (!shiftx1x) & (ax57x) & (ax56x) & (ax55x) & (ax54x)) + ((!shiftx0x) & (shiftx1x) & (!ax57x) & (!ax56x) & (ax55x) & (!ax54x)) + ((!shiftx0x) & (shiftx1x) & (!ax57x) & (!ax56x) & (ax55x) & (ax54x)) + ((!shiftx0x) & (shiftx1x) & (!ax57x) & (ax56x) & (ax55x) & (!ax54x)) + ((!shiftx0x) & (shiftx1x) & (!ax57x) & (ax56x) & (ax55x) & (ax54x)) + ((!shiftx0x) & (shiftx1x) & (ax57x) & (!ax56x) & (ax55x) & (!ax54x)) + ((!shiftx0x) & (shiftx1x) & (ax57x) & (!ax56x) & (ax55x) & (ax54x)) + ((!shiftx0x) & (shiftx1x) & (ax57x) & (ax56x) & (ax55x) & (!ax54x)) + ((!shiftx0x) & (shiftx1x) & (ax57x) & (ax56x) & (ax55x) & (ax54x)) + ((shiftx0x) & (!shiftx1x) & (!ax57x) & (ax56x) & (!ax55x) & (!ax54x)) + ((shiftx0x) & (!shiftx1x) & (!ax57x) & (ax56x) & (!ax55x) & (ax54x)) + ((shiftx0x) & (!shiftx1x) & (!ax57x) & (ax56x) & (ax55x) & (!ax54x)) + ((shiftx0x) & (!shiftx1x) & (!ax57x) & (ax56x) & (ax55x) & (ax54x)) + ((shiftx0x) & (!shiftx1x) & (ax57x) & (ax56x) & (!ax55x) & (!ax54x)) + ((shiftx0x) & (!shiftx1x) & (ax57x) & (ax56x) & (!ax55x) & (ax54x)) + ((shiftx0x) & (!shiftx1x) & (ax57x) & (ax56x) & (ax55x) & (!ax54x)) + ((shiftx0x) & (!shiftx1x) & (ax57x) & (ax56x) & (ax55x) & (ax54x)) + ((shiftx0x) & (shiftx1x) & (!ax57x) & (!ax56x) & (!ax55x) & (ax54x)) + ((shiftx0x) & (shiftx1x) & (!ax57x) & (!ax56x) & (ax55x) & (ax54x)) + ((shiftx0x) & (shiftx1x) & (!ax57x) & (ax56x) & (!ax55x) & (ax54x)) + ((shiftx0x) & (shiftx1x) & (!ax57x) & (ax56x) & (ax55x) & (ax54x)) + ((shiftx0x) & (shiftx1x) & (ax57x) & (!ax56x) & (!ax55x) & (ax54x)) + ((shiftx0x) & (shiftx1x) & (ax57x) & (!ax56x) & (ax55x) & (ax54x)) + ((shiftx0x) & (shiftx1x) & (ax57x) & (ax56x) & (!ax55x) & (ax54x)) + ((shiftx0x) & (shiftx1x) & (ax57x) & (ax56x) & (ax55x) & (ax54x)));
	assign g48 = (((!shiftx2x) & (!shiftx3x) & (g44) & (!g45) & (!g46) & (!g47)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (!g45) & (!g46) & (g47)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (!g45) & (g46) & (!g47)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (!g45) & (g46) & (g47)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (g45) & (!g46) & (!g47)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (g45) & (!g46) & (g47)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (g45) & (g46) & (!g47)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (g45) & (g46) & (g47)) + ((!shiftx2x) & (shiftx3x) & (!g44) & (!g45) & (!g46) & (g47)) + ((!shiftx2x) & (shiftx3x) & (!g44) & (!g45) & (g46) & (g47)) + ((!shiftx2x) & (shiftx3x) & (!g44) & (g45) & (!g46) & (g47)) + ((!shiftx2x) & (shiftx3x) & (!g44) & (g45) & (g46) & (g47)) + ((!shiftx2x) & (shiftx3x) & (g44) & (!g45) & (!g46) & (g47)) + ((!shiftx2x) & (shiftx3x) & (g44) & (!g45) & (g46) & (g47)) + ((!shiftx2x) & (shiftx3x) & (g44) & (g45) & (!g46) & (g47)) + ((!shiftx2x) & (shiftx3x) & (g44) & (g45) & (g46) & (g47)) + ((shiftx2x) & (!shiftx3x) & (!g44) & (g45) & (!g46) & (!g47)) + ((shiftx2x) & (!shiftx3x) & (!g44) & (g45) & (!g46) & (g47)) + ((shiftx2x) & (!shiftx3x) & (!g44) & (g45) & (g46) & (!g47)) + ((shiftx2x) & (!shiftx3x) & (!g44) & (g45) & (g46) & (g47)) + ((shiftx2x) & (!shiftx3x) & (g44) & (g45) & (!g46) & (!g47)) + ((shiftx2x) & (!shiftx3x) & (g44) & (g45) & (!g46) & (g47)) + ((shiftx2x) & (!shiftx3x) & (g44) & (g45) & (g46) & (!g47)) + ((shiftx2x) & (!shiftx3x) & (g44) & (g45) & (g46) & (g47)) + ((shiftx2x) & (shiftx3x) & (!g44) & (!g45) & (g46) & (!g47)) + ((shiftx2x) & (shiftx3x) & (!g44) & (!g45) & (g46) & (g47)) + ((shiftx2x) & (shiftx3x) & (!g44) & (g45) & (g46) & (!g47)) + ((shiftx2x) & (shiftx3x) & (!g44) & (g45) & (g46) & (g47)) + ((shiftx2x) & (shiftx3x) & (g44) & (!g45) & (g46) & (!g47)) + ((shiftx2x) & (shiftx3x) & (g44) & (!g45) & (g46) & (g47)) + ((shiftx2x) & (shiftx3x) & (g44) & (g45) & (g46) & (!g47)) + ((shiftx2x) & (shiftx3x) & (g44) & (g45) & (g46) & (g47)));
	assign g49 = (((!ax16x) & (!ax15x) & (!ax14x) & (!shiftx0x) & (!shiftx1x) & (ax17x)) + ((!ax16x) & (!ax15x) & (ax14x) & (!shiftx0x) & (!shiftx1x) & (ax17x)) + ((!ax16x) & (!ax15x) & (ax14x) & (shiftx0x) & (shiftx1x) & (!ax17x)) + ((!ax16x) & (!ax15x) & (ax14x) & (shiftx0x) & (shiftx1x) & (ax17x)) + ((!ax16x) & (ax15x) & (!ax14x) & (!shiftx0x) & (!shiftx1x) & (ax17x)) + ((!ax16x) & (ax15x) & (!ax14x) & (!shiftx0x) & (shiftx1x) & (!ax17x)) + ((!ax16x) & (ax15x) & (!ax14x) & (!shiftx0x) & (shiftx1x) & (ax17x)) + ((!ax16x) & (ax15x) & (ax14x) & (!shiftx0x) & (!shiftx1x) & (ax17x)) + ((!ax16x) & (ax15x) & (ax14x) & (!shiftx0x) & (shiftx1x) & (!ax17x)) + ((!ax16x) & (ax15x) & (ax14x) & (!shiftx0x) & (shiftx1x) & (ax17x)) + ((!ax16x) & (ax15x) & (ax14x) & (shiftx0x) & (shiftx1x) & (!ax17x)) + ((!ax16x) & (ax15x) & (ax14x) & (shiftx0x) & (shiftx1x) & (ax17x)) + ((ax16x) & (!ax15x) & (!ax14x) & (!shiftx0x) & (!shiftx1x) & (ax17x)) + ((ax16x) & (!ax15x) & (!ax14x) & (shiftx0x) & (!shiftx1x) & (!ax17x)) + ((ax16x) & (!ax15x) & (!ax14x) & (shiftx0x) & (!shiftx1x) & (ax17x)) + ((ax16x) & (!ax15x) & (ax14x) & (!shiftx0x) & (!shiftx1x) & (ax17x)) + ((ax16x) & (!ax15x) & (ax14x) & (shiftx0x) & (!shiftx1x) & (!ax17x)) + ((ax16x) & (!ax15x) & (ax14x) & (shiftx0x) & (!shiftx1x) & (ax17x)) + ((ax16x) & (!ax15x) & (ax14x) & (shiftx0x) & (shiftx1x) & (!ax17x)) + ((ax16x) & (!ax15x) & (ax14x) & (shiftx0x) & (shiftx1x) & (ax17x)) + ((ax16x) & (ax15x) & (!ax14x) & (!shiftx0x) & (!shiftx1x) & (ax17x)) + ((ax16x) & (ax15x) & (!ax14x) & (!shiftx0x) & (shiftx1x) & (!ax17x)) + ((ax16x) & (ax15x) & (!ax14x) & (!shiftx0x) & (shiftx1x) & (ax17x)) + ((ax16x) & (ax15x) & (!ax14x) & (shiftx0x) & (!shiftx1x) & (!ax17x)) + ((ax16x) & (ax15x) & (!ax14x) & (shiftx0x) & (!shiftx1x) & (ax17x)) + ((ax16x) & (ax15x) & (ax14x) & (!shiftx0x) & (!shiftx1x) & (ax17x)) + ((ax16x) & (ax15x) & (ax14x) & (!shiftx0x) & (shiftx1x) & (!ax17x)) + ((ax16x) & (ax15x) & (ax14x) & (!shiftx0x) & (shiftx1x) & (ax17x)) + ((ax16x) & (ax15x) & (ax14x) & (shiftx0x) & (!shiftx1x) & (!ax17x)) + ((ax16x) & (ax15x) & (ax14x) & (shiftx0x) & (!shiftx1x) & (ax17x)) + ((ax16x) & (ax15x) & (ax14x) & (shiftx0x) & (shiftx1x) & (!ax17x)) + ((ax16x) & (ax15x) & (ax14x) & (shiftx0x) & (shiftx1x) & (ax17x)));
	assign g50 = (((!ax13x) & (!shiftx0x) & (shiftx1x) & (!ax12x) & (ax11x) & (!ax10x)) + ((!ax13x) & (!shiftx0x) & (shiftx1x) & (!ax12x) & (ax11x) & (ax10x)) + ((!ax13x) & (!shiftx0x) & (shiftx1x) & (ax12x) & (ax11x) & (!ax10x)) + ((!ax13x) & (!shiftx0x) & (shiftx1x) & (ax12x) & (ax11x) & (ax10x)) + ((!ax13x) & (shiftx0x) & (!shiftx1x) & (ax12x) & (!ax11x) & (!ax10x)) + ((!ax13x) & (shiftx0x) & (!shiftx1x) & (ax12x) & (!ax11x) & (ax10x)) + ((!ax13x) & (shiftx0x) & (!shiftx1x) & (ax12x) & (ax11x) & (!ax10x)) + ((!ax13x) & (shiftx0x) & (!shiftx1x) & (ax12x) & (ax11x) & (ax10x)) + ((!ax13x) & (shiftx0x) & (shiftx1x) & (!ax12x) & (!ax11x) & (ax10x)) + ((!ax13x) & (shiftx0x) & (shiftx1x) & (!ax12x) & (ax11x) & (ax10x)) + ((!ax13x) & (shiftx0x) & (shiftx1x) & (ax12x) & (!ax11x) & (ax10x)) + ((!ax13x) & (shiftx0x) & (shiftx1x) & (ax12x) & (ax11x) & (ax10x)) + ((ax13x) & (!shiftx0x) & (!shiftx1x) & (!ax12x) & (!ax11x) & (!ax10x)) + ((ax13x) & (!shiftx0x) & (!shiftx1x) & (!ax12x) & (!ax11x) & (ax10x)) + ((ax13x) & (!shiftx0x) & (!shiftx1x) & (!ax12x) & (ax11x) & (!ax10x)) + ((ax13x) & (!shiftx0x) & (!shiftx1x) & (!ax12x) & (ax11x) & (ax10x)) + ((ax13x) & (!shiftx0x) & (!shiftx1x) & (ax12x) & (!ax11x) & (!ax10x)) + ((ax13x) & (!shiftx0x) & (!shiftx1x) & (ax12x) & (!ax11x) & (ax10x)) + ((ax13x) & (!shiftx0x) & (!shiftx1x) & (ax12x) & (ax11x) & (!ax10x)) + ((ax13x) & (!shiftx0x) & (!shiftx1x) & (ax12x) & (ax11x) & (ax10x)) + ((ax13x) & (!shiftx0x) & (shiftx1x) & (!ax12x) & (ax11x) & (!ax10x)) + ((ax13x) & (!shiftx0x) & (shiftx1x) & (!ax12x) & (ax11x) & (ax10x)) + ((ax13x) & (!shiftx0x) & (shiftx1x) & (ax12x) & (ax11x) & (!ax10x)) + ((ax13x) & (!shiftx0x) & (shiftx1x) & (ax12x) & (ax11x) & (ax10x)) + ((ax13x) & (shiftx0x) & (!shiftx1x) & (ax12x) & (!ax11x) & (!ax10x)) + ((ax13x) & (shiftx0x) & (!shiftx1x) & (ax12x) & (!ax11x) & (ax10x)) + ((ax13x) & (shiftx0x) & (!shiftx1x) & (ax12x) & (ax11x) & (!ax10x)) + ((ax13x) & (shiftx0x) & (!shiftx1x) & (ax12x) & (ax11x) & (ax10x)) + ((ax13x) & (shiftx0x) & (shiftx1x) & (!ax12x) & (!ax11x) & (ax10x)) + ((ax13x) & (shiftx0x) & (shiftx1x) & (!ax12x) & (ax11x) & (ax10x)) + ((ax13x) & (shiftx0x) & (shiftx1x) & (ax12x) & (!ax11x) & (ax10x)) + ((ax13x) & (shiftx0x) & (shiftx1x) & (ax12x) & (ax11x) & (ax10x)));
	assign g51 = (((!shiftx0x) & (!shiftx1x) & (!ax4x) & (!ax3x) & (!ax2x) & (ax5x)) + ((!shiftx0x) & (!shiftx1x) & (!ax4x) & (!ax3x) & (ax2x) & (ax5x)) + ((!shiftx0x) & (!shiftx1x) & (!ax4x) & (ax3x) & (!ax2x) & (ax5x)) + ((!shiftx0x) & (!shiftx1x) & (!ax4x) & (ax3x) & (ax2x) & (ax5x)) + ((!shiftx0x) & (!shiftx1x) & (ax4x) & (!ax3x) & (!ax2x) & (ax5x)) + ((!shiftx0x) & (!shiftx1x) & (ax4x) & (!ax3x) & (ax2x) & (ax5x)) + ((!shiftx0x) & (!shiftx1x) & (ax4x) & (ax3x) & (!ax2x) & (ax5x)) + ((!shiftx0x) & (!shiftx1x) & (ax4x) & (ax3x) & (ax2x) & (ax5x)) + ((!shiftx0x) & (shiftx1x) & (!ax4x) & (ax3x) & (!ax2x) & (!ax5x)) + ((!shiftx0x) & (shiftx1x) & (!ax4x) & (ax3x) & (!ax2x) & (ax5x)) + ((!shiftx0x) & (shiftx1x) & (!ax4x) & (ax3x) & (ax2x) & (!ax5x)) + ((!shiftx0x) & (shiftx1x) & (!ax4x) & (ax3x) & (ax2x) & (ax5x)) + ((!shiftx0x) & (shiftx1x) & (ax4x) & (ax3x) & (!ax2x) & (!ax5x)) + ((!shiftx0x) & (shiftx1x) & (ax4x) & (ax3x) & (!ax2x) & (ax5x)) + ((!shiftx0x) & (shiftx1x) & (ax4x) & (ax3x) & (ax2x) & (!ax5x)) + ((!shiftx0x) & (shiftx1x) & (ax4x) & (ax3x) & (ax2x) & (ax5x)) + ((shiftx0x) & (!shiftx1x) & (ax4x) & (!ax3x) & (!ax2x) & (!ax5x)) + ((shiftx0x) & (!shiftx1x) & (ax4x) & (!ax3x) & (!ax2x) & (ax5x)) + ((shiftx0x) & (!shiftx1x) & (ax4x) & (!ax3x) & (ax2x) & (!ax5x)) + ((shiftx0x) & (!shiftx1x) & (ax4x) & (!ax3x) & (ax2x) & (ax5x)) + ((shiftx0x) & (!shiftx1x) & (ax4x) & (ax3x) & (!ax2x) & (!ax5x)) + ((shiftx0x) & (!shiftx1x) & (ax4x) & (ax3x) & (!ax2x) & (ax5x)) + ((shiftx0x) & (!shiftx1x) & (ax4x) & (ax3x) & (ax2x) & (!ax5x)) + ((shiftx0x) & (!shiftx1x) & (ax4x) & (ax3x) & (ax2x) & (ax5x)) + ((shiftx0x) & (shiftx1x) & (!ax4x) & (!ax3x) & (ax2x) & (!ax5x)) + ((shiftx0x) & (shiftx1x) & (!ax4x) & (!ax3x) & (ax2x) & (ax5x)) + ((shiftx0x) & (shiftx1x) & (!ax4x) & (ax3x) & (ax2x) & (!ax5x)) + ((shiftx0x) & (shiftx1x) & (!ax4x) & (ax3x) & (ax2x) & (ax5x)) + ((shiftx0x) & (shiftx1x) & (ax4x) & (!ax3x) & (ax2x) & (!ax5x)) + ((shiftx0x) & (shiftx1x) & (ax4x) & (!ax3x) & (ax2x) & (ax5x)) + ((shiftx0x) & (shiftx1x) & (ax4x) & (ax3x) & (ax2x) & (!ax5x)) + ((shiftx0x) & (shiftx1x) & (ax4x) & (ax3x) & (ax2x) & (ax5x)));
	assign g52 = (((!shiftx0x) & (!shiftx1x) & (ax9x) & (!ax8x) & (!ax7x) & (!ax6x)) + ((!shiftx0x) & (!shiftx1x) & (ax9x) & (!ax8x) & (!ax7x) & (ax6x)) + ((!shiftx0x) & (!shiftx1x) & (ax9x) & (!ax8x) & (ax7x) & (!ax6x)) + ((!shiftx0x) & (!shiftx1x) & (ax9x) & (!ax8x) & (ax7x) & (ax6x)) + ((!shiftx0x) & (!shiftx1x) & (ax9x) & (ax8x) & (!ax7x) & (!ax6x)) + ((!shiftx0x) & (!shiftx1x) & (ax9x) & (ax8x) & (!ax7x) & (ax6x)) + ((!shiftx0x) & (!shiftx1x) & (ax9x) & (ax8x) & (ax7x) & (!ax6x)) + ((!shiftx0x) & (!shiftx1x) & (ax9x) & (ax8x) & (ax7x) & (ax6x)) + ((!shiftx0x) & (shiftx1x) & (!ax9x) & (!ax8x) & (ax7x) & (!ax6x)) + ((!shiftx0x) & (shiftx1x) & (!ax9x) & (!ax8x) & (ax7x) & (ax6x)) + ((!shiftx0x) & (shiftx1x) & (!ax9x) & (ax8x) & (ax7x) & (!ax6x)) + ((!shiftx0x) & (shiftx1x) & (!ax9x) & (ax8x) & (ax7x) & (ax6x)) + ((!shiftx0x) & (shiftx1x) & (ax9x) & (!ax8x) & (ax7x) & (!ax6x)) + ((!shiftx0x) & (shiftx1x) & (ax9x) & (!ax8x) & (ax7x) & (ax6x)) + ((!shiftx0x) & (shiftx1x) & (ax9x) & (ax8x) & (ax7x) & (!ax6x)) + ((!shiftx0x) & (shiftx1x) & (ax9x) & (ax8x) & (ax7x) & (ax6x)) + ((shiftx0x) & (!shiftx1x) & (!ax9x) & (ax8x) & (!ax7x) & (!ax6x)) + ((shiftx0x) & (!shiftx1x) & (!ax9x) & (ax8x) & (!ax7x) & (ax6x)) + ((shiftx0x) & (!shiftx1x) & (!ax9x) & (ax8x) & (ax7x) & (!ax6x)) + ((shiftx0x) & (!shiftx1x) & (!ax9x) & (ax8x) & (ax7x) & (ax6x)) + ((shiftx0x) & (!shiftx1x) & (ax9x) & (ax8x) & (!ax7x) & (!ax6x)) + ((shiftx0x) & (!shiftx1x) & (ax9x) & (ax8x) & (!ax7x) & (ax6x)) + ((shiftx0x) & (!shiftx1x) & (ax9x) & (ax8x) & (ax7x) & (!ax6x)) + ((shiftx0x) & (!shiftx1x) & (ax9x) & (ax8x) & (ax7x) & (ax6x)) + ((shiftx0x) & (shiftx1x) & (!ax9x) & (!ax8x) & (!ax7x) & (ax6x)) + ((shiftx0x) & (shiftx1x) & (!ax9x) & (!ax8x) & (ax7x) & (ax6x)) + ((shiftx0x) & (shiftx1x) & (!ax9x) & (ax8x) & (!ax7x) & (ax6x)) + ((shiftx0x) & (shiftx1x) & (!ax9x) & (ax8x) & (ax7x) & (ax6x)) + ((shiftx0x) & (shiftx1x) & (ax9x) & (!ax8x) & (!ax7x) & (ax6x)) + ((shiftx0x) & (shiftx1x) & (ax9x) & (!ax8x) & (ax7x) & (ax6x)) + ((shiftx0x) & (shiftx1x) & (ax9x) & (ax8x) & (!ax7x) & (ax6x)) + ((shiftx0x) & (shiftx1x) & (ax9x) & (ax8x) & (ax7x) & (ax6x)));
	assign g53 = (((!shiftx2x) & (!shiftx3x) & (g49) & (!g50) & (!g51) & (!g52)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (!g50) & (!g51) & (g52)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (!g50) & (g51) & (!g52)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (!g50) & (g51) & (g52)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (g50) & (!g51) & (!g52)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (g50) & (!g51) & (g52)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (g50) & (g51) & (!g52)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (g50) & (g51) & (g52)) + ((!shiftx2x) & (shiftx3x) & (!g49) & (!g50) & (!g51) & (g52)) + ((!shiftx2x) & (shiftx3x) & (!g49) & (!g50) & (g51) & (g52)) + ((!shiftx2x) & (shiftx3x) & (!g49) & (g50) & (!g51) & (g52)) + ((!shiftx2x) & (shiftx3x) & (!g49) & (g50) & (g51) & (g52)) + ((!shiftx2x) & (shiftx3x) & (g49) & (!g50) & (!g51) & (g52)) + ((!shiftx2x) & (shiftx3x) & (g49) & (!g50) & (g51) & (g52)) + ((!shiftx2x) & (shiftx3x) & (g49) & (g50) & (!g51) & (g52)) + ((!shiftx2x) & (shiftx3x) & (g49) & (g50) & (g51) & (g52)) + ((shiftx2x) & (!shiftx3x) & (!g49) & (g50) & (!g51) & (!g52)) + ((shiftx2x) & (!shiftx3x) & (!g49) & (g50) & (!g51) & (g52)) + ((shiftx2x) & (!shiftx3x) & (!g49) & (g50) & (g51) & (!g52)) + ((shiftx2x) & (!shiftx3x) & (!g49) & (g50) & (g51) & (g52)) + ((shiftx2x) & (!shiftx3x) & (g49) & (g50) & (!g51) & (!g52)) + ((shiftx2x) & (!shiftx3x) & (g49) & (g50) & (!g51) & (g52)) + ((shiftx2x) & (!shiftx3x) & (g49) & (g50) & (g51) & (!g52)) + ((shiftx2x) & (!shiftx3x) & (g49) & (g50) & (g51) & (g52)) + ((shiftx2x) & (shiftx3x) & (!g49) & (!g50) & (g51) & (!g52)) + ((shiftx2x) & (shiftx3x) & (!g49) & (!g50) & (g51) & (g52)) + ((shiftx2x) & (shiftx3x) & (!g49) & (g50) & (g51) & (!g52)) + ((shiftx2x) & (shiftx3x) & (!g49) & (g50) & (g51) & (g52)) + ((shiftx2x) & (shiftx3x) & (g49) & (!g50) & (g51) & (!g52)) + ((shiftx2x) & (shiftx3x) & (g49) & (!g50) & (g51) & (g52)) + ((shiftx2x) & (shiftx3x) & (g49) & (g50) & (g51) & (!g52)) + ((shiftx2x) & (shiftx3x) & (g49) & (g50) & (g51) & (g52)));
	assign g54 = (((!shiftx0x) & (!shiftx1x) & (ax49x) & (!ax48x) & (!ax47x) & (!ax46x)) + ((!shiftx0x) & (!shiftx1x) & (ax49x) & (!ax48x) & (!ax47x) & (ax46x)) + ((!shiftx0x) & (!shiftx1x) & (ax49x) & (!ax48x) & (ax47x) & (!ax46x)) + ((!shiftx0x) & (!shiftx1x) & (ax49x) & (!ax48x) & (ax47x) & (ax46x)) + ((!shiftx0x) & (!shiftx1x) & (ax49x) & (ax48x) & (!ax47x) & (!ax46x)) + ((!shiftx0x) & (!shiftx1x) & (ax49x) & (ax48x) & (!ax47x) & (ax46x)) + ((!shiftx0x) & (!shiftx1x) & (ax49x) & (ax48x) & (ax47x) & (!ax46x)) + ((!shiftx0x) & (!shiftx1x) & (ax49x) & (ax48x) & (ax47x) & (ax46x)) + ((!shiftx0x) & (shiftx1x) & (!ax49x) & (!ax48x) & (ax47x) & (!ax46x)) + ((!shiftx0x) & (shiftx1x) & (!ax49x) & (!ax48x) & (ax47x) & (ax46x)) + ((!shiftx0x) & (shiftx1x) & (!ax49x) & (ax48x) & (ax47x) & (!ax46x)) + ((!shiftx0x) & (shiftx1x) & (!ax49x) & (ax48x) & (ax47x) & (ax46x)) + ((!shiftx0x) & (shiftx1x) & (ax49x) & (!ax48x) & (ax47x) & (!ax46x)) + ((!shiftx0x) & (shiftx1x) & (ax49x) & (!ax48x) & (ax47x) & (ax46x)) + ((!shiftx0x) & (shiftx1x) & (ax49x) & (ax48x) & (ax47x) & (!ax46x)) + ((!shiftx0x) & (shiftx1x) & (ax49x) & (ax48x) & (ax47x) & (ax46x)) + ((shiftx0x) & (!shiftx1x) & (!ax49x) & (ax48x) & (!ax47x) & (!ax46x)) + ((shiftx0x) & (!shiftx1x) & (!ax49x) & (ax48x) & (!ax47x) & (ax46x)) + ((shiftx0x) & (!shiftx1x) & (!ax49x) & (ax48x) & (ax47x) & (!ax46x)) + ((shiftx0x) & (!shiftx1x) & (!ax49x) & (ax48x) & (ax47x) & (ax46x)) + ((shiftx0x) & (!shiftx1x) & (ax49x) & (ax48x) & (!ax47x) & (!ax46x)) + ((shiftx0x) & (!shiftx1x) & (ax49x) & (ax48x) & (!ax47x) & (ax46x)) + ((shiftx0x) & (!shiftx1x) & (ax49x) & (ax48x) & (ax47x) & (!ax46x)) + ((shiftx0x) & (!shiftx1x) & (ax49x) & (ax48x) & (ax47x) & (ax46x)) + ((shiftx0x) & (shiftx1x) & (!ax49x) & (!ax48x) & (!ax47x) & (ax46x)) + ((shiftx0x) & (shiftx1x) & (!ax49x) & (!ax48x) & (ax47x) & (ax46x)) + ((shiftx0x) & (shiftx1x) & (!ax49x) & (ax48x) & (!ax47x) & (ax46x)) + ((shiftx0x) & (shiftx1x) & (!ax49x) & (ax48x) & (ax47x) & (ax46x)) + ((shiftx0x) & (shiftx1x) & (ax49x) & (!ax48x) & (!ax47x) & (ax46x)) + ((shiftx0x) & (shiftx1x) & (ax49x) & (!ax48x) & (ax47x) & (ax46x)) + ((shiftx0x) & (shiftx1x) & (ax49x) & (ax48x) & (!ax47x) & (ax46x)) + ((shiftx0x) & (shiftx1x) & (ax49x) & (ax48x) & (ax47x) & (ax46x)));
	assign g55 = (((!ax45x) & (!ax44x) & (!ax43x) & (ax42x) & (shiftx0x) & (shiftx1x)) + ((!ax45x) & (!ax44x) & (ax43x) & (!ax42x) & (!shiftx0x) & (shiftx1x)) + ((!ax45x) & (!ax44x) & (ax43x) & (ax42x) & (!shiftx0x) & (shiftx1x)) + ((!ax45x) & (!ax44x) & (ax43x) & (ax42x) & (shiftx0x) & (shiftx1x)) + ((!ax45x) & (ax44x) & (!ax43x) & (!ax42x) & (shiftx0x) & (!shiftx1x)) + ((!ax45x) & (ax44x) & (!ax43x) & (ax42x) & (shiftx0x) & (!shiftx1x)) + ((!ax45x) & (ax44x) & (!ax43x) & (ax42x) & (shiftx0x) & (shiftx1x)) + ((!ax45x) & (ax44x) & (ax43x) & (!ax42x) & (!shiftx0x) & (shiftx1x)) + ((!ax45x) & (ax44x) & (ax43x) & (!ax42x) & (shiftx0x) & (!shiftx1x)) + ((!ax45x) & (ax44x) & (ax43x) & (ax42x) & (!shiftx0x) & (shiftx1x)) + ((!ax45x) & (ax44x) & (ax43x) & (ax42x) & (shiftx0x) & (!shiftx1x)) + ((!ax45x) & (ax44x) & (ax43x) & (ax42x) & (shiftx0x) & (shiftx1x)) + ((ax45x) & (!ax44x) & (!ax43x) & (!ax42x) & (!shiftx0x) & (!shiftx1x)) + ((ax45x) & (!ax44x) & (!ax43x) & (ax42x) & (!shiftx0x) & (!shiftx1x)) + ((ax45x) & (!ax44x) & (!ax43x) & (ax42x) & (shiftx0x) & (shiftx1x)) + ((ax45x) & (!ax44x) & (ax43x) & (!ax42x) & (!shiftx0x) & (!shiftx1x)) + ((ax45x) & (!ax44x) & (ax43x) & (!ax42x) & (!shiftx0x) & (shiftx1x)) + ((ax45x) & (!ax44x) & (ax43x) & (ax42x) & (!shiftx0x) & (!shiftx1x)) + ((ax45x) & (!ax44x) & (ax43x) & (ax42x) & (!shiftx0x) & (shiftx1x)) + ((ax45x) & (!ax44x) & (ax43x) & (ax42x) & (shiftx0x) & (shiftx1x)) + ((ax45x) & (ax44x) & (!ax43x) & (!ax42x) & (!shiftx0x) & (!shiftx1x)) + ((ax45x) & (ax44x) & (!ax43x) & (!ax42x) & (shiftx0x) & (!shiftx1x)) + ((ax45x) & (ax44x) & (!ax43x) & (ax42x) & (!shiftx0x) & (!shiftx1x)) + ((ax45x) & (ax44x) & (!ax43x) & (ax42x) & (shiftx0x) & (!shiftx1x)) + ((ax45x) & (ax44x) & (!ax43x) & (ax42x) & (shiftx0x) & (shiftx1x)) + ((ax45x) & (ax44x) & (ax43x) & (!ax42x) & (!shiftx0x) & (!shiftx1x)) + ((ax45x) & (ax44x) & (ax43x) & (!ax42x) & (!shiftx0x) & (shiftx1x)) + ((ax45x) & (ax44x) & (ax43x) & (!ax42x) & (shiftx0x) & (!shiftx1x)) + ((ax45x) & (ax44x) & (ax43x) & (ax42x) & (!shiftx0x) & (!shiftx1x)) + ((ax45x) & (ax44x) & (ax43x) & (ax42x) & (!shiftx0x) & (shiftx1x)) + ((ax45x) & (ax44x) & (ax43x) & (ax42x) & (shiftx0x) & (!shiftx1x)) + ((ax45x) & (ax44x) & (ax43x) & (ax42x) & (shiftx0x) & (shiftx1x)));
	assign g56 = (((!shiftx0x) & (!shiftx1x) & (!ax36x) & (!ax35x) & (!ax34x) & (ax37x)) + ((!shiftx0x) & (!shiftx1x) & (!ax36x) & (!ax35x) & (ax34x) & (ax37x)) + ((!shiftx0x) & (!shiftx1x) & (!ax36x) & (ax35x) & (!ax34x) & (ax37x)) + ((!shiftx0x) & (!shiftx1x) & (!ax36x) & (ax35x) & (ax34x) & (ax37x)) + ((!shiftx0x) & (!shiftx1x) & (ax36x) & (!ax35x) & (!ax34x) & (ax37x)) + ((!shiftx0x) & (!shiftx1x) & (ax36x) & (!ax35x) & (ax34x) & (ax37x)) + ((!shiftx0x) & (!shiftx1x) & (ax36x) & (ax35x) & (!ax34x) & (ax37x)) + ((!shiftx0x) & (!shiftx1x) & (ax36x) & (ax35x) & (ax34x) & (ax37x)) + ((!shiftx0x) & (shiftx1x) & (!ax36x) & (ax35x) & (!ax34x) & (!ax37x)) + ((!shiftx0x) & (shiftx1x) & (!ax36x) & (ax35x) & (!ax34x) & (ax37x)) + ((!shiftx0x) & (shiftx1x) & (!ax36x) & (ax35x) & (ax34x) & (!ax37x)) + ((!shiftx0x) & (shiftx1x) & (!ax36x) & (ax35x) & (ax34x) & (ax37x)) + ((!shiftx0x) & (shiftx1x) & (ax36x) & (ax35x) & (!ax34x) & (!ax37x)) + ((!shiftx0x) & (shiftx1x) & (ax36x) & (ax35x) & (!ax34x) & (ax37x)) + ((!shiftx0x) & (shiftx1x) & (ax36x) & (ax35x) & (ax34x) & (!ax37x)) + ((!shiftx0x) & (shiftx1x) & (ax36x) & (ax35x) & (ax34x) & (ax37x)) + ((shiftx0x) & (!shiftx1x) & (ax36x) & (!ax35x) & (!ax34x) & (!ax37x)) + ((shiftx0x) & (!shiftx1x) & (ax36x) & (!ax35x) & (!ax34x) & (ax37x)) + ((shiftx0x) & (!shiftx1x) & (ax36x) & (!ax35x) & (ax34x) & (!ax37x)) + ((shiftx0x) & (!shiftx1x) & (ax36x) & (!ax35x) & (ax34x) & (ax37x)) + ((shiftx0x) & (!shiftx1x) & (ax36x) & (ax35x) & (!ax34x) & (!ax37x)) + ((shiftx0x) & (!shiftx1x) & (ax36x) & (ax35x) & (!ax34x) & (ax37x)) + ((shiftx0x) & (!shiftx1x) & (ax36x) & (ax35x) & (ax34x) & (!ax37x)) + ((shiftx0x) & (!shiftx1x) & (ax36x) & (ax35x) & (ax34x) & (ax37x)) + ((shiftx0x) & (shiftx1x) & (!ax36x) & (!ax35x) & (ax34x) & (!ax37x)) + ((shiftx0x) & (shiftx1x) & (!ax36x) & (!ax35x) & (ax34x) & (ax37x)) + ((shiftx0x) & (shiftx1x) & (!ax36x) & (ax35x) & (ax34x) & (!ax37x)) + ((shiftx0x) & (shiftx1x) & (!ax36x) & (ax35x) & (ax34x) & (ax37x)) + ((shiftx0x) & (shiftx1x) & (ax36x) & (!ax35x) & (ax34x) & (!ax37x)) + ((shiftx0x) & (shiftx1x) & (ax36x) & (!ax35x) & (ax34x) & (ax37x)) + ((shiftx0x) & (shiftx1x) & (ax36x) & (ax35x) & (ax34x) & (!ax37x)) + ((shiftx0x) & (shiftx1x) & (ax36x) & (ax35x) & (ax34x) & (ax37x)));
	assign g57 = (((!ax41x) & (!ax40x) & (!ax39x) & (ax38x) & (shiftx0x) & (shiftx1x)) + ((!ax41x) & (!ax40x) & (ax39x) & (!ax38x) & (!shiftx0x) & (shiftx1x)) + ((!ax41x) & (!ax40x) & (ax39x) & (ax38x) & (!shiftx0x) & (shiftx1x)) + ((!ax41x) & (!ax40x) & (ax39x) & (ax38x) & (shiftx0x) & (shiftx1x)) + ((!ax41x) & (ax40x) & (!ax39x) & (!ax38x) & (shiftx0x) & (!shiftx1x)) + ((!ax41x) & (ax40x) & (!ax39x) & (ax38x) & (shiftx0x) & (!shiftx1x)) + ((!ax41x) & (ax40x) & (!ax39x) & (ax38x) & (shiftx0x) & (shiftx1x)) + ((!ax41x) & (ax40x) & (ax39x) & (!ax38x) & (!shiftx0x) & (shiftx1x)) + ((!ax41x) & (ax40x) & (ax39x) & (!ax38x) & (shiftx0x) & (!shiftx1x)) + ((!ax41x) & (ax40x) & (ax39x) & (ax38x) & (!shiftx0x) & (shiftx1x)) + ((!ax41x) & (ax40x) & (ax39x) & (ax38x) & (shiftx0x) & (!shiftx1x)) + ((!ax41x) & (ax40x) & (ax39x) & (ax38x) & (shiftx0x) & (shiftx1x)) + ((ax41x) & (!ax40x) & (!ax39x) & (!ax38x) & (!shiftx0x) & (!shiftx1x)) + ((ax41x) & (!ax40x) & (!ax39x) & (ax38x) & (!shiftx0x) & (!shiftx1x)) + ((ax41x) & (!ax40x) & (!ax39x) & (ax38x) & (shiftx0x) & (shiftx1x)) + ((ax41x) & (!ax40x) & (ax39x) & (!ax38x) & (!shiftx0x) & (!shiftx1x)) + ((ax41x) & (!ax40x) & (ax39x) & (!ax38x) & (!shiftx0x) & (shiftx1x)) + ((ax41x) & (!ax40x) & (ax39x) & (ax38x) & (!shiftx0x) & (!shiftx1x)) + ((ax41x) & (!ax40x) & (ax39x) & (ax38x) & (!shiftx0x) & (shiftx1x)) + ((ax41x) & (!ax40x) & (ax39x) & (ax38x) & (shiftx0x) & (shiftx1x)) + ((ax41x) & (ax40x) & (!ax39x) & (!ax38x) & (!shiftx0x) & (!shiftx1x)) + ((ax41x) & (ax40x) & (!ax39x) & (!ax38x) & (shiftx0x) & (!shiftx1x)) + ((ax41x) & (ax40x) & (!ax39x) & (ax38x) & (!shiftx0x) & (!shiftx1x)) + ((ax41x) & (ax40x) & (!ax39x) & (ax38x) & (shiftx0x) & (!shiftx1x)) + ((ax41x) & (ax40x) & (!ax39x) & (ax38x) & (shiftx0x) & (shiftx1x)) + ((ax41x) & (ax40x) & (ax39x) & (!ax38x) & (!shiftx0x) & (!shiftx1x)) + ((ax41x) & (ax40x) & (ax39x) & (!ax38x) & (!shiftx0x) & (shiftx1x)) + ((ax41x) & (ax40x) & (ax39x) & (!ax38x) & (shiftx0x) & (!shiftx1x)) + ((ax41x) & (ax40x) & (ax39x) & (ax38x) & (!shiftx0x) & (!shiftx1x)) + ((ax41x) & (ax40x) & (ax39x) & (ax38x) & (!shiftx0x) & (shiftx1x)) + ((ax41x) & (ax40x) & (ax39x) & (ax38x) & (shiftx0x) & (!shiftx1x)) + ((ax41x) & (ax40x) & (ax39x) & (ax38x) & (shiftx0x) & (shiftx1x)));
	assign g58 = (((!shiftx2x) & (!shiftx3x) & (g54) & (!g55) & (!g56) & (!g57)) + ((!shiftx2x) & (!shiftx3x) & (g54) & (!g55) & (!g56) & (g57)) + ((!shiftx2x) & (!shiftx3x) & (g54) & (!g55) & (g56) & (!g57)) + ((!shiftx2x) & (!shiftx3x) & (g54) & (!g55) & (g56) & (g57)) + ((!shiftx2x) & (!shiftx3x) & (g54) & (g55) & (!g56) & (!g57)) + ((!shiftx2x) & (!shiftx3x) & (g54) & (g55) & (!g56) & (g57)) + ((!shiftx2x) & (!shiftx3x) & (g54) & (g55) & (g56) & (!g57)) + ((!shiftx2x) & (!shiftx3x) & (g54) & (g55) & (g56) & (g57)) + ((!shiftx2x) & (shiftx3x) & (!g54) & (!g55) & (!g56) & (g57)) + ((!shiftx2x) & (shiftx3x) & (!g54) & (!g55) & (g56) & (g57)) + ((!shiftx2x) & (shiftx3x) & (!g54) & (g55) & (!g56) & (g57)) + ((!shiftx2x) & (shiftx3x) & (!g54) & (g55) & (g56) & (g57)) + ((!shiftx2x) & (shiftx3x) & (g54) & (!g55) & (!g56) & (g57)) + ((!shiftx2x) & (shiftx3x) & (g54) & (!g55) & (g56) & (g57)) + ((!shiftx2x) & (shiftx3x) & (g54) & (g55) & (!g56) & (g57)) + ((!shiftx2x) & (shiftx3x) & (g54) & (g55) & (g56) & (g57)) + ((shiftx2x) & (!shiftx3x) & (!g54) & (g55) & (!g56) & (!g57)) + ((shiftx2x) & (!shiftx3x) & (!g54) & (g55) & (!g56) & (g57)) + ((shiftx2x) & (!shiftx3x) & (!g54) & (g55) & (g56) & (!g57)) + ((shiftx2x) & (!shiftx3x) & (!g54) & (g55) & (g56) & (g57)) + ((shiftx2x) & (!shiftx3x) & (g54) & (g55) & (!g56) & (!g57)) + ((shiftx2x) & (!shiftx3x) & (g54) & (g55) & (!g56) & (g57)) + ((shiftx2x) & (!shiftx3x) & (g54) & (g55) & (g56) & (!g57)) + ((shiftx2x) & (!shiftx3x) & (g54) & (g55) & (g56) & (g57)) + ((shiftx2x) & (shiftx3x) & (!g54) & (!g55) & (g56) & (!g57)) + ((shiftx2x) & (shiftx3x) & (!g54) & (!g55) & (g56) & (g57)) + ((shiftx2x) & (shiftx3x) & (!g54) & (g55) & (g56) & (!g57)) + ((shiftx2x) & (shiftx3x) & (!g54) & (g55) & (g56) & (g57)) + ((shiftx2x) & (shiftx3x) & (g54) & (!g55) & (g56) & (!g57)) + ((shiftx2x) & (shiftx3x) & (g54) & (!g55) & (g56) & (g57)) + ((shiftx2x) & (shiftx3x) & (g54) & (g55) & (g56) & (!g57)) + ((shiftx2x) & (shiftx3x) & (g54) & (g55) & (g56) & (g57)));
	assign g59 = (((!shiftx0x) & (!shiftx1x) & (!ax32x) & (!ax31x) & (!ax30x) & (ax33x)) + ((!shiftx0x) & (!shiftx1x) & (!ax32x) & (!ax31x) & (ax30x) & (ax33x)) + ((!shiftx0x) & (!shiftx1x) & (!ax32x) & (ax31x) & (!ax30x) & (ax33x)) + ((!shiftx0x) & (!shiftx1x) & (!ax32x) & (ax31x) & (ax30x) & (ax33x)) + ((!shiftx0x) & (!shiftx1x) & (ax32x) & (!ax31x) & (!ax30x) & (ax33x)) + ((!shiftx0x) & (!shiftx1x) & (ax32x) & (!ax31x) & (ax30x) & (ax33x)) + ((!shiftx0x) & (!shiftx1x) & (ax32x) & (ax31x) & (!ax30x) & (ax33x)) + ((!shiftx0x) & (!shiftx1x) & (ax32x) & (ax31x) & (ax30x) & (ax33x)) + ((!shiftx0x) & (shiftx1x) & (!ax32x) & (ax31x) & (!ax30x) & (!ax33x)) + ((!shiftx0x) & (shiftx1x) & (!ax32x) & (ax31x) & (!ax30x) & (ax33x)) + ((!shiftx0x) & (shiftx1x) & (!ax32x) & (ax31x) & (ax30x) & (!ax33x)) + ((!shiftx0x) & (shiftx1x) & (!ax32x) & (ax31x) & (ax30x) & (ax33x)) + ((!shiftx0x) & (shiftx1x) & (ax32x) & (ax31x) & (!ax30x) & (!ax33x)) + ((!shiftx0x) & (shiftx1x) & (ax32x) & (ax31x) & (!ax30x) & (ax33x)) + ((!shiftx0x) & (shiftx1x) & (ax32x) & (ax31x) & (ax30x) & (!ax33x)) + ((!shiftx0x) & (shiftx1x) & (ax32x) & (ax31x) & (ax30x) & (ax33x)) + ((shiftx0x) & (!shiftx1x) & (ax32x) & (!ax31x) & (!ax30x) & (!ax33x)) + ((shiftx0x) & (!shiftx1x) & (ax32x) & (!ax31x) & (!ax30x) & (ax33x)) + ((shiftx0x) & (!shiftx1x) & (ax32x) & (!ax31x) & (ax30x) & (!ax33x)) + ((shiftx0x) & (!shiftx1x) & (ax32x) & (!ax31x) & (ax30x) & (ax33x)) + ((shiftx0x) & (!shiftx1x) & (ax32x) & (ax31x) & (!ax30x) & (!ax33x)) + ((shiftx0x) & (!shiftx1x) & (ax32x) & (ax31x) & (!ax30x) & (ax33x)) + ((shiftx0x) & (!shiftx1x) & (ax32x) & (ax31x) & (ax30x) & (!ax33x)) + ((shiftx0x) & (!shiftx1x) & (ax32x) & (ax31x) & (ax30x) & (ax33x)) + ((shiftx0x) & (shiftx1x) & (!ax32x) & (!ax31x) & (ax30x) & (!ax33x)) + ((shiftx0x) & (shiftx1x) & (!ax32x) & (!ax31x) & (ax30x) & (ax33x)) + ((shiftx0x) & (shiftx1x) & (!ax32x) & (ax31x) & (ax30x) & (!ax33x)) + ((shiftx0x) & (shiftx1x) & (!ax32x) & (ax31x) & (ax30x) & (ax33x)) + ((shiftx0x) & (shiftx1x) & (ax32x) & (!ax31x) & (ax30x) & (!ax33x)) + ((shiftx0x) & (shiftx1x) & (ax32x) & (!ax31x) & (ax30x) & (ax33x)) + ((shiftx0x) & (shiftx1x) & (ax32x) & (ax31x) & (ax30x) & (!ax33x)) + ((shiftx0x) & (shiftx1x) & (ax32x) & (ax31x) & (ax30x) & (ax33x)));
	assign g60 = (((!shiftx0x) & (!shiftx1x) & (ax29x) & (!ax28x) & (!ax27x) & (!ax26x)) + ((!shiftx0x) & (!shiftx1x) & (ax29x) & (!ax28x) & (!ax27x) & (ax26x)) + ((!shiftx0x) & (!shiftx1x) & (ax29x) & (!ax28x) & (ax27x) & (!ax26x)) + ((!shiftx0x) & (!shiftx1x) & (ax29x) & (!ax28x) & (ax27x) & (ax26x)) + ((!shiftx0x) & (!shiftx1x) & (ax29x) & (ax28x) & (!ax27x) & (!ax26x)) + ((!shiftx0x) & (!shiftx1x) & (ax29x) & (ax28x) & (!ax27x) & (ax26x)) + ((!shiftx0x) & (!shiftx1x) & (ax29x) & (ax28x) & (ax27x) & (!ax26x)) + ((!shiftx0x) & (!shiftx1x) & (ax29x) & (ax28x) & (ax27x) & (ax26x)) + ((!shiftx0x) & (shiftx1x) & (!ax29x) & (!ax28x) & (ax27x) & (!ax26x)) + ((!shiftx0x) & (shiftx1x) & (!ax29x) & (!ax28x) & (ax27x) & (ax26x)) + ((!shiftx0x) & (shiftx1x) & (!ax29x) & (ax28x) & (ax27x) & (!ax26x)) + ((!shiftx0x) & (shiftx1x) & (!ax29x) & (ax28x) & (ax27x) & (ax26x)) + ((!shiftx0x) & (shiftx1x) & (ax29x) & (!ax28x) & (ax27x) & (!ax26x)) + ((!shiftx0x) & (shiftx1x) & (ax29x) & (!ax28x) & (ax27x) & (ax26x)) + ((!shiftx0x) & (shiftx1x) & (ax29x) & (ax28x) & (ax27x) & (!ax26x)) + ((!shiftx0x) & (shiftx1x) & (ax29x) & (ax28x) & (ax27x) & (ax26x)) + ((shiftx0x) & (!shiftx1x) & (!ax29x) & (ax28x) & (!ax27x) & (!ax26x)) + ((shiftx0x) & (!shiftx1x) & (!ax29x) & (ax28x) & (!ax27x) & (ax26x)) + ((shiftx0x) & (!shiftx1x) & (!ax29x) & (ax28x) & (ax27x) & (!ax26x)) + ((shiftx0x) & (!shiftx1x) & (!ax29x) & (ax28x) & (ax27x) & (ax26x)) + ((shiftx0x) & (!shiftx1x) & (ax29x) & (ax28x) & (!ax27x) & (!ax26x)) + ((shiftx0x) & (!shiftx1x) & (ax29x) & (ax28x) & (!ax27x) & (ax26x)) + ((shiftx0x) & (!shiftx1x) & (ax29x) & (ax28x) & (ax27x) & (!ax26x)) + ((shiftx0x) & (!shiftx1x) & (ax29x) & (ax28x) & (ax27x) & (ax26x)) + ((shiftx0x) & (shiftx1x) & (!ax29x) & (!ax28x) & (!ax27x) & (ax26x)) + ((shiftx0x) & (shiftx1x) & (!ax29x) & (!ax28x) & (ax27x) & (ax26x)) + ((shiftx0x) & (shiftx1x) & (!ax29x) & (ax28x) & (!ax27x) & (ax26x)) + ((shiftx0x) & (shiftx1x) & (!ax29x) & (ax28x) & (ax27x) & (ax26x)) + ((shiftx0x) & (shiftx1x) & (ax29x) & (!ax28x) & (!ax27x) & (ax26x)) + ((shiftx0x) & (shiftx1x) & (ax29x) & (!ax28x) & (ax27x) & (ax26x)) + ((shiftx0x) & (shiftx1x) & (ax29x) & (ax28x) & (!ax27x) & (ax26x)) + ((shiftx0x) & (shiftx1x) & (ax29x) & (ax28x) & (ax27x) & (ax26x)));
	assign g61 = (((!shiftx0x) & (!shiftx1x) & (!ax20x) & (!ax19x) & (!ax18x) & (ax21x)) + ((!shiftx0x) & (!shiftx1x) & (!ax20x) & (!ax19x) & (ax18x) & (ax21x)) + ((!shiftx0x) & (!shiftx1x) & (!ax20x) & (ax19x) & (!ax18x) & (ax21x)) + ((!shiftx0x) & (!shiftx1x) & (!ax20x) & (ax19x) & (ax18x) & (ax21x)) + ((!shiftx0x) & (!shiftx1x) & (ax20x) & (!ax19x) & (!ax18x) & (ax21x)) + ((!shiftx0x) & (!shiftx1x) & (ax20x) & (!ax19x) & (ax18x) & (ax21x)) + ((!shiftx0x) & (!shiftx1x) & (ax20x) & (ax19x) & (!ax18x) & (ax21x)) + ((!shiftx0x) & (!shiftx1x) & (ax20x) & (ax19x) & (ax18x) & (ax21x)) + ((!shiftx0x) & (shiftx1x) & (!ax20x) & (ax19x) & (!ax18x) & (!ax21x)) + ((!shiftx0x) & (shiftx1x) & (!ax20x) & (ax19x) & (!ax18x) & (ax21x)) + ((!shiftx0x) & (shiftx1x) & (!ax20x) & (ax19x) & (ax18x) & (!ax21x)) + ((!shiftx0x) & (shiftx1x) & (!ax20x) & (ax19x) & (ax18x) & (ax21x)) + ((!shiftx0x) & (shiftx1x) & (ax20x) & (ax19x) & (!ax18x) & (!ax21x)) + ((!shiftx0x) & (shiftx1x) & (ax20x) & (ax19x) & (!ax18x) & (ax21x)) + ((!shiftx0x) & (shiftx1x) & (ax20x) & (ax19x) & (ax18x) & (!ax21x)) + ((!shiftx0x) & (shiftx1x) & (ax20x) & (ax19x) & (ax18x) & (ax21x)) + ((shiftx0x) & (!shiftx1x) & (ax20x) & (!ax19x) & (!ax18x) & (!ax21x)) + ((shiftx0x) & (!shiftx1x) & (ax20x) & (!ax19x) & (!ax18x) & (ax21x)) + ((shiftx0x) & (!shiftx1x) & (ax20x) & (!ax19x) & (ax18x) & (!ax21x)) + ((shiftx0x) & (!shiftx1x) & (ax20x) & (!ax19x) & (ax18x) & (ax21x)) + ((shiftx0x) & (!shiftx1x) & (ax20x) & (ax19x) & (!ax18x) & (!ax21x)) + ((shiftx0x) & (!shiftx1x) & (ax20x) & (ax19x) & (!ax18x) & (ax21x)) + ((shiftx0x) & (!shiftx1x) & (ax20x) & (ax19x) & (ax18x) & (!ax21x)) + ((shiftx0x) & (!shiftx1x) & (ax20x) & (ax19x) & (ax18x) & (ax21x)) + ((shiftx0x) & (shiftx1x) & (!ax20x) & (!ax19x) & (ax18x) & (!ax21x)) + ((shiftx0x) & (shiftx1x) & (!ax20x) & (!ax19x) & (ax18x) & (ax21x)) + ((shiftx0x) & (shiftx1x) & (!ax20x) & (ax19x) & (ax18x) & (!ax21x)) + ((shiftx0x) & (shiftx1x) & (!ax20x) & (ax19x) & (ax18x) & (ax21x)) + ((shiftx0x) & (shiftx1x) & (ax20x) & (!ax19x) & (ax18x) & (!ax21x)) + ((shiftx0x) & (shiftx1x) & (ax20x) & (!ax19x) & (ax18x) & (ax21x)) + ((shiftx0x) & (shiftx1x) & (ax20x) & (ax19x) & (ax18x) & (!ax21x)) + ((shiftx0x) & (shiftx1x) & (ax20x) & (ax19x) & (ax18x) & (ax21x)));
	assign g62 = (((!shiftx0x) & (!shiftx1x) & (ax25x) & (!ax24x) & (!ax23x) & (!ax22x)) + ((!shiftx0x) & (!shiftx1x) & (ax25x) & (!ax24x) & (!ax23x) & (ax22x)) + ((!shiftx0x) & (!shiftx1x) & (ax25x) & (!ax24x) & (ax23x) & (!ax22x)) + ((!shiftx0x) & (!shiftx1x) & (ax25x) & (!ax24x) & (ax23x) & (ax22x)) + ((!shiftx0x) & (!shiftx1x) & (ax25x) & (ax24x) & (!ax23x) & (!ax22x)) + ((!shiftx0x) & (!shiftx1x) & (ax25x) & (ax24x) & (!ax23x) & (ax22x)) + ((!shiftx0x) & (!shiftx1x) & (ax25x) & (ax24x) & (ax23x) & (!ax22x)) + ((!shiftx0x) & (!shiftx1x) & (ax25x) & (ax24x) & (ax23x) & (ax22x)) + ((!shiftx0x) & (shiftx1x) & (!ax25x) & (!ax24x) & (ax23x) & (!ax22x)) + ((!shiftx0x) & (shiftx1x) & (!ax25x) & (!ax24x) & (ax23x) & (ax22x)) + ((!shiftx0x) & (shiftx1x) & (!ax25x) & (ax24x) & (ax23x) & (!ax22x)) + ((!shiftx0x) & (shiftx1x) & (!ax25x) & (ax24x) & (ax23x) & (ax22x)) + ((!shiftx0x) & (shiftx1x) & (ax25x) & (!ax24x) & (ax23x) & (!ax22x)) + ((!shiftx0x) & (shiftx1x) & (ax25x) & (!ax24x) & (ax23x) & (ax22x)) + ((!shiftx0x) & (shiftx1x) & (ax25x) & (ax24x) & (ax23x) & (!ax22x)) + ((!shiftx0x) & (shiftx1x) & (ax25x) & (ax24x) & (ax23x) & (ax22x)) + ((shiftx0x) & (!shiftx1x) & (!ax25x) & (ax24x) & (!ax23x) & (!ax22x)) + ((shiftx0x) & (!shiftx1x) & (!ax25x) & (ax24x) & (!ax23x) & (ax22x)) + ((shiftx0x) & (!shiftx1x) & (!ax25x) & (ax24x) & (ax23x) & (!ax22x)) + ((shiftx0x) & (!shiftx1x) & (!ax25x) & (ax24x) & (ax23x) & (ax22x)) + ((shiftx0x) & (!shiftx1x) & (ax25x) & (ax24x) & (!ax23x) & (!ax22x)) + ((shiftx0x) & (!shiftx1x) & (ax25x) & (ax24x) & (!ax23x) & (ax22x)) + ((shiftx0x) & (!shiftx1x) & (ax25x) & (ax24x) & (ax23x) & (!ax22x)) + ((shiftx0x) & (!shiftx1x) & (ax25x) & (ax24x) & (ax23x) & (ax22x)) + ((shiftx0x) & (shiftx1x) & (!ax25x) & (!ax24x) & (!ax23x) & (ax22x)) + ((shiftx0x) & (shiftx1x) & (!ax25x) & (!ax24x) & (ax23x) & (ax22x)) + ((shiftx0x) & (shiftx1x) & (!ax25x) & (ax24x) & (!ax23x) & (ax22x)) + ((shiftx0x) & (shiftx1x) & (!ax25x) & (ax24x) & (ax23x) & (ax22x)) + ((shiftx0x) & (shiftx1x) & (ax25x) & (!ax24x) & (!ax23x) & (ax22x)) + ((shiftx0x) & (shiftx1x) & (ax25x) & (!ax24x) & (ax23x) & (ax22x)) + ((shiftx0x) & (shiftx1x) & (ax25x) & (ax24x) & (!ax23x) & (ax22x)) + ((shiftx0x) & (shiftx1x) & (ax25x) & (ax24x) & (ax23x) & (ax22x)));
	assign g63 = (((!shiftx2x) & (!shiftx3x) & (g59) & (!g60) & (!g61) & (!g62)) + ((!shiftx2x) & (!shiftx3x) & (g59) & (!g60) & (!g61) & (g62)) + ((!shiftx2x) & (!shiftx3x) & (g59) & (!g60) & (g61) & (!g62)) + ((!shiftx2x) & (!shiftx3x) & (g59) & (!g60) & (g61) & (g62)) + ((!shiftx2x) & (!shiftx3x) & (g59) & (g60) & (!g61) & (!g62)) + ((!shiftx2x) & (!shiftx3x) & (g59) & (g60) & (!g61) & (g62)) + ((!shiftx2x) & (!shiftx3x) & (g59) & (g60) & (g61) & (!g62)) + ((!shiftx2x) & (!shiftx3x) & (g59) & (g60) & (g61) & (g62)) + ((!shiftx2x) & (shiftx3x) & (!g59) & (!g60) & (!g61) & (g62)) + ((!shiftx2x) & (shiftx3x) & (!g59) & (!g60) & (g61) & (g62)) + ((!shiftx2x) & (shiftx3x) & (!g59) & (g60) & (!g61) & (g62)) + ((!shiftx2x) & (shiftx3x) & (!g59) & (g60) & (g61) & (g62)) + ((!shiftx2x) & (shiftx3x) & (g59) & (!g60) & (!g61) & (g62)) + ((!shiftx2x) & (shiftx3x) & (g59) & (!g60) & (g61) & (g62)) + ((!shiftx2x) & (shiftx3x) & (g59) & (g60) & (!g61) & (g62)) + ((!shiftx2x) & (shiftx3x) & (g59) & (g60) & (g61) & (g62)) + ((shiftx2x) & (!shiftx3x) & (!g59) & (g60) & (!g61) & (!g62)) + ((shiftx2x) & (!shiftx3x) & (!g59) & (g60) & (!g61) & (g62)) + ((shiftx2x) & (!shiftx3x) & (!g59) & (g60) & (g61) & (!g62)) + ((shiftx2x) & (!shiftx3x) & (!g59) & (g60) & (g61) & (g62)) + ((shiftx2x) & (!shiftx3x) & (g59) & (g60) & (!g61) & (!g62)) + ((shiftx2x) & (!shiftx3x) & (g59) & (g60) & (!g61) & (g62)) + ((shiftx2x) & (!shiftx3x) & (g59) & (g60) & (g61) & (!g62)) + ((shiftx2x) & (!shiftx3x) & (g59) & (g60) & (g61) & (g62)) + ((shiftx2x) & (shiftx3x) & (!g59) & (!g60) & (g61) & (!g62)) + ((shiftx2x) & (shiftx3x) & (!g59) & (!g60) & (g61) & (g62)) + ((shiftx2x) & (shiftx3x) & (!g59) & (g60) & (g61) & (!g62)) + ((shiftx2x) & (shiftx3x) & (!g59) & (g60) & (g61) & (g62)) + ((shiftx2x) & (shiftx3x) & (g59) & (!g60) & (g61) & (!g62)) + ((shiftx2x) & (shiftx3x) & (g59) & (!g60) & (g61) & (g62)) + ((shiftx2x) & (shiftx3x) & (g59) & (g60) & (g61) & (!g62)) + ((shiftx2x) & (shiftx3x) & (g59) & (g60) & (g61) & (g62)));
	assign g64 = (((!shiftx4x) & (!shiftx5x) & (g48) & (!g53) & (!g58) & (!g63)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (!g53) & (!g58) & (g63)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (!g53) & (g58) & (!g63)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (!g53) & (g58) & (g63)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (g53) & (!g58) & (!g63)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (g53) & (!g58) & (g63)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (g53) & (g58) & (!g63)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (g53) & (g58) & (g63)) + ((!shiftx4x) & (shiftx5x) & (!g48) & (!g53) & (!g58) & (g63)) + ((!shiftx4x) & (shiftx5x) & (!g48) & (!g53) & (g58) & (g63)) + ((!shiftx4x) & (shiftx5x) & (!g48) & (g53) & (!g58) & (g63)) + ((!shiftx4x) & (shiftx5x) & (!g48) & (g53) & (g58) & (g63)) + ((!shiftx4x) & (shiftx5x) & (g48) & (!g53) & (!g58) & (g63)) + ((!shiftx4x) & (shiftx5x) & (g48) & (!g53) & (g58) & (g63)) + ((!shiftx4x) & (shiftx5x) & (g48) & (g53) & (!g58) & (g63)) + ((!shiftx4x) & (shiftx5x) & (g48) & (g53) & (g58) & (g63)) + ((shiftx4x) & (!shiftx5x) & (!g48) & (!g53) & (g58) & (!g63)) + ((shiftx4x) & (!shiftx5x) & (!g48) & (!g53) & (g58) & (g63)) + ((shiftx4x) & (!shiftx5x) & (!g48) & (g53) & (g58) & (!g63)) + ((shiftx4x) & (!shiftx5x) & (!g48) & (g53) & (g58) & (g63)) + ((shiftx4x) & (!shiftx5x) & (g48) & (!g53) & (g58) & (!g63)) + ((shiftx4x) & (!shiftx5x) & (g48) & (!g53) & (g58) & (g63)) + ((shiftx4x) & (!shiftx5x) & (g48) & (g53) & (g58) & (!g63)) + ((shiftx4x) & (!shiftx5x) & (g48) & (g53) & (g58) & (g63)) + ((shiftx4x) & (shiftx5x) & (!g48) & (g53) & (!g58) & (!g63)) + ((shiftx4x) & (shiftx5x) & (!g48) & (g53) & (!g58) & (g63)) + ((shiftx4x) & (shiftx5x) & (!g48) & (g53) & (g58) & (!g63)) + ((shiftx4x) & (shiftx5x) & (!g48) & (g53) & (g58) & (g63)) + ((shiftx4x) & (shiftx5x) & (g48) & (g53) & (!g58) & (!g63)) + ((shiftx4x) & (shiftx5x) & (g48) & (g53) & (!g58) & (g63)) + ((shiftx4x) & (shiftx5x) & (g48) & (g53) & (g58) & (!g63)) + ((shiftx4x) & (shiftx5x) & (g48) & (g53) & (g58) & (g63)));
	assign g65 = (((!shiftx0x) & (!shiftx1x) & (!ax80x) & (!ax79x) & (!ax78x) & (ax81x)) + ((!shiftx0x) & (!shiftx1x) & (!ax80x) & (!ax79x) & (ax78x) & (ax81x)) + ((!shiftx0x) & (!shiftx1x) & (!ax80x) & (ax79x) & (!ax78x) & (ax81x)) + ((!shiftx0x) & (!shiftx1x) & (!ax80x) & (ax79x) & (ax78x) & (ax81x)) + ((!shiftx0x) & (!shiftx1x) & (ax80x) & (!ax79x) & (!ax78x) & (ax81x)) + ((!shiftx0x) & (!shiftx1x) & (ax80x) & (!ax79x) & (ax78x) & (ax81x)) + ((!shiftx0x) & (!shiftx1x) & (ax80x) & (ax79x) & (!ax78x) & (ax81x)) + ((!shiftx0x) & (!shiftx1x) & (ax80x) & (ax79x) & (ax78x) & (ax81x)) + ((!shiftx0x) & (shiftx1x) & (!ax80x) & (ax79x) & (!ax78x) & (!ax81x)) + ((!shiftx0x) & (shiftx1x) & (!ax80x) & (ax79x) & (!ax78x) & (ax81x)) + ((!shiftx0x) & (shiftx1x) & (!ax80x) & (ax79x) & (ax78x) & (!ax81x)) + ((!shiftx0x) & (shiftx1x) & (!ax80x) & (ax79x) & (ax78x) & (ax81x)) + ((!shiftx0x) & (shiftx1x) & (ax80x) & (ax79x) & (!ax78x) & (!ax81x)) + ((!shiftx0x) & (shiftx1x) & (ax80x) & (ax79x) & (!ax78x) & (ax81x)) + ((!shiftx0x) & (shiftx1x) & (ax80x) & (ax79x) & (ax78x) & (!ax81x)) + ((!shiftx0x) & (shiftx1x) & (ax80x) & (ax79x) & (ax78x) & (ax81x)) + ((shiftx0x) & (!shiftx1x) & (ax80x) & (!ax79x) & (!ax78x) & (!ax81x)) + ((shiftx0x) & (!shiftx1x) & (ax80x) & (!ax79x) & (!ax78x) & (ax81x)) + ((shiftx0x) & (!shiftx1x) & (ax80x) & (!ax79x) & (ax78x) & (!ax81x)) + ((shiftx0x) & (!shiftx1x) & (ax80x) & (!ax79x) & (ax78x) & (ax81x)) + ((shiftx0x) & (!shiftx1x) & (ax80x) & (ax79x) & (!ax78x) & (!ax81x)) + ((shiftx0x) & (!shiftx1x) & (ax80x) & (ax79x) & (!ax78x) & (ax81x)) + ((shiftx0x) & (!shiftx1x) & (ax80x) & (ax79x) & (ax78x) & (!ax81x)) + ((shiftx0x) & (!shiftx1x) & (ax80x) & (ax79x) & (ax78x) & (ax81x)) + ((shiftx0x) & (shiftx1x) & (!ax80x) & (!ax79x) & (ax78x) & (!ax81x)) + ((shiftx0x) & (shiftx1x) & (!ax80x) & (!ax79x) & (ax78x) & (ax81x)) + ((shiftx0x) & (shiftx1x) & (!ax80x) & (ax79x) & (ax78x) & (!ax81x)) + ((shiftx0x) & (shiftx1x) & (!ax80x) & (ax79x) & (ax78x) & (ax81x)) + ((shiftx0x) & (shiftx1x) & (ax80x) & (!ax79x) & (ax78x) & (!ax81x)) + ((shiftx0x) & (shiftx1x) & (ax80x) & (!ax79x) & (ax78x) & (ax81x)) + ((shiftx0x) & (shiftx1x) & (ax80x) & (ax79x) & (ax78x) & (!ax81x)) + ((shiftx0x) & (shiftx1x) & (ax80x) & (ax79x) & (ax78x) & (ax81x)));
	assign g66 = (((!shiftx0x) & (!shiftx1x) & (ax77x) & (!ax76x) & (!ax75x) & (!ax74x)) + ((!shiftx0x) & (!shiftx1x) & (ax77x) & (!ax76x) & (!ax75x) & (ax74x)) + ((!shiftx0x) & (!shiftx1x) & (ax77x) & (!ax76x) & (ax75x) & (!ax74x)) + ((!shiftx0x) & (!shiftx1x) & (ax77x) & (!ax76x) & (ax75x) & (ax74x)) + ((!shiftx0x) & (!shiftx1x) & (ax77x) & (ax76x) & (!ax75x) & (!ax74x)) + ((!shiftx0x) & (!shiftx1x) & (ax77x) & (ax76x) & (!ax75x) & (ax74x)) + ((!shiftx0x) & (!shiftx1x) & (ax77x) & (ax76x) & (ax75x) & (!ax74x)) + ((!shiftx0x) & (!shiftx1x) & (ax77x) & (ax76x) & (ax75x) & (ax74x)) + ((!shiftx0x) & (shiftx1x) & (!ax77x) & (!ax76x) & (ax75x) & (!ax74x)) + ((!shiftx0x) & (shiftx1x) & (!ax77x) & (!ax76x) & (ax75x) & (ax74x)) + ((!shiftx0x) & (shiftx1x) & (!ax77x) & (ax76x) & (ax75x) & (!ax74x)) + ((!shiftx0x) & (shiftx1x) & (!ax77x) & (ax76x) & (ax75x) & (ax74x)) + ((!shiftx0x) & (shiftx1x) & (ax77x) & (!ax76x) & (ax75x) & (!ax74x)) + ((!shiftx0x) & (shiftx1x) & (ax77x) & (!ax76x) & (ax75x) & (ax74x)) + ((!shiftx0x) & (shiftx1x) & (ax77x) & (ax76x) & (ax75x) & (!ax74x)) + ((!shiftx0x) & (shiftx1x) & (ax77x) & (ax76x) & (ax75x) & (ax74x)) + ((shiftx0x) & (!shiftx1x) & (!ax77x) & (ax76x) & (!ax75x) & (!ax74x)) + ((shiftx0x) & (!shiftx1x) & (!ax77x) & (ax76x) & (!ax75x) & (ax74x)) + ((shiftx0x) & (!shiftx1x) & (!ax77x) & (ax76x) & (ax75x) & (!ax74x)) + ((shiftx0x) & (!shiftx1x) & (!ax77x) & (ax76x) & (ax75x) & (ax74x)) + ((shiftx0x) & (!shiftx1x) & (ax77x) & (ax76x) & (!ax75x) & (!ax74x)) + ((shiftx0x) & (!shiftx1x) & (ax77x) & (ax76x) & (!ax75x) & (ax74x)) + ((shiftx0x) & (!shiftx1x) & (ax77x) & (ax76x) & (ax75x) & (!ax74x)) + ((shiftx0x) & (!shiftx1x) & (ax77x) & (ax76x) & (ax75x) & (ax74x)) + ((shiftx0x) & (shiftx1x) & (!ax77x) & (!ax76x) & (!ax75x) & (ax74x)) + ((shiftx0x) & (shiftx1x) & (!ax77x) & (!ax76x) & (ax75x) & (ax74x)) + ((shiftx0x) & (shiftx1x) & (!ax77x) & (ax76x) & (!ax75x) & (ax74x)) + ((shiftx0x) & (shiftx1x) & (!ax77x) & (ax76x) & (ax75x) & (ax74x)) + ((shiftx0x) & (shiftx1x) & (ax77x) & (!ax76x) & (!ax75x) & (ax74x)) + ((shiftx0x) & (shiftx1x) & (ax77x) & (!ax76x) & (ax75x) & (ax74x)) + ((shiftx0x) & (shiftx1x) & (ax77x) & (ax76x) & (!ax75x) & (ax74x)) + ((shiftx0x) & (shiftx1x) & (ax77x) & (ax76x) & (ax75x) & (ax74x)));
	assign g67 = (((!shiftx0x) & (!shiftx1x) & (!ax68x) & (!ax67x) & (!ax66x) & (ax69x)) + ((!shiftx0x) & (!shiftx1x) & (!ax68x) & (!ax67x) & (ax66x) & (ax69x)) + ((!shiftx0x) & (!shiftx1x) & (!ax68x) & (ax67x) & (!ax66x) & (ax69x)) + ((!shiftx0x) & (!shiftx1x) & (!ax68x) & (ax67x) & (ax66x) & (ax69x)) + ((!shiftx0x) & (!shiftx1x) & (ax68x) & (!ax67x) & (!ax66x) & (ax69x)) + ((!shiftx0x) & (!shiftx1x) & (ax68x) & (!ax67x) & (ax66x) & (ax69x)) + ((!shiftx0x) & (!shiftx1x) & (ax68x) & (ax67x) & (!ax66x) & (ax69x)) + ((!shiftx0x) & (!shiftx1x) & (ax68x) & (ax67x) & (ax66x) & (ax69x)) + ((!shiftx0x) & (shiftx1x) & (!ax68x) & (ax67x) & (!ax66x) & (!ax69x)) + ((!shiftx0x) & (shiftx1x) & (!ax68x) & (ax67x) & (!ax66x) & (ax69x)) + ((!shiftx0x) & (shiftx1x) & (!ax68x) & (ax67x) & (ax66x) & (!ax69x)) + ((!shiftx0x) & (shiftx1x) & (!ax68x) & (ax67x) & (ax66x) & (ax69x)) + ((!shiftx0x) & (shiftx1x) & (ax68x) & (ax67x) & (!ax66x) & (!ax69x)) + ((!shiftx0x) & (shiftx1x) & (ax68x) & (ax67x) & (!ax66x) & (ax69x)) + ((!shiftx0x) & (shiftx1x) & (ax68x) & (ax67x) & (ax66x) & (!ax69x)) + ((!shiftx0x) & (shiftx1x) & (ax68x) & (ax67x) & (ax66x) & (ax69x)) + ((shiftx0x) & (!shiftx1x) & (ax68x) & (!ax67x) & (!ax66x) & (!ax69x)) + ((shiftx0x) & (!shiftx1x) & (ax68x) & (!ax67x) & (!ax66x) & (ax69x)) + ((shiftx0x) & (!shiftx1x) & (ax68x) & (!ax67x) & (ax66x) & (!ax69x)) + ((shiftx0x) & (!shiftx1x) & (ax68x) & (!ax67x) & (ax66x) & (ax69x)) + ((shiftx0x) & (!shiftx1x) & (ax68x) & (ax67x) & (!ax66x) & (!ax69x)) + ((shiftx0x) & (!shiftx1x) & (ax68x) & (ax67x) & (!ax66x) & (ax69x)) + ((shiftx0x) & (!shiftx1x) & (ax68x) & (ax67x) & (ax66x) & (!ax69x)) + ((shiftx0x) & (!shiftx1x) & (ax68x) & (ax67x) & (ax66x) & (ax69x)) + ((shiftx0x) & (shiftx1x) & (!ax68x) & (!ax67x) & (ax66x) & (!ax69x)) + ((shiftx0x) & (shiftx1x) & (!ax68x) & (!ax67x) & (ax66x) & (ax69x)) + ((shiftx0x) & (shiftx1x) & (!ax68x) & (ax67x) & (ax66x) & (!ax69x)) + ((shiftx0x) & (shiftx1x) & (!ax68x) & (ax67x) & (ax66x) & (ax69x)) + ((shiftx0x) & (shiftx1x) & (ax68x) & (!ax67x) & (ax66x) & (!ax69x)) + ((shiftx0x) & (shiftx1x) & (ax68x) & (!ax67x) & (ax66x) & (ax69x)) + ((shiftx0x) & (shiftx1x) & (ax68x) & (ax67x) & (ax66x) & (!ax69x)) + ((shiftx0x) & (shiftx1x) & (ax68x) & (ax67x) & (ax66x) & (ax69x)));
	assign g68 = (((!shiftx0x) & (!shiftx1x) & (ax73x) & (!ax72x) & (!ax71x) & (!ax70x)) + ((!shiftx0x) & (!shiftx1x) & (ax73x) & (!ax72x) & (!ax71x) & (ax70x)) + ((!shiftx0x) & (!shiftx1x) & (ax73x) & (!ax72x) & (ax71x) & (!ax70x)) + ((!shiftx0x) & (!shiftx1x) & (ax73x) & (!ax72x) & (ax71x) & (ax70x)) + ((!shiftx0x) & (!shiftx1x) & (ax73x) & (ax72x) & (!ax71x) & (!ax70x)) + ((!shiftx0x) & (!shiftx1x) & (ax73x) & (ax72x) & (!ax71x) & (ax70x)) + ((!shiftx0x) & (!shiftx1x) & (ax73x) & (ax72x) & (ax71x) & (!ax70x)) + ((!shiftx0x) & (!shiftx1x) & (ax73x) & (ax72x) & (ax71x) & (ax70x)) + ((!shiftx0x) & (shiftx1x) & (!ax73x) & (!ax72x) & (ax71x) & (!ax70x)) + ((!shiftx0x) & (shiftx1x) & (!ax73x) & (!ax72x) & (ax71x) & (ax70x)) + ((!shiftx0x) & (shiftx1x) & (!ax73x) & (ax72x) & (ax71x) & (!ax70x)) + ((!shiftx0x) & (shiftx1x) & (!ax73x) & (ax72x) & (ax71x) & (ax70x)) + ((!shiftx0x) & (shiftx1x) & (ax73x) & (!ax72x) & (ax71x) & (!ax70x)) + ((!shiftx0x) & (shiftx1x) & (ax73x) & (!ax72x) & (ax71x) & (ax70x)) + ((!shiftx0x) & (shiftx1x) & (ax73x) & (ax72x) & (ax71x) & (!ax70x)) + ((!shiftx0x) & (shiftx1x) & (ax73x) & (ax72x) & (ax71x) & (ax70x)) + ((shiftx0x) & (!shiftx1x) & (!ax73x) & (ax72x) & (!ax71x) & (!ax70x)) + ((shiftx0x) & (!shiftx1x) & (!ax73x) & (ax72x) & (!ax71x) & (ax70x)) + ((shiftx0x) & (!shiftx1x) & (!ax73x) & (ax72x) & (ax71x) & (!ax70x)) + ((shiftx0x) & (!shiftx1x) & (!ax73x) & (ax72x) & (ax71x) & (ax70x)) + ((shiftx0x) & (!shiftx1x) & (ax73x) & (ax72x) & (!ax71x) & (!ax70x)) + ((shiftx0x) & (!shiftx1x) & (ax73x) & (ax72x) & (!ax71x) & (ax70x)) + ((shiftx0x) & (!shiftx1x) & (ax73x) & (ax72x) & (ax71x) & (!ax70x)) + ((shiftx0x) & (!shiftx1x) & (ax73x) & (ax72x) & (ax71x) & (ax70x)) + ((shiftx0x) & (shiftx1x) & (!ax73x) & (!ax72x) & (!ax71x) & (ax70x)) + ((shiftx0x) & (shiftx1x) & (!ax73x) & (!ax72x) & (ax71x) & (ax70x)) + ((shiftx0x) & (shiftx1x) & (!ax73x) & (ax72x) & (!ax71x) & (ax70x)) + ((shiftx0x) & (shiftx1x) & (!ax73x) & (ax72x) & (ax71x) & (ax70x)) + ((shiftx0x) & (shiftx1x) & (ax73x) & (!ax72x) & (!ax71x) & (ax70x)) + ((shiftx0x) & (shiftx1x) & (ax73x) & (!ax72x) & (ax71x) & (ax70x)) + ((shiftx0x) & (shiftx1x) & (ax73x) & (ax72x) & (!ax71x) & (ax70x)) + ((shiftx0x) & (shiftx1x) & (ax73x) & (ax72x) & (ax71x) & (ax70x)));
	assign g69 = (((!shiftx2x) & (!shiftx3x) & (g65) & (!g66) & (!g67) & (!g68)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (!g66) & (!g67) & (g68)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (!g66) & (g67) & (!g68)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (!g66) & (g67) & (g68)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (g66) & (!g67) & (!g68)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (g66) & (!g67) & (g68)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (g66) & (g67) & (!g68)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (g66) & (g67) & (g68)) + ((!shiftx2x) & (shiftx3x) & (!g65) & (!g66) & (!g67) & (g68)) + ((!shiftx2x) & (shiftx3x) & (!g65) & (!g66) & (g67) & (g68)) + ((!shiftx2x) & (shiftx3x) & (!g65) & (g66) & (!g67) & (g68)) + ((!shiftx2x) & (shiftx3x) & (!g65) & (g66) & (g67) & (g68)) + ((!shiftx2x) & (shiftx3x) & (g65) & (!g66) & (!g67) & (g68)) + ((!shiftx2x) & (shiftx3x) & (g65) & (!g66) & (g67) & (g68)) + ((!shiftx2x) & (shiftx3x) & (g65) & (g66) & (!g67) & (g68)) + ((!shiftx2x) & (shiftx3x) & (g65) & (g66) & (g67) & (g68)) + ((shiftx2x) & (!shiftx3x) & (!g65) & (g66) & (!g67) & (!g68)) + ((shiftx2x) & (!shiftx3x) & (!g65) & (g66) & (!g67) & (g68)) + ((shiftx2x) & (!shiftx3x) & (!g65) & (g66) & (g67) & (!g68)) + ((shiftx2x) & (!shiftx3x) & (!g65) & (g66) & (g67) & (g68)) + ((shiftx2x) & (!shiftx3x) & (g65) & (g66) & (!g67) & (!g68)) + ((shiftx2x) & (!shiftx3x) & (g65) & (g66) & (!g67) & (g68)) + ((shiftx2x) & (!shiftx3x) & (g65) & (g66) & (g67) & (!g68)) + ((shiftx2x) & (!shiftx3x) & (g65) & (g66) & (g67) & (g68)) + ((shiftx2x) & (shiftx3x) & (!g65) & (!g66) & (g67) & (!g68)) + ((shiftx2x) & (shiftx3x) & (!g65) & (!g66) & (g67) & (g68)) + ((shiftx2x) & (shiftx3x) & (!g65) & (g66) & (g67) & (!g68)) + ((shiftx2x) & (shiftx3x) & (!g65) & (g66) & (g67) & (g68)) + ((shiftx2x) & (shiftx3x) & (g65) & (!g66) & (g67) & (!g68)) + ((shiftx2x) & (shiftx3x) & (g65) & (!g66) & (g67) & (g68)) + ((shiftx2x) & (shiftx3x) & (g65) & (g66) & (g67) & (!g68)) + ((shiftx2x) & (shiftx3x) & (g65) & (g66) & (g67) & (g68)));
	assign g70 = (((!shiftx0x) & (!shiftx1x) & (!ax96x) & (!ax95x) & (!ax94x) & (ax97x)) + ((!shiftx0x) & (!shiftx1x) & (!ax96x) & (!ax95x) & (ax94x) & (ax97x)) + ((!shiftx0x) & (!shiftx1x) & (!ax96x) & (ax95x) & (!ax94x) & (ax97x)) + ((!shiftx0x) & (!shiftx1x) & (!ax96x) & (ax95x) & (ax94x) & (ax97x)) + ((!shiftx0x) & (!shiftx1x) & (ax96x) & (!ax95x) & (!ax94x) & (ax97x)) + ((!shiftx0x) & (!shiftx1x) & (ax96x) & (!ax95x) & (ax94x) & (ax97x)) + ((!shiftx0x) & (!shiftx1x) & (ax96x) & (ax95x) & (!ax94x) & (ax97x)) + ((!shiftx0x) & (!shiftx1x) & (ax96x) & (ax95x) & (ax94x) & (ax97x)) + ((!shiftx0x) & (shiftx1x) & (!ax96x) & (ax95x) & (!ax94x) & (!ax97x)) + ((!shiftx0x) & (shiftx1x) & (!ax96x) & (ax95x) & (!ax94x) & (ax97x)) + ((!shiftx0x) & (shiftx1x) & (!ax96x) & (ax95x) & (ax94x) & (!ax97x)) + ((!shiftx0x) & (shiftx1x) & (!ax96x) & (ax95x) & (ax94x) & (ax97x)) + ((!shiftx0x) & (shiftx1x) & (ax96x) & (ax95x) & (!ax94x) & (!ax97x)) + ((!shiftx0x) & (shiftx1x) & (ax96x) & (ax95x) & (!ax94x) & (ax97x)) + ((!shiftx0x) & (shiftx1x) & (ax96x) & (ax95x) & (ax94x) & (!ax97x)) + ((!shiftx0x) & (shiftx1x) & (ax96x) & (ax95x) & (ax94x) & (ax97x)) + ((shiftx0x) & (!shiftx1x) & (ax96x) & (!ax95x) & (!ax94x) & (!ax97x)) + ((shiftx0x) & (!shiftx1x) & (ax96x) & (!ax95x) & (!ax94x) & (ax97x)) + ((shiftx0x) & (!shiftx1x) & (ax96x) & (!ax95x) & (ax94x) & (!ax97x)) + ((shiftx0x) & (!shiftx1x) & (ax96x) & (!ax95x) & (ax94x) & (ax97x)) + ((shiftx0x) & (!shiftx1x) & (ax96x) & (ax95x) & (!ax94x) & (!ax97x)) + ((shiftx0x) & (!shiftx1x) & (ax96x) & (ax95x) & (!ax94x) & (ax97x)) + ((shiftx0x) & (!shiftx1x) & (ax96x) & (ax95x) & (ax94x) & (!ax97x)) + ((shiftx0x) & (!shiftx1x) & (ax96x) & (ax95x) & (ax94x) & (ax97x)) + ((shiftx0x) & (shiftx1x) & (!ax96x) & (!ax95x) & (ax94x) & (!ax97x)) + ((shiftx0x) & (shiftx1x) & (!ax96x) & (!ax95x) & (ax94x) & (ax97x)) + ((shiftx0x) & (shiftx1x) & (!ax96x) & (ax95x) & (ax94x) & (!ax97x)) + ((shiftx0x) & (shiftx1x) & (!ax96x) & (ax95x) & (ax94x) & (ax97x)) + ((shiftx0x) & (shiftx1x) & (ax96x) & (!ax95x) & (ax94x) & (!ax97x)) + ((shiftx0x) & (shiftx1x) & (ax96x) & (!ax95x) & (ax94x) & (ax97x)) + ((shiftx0x) & (shiftx1x) & (ax96x) & (ax95x) & (ax94x) & (!ax97x)) + ((shiftx0x) & (shiftx1x) & (ax96x) & (ax95x) & (ax94x) & (ax97x)));
	assign g71 = (((!shiftx0x) & (!shiftx1x) & (ax93x) & (!ax92x) & (!ax91x) & (!ax90x)) + ((!shiftx0x) & (!shiftx1x) & (ax93x) & (!ax92x) & (!ax91x) & (ax90x)) + ((!shiftx0x) & (!shiftx1x) & (ax93x) & (!ax92x) & (ax91x) & (!ax90x)) + ((!shiftx0x) & (!shiftx1x) & (ax93x) & (!ax92x) & (ax91x) & (ax90x)) + ((!shiftx0x) & (!shiftx1x) & (ax93x) & (ax92x) & (!ax91x) & (!ax90x)) + ((!shiftx0x) & (!shiftx1x) & (ax93x) & (ax92x) & (!ax91x) & (ax90x)) + ((!shiftx0x) & (!shiftx1x) & (ax93x) & (ax92x) & (ax91x) & (!ax90x)) + ((!shiftx0x) & (!shiftx1x) & (ax93x) & (ax92x) & (ax91x) & (ax90x)) + ((!shiftx0x) & (shiftx1x) & (!ax93x) & (!ax92x) & (ax91x) & (!ax90x)) + ((!shiftx0x) & (shiftx1x) & (!ax93x) & (!ax92x) & (ax91x) & (ax90x)) + ((!shiftx0x) & (shiftx1x) & (!ax93x) & (ax92x) & (ax91x) & (!ax90x)) + ((!shiftx0x) & (shiftx1x) & (!ax93x) & (ax92x) & (ax91x) & (ax90x)) + ((!shiftx0x) & (shiftx1x) & (ax93x) & (!ax92x) & (ax91x) & (!ax90x)) + ((!shiftx0x) & (shiftx1x) & (ax93x) & (!ax92x) & (ax91x) & (ax90x)) + ((!shiftx0x) & (shiftx1x) & (ax93x) & (ax92x) & (ax91x) & (!ax90x)) + ((!shiftx0x) & (shiftx1x) & (ax93x) & (ax92x) & (ax91x) & (ax90x)) + ((shiftx0x) & (!shiftx1x) & (!ax93x) & (ax92x) & (!ax91x) & (!ax90x)) + ((shiftx0x) & (!shiftx1x) & (!ax93x) & (ax92x) & (!ax91x) & (ax90x)) + ((shiftx0x) & (!shiftx1x) & (!ax93x) & (ax92x) & (ax91x) & (!ax90x)) + ((shiftx0x) & (!shiftx1x) & (!ax93x) & (ax92x) & (ax91x) & (ax90x)) + ((shiftx0x) & (!shiftx1x) & (ax93x) & (ax92x) & (!ax91x) & (!ax90x)) + ((shiftx0x) & (!shiftx1x) & (ax93x) & (ax92x) & (!ax91x) & (ax90x)) + ((shiftx0x) & (!shiftx1x) & (ax93x) & (ax92x) & (ax91x) & (!ax90x)) + ((shiftx0x) & (!shiftx1x) & (ax93x) & (ax92x) & (ax91x) & (ax90x)) + ((shiftx0x) & (shiftx1x) & (!ax93x) & (!ax92x) & (!ax91x) & (ax90x)) + ((shiftx0x) & (shiftx1x) & (!ax93x) & (!ax92x) & (ax91x) & (ax90x)) + ((shiftx0x) & (shiftx1x) & (!ax93x) & (ax92x) & (!ax91x) & (ax90x)) + ((shiftx0x) & (shiftx1x) & (!ax93x) & (ax92x) & (ax91x) & (ax90x)) + ((shiftx0x) & (shiftx1x) & (ax93x) & (!ax92x) & (!ax91x) & (ax90x)) + ((shiftx0x) & (shiftx1x) & (ax93x) & (!ax92x) & (ax91x) & (ax90x)) + ((shiftx0x) & (shiftx1x) & (ax93x) & (ax92x) & (!ax91x) & (ax90x)) + ((shiftx0x) & (shiftx1x) & (ax93x) & (ax92x) & (ax91x) & (ax90x)));
	assign g72 = (((!shiftx0x) & (!shiftx1x) & (!ax84x) & (!ax83x) & (!ax82x) & (ax85x)) + ((!shiftx0x) & (!shiftx1x) & (!ax84x) & (!ax83x) & (ax82x) & (ax85x)) + ((!shiftx0x) & (!shiftx1x) & (!ax84x) & (ax83x) & (!ax82x) & (ax85x)) + ((!shiftx0x) & (!shiftx1x) & (!ax84x) & (ax83x) & (ax82x) & (ax85x)) + ((!shiftx0x) & (!shiftx1x) & (ax84x) & (!ax83x) & (!ax82x) & (ax85x)) + ((!shiftx0x) & (!shiftx1x) & (ax84x) & (!ax83x) & (ax82x) & (ax85x)) + ((!shiftx0x) & (!shiftx1x) & (ax84x) & (ax83x) & (!ax82x) & (ax85x)) + ((!shiftx0x) & (!shiftx1x) & (ax84x) & (ax83x) & (ax82x) & (ax85x)) + ((!shiftx0x) & (shiftx1x) & (!ax84x) & (ax83x) & (!ax82x) & (!ax85x)) + ((!shiftx0x) & (shiftx1x) & (!ax84x) & (ax83x) & (!ax82x) & (ax85x)) + ((!shiftx0x) & (shiftx1x) & (!ax84x) & (ax83x) & (ax82x) & (!ax85x)) + ((!shiftx0x) & (shiftx1x) & (!ax84x) & (ax83x) & (ax82x) & (ax85x)) + ((!shiftx0x) & (shiftx1x) & (ax84x) & (ax83x) & (!ax82x) & (!ax85x)) + ((!shiftx0x) & (shiftx1x) & (ax84x) & (ax83x) & (!ax82x) & (ax85x)) + ((!shiftx0x) & (shiftx1x) & (ax84x) & (ax83x) & (ax82x) & (!ax85x)) + ((!shiftx0x) & (shiftx1x) & (ax84x) & (ax83x) & (ax82x) & (ax85x)) + ((shiftx0x) & (!shiftx1x) & (ax84x) & (!ax83x) & (!ax82x) & (!ax85x)) + ((shiftx0x) & (!shiftx1x) & (ax84x) & (!ax83x) & (!ax82x) & (ax85x)) + ((shiftx0x) & (!shiftx1x) & (ax84x) & (!ax83x) & (ax82x) & (!ax85x)) + ((shiftx0x) & (!shiftx1x) & (ax84x) & (!ax83x) & (ax82x) & (ax85x)) + ((shiftx0x) & (!shiftx1x) & (ax84x) & (ax83x) & (!ax82x) & (!ax85x)) + ((shiftx0x) & (!shiftx1x) & (ax84x) & (ax83x) & (!ax82x) & (ax85x)) + ((shiftx0x) & (!shiftx1x) & (ax84x) & (ax83x) & (ax82x) & (!ax85x)) + ((shiftx0x) & (!shiftx1x) & (ax84x) & (ax83x) & (ax82x) & (ax85x)) + ((shiftx0x) & (shiftx1x) & (!ax84x) & (!ax83x) & (ax82x) & (!ax85x)) + ((shiftx0x) & (shiftx1x) & (!ax84x) & (!ax83x) & (ax82x) & (ax85x)) + ((shiftx0x) & (shiftx1x) & (!ax84x) & (ax83x) & (ax82x) & (!ax85x)) + ((shiftx0x) & (shiftx1x) & (!ax84x) & (ax83x) & (ax82x) & (ax85x)) + ((shiftx0x) & (shiftx1x) & (ax84x) & (!ax83x) & (ax82x) & (!ax85x)) + ((shiftx0x) & (shiftx1x) & (ax84x) & (!ax83x) & (ax82x) & (ax85x)) + ((shiftx0x) & (shiftx1x) & (ax84x) & (ax83x) & (ax82x) & (!ax85x)) + ((shiftx0x) & (shiftx1x) & (ax84x) & (ax83x) & (ax82x) & (ax85x)));
	assign g73 = (((!shiftx0x) & (!shiftx1x) & (ax89x) & (!ax88x) & (!ax87x) & (!ax86x)) + ((!shiftx0x) & (!shiftx1x) & (ax89x) & (!ax88x) & (!ax87x) & (ax86x)) + ((!shiftx0x) & (!shiftx1x) & (ax89x) & (!ax88x) & (ax87x) & (!ax86x)) + ((!shiftx0x) & (!shiftx1x) & (ax89x) & (!ax88x) & (ax87x) & (ax86x)) + ((!shiftx0x) & (!shiftx1x) & (ax89x) & (ax88x) & (!ax87x) & (!ax86x)) + ((!shiftx0x) & (!shiftx1x) & (ax89x) & (ax88x) & (!ax87x) & (ax86x)) + ((!shiftx0x) & (!shiftx1x) & (ax89x) & (ax88x) & (ax87x) & (!ax86x)) + ((!shiftx0x) & (!shiftx1x) & (ax89x) & (ax88x) & (ax87x) & (ax86x)) + ((!shiftx0x) & (shiftx1x) & (!ax89x) & (!ax88x) & (ax87x) & (!ax86x)) + ((!shiftx0x) & (shiftx1x) & (!ax89x) & (!ax88x) & (ax87x) & (ax86x)) + ((!shiftx0x) & (shiftx1x) & (!ax89x) & (ax88x) & (ax87x) & (!ax86x)) + ((!shiftx0x) & (shiftx1x) & (!ax89x) & (ax88x) & (ax87x) & (ax86x)) + ((!shiftx0x) & (shiftx1x) & (ax89x) & (!ax88x) & (ax87x) & (!ax86x)) + ((!shiftx0x) & (shiftx1x) & (ax89x) & (!ax88x) & (ax87x) & (ax86x)) + ((!shiftx0x) & (shiftx1x) & (ax89x) & (ax88x) & (ax87x) & (!ax86x)) + ((!shiftx0x) & (shiftx1x) & (ax89x) & (ax88x) & (ax87x) & (ax86x)) + ((shiftx0x) & (!shiftx1x) & (!ax89x) & (ax88x) & (!ax87x) & (!ax86x)) + ((shiftx0x) & (!shiftx1x) & (!ax89x) & (ax88x) & (!ax87x) & (ax86x)) + ((shiftx0x) & (!shiftx1x) & (!ax89x) & (ax88x) & (ax87x) & (!ax86x)) + ((shiftx0x) & (!shiftx1x) & (!ax89x) & (ax88x) & (ax87x) & (ax86x)) + ((shiftx0x) & (!shiftx1x) & (ax89x) & (ax88x) & (!ax87x) & (!ax86x)) + ((shiftx0x) & (!shiftx1x) & (ax89x) & (ax88x) & (!ax87x) & (ax86x)) + ((shiftx0x) & (!shiftx1x) & (ax89x) & (ax88x) & (ax87x) & (!ax86x)) + ((shiftx0x) & (!shiftx1x) & (ax89x) & (ax88x) & (ax87x) & (ax86x)) + ((shiftx0x) & (shiftx1x) & (!ax89x) & (!ax88x) & (!ax87x) & (ax86x)) + ((shiftx0x) & (shiftx1x) & (!ax89x) & (!ax88x) & (ax87x) & (ax86x)) + ((shiftx0x) & (shiftx1x) & (!ax89x) & (ax88x) & (!ax87x) & (ax86x)) + ((shiftx0x) & (shiftx1x) & (!ax89x) & (ax88x) & (ax87x) & (ax86x)) + ((shiftx0x) & (shiftx1x) & (ax89x) & (!ax88x) & (!ax87x) & (ax86x)) + ((shiftx0x) & (shiftx1x) & (ax89x) & (!ax88x) & (ax87x) & (ax86x)) + ((shiftx0x) & (shiftx1x) & (ax89x) & (ax88x) & (!ax87x) & (ax86x)) + ((shiftx0x) & (shiftx1x) & (ax89x) & (ax88x) & (ax87x) & (ax86x)));
	assign g74 = (((!shiftx2x) & (!shiftx3x) & (g70) & (!g71) & (!g72) & (!g73)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (!g71) & (!g72) & (g73)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (!g71) & (g72) & (!g73)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (!g71) & (g72) & (g73)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (g71) & (!g72) & (!g73)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (g71) & (!g72) & (g73)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (g71) & (g72) & (!g73)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (g71) & (g72) & (g73)) + ((!shiftx2x) & (shiftx3x) & (!g70) & (!g71) & (!g72) & (g73)) + ((!shiftx2x) & (shiftx3x) & (!g70) & (!g71) & (g72) & (g73)) + ((!shiftx2x) & (shiftx3x) & (!g70) & (g71) & (!g72) & (g73)) + ((!shiftx2x) & (shiftx3x) & (!g70) & (g71) & (g72) & (g73)) + ((!shiftx2x) & (shiftx3x) & (g70) & (!g71) & (!g72) & (g73)) + ((!shiftx2x) & (shiftx3x) & (g70) & (!g71) & (g72) & (g73)) + ((!shiftx2x) & (shiftx3x) & (g70) & (g71) & (!g72) & (g73)) + ((!shiftx2x) & (shiftx3x) & (g70) & (g71) & (g72) & (g73)) + ((shiftx2x) & (!shiftx3x) & (!g70) & (g71) & (!g72) & (!g73)) + ((shiftx2x) & (!shiftx3x) & (!g70) & (g71) & (!g72) & (g73)) + ((shiftx2x) & (!shiftx3x) & (!g70) & (g71) & (g72) & (!g73)) + ((shiftx2x) & (!shiftx3x) & (!g70) & (g71) & (g72) & (g73)) + ((shiftx2x) & (!shiftx3x) & (g70) & (g71) & (!g72) & (!g73)) + ((shiftx2x) & (!shiftx3x) & (g70) & (g71) & (!g72) & (g73)) + ((shiftx2x) & (!shiftx3x) & (g70) & (g71) & (g72) & (!g73)) + ((shiftx2x) & (!shiftx3x) & (g70) & (g71) & (g72) & (g73)) + ((shiftx2x) & (shiftx3x) & (!g70) & (!g71) & (g72) & (!g73)) + ((shiftx2x) & (shiftx3x) & (!g70) & (!g71) & (g72) & (g73)) + ((shiftx2x) & (shiftx3x) & (!g70) & (g71) & (g72) & (!g73)) + ((shiftx2x) & (shiftx3x) & (!g70) & (g71) & (g72) & (g73)) + ((shiftx2x) & (shiftx3x) & (g70) & (!g71) & (g72) & (!g73)) + ((shiftx2x) & (shiftx3x) & (g70) & (!g71) & (g72) & (g73)) + ((shiftx2x) & (shiftx3x) & (g70) & (g71) & (g72) & (!g73)) + ((shiftx2x) & (shiftx3x) & (g70) & (g71) & (g72) & (g73)));
	assign g75 = (((!shiftx0x) & (!shiftx1x) & (ax1x) & (!ax0x) & (!ax127x) & (!ax126x)) + ((!shiftx0x) & (!shiftx1x) & (ax1x) & (!ax0x) & (!ax127x) & (ax126x)) + ((!shiftx0x) & (!shiftx1x) & (ax1x) & (!ax0x) & (ax127x) & (!ax126x)) + ((!shiftx0x) & (!shiftx1x) & (ax1x) & (!ax0x) & (ax127x) & (ax126x)) + ((!shiftx0x) & (!shiftx1x) & (ax1x) & (ax0x) & (!ax127x) & (!ax126x)) + ((!shiftx0x) & (!shiftx1x) & (ax1x) & (ax0x) & (!ax127x) & (ax126x)) + ((!shiftx0x) & (!shiftx1x) & (ax1x) & (ax0x) & (ax127x) & (!ax126x)) + ((!shiftx0x) & (!shiftx1x) & (ax1x) & (ax0x) & (ax127x) & (ax126x)) + ((!shiftx0x) & (shiftx1x) & (!ax1x) & (!ax0x) & (ax127x) & (!ax126x)) + ((!shiftx0x) & (shiftx1x) & (!ax1x) & (!ax0x) & (ax127x) & (ax126x)) + ((!shiftx0x) & (shiftx1x) & (!ax1x) & (ax0x) & (ax127x) & (!ax126x)) + ((!shiftx0x) & (shiftx1x) & (!ax1x) & (ax0x) & (ax127x) & (ax126x)) + ((!shiftx0x) & (shiftx1x) & (ax1x) & (!ax0x) & (ax127x) & (!ax126x)) + ((!shiftx0x) & (shiftx1x) & (ax1x) & (!ax0x) & (ax127x) & (ax126x)) + ((!shiftx0x) & (shiftx1x) & (ax1x) & (ax0x) & (ax127x) & (!ax126x)) + ((!shiftx0x) & (shiftx1x) & (ax1x) & (ax0x) & (ax127x) & (ax126x)) + ((shiftx0x) & (!shiftx1x) & (!ax1x) & (ax0x) & (!ax127x) & (!ax126x)) + ((shiftx0x) & (!shiftx1x) & (!ax1x) & (ax0x) & (!ax127x) & (ax126x)) + ((shiftx0x) & (!shiftx1x) & (!ax1x) & (ax0x) & (ax127x) & (!ax126x)) + ((shiftx0x) & (!shiftx1x) & (!ax1x) & (ax0x) & (ax127x) & (ax126x)) + ((shiftx0x) & (!shiftx1x) & (ax1x) & (ax0x) & (!ax127x) & (!ax126x)) + ((shiftx0x) & (!shiftx1x) & (ax1x) & (ax0x) & (!ax127x) & (ax126x)) + ((shiftx0x) & (!shiftx1x) & (ax1x) & (ax0x) & (ax127x) & (!ax126x)) + ((shiftx0x) & (!shiftx1x) & (ax1x) & (ax0x) & (ax127x) & (ax126x)) + ((shiftx0x) & (shiftx1x) & (!ax1x) & (!ax0x) & (!ax127x) & (ax126x)) + ((shiftx0x) & (shiftx1x) & (!ax1x) & (!ax0x) & (ax127x) & (ax126x)) + ((shiftx0x) & (shiftx1x) & (!ax1x) & (ax0x) & (!ax127x) & (ax126x)) + ((shiftx0x) & (shiftx1x) & (!ax1x) & (ax0x) & (ax127x) & (ax126x)) + ((shiftx0x) & (shiftx1x) & (ax1x) & (!ax0x) & (!ax127x) & (ax126x)) + ((shiftx0x) & (shiftx1x) & (ax1x) & (!ax0x) & (ax127x) & (ax126x)) + ((shiftx0x) & (shiftx1x) & (ax1x) & (ax0x) & (!ax127x) & (ax126x)) + ((shiftx0x) & (shiftx1x) & (ax1x) & (ax0x) & (ax127x) & (ax126x)));
	assign g76 = (((!shiftx0x) & (!shiftx1x) & (ax125x) & (!ax124x) & (!ax123x) & (!ax122x)) + ((!shiftx0x) & (!shiftx1x) & (ax125x) & (!ax124x) & (!ax123x) & (ax122x)) + ((!shiftx0x) & (!shiftx1x) & (ax125x) & (!ax124x) & (ax123x) & (!ax122x)) + ((!shiftx0x) & (!shiftx1x) & (ax125x) & (!ax124x) & (ax123x) & (ax122x)) + ((!shiftx0x) & (!shiftx1x) & (ax125x) & (ax124x) & (!ax123x) & (!ax122x)) + ((!shiftx0x) & (!shiftx1x) & (ax125x) & (ax124x) & (!ax123x) & (ax122x)) + ((!shiftx0x) & (!shiftx1x) & (ax125x) & (ax124x) & (ax123x) & (!ax122x)) + ((!shiftx0x) & (!shiftx1x) & (ax125x) & (ax124x) & (ax123x) & (ax122x)) + ((!shiftx0x) & (shiftx1x) & (!ax125x) & (!ax124x) & (ax123x) & (!ax122x)) + ((!shiftx0x) & (shiftx1x) & (!ax125x) & (!ax124x) & (ax123x) & (ax122x)) + ((!shiftx0x) & (shiftx1x) & (!ax125x) & (ax124x) & (ax123x) & (!ax122x)) + ((!shiftx0x) & (shiftx1x) & (!ax125x) & (ax124x) & (ax123x) & (ax122x)) + ((!shiftx0x) & (shiftx1x) & (ax125x) & (!ax124x) & (ax123x) & (!ax122x)) + ((!shiftx0x) & (shiftx1x) & (ax125x) & (!ax124x) & (ax123x) & (ax122x)) + ((!shiftx0x) & (shiftx1x) & (ax125x) & (ax124x) & (ax123x) & (!ax122x)) + ((!shiftx0x) & (shiftx1x) & (ax125x) & (ax124x) & (ax123x) & (ax122x)) + ((shiftx0x) & (!shiftx1x) & (!ax125x) & (ax124x) & (!ax123x) & (!ax122x)) + ((shiftx0x) & (!shiftx1x) & (!ax125x) & (ax124x) & (!ax123x) & (ax122x)) + ((shiftx0x) & (!shiftx1x) & (!ax125x) & (ax124x) & (ax123x) & (!ax122x)) + ((shiftx0x) & (!shiftx1x) & (!ax125x) & (ax124x) & (ax123x) & (ax122x)) + ((shiftx0x) & (!shiftx1x) & (ax125x) & (ax124x) & (!ax123x) & (!ax122x)) + ((shiftx0x) & (!shiftx1x) & (ax125x) & (ax124x) & (!ax123x) & (ax122x)) + ((shiftx0x) & (!shiftx1x) & (ax125x) & (ax124x) & (ax123x) & (!ax122x)) + ((shiftx0x) & (!shiftx1x) & (ax125x) & (ax124x) & (ax123x) & (ax122x)) + ((shiftx0x) & (shiftx1x) & (!ax125x) & (!ax124x) & (!ax123x) & (ax122x)) + ((shiftx0x) & (shiftx1x) & (!ax125x) & (!ax124x) & (ax123x) & (ax122x)) + ((shiftx0x) & (shiftx1x) & (!ax125x) & (ax124x) & (!ax123x) & (ax122x)) + ((shiftx0x) & (shiftx1x) & (!ax125x) & (ax124x) & (ax123x) & (ax122x)) + ((shiftx0x) & (shiftx1x) & (ax125x) & (!ax124x) & (!ax123x) & (ax122x)) + ((shiftx0x) & (shiftx1x) & (ax125x) & (!ax124x) & (ax123x) & (ax122x)) + ((shiftx0x) & (shiftx1x) & (ax125x) & (ax124x) & (!ax123x) & (ax122x)) + ((shiftx0x) & (shiftx1x) & (ax125x) & (ax124x) & (ax123x) & (ax122x)));
	assign g77 = (((!shiftx0x) & (!shiftx1x) & (!ax116x) & (!ax115x) & (!ax114x) & (ax117x)) + ((!shiftx0x) & (!shiftx1x) & (!ax116x) & (!ax115x) & (ax114x) & (ax117x)) + ((!shiftx0x) & (!shiftx1x) & (!ax116x) & (ax115x) & (!ax114x) & (ax117x)) + ((!shiftx0x) & (!shiftx1x) & (!ax116x) & (ax115x) & (ax114x) & (ax117x)) + ((!shiftx0x) & (!shiftx1x) & (ax116x) & (!ax115x) & (!ax114x) & (ax117x)) + ((!shiftx0x) & (!shiftx1x) & (ax116x) & (!ax115x) & (ax114x) & (ax117x)) + ((!shiftx0x) & (!shiftx1x) & (ax116x) & (ax115x) & (!ax114x) & (ax117x)) + ((!shiftx0x) & (!shiftx1x) & (ax116x) & (ax115x) & (ax114x) & (ax117x)) + ((!shiftx0x) & (shiftx1x) & (!ax116x) & (ax115x) & (!ax114x) & (!ax117x)) + ((!shiftx0x) & (shiftx1x) & (!ax116x) & (ax115x) & (!ax114x) & (ax117x)) + ((!shiftx0x) & (shiftx1x) & (!ax116x) & (ax115x) & (ax114x) & (!ax117x)) + ((!shiftx0x) & (shiftx1x) & (!ax116x) & (ax115x) & (ax114x) & (ax117x)) + ((!shiftx0x) & (shiftx1x) & (ax116x) & (ax115x) & (!ax114x) & (!ax117x)) + ((!shiftx0x) & (shiftx1x) & (ax116x) & (ax115x) & (!ax114x) & (ax117x)) + ((!shiftx0x) & (shiftx1x) & (ax116x) & (ax115x) & (ax114x) & (!ax117x)) + ((!shiftx0x) & (shiftx1x) & (ax116x) & (ax115x) & (ax114x) & (ax117x)) + ((shiftx0x) & (!shiftx1x) & (ax116x) & (!ax115x) & (!ax114x) & (!ax117x)) + ((shiftx0x) & (!shiftx1x) & (ax116x) & (!ax115x) & (!ax114x) & (ax117x)) + ((shiftx0x) & (!shiftx1x) & (ax116x) & (!ax115x) & (ax114x) & (!ax117x)) + ((shiftx0x) & (!shiftx1x) & (ax116x) & (!ax115x) & (ax114x) & (ax117x)) + ((shiftx0x) & (!shiftx1x) & (ax116x) & (ax115x) & (!ax114x) & (!ax117x)) + ((shiftx0x) & (!shiftx1x) & (ax116x) & (ax115x) & (!ax114x) & (ax117x)) + ((shiftx0x) & (!shiftx1x) & (ax116x) & (ax115x) & (ax114x) & (!ax117x)) + ((shiftx0x) & (!shiftx1x) & (ax116x) & (ax115x) & (ax114x) & (ax117x)) + ((shiftx0x) & (shiftx1x) & (!ax116x) & (!ax115x) & (ax114x) & (!ax117x)) + ((shiftx0x) & (shiftx1x) & (!ax116x) & (!ax115x) & (ax114x) & (ax117x)) + ((shiftx0x) & (shiftx1x) & (!ax116x) & (ax115x) & (ax114x) & (!ax117x)) + ((shiftx0x) & (shiftx1x) & (!ax116x) & (ax115x) & (ax114x) & (ax117x)) + ((shiftx0x) & (shiftx1x) & (ax116x) & (!ax115x) & (ax114x) & (!ax117x)) + ((shiftx0x) & (shiftx1x) & (ax116x) & (!ax115x) & (ax114x) & (ax117x)) + ((shiftx0x) & (shiftx1x) & (ax116x) & (ax115x) & (ax114x) & (!ax117x)) + ((shiftx0x) & (shiftx1x) & (ax116x) & (ax115x) & (ax114x) & (ax117x)));
	assign g78 = (((!shiftx0x) & (!shiftx1x) & (ax121x) & (!ax120x) & (!ax119x) & (!ax118x)) + ((!shiftx0x) & (!shiftx1x) & (ax121x) & (!ax120x) & (!ax119x) & (ax118x)) + ((!shiftx0x) & (!shiftx1x) & (ax121x) & (!ax120x) & (ax119x) & (!ax118x)) + ((!shiftx0x) & (!shiftx1x) & (ax121x) & (!ax120x) & (ax119x) & (ax118x)) + ((!shiftx0x) & (!shiftx1x) & (ax121x) & (ax120x) & (!ax119x) & (!ax118x)) + ((!shiftx0x) & (!shiftx1x) & (ax121x) & (ax120x) & (!ax119x) & (ax118x)) + ((!shiftx0x) & (!shiftx1x) & (ax121x) & (ax120x) & (ax119x) & (!ax118x)) + ((!shiftx0x) & (!shiftx1x) & (ax121x) & (ax120x) & (ax119x) & (ax118x)) + ((!shiftx0x) & (shiftx1x) & (!ax121x) & (!ax120x) & (ax119x) & (!ax118x)) + ((!shiftx0x) & (shiftx1x) & (!ax121x) & (!ax120x) & (ax119x) & (ax118x)) + ((!shiftx0x) & (shiftx1x) & (!ax121x) & (ax120x) & (ax119x) & (!ax118x)) + ((!shiftx0x) & (shiftx1x) & (!ax121x) & (ax120x) & (ax119x) & (ax118x)) + ((!shiftx0x) & (shiftx1x) & (ax121x) & (!ax120x) & (ax119x) & (!ax118x)) + ((!shiftx0x) & (shiftx1x) & (ax121x) & (!ax120x) & (ax119x) & (ax118x)) + ((!shiftx0x) & (shiftx1x) & (ax121x) & (ax120x) & (ax119x) & (!ax118x)) + ((!shiftx0x) & (shiftx1x) & (ax121x) & (ax120x) & (ax119x) & (ax118x)) + ((shiftx0x) & (!shiftx1x) & (!ax121x) & (ax120x) & (!ax119x) & (!ax118x)) + ((shiftx0x) & (!shiftx1x) & (!ax121x) & (ax120x) & (!ax119x) & (ax118x)) + ((shiftx0x) & (!shiftx1x) & (!ax121x) & (ax120x) & (ax119x) & (!ax118x)) + ((shiftx0x) & (!shiftx1x) & (!ax121x) & (ax120x) & (ax119x) & (ax118x)) + ((shiftx0x) & (!shiftx1x) & (ax121x) & (ax120x) & (!ax119x) & (!ax118x)) + ((shiftx0x) & (!shiftx1x) & (ax121x) & (ax120x) & (!ax119x) & (ax118x)) + ((shiftx0x) & (!shiftx1x) & (ax121x) & (ax120x) & (ax119x) & (!ax118x)) + ((shiftx0x) & (!shiftx1x) & (ax121x) & (ax120x) & (ax119x) & (ax118x)) + ((shiftx0x) & (shiftx1x) & (!ax121x) & (!ax120x) & (!ax119x) & (ax118x)) + ((shiftx0x) & (shiftx1x) & (!ax121x) & (!ax120x) & (ax119x) & (ax118x)) + ((shiftx0x) & (shiftx1x) & (!ax121x) & (ax120x) & (!ax119x) & (ax118x)) + ((shiftx0x) & (shiftx1x) & (!ax121x) & (ax120x) & (ax119x) & (ax118x)) + ((shiftx0x) & (shiftx1x) & (ax121x) & (!ax120x) & (!ax119x) & (ax118x)) + ((shiftx0x) & (shiftx1x) & (ax121x) & (!ax120x) & (ax119x) & (ax118x)) + ((shiftx0x) & (shiftx1x) & (ax121x) & (ax120x) & (!ax119x) & (ax118x)) + ((shiftx0x) & (shiftx1x) & (ax121x) & (ax120x) & (ax119x) & (ax118x)));
	assign g79 = (((!shiftx2x) & (!shiftx3x) & (g75) & (!g76) & (!g77) & (!g78)) + ((!shiftx2x) & (!shiftx3x) & (g75) & (!g76) & (!g77) & (g78)) + ((!shiftx2x) & (!shiftx3x) & (g75) & (!g76) & (g77) & (!g78)) + ((!shiftx2x) & (!shiftx3x) & (g75) & (!g76) & (g77) & (g78)) + ((!shiftx2x) & (!shiftx3x) & (g75) & (g76) & (!g77) & (!g78)) + ((!shiftx2x) & (!shiftx3x) & (g75) & (g76) & (!g77) & (g78)) + ((!shiftx2x) & (!shiftx3x) & (g75) & (g76) & (g77) & (!g78)) + ((!shiftx2x) & (!shiftx3x) & (g75) & (g76) & (g77) & (g78)) + ((!shiftx2x) & (shiftx3x) & (!g75) & (!g76) & (!g77) & (g78)) + ((!shiftx2x) & (shiftx3x) & (!g75) & (!g76) & (g77) & (g78)) + ((!shiftx2x) & (shiftx3x) & (!g75) & (g76) & (!g77) & (g78)) + ((!shiftx2x) & (shiftx3x) & (!g75) & (g76) & (g77) & (g78)) + ((!shiftx2x) & (shiftx3x) & (g75) & (!g76) & (!g77) & (g78)) + ((!shiftx2x) & (shiftx3x) & (g75) & (!g76) & (g77) & (g78)) + ((!shiftx2x) & (shiftx3x) & (g75) & (g76) & (!g77) & (g78)) + ((!shiftx2x) & (shiftx3x) & (g75) & (g76) & (g77) & (g78)) + ((shiftx2x) & (!shiftx3x) & (!g75) & (g76) & (!g77) & (!g78)) + ((shiftx2x) & (!shiftx3x) & (!g75) & (g76) & (!g77) & (g78)) + ((shiftx2x) & (!shiftx3x) & (!g75) & (g76) & (g77) & (!g78)) + ((shiftx2x) & (!shiftx3x) & (!g75) & (g76) & (g77) & (g78)) + ((shiftx2x) & (!shiftx3x) & (g75) & (g76) & (!g77) & (!g78)) + ((shiftx2x) & (!shiftx3x) & (g75) & (g76) & (!g77) & (g78)) + ((shiftx2x) & (!shiftx3x) & (g75) & (g76) & (g77) & (!g78)) + ((shiftx2x) & (!shiftx3x) & (g75) & (g76) & (g77) & (g78)) + ((shiftx2x) & (shiftx3x) & (!g75) & (!g76) & (g77) & (!g78)) + ((shiftx2x) & (shiftx3x) & (!g75) & (!g76) & (g77) & (g78)) + ((shiftx2x) & (shiftx3x) & (!g75) & (g76) & (g77) & (!g78)) + ((shiftx2x) & (shiftx3x) & (!g75) & (g76) & (g77) & (g78)) + ((shiftx2x) & (shiftx3x) & (g75) & (!g76) & (g77) & (!g78)) + ((shiftx2x) & (shiftx3x) & (g75) & (!g76) & (g77) & (g78)) + ((shiftx2x) & (shiftx3x) & (g75) & (g76) & (g77) & (!g78)) + ((shiftx2x) & (shiftx3x) & (g75) & (g76) & (g77) & (g78)));
	assign g80 = (((!shiftx0x) & (!shiftx1x) & (ax113x) & (!ax112x) & (!ax111x) & (!ax110x)) + ((!shiftx0x) & (!shiftx1x) & (ax113x) & (!ax112x) & (!ax111x) & (ax110x)) + ((!shiftx0x) & (!shiftx1x) & (ax113x) & (!ax112x) & (ax111x) & (!ax110x)) + ((!shiftx0x) & (!shiftx1x) & (ax113x) & (!ax112x) & (ax111x) & (ax110x)) + ((!shiftx0x) & (!shiftx1x) & (ax113x) & (ax112x) & (!ax111x) & (!ax110x)) + ((!shiftx0x) & (!shiftx1x) & (ax113x) & (ax112x) & (!ax111x) & (ax110x)) + ((!shiftx0x) & (!shiftx1x) & (ax113x) & (ax112x) & (ax111x) & (!ax110x)) + ((!shiftx0x) & (!shiftx1x) & (ax113x) & (ax112x) & (ax111x) & (ax110x)) + ((!shiftx0x) & (shiftx1x) & (!ax113x) & (!ax112x) & (ax111x) & (!ax110x)) + ((!shiftx0x) & (shiftx1x) & (!ax113x) & (!ax112x) & (ax111x) & (ax110x)) + ((!shiftx0x) & (shiftx1x) & (!ax113x) & (ax112x) & (ax111x) & (!ax110x)) + ((!shiftx0x) & (shiftx1x) & (!ax113x) & (ax112x) & (ax111x) & (ax110x)) + ((!shiftx0x) & (shiftx1x) & (ax113x) & (!ax112x) & (ax111x) & (!ax110x)) + ((!shiftx0x) & (shiftx1x) & (ax113x) & (!ax112x) & (ax111x) & (ax110x)) + ((!shiftx0x) & (shiftx1x) & (ax113x) & (ax112x) & (ax111x) & (!ax110x)) + ((!shiftx0x) & (shiftx1x) & (ax113x) & (ax112x) & (ax111x) & (ax110x)) + ((shiftx0x) & (!shiftx1x) & (!ax113x) & (ax112x) & (!ax111x) & (!ax110x)) + ((shiftx0x) & (!shiftx1x) & (!ax113x) & (ax112x) & (!ax111x) & (ax110x)) + ((shiftx0x) & (!shiftx1x) & (!ax113x) & (ax112x) & (ax111x) & (!ax110x)) + ((shiftx0x) & (!shiftx1x) & (!ax113x) & (ax112x) & (ax111x) & (ax110x)) + ((shiftx0x) & (!shiftx1x) & (ax113x) & (ax112x) & (!ax111x) & (!ax110x)) + ((shiftx0x) & (!shiftx1x) & (ax113x) & (ax112x) & (!ax111x) & (ax110x)) + ((shiftx0x) & (!shiftx1x) & (ax113x) & (ax112x) & (ax111x) & (!ax110x)) + ((shiftx0x) & (!shiftx1x) & (ax113x) & (ax112x) & (ax111x) & (ax110x)) + ((shiftx0x) & (shiftx1x) & (!ax113x) & (!ax112x) & (!ax111x) & (ax110x)) + ((shiftx0x) & (shiftx1x) & (!ax113x) & (!ax112x) & (ax111x) & (ax110x)) + ((shiftx0x) & (shiftx1x) & (!ax113x) & (ax112x) & (!ax111x) & (ax110x)) + ((shiftx0x) & (shiftx1x) & (!ax113x) & (ax112x) & (ax111x) & (ax110x)) + ((shiftx0x) & (shiftx1x) & (ax113x) & (!ax112x) & (!ax111x) & (ax110x)) + ((shiftx0x) & (shiftx1x) & (ax113x) & (!ax112x) & (ax111x) & (ax110x)) + ((shiftx0x) & (shiftx1x) & (ax113x) & (ax112x) & (!ax111x) & (ax110x)) + ((shiftx0x) & (shiftx1x) & (ax113x) & (ax112x) & (ax111x) & (ax110x)));
	assign g81 = (((!shiftx0x) & (!shiftx1x) & (ax109x) & (!ax108x) & (!ax107x) & (!ax106x)) + ((!shiftx0x) & (!shiftx1x) & (ax109x) & (!ax108x) & (!ax107x) & (ax106x)) + ((!shiftx0x) & (!shiftx1x) & (ax109x) & (!ax108x) & (ax107x) & (!ax106x)) + ((!shiftx0x) & (!shiftx1x) & (ax109x) & (!ax108x) & (ax107x) & (ax106x)) + ((!shiftx0x) & (!shiftx1x) & (ax109x) & (ax108x) & (!ax107x) & (!ax106x)) + ((!shiftx0x) & (!shiftx1x) & (ax109x) & (ax108x) & (!ax107x) & (ax106x)) + ((!shiftx0x) & (!shiftx1x) & (ax109x) & (ax108x) & (ax107x) & (!ax106x)) + ((!shiftx0x) & (!shiftx1x) & (ax109x) & (ax108x) & (ax107x) & (ax106x)) + ((!shiftx0x) & (shiftx1x) & (!ax109x) & (!ax108x) & (ax107x) & (!ax106x)) + ((!shiftx0x) & (shiftx1x) & (!ax109x) & (!ax108x) & (ax107x) & (ax106x)) + ((!shiftx0x) & (shiftx1x) & (!ax109x) & (ax108x) & (ax107x) & (!ax106x)) + ((!shiftx0x) & (shiftx1x) & (!ax109x) & (ax108x) & (ax107x) & (ax106x)) + ((!shiftx0x) & (shiftx1x) & (ax109x) & (!ax108x) & (ax107x) & (!ax106x)) + ((!shiftx0x) & (shiftx1x) & (ax109x) & (!ax108x) & (ax107x) & (ax106x)) + ((!shiftx0x) & (shiftx1x) & (ax109x) & (ax108x) & (ax107x) & (!ax106x)) + ((!shiftx0x) & (shiftx1x) & (ax109x) & (ax108x) & (ax107x) & (ax106x)) + ((shiftx0x) & (!shiftx1x) & (!ax109x) & (ax108x) & (!ax107x) & (!ax106x)) + ((shiftx0x) & (!shiftx1x) & (!ax109x) & (ax108x) & (!ax107x) & (ax106x)) + ((shiftx0x) & (!shiftx1x) & (!ax109x) & (ax108x) & (ax107x) & (!ax106x)) + ((shiftx0x) & (!shiftx1x) & (!ax109x) & (ax108x) & (ax107x) & (ax106x)) + ((shiftx0x) & (!shiftx1x) & (ax109x) & (ax108x) & (!ax107x) & (!ax106x)) + ((shiftx0x) & (!shiftx1x) & (ax109x) & (ax108x) & (!ax107x) & (ax106x)) + ((shiftx0x) & (!shiftx1x) & (ax109x) & (ax108x) & (ax107x) & (!ax106x)) + ((shiftx0x) & (!shiftx1x) & (ax109x) & (ax108x) & (ax107x) & (ax106x)) + ((shiftx0x) & (shiftx1x) & (!ax109x) & (!ax108x) & (!ax107x) & (ax106x)) + ((shiftx0x) & (shiftx1x) & (!ax109x) & (!ax108x) & (ax107x) & (ax106x)) + ((shiftx0x) & (shiftx1x) & (!ax109x) & (ax108x) & (!ax107x) & (ax106x)) + ((shiftx0x) & (shiftx1x) & (!ax109x) & (ax108x) & (ax107x) & (ax106x)) + ((shiftx0x) & (shiftx1x) & (ax109x) & (!ax108x) & (!ax107x) & (ax106x)) + ((shiftx0x) & (shiftx1x) & (ax109x) & (!ax108x) & (ax107x) & (ax106x)) + ((shiftx0x) & (shiftx1x) & (ax109x) & (ax108x) & (!ax107x) & (ax106x)) + ((shiftx0x) & (shiftx1x) & (ax109x) & (ax108x) & (ax107x) & (ax106x)));
	assign g82 = (((!shiftx0x) & (!shiftx1x) & (!ax100x) & (!ax99x) & (!ax98x) & (ax101x)) + ((!shiftx0x) & (!shiftx1x) & (!ax100x) & (!ax99x) & (ax98x) & (ax101x)) + ((!shiftx0x) & (!shiftx1x) & (!ax100x) & (ax99x) & (!ax98x) & (ax101x)) + ((!shiftx0x) & (!shiftx1x) & (!ax100x) & (ax99x) & (ax98x) & (ax101x)) + ((!shiftx0x) & (!shiftx1x) & (ax100x) & (!ax99x) & (!ax98x) & (ax101x)) + ((!shiftx0x) & (!shiftx1x) & (ax100x) & (!ax99x) & (ax98x) & (ax101x)) + ((!shiftx0x) & (!shiftx1x) & (ax100x) & (ax99x) & (!ax98x) & (ax101x)) + ((!shiftx0x) & (!shiftx1x) & (ax100x) & (ax99x) & (ax98x) & (ax101x)) + ((!shiftx0x) & (shiftx1x) & (!ax100x) & (ax99x) & (!ax98x) & (!ax101x)) + ((!shiftx0x) & (shiftx1x) & (!ax100x) & (ax99x) & (!ax98x) & (ax101x)) + ((!shiftx0x) & (shiftx1x) & (!ax100x) & (ax99x) & (ax98x) & (!ax101x)) + ((!shiftx0x) & (shiftx1x) & (!ax100x) & (ax99x) & (ax98x) & (ax101x)) + ((!shiftx0x) & (shiftx1x) & (ax100x) & (ax99x) & (!ax98x) & (!ax101x)) + ((!shiftx0x) & (shiftx1x) & (ax100x) & (ax99x) & (!ax98x) & (ax101x)) + ((!shiftx0x) & (shiftx1x) & (ax100x) & (ax99x) & (ax98x) & (!ax101x)) + ((!shiftx0x) & (shiftx1x) & (ax100x) & (ax99x) & (ax98x) & (ax101x)) + ((shiftx0x) & (!shiftx1x) & (ax100x) & (!ax99x) & (!ax98x) & (!ax101x)) + ((shiftx0x) & (!shiftx1x) & (ax100x) & (!ax99x) & (!ax98x) & (ax101x)) + ((shiftx0x) & (!shiftx1x) & (ax100x) & (!ax99x) & (ax98x) & (!ax101x)) + ((shiftx0x) & (!shiftx1x) & (ax100x) & (!ax99x) & (ax98x) & (ax101x)) + ((shiftx0x) & (!shiftx1x) & (ax100x) & (ax99x) & (!ax98x) & (!ax101x)) + ((shiftx0x) & (!shiftx1x) & (ax100x) & (ax99x) & (!ax98x) & (ax101x)) + ((shiftx0x) & (!shiftx1x) & (ax100x) & (ax99x) & (ax98x) & (!ax101x)) + ((shiftx0x) & (!shiftx1x) & (ax100x) & (ax99x) & (ax98x) & (ax101x)) + ((shiftx0x) & (shiftx1x) & (!ax100x) & (!ax99x) & (ax98x) & (!ax101x)) + ((shiftx0x) & (shiftx1x) & (!ax100x) & (!ax99x) & (ax98x) & (ax101x)) + ((shiftx0x) & (shiftx1x) & (!ax100x) & (ax99x) & (ax98x) & (!ax101x)) + ((shiftx0x) & (shiftx1x) & (!ax100x) & (ax99x) & (ax98x) & (ax101x)) + ((shiftx0x) & (shiftx1x) & (ax100x) & (!ax99x) & (ax98x) & (!ax101x)) + ((shiftx0x) & (shiftx1x) & (ax100x) & (!ax99x) & (ax98x) & (ax101x)) + ((shiftx0x) & (shiftx1x) & (ax100x) & (ax99x) & (ax98x) & (!ax101x)) + ((shiftx0x) & (shiftx1x) & (ax100x) & (ax99x) & (ax98x) & (ax101x)));
	assign g83 = (((!shiftx0x) & (!shiftx1x) & (ax105x) & (!ax104x) & (!ax103x) & (!ax102x)) + ((!shiftx0x) & (!shiftx1x) & (ax105x) & (!ax104x) & (!ax103x) & (ax102x)) + ((!shiftx0x) & (!shiftx1x) & (ax105x) & (!ax104x) & (ax103x) & (!ax102x)) + ((!shiftx0x) & (!shiftx1x) & (ax105x) & (!ax104x) & (ax103x) & (ax102x)) + ((!shiftx0x) & (!shiftx1x) & (ax105x) & (ax104x) & (!ax103x) & (!ax102x)) + ((!shiftx0x) & (!shiftx1x) & (ax105x) & (ax104x) & (!ax103x) & (ax102x)) + ((!shiftx0x) & (!shiftx1x) & (ax105x) & (ax104x) & (ax103x) & (!ax102x)) + ((!shiftx0x) & (!shiftx1x) & (ax105x) & (ax104x) & (ax103x) & (ax102x)) + ((!shiftx0x) & (shiftx1x) & (!ax105x) & (!ax104x) & (ax103x) & (!ax102x)) + ((!shiftx0x) & (shiftx1x) & (!ax105x) & (!ax104x) & (ax103x) & (ax102x)) + ((!shiftx0x) & (shiftx1x) & (!ax105x) & (ax104x) & (ax103x) & (!ax102x)) + ((!shiftx0x) & (shiftx1x) & (!ax105x) & (ax104x) & (ax103x) & (ax102x)) + ((!shiftx0x) & (shiftx1x) & (ax105x) & (!ax104x) & (ax103x) & (!ax102x)) + ((!shiftx0x) & (shiftx1x) & (ax105x) & (!ax104x) & (ax103x) & (ax102x)) + ((!shiftx0x) & (shiftx1x) & (ax105x) & (ax104x) & (ax103x) & (!ax102x)) + ((!shiftx0x) & (shiftx1x) & (ax105x) & (ax104x) & (ax103x) & (ax102x)) + ((shiftx0x) & (!shiftx1x) & (!ax105x) & (ax104x) & (!ax103x) & (!ax102x)) + ((shiftx0x) & (!shiftx1x) & (!ax105x) & (ax104x) & (!ax103x) & (ax102x)) + ((shiftx0x) & (!shiftx1x) & (!ax105x) & (ax104x) & (ax103x) & (!ax102x)) + ((shiftx0x) & (!shiftx1x) & (!ax105x) & (ax104x) & (ax103x) & (ax102x)) + ((shiftx0x) & (!shiftx1x) & (ax105x) & (ax104x) & (!ax103x) & (!ax102x)) + ((shiftx0x) & (!shiftx1x) & (ax105x) & (ax104x) & (!ax103x) & (ax102x)) + ((shiftx0x) & (!shiftx1x) & (ax105x) & (ax104x) & (ax103x) & (!ax102x)) + ((shiftx0x) & (!shiftx1x) & (ax105x) & (ax104x) & (ax103x) & (ax102x)) + ((shiftx0x) & (shiftx1x) & (!ax105x) & (!ax104x) & (!ax103x) & (ax102x)) + ((shiftx0x) & (shiftx1x) & (!ax105x) & (!ax104x) & (ax103x) & (ax102x)) + ((shiftx0x) & (shiftx1x) & (!ax105x) & (ax104x) & (!ax103x) & (ax102x)) + ((shiftx0x) & (shiftx1x) & (!ax105x) & (ax104x) & (ax103x) & (ax102x)) + ((shiftx0x) & (shiftx1x) & (ax105x) & (!ax104x) & (!ax103x) & (ax102x)) + ((shiftx0x) & (shiftx1x) & (ax105x) & (!ax104x) & (ax103x) & (ax102x)) + ((shiftx0x) & (shiftx1x) & (ax105x) & (ax104x) & (!ax103x) & (ax102x)) + ((shiftx0x) & (shiftx1x) & (ax105x) & (ax104x) & (ax103x) & (ax102x)));
	assign g84 = (((!shiftx2x) & (!shiftx3x) & (g80) & (!g81) & (!g82) & (!g83)) + ((!shiftx2x) & (!shiftx3x) & (g80) & (!g81) & (!g82) & (g83)) + ((!shiftx2x) & (!shiftx3x) & (g80) & (!g81) & (g82) & (!g83)) + ((!shiftx2x) & (!shiftx3x) & (g80) & (!g81) & (g82) & (g83)) + ((!shiftx2x) & (!shiftx3x) & (g80) & (g81) & (!g82) & (!g83)) + ((!shiftx2x) & (!shiftx3x) & (g80) & (g81) & (!g82) & (g83)) + ((!shiftx2x) & (!shiftx3x) & (g80) & (g81) & (g82) & (!g83)) + ((!shiftx2x) & (!shiftx3x) & (g80) & (g81) & (g82) & (g83)) + ((!shiftx2x) & (shiftx3x) & (!g80) & (!g81) & (!g82) & (g83)) + ((!shiftx2x) & (shiftx3x) & (!g80) & (!g81) & (g82) & (g83)) + ((!shiftx2x) & (shiftx3x) & (!g80) & (g81) & (!g82) & (g83)) + ((!shiftx2x) & (shiftx3x) & (!g80) & (g81) & (g82) & (g83)) + ((!shiftx2x) & (shiftx3x) & (g80) & (!g81) & (!g82) & (g83)) + ((!shiftx2x) & (shiftx3x) & (g80) & (!g81) & (g82) & (g83)) + ((!shiftx2x) & (shiftx3x) & (g80) & (g81) & (!g82) & (g83)) + ((!shiftx2x) & (shiftx3x) & (g80) & (g81) & (g82) & (g83)) + ((shiftx2x) & (!shiftx3x) & (!g80) & (g81) & (!g82) & (!g83)) + ((shiftx2x) & (!shiftx3x) & (!g80) & (g81) & (!g82) & (g83)) + ((shiftx2x) & (!shiftx3x) & (!g80) & (g81) & (g82) & (!g83)) + ((shiftx2x) & (!shiftx3x) & (!g80) & (g81) & (g82) & (g83)) + ((shiftx2x) & (!shiftx3x) & (g80) & (g81) & (!g82) & (!g83)) + ((shiftx2x) & (!shiftx3x) & (g80) & (g81) & (!g82) & (g83)) + ((shiftx2x) & (!shiftx3x) & (g80) & (g81) & (g82) & (!g83)) + ((shiftx2x) & (!shiftx3x) & (g80) & (g81) & (g82) & (g83)) + ((shiftx2x) & (shiftx3x) & (!g80) & (!g81) & (g82) & (!g83)) + ((shiftx2x) & (shiftx3x) & (!g80) & (!g81) & (g82) & (g83)) + ((shiftx2x) & (shiftx3x) & (!g80) & (g81) & (g82) & (!g83)) + ((shiftx2x) & (shiftx3x) & (!g80) & (g81) & (g82) & (g83)) + ((shiftx2x) & (shiftx3x) & (g80) & (!g81) & (g82) & (!g83)) + ((shiftx2x) & (shiftx3x) & (g80) & (!g81) & (g82) & (g83)) + ((shiftx2x) & (shiftx3x) & (g80) & (g81) & (g82) & (!g83)) + ((shiftx2x) & (shiftx3x) & (g80) & (g81) & (g82) & (g83)));
	assign g85 = (((!shiftx4x) & (!shiftx5x) & (!g69) & (!g74) & (g79) & (!g84)) + ((!shiftx4x) & (!shiftx5x) & (!g69) & (!g74) & (g79) & (g84)) + ((!shiftx4x) & (!shiftx5x) & (!g69) & (g74) & (g79) & (!g84)) + ((!shiftx4x) & (!shiftx5x) & (!g69) & (g74) & (g79) & (g84)) + ((!shiftx4x) & (!shiftx5x) & (g69) & (!g74) & (g79) & (!g84)) + ((!shiftx4x) & (!shiftx5x) & (g69) & (!g74) & (g79) & (g84)) + ((!shiftx4x) & (!shiftx5x) & (g69) & (g74) & (g79) & (!g84)) + ((!shiftx4x) & (!shiftx5x) & (g69) & (g74) & (g79) & (g84)) + ((!shiftx4x) & (shiftx5x) & (!g69) & (g74) & (!g79) & (!g84)) + ((!shiftx4x) & (shiftx5x) & (!g69) & (g74) & (!g79) & (g84)) + ((!shiftx4x) & (shiftx5x) & (!g69) & (g74) & (g79) & (!g84)) + ((!shiftx4x) & (shiftx5x) & (!g69) & (g74) & (g79) & (g84)) + ((!shiftx4x) & (shiftx5x) & (g69) & (g74) & (!g79) & (!g84)) + ((!shiftx4x) & (shiftx5x) & (g69) & (g74) & (!g79) & (g84)) + ((!shiftx4x) & (shiftx5x) & (g69) & (g74) & (g79) & (!g84)) + ((!shiftx4x) & (shiftx5x) & (g69) & (g74) & (g79) & (g84)) + ((shiftx4x) & (!shiftx5x) & (!g69) & (!g74) & (!g79) & (g84)) + ((shiftx4x) & (!shiftx5x) & (!g69) & (!g74) & (g79) & (g84)) + ((shiftx4x) & (!shiftx5x) & (!g69) & (g74) & (!g79) & (g84)) + ((shiftx4x) & (!shiftx5x) & (!g69) & (g74) & (g79) & (g84)) + ((shiftx4x) & (!shiftx5x) & (g69) & (!g74) & (!g79) & (g84)) + ((shiftx4x) & (!shiftx5x) & (g69) & (!g74) & (g79) & (g84)) + ((shiftx4x) & (!shiftx5x) & (g69) & (g74) & (!g79) & (g84)) + ((shiftx4x) & (!shiftx5x) & (g69) & (g74) & (g79) & (g84)) + ((shiftx4x) & (shiftx5x) & (g69) & (!g74) & (!g79) & (!g84)) + ((shiftx4x) & (shiftx5x) & (g69) & (!g74) & (!g79) & (g84)) + ((shiftx4x) & (shiftx5x) & (g69) & (!g74) & (g79) & (!g84)) + ((shiftx4x) & (shiftx5x) & (g69) & (!g74) & (g79) & (g84)) + ((shiftx4x) & (shiftx5x) & (g69) & (g74) & (!g79) & (!g84)) + ((shiftx4x) & (shiftx5x) & (g69) & (g74) & (!g79) & (g84)) + ((shiftx4x) & (shiftx5x) & (g69) & (g74) & (g79) & (!g84)) + ((shiftx4x) & (shiftx5x) & (g69) & (g74) & (g79) & (g84)));
	assign resultx1x = (((!sk[85]) & (shiftx6x) & (!g64) & (!g85)) + ((!sk[85]) & (shiftx6x) & (!g64) & (g85)) + ((!sk[85]) & (shiftx6x) & (g64) & (!g85)) + ((!sk[85]) & (shiftx6x) & (g64) & (g85)) + ((sk[85]) & (!shiftx6x) & (!g64) & (g85)) + ((sk[85]) & (!shiftx6x) & (g64) & (g85)) + ((sk[85]) & (shiftx6x) & (g64) & (!g85)) + ((sk[85]) & (shiftx6x) & (g64) & (g85)));
	assign g87 = (((!ax66x) & (!ax65x) & (!ax64x) & (ax63x) & (shiftx0x) & (shiftx1x)) + ((!ax66x) & (!ax65x) & (ax64x) & (!ax63x) & (!shiftx0x) & (shiftx1x)) + ((!ax66x) & (!ax65x) & (ax64x) & (ax63x) & (!shiftx0x) & (shiftx1x)) + ((!ax66x) & (!ax65x) & (ax64x) & (ax63x) & (shiftx0x) & (shiftx1x)) + ((!ax66x) & (ax65x) & (!ax64x) & (!ax63x) & (shiftx0x) & (!shiftx1x)) + ((!ax66x) & (ax65x) & (!ax64x) & (ax63x) & (shiftx0x) & (!shiftx1x)) + ((!ax66x) & (ax65x) & (!ax64x) & (ax63x) & (shiftx0x) & (shiftx1x)) + ((!ax66x) & (ax65x) & (ax64x) & (!ax63x) & (!shiftx0x) & (shiftx1x)) + ((!ax66x) & (ax65x) & (ax64x) & (!ax63x) & (shiftx0x) & (!shiftx1x)) + ((!ax66x) & (ax65x) & (ax64x) & (ax63x) & (!shiftx0x) & (shiftx1x)) + ((!ax66x) & (ax65x) & (ax64x) & (ax63x) & (shiftx0x) & (!shiftx1x)) + ((!ax66x) & (ax65x) & (ax64x) & (ax63x) & (shiftx0x) & (shiftx1x)) + ((ax66x) & (!ax65x) & (!ax64x) & (!ax63x) & (!shiftx0x) & (!shiftx1x)) + ((ax66x) & (!ax65x) & (!ax64x) & (ax63x) & (!shiftx0x) & (!shiftx1x)) + ((ax66x) & (!ax65x) & (!ax64x) & (ax63x) & (shiftx0x) & (shiftx1x)) + ((ax66x) & (!ax65x) & (ax64x) & (!ax63x) & (!shiftx0x) & (!shiftx1x)) + ((ax66x) & (!ax65x) & (ax64x) & (!ax63x) & (!shiftx0x) & (shiftx1x)) + ((ax66x) & (!ax65x) & (ax64x) & (ax63x) & (!shiftx0x) & (!shiftx1x)) + ((ax66x) & (!ax65x) & (ax64x) & (ax63x) & (!shiftx0x) & (shiftx1x)) + ((ax66x) & (!ax65x) & (ax64x) & (ax63x) & (shiftx0x) & (shiftx1x)) + ((ax66x) & (ax65x) & (!ax64x) & (!ax63x) & (!shiftx0x) & (!shiftx1x)) + ((ax66x) & (ax65x) & (!ax64x) & (!ax63x) & (shiftx0x) & (!shiftx1x)) + ((ax66x) & (ax65x) & (!ax64x) & (ax63x) & (!shiftx0x) & (!shiftx1x)) + ((ax66x) & (ax65x) & (!ax64x) & (ax63x) & (shiftx0x) & (!shiftx1x)) + ((ax66x) & (ax65x) & (!ax64x) & (ax63x) & (shiftx0x) & (shiftx1x)) + ((ax66x) & (ax65x) & (ax64x) & (!ax63x) & (!shiftx0x) & (!shiftx1x)) + ((ax66x) & (ax65x) & (ax64x) & (!ax63x) & (!shiftx0x) & (shiftx1x)) + ((ax66x) & (ax65x) & (ax64x) & (!ax63x) & (shiftx0x) & (!shiftx1x)) + ((ax66x) & (ax65x) & (ax64x) & (ax63x) & (!shiftx0x) & (!shiftx1x)) + ((ax66x) & (ax65x) & (ax64x) & (ax63x) & (!shiftx0x) & (shiftx1x)) + ((ax66x) & (ax65x) & (ax64x) & (ax63x) & (shiftx0x) & (!shiftx1x)) + ((ax66x) & (ax65x) & (ax64x) & (ax63x) & (shiftx0x) & (shiftx1x)));
	assign g88 = (((!ax62x) & (!ax61x) & (!ax60x) & (ax59x) & (shiftx0x) & (shiftx1x)) + ((!ax62x) & (!ax61x) & (ax60x) & (!ax59x) & (!shiftx0x) & (shiftx1x)) + ((!ax62x) & (!ax61x) & (ax60x) & (ax59x) & (!shiftx0x) & (shiftx1x)) + ((!ax62x) & (!ax61x) & (ax60x) & (ax59x) & (shiftx0x) & (shiftx1x)) + ((!ax62x) & (ax61x) & (!ax60x) & (!ax59x) & (shiftx0x) & (!shiftx1x)) + ((!ax62x) & (ax61x) & (!ax60x) & (ax59x) & (shiftx0x) & (!shiftx1x)) + ((!ax62x) & (ax61x) & (!ax60x) & (ax59x) & (shiftx0x) & (shiftx1x)) + ((!ax62x) & (ax61x) & (ax60x) & (!ax59x) & (!shiftx0x) & (shiftx1x)) + ((!ax62x) & (ax61x) & (ax60x) & (!ax59x) & (shiftx0x) & (!shiftx1x)) + ((!ax62x) & (ax61x) & (ax60x) & (ax59x) & (!shiftx0x) & (shiftx1x)) + ((!ax62x) & (ax61x) & (ax60x) & (ax59x) & (shiftx0x) & (!shiftx1x)) + ((!ax62x) & (ax61x) & (ax60x) & (ax59x) & (shiftx0x) & (shiftx1x)) + ((ax62x) & (!ax61x) & (!ax60x) & (!ax59x) & (!shiftx0x) & (!shiftx1x)) + ((ax62x) & (!ax61x) & (!ax60x) & (ax59x) & (!shiftx0x) & (!shiftx1x)) + ((ax62x) & (!ax61x) & (!ax60x) & (ax59x) & (shiftx0x) & (shiftx1x)) + ((ax62x) & (!ax61x) & (ax60x) & (!ax59x) & (!shiftx0x) & (!shiftx1x)) + ((ax62x) & (!ax61x) & (ax60x) & (!ax59x) & (!shiftx0x) & (shiftx1x)) + ((ax62x) & (!ax61x) & (ax60x) & (ax59x) & (!shiftx0x) & (!shiftx1x)) + ((ax62x) & (!ax61x) & (ax60x) & (ax59x) & (!shiftx0x) & (shiftx1x)) + ((ax62x) & (!ax61x) & (ax60x) & (ax59x) & (shiftx0x) & (shiftx1x)) + ((ax62x) & (ax61x) & (!ax60x) & (!ax59x) & (!shiftx0x) & (!shiftx1x)) + ((ax62x) & (ax61x) & (!ax60x) & (!ax59x) & (shiftx0x) & (!shiftx1x)) + ((ax62x) & (ax61x) & (!ax60x) & (ax59x) & (!shiftx0x) & (!shiftx1x)) + ((ax62x) & (ax61x) & (!ax60x) & (ax59x) & (shiftx0x) & (!shiftx1x)) + ((ax62x) & (ax61x) & (!ax60x) & (ax59x) & (shiftx0x) & (shiftx1x)) + ((ax62x) & (ax61x) & (ax60x) & (!ax59x) & (!shiftx0x) & (!shiftx1x)) + ((ax62x) & (ax61x) & (ax60x) & (!ax59x) & (!shiftx0x) & (shiftx1x)) + ((ax62x) & (ax61x) & (ax60x) & (!ax59x) & (shiftx0x) & (!shiftx1x)) + ((ax62x) & (ax61x) & (ax60x) & (ax59x) & (!shiftx0x) & (!shiftx1x)) + ((ax62x) & (ax61x) & (ax60x) & (ax59x) & (!shiftx0x) & (shiftx1x)) + ((ax62x) & (ax61x) & (ax60x) & (ax59x) & (shiftx0x) & (!shiftx1x)) + ((ax62x) & (ax61x) & (ax60x) & (ax59x) & (shiftx0x) & (shiftx1x)));
	assign g89 = (((!ax54x) & (!ax53x) & (!ax52x) & (ax51x) & (shiftx0x) & (shiftx1x)) + ((!ax54x) & (!ax53x) & (ax52x) & (!ax51x) & (!shiftx0x) & (shiftx1x)) + ((!ax54x) & (!ax53x) & (ax52x) & (ax51x) & (!shiftx0x) & (shiftx1x)) + ((!ax54x) & (!ax53x) & (ax52x) & (ax51x) & (shiftx0x) & (shiftx1x)) + ((!ax54x) & (ax53x) & (!ax52x) & (!ax51x) & (shiftx0x) & (!shiftx1x)) + ((!ax54x) & (ax53x) & (!ax52x) & (ax51x) & (shiftx0x) & (!shiftx1x)) + ((!ax54x) & (ax53x) & (!ax52x) & (ax51x) & (shiftx0x) & (shiftx1x)) + ((!ax54x) & (ax53x) & (ax52x) & (!ax51x) & (!shiftx0x) & (shiftx1x)) + ((!ax54x) & (ax53x) & (ax52x) & (!ax51x) & (shiftx0x) & (!shiftx1x)) + ((!ax54x) & (ax53x) & (ax52x) & (ax51x) & (!shiftx0x) & (shiftx1x)) + ((!ax54x) & (ax53x) & (ax52x) & (ax51x) & (shiftx0x) & (!shiftx1x)) + ((!ax54x) & (ax53x) & (ax52x) & (ax51x) & (shiftx0x) & (shiftx1x)) + ((ax54x) & (!ax53x) & (!ax52x) & (!ax51x) & (!shiftx0x) & (!shiftx1x)) + ((ax54x) & (!ax53x) & (!ax52x) & (ax51x) & (!shiftx0x) & (!shiftx1x)) + ((ax54x) & (!ax53x) & (!ax52x) & (ax51x) & (shiftx0x) & (shiftx1x)) + ((ax54x) & (!ax53x) & (ax52x) & (!ax51x) & (!shiftx0x) & (!shiftx1x)) + ((ax54x) & (!ax53x) & (ax52x) & (!ax51x) & (!shiftx0x) & (shiftx1x)) + ((ax54x) & (!ax53x) & (ax52x) & (ax51x) & (!shiftx0x) & (!shiftx1x)) + ((ax54x) & (!ax53x) & (ax52x) & (ax51x) & (!shiftx0x) & (shiftx1x)) + ((ax54x) & (!ax53x) & (ax52x) & (ax51x) & (shiftx0x) & (shiftx1x)) + ((ax54x) & (ax53x) & (!ax52x) & (!ax51x) & (!shiftx0x) & (!shiftx1x)) + ((ax54x) & (ax53x) & (!ax52x) & (!ax51x) & (shiftx0x) & (!shiftx1x)) + ((ax54x) & (ax53x) & (!ax52x) & (ax51x) & (!shiftx0x) & (!shiftx1x)) + ((ax54x) & (ax53x) & (!ax52x) & (ax51x) & (shiftx0x) & (!shiftx1x)) + ((ax54x) & (ax53x) & (!ax52x) & (ax51x) & (shiftx0x) & (shiftx1x)) + ((ax54x) & (ax53x) & (ax52x) & (!ax51x) & (!shiftx0x) & (!shiftx1x)) + ((ax54x) & (ax53x) & (ax52x) & (!ax51x) & (!shiftx0x) & (shiftx1x)) + ((ax54x) & (ax53x) & (ax52x) & (!ax51x) & (shiftx0x) & (!shiftx1x)) + ((ax54x) & (ax53x) & (ax52x) & (ax51x) & (!shiftx0x) & (!shiftx1x)) + ((ax54x) & (ax53x) & (ax52x) & (ax51x) & (!shiftx0x) & (shiftx1x)) + ((ax54x) & (ax53x) & (ax52x) & (ax51x) & (shiftx0x) & (!shiftx1x)) + ((ax54x) & (ax53x) & (ax52x) & (ax51x) & (shiftx0x) & (shiftx1x)));
	assign g90 = (((!ax58x) & (!ax57x) & (!ax56x) & (ax55x) & (shiftx0x) & (shiftx1x)) + ((!ax58x) & (!ax57x) & (ax56x) & (!ax55x) & (!shiftx0x) & (shiftx1x)) + ((!ax58x) & (!ax57x) & (ax56x) & (ax55x) & (!shiftx0x) & (shiftx1x)) + ((!ax58x) & (!ax57x) & (ax56x) & (ax55x) & (shiftx0x) & (shiftx1x)) + ((!ax58x) & (ax57x) & (!ax56x) & (!ax55x) & (shiftx0x) & (!shiftx1x)) + ((!ax58x) & (ax57x) & (!ax56x) & (ax55x) & (shiftx0x) & (!shiftx1x)) + ((!ax58x) & (ax57x) & (!ax56x) & (ax55x) & (shiftx0x) & (shiftx1x)) + ((!ax58x) & (ax57x) & (ax56x) & (!ax55x) & (!shiftx0x) & (shiftx1x)) + ((!ax58x) & (ax57x) & (ax56x) & (!ax55x) & (shiftx0x) & (!shiftx1x)) + ((!ax58x) & (ax57x) & (ax56x) & (ax55x) & (!shiftx0x) & (shiftx1x)) + ((!ax58x) & (ax57x) & (ax56x) & (ax55x) & (shiftx0x) & (!shiftx1x)) + ((!ax58x) & (ax57x) & (ax56x) & (ax55x) & (shiftx0x) & (shiftx1x)) + ((ax58x) & (!ax57x) & (!ax56x) & (!ax55x) & (!shiftx0x) & (!shiftx1x)) + ((ax58x) & (!ax57x) & (!ax56x) & (ax55x) & (!shiftx0x) & (!shiftx1x)) + ((ax58x) & (!ax57x) & (!ax56x) & (ax55x) & (shiftx0x) & (shiftx1x)) + ((ax58x) & (!ax57x) & (ax56x) & (!ax55x) & (!shiftx0x) & (!shiftx1x)) + ((ax58x) & (!ax57x) & (ax56x) & (!ax55x) & (!shiftx0x) & (shiftx1x)) + ((ax58x) & (!ax57x) & (ax56x) & (ax55x) & (!shiftx0x) & (!shiftx1x)) + ((ax58x) & (!ax57x) & (ax56x) & (ax55x) & (!shiftx0x) & (shiftx1x)) + ((ax58x) & (!ax57x) & (ax56x) & (ax55x) & (shiftx0x) & (shiftx1x)) + ((ax58x) & (ax57x) & (!ax56x) & (!ax55x) & (!shiftx0x) & (!shiftx1x)) + ((ax58x) & (ax57x) & (!ax56x) & (!ax55x) & (shiftx0x) & (!shiftx1x)) + ((ax58x) & (ax57x) & (!ax56x) & (ax55x) & (!shiftx0x) & (!shiftx1x)) + ((ax58x) & (ax57x) & (!ax56x) & (ax55x) & (shiftx0x) & (!shiftx1x)) + ((ax58x) & (ax57x) & (!ax56x) & (ax55x) & (shiftx0x) & (shiftx1x)) + ((ax58x) & (ax57x) & (ax56x) & (!ax55x) & (!shiftx0x) & (!shiftx1x)) + ((ax58x) & (ax57x) & (ax56x) & (!ax55x) & (!shiftx0x) & (shiftx1x)) + ((ax58x) & (ax57x) & (ax56x) & (!ax55x) & (shiftx0x) & (!shiftx1x)) + ((ax58x) & (ax57x) & (ax56x) & (ax55x) & (!shiftx0x) & (!shiftx1x)) + ((ax58x) & (ax57x) & (ax56x) & (ax55x) & (!shiftx0x) & (shiftx1x)) + ((ax58x) & (ax57x) & (ax56x) & (ax55x) & (shiftx0x) & (!shiftx1x)) + ((ax58x) & (ax57x) & (ax56x) & (ax55x) & (shiftx0x) & (shiftx1x)));
	assign g91 = (((!shiftx2x) & (!shiftx3x) & (g87) & (!g88) & (!g89) & (!g90)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (!g88) & (!g89) & (g90)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (!g88) & (g89) & (!g90)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (!g88) & (g89) & (g90)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (g88) & (!g89) & (!g90)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (g88) & (!g89) & (g90)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (g88) & (g89) & (!g90)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (g88) & (g89) & (g90)) + ((!shiftx2x) & (shiftx3x) & (!g87) & (!g88) & (!g89) & (g90)) + ((!shiftx2x) & (shiftx3x) & (!g87) & (!g88) & (g89) & (g90)) + ((!shiftx2x) & (shiftx3x) & (!g87) & (g88) & (!g89) & (g90)) + ((!shiftx2x) & (shiftx3x) & (!g87) & (g88) & (g89) & (g90)) + ((!shiftx2x) & (shiftx3x) & (g87) & (!g88) & (!g89) & (g90)) + ((!shiftx2x) & (shiftx3x) & (g87) & (!g88) & (g89) & (g90)) + ((!shiftx2x) & (shiftx3x) & (g87) & (g88) & (!g89) & (g90)) + ((!shiftx2x) & (shiftx3x) & (g87) & (g88) & (g89) & (g90)) + ((shiftx2x) & (!shiftx3x) & (!g87) & (g88) & (!g89) & (!g90)) + ((shiftx2x) & (!shiftx3x) & (!g87) & (g88) & (!g89) & (g90)) + ((shiftx2x) & (!shiftx3x) & (!g87) & (g88) & (g89) & (!g90)) + ((shiftx2x) & (!shiftx3x) & (!g87) & (g88) & (g89) & (g90)) + ((shiftx2x) & (!shiftx3x) & (g87) & (g88) & (!g89) & (!g90)) + ((shiftx2x) & (!shiftx3x) & (g87) & (g88) & (!g89) & (g90)) + ((shiftx2x) & (!shiftx3x) & (g87) & (g88) & (g89) & (!g90)) + ((shiftx2x) & (!shiftx3x) & (g87) & (g88) & (g89) & (g90)) + ((shiftx2x) & (shiftx3x) & (!g87) & (!g88) & (g89) & (!g90)) + ((shiftx2x) & (shiftx3x) & (!g87) & (!g88) & (g89) & (g90)) + ((shiftx2x) & (shiftx3x) & (!g87) & (g88) & (g89) & (!g90)) + ((shiftx2x) & (shiftx3x) & (!g87) & (g88) & (g89) & (g90)) + ((shiftx2x) & (shiftx3x) & (g87) & (!g88) & (g89) & (!g90)) + ((shiftx2x) & (shiftx3x) & (g87) & (!g88) & (g89) & (g90)) + ((shiftx2x) & (shiftx3x) & (g87) & (g88) & (g89) & (!g90)) + ((shiftx2x) & (shiftx3x) & (g87) & (g88) & (g89) & (g90)));
	assign g92 = (((!ax18x) & (!ax17x) & (!ax16x) & (ax15x) & (shiftx0x) & (shiftx1x)) + ((!ax18x) & (!ax17x) & (ax16x) & (!ax15x) & (!shiftx0x) & (shiftx1x)) + ((!ax18x) & (!ax17x) & (ax16x) & (ax15x) & (!shiftx0x) & (shiftx1x)) + ((!ax18x) & (!ax17x) & (ax16x) & (ax15x) & (shiftx0x) & (shiftx1x)) + ((!ax18x) & (ax17x) & (!ax16x) & (!ax15x) & (shiftx0x) & (!shiftx1x)) + ((!ax18x) & (ax17x) & (!ax16x) & (ax15x) & (shiftx0x) & (!shiftx1x)) + ((!ax18x) & (ax17x) & (!ax16x) & (ax15x) & (shiftx0x) & (shiftx1x)) + ((!ax18x) & (ax17x) & (ax16x) & (!ax15x) & (!shiftx0x) & (shiftx1x)) + ((!ax18x) & (ax17x) & (ax16x) & (!ax15x) & (shiftx0x) & (!shiftx1x)) + ((!ax18x) & (ax17x) & (ax16x) & (ax15x) & (!shiftx0x) & (shiftx1x)) + ((!ax18x) & (ax17x) & (ax16x) & (ax15x) & (shiftx0x) & (!shiftx1x)) + ((!ax18x) & (ax17x) & (ax16x) & (ax15x) & (shiftx0x) & (shiftx1x)) + ((ax18x) & (!ax17x) & (!ax16x) & (!ax15x) & (!shiftx0x) & (!shiftx1x)) + ((ax18x) & (!ax17x) & (!ax16x) & (ax15x) & (!shiftx0x) & (!shiftx1x)) + ((ax18x) & (!ax17x) & (!ax16x) & (ax15x) & (shiftx0x) & (shiftx1x)) + ((ax18x) & (!ax17x) & (ax16x) & (!ax15x) & (!shiftx0x) & (!shiftx1x)) + ((ax18x) & (!ax17x) & (ax16x) & (!ax15x) & (!shiftx0x) & (shiftx1x)) + ((ax18x) & (!ax17x) & (ax16x) & (ax15x) & (!shiftx0x) & (!shiftx1x)) + ((ax18x) & (!ax17x) & (ax16x) & (ax15x) & (!shiftx0x) & (shiftx1x)) + ((ax18x) & (!ax17x) & (ax16x) & (ax15x) & (shiftx0x) & (shiftx1x)) + ((ax18x) & (ax17x) & (!ax16x) & (!ax15x) & (!shiftx0x) & (!shiftx1x)) + ((ax18x) & (ax17x) & (!ax16x) & (!ax15x) & (shiftx0x) & (!shiftx1x)) + ((ax18x) & (ax17x) & (!ax16x) & (ax15x) & (!shiftx0x) & (!shiftx1x)) + ((ax18x) & (ax17x) & (!ax16x) & (ax15x) & (shiftx0x) & (!shiftx1x)) + ((ax18x) & (ax17x) & (!ax16x) & (ax15x) & (shiftx0x) & (shiftx1x)) + ((ax18x) & (ax17x) & (ax16x) & (!ax15x) & (!shiftx0x) & (!shiftx1x)) + ((ax18x) & (ax17x) & (ax16x) & (!ax15x) & (!shiftx0x) & (shiftx1x)) + ((ax18x) & (ax17x) & (ax16x) & (!ax15x) & (shiftx0x) & (!shiftx1x)) + ((ax18x) & (ax17x) & (ax16x) & (ax15x) & (!shiftx0x) & (!shiftx1x)) + ((ax18x) & (ax17x) & (ax16x) & (ax15x) & (!shiftx0x) & (shiftx1x)) + ((ax18x) & (ax17x) & (ax16x) & (ax15x) & (shiftx0x) & (!shiftx1x)) + ((ax18x) & (ax17x) & (ax16x) & (ax15x) & (shiftx0x) & (shiftx1x)));
	assign g93 = (((!ax14x) & (!ax13x) & (!ax12x) & (ax11x) & (shiftx0x) & (shiftx1x)) + ((!ax14x) & (!ax13x) & (ax12x) & (!ax11x) & (!shiftx0x) & (shiftx1x)) + ((!ax14x) & (!ax13x) & (ax12x) & (ax11x) & (!shiftx0x) & (shiftx1x)) + ((!ax14x) & (!ax13x) & (ax12x) & (ax11x) & (shiftx0x) & (shiftx1x)) + ((!ax14x) & (ax13x) & (!ax12x) & (!ax11x) & (shiftx0x) & (!shiftx1x)) + ((!ax14x) & (ax13x) & (!ax12x) & (ax11x) & (shiftx0x) & (!shiftx1x)) + ((!ax14x) & (ax13x) & (!ax12x) & (ax11x) & (shiftx0x) & (shiftx1x)) + ((!ax14x) & (ax13x) & (ax12x) & (!ax11x) & (!shiftx0x) & (shiftx1x)) + ((!ax14x) & (ax13x) & (ax12x) & (!ax11x) & (shiftx0x) & (!shiftx1x)) + ((!ax14x) & (ax13x) & (ax12x) & (ax11x) & (!shiftx0x) & (shiftx1x)) + ((!ax14x) & (ax13x) & (ax12x) & (ax11x) & (shiftx0x) & (!shiftx1x)) + ((!ax14x) & (ax13x) & (ax12x) & (ax11x) & (shiftx0x) & (shiftx1x)) + ((ax14x) & (!ax13x) & (!ax12x) & (!ax11x) & (!shiftx0x) & (!shiftx1x)) + ((ax14x) & (!ax13x) & (!ax12x) & (ax11x) & (!shiftx0x) & (!shiftx1x)) + ((ax14x) & (!ax13x) & (!ax12x) & (ax11x) & (shiftx0x) & (shiftx1x)) + ((ax14x) & (!ax13x) & (ax12x) & (!ax11x) & (!shiftx0x) & (!shiftx1x)) + ((ax14x) & (!ax13x) & (ax12x) & (!ax11x) & (!shiftx0x) & (shiftx1x)) + ((ax14x) & (!ax13x) & (ax12x) & (ax11x) & (!shiftx0x) & (!shiftx1x)) + ((ax14x) & (!ax13x) & (ax12x) & (ax11x) & (!shiftx0x) & (shiftx1x)) + ((ax14x) & (!ax13x) & (ax12x) & (ax11x) & (shiftx0x) & (shiftx1x)) + ((ax14x) & (ax13x) & (!ax12x) & (!ax11x) & (!shiftx0x) & (!shiftx1x)) + ((ax14x) & (ax13x) & (!ax12x) & (!ax11x) & (shiftx0x) & (!shiftx1x)) + ((ax14x) & (ax13x) & (!ax12x) & (ax11x) & (!shiftx0x) & (!shiftx1x)) + ((ax14x) & (ax13x) & (!ax12x) & (ax11x) & (shiftx0x) & (!shiftx1x)) + ((ax14x) & (ax13x) & (!ax12x) & (ax11x) & (shiftx0x) & (shiftx1x)) + ((ax14x) & (ax13x) & (ax12x) & (!ax11x) & (!shiftx0x) & (!shiftx1x)) + ((ax14x) & (ax13x) & (ax12x) & (!ax11x) & (!shiftx0x) & (shiftx1x)) + ((ax14x) & (ax13x) & (ax12x) & (!ax11x) & (shiftx0x) & (!shiftx1x)) + ((ax14x) & (ax13x) & (ax12x) & (ax11x) & (!shiftx0x) & (!shiftx1x)) + ((ax14x) & (ax13x) & (ax12x) & (ax11x) & (!shiftx0x) & (shiftx1x)) + ((ax14x) & (ax13x) & (ax12x) & (ax11x) & (shiftx0x) & (!shiftx1x)) + ((ax14x) & (ax13x) & (ax12x) & (ax11x) & (shiftx0x) & (shiftx1x)));
	assign g94 = (((!ax6x) & (!ax5x) & (!ax4x) & (ax3x) & (shiftx0x) & (shiftx1x)) + ((!ax6x) & (!ax5x) & (ax4x) & (!ax3x) & (!shiftx0x) & (shiftx1x)) + ((!ax6x) & (!ax5x) & (ax4x) & (ax3x) & (!shiftx0x) & (shiftx1x)) + ((!ax6x) & (!ax5x) & (ax4x) & (ax3x) & (shiftx0x) & (shiftx1x)) + ((!ax6x) & (ax5x) & (!ax4x) & (!ax3x) & (shiftx0x) & (!shiftx1x)) + ((!ax6x) & (ax5x) & (!ax4x) & (ax3x) & (shiftx0x) & (!shiftx1x)) + ((!ax6x) & (ax5x) & (!ax4x) & (ax3x) & (shiftx0x) & (shiftx1x)) + ((!ax6x) & (ax5x) & (ax4x) & (!ax3x) & (!shiftx0x) & (shiftx1x)) + ((!ax6x) & (ax5x) & (ax4x) & (!ax3x) & (shiftx0x) & (!shiftx1x)) + ((!ax6x) & (ax5x) & (ax4x) & (ax3x) & (!shiftx0x) & (shiftx1x)) + ((!ax6x) & (ax5x) & (ax4x) & (ax3x) & (shiftx0x) & (!shiftx1x)) + ((!ax6x) & (ax5x) & (ax4x) & (ax3x) & (shiftx0x) & (shiftx1x)) + ((ax6x) & (!ax5x) & (!ax4x) & (!ax3x) & (!shiftx0x) & (!shiftx1x)) + ((ax6x) & (!ax5x) & (!ax4x) & (ax3x) & (!shiftx0x) & (!shiftx1x)) + ((ax6x) & (!ax5x) & (!ax4x) & (ax3x) & (shiftx0x) & (shiftx1x)) + ((ax6x) & (!ax5x) & (ax4x) & (!ax3x) & (!shiftx0x) & (!shiftx1x)) + ((ax6x) & (!ax5x) & (ax4x) & (!ax3x) & (!shiftx0x) & (shiftx1x)) + ((ax6x) & (!ax5x) & (ax4x) & (ax3x) & (!shiftx0x) & (!shiftx1x)) + ((ax6x) & (!ax5x) & (ax4x) & (ax3x) & (!shiftx0x) & (shiftx1x)) + ((ax6x) & (!ax5x) & (ax4x) & (ax3x) & (shiftx0x) & (shiftx1x)) + ((ax6x) & (ax5x) & (!ax4x) & (!ax3x) & (!shiftx0x) & (!shiftx1x)) + ((ax6x) & (ax5x) & (!ax4x) & (!ax3x) & (shiftx0x) & (!shiftx1x)) + ((ax6x) & (ax5x) & (!ax4x) & (ax3x) & (!shiftx0x) & (!shiftx1x)) + ((ax6x) & (ax5x) & (!ax4x) & (ax3x) & (shiftx0x) & (!shiftx1x)) + ((ax6x) & (ax5x) & (!ax4x) & (ax3x) & (shiftx0x) & (shiftx1x)) + ((ax6x) & (ax5x) & (ax4x) & (!ax3x) & (!shiftx0x) & (!shiftx1x)) + ((ax6x) & (ax5x) & (ax4x) & (!ax3x) & (!shiftx0x) & (shiftx1x)) + ((ax6x) & (ax5x) & (ax4x) & (!ax3x) & (shiftx0x) & (!shiftx1x)) + ((ax6x) & (ax5x) & (ax4x) & (ax3x) & (!shiftx0x) & (!shiftx1x)) + ((ax6x) & (ax5x) & (ax4x) & (ax3x) & (!shiftx0x) & (shiftx1x)) + ((ax6x) & (ax5x) & (ax4x) & (ax3x) & (shiftx0x) & (!shiftx1x)) + ((ax6x) & (ax5x) & (ax4x) & (ax3x) & (shiftx0x) & (shiftx1x)));
	assign g95 = (((!ax10x) & (!ax9x) & (!ax8x) & (ax7x) & (shiftx0x) & (shiftx1x)) + ((!ax10x) & (!ax9x) & (ax8x) & (!ax7x) & (!shiftx0x) & (shiftx1x)) + ((!ax10x) & (!ax9x) & (ax8x) & (ax7x) & (!shiftx0x) & (shiftx1x)) + ((!ax10x) & (!ax9x) & (ax8x) & (ax7x) & (shiftx0x) & (shiftx1x)) + ((!ax10x) & (ax9x) & (!ax8x) & (!ax7x) & (shiftx0x) & (!shiftx1x)) + ((!ax10x) & (ax9x) & (!ax8x) & (ax7x) & (shiftx0x) & (!shiftx1x)) + ((!ax10x) & (ax9x) & (!ax8x) & (ax7x) & (shiftx0x) & (shiftx1x)) + ((!ax10x) & (ax9x) & (ax8x) & (!ax7x) & (!shiftx0x) & (shiftx1x)) + ((!ax10x) & (ax9x) & (ax8x) & (!ax7x) & (shiftx0x) & (!shiftx1x)) + ((!ax10x) & (ax9x) & (ax8x) & (ax7x) & (!shiftx0x) & (shiftx1x)) + ((!ax10x) & (ax9x) & (ax8x) & (ax7x) & (shiftx0x) & (!shiftx1x)) + ((!ax10x) & (ax9x) & (ax8x) & (ax7x) & (shiftx0x) & (shiftx1x)) + ((ax10x) & (!ax9x) & (!ax8x) & (!ax7x) & (!shiftx0x) & (!shiftx1x)) + ((ax10x) & (!ax9x) & (!ax8x) & (ax7x) & (!shiftx0x) & (!shiftx1x)) + ((ax10x) & (!ax9x) & (!ax8x) & (ax7x) & (shiftx0x) & (shiftx1x)) + ((ax10x) & (!ax9x) & (ax8x) & (!ax7x) & (!shiftx0x) & (!shiftx1x)) + ((ax10x) & (!ax9x) & (ax8x) & (!ax7x) & (!shiftx0x) & (shiftx1x)) + ((ax10x) & (!ax9x) & (ax8x) & (ax7x) & (!shiftx0x) & (!shiftx1x)) + ((ax10x) & (!ax9x) & (ax8x) & (ax7x) & (!shiftx0x) & (shiftx1x)) + ((ax10x) & (!ax9x) & (ax8x) & (ax7x) & (shiftx0x) & (shiftx1x)) + ((ax10x) & (ax9x) & (!ax8x) & (!ax7x) & (!shiftx0x) & (!shiftx1x)) + ((ax10x) & (ax9x) & (!ax8x) & (!ax7x) & (shiftx0x) & (!shiftx1x)) + ((ax10x) & (ax9x) & (!ax8x) & (ax7x) & (!shiftx0x) & (!shiftx1x)) + ((ax10x) & (ax9x) & (!ax8x) & (ax7x) & (shiftx0x) & (!shiftx1x)) + ((ax10x) & (ax9x) & (!ax8x) & (ax7x) & (shiftx0x) & (shiftx1x)) + ((ax10x) & (ax9x) & (ax8x) & (!ax7x) & (!shiftx0x) & (!shiftx1x)) + ((ax10x) & (ax9x) & (ax8x) & (!ax7x) & (!shiftx0x) & (shiftx1x)) + ((ax10x) & (ax9x) & (ax8x) & (!ax7x) & (shiftx0x) & (!shiftx1x)) + ((ax10x) & (ax9x) & (ax8x) & (ax7x) & (!shiftx0x) & (!shiftx1x)) + ((ax10x) & (ax9x) & (ax8x) & (ax7x) & (!shiftx0x) & (shiftx1x)) + ((ax10x) & (ax9x) & (ax8x) & (ax7x) & (shiftx0x) & (!shiftx1x)) + ((ax10x) & (ax9x) & (ax8x) & (ax7x) & (shiftx0x) & (shiftx1x)));
	assign g96 = (((!shiftx2x) & (!shiftx3x) & (g92) & (!g93) & (!g94) & (!g95)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (!g93) & (!g94) & (g95)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (!g93) & (g94) & (!g95)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (!g93) & (g94) & (g95)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (g93) & (!g94) & (!g95)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (g93) & (!g94) & (g95)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (g93) & (g94) & (!g95)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (g93) & (g94) & (g95)) + ((!shiftx2x) & (shiftx3x) & (!g92) & (!g93) & (!g94) & (g95)) + ((!shiftx2x) & (shiftx3x) & (!g92) & (!g93) & (g94) & (g95)) + ((!shiftx2x) & (shiftx3x) & (!g92) & (g93) & (!g94) & (g95)) + ((!shiftx2x) & (shiftx3x) & (!g92) & (g93) & (g94) & (g95)) + ((!shiftx2x) & (shiftx3x) & (g92) & (!g93) & (!g94) & (g95)) + ((!shiftx2x) & (shiftx3x) & (g92) & (!g93) & (g94) & (g95)) + ((!shiftx2x) & (shiftx3x) & (g92) & (g93) & (!g94) & (g95)) + ((!shiftx2x) & (shiftx3x) & (g92) & (g93) & (g94) & (g95)) + ((shiftx2x) & (!shiftx3x) & (!g92) & (g93) & (!g94) & (!g95)) + ((shiftx2x) & (!shiftx3x) & (!g92) & (g93) & (!g94) & (g95)) + ((shiftx2x) & (!shiftx3x) & (!g92) & (g93) & (g94) & (!g95)) + ((shiftx2x) & (!shiftx3x) & (!g92) & (g93) & (g94) & (g95)) + ((shiftx2x) & (!shiftx3x) & (g92) & (g93) & (!g94) & (!g95)) + ((shiftx2x) & (!shiftx3x) & (g92) & (g93) & (!g94) & (g95)) + ((shiftx2x) & (!shiftx3x) & (g92) & (g93) & (g94) & (!g95)) + ((shiftx2x) & (!shiftx3x) & (g92) & (g93) & (g94) & (g95)) + ((shiftx2x) & (shiftx3x) & (!g92) & (!g93) & (g94) & (!g95)) + ((shiftx2x) & (shiftx3x) & (!g92) & (!g93) & (g94) & (g95)) + ((shiftx2x) & (shiftx3x) & (!g92) & (g93) & (g94) & (!g95)) + ((shiftx2x) & (shiftx3x) & (!g92) & (g93) & (g94) & (g95)) + ((shiftx2x) & (shiftx3x) & (g92) & (!g93) & (g94) & (!g95)) + ((shiftx2x) & (shiftx3x) & (g92) & (!g93) & (g94) & (g95)) + ((shiftx2x) & (shiftx3x) & (g92) & (g93) & (g94) & (!g95)) + ((shiftx2x) & (shiftx3x) & (g92) & (g93) & (g94) & (g95)));
	assign g97 = (((!ax50x) & (!ax49x) & (!ax48x) & (ax47x) & (shiftx0x) & (shiftx1x)) + ((!ax50x) & (!ax49x) & (ax48x) & (!ax47x) & (!shiftx0x) & (shiftx1x)) + ((!ax50x) & (!ax49x) & (ax48x) & (ax47x) & (!shiftx0x) & (shiftx1x)) + ((!ax50x) & (!ax49x) & (ax48x) & (ax47x) & (shiftx0x) & (shiftx1x)) + ((!ax50x) & (ax49x) & (!ax48x) & (!ax47x) & (shiftx0x) & (!shiftx1x)) + ((!ax50x) & (ax49x) & (!ax48x) & (ax47x) & (shiftx0x) & (!shiftx1x)) + ((!ax50x) & (ax49x) & (!ax48x) & (ax47x) & (shiftx0x) & (shiftx1x)) + ((!ax50x) & (ax49x) & (ax48x) & (!ax47x) & (!shiftx0x) & (shiftx1x)) + ((!ax50x) & (ax49x) & (ax48x) & (!ax47x) & (shiftx0x) & (!shiftx1x)) + ((!ax50x) & (ax49x) & (ax48x) & (ax47x) & (!shiftx0x) & (shiftx1x)) + ((!ax50x) & (ax49x) & (ax48x) & (ax47x) & (shiftx0x) & (!shiftx1x)) + ((!ax50x) & (ax49x) & (ax48x) & (ax47x) & (shiftx0x) & (shiftx1x)) + ((ax50x) & (!ax49x) & (!ax48x) & (!ax47x) & (!shiftx0x) & (!shiftx1x)) + ((ax50x) & (!ax49x) & (!ax48x) & (ax47x) & (!shiftx0x) & (!shiftx1x)) + ((ax50x) & (!ax49x) & (!ax48x) & (ax47x) & (shiftx0x) & (shiftx1x)) + ((ax50x) & (!ax49x) & (ax48x) & (!ax47x) & (!shiftx0x) & (!shiftx1x)) + ((ax50x) & (!ax49x) & (ax48x) & (!ax47x) & (!shiftx0x) & (shiftx1x)) + ((ax50x) & (!ax49x) & (ax48x) & (ax47x) & (!shiftx0x) & (!shiftx1x)) + ((ax50x) & (!ax49x) & (ax48x) & (ax47x) & (!shiftx0x) & (shiftx1x)) + ((ax50x) & (!ax49x) & (ax48x) & (ax47x) & (shiftx0x) & (shiftx1x)) + ((ax50x) & (ax49x) & (!ax48x) & (!ax47x) & (!shiftx0x) & (!shiftx1x)) + ((ax50x) & (ax49x) & (!ax48x) & (!ax47x) & (shiftx0x) & (!shiftx1x)) + ((ax50x) & (ax49x) & (!ax48x) & (ax47x) & (!shiftx0x) & (!shiftx1x)) + ((ax50x) & (ax49x) & (!ax48x) & (ax47x) & (shiftx0x) & (!shiftx1x)) + ((ax50x) & (ax49x) & (!ax48x) & (ax47x) & (shiftx0x) & (shiftx1x)) + ((ax50x) & (ax49x) & (ax48x) & (!ax47x) & (!shiftx0x) & (!shiftx1x)) + ((ax50x) & (ax49x) & (ax48x) & (!ax47x) & (!shiftx0x) & (shiftx1x)) + ((ax50x) & (ax49x) & (ax48x) & (!ax47x) & (shiftx0x) & (!shiftx1x)) + ((ax50x) & (ax49x) & (ax48x) & (ax47x) & (!shiftx0x) & (!shiftx1x)) + ((ax50x) & (ax49x) & (ax48x) & (ax47x) & (!shiftx0x) & (shiftx1x)) + ((ax50x) & (ax49x) & (ax48x) & (ax47x) & (shiftx0x) & (!shiftx1x)) + ((ax50x) & (ax49x) & (ax48x) & (ax47x) & (shiftx0x) & (shiftx1x)));
	assign g98 = (((!ax46x) & (!ax45x) & (!ax44x) & (ax43x) & (shiftx0x) & (shiftx1x)) + ((!ax46x) & (!ax45x) & (ax44x) & (!ax43x) & (!shiftx0x) & (shiftx1x)) + ((!ax46x) & (!ax45x) & (ax44x) & (ax43x) & (!shiftx0x) & (shiftx1x)) + ((!ax46x) & (!ax45x) & (ax44x) & (ax43x) & (shiftx0x) & (shiftx1x)) + ((!ax46x) & (ax45x) & (!ax44x) & (!ax43x) & (shiftx0x) & (!shiftx1x)) + ((!ax46x) & (ax45x) & (!ax44x) & (ax43x) & (shiftx0x) & (!shiftx1x)) + ((!ax46x) & (ax45x) & (!ax44x) & (ax43x) & (shiftx0x) & (shiftx1x)) + ((!ax46x) & (ax45x) & (ax44x) & (!ax43x) & (!shiftx0x) & (shiftx1x)) + ((!ax46x) & (ax45x) & (ax44x) & (!ax43x) & (shiftx0x) & (!shiftx1x)) + ((!ax46x) & (ax45x) & (ax44x) & (ax43x) & (!shiftx0x) & (shiftx1x)) + ((!ax46x) & (ax45x) & (ax44x) & (ax43x) & (shiftx0x) & (!shiftx1x)) + ((!ax46x) & (ax45x) & (ax44x) & (ax43x) & (shiftx0x) & (shiftx1x)) + ((ax46x) & (!ax45x) & (!ax44x) & (!ax43x) & (!shiftx0x) & (!shiftx1x)) + ((ax46x) & (!ax45x) & (!ax44x) & (ax43x) & (!shiftx0x) & (!shiftx1x)) + ((ax46x) & (!ax45x) & (!ax44x) & (ax43x) & (shiftx0x) & (shiftx1x)) + ((ax46x) & (!ax45x) & (ax44x) & (!ax43x) & (!shiftx0x) & (!shiftx1x)) + ((ax46x) & (!ax45x) & (ax44x) & (!ax43x) & (!shiftx0x) & (shiftx1x)) + ((ax46x) & (!ax45x) & (ax44x) & (ax43x) & (!shiftx0x) & (!shiftx1x)) + ((ax46x) & (!ax45x) & (ax44x) & (ax43x) & (!shiftx0x) & (shiftx1x)) + ((ax46x) & (!ax45x) & (ax44x) & (ax43x) & (shiftx0x) & (shiftx1x)) + ((ax46x) & (ax45x) & (!ax44x) & (!ax43x) & (!shiftx0x) & (!shiftx1x)) + ((ax46x) & (ax45x) & (!ax44x) & (!ax43x) & (shiftx0x) & (!shiftx1x)) + ((ax46x) & (ax45x) & (!ax44x) & (ax43x) & (!shiftx0x) & (!shiftx1x)) + ((ax46x) & (ax45x) & (!ax44x) & (ax43x) & (shiftx0x) & (!shiftx1x)) + ((ax46x) & (ax45x) & (!ax44x) & (ax43x) & (shiftx0x) & (shiftx1x)) + ((ax46x) & (ax45x) & (ax44x) & (!ax43x) & (!shiftx0x) & (!shiftx1x)) + ((ax46x) & (ax45x) & (ax44x) & (!ax43x) & (!shiftx0x) & (shiftx1x)) + ((ax46x) & (ax45x) & (ax44x) & (!ax43x) & (shiftx0x) & (!shiftx1x)) + ((ax46x) & (ax45x) & (ax44x) & (ax43x) & (!shiftx0x) & (!shiftx1x)) + ((ax46x) & (ax45x) & (ax44x) & (ax43x) & (!shiftx0x) & (shiftx1x)) + ((ax46x) & (ax45x) & (ax44x) & (ax43x) & (shiftx0x) & (!shiftx1x)) + ((ax46x) & (ax45x) & (ax44x) & (ax43x) & (shiftx0x) & (shiftx1x)));
	assign g99 = (((!ax38x) & (!ax37x) & (!ax36x) & (ax35x) & (shiftx0x) & (shiftx1x)) + ((!ax38x) & (!ax37x) & (ax36x) & (!ax35x) & (!shiftx0x) & (shiftx1x)) + ((!ax38x) & (!ax37x) & (ax36x) & (ax35x) & (!shiftx0x) & (shiftx1x)) + ((!ax38x) & (!ax37x) & (ax36x) & (ax35x) & (shiftx0x) & (shiftx1x)) + ((!ax38x) & (ax37x) & (!ax36x) & (!ax35x) & (shiftx0x) & (!shiftx1x)) + ((!ax38x) & (ax37x) & (!ax36x) & (ax35x) & (shiftx0x) & (!shiftx1x)) + ((!ax38x) & (ax37x) & (!ax36x) & (ax35x) & (shiftx0x) & (shiftx1x)) + ((!ax38x) & (ax37x) & (ax36x) & (!ax35x) & (!shiftx0x) & (shiftx1x)) + ((!ax38x) & (ax37x) & (ax36x) & (!ax35x) & (shiftx0x) & (!shiftx1x)) + ((!ax38x) & (ax37x) & (ax36x) & (ax35x) & (!shiftx0x) & (shiftx1x)) + ((!ax38x) & (ax37x) & (ax36x) & (ax35x) & (shiftx0x) & (!shiftx1x)) + ((!ax38x) & (ax37x) & (ax36x) & (ax35x) & (shiftx0x) & (shiftx1x)) + ((ax38x) & (!ax37x) & (!ax36x) & (!ax35x) & (!shiftx0x) & (!shiftx1x)) + ((ax38x) & (!ax37x) & (!ax36x) & (ax35x) & (!shiftx0x) & (!shiftx1x)) + ((ax38x) & (!ax37x) & (!ax36x) & (ax35x) & (shiftx0x) & (shiftx1x)) + ((ax38x) & (!ax37x) & (ax36x) & (!ax35x) & (!shiftx0x) & (!shiftx1x)) + ((ax38x) & (!ax37x) & (ax36x) & (!ax35x) & (!shiftx0x) & (shiftx1x)) + ((ax38x) & (!ax37x) & (ax36x) & (ax35x) & (!shiftx0x) & (!shiftx1x)) + ((ax38x) & (!ax37x) & (ax36x) & (ax35x) & (!shiftx0x) & (shiftx1x)) + ((ax38x) & (!ax37x) & (ax36x) & (ax35x) & (shiftx0x) & (shiftx1x)) + ((ax38x) & (ax37x) & (!ax36x) & (!ax35x) & (!shiftx0x) & (!shiftx1x)) + ((ax38x) & (ax37x) & (!ax36x) & (!ax35x) & (shiftx0x) & (!shiftx1x)) + ((ax38x) & (ax37x) & (!ax36x) & (ax35x) & (!shiftx0x) & (!shiftx1x)) + ((ax38x) & (ax37x) & (!ax36x) & (ax35x) & (shiftx0x) & (!shiftx1x)) + ((ax38x) & (ax37x) & (!ax36x) & (ax35x) & (shiftx0x) & (shiftx1x)) + ((ax38x) & (ax37x) & (ax36x) & (!ax35x) & (!shiftx0x) & (!shiftx1x)) + ((ax38x) & (ax37x) & (ax36x) & (!ax35x) & (!shiftx0x) & (shiftx1x)) + ((ax38x) & (ax37x) & (ax36x) & (!ax35x) & (shiftx0x) & (!shiftx1x)) + ((ax38x) & (ax37x) & (ax36x) & (ax35x) & (!shiftx0x) & (!shiftx1x)) + ((ax38x) & (ax37x) & (ax36x) & (ax35x) & (!shiftx0x) & (shiftx1x)) + ((ax38x) & (ax37x) & (ax36x) & (ax35x) & (shiftx0x) & (!shiftx1x)) + ((ax38x) & (ax37x) & (ax36x) & (ax35x) & (shiftx0x) & (shiftx1x)));
	assign g100 = (((!ax42x) & (!ax41x) & (!ax40x) & (ax39x) & (shiftx0x) & (shiftx1x)) + ((!ax42x) & (!ax41x) & (ax40x) & (!ax39x) & (!shiftx0x) & (shiftx1x)) + ((!ax42x) & (!ax41x) & (ax40x) & (ax39x) & (!shiftx0x) & (shiftx1x)) + ((!ax42x) & (!ax41x) & (ax40x) & (ax39x) & (shiftx0x) & (shiftx1x)) + ((!ax42x) & (ax41x) & (!ax40x) & (!ax39x) & (shiftx0x) & (!shiftx1x)) + ((!ax42x) & (ax41x) & (!ax40x) & (ax39x) & (shiftx0x) & (!shiftx1x)) + ((!ax42x) & (ax41x) & (!ax40x) & (ax39x) & (shiftx0x) & (shiftx1x)) + ((!ax42x) & (ax41x) & (ax40x) & (!ax39x) & (!shiftx0x) & (shiftx1x)) + ((!ax42x) & (ax41x) & (ax40x) & (!ax39x) & (shiftx0x) & (!shiftx1x)) + ((!ax42x) & (ax41x) & (ax40x) & (ax39x) & (!shiftx0x) & (shiftx1x)) + ((!ax42x) & (ax41x) & (ax40x) & (ax39x) & (shiftx0x) & (!shiftx1x)) + ((!ax42x) & (ax41x) & (ax40x) & (ax39x) & (shiftx0x) & (shiftx1x)) + ((ax42x) & (!ax41x) & (!ax40x) & (!ax39x) & (!shiftx0x) & (!shiftx1x)) + ((ax42x) & (!ax41x) & (!ax40x) & (ax39x) & (!shiftx0x) & (!shiftx1x)) + ((ax42x) & (!ax41x) & (!ax40x) & (ax39x) & (shiftx0x) & (shiftx1x)) + ((ax42x) & (!ax41x) & (ax40x) & (!ax39x) & (!shiftx0x) & (!shiftx1x)) + ((ax42x) & (!ax41x) & (ax40x) & (!ax39x) & (!shiftx0x) & (shiftx1x)) + ((ax42x) & (!ax41x) & (ax40x) & (ax39x) & (!shiftx0x) & (!shiftx1x)) + ((ax42x) & (!ax41x) & (ax40x) & (ax39x) & (!shiftx0x) & (shiftx1x)) + ((ax42x) & (!ax41x) & (ax40x) & (ax39x) & (shiftx0x) & (shiftx1x)) + ((ax42x) & (ax41x) & (!ax40x) & (!ax39x) & (!shiftx0x) & (!shiftx1x)) + ((ax42x) & (ax41x) & (!ax40x) & (!ax39x) & (shiftx0x) & (!shiftx1x)) + ((ax42x) & (ax41x) & (!ax40x) & (ax39x) & (!shiftx0x) & (!shiftx1x)) + ((ax42x) & (ax41x) & (!ax40x) & (ax39x) & (shiftx0x) & (!shiftx1x)) + ((ax42x) & (ax41x) & (!ax40x) & (ax39x) & (shiftx0x) & (shiftx1x)) + ((ax42x) & (ax41x) & (ax40x) & (!ax39x) & (!shiftx0x) & (!shiftx1x)) + ((ax42x) & (ax41x) & (ax40x) & (!ax39x) & (!shiftx0x) & (shiftx1x)) + ((ax42x) & (ax41x) & (ax40x) & (!ax39x) & (shiftx0x) & (!shiftx1x)) + ((ax42x) & (ax41x) & (ax40x) & (ax39x) & (!shiftx0x) & (!shiftx1x)) + ((ax42x) & (ax41x) & (ax40x) & (ax39x) & (!shiftx0x) & (shiftx1x)) + ((ax42x) & (ax41x) & (ax40x) & (ax39x) & (shiftx0x) & (!shiftx1x)) + ((ax42x) & (ax41x) & (ax40x) & (ax39x) & (shiftx0x) & (shiftx1x)));
	assign g101 = (((!shiftx2x) & (!shiftx3x) & (g97) & (!g98) & (!g99) & (!g100)) + ((!shiftx2x) & (!shiftx3x) & (g97) & (!g98) & (!g99) & (g100)) + ((!shiftx2x) & (!shiftx3x) & (g97) & (!g98) & (g99) & (!g100)) + ((!shiftx2x) & (!shiftx3x) & (g97) & (!g98) & (g99) & (g100)) + ((!shiftx2x) & (!shiftx3x) & (g97) & (g98) & (!g99) & (!g100)) + ((!shiftx2x) & (!shiftx3x) & (g97) & (g98) & (!g99) & (g100)) + ((!shiftx2x) & (!shiftx3x) & (g97) & (g98) & (g99) & (!g100)) + ((!shiftx2x) & (!shiftx3x) & (g97) & (g98) & (g99) & (g100)) + ((!shiftx2x) & (shiftx3x) & (!g97) & (!g98) & (!g99) & (g100)) + ((!shiftx2x) & (shiftx3x) & (!g97) & (!g98) & (g99) & (g100)) + ((!shiftx2x) & (shiftx3x) & (!g97) & (g98) & (!g99) & (g100)) + ((!shiftx2x) & (shiftx3x) & (!g97) & (g98) & (g99) & (g100)) + ((!shiftx2x) & (shiftx3x) & (g97) & (!g98) & (!g99) & (g100)) + ((!shiftx2x) & (shiftx3x) & (g97) & (!g98) & (g99) & (g100)) + ((!shiftx2x) & (shiftx3x) & (g97) & (g98) & (!g99) & (g100)) + ((!shiftx2x) & (shiftx3x) & (g97) & (g98) & (g99) & (g100)) + ((shiftx2x) & (!shiftx3x) & (!g97) & (g98) & (!g99) & (!g100)) + ((shiftx2x) & (!shiftx3x) & (!g97) & (g98) & (!g99) & (g100)) + ((shiftx2x) & (!shiftx3x) & (!g97) & (g98) & (g99) & (!g100)) + ((shiftx2x) & (!shiftx3x) & (!g97) & (g98) & (g99) & (g100)) + ((shiftx2x) & (!shiftx3x) & (g97) & (g98) & (!g99) & (!g100)) + ((shiftx2x) & (!shiftx3x) & (g97) & (g98) & (!g99) & (g100)) + ((shiftx2x) & (!shiftx3x) & (g97) & (g98) & (g99) & (!g100)) + ((shiftx2x) & (!shiftx3x) & (g97) & (g98) & (g99) & (g100)) + ((shiftx2x) & (shiftx3x) & (!g97) & (!g98) & (g99) & (!g100)) + ((shiftx2x) & (shiftx3x) & (!g97) & (!g98) & (g99) & (g100)) + ((shiftx2x) & (shiftx3x) & (!g97) & (g98) & (g99) & (!g100)) + ((shiftx2x) & (shiftx3x) & (!g97) & (g98) & (g99) & (g100)) + ((shiftx2x) & (shiftx3x) & (g97) & (!g98) & (g99) & (!g100)) + ((shiftx2x) & (shiftx3x) & (g97) & (!g98) & (g99) & (g100)) + ((shiftx2x) & (shiftx3x) & (g97) & (g98) & (g99) & (!g100)) + ((shiftx2x) & (shiftx3x) & (g97) & (g98) & (g99) & (g100)));
	assign g102 = (((!ax34x) & (!ax33x) & (!ax32x) & (ax31x) & (shiftx0x) & (shiftx1x)) + ((!ax34x) & (!ax33x) & (ax32x) & (!ax31x) & (!shiftx0x) & (shiftx1x)) + ((!ax34x) & (!ax33x) & (ax32x) & (ax31x) & (!shiftx0x) & (shiftx1x)) + ((!ax34x) & (!ax33x) & (ax32x) & (ax31x) & (shiftx0x) & (shiftx1x)) + ((!ax34x) & (ax33x) & (!ax32x) & (!ax31x) & (shiftx0x) & (!shiftx1x)) + ((!ax34x) & (ax33x) & (!ax32x) & (ax31x) & (shiftx0x) & (!shiftx1x)) + ((!ax34x) & (ax33x) & (!ax32x) & (ax31x) & (shiftx0x) & (shiftx1x)) + ((!ax34x) & (ax33x) & (ax32x) & (!ax31x) & (!shiftx0x) & (shiftx1x)) + ((!ax34x) & (ax33x) & (ax32x) & (!ax31x) & (shiftx0x) & (!shiftx1x)) + ((!ax34x) & (ax33x) & (ax32x) & (ax31x) & (!shiftx0x) & (shiftx1x)) + ((!ax34x) & (ax33x) & (ax32x) & (ax31x) & (shiftx0x) & (!shiftx1x)) + ((!ax34x) & (ax33x) & (ax32x) & (ax31x) & (shiftx0x) & (shiftx1x)) + ((ax34x) & (!ax33x) & (!ax32x) & (!ax31x) & (!shiftx0x) & (!shiftx1x)) + ((ax34x) & (!ax33x) & (!ax32x) & (ax31x) & (!shiftx0x) & (!shiftx1x)) + ((ax34x) & (!ax33x) & (!ax32x) & (ax31x) & (shiftx0x) & (shiftx1x)) + ((ax34x) & (!ax33x) & (ax32x) & (!ax31x) & (!shiftx0x) & (!shiftx1x)) + ((ax34x) & (!ax33x) & (ax32x) & (!ax31x) & (!shiftx0x) & (shiftx1x)) + ((ax34x) & (!ax33x) & (ax32x) & (ax31x) & (!shiftx0x) & (!shiftx1x)) + ((ax34x) & (!ax33x) & (ax32x) & (ax31x) & (!shiftx0x) & (shiftx1x)) + ((ax34x) & (!ax33x) & (ax32x) & (ax31x) & (shiftx0x) & (shiftx1x)) + ((ax34x) & (ax33x) & (!ax32x) & (!ax31x) & (!shiftx0x) & (!shiftx1x)) + ((ax34x) & (ax33x) & (!ax32x) & (!ax31x) & (shiftx0x) & (!shiftx1x)) + ((ax34x) & (ax33x) & (!ax32x) & (ax31x) & (!shiftx0x) & (!shiftx1x)) + ((ax34x) & (ax33x) & (!ax32x) & (ax31x) & (shiftx0x) & (!shiftx1x)) + ((ax34x) & (ax33x) & (!ax32x) & (ax31x) & (shiftx0x) & (shiftx1x)) + ((ax34x) & (ax33x) & (ax32x) & (!ax31x) & (!shiftx0x) & (!shiftx1x)) + ((ax34x) & (ax33x) & (ax32x) & (!ax31x) & (!shiftx0x) & (shiftx1x)) + ((ax34x) & (ax33x) & (ax32x) & (!ax31x) & (shiftx0x) & (!shiftx1x)) + ((ax34x) & (ax33x) & (ax32x) & (ax31x) & (!shiftx0x) & (!shiftx1x)) + ((ax34x) & (ax33x) & (ax32x) & (ax31x) & (!shiftx0x) & (shiftx1x)) + ((ax34x) & (ax33x) & (ax32x) & (ax31x) & (shiftx0x) & (!shiftx1x)) + ((ax34x) & (ax33x) & (ax32x) & (ax31x) & (shiftx0x) & (shiftx1x)));
	assign g103 = (((!ax30x) & (!ax29x) & (!ax28x) & (ax27x) & (shiftx0x) & (shiftx1x)) + ((!ax30x) & (!ax29x) & (ax28x) & (!ax27x) & (!shiftx0x) & (shiftx1x)) + ((!ax30x) & (!ax29x) & (ax28x) & (ax27x) & (!shiftx0x) & (shiftx1x)) + ((!ax30x) & (!ax29x) & (ax28x) & (ax27x) & (shiftx0x) & (shiftx1x)) + ((!ax30x) & (ax29x) & (!ax28x) & (!ax27x) & (shiftx0x) & (!shiftx1x)) + ((!ax30x) & (ax29x) & (!ax28x) & (ax27x) & (shiftx0x) & (!shiftx1x)) + ((!ax30x) & (ax29x) & (!ax28x) & (ax27x) & (shiftx0x) & (shiftx1x)) + ((!ax30x) & (ax29x) & (ax28x) & (!ax27x) & (!shiftx0x) & (shiftx1x)) + ((!ax30x) & (ax29x) & (ax28x) & (!ax27x) & (shiftx0x) & (!shiftx1x)) + ((!ax30x) & (ax29x) & (ax28x) & (ax27x) & (!shiftx0x) & (shiftx1x)) + ((!ax30x) & (ax29x) & (ax28x) & (ax27x) & (shiftx0x) & (!shiftx1x)) + ((!ax30x) & (ax29x) & (ax28x) & (ax27x) & (shiftx0x) & (shiftx1x)) + ((ax30x) & (!ax29x) & (!ax28x) & (!ax27x) & (!shiftx0x) & (!shiftx1x)) + ((ax30x) & (!ax29x) & (!ax28x) & (ax27x) & (!shiftx0x) & (!shiftx1x)) + ((ax30x) & (!ax29x) & (!ax28x) & (ax27x) & (shiftx0x) & (shiftx1x)) + ((ax30x) & (!ax29x) & (ax28x) & (!ax27x) & (!shiftx0x) & (!shiftx1x)) + ((ax30x) & (!ax29x) & (ax28x) & (!ax27x) & (!shiftx0x) & (shiftx1x)) + ((ax30x) & (!ax29x) & (ax28x) & (ax27x) & (!shiftx0x) & (!shiftx1x)) + ((ax30x) & (!ax29x) & (ax28x) & (ax27x) & (!shiftx0x) & (shiftx1x)) + ((ax30x) & (!ax29x) & (ax28x) & (ax27x) & (shiftx0x) & (shiftx1x)) + ((ax30x) & (ax29x) & (!ax28x) & (!ax27x) & (!shiftx0x) & (!shiftx1x)) + ((ax30x) & (ax29x) & (!ax28x) & (!ax27x) & (shiftx0x) & (!shiftx1x)) + ((ax30x) & (ax29x) & (!ax28x) & (ax27x) & (!shiftx0x) & (!shiftx1x)) + ((ax30x) & (ax29x) & (!ax28x) & (ax27x) & (shiftx0x) & (!shiftx1x)) + ((ax30x) & (ax29x) & (!ax28x) & (ax27x) & (shiftx0x) & (shiftx1x)) + ((ax30x) & (ax29x) & (ax28x) & (!ax27x) & (!shiftx0x) & (!shiftx1x)) + ((ax30x) & (ax29x) & (ax28x) & (!ax27x) & (!shiftx0x) & (shiftx1x)) + ((ax30x) & (ax29x) & (ax28x) & (!ax27x) & (shiftx0x) & (!shiftx1x)) + ((ax30x) & (ax29x) & (ax28x) & (ax27x) & (!shiftx0x) & (!shiftx1x)) + ((ax30x) & (ax29x) & (ax28x) & (ax27x) & (!shiftx0x) & (shiftx1x)) + ((ax30x) & (ax29x) & (ax28x) & (ax27x) & (shiftx0x) & (!shiftx1x)) + ((ax30x) & (ax29x) & (ax28x) & (ax27x) & (shiftx0x) & (shiftx1x)));
	assign g104 = (((!ax22x) & (!ax21x) & (!ax20x) & (ax19x) & (shiftx0x) & (shiftx1x)) + ((!ax22x) & (!ax21x) & (ax20x) & (!ax19x) & (!shiftx0x) & (shiftx1x)) + ((!ax22x) & (!ax21x) & (ax20x) & (ax19x) & (!shiftx0x) & (shiftx1x)) + ((!ax22x) & (!ax21x) & (ax20x) & (ax19x) & (shiftx0x) & (shiftx1x)) + ((!ax22x) & (ax21x) & (!ax20x) & (!ax19x) & (shiftx0x) & (!shiftx1x)) + ((!ax22x) & (ax21x) & (!ax20x) & (ax19x) & (shiftx0x) & (!shiftx1x)) + ((!ax22x) & (ax21x) & (!ax20x) & (ax19x) & (shiftx0x) & (shiftx1x)) + ((!ax22x) & (ax21x) & (ax20x) & (!ax19x) & (!shiftx0x) & (shiftx1x)) + ((!ax22x) & (ax21x) & (ax20x) & (!ax19x) & (shiftx0x) & (!shiftx1x)) + ((!ax22x) & (ax21x) & (ax20x) & (ax19x) & (!shiftx0x) & (shiftx1x)) + ((!ax22x) & (ax21x) & (ax20x) & (ax19x) & (shiftx0x) & (!shiftx1x)) + ((!ax22x) & (ax21x) & (ax20x) & (ax19x) & (shiftx0x) & (shiftx1x)) + ((ax22x) & (!ax21x) & (!ax20x) & (!ax19x) & (!shiftx0x) & (!shiftx1x)) + ((ax22x) & (!ax21x) & (!ax20x) & (ax19x) & (!shiftx0x) & (!shiftx1x)) + ((ax22x) & (!ax21x) & (!ax20x) & (ax19x) & (shiftx0x) & (shiftx1x)) + ((ax22x) & (!ax21x) & (ax20x) & (!ax19x) & (!shiftx0x) & (!shiftx1x)) + ((ax22x) & (!ax21x) & (ax20x) & (!ax19x) & (!shiftx0x) & (shiftx1x)) + ((ax22x) & (!ax21x) & (ax20x) & (ax19x) & (!shiftx0x) & (!shiftx1x)) + ((ax22x) & (!ax21x) & (ax20x) & (ax19x) & (!shiftx0x) & (shiftx1x)) + ((ax22x) & (!ax21x) & (ax20x) & (ax19x) & (shiftx0x) & (shiftx1x)) + ((ax22x) & (ax21x) & (!ax20x) & (!ax19x) & (!shiftx0x) & (!shiftx1x)) + ((ax22x) & (ax21x) & (!ax20x) & (!ax19x) & (shiftx0x) & (!shiftx1x)) + ((ax22x) & (ax21x) & (!ax20x) & (ax19x) & (!shiftx0x) & (!shiftx1x)) + ((ax22x) & (ax21x) & (!ax20x) & (ax19x) & (shiftx0x) & (!shiftx1x)) + ((ax22x) & (ax21x) & (!ax20x) & (ax19x) & (shiftx0x) & (shiftx1x)) + ((ax22x) & (ax21x) & (ax20x) & (!ax19x) & (!shiftx0x) & (!shiftx1x)) + ((ax22x) & (ax21x) & (ax20x) & (!ax19x) & (!shiftx0x) & (shiftx1x)) + ((ax22x) & (ax21x) & (ax20x) & (!ax19x) & (shiftx0x) & (!shiftx1x)) + ((ax22x) & (ax21x) & (ax20x) & (ax19x) & (!shiftx0x) & (!shiftx1x)) + ((ax22x) & (ax21x) & (ax20x) & (ax19x) & (!shiftx0x) & (shiftx1x)) + ((ax22x) & (ax21x) & (ax20x) & (ax19x) & (shiftx0x) & (!shiftx1x)) + ((ax22x) & (ax21x) & (ax20x) & (ax19x) & (shiftx0x) & (shiftx1x)));
	assign g105 = (((!ax26x) & (!ax25x) & (!ax24x) & (ax23x) & (shiftx0x) & (shiftx1x)) + ((!ax26x) & (!ax25x) & (ax24x) & (!ax23x) & (!shiftx0x) & (shiftx1x)) + ((!ax26x) & (!ax25x) & (ax24x) & (ax23x) & (!shiftx0x) & (shiftx1x)) + ((!ax26x) & (!ax25x) & (ax24x) & (ax23x) & (shiftx0x) & (shiftx1x)) + ((!ax26x) & (ax25x) & (!ax24x) & (!ax23x) & (shiftx0x) & (!shiftx1x)) + ((!ax26x) & (ax25x) & (!ax24x) & (ax23x) & (shiftx0x) & (!shiftx1x)) + ((!ax26x) & (ax25x) & (!ax24x) & (ax23x) & (shiftx0x) & (shiftx1x)) + ((!ax26x) & (ax25x) & (ax24x) & (!ax23x) & (!shiftx0x) & (shiftx1x)) + ((!ax26x) & (ax25x) & (ax24x) & (!ax23x) & (shiftx0x) & (!shiftx1x)) + ((!ax26x) & (ax25x) & (ax24x) & (ax23x) & (!shiftx0x) & (shiftx1x)) + ((!ax26x) & (ax25x) & (ax24x) & (ax23x) & (shiftx0x) & (!shiftx1x)) + ((!ax26x) & (ax25x) & (ax24x) & (ax23x) & (shiftx0x) & (shiftx1x)) + ((ax26x) & (!ax25x) & (!ax24x) & (!ax23x) & (!shiftx0x) & (!shiftx1x)) + ((ax26x) & (!ax25x) & (!ax24x) & (ax23x) & (!shiftx0x) & (!shiftx1x)) + ((ax26x) & (!ax25x) & (!ax24x) & (ax23x) & (shiftx0x) & (shiftx1x)) + ((ax26x) & (!ax25x) & (ax24x) & (!ax23x) & (!shiftx0x) & (!shiftx1x)) + ((ax26x) & (!ax25x) & (ax24x) & (!ax23x) & (!shiftx0x) & (shiftx1x)) + ((ax26x) & (!ax25x) & (ax24x) & (ax23x) & (!shiftx0x) & (!shiftx1x)) + ((ax26x) & (!ax25x) & (ax24x) & (ax23x) & (!shiftx0x) & (shiftx1x)) + ((ax26x) & (!ax25x) & (ax24x) & (ax23x) & (shiftx0x) & (shiftx1x)) + ((ax26x) & (ax25x) & (!ax24x) & (!ax23x) & (!shiftx0x) & (!shiftx1x)) + ((ax26x) & (ax25x) & (!ax24x) & (!ax23x) & (shiftx0x) & (!shiftx1x)) + ((ax26x) & (ax25x) & (!ax24x) & (ax23x) & (!shiftx0x) & (!shiftx1x)) + ((ax26x) & (ax25x) & (!ax24x) & (ax23x) & (shiftx0x) & (!shiftx1x)) + ((ax26x) & (ax25x) & (!ax24x) & (ax23x) & (shiftx0x) & (shiftx1x)) + ((ax26x) & (ax25x) & (ax24x) & (!ax23x) & (!shiftx0x) & (!shiftx1x)) + ((ax26x) & (ax25x) & (ax24x) & (!ax23x) & (!shiftx0x) & (shiftx1x)) + ((ax26x) & (ax25x) & (ax24x) & (!ax23x) & (shiftx0x) & (!shiftx1x)) + ((ax26x) & (ax25x) & (ax24x) & (ax23x) & (!shiftx0x) & (!shiftx1x)) + ((ax26x) & (ax25x) & (ax24x) & (ax23x) & (!shiftx0x) & (shiftx1x)) + ((ax26x) & (ax25x) & (ax24x) & (ax23x) & (shiftx0x) & (!shiftx1x)) + ((ax26x) & (ax25x) & (ax24x) & (ax23x) & (shiftx0x) & (shiftx1x)));
	assign g106 = (((!shiftx2x) & (!shiftx3x) & (g102) & (!g103) & (!g104) & (!g105)) + ((!shiftx2x) & (!shiftx3x) & (g102) & (!g103) & (!g104) & (g105)) + ((!shiftx2x) & (!shiftx3x) & (g102) & (!g103) & (g104) & (!g105)) + ((!shiftx2x) & (!shiftx3x) & (g102) & (!g103) & (g104) & (g105)) + ((!shiftx2x) & (!shiftx3x) & (g102) & (g103) & (!g104) & (!g105)) + ((!shiftx2x) & (!shiftx3x) & (g102) & (g103) & (!g104) & (g105)) + ((!shiftx2x) & (!shiftx3x) & (g102) & (g103) & (g104) & (!g105)) + ((!shiftx2x) & (!shiftx3x) & (g102) & (g103) & (g104) & (g105)) + ((!shiftx2x) & (shiftx3x) & (!g102) & (!g103) & (!g104) & (g105)) + ((!shiftx2x) & (shiftx3x) & (!g102) & (!g103) & (g104) & (g105)) + ((!shiftx2x) & (shiftx3x) & (!g102) & (g103) & (!g104) & (g105)) + ((!shiftx2x) & (shiftx3x) & (!g102) & (g103) & (g104) & (g105)) + ((!shiftx2x) & (shiftx3x) & (g102) & (!g103) & (!g104) & (g105)) + ((!shiftx2x) & (shiftx3x) & (g102) & (!g103) & (g104) & (g105)) + ((!shiftx2x) & (shiftx3x) & (g102) & (g103) & (!g104) & (g105)) + ((!shiftx2x) & (shiftx3x) & (g102) & (g103) & (g104) & (g105)) + ((shiftx2x) & (!shiftx3x) & (!g102) & (g103) & (!g104) & (!g105)) + ((shiftx2x) & (!shiftx3x) & (!g102) & (g103) & (!g104) & (g105)) + ((shiftx2x) & (!shiftx3x) & (!g102) & (g103) & (g104) & (!g105)) + ((shiftx2x) & (!shiftx3x) & (!g102) & (g103) & (g104) & (g105)) + ((shiftx2x) & (!shiftx3x) & (g102) & (g103) & (!g104) & (!g105)) + ((shiftx2x) & (!shiftx3x) & (g102) & (g103) & (!g104) & (g105)) + ((shiftx2x) & (!shiftx3x) & (g102) & (g103) & (g104) & (!g105)) + ((shiftx2x) & (!shiftx3x) & (g102) & (g103) & (g104) & (g105)) + ((shiftx2x) & (shiftx3x) & (!g102) & (!g103) & (g104) & (!g105)) + ((shiftx2x) & (shiftx3x) & (!g102) & (!g103) & (g104) & (g105)) + ((shiftx2x) & (shiftx3x) & (!g102) & (g103) & (g104) & (!g105)) + ((shiftx2x) & (shiftx3x) & (!g102) & (g103) & (g104) & (g105)) + ((shiftx2x) & (shiftx3x) & (g102) & (!g103) & (g104) & (!g105)) + ((shiftx2x) & (shiftx3x) & (g102) & (!g103) & (g104) & (g105)) + ((shiftx2x) & (shiftx3x) & (g102) & (g103) & (g104) & (!g105)) + ((shiftx2x) & (shiftx3x) & (g102) & (g103) & (g104) & (g105)));
	assign g107 = (((!shiftx4x) & (!shiftx5x) & (g91) & (!g96) & (!g101) & (!g106)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (!g96) & (!g101) & (g106)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (!g96) & (g101) & (!g106)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (!g96) & (g101) & (g106)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (g96) & (!g101) & (!g106)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (g96) & (!g101) & (g106)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (g96) & (g101) & (!g106)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (g96) & (g101) & (g106)) + ((!shiftx4x) & (shiftx5x) & (!g91) & (!g96) & (!g101) & (g106)) + ((!shiftx4x) & (shiftx5x) & (!g91) & (!g96) & (g101) & (g106)) + ((!shiftx4x) & (shiftx5x) & (!g91) & (g96) & (!g101) & (g106)) + ((!shiftx4x) & (shiftx5x) & (!g91) & (g96) & (g101) & (g106)) + ((!shiftx4x) & (shiftx5x) & (g91) & (!g96) & (!g101) & (g106)) + ((!shiftx4x) & (shiftx5x) & (g91) & (!g96) & (g101) & (g106)) + ((!shiftx4x) & (shiftx5x) & (g91) & (g96) & (!g101) & (g106)) + ((!shiftx4x) & (shiftx5x) & (g91) & (g96) & (g101) & (g106)) + ((shiftx4x) & (!shiftx5x) & (!g91) & (!g96) & (g101) & (!g106)) + ((shiftx4x) & (!shiftx5x) & (!g91) & (!g96) & (g101) & (g106)) + ((shiftx4x) & (!shiftx5x) & (!g91) & (g96) & (g101) & (!g106)) + ((shiftx4x) & (!shiftx5x) & (!g91) & (g96) & (g101) & (g106)) + ((shiftx4x) & (!shiftx5x) & (g91) & (!g96) & (g101) & (!g106)) + ((shiftx4x) & (!shiftx5x) & (g91) & (!g96) & (g101) & (g106)) + ((shiftx4x) & (!shiftx5x) & (g91) & (g96) & (g101) & (!g106)) + ((shiftx4x) & (!shiftx5x) & (g91) & (g96) & (g101) & (g106)) + ((shiftx4x) & (shiftx5x) & (!g91) & (g96) & (!g101) & (!g106)) + ((shiftx4x) & (shiftx5x) & (!g91) & (g96) & (!g101) & (g106)) + ((shiftx4x) & (shiftx5x) & (!g91) & (g96) & (g101) & (!g106)) + ((shiftx4x) & (shiftx5x) & (!g91) & (g96) & (g101) & (g106)) + ((shiftx4x) & (shiftx5x) & (g91) & (g96) & (!g101) & (!g106)) + ((shiftx4x) & (shiftx5x) & (g91) & (g96) & (!g101) & (g106)) + ((shiftx4x) & (shiftx5x) & (g91) & (g96) & (g101) & (!g106)) + ((shiftx4x) & (shiftx5x) & (g91) & (g96) & (g101) & (g106)));
	assign g108 = (((!ax82x) & (!ax81x) & (!ax80x) & (ax79x) & (shiftx0x) & (shiftx1x)) + ((!ax82x) & (!ax81x) & (ax80x) & (!ax79x) & (!shiftx0x) & (shiftx1x)) + ((!ax82x) & (!ax81x) & (ax80x) & (ax79x) & (!shiftx0x) & (shiftx1x)) + ((!ax82x) & (!ax81x) & (ax80x) & (ax79x) & (shiftx0x) & (shiftx1x)) + ((!ax82x) & (ax81x) & (!ax80x) & (!ax79x) & (shiftx0x) & (!shiftx1x)) + ((!ax82x) & (ax81x) & (!ax80x) & (ax79x) & (shiftx0x) & (!shiftx1x)) + ((!ax82x) & (ax81x) & (!ax80x) & (ax79x) & (shiftx0x) & (shiftx1x)) + ((!ax82x) & (ax81x) & (ax80x) & (!ax79x) & (!shiftx0x) & (shiftx1x)) + ((!ax82x) & (ax81x) & (ax80x) & (!ax79x) & (shiftx0x) & (!shiftx1x)) + ((!ax82x) & (ax81x) & (ax80x) & (ax79x) & (!shiftx0x) & (shiftx1x)) + ((!ax82x) & (ax81x) & (ax80x) & (ax79x) & (shiftx0x) & (!shiftx1x)) + ((!ax82x) & (ax81x) & (ax80x) & (ax79x) & (shiftx0x) & (shiftx1x)) + ((ax82x) & (!ax81x) & (!ax80x) & (!ax79x) & (!shiftx0x) & (!shiftx1x)) + ((ax82x) & (!ax81x) & (!ax80x) & (ax79x) & (!shiftx0x) & (!shiftx1x)) + ((ax82x) & (!ax81x) & (!ax80x) & (ax79x) & (shiftx0x) & (shiftx1x)) + ((ax82x) & (!ax81x) & (ax80x) & (!ax79x) & (!shiftx0x) & (!shiftx1x)) + ((ax82x) & (!ax81x) & (ax80x) & (!ax79x) & (!shiftx0x) & (shiftx1x)) + ((ax82x) & (!ax81x) & (ax80x) & (ax79x) & (!shiftx0x) & (!shiftx1x)) + ((ax82x) & (!ax81x) & (ax80x) & (ax79x) & (!shiftx0x) & (shiftx1x)) + ((ax82x) & (!ax81x) & (ax80x) & (ax79x) & (shiftx0x) & (shiftx1x)) + ((ax82x) & (ax81x) & (!ax80x) & (!ax79x) & (!shiftx0x) & (!shiftx1x)) + ((ax82x) & (ax81x) & (!ax80x) & (!ax79x) & (shiftx0x) & (!shiftx1x)) + ((ax82x) & (ax81x) & (!ax80x) & (ax79x) & (!shiftx0x) & (!shiftx1x)) + ((ax82x) & (ax81x) & (!ax80x) & (ax79x) & (shiftx0x) & (!shiftx1x)) + ((ax82x) & (ax81x) & (!ax80x) & (ax79x) & (shiftx0x) & (shiftx1x)) + ((ax82x) & (ax81x) & (ax80x) & (!ax79x) & (!shiftx0x) & (!shiftx1x)) + ((ax82x) & (ax81x) & (ax80x) & (!ax79x) & (!shiftx0x) & (shiftx1x)) + ((ax82x) & (ax81x) & (ax80x) & (!ax79x) & (shiftx0x) & (!shiftx1x)) + ((ax82x) & (ax81x) & (ax80x) & (ax79x) & (!shiftx0x) & (!shiftx1x)) + ((ax82x) & (ax81x) & (ax80x) & (ax79x) & (!shiftx0x) & (shiftx1x)) + ((ax82x) & (ax81x) & (ax80x) & (ax79x) & (shiftx0x) & (!shiftx1x)) + ((ax82x) & (ax81x) & (ax80x) & (ax79x) & (shiftx0x) & (shiftx1x)));
	assign g109 = (((!ax78x) & (!ax77x) & (!ax76x) & (ax75x) & (shiftx0x) & (shiftx1x)) + ((!ax78x) & (!ax77x) & (ax76x) & (!ax75x) & (!shiftx0x) & (shiftx1x)) + ((!ax78x) & (!ax77x) & (ax76x) & (ax75x) & (!shiftx0x) & (shiftx1x)) + ((!ax78x) & (!ax77x) & (ax76x) & (ax75x) & (shiftx0x) & (shiftx1x)) + ((!ax78x) & (ax77x) & (!ax76x) & (!ax75x) & (shiftx0x) & (!shiftx1x)) + ((!ax78x) & (ax77x) & (!ax76x) & (ax75x) & (shiftx0x) & (!shiftx1x)) + ((!ax78x) & (ax77x) & (!ax76x) & (ax75x) & (shiftx0x) & (shiftx1x)) + ((!ax78x) & (ax77x) & (ax76x) & (!ax75x) & (!shiftx0x) & (shiftx1x)) + ((!ax78x) & (ax77x) & (ax76x) & (!ax75x) & (shiftx0x) & (!shiftx1x)) + ((!ax78x) & (ax77x) & (ax76x) & (ax75x) & (!shiftx0x) & (shiftx1x)) + ((!ax78x) & (ax77x) & (ax76x) & (ax75x) & (shiftx0x) & (!shiftx1x)) + ((!ax78x) & (ax77x) & (ax76x) & (ax75x) & (shiftx0x) & (shiftx1x)) + ((ax78x) & (!ax77x) & (!ax76x) & (!ax75x) & (!shiftx0x) & (!shiftx1x)) + ((ax78x) & (!ax77x) & (!ax76x) & (ax75x) & (!shiftx0x) & (!shiftx1x)) + ((ax78x) & (!ax77x) & (!ax76x) & (ax75x) & (shiftx0x) & (shiftx1x)) + ((ax78x) & (!ax77x) & (ax76x) & (!ax75x) & (!shiftx0x) & (!shiftx1x)) + ((ax78x) & (!ax77x) & (ax76x) & (!ax75x) & (!shiftx0x) & (shiftx1x)) + ((ax78x) & (!ax77x) & (ax76x) & (ax75x) & (!shiftx0x) & (!shiftx1x)) + ((ax78x) & (!ax77x) & (ax76x) & (ax75x) & (!shiftx0x) & (shiftx1x)) + ((ax78x) & (!ax77x) & (ax76x) & (ax75x) & (shiftx0x) & (shiftx1x)) + ((ax78x) & (ax77x) & (!ax76x) & (!ax75x) & (!shiftx0x) & (!shiftx1x)) + ((ax78x) & (ax77x) & (!ax76x) & (!ax75x) & (shiftx0x) & (!shiftx1x)) + ((ax78x) & (ax77x) & (!ax76x) & (ax75x) & (!shiftx0x) & (!shiftx1x)) + ((ax78x) & (ax77x) & (!ax76x) & (ax75x) & (shiftx0x) & (!shiftx1x)) + ((ax78x) & (ax77x) & (!ax76x) & (ax75x) & (shiftx0x) & (shiftx1x)) + ((ax78x) & (ax77x) & (ax76x) & (!ax75x) & (!shiftx0x) & (!shiftx1x)) + ((ax78x) & (ax77x) & (ax76x) & (!ax75x) & (!shiftx0x) & (shiftx1x)) + ((ax78x) & (ax77x) & (ax76x) & (!ax75x) & (shiftx0x) & (!shiftx1x)) + ((ax78x) & (ax77x) & (ax76x) & (ax75x) & (!shiftx0x) & (!shiftx1x)) + ((ax78x) & (ax77x) & (ax76x) & (ax75x) & (!shiftx0x) & (shiftx1x)) + ((ax78x) & (ax77x) & (ax76x) & (ax75x) & (shiftx0x) & (!shiftx1x)) + ((ax78x) & (ax77x) & (ax76x) & (ax75x) & (shiftx0x) & (shiftx1x)));
	assign g110 = (((!ax70x) & (!ax69x) & (!ax68x) & (ax67x) & (shiftx0x) & (shiftx1x)) + ((!ax70x) & (!ax69x) & (ax68x) & (!ax67x) & (!shiftx0x) & (shiftx1x)) + ((!ax70x) & (!ax69x) & (ax68x) & (ax67x) & (!shiftx0x) & (shiftx1x)) + ((!ax70x) & (!ax69x) & (ax68x) & (ax67x) & (shiftx0x) & (shiftx1x)) + ((!ax70x) & (ax69x) & (!ax68x) & (!ax67x) & (shiftx0x) & (!shiftx1x)) + ((!ax70x) & (ax69x) & (!ax68x) & (ax67x) & (shiftx0x) & (!shiftx1x)) + ((!ax70x) & (ax69x) & (!ax68x) & (ax67x) & (shiftx0x) & (shiftx1x)) + ((!ax70x) & (ax69x) & (ax68x) & (!ax67x) & (!shiftx0x) & (shiftx1x)) + ((!ax70x) & (ax69x) & (ax68x) & (!ax67x) & (shiftx0x) & (!shiftx1x)) + ((!ax70x) & (ax69x) & (ax68x) & (ax67x) & (!shiftx0x) & (shiftx1x)) + ((!ax70x) & (ax69x) & (ax68x) & (ax67x) & (shiftx0x) & (!shiftx1x)) + ((!ax70x) & (ax69x) & (ax68x) & (ax67x) & (shiftx0x) & (shiftx1x)) + ((ax70x) & (!ax69x) & (!ax68x) & (!ax67x) & (!shiftx0x) & (!shiftx1x)) + ((ax70x) & (!ax69x) & (!ax68x) & (ax67x) & (!shiftx0x) & (!shiftx1x)) + ((ax70x) & (!ax69x) & (!ax68x) & (ax67x) & (shiftx0x) & (shiftx1x)) + ((ax70x) & (!ax69x) & (ax68x) & (!ax67x) & (!shiftx0x) & (!shiftx1x)) + ((ax70x) & (!ax69x) & (ax68x) & (!ax67x) & (!shiftx0x) & (shiftx1x)) + ((ax70x) & (!ax69x) & (ax68x) & (ax67x) & (!shiftx0x) & (!shiftx1x)) + ((ax70x) & (!ax69x) & (ax68x) & (ax67x) & (!shiftx0x) & (shiftx1x)) + ((ax70x) & (!ax69x) & (ax68x) & (ax67x) & (shiftx0x) & (shiftx1x)) + ((ax70x) & (ax69x) & (!ax68x) & (!ax67x) & (!shiftx0x) & (!shiftx1x)) + ((ax70x) & (ax69x) & (!ax68x) & (!ax67x) & (shiftx0x) & (!shiftx1x)) + ((ax70x) & (ax69x) & (!ax68x) & (ax67x) & (!shiftx0x) & (!shiftx1x)) + ((ax70x) & (ax69x) & (!ax68x) & (ax67x) & (shiftx0x) & (!shiftx1x)) + ((ax70x) & (ax69x) & (!ax68x) & (ax67x) & (shiftx0x) & (shiftx1x)) + ((ax70x) & (ax69x) & (ax68x) & (!ax67x) & (!shiftx0x) & (!shiftx1x)) + ((ax70x) & (ax69x) & (ax68x) & (!ax67x) & (!shiftx0x) & (shiftx1x)) + ((ax70x) & (ax69x) & (ax68x) & (!ax67x) & (shiftx0x) & (!shiftx1x)) + ((ax70x) & (ax69x) & (ax68x) & (ax67x) & (!shiftx0x) & (!shiftx1x)) + ((ax70x) & (ax69x) & (ax68x) & (ax67x) & (!shiftx0x) & (shiftx1x)) + ((ax70x) & (ax69x) & (ax68x) & (ax67x) & (shiftx0x) & (!shiftx1x)) + ((ax70x) & (ax69x) & (ax68x) & (ax67x) & (shiftx0x) & (shiftx1x)));
	assign g111 = (((!ax74x) & (!ax73x) & (!ax72x) & (ax71x) & (shiftx0x) & (shiftx1x)) + ((!ax74x) & (!ax73x) & (ax72x) & (!ax71x) & (!shiftx0x) & (shiftx1x)) + ((!ax74x) & (!ax73x) & (ax72x) & (ax71x) & (!shiftx0x) & (shiftx1x)) + ((!ax74x) & (!ax73x) & (ax72x) & (ax71x) & (shiftx0x) & (shiftx1x)) + ((!ax74x) & (ax73x) & (!ax72x) & (!ax71x) & (shiftx0x) & (!shiftx1x)) + ((!ax74x) & (ax73x) & (!ax72x) & (ax71x) & (shiftx0x) & (!shiftx1x)) + ((!ax74x) & (ax73x) & (!ax72x) & (ax71x) & (shiftx0x) & (shiftx1x)) + ((!ax74x) & (ax73x) & (ax72x) & (!ax71x) & (!shiftx0x) & (shiftx1x)) + ((!ax74x) & (ax73x) & (ax72x) & (!ax71x) & (shiftx0x) & (!shiftx1x)) + ((!ax74x) & (ax73x) & (ax72x) & (ax71x) & (!shiftx0x) & (shiftx1x)) + ((!ax74x) & (ax73x) & (ax72x) & (ax71x) & (shiftx0x) & (!shiftx1x)) + ((!ax74x) & (ax73x) & (ax72x) & (ax71x) & (shiftx0x) & (shiftx1x)) + ((ax74x) & (!ax73x) & (!ax72x) & (!ax71x) & (!shiftx0x) & (!shiftx1x)) + ((ax74x) & (!ax73x) & (!ax72x) & (ax71x) & (!shiftx0x) & (!shiftx1x)) + ((ax74x) & (!ax73x) & (!ax72x) & (ax71x) & (shiftx0x) & (shiftx1x)) + ((ax74x) & (!ax73x) & (ax72x) & (!ax71x) & (!shiftx0x) & (!shiftx1x)) + ((ax74x) & (!ax73x) & (ax72x) & (!ax71x) & (!shiftx0x) & (shiftx1x)) + ((ax74x) & (!ax73x) & (ax72x) & (ax71x) & (!shiftx0x) & (!shiftx1x)) + ((ax74x) & (!ax73x) & (ax72x) & (ax71x) & (!shiftx0x) & (shiftx1x)) + ((ax74x) & (!ax73x) & (ax72x) & (ax71x) & (shiftx0x) & (shiftx1x)) + ((ax74x) & (ax73x) & (!ax72x) & (!ax71x) & (!shiftx0x) & (!shiftx1x)) + ((ax74x) & (ax73x) & (!ax72x) & (!ax71x) & (shiftx0x) & (!shiftx1x)) + ((ax74x) & (ax73x) & (!ax72x) & (ax71x) & (!shiftx0x) & (!shiftx1x)) + ((ax74x) & (ax73x) & (!ax72x) & (ax71x) & (shiftx0x) & (!shiftx1x)) + ((ax74x) & (ax73x) & (!ax72x) & (ax71x) & (shiftx0x) & (shiftx1x)) + ((ax74x) & (ax73x) & (ax72x) & (!ax71x) & (!shiftx0x) & (!shiftx1x)) + ((ax74x) & (ax73x) & (ax72x) & (!ax71x) & (!shiftx0x) & (shiftx1x)) + ((ax74x) & (ax73x) & (ax72x) & (!ax71x) & (shiftx0x) & (!shiftx1x)) + ((ax74x) & (ax73x) & (ax72x) & (ax71x) & (!shiftx0x) & (!shiftx1x)) + ((ax74x) & (ax73x) & (ax72x) & (ax71x) & (!shiftx0x) & (shiftx1x)) + ((ax74x) & (ax73x) & (ax72x) & (ax71x) & (shiftx0x) & (!shiftx1x)) + ((ax74x) & (ax73x) & (ax72x) & (ax71x) & (shiftx0x) & (shiftx1x)));
	assign g112 = (((!shiftx2x) & (!shiftx3x) & (g108) & (!g109) & (!g110) & (!g111)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (!g109) & (!g110) & (g111)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (!g109) & (g110) & (!g111)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (!g109) & (g110) & (g111)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (g109) & (!g110) & (!g111)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (g109) & (!g110) & (g111)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (g109) & (g110) & (!g111)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (g109) & (g110) & (g111)) + ((!shiftx2x) & (shiftx3x) & (!g108) & (!g109) & (!g110) & (g111)) + ((!shiftx2x) & (shiftx3x) & (!g108) & (!g109) & (g110) & (g111)) + ((!shiftx2x) & (shiftx3x) & (!g108) & (g109) & (!g110) & (g111)) + ((!shiftx2x) & (shiftx3x) & (!g108) & (g109) & (g110) & (g111)) + ((!shiftx2x) & (shiftx3x) & (g108) & (!g109) & (!g110) & (g111)) + ((!shiftx2x) & (shiftx3x) & (g108) & (!g109) & (g110) & (g111)) + ((!shiftx2x) & (shiftx3x) & (g108) & (g109) & (!g110) & (g111)) + ((!shiftx2x) & (shiftx3x) & (g108) & (g109) & (g110) & (g111)) + ((shiftx2x) & (!shiftx3x) & (!g108) & (g109) & (!g110) & (!g111)) + ((shiftx2x) & (!shiftx3x) & (!g108) & (g109) & (!g110) & (g111)) + ((shiftx2x) & (!shiftx3x) & (!g108) & (g109) & (g110) & (!g111)) + ((shiftx2x) & (!shiftx3x) & (!g108) & (g109) & (g110) & (g111)) + ((shiftx2x) & (!shiftx3x) & (g108) & (g109) & (!g110) & (!g111)) + ((shiftx2x) & (!shiftx3x) & (g108) & (g109) & (!g110) & (g111)) + ((shiftx2x) & (!shiftx3x) & (g108) & (g109) & (g110) & (!g111)) + ((shiftx2x) & (!shiftx3x) & (g108) & (g109) & (g110) & (g111)) + ((shiftx2x) & (shiftx3x) & (!g108) & (!g109) & (g110) & (!g111)) + ((shiftx2x) & (shiftx3x) & (!g108) & (!g109) & (g110) & (g111)) + ((shiftx2x) & (shiftx3x) & (!g108) & (g109) & (g110) & (!g111)) + ((shiftx2x) & (shiftx3x) & (!g108) & (g109) & (g110) & (g111)) + ((shiftx2x) & (shiftx3x) & (g108) & (!g109) & (g110) & (!g111)) + ((shiftx2x) & (shiftx3x) & (g108) & (!g109) & (g110) & (g111)) + ((shiftx2x) & (shiftx3x) & (g108) & (g109) & (g110) & (!g111)) + ((shiftx2x) & (shiftx3x) & (g108) & (g109) & (g110) & (g111)));
	assign g113 = (((!ax98x) & (!ax97x) & (!ax96x) & (ax95x) & (shiftx0x) & (shiftx1x)) + ((!ax98x) & (!ax97x) & (ax96x) & (!ax95x) & (!shiftx0x) & (shiftx1x)) + ((!ax98x) & (!ax97x) & (ax96x) & (ax95x) & (!shiftx0x) & (shiftx1x)) + ((!ax98x) & (!ax97x) & (ax96x) & (ax95x) & (shiftx0x) & (shiftx1x)) + ((!ax98x) & (ax97x) & (!ax96x) & (!ax95x) & (shiftx0x) & (!shiftx1x)) + ((!ax98x) & (ax97x) & (!ax96x) & (ax95x) & (shiftx0x) & (!shiftx1x)) + ((!ax98x) & (ax97x) & (!ax96x) & (ax95x) & (shiftx0x) & (shiftx1x)) + ((!ax98x) & (ax97x) & (ax96x) & (!ax95x) & (!shiftx0x) & (shiftx1x)) + ((!ax98x) & (ax97x) & (ax96x) & (!ax95x) & (shiftx0x) & (!shiftx1x)) + ((!ax98x) & (ax97x) & (ax96x) & (ax95x) & (!shiftx0x) & (shiftx1x)) + ((!ax98x) & (ax97x) & (ax96x) & (ax95x) & (shiftx0x) & (!shiftx1x)) + ((!ax98x) & (ax97x) & (ax96x) & (ax95x) & (shiftx0x) & (shiftx1x)) + ((ax98x) & (!ax97x) & (!ax96x) & (!ax95x) & (!shiftx0x) & (!shiftx1x)) + ((ax98x) & (!ax97x) & (!ax96x) & (ax95x) & (!shiftx0x) & (!shiftx1x)) + ((ax98x) & (!ax97x) & (!ax96x) & (ax95x) & (shiftx0x) & (shiftx1x)) + ((ax98x) & (!ax97x) & (ax96x) & (!ax95x) & (!shiftx0x) & (!shiftx1x)) + ((ax98x) & (!ax97x) & (ax96x) & (!ax95x) & (!shiftx0x) & (shiftx1x)) + ((ax98x) & (!ax97x) & (ax96x) & (ax95x) & (!shiftx0x) & (!shiftx1x)) + ((ax98x) & (!ax97x) & (ax96x) & (ax95x) & (!shiftx0x) & (shiftx1x)) + ((ax98x) & (!ax97x) & (ax96x) & (ax95x) & (shiftx0x) & (shiftx1x)) + ((ax98x) & (ax97x) & (!ax96x) & (!ax95x) & (!shiftx0x) & (!shiftx1x)) + ((ax98x) & (ax97x) & (!ax96x) & (!ax95x) & (shiftx0x) & (!shiftx1x)) + ((ax98x) & (ax97x) & (!ax96x) & (ax95x) & (!shiftx0x) & (!shiftx1x)) + ((ax98x) & (ax97x) & (!ax96x) & (ax95x) & (shiftx0x) & (!shiftx1x)) + ((ax98x) & (ax97x) & (!ax96x) & (ax95x) & (shiftx0x) & (shiftx1x)) + ((ax98x) & (ax97x) & (ax96x) & (!ax95x) & (!shiftx0x) & (!shiftx1x)) + ((ax98x) & (ax97x) & (ax96x) & (!ax95x) & (!shiftx0x) & (shiftx1x)) + ((ax98x) & (ax97x) & (ax96x) & (!ax95x) & (shiftx0x) & (!shiftx1x)) + ((ax98x) & (ax97x) & (ax96x) & (ax95x) & (!shiftx0x) & (!shiftx1x)) + ((ax98x) & (ax97x) & (ax96x) & (ax95x) & (!shiftx0x) & (shiftx1x)) + ((ax98x) & (ax97x) & (ax96x) & (ax95x) & (shiftx0x) & (!shiftx1x)) + ((ax98x) & (ax97x) & (ax96x) & (ax95x) & (shiftx0x) & (shiftx1x)));
	assign g114 = (((!ax94x) & (!ax93x) & (!ax92x) & (ax91x) & (shiftx0x) & (shiftx1x)) + ((!ax94x) & (!ax93x) & (ax92x) & (!ax91x) & (!shiftx0x) & (shiftx1x)) + ((!ax94x) & (!ax93x) & (ax92x) & (ax91x) & (!shiftx0x) & (shiftx1x)) + ((!ax94x) & (!ax93x) & (ax92x) & (ax91x) & (shiftx0x) & (shiftx1x)) + ((!ax94x) & (ax93x) & (!ax92x) & (!ax91x) & (shiftx0x) & (!shiftx1x)) + ((!ax94x) & (ax93x) & (!ax92x) & (ax91x) & (shiftx0x) & (!shiftx1x)) + ((!ax94x) & (ax93x) & (!ax92x) & (ax91x) & (shiftx0x) & (shiftx1x)) + ((!ax94x) & (ax93x) & (ax92x) & (!ax91x) & (!shiftx0x) & (shiftx1x)) + ((!ax94x) & (ax93x) & (ax92x) & (!ax91x) & (shiftx0x) & (!shiftx1x)) + ((!ax94x) & (ax93x) & (ax92x) & (ax91x) & (!shiftx0x) & (shiftx1x)) + ((!ax94x) & (ax93x) & (ax92x) & (ax91x) & (shiftx0x) & (!shiftx1x)) + ((!ax94x) & (ax93x) & (ax92x) & (ax91x) & (shiftx0x) & (shiftx1x)) + ((ax94x) & (!ax93x) & (!ax92x) & (!ax91x) & (!shiftx0x) & (!shiftx1x)) + ((ax94x) & (!ax93x) & (!ax92x) & (ax91x) & (!shiftx0x) & (!shiftx1x)) + ((ax94x) & (!ax93x) & (!ax92x) & (ax91x) & (shiftx0x) & (shiftx1x)) + ((ax94x) & (!ax93x) & (ax92x) & (!ax91x) & (!shiftx0x) & (!shiftx1x)) + ((ax94x) & (!ax93x) & (ax92x) & (!ax91x) & (!shiftx0x) & (shiftx1x)) + ((ax94x) & (!ax93x) & (ax92x) & (ax91x) & (!shiftx0x) & (!shiftx1x)) + ((ax94x) & (!ax93x) & (ax92x) & (ax91x) & (!shiftx0x) & (shiftx1x)) + ((ax94x) & (!ax93x) & (ax92x) & (ax91x) & (shiftx0x) & (shiftx1x)) + ((ax94x) & (ax93x) & (!ax92x) & (!ax91x) & (!shiftx0x) & (!shiftx1x)) + ((ax94x) & (ax93x) & (!ax92x) & (!ax91x) & (shiftx0x) & (!shiftx1x)) + ((ax94x) & (ax93x) & (!ax92x) & (ax91x) & (!shiftx0x) & (!shiftx1x)) + ((ax94x) & (ax93x) & (!ax92x) & (ax91x) & (shiftx0x) & (!shiftx1x)) + ((ax94x) & (ax93x) & (!ax92x) & (ax91x) & (shiftx0x) & (shiftx1x)) + ((ax94x) & (ax93x) & (ax92x) & (!ax91x) & (!shiftx0x) & (!shiftx1x)) + ((ax94x) & (ax93x) & (ax92x) & (!ax91x) & (!shiftx0x) & (shiftx1x)) + ((ax94x) & (ax93x) & (ax92x) & (!ax91x) & (shiftx0x) & (!shiftx1x)) + ((ax94x) & (ax93x) & (ax92x) & (ax91x) & (!shiftx0x) & (!shiftx1x)) + ((ax94x) & (ax93x) & (ax92x) & (ax91x) & (!shiftx0x) & (shiftx1x)) + ((ax94x) & (ax93x) & (ax92x) & (ax91x) & (shiftx0x) & (!shiftx1x)) + ((ax94x) & (ax93x) & (ax92x) & (ax91x) & (shiftx0x) & (shiftx1x)));
	assign g115 = (((!ax86x) & (!ax85x) & (!ax84x) & (ax83x) & (shiftx0x) & (shiftx1x)) + ((!ax86x) & (!ax85x) & (ax84x) & (!ax83x) & (!shiftx0x) & (shiftx1x)) + ((!ax86x) & (!ax85x) & (ax84x) & (ax83x) & (!shiftx0x) & (shiftx1x)) + ((!ax86x) & (!ax85x) & (ax84x) & (ax83x) & (shiftx0x) & (shiftx1x)) + ((!ax86x) & (ax85x) & (!ax84x) & (!ax83x) & (shiftx0x) & (!shiftx1x)) + ((!ax86x) & (ax85x) & (!ax84x) & (ax83x) & (shiftx0x) & (!shiftx1x)) + ((!ax86x) & (ax85x) & (!ax84x) & (ax83x) & (shiftx0x) & (shiftx1x)) + ((!ax86x) & (ax85x) & (ax84x) & (!ax83x) & (!shiftx0x) & (shiftx1x)) + ((!ax86x) & (ax85x) & (ax84x) & (!ax83x) & (shiftx0x) & (!shiftx1x)) + ((!ax86x) & (ax85x) & (ax84x) & (ax83x) & (!shiftx0x) & (shiftx1x)) + ((!ax86x) & (ax85x) & (ax84x) & (ax83x) & (shiftx0x) & (!shiftx1x)) + ((!ax86x) & (ax85x) & (ax84x) & (ax83x) & (shiftx0x) & (shiftx1x)) + ((ax86x) & (!ax85x) & (!ax84x) & (!ax83x) & (!shiftx0x) & (!shiftx1x)) + ((ax86x) & (!ax85x) & (!ax84x) & (ax83x) & (!shiftx0x) & (!shiftx1x)) + ((ax86x) & (!ax85x) & (!ax84x) & (ax83x) & (shiftx0x) & (shiftx1x)) + ((ax86x) & (!ax85x) & (ax84x) & (!ax83x) & (!shiftx0x) & (!shiftx1x)) + ((ax86x) & (!ax85x) & (ax84x) & (!ax83x) & (!shiftx0x) & (shiftx1x)) + ((ax86x) & (!ax85x) & (ax84x) & (ax83x) & (!shiftx0x) & (!shiftx1x)) + ((ax86x) & (!ax85x) & (ax84x) & (ax83x) & (!shiftx0x) & (shiftx1x)) + ((ax86x) & (!ax85x) & (ax84x) & (ax83x) & (shiftx0x) & (shiftx1x)) + ((ax86x) & (ax85x) & (!ax84x) & (!ax83x) & (!shiftx0x) & (!shiftx1x)) + ((ax86x) & (ax85x) & (!ax84x) & (!ax83x) & (shiftx0x) & (!shiftx1x)) + ((ax86x) & (ax85x) & (!ax84x) & (ax83x) & (!shiftx0x) & (!shiftx1x)) + ((ax86x) & (ax85x) & (!ax84x) & (ax83x) & (shiftx0x) & (!shiftx1x)) + ((ax86x) & (ax85x) & (!ax84x) & (ax83x) & (shiftx0x) & (shiftx1x)) + ((ax86x) & (ax85x) & (ax84x) & (!ax83x) & (!shiftx0x) & (!shiftx1x)) + ((ax86x) & (ax85x) & (ax84x) & (!ax83x) & (!shiftx0x) & (shiftx1x)) + ((ax86x) & (ax85x) & (ax84x) & (!ax83x) & (shiftx0x) & (!shiftx1x)) + ((ax86x) & (ax85x) & (ax84x) & (ax83x) & (!shiftx0x) & (!shiftx1x)) + ((ax86x) & (ax85x) & (ax84x) & (ax83x) & (!shiftx0x) & (shiftx1x)) + ((ax86x) & (ax85x) & (ax84x) & (ax83x) & (shiftx0x) & (!shiftx1x)) + ((ax86x) & (ax85x) & (ax84x) & (ax83x) & (shiftx0x) & (shiftx1x)));
	assign g116 = (((!ax90x) & (!ax89x) & (!ax88x) & (ax87x) & (shiftx0x) & (shiftx1x)) + ((!ax90x) & (!ax89x) & (ax88x) & (!ax87x) & (!shiftx0x) & (shiftx1x)) + ((!ax90x) & (!ax89x) & (ax88x) & (ax87x) & (!shiftx0x) & (shiftx1x)) + ((!ax90x) & (!ax89x) & (ax88x) & (ax87x) & (shiftx0x) & (shiftx1x)) + ((!ax90x) & (ax89x) & (!ax88x) & (!ax87x) & (shiftx0x) & (!shiftx1x)) + ((!ax90x) & (ax89x) & (!ax88x) & (ax87x) & (shiftx0x) & (!shiftx1x)) + ((!ax90x) & (ax89x) & (!ax88x) & (ax87x) & (shiftx0x) & (shiftx1x)) + ((!ax90x) & (ax89x) & (ax88x) & (!ax87x) & (!shiftx0x) & (shiftx1x)) + ((!ax90x) & (ax89x) & (ax88x) & (!ax87x) & (shiftx0x) & (!shiftx1x)) + ((!ax90x) & (ax89x) & (ax88x) & (ax87x) & (!shiftx0x) & (shiftx1x)) + ((!ax90x) & (ax89x) & (ax88x) & (ax87x) & (shiftx0x) & (!shiftx1x)) + ((!ax90x) & (ax89x) & (ax88x) & (ax87x) & (shiftx0x) & (shiftx1x)) + ((ax90x) & (!ax89x) & (!ax88x) & (!ax87x) & (!shiftx0x) & (!shiftx1x)) + ((ax90x) & (!ax89x) & (!ax88x) & (ax87x) & (!shiftx0x) & (!shiftx1x)) + ((ax90x) & (!ax89x) & (!ax88x) & (ax87x) & (shiftx0x) & (shiftx1x)) + ((ax90x) & (!ax89x) & (ax88x) & (!ax87x) & (!shiftx0x) & (!shiftx1x)) + ((ax90x) & (!ax89x) & (ax88x) & (!ax87x) & (!shiftx0x) & (shiftx1x)) + ((ax90x) & (!ax89x) & (ax88x) & (ax87x) & (!shiftx0x) & (!shiftx1x)) + ((ax90x) & (!ax89x) & (ax88x) & (ax87x) & (!shiftx0x) & (shiftx1x)) + ((ax90x) & (!ax89x) & (ax88x) & (ax87x) & (shiftx0x) & (shiftx1x)) + ((ax90x) & (ax89x) & (!ax88x) & (!ax87x) & (!shiftx0x) & (!shiftx1x)) + ((ax90x) & (ax89x) & (!ax88x) & (!ax87x) & (shiftx0x) & (!shiftx1x)) + ((ax90x) & (ax89x) & (!ax88x) & (ax87x) & (!shiftx0x) & (!shiftx1x)) + ((ax90x) & (ax89x) & (!ax88x) & (ax87x) & (shiftx0x) & (!shiftx1x)) + ((ax90x) & (ax89x) & (!ax88x) & (ax87x) & (shiftx0x) & (shiftx1x)) + ((ax90x) & (ax89x) & (ax88x) & (!ax87x) & (!shiftx0x) & (!shiftx1x)) + ((ax90x) & (ax89x) & (ax88x) & (!ax87x) & (!shiftx0x) & (shiftx1x)) + ((ax90x) & (ax89x) & (ax88x) & (!ax87x) & (shiftx0x) & (!shiftx1x)) + ((ax90x) & (ax89x) & (ax88x) & (ax87x) & (!shiftx0x) & (!shiftx1x)) + ((ax90x) & (ax89x) & (ax88x) & (ax87x) & (!shiftx0x) & (shiftx1x)) + ((ax90x) & (ax89x) & (ax88x) & (ax87x) & (shiftx0x) & (!shiftx1x)) + ((ax90x) & (ax89x) & (ax88x) & (ax87x) & (shiftx0x) & (shiftx1x)));
	assign g117 = (((!shiftx2x) & (!shiftx3x) & (g113) & (!g114) & (!g115) & (!g116)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (!g114) & (!g115) & (g116)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (!g114) & (g115) & (!g116)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (!g114) & (g115) & (g116)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (g114) & (!g115) & (!g116)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (g114) & (!g115) & (g116)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (g114) & (g115) & (!g116)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (g114) & (g115) & (g116)) + ((!shiftx2x) & (shiftx3x) & (!g113) & (!g114) & (!g115) & (g116)) + ((!shiftx2x) & (shiftx3x) & (!g113) & (!g114) & (g115) & (g116)) + ((!shiftx2x) & (shiftx3x) & (!g113) & (g114) & (!g115) & (g116)) + ((!shiftx2x) & (shiftx3x) & (!g113) & (g114) & (g115) & (g116)) + ((!shiftx2x) & (shiftx3x) & (g113) & (!g114) & (!g115) & (g116)) + ((!shiftx2x) & (shiftx3x) & (g113) & (!g114) & (g115) & (g116)) + ((!shiftx2x) & (shiftx3x) & (g113) & (g114) & (!g115) & (g116)) + ((!shiftx2x) & (shiftx3x) & (g113) & (g114) & (g115) & (g116)) + ((shiftx2x) & (!shiftx3x) & (!g113) & (g114) & (!g115) & (!g116)) + ((shiftx2x) & (!shiftx3x) & (!g113) & (g114) & (!g115) & (g116)) + ((shiftx2x) & (!shiftx3x) & (!g113) & (g114) & (g115) & (!g116)) + ((shiftx2x) & (!shiftx3x) & (!g113) & (g114) & (g115) & (g116)) + ((shiftx2x) & (!shiftx3x) & (g113) & (g114) & (!g115) & (!g116)) + ((shiftx2x) & (!shiftx3x) & (g113) & (g114) & (!g115) & (g116)) + ((shiftx2x) & (!shiftx3x) & (g113) & (g114) & (g115) & (!g116)) + ((shiftx2x) & (!shiftx3x) & (g113) & (g114) & (g115) & (g116)) + ((shiftx2x) & (shiftx3x) & (!g113) & (!g114) & (g115) & (!g116)) + ((shiftx2x) & (shiftx3x) & (!g113) & (!g114) & (g115) & (g116)) + ((shiftx2x) & (shiftx3x) & (!g113) & (g114) & (g115) & (!g116)) + ((shiftx2x) & (shiftx3x) & (!g113) & (g114) & (g115) & (g116)) + ((shiftx2x) & (shiftx3x) & (g113) & (!g114) & (g115) & (!g116)) + ((shiftx2x) & (shiftx3x) & (g113) & (!g114) & (g115) & (g116)) + ((shiftx2x) & (shiftx3x) & (g113) & (g114) & (g115) & (!g116)) + ((shiftx2x) & (shiftx3x) & (g113) & (g114) & (g115) & (g116)));
	assign g118 = (((!ax2x) & (!ax1x) & (!ax0x) & (ax127x) & (shiftx0x) & (shiftx1x)) + ((!ax2x) & (!ax1x) & (ax0x) & (!ax127x) & (!shiftx0x) & (shiftx1x)) + ((!ax2x) & (!ax1x) & (ax0x) & (ax127x) & (!shiftx0x) & (shiftx1x)) + ((!ax2x) & (!ax1x) & (ax0x) & (ax127x) & (shiftx0x) & (shiftx1x)) + ((!ax2x) & (ax1x) & (!ax0x) & (!ax127x) & (shiftx0x) & (!shiftx1x)) + ((!ax2x) & (ax1x) & (!ax0x) & (ax127x) & (shiftx0x) & (!shiftx1x)) + ((!ax2x) & (ax1x) & (!ax0x) & (ax127x) & (shiftx0x) & (shiftx1x)) + ((!ax2x) & (ax1x) & (ax0x) & (!ax127x) & (!shiftx0x) & (shiftx1x)) + ((!ax2x) & (ax1x) & (ax0x) & (!ax127x) & (shiftx0x) & (!shiftx1x)) + ((!ax2x) & (ax1x) & (ax0x) & (ax127x) & (!shiftx0x) & (shiftx1x)) + ((!ax2x) & (ax1x) & (ax0x) & (ax127x) & (shiftx0x) & (!shiftx1x)) + ((!ax2x) & (ax1x) & (ax0x) & (ax127x) & (shiftx0x) & (shiftx1x)) + ((ax2x) & (!ax1x) & (!ax0x) & (!ax127x) & (!shiftx0x) & (!shiftx1x)) + ((ax2x) & (!ax1x) & (!ax0x) & (ax127x) & (!shiftx0x) & (!shiftx1x)) + ((ax2x) & (!ax1x) & (!ax0x) & (ax127x) & (shiftx0x) & (shiftx1x)) + ((ax2x) & (!ax1x) & (ax0x) & (!ax127x) & (!shiftx0x) & (!shiftx1x)) + ((ax2x) & (!ax1x) & (ax0x) & (!ax127x) & (!shiftx0x) & (shiftx1x)) + ((ax2x) & (!ax1x) & (ax0x) & (ax127x) & (!shiftx0x) & (!shiftx1x)) + ((ax2x) & (!ax1x) & (ax0x) & (ax127x) & (!shiftx0x) & (shiftx1x)) + ((ax2x) & (!ax1x) & (ax0x) & (ax127x) & (shiftx0x) & (shiftx1x)) + ((ax2x) & (ax1x) & (!ax0x) & (!ax127x) & (!shiftx0x) & (!shiftx1x)) + ((ax2x) & (ax1x) & (!ax0x) & (!ax127x) & (shiftx0x) & (!shiftx1x)) + ((ax2x) & (ax1x) & (!ax0x) & (ax127x) & (!shiftx0x) & (!shiftx1x)) + ((ax2x) & (ax1x) & (!ax0x) & (ax127x) & (shiftx0x) & (!shiftx1x)) + ((ax2x) & (ax1x) & (!ax0x) & (ax127x) & (shiftx0x) & (shiftx1x)) + ((ax2x) & (ax1x) & (ax0x) & (!ax127x) & (!shiftx0x) & (!shiftx1x)) + ((ax2x) & (ax1x) & (ax0x) & (!ax127x) & (!shiftx0x) & (shiftx1x)) + ((ax2x) & (ax1x) & (ax0x) & (!ax127x) & (shiftx0x) & (!shiftx1x)) + ((ax2x) & (ax1x) & (ax0x) & (ax127x) & (!shiftx0x) & (!shiftx1x)) + ((ax2x) & (ax1x) & (ax0x) & (ax127x) & (!shiftx0x) & (shiftx1x)) + ((ax2x) & (ax1x) & (ax0x) & (ax127x) & (shiftx0x) & (!shiftx1x)) + ((ax2x) & (ax1x) & (ax0x) & (ax127x) & (shiftx0x) & (shiftx1x)));
	assign g119 = (((!ax126x) & (!ax125x) & (!ax124x) & (ax123x) & (shiftx0x) & (shiftx1x)) + ((!ax126x) & (!ax125x) & (ax124x) & (!ax123x) & (!shiftx0x) & (shiftx1x)) + ((!ax126x) & (!ax125x) & (ax124x) & (ax123x) & (!shiftx0x) & (shiftx1x)) + ((!ax126x) & (!ax125x) & (ax124x) & (ax123x) & (shiftx0x) & (shiftx1x)) + ((!ax126x) & (ax125x) & (!ax124x) & (!ax123x) & (shiftx0x) & (!shiftx1x)) + ((!ax126x) & (ax125x) & (!ax124x) & (ax123x) & (shiftx0x) & (!shiftx1x)) + ((!ax126x) & (ax125x) & (!ax124x) & (ax123x) & (shiftx0x) & (shiftx1x)) + ((!ax126x) & (ax125x) & (ax124x) & (!ax123x) & (!shiftx0x) & (shiftx1x)) + ((!ax126x) & (ax125x) & (ax124x) & (!ax123x) & (shiftx0x) & (!shiftx1x)) + ((!ax126x) & (ax125x) & (ax124x) & (ax123x) & (!shiftx0x) & (shiftx1x)) + ((!ax126x) & (ax125x) & (ax124x) & (ax123x) & (shiftx0x) & (!shiftx1x)) + ((!ax126x) & (ax125x) & (ax124x) & (ax123x) & (shiftx0x) & (shiftx1x)) + ((ax126x) & (!ax125x) & (!ax124x) & (!ax123x) & (!shiftx0x) & (!shiftx1x)) + ((ax126x) & (!ax125x) & (!ax124x) & (ax123x) & (!shiftx0x) & (!shiftx1x)) + ((ax126x) & (!ax125x) & (!ax124x) & (ax123x) & (shiftx0x) & (shiftx1x)) + ((ax126x) & (!ax125x) & (ax124x) & (!ax123x) & (!shiftx0x) & (!shiftx1x)) + ((ax126x) & (!ax125x) & (ax124x) & (!ax123x) & (!shiftx0x) & (shiftx1x)) + ((ax126x) & (!ax125x) & (ax124x) & (ax123x) & (!shiftx0x) & (!shiftx1x)) + ((ax126x) & (!ax125x) & (ax124x) & (ax123x) & (!shiftx0x) & (shiftx1x)) + ((ax126x) & (!ax125x) & (ax124x) & (ax123x) & (shiftx0x) & (shiftx1x)) + ((ax126x) & (ax125x) & (!ax124x) & (!ax123x) & (!shiftx0x) & (!shiftx1x)) + ((ax126x) & (ax125x) & (!ax124x) & (!ax123x) & (shiftx0x) & (!shiftx1x)) + ((ax126x) & (ax125x) & (!ax124x) & (ax123x) & (!shiftx0x) & (!shiftx1x)) + ((ax126x) & (ax125x) & (!ax124x) & (ax123x) & (shiftx0x) & (!shiftx1x)) + ((ax126x) & (ax125x) & (!ax124x) & (ax123x) & (shiftx0x) & (shiftx1x)) + ((ax126x) & (ax125x) & (ax124x) & (!ax123x) & (!shiftx0x) & (!shiftx1x)) + ((ax126x) & (ax125x) & (ax124x) & (!ax123x) & (!shiftx0x) & (shiftx1x)) + ((ax126x) & (ax125x) & (ax124x) & (!ax123x) & (shiftx0x) & (!shiftx1x)) + ((ax126x) & (ax125x) & (ax124x) & (ax123x) & (!shiftx0x) & (!shiftx1x)) + ((ax126x) & (ax125x) & (ax124x) & (ax123x) & (!shiftx0x) & (shiftx1x)) + ((ax126x) & (ax125x) & (ax124x) & (ax123x) & (shiftx0x) & (!shiftx1x)) + ((ax126x) & (ax125x) & (ax124x) & (ax123x) & (shiftx0x) & (shiftx1x)));
	assign g120 = (((!ax118x) & (!ax117x) & (!ax116x) & (ax115x) & (shiftx0x) & (shiftx1x)) + ((!ax118x) & (!ax117x) & (ax116x) & (!ax115x) & (!shiftx0x) & (shiftx1x)) + ((!ax118x) & (!ax117x) & (ax116x) & (ax115x) & (!shiftx0x) & (shiftx1x)) + ((!ax118x) & (!ax117x) & (ax116x) & (ax115x) & (shiftx0x) & (shiftx1x)) + ((!ax118x) & (ax117x) & (!ax116x) & (!ax115x) & (shiftx0x) & (!shiftx1x)) + ((!ax118x) & (ax117x) & (!ax116x) & (ax115x) & (shiftx0x) & (!shiftx1x)) + ((!ax118x) & (ax117x) & (!ax116x) & (ax115x) & (shiftx0x) & (shiftx1x)) + ((!ax118x) & (ax117x) & (ax116x) & (!ax115x) & (!shiftx0x) & (shiftx1x)) + ((!ax118x) & (ax117x) & (ax116x) & (!ax115x) & (shiftx0x) & (!shiftx1x)) + ((!ax118x) & (ax117x) & (ax116x) & (ax115x) & (!shiftx0x) & (shiftx1x)) + ((!ax118x) & (ax117x) & (ax116x) & (ax115x) & (shiftx0x) & (!shiftx1x)) + ((!ax118x) & (ax117x) & (ax116x) & (ax115x) & (shiftx0x) & (shiftx1x)) + ((ax118x) & (!ax117x) & (!ax116x) & (!ax115x) & (!shiftx0x) & (!shiftx1x)) + ((ax118x) & (!ax117x) & (!ax116x) & (ax115x) & (!shiftx0x) & (!shiftx1x)) + ((ax118x) & (!ax117x) & (!ax116x) & (ax115x) & (shiftx0x) & (shiftx1x)) + ((ax118x) & (!ax117x) & (ax116x) & (!ax115x) & (!shiftx0x) & (!shiftx1x)) + ((ax118x) & (!ax117x) & (ax116x) & (!ax115x) & (!shiftx0x) & (shiftx1x)) + ((ax118x) & (!ax117x) & (ax116x) & (ax115x) & (!shiftx0x) & (!shiftx1x)) + ((ax118x) & (!ax117x) & (ax116x) & (ax115x) & (!shiftx0x) & (shiftx1x)) + ((ax118x) & (!ax117x) & (ax116x) & (ax115x) & (shiftx0x) & (shiftx1x)) + ((ax118x) & (ax117x) & (!ax116x) & (!ax115x) & (!shiftx0x) & (!shiftx1x)) + ((ax118x) & (ax117x) & (!ax116x) & (!ax115x) & (shiftx0x) & (!shiftx1x)) + ((ax118x) & (ax117x) & (!ax116x) & (ax115x) & (!shiftx0x) & (!shiftx1x)) + ((ax118x) & (ax117x) & (!ax116x) & (ax115x) & (shiftx0x) & (!shiftx1x)) + ((ax118x) & (ax117x) & (!ax116x) & (ax115x) & (shiftx0x) & (shiftx1x)) + ((ax118x) & (ax117x) & (ax116x) & (!ax115x) & (!shiftx0x) & (!shiftx1x)) + ((ax118x) & (ax117x) & (ax116x) & (!ax115x) & (!shiftx0x) & (shiftx1x)) + ((ax118x) & (ax117x) & (ax116x) & (!ax115x) & (shiftx0x) & (!shiftx1x)) + ((ax118x) & (ax117x) & (ax116x) & (ax115x) & (!shiftx0x) & (!shiftx1x)) + ((ax118x) & (ax117x) & (ax116x) & (ax115x) & (!shiftx0x) & (shiftx1x)) + ((ax118x) & (ax117x) & (ax116x) & (ax115x) & (shiftx0x) & (!shiftx1x)) + ((ax118x) & (ax117x) & (ax116x) & (ax115x) & (shiftx0x) & (shiftx1x)));
	assign g121 = (((!ax122x) & (!ax121x) & (!ax120x) & (ax119x) & (shiftx0x) & (shiftx1x)) + ((!ax122x) & (!ax121x) & (ax120x) & (!ax119x) & (!shiftx0x) & (shiftx1x)) + ((!ax122x) & (!ax121x) & (ax120x) & (ax119x) & (!shiftx0x) & (shiftx1x)) + ((!ax122x) & (!ax121x) & (ax120x) & (ax119x) & (shiftx0x) & (shiftx1x)) + ((!ax122x) & (ax121x) & (!ax120x) & (!ax119x) & (shiftx0x) & (!shiftx1x)) + ((!ax122x) & (ax121x) & (!ax120x) & (ax119x) & (shiftx0x) & (!shiftx1x)) + ((!ax122x) & (ax121x) & (!ax120x) & (ax119x) & (shiftx0x) & (shiftx1x)) + ((!ax122x) & (ax121x) & (ax120x) & (!ax119x) & (!shiftx0x) & (shiftx1x)) + ((!ax122x) & (ax121x) & (ax120x) & (!ax119x) & (shiftx0x) & (!shiftx1x)) + ((!ax122x) & (ax121x) & (ax120x) & (ax119x) & (!shiftx0x) & (shiftx1x)) + ((!ax122x) & (ax121x) & (ax120x) & (ax119x) & (shiftx0x) & (!shiftx1x)) + ((!ax122x) & (ax121x) & (ax120x) & (ax119x) & (shiftx0x) & (shiftx1x)) + ((ax122x) & (!ax121x) & (!ax120x) & (!ax119x) & (!shiftx0x) & (!shiftx1x)) + ((ax122x) & (!ax121x) & (!ax120x) & (ax119x) & (!shiftx0x) & (!shiftx1x)) + ((ax122x) & (!ax121x) & (!ax120x) & (ax119x) & (shiftx0x) & (shiftx1x)) + ((ax122x) & (!ax121x) & (ax120x) & (!ax119x) & (!shiftx0x) & (!shiftx1x)) + ((ax122x) & (!ax121x) & (ax120x) & (!ax119x) & (!shiftx0x) & (shiftx1x)) + ((ax122x) & (!ax121x) & (ax120x) & (ax119x) & (!shiftx0x) & (!shiftx1x)) + ((ax122x) & (!ax121x) & (ax120x) & (ax119x) & (!shiftx0x) & (shiftx1x)) + ((ax122x) & (!ax121x) & (ax120x) & (ax119x) & (shiftx0x) & (shiftx1x)) + ((ax122x) & (ax121x) & (!ax120x) & (!ax119x) & (!shiftx0x) & (!shiftx1x)) + ((ax122x) & (ax121x) & (!ax120x) & (!ax119x) & (shiftx0x) & (!shiftx1x)) + ((ax122x) & (ax121x) & (!ax120x) & (ax119x) & (!shiftx0x) & (!shiftx1x)) + ((ax122x) & (ax121x) & (!ax120x) & (ax119x) & (shiftx0x) & (!shiftx1x)) + ((ax122x) & (ax121x) & (!ax120x) & (ax119x) & (shiftx0x) & (shiftx1x)) + ((ax122x) & (ax121x) & (ax120x) & (!ax119x) & (!shiftx0x) & (!shiftx1x)) + ((ax122x) & (ax121x) & (ax120x) & (!ax119x) & (!shiftx0x) & (shiftx1x)) + ((ax122x) & (ax121x) & (ax120x) & (!ax119x) & (shiftx0x) & (!shiftx1x)) + ((ax122x) & (ax121x) & (ax120x) & (ax119x) & (!shiftx0x) & (!shiftx1x)) + ((ax122x) & (ax121x) & (ax120x) & (ax119x) & (!shiftx0x) & (shiftx1x)) + ((ax122x) & (ax121x) & (ax120x) & (ax119x) & (shiftx0x) & (!shiftx1x)) + ((ax122x) & (ax121x) & (ax120x) & (ax119x) & (shiftx0x) & (shiftx1x)));
	assign g122 = (((!shiftx2x) & (!shiftx3x) & (g118) & (!g119) & (!g120) & (!g121)) + ((!shiftx2x) & (!shiftx3x) & (g118) & (!g119) & (!g120) & (g121)) + ((!shiftx2x) & (!shiftx3x) & (g118) & (!g119) & (g120) & (!g121)) + ((!shiftx2x) & (!shiftx3x) & (g118) & (!g119) & (g120) & (g121)) + ((!shiftx2x) & (!shiftx3x) & (g118) & (g119) & (!g120) & (!g121)) + ((!shiftx2x) & (!shiftx3x) & (g118) & (g119) & (!g120) & (g121)) + ((!shiftx2x) & (!shiftx3x) & (g118) & (g119) & (g120) & (!g121)) + ((!shiftx2x) & (!shiftx3x) & (g118) & (g119) & (g120) & (g121)) + ((!shiftx2x) & (shiftx3x) & (!g118) & (!g119) & (!g120) & (g121)) + ((!shiftx2x) & (shiftx3x) & (!g118) & (!g119) & (g120) & (g121)) + ((!shiftx2x) & (shiftx3x) & (!g118) & (g119) & (!g120) & (g121)) + ((!shiftx2x) & (shiftx3x) & (!g118) & (g119) & (g120) & (g121)) + ((!shiftx2x) & (shiftx3x) & (g118) & (!g119) & (!g120) & (g121)) + ((!shiftx2x) & (shiftx3x) & (g118) & (!g119) & (g120) & (g121)) + ((!shiftx2x) & (shiftx3x) & (g118) & (g119) & (!g120) & (g121)) + ((!shiftx2x) & (shiftx3x) & (g118) & (g119) & (g120) & (g121)) + ((shiftx2x) & (!shiftx3x) & (!g118) & (g119) & (!g120) & (!g121)) + ((shiftx2x) & (!shiftx3x) & (!g118) & (g119) & (!g120) & (g121)) + ((shiftx2x) & (!shiftx3x) & (!g118) & (g119) & (g120) & (!g121)) + ((shiftx2x) & (!shiftx3x) & (!g118) & (g119) & (g120) & (g121)) + ((shiftx2x) & (!shiftx3x) & (g118) & (g119) & (!g120) & (!g121)) + ((shiftx2x) & (!shiftx3x) & (g118) & (g119) & (!g120) & (g121)) + ((shiftx2x) & (!shiftx3x) & (g118) & (g119) & (g120) & (!g121)) + ((shiftx2x) & (!shiftx3x) & (g118) & (g119) & (g120) & (g121)) + ((shiftx2x) & (shiftx3x) & (!g118) & (!g119) & (g120) & (!g121)) + ((shiftx2x) & (shiftx3x) & (!g118) & (!g119) & (g120) & (g121)) + ((shiftx2x) & (shiftx3x) & (!g118) & (g119) & (g120) & (!g121)) + ((shiftx2x) & (shiftx3x) & (!g118) & (g119) & (g120) & (g121)) + ((shiftx2x) & (shiftx3x) & (g118) & (!g119) & (g120) & (!g121)) + ((shiftx2x) & (shiftx3x) & (g118) & (!g119) & (g120) & (g121)) + ((shiftx2x) & (shiftx3x) & (g118) & (g119) & (g120) & (!g121)) + ((shiftx2x) & (shiftx3x) & (g118) & (g119) & (g120) & (g121)));
	assign g123 = (((!ax114x) & (!ax113x) & (!ax112x) & (ax111x) & (shiftx0x) & (shiftx1x)) + ((!ax114x) & (!ax113x) & (ax112x) & (!ax111x) & (!shiftx0x) & (shiftx1x)) + ((!ax114x) & (!ax113x) & (ax112x) & (ax111x) & (!shiftx0x) & (shiftx1x)) + ((!ax114x) & (!ax113x) & (ax112x) & (ax111x) & (shiftx0x) & (shiftx1x)) + ((!ax114x) & (ax113x) & (!ax112x) & (!ax111x) & (shiftx0x) & (!shiftx1x)) + ((!ax114x) & (ax113x) & (!ax112x) & (ax111x) & (shiftx0x) & (!shiftx1x)) + ((!ax114x) & (ax113x) & (!ax112x) & (ax111x) & (shiftx0x) & (shiftx1x)) + ((!ax114x) & (ax113x) & (ax112x) & (!ax111x) & (!shiftx0x) & (shiftx1x)) + ((!ax114x) & (ax113x) & (ax112x) & (!ax111x) & (shiftx0x) & (!shiftx1x)) + ((!ax114x) & (ax113x) & (ax112x) & (ax111x) & (!shiftx0x) & (shiftx1x)) + ((!ax114x) & (ax113x) & (ax112x) & (ax111x) & (shiftx0x) & (!shiftx1x)) + ((!ax114x) & (ax113x) & (ax112x) & (ax111x) & (shiftx0x) & (shiftx1x)) + ((ax114x) & (!ax113x) & (!ax112x) & (!ax111x) & (!shiftx0x) & (!shiftx1x)) + ((ax114x) & (!ax113x) & (!ax112x) & (ax111x) & (!shiftx0x) & (!shiftx1x)) + ((ax114x) & (!ax113x) & (!ax112x) & (ax111x) & (shiftx0x) & (shiftx1x)) + ((ax114x) & (!ax113x) & (ax112x) & (!ax111x) & (!shiftx0x) & (!shiftx1x)) + ((ax114x) & (!ax113x) & (ax112x) & (!ax111x) & (!shiftx0x) & (shiftx1x)) + ((ax114x) & (!ax113x) & (ax112x) & (ax111x) & (!shiftx0x) & (!shiftx1x)) + ((ax114x) & (!ax113x) & (ax112x) & (ax111x) & (!shiftx0x) & (shiftx1x)) + ((ax114x) & (!ax113x) & (ax112x) & (ax111x) & (shiftx0x) & (shiftx1x)) + ((ax114x) & (ax113x) & (!ax112x) & (!ax111x) & (!shiftx0x) & (!shiftx1x)) + ((ax114x) & (ax113x) & (!ax112x) & (!ax111x) & (shiftx0x) & (!shiftx1x)) + ((ax114x) & (ax113x) & (!ax112x) & (ax111x) & (!shiftx0x) & (!shiftx1x)) + ((ax114x) & (ax113x) & (!ax112x) & (ax111x) & (shiftx0x) & (!shiftx1x)) + ((ax114x) & (ax113x) & (!ax112x) & (ax111x) & (shiftx0x) & (shiftx1x)) + ((ax114x) & (ax113x) & (ax112x) & (!ax111x) & (!shiftx0x) & (!shiftx1x)) + ((ax114x) & (ax113x) & (ax112x) & (!ax111x) & (!shiftx0x) & (shiftx1x)) + ((ax114x) & (ax113x) & (ax112x) & (!ax111x) & (shiftx0x) & (!shiftx1x)) + ((ax114x) & (ax113x) & (ax112x) & (ax111x) & (!shiftx0x) & (!shiftx1x)) + ((ax114x) & (ax113x) & (ax112x) & (ax111x) & (!shiftx0x) & (shiftx1x)) + ((ax114x) & (ax113x) & (ax112x) & (ax111x) & (shiftx0x) & (!shiftx1x)) + ((ax114x) & (ax113x) & (ax112x) & (ax111x) & (shiftx0x) & (shiftx1x)));
	assign g124 = (((!ax110x) & (!ax109x) & (!ax108x) & (ax107x) & (shiftx0x) & (shiftx1x)) + ((!ax110x) & (!ax109x) & (ax108x) & (!ax107x) & (!shiftx0x) & (shiftx1x)) + ((!ax110x) & (!ax109x) & (ax108x) & (ax107x) & (!shiftx0x) & (shiftx1x)) + ((!ax110x) & (!ax109x) & (ax108x) & (ax107x) & (shiftx0x) & (shiftx1x)) + ((!ax110x) & (ax109x) & (!ax108x) & (!ax107x) & (shiftx0x) & (!shiftx1x)) + ((!ax110x) & (ax109x) & (!ax108x) & (ax107x) & (shiftx0x) & (!shiftx1x)) + ((!ax110x) & (ax109x) & (!ax108x) & (ax107x) & (shiftx0x) & (shiftx1x)) + ((!ax110x) & (ax109x) & (ax108x) & (!ax107x) & (!shiftx0x) & (shiftx1x)) + ((!ax110x) & (ax109x) & (ax108x) & (!ax107x) & (shiftx0x) & (!shiftx1x)) + ((!ax110x) & (ax109x) & (ax108x) & (ax107x) & (!shiftx0x) & (shiftx1x)) + ((!ax110x) & (ax109x) & (ax108x) & (ax107x) & (shiftx0x) & (!shiftx1x)) + ((!ax110x) & (ax109x) & (ax108x) & (ax107x) & (shiftx0x) & (shiftx1x)) + ((ax110x) & (!ax109x) & (!ax108x) & (!ax107x) & (!shiftx0x) & (!shiftx1x)) + ((ax110x) & (!ax109x) & (!ax108x) & (ax107x) & (!shiftx0x) & (!shiftx1x)) + ((ax110x) & (!ax109x) & (!ax108x) & (ax107x) & (shiftx0x) & (shiftx1x)) + ((ax110x) & (!ax109x) & (ax108x) & (!ax107x) & (!shiftx0x) & (!shiftx1x)) + ((ax110x) & (!ax109x) & (ax108x) & (!ax107x) & (!shiftx0x) & (shiftx1x)) + ((ax110x) & (!ax109x) & (ax108x) & (ax107x) & (!shiftx0x) & (!shiftx1x)) + ((ax110x) & (!ax109x) & (ax108x) & (ax107x) & (!shiftx0x) & (shiftx1x)) + ((ax110x) & (!ax109x) & (ax108x) & (ax107x) & (shiftx0x) & (shiftx1x)) + ((ax110x) & (ax109x) & (!ax108x) & (!ax107x) & (!shiftx0x) & (!shiftx1x)) + ((ax110x) & (ax109x) & (!ax108x) & (!ax107x) & (shiftx0x) & (!shiftx1x)) + ((ax110x) & (ax109x) & (!ax108x) & (ax107x) & (!shiftx0x) & (!shiftx1x)) + ((ax110x) & (ax109x) & (!ax108x) & (ax107x) & (shiftx0x) & (!shiftx1x)) + ((ax110x) & (ax109x) & (!ax108x) & (ax107x) & (shiftx0x) & (shiftx1x)) + ((ax110x) & (ax109x) & (ax108x) & (!ax107x) & (!shiftx0x) & (!shiftx1x)) + ((ax110x) & (ax109x) & (ax108x) & (!ax107x) & (!shiftx0x) & (shiftx1x)) + ((ax110x) & (ax109x) & (ax108x) & (!ax107x) & (shiftx0x) & (!shiftx1x)) + ((ax110x) & (ax109x) & (ax108x) & (ax107x) & (!shiftx0x) & (!shiftx1x)) + ((ax110x) & (ax109x) & (ax108x) & (ax107x) & (!shiftx0x) & (shiftx1x)) + ((ax110x) & (ax109x) & (ax108x) & (ax107x) & (shiftx0x) & (!shiftx1x)) + ((ax110x) & (ax109x) & (ax108x) & (ax107x) & (shiftx0x) & (shiftx1x)));
	assign g125 = (((!ax102x) & (!ax101x) & (!ax100x) & (ax99x) & (shiftx0x) & (shiftx1x)) + ((!ax102x) & (!ax101x) & (ax100x) & (!ax99x) & (!shiftx0x) & (shiftx1x)) + ((!ax102x) & (!ax101x) & (ax100x) & (ax99x) & (!shiftx0x) & (shiftx1x)) + ((!ax102x) & (!ax101x) & (ax100x) & (ax99x) & (shiftx0x) & (shiftx1x)) + ((!ax102x) & (ax101x) & (!ax100x) & (!ax99x) & (shiftx0x) & (!shiftx1x)) + ((!ax102x) & (ax101x) & (!ax100x) & (ax99x) & (shiftx0x) & (!shiftx1x)) + ((!ax102x) & (ax101x) & (!ax100x) & (ax99x) & (shiftx0x) & (shiftx1x)) + ((!ax102x) & (ax101x) & (ax100x) & (!ax99x) & (!shiftx0x) & (shiftx1x)) + ((!ax102x) & (ax101x) & (ax100x) & (!ax99x) & (shiftx0x) & (!shiftx1x)) + ((!ax102x) & (ax101x) & (ax100x) & (ax99x) & (!shiftx0x) & (shiftx1x)) + ((!ax102x) & (ax101x) & (ax100x) & (ax99x) & (shiftx0x) & (!shiftx1x)) + ((!ax102x) & (ax101x) & (ax100x) & (ax99x) & (shiftx0x) & (shiftx1x)) + ((ax102x) & (!ax101x) & (!ax100x) & (!ax99x) & (!shiftx0x) & (!shiftx1x)) + ((ax102x) & (!ax101x) & (!ax100x) & (ax99x) & (!shiftx0x) & (!shiftx1x)) + ((ax102x) & (!ax101x) & (!ax100x) & (ax99x) & (shiftx0x) & (shiftx1x)) + ((ax102x) & (!ax101x) & (ax100x) & (!ax99x) & (!shiftx0x) & (!shiftx1x)) + ((ax102x) & (!ax101x) & (ax100x) & (!ax99x) & (!shiftx0x) & (shiftx1x)) + ((ax102x) & (!ax101x) & (ax100x) & (ax99x) & (!shiftx0x) & (!shiftx1x)) + ((ax102x) & (!ax101x) & (ax100x) & (ax99x) & (!shiftx0x) & (shiftx1x)) + ((ax102x) & (!ax101x) & (ax100x) & (ax99x) & (shiftx0x) & (shiftx1x)) + ((ax102x) & (ax101x) & (!ax100x) & (!ax99x) & (!shiftx0x) & (!shiftx1x)) + ((ax102x) & (ax101x) & (!ax100x) & (!ax99x) & (shiftx0x) & (!shiftx1x)) + ((ax102x) & (ax101x) & (!ax100x) & (ax99x) & (!shiftx0x) & (!shiftx1x)) + ((ax102x) & (ax101x) & (!ax100x) & (ax99x) & (shiftx0x) & (!shiftx1x)) + ((ax102x) & (ax101x) & (!ax100x) & (ax99x) & (shiftx0x) & (shiftx1x)) + ((ax102x) & (ax101x) & (ax100x) & (!ax99x) & (!shiftx0x) & (!shiftx1x)) + ((ax102x) & (ax101x) & (ax100x) & (!ax99x) & (!shiftx0x) & (shiftx1x)) + ((ax102x) & (ax101x) & (ax100x) & (!ax99x) & (shiftx0x) & (!shiftx1x)) + ((ax102x) & (ax101x) & (ax100x) & (ax99x) & (!shiftx0x) & (!shiftx1x)) + ((ax102x) & (ax101x) & (ax100x) & (ax99x) & (!shiftx0x) & (shiftx1x)) + ((ax102x) & (ax101x) & (ax100x) & (ax99x) & (shiftx0x) & (!shiftx1x)) + ((ax102x) & (ax101x) & (ax100x) & (ax99x) & (shiftx0x) & (shiftx1x)));
	assign g126 = (((!ax106x) & (!ax105x) & (!ax104x) & (ax103x) & (shiftx0x) & (shiftx1x)) + ((!ax106x) & (!ax105x) & (ax104x) & (!ax103x) & (!shiftx0x) & (shiftx1x)) + ((!ax106x) & (!ax105x) & (ax104x) & (ax103x) & (!shiftx0x) & (shiftx1x)) + ((!ax106x) & (!ax105x) & (ax104x) & (ax103x) & (shiftx0x) & (shiftx1x)) + ((!ax106x) & (ax105x) & (!ax104x) & (!ax103x) & (shiftx0x) & (!shiftx1x)) + ((!ax106x) & (ax105x) & (!ax104x) & (ax103x) & (shiftx0x) & (!shiftx1x)) + ((!ax106x) & (ax105x) & (!ax104x) & (ax103x) & (shiftx0x) & (shiftx1x)) + ((!ax106x) & (ax105x) & (ax104x) & (!ax103x) & (!shiftx0x) & (shiftx1x)) + ((!ax106x) & (ax105x) & (ax104x) & (!ax103x) & (shiftx0x) & (!shiftx1x)) + ((!ax106x) & (ax105x) & (ax104x) & (ax103x) & (!shiftx0x) & (shiftx1x)) + ((!ax106x) & (ax105x) & (ax104x) & (ax103x) & (shiftx0x) & (!shiftx1x)) + ((!ax106x) & (ax105x) & (ax104x) & (ax103x) & (shiftx0x) & (shiftx1x)) + ((ax106x) & (!ax105x) & (!ax104x) & (!ax103x) & (!shiftx0x) & (!shiftx1x)) + ((ax106x) & (!ax105x) & (!ax104x) & (ax103x) & (!shiftx0x) & (!shiftx1x)) + ((ax106x) & (!ax105x) & (!ax104x) & (ax103x) & (shiftx0x) & (shiftx1x)) + ((ax106x) & (!ax105x) & (ax104x) & (!ax103x) & (!shiftx0x) & (!shiftx1x)) + ((ax106x) & (!ax105x) & (ax104x) & (!ax103x) & (!shiftx0x) & (shiftx1x)) + ((ax106x) & (!ax105x) & (ax104x) & (ax103x) & (!shiftx0x) & (!shiftx1x)) + ((ax106x) & (!ax105x) & (ax104x) & (ax103x) & (!shiftx0x) & (shiftx1x)) + ((ax106x) & (!ax105x) & (ax104x) & (ax103x) & (shiftx0x) & (shiftx1x)) + ((ax106x) & (ax105x) & (!ax104x) & (!ax103x) & (!shiftx0x) & (!shiftx1x)) + ((ax106x) & (ax105x) & (!ax104x) & (!ax103x) & (shiftx0x) & (!shiftx1x)) + ((ax106x) & (ax105x) & (!ax104x) & (ax103x) & (!shiftx0x) & (!shiftx1x)) + ((ax106x) & (ax105x) & (!ax104x) & (ax103x) & (shiftx0x) & (!shiftx1x)) + ((ax106x) & (ax105x) & (!ax104x) & (ax103x) & (shiftx0x) & (shiftx1x)) + ((ax106x) & (ax105x) & (ax104x) & (!ax103x) & (!shiftx0x) & (!shiftx1x)) + ((ax106x) & (ax105x) & (ax104x) & (!ax103x) & (!shiftx0x) & (shiftx1x)) + ((ax106x) & (ax105x) & (ax104x) & (!ax103x) & (shiftx0x) & (!shiftx1x)) + ((ax106x) & (ax105x) & (ax104x) & (ax103x) & (!shiftx0x) & (!shiftx1x)) + ((ax106x) & (ax105x) & (ax104x) & (ax103x) & (!shiftx0x) & (shiftx1x)) + ((ax106x) & (ax105x) & (ax104x) & (ax103x) & (shiftx0x) & (!shiftx1x)) + ((ax106x) & (ax105x) & (ax104x) & (ax103x) & (shiftx0x) & (shiftx1x)));
	assign g127 = (((!shiftx2x) & (!shiftx3x) & (g123) & (!g124) & (!g125) & (!g126)) + ((!shiftx2x) & (!shiftx3x) & (g123) & (!g124) & (!g125) & (g126)) + ((!shiftx2x) & (!shiftx3x) & (g123) & (!g124) & (g125) & (!g126)) + ((!shiftx2x) & (!shiftx3x) & (g123) & (!g124) & (g125) & (g126)) + ((!shiftx2x) & (!shiftx3x) & (g123) & (g124) & (!g125) & (!g126)) + ((!shiftx2x) & (!shiftx3x) & (g123) & (g124) & (!g125) & (g126)) + ((!shiftx2x) & (!shiftx3x) & (g123) & (g124) & (g125) & (!g126)) + ((!shiftx2x) & (!shiftx3x) & (g123) & (g124) & (g125) & (g126)) + ((!shiftx2x) & (shiftx3x) & (!g123) & (!g124) & (!g125) & (g126)) + ((!shiftx2x) & (shiftx3x) & (!g123) & (!g124) & (g125) & (g126)) + ((!shiftx2x) & (shiftx3x) & (!g123) & (g124) & (!g125) & (g126)) + ((!shiftx2x) & (shiftx3x) & (!g123) & (g124) & (g125) & (g126)) + ((!shiftx2x) & (shiftx3x) & (g123) & (!g124) & (!g125) & (g126)) + ((!shiftx2x) & (shiftx3x) & (g123) & (!g124) & (g125) & (g126)) + ((!shiftx2x) & (shiftx3x) & (g123) & (g124) & (!g125) & (g126)) + ((!shiftx2x) & (shiftx3x) & (g123) & (g124) & (g125) & (g126)) + ((shiftx2x) & (!shiftx3x) & (!g123) & (g124) & (!g125) & (!g126)) + ((shiftx2x) & (!shiftx3x) & (!g123) & (g124) & (!g125) & (g126)) + ((shiftx2x) & (!shiftx3x) & (!g123) & (g124) & (g125) & (!g126)) + ((shiftx2x) & (!shiftx3x) & (!g123) & (g124) & (g125) & (g126)) + ((shiftx2x) & (!shiftx3x) & (g123) & (g124) & (!g125) & (!g126)) + ((shiftx2x) & (!shiftx3x) & (g123) & (g124) & (!g125) & (g126)) + ((shiftx2x) & (!shiftx3x) & (g123) & (g124) & (g125) & (!g126)) + ((shiftx2x) & (!shiftx3x) & (g123) & (g124) & (g125) & (g126)) + ((shiftx2x) & (shiftx3x) & (!g123) & (!g124) & (g125) & (!g126)) + ((shiftx2x) & (shiftx3x) & (!g123) & (!g124) & (g125) & (g126)) + ((shiftx2x) & (shiftx3x) & (!g123) & (g124) & (g125) & (!g126)) + ((shiftx2x) & (shiftx3x) & (!g123) & (g124) & (g125) & (g126)) + ((shiftx2x) & (shiftx3x) & (g123) & (!g124) & (g125) & (!g126)) + ((shiftx2x) & (shiftx3x) & (g123) & (!g124) & (g125) & (g126)) + ((shiftx2x) & (shiftx3x) & (g123) & (g124) & (g125) & (!g126)) + ((shiftx2x) & (shiftx3x) & (g123) & (g124) & (g125) & (g126)));
	assign g128 = (((!shiftx4x) & (!shiftx5x) & (!g112) & (!g117) & (g122) & (!g127)) + ((!shiftx4x) & (!shiftx5x) & (!g112) & (!g117) & (g122) & (g127)) + ((!shiftx4x) & (!shiftx5x) & (!g112) & (g117) & (g122) & (!g127)) + ((!shiftx4x) & (!shiftx5x) & (!g112) & (g117) & (g122) & (g127)) + ((!shiftx4x) & (!shiftx5x) & (g112) & (!g117) & (g122) & (!g127)) + ((!shiftx4x) & (!shiftx5x) & (g112) & (!g117) & (g122) & (g127)) + ((!shiftx4x) & (!shiftx5x) & (g112) & (g117) & (g122) & (!g127)) + ((!shiftx4x) & (!shiftx5x) & (g112) & (g117) & (g122) & (g127)) + ((!shiftx4x) & (shiftx5x) & (!g112) & (g117) & (!g122) & (!g127)) + ((!shiftx4x) & (shiftx5x) & (!g112) & (g117) & (!g122) & (g127)) + ((!shiftx4x) & (shiftx5x) & (!g112) & (g117) & (g122) & (!g127)) + ((!shiftx4x) & (shiftx5x) & (!g112) & (g117) & (g122) & (g127)) + ((!shiftx4x) & (shiftx5x) & (g112) & (g117) & (!g122) & (!g127)) + ((!shiftx4x) & (shiftx5x) & (g112) & (g117) & (!g122) & (g127)) + ((!shiftx4x) & (shiftx5x) & (g112) & (g117) & (g122) & (!g127)) + ((!shiftx4x) & (shiftx5x) & (g112) & (g117) & (g122) & (g127)) + ((shiftx4x) & (!shiftx5x) & (!g112) & (!g117) & (!g122) & (g127)) + ((shiftx4x) & (!shiftx5x) & (!g112) & (!g117) & (g122) & (g127)) + ((shiftx4x) & (!shiftx5x) & (!g112) & (g117) & (!g122) & (g127)) + ((shiftx4x) & (!shiftx5x) & (!g112) & (g117) & (g122) & (g127)) + ((shiftx4x) & (!shiftx5x) & (g112) & (!g117) & (!g122) & (g127)) + ((shiftx4x) & (!shiftx5x) & (g112) & (!g117) & (g122) & (g127)) + ((shiftx4x) & (!shiftx5x) & (g112) & (g117) & (!g122) & (g127)) + ((shiftx4x) & (!shiftx5x) & (g112) & (g117) & (g122) & (g127)) + ((shiftx4x) & (shiftx5x) & (g112) & (!g117) & (!g122) & (!g127)) + ((shiftx4x) & (shiftx5x) & (g112) & (!g117) & (!g122) & (g127)) + ((shiftx4x) & (shiftx5x) & (g112) & (!g117) & (g122) & (!g127)) + ((shiftx4x) & (shiftx5x) & (g112) & (!g117) & (g122) & (g127)) + ((shiftx4x) & (shiftx5x) & (g112) & (g117) & (!g122) & (!g127)) + ((shiftx4x) & (shiftx5x) & (g112) & (g117) & (!g122) & (g127)) + ((shiftx4x) & (shiftx5x) & (g112) & (g117) & (g122) & (!g127)) + ((shiftx4x) & (shiftx5x) & (g112) & (g117) & (g122) & (g127)));
	assign resultx2x = (((!shiftx6x) & (sk[0]) & (!g107) & (g128)) + ((!shiftx6x) & (sk[0]) & (g107) & (g128)) + ((shiftx6x) & (!sk[0]) & (!g107) & (!g128)) + ((shiftx6x) & (!sk[0]) & (!g107) & (g128)) + ((shiftx6x) & (!sk[0]) & (g107) & (!g128)) + ((shiftx6x) & (!sk[0]) & (g107) & (g128)) + ((shiftx6x) & (sk[0]) & (g107) & (!g128)) + ((shiftx6x) & (sk[0]) & (g107) & (g128)));
	assign g130 = (((!shiftx0x) & (!shiftx1x) & (!ax64x) & (ax67x) & (!ax66x) & (!ax65x)) + ((!shiftx0x) & (!shiftx1x) & (!ax64x) & (ax67x) & (!ax66x) & (ax65x)) + ((!shiftx0x) & (!shiftx1x) & (!ax64x) & (ax67x) & (ax66x) & (!ax65x)) + ((!shiftx0x) & (!shiftx1x) & (!ax64x) & (ax67x) & (ax66x) & (ax65x)) + ((!shiftx0x) & (!shiftx1x) & (ax64x) & (ax67x) & (!ax66x) & (!ax65x)) + ((!shiftx0x) & (!shiftx1x) & (ax64x) & (ax67x) & (!ax66x) & (ax65x)) + ((!shiftx0x) & (!shiftx1x) & (ax64x) & (ax67x) & (ax66x) & (!ax65x)) + ((!shiftx0x) & (!shiftx1x) & (ax64x) & (ax67x) & (ax66x) & (ax65x)) + ((!shiftx0x) & (shiftx1x) & (!ax64x) & (!ax67x) & (!ax66x) & (ax65x)) + ((!shiftx0x) & (shiftx1x) & (!ax64x) & (!ax67x) & (ax66x) & (ax65x)) + ((!shiftx0x) & (shiftx1x) & (!ax64x) & (ax67x) & (!ax66x) & (ax65x)) + ((!shiftx0x) & (shiftx1x) & (!ax64x) & (ax67x) & (ax66x) & (ax65x)) + ((!shiftx0x) & (shiftx1x) & (ax64x) & (!ax67x) & (!ax66x) & (ax65x)) + ((!shiftx0x) & (shiftx1x) & (ax64x) & (!ax67x) & (ax66x) & (ax65x)) + ((!shiftx0x) & (shiftx1x) & (ax64x) & (ax67x) & (!ax66x) & (ax65x)) + ((!shiftx0x) & (shiftx1x) & (ax64x) & (ax67x) & (ax66x) & (ax65x)) + ((shiftx0x) & (!shiftx1x) & (!ax64x) & (!ax67x) & (ax66x) & (!ax65x)) + ((shiftx0x) & (!shiftx1x) & (!ax64x) & (!ax67x) & (ax66x) & (ax65x)) + ((shiftx0x) & (!shiftx1x) & (!ax64x) & (ax67x) & (ax66x) & (!ax65x)) + ((shiftx0x) & (!shiftx1x) & (!ax64x) & (ax67x) & (ax66x) & (ax65x)) + ((shiftx0x) & (!shiftx1x) & (ax64x) & (!ax67x) & (ax66x) & (!ax65x)) + ((shiftx0x) & (!shiftx1x) & (ax64x) & (!ax67x) & (ax66x) & (ax65x)) + ((shiftx0x) & (!shiftx1x) & (ax64x) & (ax67x) & (ax66x) & (!ax65x)) + ((shiftx0x) & (!shiftx1x) & (ax64x) & (ax67x) & (ax66x) & (ax65x)) + ((shiftx0x) & (shiftx1x) & (ax64x) & (!ax67x) & (!ax66x) & (!ax65x)) + ((shiftx0x) & (shiftx1x) & (ax64x) & (!ax67x) & (!ax66x) & (ax65x)) + ((shiftx0x) & (shiftx1x) & (ax64x) & (!ax67x) & (ax66x) & (!ax65x)) + ((shiftx0x) & (shiftx1x) & (ax64x) & (!ax67x) & (ax66x) & (ax65x)) + ((shiftx0x) & (shiftx1x) & (ax64x) & (ax67x) & (!ax66x) & (!ax65x)) + ((shiftx0x) & (shiftx1x) & (ax64x) & (ax67x) & (!ax66x) & (ax65x)) + ((shiftx0x) & (shiftx1x) & (ax64x) & (ax67x) & (ax66x) & (!ax65x)) + ((shiftx0x) & (shiftx1x) & (ax64x) & (ax67x) & (ax66x) & (ax65x)));
	assign g131 = (((!shiftx0x) & (!shiftx1x) & (ax63x) & (!ax62x) & (!ax61x) & (!ax60x)) + ((!shiftx0x) & (!shiftx1x) & (ax63x) & (!ax62x) & (!ax61x) & (ax60x)) + ((!shiftx0x) & (!shiftx1x) & (ax63x) & (!ax62x) & (ax61x) & (!ax60x)) + ((!shiftx0x) & (!shiftx1x) & (ax63x) & (!ax62x) & (ax61x) & (ax60x)) + ((!shiftx0x) & (!shiftx1x) & (ax63x) & (ax62x) & (!ax61x) & (!ax60x)) + ((!shiftx0x) & (!shiftx1x) & (ax63x) & (ax62x) & (!ax61x) & (ax60x)) + ((!shiftx0x) & (!shiftx1x) & (ax63x) & (ax62x) & (ax61x) & (!ax60x)) + ((!shiftx0x) & (!shiftx1x) & (ax63x) & (ax62x) & (ax61x) & (ax60x)) + ((!shiftx0x) & (shiftx1x) & (!ax63x) & (!ax62x) & (ax61x) & (!ax60x)) + ((!shiftx0x) & (shiftx1x) & (!ax63x) & (!ax62x) & (ax61x) & (ax60x)) + ((!shiftx0x) & (shiftx1x) & (!ax63x) & (ax62x) & (ax61x) & (!ax60x)) + ((!shiftx0x) & (shiftx1x) & (!ax63x) & (ax62x) & (ax61x) & (ax60x)) + ((!shiftx0x) & (shiftx1x) & (ax63x) & (!ax62x) & (ax61x) & (!ax60x)) + ((!shiftx0x) & (shiftx1x) & (ax63x) & (!ax62x) & (ax61x) & (ax60x)) + ((!shiftx0x) & (shiftx1x) & (ax63x) & (ax62x) & (ax61x) & (!ax60x)) + ((!shiftx0x) & (shiftx1x) & (ax63x) & (ax62x) & (ax61x) & (ax60x)) + ((shiftx0x) & (!shiftx1x) & (!ax63x) & (ax62x) & (!ax61x) & (!ax60x)) + ((shiftx0x) & (!shiftx1x) & (!ax63x) & (ax62x) & (!ax61x) & (ax60x)) + ((shiftx0x) & (!shiftx1x) & (!ax63x) & (ax62x) & (ax61x) & (!ax60x)) + ((shiftx0x) & (!shiftx1x) & (!ax63x) & (ax62x) & (ax61x) & (ax60x)) + ((shiftx0x) & (!shiftx1x) & (ax63x) & (ax62x) & (!ax61x) & (!ax60x)) + ((shiftx0x) & (!shiftx1x) & (ax63x) & (ax62x) & (!ax61x) & (ax60x)) + ((shiftx0x) & (!shiftx1x) & (ax63x) & (ax62x) & (ax61x) & (!ax60x)) + ((shiftx0x) & (!shiftx1x) & (ax63x) & (ax62x) & (ax61x) & (ax60x)) + ((shiftx0x) & (shiftx1x) & (!ax63x) & (!ax62x) & (!ax61x) & (ax60x)) + ((shiftx0x) & (shiftx1x) & (!ax63x) & (!ax62x) & (ax61x) & (ax60x)) + ((shiftx0x) & (shiftx1x) & (!ax63x) & (ax62x) & (!ax61x) & (ax60x)) + ((shiftx0x) & (shiftx1x) & (!ax63x) & (ax62x) & (ax61x) & (ax60x)) + ((shiftx0x) & (shiftx1x) & (ax63x) & (!ax62x) & (!ax61x) & (ax60x)) + ((shiftx0x) & (shiftx1x) & (ax63x) & (!ax62x) & (ax61x) & (ax60x)) + ((shiftx0x) & (shiftx1x) & (ax63x) & (ax62x) & (!ax61x) & (ax60x)) + ((shiftx0x) & (shiftx1x) & (ax63x) & (ax62x) & (ax61x) & (ax60x)));
	assign g132 = (((!shiftx0x) & (!shiftx1x) & (!ax52x) & (ax55x) & (!ax54x) & (!ax53x)) + ((!shiftx0x) & (!shiftx1x) & (!ax52x) & (ax55x) & (!ax54x) & (ax53x)) + ((!shiftx0x) & (!shiftx1x) & (!ax52x) & (ax55x) & (ax54x) & (!ax53x)) + ((!shiftx0x) & (!shiftx1x) & (!ax52x) & (ax55x) & (ax54x) & (ax53x)) + ((!shiftx0x) & (!shiftx1x) & (ax52x) & (ax55x) & (!ax54x) & (!ax53x)) + ((!shiftx0x) & (!shiftx1x) & (ax52x) & (ax55x) & (!ax54x) & (ax53x)) + ((!shiftx0x) & (!shiftx1x) & (ax52x) & (ax55x) & (ax54x) & (!ax53x)) + ((!shiftx0x) & (!shiftx1x) & (ax52x) & (ax55x) & (ax54x) & (ax53x)) + ((!shiftx0x) & (shiftx1x) & (!ax52x) & (!ax55x) & (!ax54x) & (ax53x)) + ((!shiftx0x) & (shiftx1x) & (!ax52x) & (!ax55x) & (ax54x) & (ax53x)) + ((!shiftx0x) & (shiftx1x) & (!ax52x) & (ax55x) & (!ax54x) & (ax53x)) + ((!shiftx0x) & (shiftx1x) & (!ax52x) & (ax55x) & (ax54x) & (ax53x)) + ((!shiftx0x) & (shiftx1x) & (ax52x) & (!ax55x) & (!ax54x) & (ax53x)) + ((!shiftx0x) & (shiftx1x) & (ax52x) & (!ax55x) & (ax54x) & (ax53x)) + ((!shiftx0x) & (shiftx1x) & (ax52x) & (ax55x) & (!ax54x) & (ax53x)) + ((!shiftx0x) & (shiftx1x) & (ax52x) & (ax55x) & (ax54x) & (ax53x)) + ((shiftx0x) & (!shiftx1x) & (!ax52x) & (!ax55x) & (ax54x) & (!ax53x)) + ((shiftx0x) & (!shiftx1x) & (!ax52x) & (!ax55x) & (ax54x) & (ax53x)) + ((shiftx0x) & (!shiftx1x) & (!ax52x) & (ax55x) & (ax54x) & (!ax53x)) + ((shiftx0x) & (!shiftx1x) & (!ax52x) & (ax55x) & (ax54x) & (ax53x)) + ((shiftx0x) & (!shiftx1x) & (ax52x) & (!ax55x) & (ax54x) & (!ax53x)) + ((shiftx0x) & (!shiftx1x) & (ax52x) & (!ax55x) & (ax54x) & (ax53x)) + ((shiftx0x) & (!shiftx1x) & (ax52x) & (ax55x) & (ax54x) & (!ax53x)) + ((shiftx0x) & (!shiftx1x) & (ax52x) & (ax55x) & (ax54x) & (ax53x)) + ((shiftx0x) & (shiftx1x) & (ax52x) & (!ax55x) & (!ax54x) & (!ax53x)) + ((shiftx0x) & (shiftx1x) & (ax52x) & (!ax55x) & (!ax54x) & (ax53x)) + ((shiftx0x) & (shiftx1x) & (ax52x) & (!ax55x) & (ax54x) & (!ax53x)) + ((shiftx0x) & (shiftx1x) & (ax52x) & (!ax55x) & (ax54x) & (ax53x)) + ((shiftx0x) & (shiftx1x) & (ax52x) & (ax55x) & (!ax54x) & (!ax53x)) + ((shiftx0x) & (shiftx1x) & (ax52x) & (ax55x) & (!ax54x) & (ax53x)) + ((shiftx0x) & (shiftx1x) & (ax52x) & (ax55x) & (ax54x) & (!ax53x)) + ((shiftx0x) & (shiftx1x) & (ax52x) & (ax55x) & (ax54x) & (ax53x)));
	assign g133 = (((!shiftx0x) & (!shiftx1x) & (ax59x) & (!ax58x) & (!ax57x) & (!ax56x)) + ((!shiftx0x) & (!shiftx1x) & (ax59x) & (!ax58x) & (!ax57x) & (ax56x)) + ((!shiftx0x) & (!shiftx1x) & (ax59x) & (!ax58x) & (ax57x) & (!ax56x)) + ((!shiftx0x) & (!shiftx1x) & (ax59x) & (!ax58x) & (ax57x) & (ax56x)) + ((!shiftx0x) & (!shiftx1x) & (ax59x) & (ax58x) & (!ax57x) & (!ax56x)) + ((!shiftx0x) & (!shiftx1x) & (ax59x) & (ax58x) & (!ax57x) & (ax56x)) + ((!shiftx0x) & (!shiftx1x) & (ax59x) & (ax58x) & (ax57x) & (!ax56x)) + ((!shiftx0x) & (!shiftx1x) & (ax59x) & (ax58x) & (ax57x) & (ax56x)) + ((!shiftx0x) & (shiftx1x) & (!ax59x) & (!ax58x) & (ax57x) & (!ax56x)) + ((!shiftx0x) & (shiftx1x) & (!ax59x) & (!ax58x) & (ax57x) & (ax56x)) + ((!shiftx0x) & (shiftx1x) & (!ax59x) & (ax58x) & (ax57x) & (!ax56x)) + ((!shiftx0x) & (shiftx1x) & (!ax59x) & (ax58x) & (ax57x) & (ax56x)) + ((!shiftx0x) & (shiftx1x) & (ax59x) & (!ax58x) & (ax57x) & (!ax56x)) + ((!shiftx0x) & (shiftx1x) & (ax59x) & (!ax58x) & (ax57x) & (ax56x)) + ((!shiftx0x) & (shiftx1x) & (ax59x) & (ax58x) & (ax57x) & (!ax56x)) + ((!shiftx0x) & (shiftx1x) & (ax59x) & (ax58x) & (ax57x) & (ax56x)) + ((shiftx0x) & (!shiftx1x) & (!ax59x) & (ax58x) & (!ax57x) & (!ax56x)) + ((shiftx0x) & (!shiftx1x) & (!ax59x) & (ax58x) & (!ax57x) & (ax56x)) + ((shiftx0x) & (!shiftx1x) & (!ax59x) & (ax58x) & (ax57x) & (!ax56x)) + ((shiftx0x) & (!shiftx1x) & (!ax59x) & (ax58x) & (ax57x) & (ax56x)) + ((shiftx0x) & (!shiftx1x) & (ax59x) & (ax58x) & (!ax57x) & (!ax56x)) + ((shiftx0x) & (!shiftx1x) & (ax59x) & (ax58x) & (!ax57x) & (ax56x)) + ((shiftx0x) & (!shiftx1x) & (ax59x) & (ax58x) & (ax57x) & (!ax56x)) + ((shiftx0x) & (!shiftx1x) & (ax59x) & (ax58x) & (ax57x) & (ax56x)) + ((shiftx0x) & (shiftx1x) & (!ax59x) & (!ax58x) & (!ax57x) & (ax56x)) + ((shiftx0x) & (shiftx1x) & (!ax59x) & (!ax58x) & (ax57x) & (ax56x)) + ((shiftx0x) & (shiftx1x) & (!ax59x) & (ax58x) & (!ax57x) & (ax56x)) + ((shiftx0x) & (shiftx1x) & (!ax59x) & (ax58x) & (ax57x) & (ax56x)) + ((shiftx0x) & (shiftx1x) & (ax59x) & (!ax58x) & (!ax57x) & (ax56x)) + ((shiftx0x) & (shiftx1x) & (ax59x) & (!ax58x) & (ax57x) & (ax56x)) + ((shiftx0x) & (shiftx1x) & (ax59x) & (ax58x) & (!ax57x) & (ax56x)) + ((shiftx0x) & (shiftx1x) & (ax59x) & (ax58x) & (ax57x) & (ax56x)));
	assign g134 = (((!shiftx2x) & (!shiftx3x) & (g130) & (!g131) & (!g132) & (!g133)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (!g131) & (!g132) & (g133)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (!g131) & (g132) & (!g133)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (!g131) & (g132) & (g133)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (g131) & (!g132) & (!g133)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (g131) & (!g132) & (g133)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (g131) & (g132) & (!g133)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (g131) & (g132) & (g133)) + ((!shiftx2x) & (shiftx3x) & (!g130) & (!g131) & (!g132) & (g133)) + ((!shiftx2x) & (shiftx3x) & (!g130) & (!g131) & (g132) & (g133)) + ((!shiftx2x) & (shiftx3x) & (!g130) & (g131) & (!g132) & (g133)) + ((!shiftx2x) & (shiftx3x) & (!g130) & (g131) & (g132) & (g133)) + ((!shiftx2x) & (shiftx3x) & (g130) & (!g131) & (!g132) & (g133)) + ((!shiftx2x) & (shiftx3x) & (g130) & (!g131) & (g132) & (g133)) + ((!shiftx2x) & (shiftx3x) & (g130) & (g131) & (!g132) & (g133)) + ((!shiftx2x) & (shiftx3x) & (g130) & (g131) & (g132) & (g133)) + ((shiftx2x) & (!shiftx3x) & (!g130) & (g131) & (!g132) & (!g133)) + ((shiftx2x) & (!shiftx3x) & (!g130) & (g131) & (!g132) & (g133)) + ((shiftx2x) & (!shiftx3x) & (!g130) & (g131) & (g132) & (!g133)) + ((shiftx2x) & (!shiftx3x) & (!g130) & (g131) & (g132) & (g133)) + ((shiftx2x) & (!shiftx3x) & (g130) & (g131) & (!g132) & (!g133)) + ((shiftx2x) & (!shiftx3x) & (g130) & (g131) & (!g132) & (g133)) + ((shiftx2x) & (!shiftx3x) & (g130) & (g131) & (g132) & (!g133)) + ((shiftx2x) & (!shiftx3x) & (g130) & (g131) & (g132) & (g133)) + ((shiftx2x) & (shiftx3x) & (!g130) & (!g131) & (g132) & (!g133)) + ((shiftx2x) & (shiftx3x) & (!g130) & (!g131) & (g132) & (g133)) + ((shiftx2x) & (shiftx3x) & (!g130) & (g131) & (g132) & (!g133)) + ((shiftx2x) & (shiftx3x) & (!g130) & (g131) & (g132) & (g133)) + ((shiftx2x) & (shiftx3x) & (g130) & (!g131) & (g132) & (!g133)) + ((shiftx2x) & (shiftx3x) & (g130) & (!g131) & (g132) & (g133)) + ((shiftx2x) & (shiftx3x) & (g130) & (g131) & (g132) & (!g133)) + ((shiftx2x) & (shiftx3x) & (g130) & (g131) & (g132) & (g133)));
	assign g135 = (((!shiftx0x) & (!shiftx1x) & (ax51x) & (!ax50x) & (!ax49x) & (!ax48x)) + ((!shiftx0x) & (!shiftx1x) & (ax51x) & (!ax50x) & (!ax49x) & (ax48x)) + ((!shiftx0x) & (!shiftx1x) & (ax51x) & (!ax50x) & (ax49x) & (!ax48x)) + ((!shiftx0x) & (!shiftx1x) & (ax51x) & (!ax50x) & (ax49x) & (ax48x)) + ((!shiftx0x) & (!shiftx1x) & (ax51x) & (ax50x) & (!ax49x) & (!ax48x)) + ((!shiftx0x) & (!shiftx1x) & (ax51x) & (ax50x) & (!ax49x) & (ax48x)) + ((!shiftx0x) & (!shiftx1x) & (ax51x) & (ax50x) & (ax49x) & (!ax48x)) + ((!shiftx0x) & (!shiftx1x) & (ax51x) & (ax50x) & (ax49x) & (ax48x)) + ((!shiftx0x) & (shiftx1x) & (!ax51x) & (!ax50x) & (ax49x) & (!ax48x)) + ((!shiftx0x) & (shiftx1x) & (!ax51x) & (!ax50x) & (ax49x) & (ax48x)) + ((!shiftx0x) & (shiftx1x) & (!ax51x) & (ax50x) & (ax49x) & (!ax48x)) + ((!shiftx0x) & (shiftx1x) & (!ax51x) & (ax50x) & (ax49x) & (ax48x)) + ((!shiftx0x) & (shiftx1x) & (ax51x) & (!ax50x) & (ax49x) & (!ax48x)) + ((!shiftx0x) & (shiftx1x) & (ax51x) & (!ax50x) & (ax49x) & (ax48x)) + ((!shiftx0x) & (shiftx1x) & (ax51x) & (ax50x) & (ax49x) & (!ax48x)) + ((!shiftx0x) & (shiftx1x) & (ax51x) & (ax50x) & (ax49x) & (ax48x)) + ((shiftx0x) & (!shiftx1x) & (!ax51x) & (ax50x) & (!ax49x) & (!ax48x)) + ((shiftx0x) & (!shiftx1x) & (!ax51x) & (ax50x) & (!ax49x) & (ax48x)) + ((shiftx0x) & (!shiftx1x) & (!ax51x) & (ax50x) & (ax49x) & (!ax48x)) + ((shiftx0x) & (!shiftx1x) & (!ax51x) & (ax50x) & (ax49x) & (ax48x)) + ((shiftx0x) & (!shiftx1x) & (ax51x) & (ax50x) & (!ax49x) & (!ax48x)) + ((shiftx0x) & (!shiftx1x) & (ax51x) & (ax50x) & (!ax49x) & (ax48x)) + ((shiftx0x) & (!shiftx1x) & (ax51x) & (ax50x) & (ax49x) & (!ax48x)) + ((shiftx0x) & (!shiftx1x) & (ax51x) & (ax50x) & (ax49x) & (ax48x)) + ((shiftx0x) & (shiftx1x) & (!ax51x) & (!ax50x) & (!ax49x) & (ax48x)) + ((shiftx0x) & (shiftx1x) & (!ax51x) & (!ax50x) & (ax49x) & (ax48x)) + ((shiftx0x) & (shiftx1x) & (!ax51x) & (ax50x) & (!ax49x) & (ax48x)) + ((shiftx0x) & (shiftx1x) & (!ax51x) & (ax50x) & (ax49x) & (ax48x)) + ((shiftx0x) & (shiftx1x) & (ax51x) & (!ax50x) & (!ax49x) & (ax48x)) + ((shiftx0x) & (shiftx1x) & (ax51x) & (!ax50x) & (ax49x) & (ax48x)) + ((shiftx0x) & (shiftx1x) & (ax51x) & (ax50x) & (!ax49x) & (ax48x)) + ((shiftx0x) & (shiftx1x) & (ax51x) & (ax50x) & (ax49x) & (ax48x)));
	assign g136 = (((!ax47x) & (!ax46x) & (!ax45x) & (ax44x) & (shiftx0x) & (shiftx1x)) + ((!ax47x) & (!ax46x) & (ax45x) & (!ax44x) & (!shiftx0x) & (shiftx1x)) + ((!ax47x) & (!ax46x) & (ax45x) & (ax44x) & (!shiftx0x) & (shiftx1x)) + ((!ax47x) & (!ax46x) & (ax45x) & (ax44x) & (shiftx0x) & (shiftx1x)) + ((!ax47x) & (ax46x) & (!ax45x) & (!ax44x) & (shiftx0x) & (!shiftx1x)) + ((!ax47x) & (ax46x) & (!ax45x) & (ax44x) & (shiftx0x) & (!shiftx1x)) + ((!ax47x) & (ax46x) & (!ax45x) & (ax44x) & (shiftx0x) & (shiftx1x)) + ((!ax47x) & (ax46x) & (ax45x) & (!ax44x) & (!shiftx0x) & (shiftx1x)) + ((!ax47x) & (ax46x) & (ax45x) & (!ax44x) & (shiftx0x) & (!shiftx1x)) + ((!ax47x) & (ax46x) & (ax45x) & (ax44x) & (!shiftx0x) & (shiftx1x)) + ((!ax47x) & (ax46x) & (ax45x) & (ax44x) & (shiftx0x) & (!shiftx1x)) + ((!ax47x) & (ax46x) & (ax45x) & (ax44x) & (shiftx0x) & (shiftx1x)) + ((ax47x) & (!ax46x) & (!ax45x) & (!ax44x) & (!shiftx0x) & (!shiftx1x)) + ((ax47x) & (!ax46x) & (!ax45x) & (ax44x) & (!shiftx0x) & (!shiftx1x)) + ((ax47x) & (!ax46x) & (!ax45x) & (ax44x) & (shiftx0x) & (shiftx1x)) + ((ax47x) & (!ax46x) & (ax45x) & (!ax44x) & (!shiftx0x) & (!shiftx1x)) + ((ax47x) & (!ax46x) & (ax45x) & (!ax44x) & (!shiftx0x) & (shiftx1x)) + ((ax47x) & (!ax46x) & (ax45x) & (ax44x) & (!shiftx0x) & (!shiftx1x)) + ((ax47x) & (!ax46x) & (ax45x) & (ax44x) & (!shiftx0x) & (shiftx1x)) + ((ax47x) & (!ax46x) & (ax45x) & (ax44x) & (shiftx0x) & (shiftx1x)) + ((ax47x) & (ax46x) & (!ax45x) & (!ax44x) & (!shiftx0x) & (!shiftx1x)) + ((ax47x) & (ax46x) & (!ax45x) & (!ax44x) & (shiftx0x) & (!shiftx1x)) + ((ax47x) & (ax46x) & (!ax45x) & (ax44x) & (!shiftx0x) & (!shiftx1x)) + ((ax47x) & (ax46x) & (!ax45x) & (ax44x) & (shiftx0x) & (!shiftx1x)) + ((ax47x) & (ax46x) & (!ax45x) & (ax44x) & (shiftx0x) & (shiftx1x)) + ((ax47x) & (ax46x) & (ax45x) & (!ax44x) & (!shiftx0x) & (!shiftx1x)) + ((ax47x) & (ax46x) & (ax45x) & (!ax44x) & (!shiftx0x) & (shiftx1x)) + ((ax47x) & (ax46x) & (ax45x) & (!ax44x) & (shiftx0x) & (!shiftx1x)) + ((ax47x) & (ax46x) & (ax45x) & (ax44x) & (!shiftx0x) & (!shiftx1x)) + ((ax47x) & (ax46x) & (ax45x) & (ax44x) & (!shiftx0x) & (shiftx1x)) + ((ax47x) & (ax46x) & (ax45x) & (ax44x) & (shiftx0x) & (!shiftx1x)) + ((ax47x) & (ax46x) & (ax45x) & (ax44x) & (shiftx0x) & (shiftx1x)));
	assign g137 = (((!shiftx0x) & (!shiftx1x) & (!ax36x) & (!ax38x) & (ax39x) & (!ax37x)) + ((!shiftx0x) & (!shiftx1x) & (!ax36x) & (!ax38x) & (ax39x) & (ax37x)) + ((!shiftx0x) & (!shiftx1x) & (!ax36x) & (ax38x) & (ax39x) & (!ax37x)) + ((!shiftx0x) & (!shiftx1x) & (!ax36x) & (ax38x) & (ax39x) & (ax37x)) + ((!shiftx0x) & (!shiftx1x) & (ax36x) & (!ax38x) & (ax39x) & (!ax37x)) + ((!shiftx0x) & (!shiftx1x) & (ax36x) & (!ax38x) & (ax39x) & (ax37x)) + ((!shiftx0x) & (!shiftx1x) & (ax36x) & (ax38x) & (ax39x) & (!ax37x)) + ((!shiftx0x) & (!shiftx1x) & (ax36x) & (ax38x) & (ax39x) & (ax37x)) + ((!shiftx0x) & (shiftx1x) & (!ax36x) & (!ax38x) & (!ax39x) & (ax37x)) + ((!shiftx0x) & (shiftx1x) & (!ax36x) & (!ax38x) & (ax39x) & (ax37x)) + ((!shiftx0x) & (shiftx1x) & (!ax36x) & (ax38x) & (!ax39x) & (ax37x)) + ((!shiftx0x) & (shiftx1x) & (!ax36x) & (ax38x) & (ax39x) & (ax37x)) + ((!shiftx0x) & (shiftx1x) & (ax36x) & (!ax38x) & (!ax39x) & (ax37x)) + ((!shiftx0x) & (shiftx1x) & (ax36x) & (!ax38x) & (ax39x) & (ax37x)) + ((!shiftx0x) & (shiftx1x) & (ax36x) & (ax38x) & (!ax39x) & (ax37x)) + ((!shiftx0x) & (shiftx1x) & (ax36x) & (ax38x) & (ax39x) & (ax37x)) + ((shiftx0x) & (!shiftx1x) & (!ax36x) & (ax38x) & (!ax39x) & (!ax37x)) + ((shiftx0x) & (!shiftx1x) & (!ax36x) & (ax38x) & (!ax39x) & (ax37x)) + ((shiftx0x) & (!shiftx1x) & (!ax36x) & (ax38x) & (ax39x) & (!ax37x)) + ((shiftx0x) & (!shiftx1x) & (!ax36x) & (ax38x) & (ax39x) & (ax37x)) + ((shiftx0x) & (!shiftx1x) & (ax36x) & (ax38x) & (!ax39x) & (!ax37x)) + ((shiftx0x) & (!shiftx1x) & (ax36x) & (ax38x) & (!ax39x) & (ax37x)) + ((shiftx0x) & (!shiftx1x) & (ax36x) & (ax38x) & (ax39x) & (!ax37x)) + ((shiftx0x) & (!shiftx1x) & (ax36x) & (ax38x) & (ax39x) & (ax37x)) + ((shiftx0x) & (shiftx1x) & (ax36x) & (!ax38x) & (!ax39x) & (!ax37x)) + ((shiftx0x) & (shiftx1x) & (ax36x) & (!ax38x) & (!ax39x) & (ax37x)) + ((shiftx0x) & (shiftx1x) & (ax36x) & (!ax38x) & (ax39x) & (!ax37x)) + ((shiftx0x) & (shiftx1x) & (ax36x) & (!ax38x) & (ax39x) & (ax37x)) + ((shiftx0x) & (shiftx1x) & (ax36x) & (ax38x) & (!ax39x) & (!ax37x)) + ((shiftx0x) & (shiftx1x) & (ax36x) & (ax38x) & (!ax39x) & (ax37x)) + ((shiftx0x) & (shiftx1x) & (ax36x) & (ax38x) & (ax39x) & (!ax37x)) + ((shiftx0x) & (shiftx1x) & (ax36x) & (ax38x) & (ax39x) & (ax37x)));
	assign g138 = (((!ax43x) & (!ax41x) & (!ax42x) & (ax40x) & (shiftx1x) & (shiftx0x)) + ((!ax43x) & (!ax41x) & (ax42x) & (!ax40x) & (!shiftx1x) & (shiftx0x)) + ((!ax43x) & (!ax41x) & (ax42x) & (ax40x) & (!shiftx1x) & (shiftx0x)) + ((!ax43x) & (!ax41x) & (ax42x) & (ax40x) & (shiftx1x) & (shiftx0x)) + ((!ax43x) & (ax41x) & (!ax42x) & (!ax40x) & (shiftx1x) & (!shiftx0x)) + ((!ax43x) & (ax41x) & (!ax42x) & (ax40x) & (shiftx1x) & (!shiftx0x)) + ((!ax43x) & (ax41x) & (!ax42x) & (ax40x) & (shiftx1x) & (shiftx0x)) + ((!ax43x) & (ax41x) & (ax42x) & (!ax40x) & (!shiftx1x) & (shiftx0x)) + ((!ax43x) & (ax41x) & (ax42x) & (!ax40x) & (shiftx1x) & (!shiftx0x)) + ((!ax43x) & (ax41x) & (ax42x) & (ax40x) & (!shiftx1x) & (shiftx0x)) + ((!ax43x) & (ax41x) & (ax42x) & (ax40x) & (shiftx1x) & (!shiftx0x)) + ((!ax43x) & (ax41x) & (ax42x) & (ax40x) & (shiftx1x) & (shiftx0x)) + ((ax43x) & (!ax41x) & (!ax42x) & (!ax40x) & (!shiftx1x) & (!shiftx0x)) + ((ax43x) & (!ax41x) & (!ax42x) & (ax40x) & (!shiftx1x) & (!shiftx0x)) + ((ax43x) & (!ax41x) & (!ax42x) & (ax40x) & (shiftx1x) & (shiftx0x)) + ((ax43x) & (!ax41x) & (ax42x) & (!ax40x) & (!shiftx1x) & (!shiftx0x)) + ((ax43x) & (!ax41x) & (ax42x) & (!ax40x) & (!shiftx1x) & (shiftx0x)) + ((ax43x) & (!ax41x) & (ax42x) & (ax40x) & (!shiftx1x) & (!shiftx0x)) + ((ax43x) & (!ax41x) & (ax42x) & (ax40x) & (!shiftx1x) & (shiftx0x)) + ((ax43x) & (!ax41x) & (ax42x) & (ax40x) & (shiftx1x) & (shiftx0x)) + ((ax43x) & (ax41x) & (!ax42x) & (!ax40x) & (!shiftx1x) & (!shiftx0x)) + ((ax43x) & (ax41x) & (!ax42x) & (!ax40x) & (shiftx1x) & (!shiftx0x)) + ((ax43x) & (ax41x) & (!ax42x) & (ax40x) & (!shiftx1x) & (!shiftx0x)) + ((ax43x) & (ax41x) & (!ax42x) & (ax40x) & (shiftx1x) & (!shiftx0x)) + ((ax43x) & (ax41x) & (!ax42x) & (ax40x) & (shiftx1x) & (shiftx0x)) + ((ax43x) & (ax41x) & (ax42x) & (!ax40x) & (!shiftx1x) & (!shiftx0x)) + ((ax43x) & (ax41x) & (ax42x) & (!ax40x) & (!shiftx1x) & (shiftx0x)) + ((ax43x) & (ax41x) & (ax42x) & (!ax40x) & (shiftx1x) & (!shiftx0x)) + ((ax43x) & (ax41x) & (ax42x) & (ax40x) & (!shiftx1x) & (!shiftx0x)) + ((ax43x) & (ax41x) & (ax42x) & (ax40x) & (!shiftx1x) & (shiftx0x)) + ((ax43x) & (ax41x) & (ax42x) & (ax40x) & (shiftx1x) & (!shiftx0x)) + ((ax43x) & (ax41x) & (ax42x) & (ax40x) & (shiftx1x) & (shiftx0x)));
	assign g139 = (((!shiftx2x) & (!shiftx3x) & (g135) & (!g136) & (!g137) & (!g138)) + ((!shiftx2x) & (!shiftx3x) & (g135) & (!g136) & (!g137) & (g138)) + ((!shiftx2x) & (!shiftx3x) & (g135) & (!g136) & (g137) & (!g138)) + ((!shiftx2x) & (!shiftx3x) & (g135) & (!g136) & (g137) & (g138)) + ((!shiftx2x) & (!shiftx3x) & (g135) & (g136) & (!g137) & (!g138)) + ((!shiftx2x) & (!shiftx3x) & (g135) & (g136) & (!g137) & (g138)) + ((!shiftx2x) & (!shiftx3x) & (g135) & (g136) & (g137) & (!g138)) + ((!shiftx2x) & (!shiftx3x) & (g135) & (g136) & (g137) & (g138)) + ((!shiftx2x) & (shiftx3x) & (!g135) & (!g136) & (!g137) & (g138)) + ((!shiftx2x) & (shiftx3x) & (!g135) & (!g136) & (g137) & (g138)) + ((!shiftx2x) & (shiftx3x) & (!g135) & (g136) & (!g137) & (g138)) + ((!shiftx2x) & (shiftx3x) & (!g135) & (g136) & (g137) & (g138)) + ((!shiftx2x) & (shiftx3x) & (g135) & (!g136) & (!g137) & (g138)) + ((!shiftx2x) & (shiftx3x) & (g135) & (!g136) & (g137) & (g138)) + ((!shiftx2x) & (shiftx3x) & (g135) & (g136) & (!g137) & (g138)) + ((!shiftx2x) & (shiftx3x) & (g135) & (g136) & (g137) & (g138)) + ((shiftx2x) & (!shiftx3x) & (!g135) & (g136) & (!g137) & (!g138)) + ((shiftx2x) & (!shiftx3x) & (!g135) & (g136) & (!g137) & (g138)) + ((shiftx2x) & (!shiftx3x) & (!g135) & (g136) & (g137) & (!g138)) + ((shiftx2x) & (!shiftx3x) & (!g135) & (g136) & (g137) & (g138)) + ((shiftx2x) & (!shiftx3x) & (g135) & (g136) & (!g137) & (!g138)) + ((shiftx2x) & (!shiftx3x) & (g135) & (g136) & (!g137) & (g138)) + ((shiftx2x) & (!shiftx3x) & (g135) & (g136) & (g137) & (!g138)) + ((shiftx2x) & (!shiftx3x) & (g135) & (g136) & (g137) & (g138)) + ((shiftx2x) & (shiftx3x) & (!g135) & (!g136) & (g137) & (!g138)) + ((shiftx2x) & (shiftx3x) & (!g135) & (!g136) & (g137) & (g138)) + ((shiftx2x) & (shiftx3x) & (!g135) & (g136) & (g137) & (!g138)) + ((shiftx2x) & (shiftx3x) & (!g135) & (g136) & (g137) & (g138)) + ((shiftx2x) & (shiftx3x) & (g135) & (!g136) & (g137) & (!g138)) + ((shiftx2x) & (shiftx3x) & (g135) & (!g136) & (g137) & (g138)) + ((shiftx2x) & (shiftx3x) & (g135) & (g136) & (g137) & (!g138)) + ((shiftx2x) & (shiftx3x) & (g135) & (g136) & (g137) & (g138)));
	assign g140 = (((!ax16x) & (!shiftx0x) & (!shiftx1x) & (ax19x) & (!ax18x) & (!ax17x)) + ((!ax16x) & (!shiftx0x) & (!shiftx1x) & (ax19x) & (!ax18x) & (ax17x)) + ((!ax16x) & (!shiftx0x) & (!shiftx1x) & (ax19x) & (ax18x) & (!ax17x)) + ((!ax16x) & (!shiftx0x) & (!shiftx1x) & (ax19x) & (ax18x) & (ax17x)) + ((!ax16x) & (!shiftx0x) & (shiftx1x) & (!ax19x) & (!ax18x) & (ax17x)) + ((!ax16x) & (!shiftx0x) & (shiftx1x) & (!ax19x) & (ax18x) & (ax17x)) + ((!ax16x) & (!shiftx0x) & (shiftx1x) & (ax19x) & (!ax18x) & (ax17x)) + ((!ax16x) & (!shiftx0x) & (shiftx1x) & (ax19x) & (ax18x) & (ax17x)) + ((!ax16x) & (shiftx0x) & (!shiftx1x) & (!ax19x) & (ax18x) & (!ax17x)) + ((!ax16x) & (shiftx0x) & (!shiftx1x) & (!ax19x) & (ax18x) & (ax17x)) + ((!ax16x) & (shiftx0x) & (!shiftx1x) & (ax19x) & (ax18x) & (!ax17x)) + ((!ax16x) & (shiftx0x) & (!shiftx1x) & (ax19x) & (ax18x) & (ax17x)) + ((ax16x) & (!shiftx0x) & (!shiftx1x) & (ax19x) & (!ax18x) & (!ax17x)) + ((ax16x) & (!shiftx0x) & (!shiftx1x) & (ax19x) & (!ax18x) & (ax17x)) + ((ax16x) & (!shiftx0x) & (!shiftx1x) & (ax19x) & (ax18x) & (!ax17x)) + ((ax16x) & (!shiftx0x) & (!shiftx1x) & (ax19x) & (ax18x) & (ax17x)) + ((ax16x) & (!shiftx0x) & (shiftx1x) & (!ax19x) & (!ax18x) & (ax17x)) + ((ax16x) & (!shiftx0x) & (shiftx1x) & (!ax19x) & (ax18x) & (ax17x)) + ((ax16x) & (!shiftx0x) & (shiftx1x) & (ax19x) & (!ax18x) & (ax17x)) + ((ax16x) & (!shiftx0x) & (shiftx1x) & (ax19x) & (ax18x) & (ax17x)) + ((ax16x) & (shiftx0x) & (!shiftx1x) & (!ax19x) & (ax18x) & (!ax17x)) + ((ax16x) & (shiftx0x) & (!shiftx1x) & (!ax19x) & (ax18x) & (ax17x)) + ((ax16x) & (shiftx0x) & (!shiftx1x) & (ax19x) & (ax18x) & (!ax17x)) + ((ax16x) & (shiftx0x) & (!shiftx1x) & (ax19x) & (ax18x) & (ax17x)) + ((ax16x) & (shiftx0x) & (shiftx1x) & (!ax19x) & (!ax18x) & (!ax17x)) + ((ax16x) & (shiftx0x) & (shiftx1x) & (!ax19x) & (!ax18x) & (ax17x)) + ((ax16x) & (shiftx0x) & (shiftx1x) & (!ax19x) & (ax18x) & (!ax17x)) + ((ax16x) & (shiftx0x) & (shiftx1x) & (!ax19x) & (ax18x) & (ax17x)) + ((ax16x) & (shiftx0x) & (shiftx1x) & (ax19x) & (!ax18x) & (!ax17x)) + ((ax16x) & (shiftx0x) & (shiftx1x) & (ax19x) & (!ax18x) & (ax17x)) + ((ax16x) & (shiftx0x) & (shiftx1x) & (ax19x) & (ax18x) & (!ax17x)) + ((ax16x) & (shiftx0x) & (shiftx1x) & (ax19x) & (ax18x) & (ax17x)));
	assign g141 = (((!ax15x) & (!ax14x) & (!ax13x) & (shiftx0x) & (shiftx1x) & (ax12x)) + ((!ax15x) & (!ax14x) & (ax13x) & (!shiftx0x) & (shiftx1x) & (!ax12x)) + ((!ax15x) & (!ax14x) & (ax13x) & (!shiftx0x) & (shiftx1x) & (ax12x)) + ((!ax15x) & (!ax14x) & (ax13x) & (shiftx0x) & (shiftx1x) & (ax12x)) + ((!ax15x) & (ax14x) & (!ax13x) & (shiftx0x) & (!shiftx1x) & (!ax12x)) + ((!ax15x) & (ax14x) & (!ax13x) & (shiftx0x) & (!shiftx1x) & (ax12x)) + ((!ax15x) & (ax14x) & (!ax13x) & (shiftx0x) & (shiftx1x) & (ax12x)) + ((!ax15x) & (ax14x) & (ax13x) & (!shiftx0x) & (shiftx1x) & (!ax12x)) + ((!ax15x) & (ax14x) & (ax13x) & (!shiftx0x) & (shiftx1x) & (ax12x)) + ((!ax15x) & (ax14x) & (ax13x) & (shiftx0x) & (!shiftx1x) & (!ax12x)) + ((!ax15x) & (ax14x) & (ax13x) & (shiftx0x) & (!shiftx1x) & (ax12x)) + ((!ax15x) & (ax14x) & (ax13x) & (shiftx0x) & (shiftx1x) & (ax12x)) + ((ax15x) & (!ax14x) & (!ax13x) & (!shiftx0x) & (!shiftx1x) & (!ax12x)) + ((ax15x) & (!ax14x) & (!ax13x) & (!shiftx0x) & (!shiftx1x) & (ax12x)) + ((ax15x) & (!ax14x) & (!ax13x) & (shiftx0x) & (shiftx1x) & (ax12x)) + ((ax15x) & (!ax14x) & (ax13x) & (!shiftx0x) & (!shiftx1x) & (!ax12x)) + ((ax15x) & (!ax14x) & (ax13x) & (!shiftx0x) & (!shiftx1x) & (ax12x)) + ((ax15x) & (!ax14x) & (ax13x) & (!shiftx0x) & (shiftx1x) & (!ax12x)) + ((ax15x) & (!ax14x) & (ax13x) & (!shiftx0x) & (shiftx1x) & (ax12x)) + ((ax15x) & (!ax14x) & (ax13x) & (shiftx0x) & (shiftx1x) & (ax12x)) + ((ax15x) & (ax14x) & (!ax13x) & (!shiftx0x) & (!shiftx1x) & (!ax12x)) + ((ax15x) & (ax14x) & (!ax13x) & (!shiftx0x) & (!shiftx1x) & (ax12x)) + ((ax15x) & (ax14x) & (!ax13x) & (shiftx0x) & (!shiftx1x) & (!ax12x)) + ((ax15x) & (ax14x) & (!ax13x) & (shiftx0x) & (!shiftx1x) & (ax12x)) + ((ax15x) & (ax14x) & (!ax13x) & (shiftx0x) & (shiftx1x) & (ax12x)) + ((ax15x) & (ax14x) & (ax13x) & (!shiftx0x) & (!shiftx1x) & (!ax12x)) + ((ax15x) & (ax14x) & (ax13x) & (!shiftx0x) & (!shiftx1x) & (ax12x)) + ((ax15x) & (ax14x) & (ax13x) & (!shiftx0x) & (shiftx1x) & (!ax12x)) + ((ax15x) & (ax14x) & (ax13x) & (!shiftx0x) & (shiftx1x) & (ax12x)) + ((ax15x) & (ax14x) & (ax13x) & (shiftx0x) & (!shiftx1x) & (!ax12x)) + ((ax15x) & (ax14x) & (ax13x) & (shiftx0x) & (!shiftx1x) & (ax12x)) + ((ax15x) & (ax14x) & (ax13x) & (shiftx0x) & (shiftx1x) & (ax12x)));
	assign g142 = (((!shiftx0x) & (!shiftx1x) & (!ax4x) & (ax7x) & (!ax6x) & (!ax5x)) + ((!shiftx0x) & (!shiftx1x) & (!ax4x) & (ax7x) & (!ax6x) & (ax5x)) + ((!shiftx0x) & (!shiftx1x) & (!ax4x) & (ax7x) & (ax6x) & (!ax5x)) + ((!shiftx0x) & (!shiftx1x) & (!ax4x) & (ax7x) & (ax6x) & (ax5x)) + ((!shiftx0x) & (!shiftx1x) & (ax4x) & (ax7x) & (!ax6x) & (!ax5x)) + ((!shiftx0x) & (!shiftx1x) & (ax4x) & (ax7x) & (!ax6x) & (ax5x)) + ((!shiftx0x) & (!shiftx1x) & (ax4x) & (ax7x) & (ax6x) & (!ax5x)) + ((!shiftx0x) & (!shiftx1x) & (ax4x) & (ax7x) & (ax6x) & (ax5x)) + ((!shiftx0x) & (shiftx1x) & (!ax4x) & (!ax7x) & (!ax6x) & (ax5x)) + ((!shiftx0x) & (shiftx1x) & (!ax4x) & (!ax7x) & (ax6x) & (ax5x)) + ((!shiftx0x) & (shiftx1x) & (!ax4x) & (ax7x) & (!ax6x) & (ax5x)) + ((!shiftx0x) & (shiftx1x) & (!ax4x) & (ax7x) & (ax6x) & (ax5x)) + ((!shiftx0x) & (shiftx1x) & (ax4x) & (!ax7x) & (!ax6x) & (ax5x)) + ((!shiftx0x) & (shiftx1x) & (ax4x) & (!ax7x) & (ax6x) & (ax5x)) + ((!shiftx0x) & (shiftx1x) & (ax4x) & (ax7x) & (!ax6x) & (ax5x)) + ((!shiftx0x) & (shiftx1x) & (ax4x) & (ax7x) & (ax6x) & (ax5x)) + ((shiftx0x) & (!shiftx1x) & (!ax4x) & (!ax7x) & (ax6x) & (!ax5x)) + ((shiftx0x) & (!shiftx1x) & (!ax4x) & (!ax7x) & (ax6x) & (ax5x)) + ((shiftx0x) & (!shiftx1x) & (!ax4x) & (ax7x) & (ax6x) & (!ax5x)) + ((shiftx0x) & (!shiftx1x) & (!ax4x) & (ax7x) & (ax6x) & (ax5x)) + ((shiftx0x) & (!shiftx1x) & (ax4x) & (!ax7x) & (ax6x) & (!ax5x)) + ((shiftx0x) & (!shiftx1x) & (ax4x) & (!ax7x) & (ax6x) & (ax5x)) + ((shiftx0x) & (!shiftx1x) & (ax4x) & (ax7x) & (ax6x) & (!ax5x)) + ((shiftx0x) & (!shiftx1x) & (ax4x) & (ax7x) & (ax6x) & (ax5x)) + ((shiftx0x) & (shiftx1x) & (ax4x) & (!ax7x) & (!ax6x) & (!ax5x)) + ((shiftx0x) & (shiftx1x) & (ax4x) & (!ax7x) & (!ax6x) & (ax5x)) + ((shiftx0x) & (shiftx1x) & (ax4x) & (!ax7x) & (ax6x) & (!ax5x)) + ((shiftx0x) & (shiftx1x) & (ax4x) & (!ax7x) & (ax6x) & (ax5x)) + ((shiftx0x) & (shiftx1x) & (ax4x) & (ax7x) & (!ax6x) & (!ax5x)) + ((shiftx0x) & (shiftx1x) & (ax4x) & (ax7x) & (!ax6x) & (ax5x)) + ((shiftx0x) & (shiftx1x) & (ax4x) & (ax7x) & (ax6x) & (!ax5x)) + ((shiftx0x) & (shiftx1x) & (ax4x) & (ax7x) & (ax6x) & (ax5x)));
	assign g143 = (((!shiftx0x) & (!shiftx1x) & (ax11x) & (!ax10x) & (!ax9x) & (!ax8x)) + ((!shiftx0x) & (!shiftx1x) & (ax11x) & (!ax10x) & (!ax9x) & (ax8x)) + ((!shiftx0x) & (!shiftx1x) & (ax11x) & (!ax10x) & (ax9x) & (!ax8x)) + ((!shiftx0x) & (!shiftx1x) & (ax11x) & (!ax10x) & (ax9x) & (ax8x)) + ((!shiftx0x) & (!shiftx1x) & (ax11x) & (ax10x) & (!ax9x) & (!ax8x)) + ((!shiftx0x) & (!shiftx1x) & (ax11x) & (ax10x) & (!ax9x) & (ax8x)) + ((!shiftx0x) & (!shiftx1x) & (ax11x) & (ax10x) & (ax9x) & (!ax8x)) + ((!shiftx0x) & (!shiftx1x) & (ax11x) & (ax10x) & (ax9x) & (ax8x)) + ((!shiftx0x) & (shiftx1x) & (!ax11x) & (!ax10x) & (ax9x) & (!ax8x)) + ((!shiftx0x) & (shiftx1x) & (!ax11x) & (!ax10x) & (ax9x) & (ax8x)) + ((!shiftx0x) & (shiftx1x) & (!ax11x) & (ax10x) & (ax9x) & (!ax8x)) + ((!shiftx0x) & (shiftx1x) & (!ax11x) & (ax10x) & (ax9x) & (ax8x)) + ((!shiftx0x) & (shiftx1x) & (ax11x) & (!ax10x) & (ax9x) & (!ax8x)) + ((!shiftx0x) & (shiftx1x) & (ax11x) & (!ax10x) & (ax9x) & (ax8x)) + ((!shiftx0x) & (shiftx1x) & (ax11x) & (ax10x) & (ax9x) & (!ax8x)) + ((!shiftx0x) & (shiftx1x) & (ax11x) & (ax10x) & (ax9x) & (ax8x)) + ((shiftx0x) & (!shiftx1x) & (!ax11x) & (ax10x) & (!ax9x) & (!ax8x)) + ((shiftx0x) & (!shiftx1x) & (!ax11x) & (ax10x) & (!ax9x) & (ax8x)) + ((shiftx0x) & (!shiftx1x) & (!ax11x) & (ax10x) & (ax9x) & (!ax8x)) + ((shiftx0x) & (!shiftx1x) & (!ax11x) & (ax10x) & (ax9x) & (ax8x)) + ((shiftx0x) & (!shiftx1x) & (ax11x) & (ax10x) & (!ax9x) & (!ax8x)) + ((shiftx0x) & (!shiftx1x) & (ax11x) & (ax10x) & (!ax9x) & (ax8x)) + ((shiftx0x) & (!shiftx1x) & (ax11x) & (ax10x) & (ax9x) & (!ax8x)) + ((shiftx0x) & (!shiftx1x) & (ax11x) & (ax10x) & (ax9x) & (ax8x)) + ((shiftx0x) & (shiftx1x) & (!ax11x) & (!ax10x) & (!ax9x) & (ax8x)) + ((shiftx0x) & (shiftx1x) & (!ax11x) & (!ax10x) & (ax9x) & (ax8x)) + ((shiftx0x) & (shiftx1x) & (!ax11x) & (ax10x) & (!ax9x) & (ax8x)) + ((shiftx0x) & (shiftx1x) & (!ax11x) & (ax10x) & (ax9x) & (ax8x)) + ((shiftx0x) & (shiftx1x) & (ax11x) & (!ax10x) & (!ax9x) & (ax8x)) + ((shiftx0x) & (shiftx1x) & (ax11x) & (!ax10x) & (ax9x) & (ax8x)) + ((shiftx0x) & (shiftx1x) & (ax11x) & (ax10x) & (!ax9x) & (ax8x)) + ((shiftx0x) & (shiftx1x) & (ax11x) & (ax10x) & (ax9x) & (ax8x)));
	assign g144 = (((!shiftx2x) & (!shiftx3x) & (g140) & (!g141) & (!g142) & (!g143)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (!g141) & (!g142) & (g143)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (!g141) & (g142) & (!g143)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (!g141) & (g142) & (g143)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (g141) & (!g142) & (!g143)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (g141) & (!g142) & (g143)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (g141) & (g142) & (!g143)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (g141) & (g142) & (g143)) + ((!shiftx2x) & (shiftx3x) & (!g140) & (!g141) & (!g142) & (g143)) + ((!shiftx2x) & (shiftx3x) & (!g140) & (!g141) & (g142) & (g143)) + ((!shiftx2x) & (shiftx3x) & (!g140) & (g141) & (!g142) & (g143)) + ((!shiftx2x) & (shiftx3x) & (!g140) & (g141) & (g142) & (g143)) + ((!shiftx2x) & (shiftx3x) & (g140) & (!g141) & (!g142) & (g143)) + ((!shiftx2x) & (shiftx3x) & (g140) & (!g141) & (g142) & (g143)) + ((!shiftx2x) & (shiftx3x) & (g140) & (g141) & (!g142) & (g143)) + ((!shiftx2x) & (shiftx3x) & (g140) & (g141) & (g142) & (g143)) + ((shiftx2x) & (!shiftx3x) & (!g140) & (g141) & (!g142) & (!g143)) + ((shiftx2x) & (!shiftx3x) & (!g140) & (g141) & (!g142) & (g143)) + ((shiftx2x) & (!shiftx3x) & (!g140) & (g141) & (g142) & (!g143)) + ((shiftx2x) & (!shiftx3x) & (!g140) & (g141) & (g142) & (g143)) + ((shiftx2x) & (!shiftx3x) & (g140) & (g141) & (!g142) & (!g143)) + ((shiftx2x) & (!shiftx3x) & (g140) & (g141) & (!g142) & (g143)) + ((shiftx2x) & (!shiftx3x) & (g140) & (g141) & (g142) & (!g143)) + ((shiftx2x) & (!shiftx3x) & (g140) & (g141) & (g142) & (g143)) + ((shiftx2x) & (shiftx3x) & (!g140) & (!g141) & (g142) & (!g143)) + ((shiftx2x) & (shiftx3x) & (!g140) & (!g141) & (g142) & (g143)) + ((shiftx2x) & (shiftx3x) & (!g140) & (g141) & (g142) & (!g143)) + ((shiftx2x) & (shiftx3x) & (!g140) & (g141) & (g142) & (g143)) + ((shiftx2x) & (shiftx3x) & (g140) & (!g141) & (g142) & (!g143)) + ((shiftx2x) & (shiftx3x) & (g140) & (!g141) & (g142) & (g143)) + ((shiftx2x) & (shiftx3x) & (g140) & (g141) & (g142) & (!g143)) + ((shiftx2x) & (shiftx3x) & (g140) & (g141) & (g142) & (g143)));
	assign g145 = (((!shiftx0x) & (!shiftx1x) & (!ax32x) & (ax35x) & (!ax34x) & (!ax33x)) + ((!shiftx0x) & (!shiftx1x) & (!ax32x) & (ax35x) & (!ax34x) & (ax33x)) + ((!shiftx0x) & (!shiftx1x) & (!ax32x) & (ax35x) & (ax34x) & (!ax33x)) + ((!shiftx0x) & (!shiftx1x) & (!ax32x) & (ax35x) & (ax34x) & (ax33x)) + ((!shiftx0x) & (!shiftx1x) & (ax32x) & (ax35x) & (!ax34x) & (!ax33x)) + ((!shiftx0x) & (!shiftx1x) & (ax32x) & (ax35x) & (!ax34x) & (ax33x)) + ((!shiftx0x) & (!shiftx1x) & (ax32x) & (ax35x) & (ax34x) & (!ax33x)) + ((!shiftx0x) & (!shiftx1x) & (ax32x) & (ax35x) & (ax34x) & (ax33x)) + ((!shiftx0x) & (shiftx1x) & (!ax32x) & (!ax35x) & (!ax34x) & (ax33x)) + ((!shiftx0x) & (shiftx1x) & (!ax32x) & (!ax35x) & (ax34x) & (ax33x)) + ((!shiftx0x) & (shiftx1x) & (!ax32x) & (ax35x) & (!ax34x) & (ax33x)) + ((!shiftx0x) & (shiftx1x) & (!ax32x) & (ax35x) & (ax34x) & (ax33x)) + ((!shiftx0x) & (shiftx1x) & (ax32x) & (!ax35x) & (!ax34x) & (ax33x)) + ((!shiftx0x) & (shiftx1x) & (ax32x) & (!ax35x) & (ax34x) & (ax33x)) + ((!shiftx0x) & (shiftx1x) & (ax32x) & (ax35x) & (!ax34x) & (ax33x)) + ((!shiftx0x) & (shiftx1x) & (ax32x) & (ax35x) & (ax34x) & (ax33x)) + ((shiftx0x) & (!shiftx1x) & (!ax32x) & (!ax35x) & (ax34x) & (!ax33x)) + ((shiftx0x) & (!shiftx1x) & (!ax32x) & (!ax35x) & (ax34x) & (ax33x)) + ((shiftx0x) & (!shiftx1x) & (!ax32x) & (ax35x) & (ax34x) & (!ax33x)) + ((shiftx0x) & (!shiftx1x) & (!ax32x) & (ax35x) & (ax34x) & (ax33x)) + ((shiftx0x) & (!shiftx1x) & (ax32x) & (!ax35x) & (ax34x) & (!ax33x)) + ((shiftx0x) & (!shiftx1x) & (ax32x) & (!ax35x) & (ax34x) & (ax33x)) + ((shiftx0x) & (!shiftx1x) & (ax32x) & (ax35x) & (ax34x) & (!ax33x)) + ((shiftx0x) & (!shiftx1x) & (ax32x) & (ax35x) & (ax34x) & (ax33x)) + ((shiftx0x) & (shiftx1x) & (ax32x) & (!ax35x) & (!ax34x) & (!ax33x)) + ((shiftx0x) & (shiftx1x) & (ax32x) & (!ax35x) & (!ax34x) & (ax33x)) + ((shiftx0x) & (shiftx1x) & (ax32x) & (!ax35x) & (ax34x) & (!ax33x)) + ((shiftx0x) & (shiftx1x) & (ax32x) & (!ax35x) & (ax34x) & (ax33x)) + ((shiftx0x) & (shiftx1x) & (ax32x) & (ax35x) & (!ax34x) & (!ax33x)) + ((shiftx0x) & (shiftx1x) & (ax32x) & (ax35x) & (!ax34x) & (ax33x)) + ((shiftx0x) & (shiftx1x) & (ax32x) & (ax35x) & (ax34x) & (!ax33x)) + ((shiftx0x) & (shiftx1x) & (ax32x) & (ax35x) & (ax34x) & (ax33x)));
	assign g146 = (((!shiftx0x) & (!shiftx1x) & (ax31x) & (!ax30x) & (!ax29x) & (!ax28x)) + ((!shiftx0x) & (!shiftx1x) & (ax31x) & (!ax30x) & (!ax29x) & (ax28x)) + ((!shiftx0x) & (!shiftx1x) & (ax31x) & (!ax30x) & (ax29x) & (!ax28x)) + ((!shiftx0x) & (!shiftx1x) & (ax31x) & (!ax30x) & (ax29x) & (ax28x)) + ((!shiftx0x) & (!shiftx1x) & (ax31x) & (ax30x) & (!ax29x) & (!ax28x)) + ((!shiftx0x) & (!shiftx1x) & (ax31x) & (ax30x) & (!ax29x) & (ax28x)) + ((!shiftx0x) & (!shiftx1x) & (ax31x) & (ax30x) & (ax29x) & (!ax28x)) + ((!shiftx0x) & (!shiftx1x) & (ax31x) & (ax30x) & (ax29x) & (ax28x)) + ((!shiftx0x) & (shiftx1x) & (!ax31x) & (!ax30x) & (ax29x) & (!ax28x)) + ((!shiftx0x) & (shiftx1x) & (!ax31x) & (!ax30x) & (ax29x) & (ax28x)) + ((!shiftx0x) & (shiftx1x) & (!ax31x) & (ax30x) & (ax29x) & (!ax28x)) + ((!shiftx0x) & (shiftx1x) & (!ax31x) & (ax30x) & (ax29x) & (ax28x)) + ((!shiftx0x) & (shiftx1x) & (ax31x) & (!ax30x) & (ax29x) & (!ax28x)) + ((!shiftx0x) & (shiftx1x) & (ax31x) & (!ax30x) & (ax29x) & (ax28x)) + ((!shiftx0x) & (shiftx1x) & (ax31x) & (ax30x) & (ax29x) & (!ax28x)) + ((!shiftx0x) & (shiftx1x) & (ax31x) & (ax30x) & (ax29x) & (ax28x)) + ((shiftx0x) & (!shiftx1x) & (!ax31x) & (ax30x) & (!ax29x) & (!ax28x)) + ((shiftx0x) & (!shiftx1x) & (!ax31x) & (ax30x) & (!ax29x) & (ax28x)) + ((shiftx0x) & (!shiftx1x) & (!ax31x) & (ax30x) & (ax29x) & (!ax28x)) + ((shiftx0x) & (!shiftx1x) & (!ax31x) & (ax30x) & (ax29x) & (ax28x)) + ((shiftx0x) & (!shiftx1x) & (ax31x) & (ax30x) & (!ax29x) & (!ax28x)) + ((shiftx0x) & (!shiftx1x) & (ax31x) & (ax30x) & (!ax29x) & (ax28x)) + ((shiftx0x) & (!shiftx1x) & (ax31x) & (ax30x) & (ax29x) & (!ax28x)) + ((shiftx0x) & (!shiftx1x) & (ax31x) & (ax30x) & (ax29x) & (ax28x)) + ((shiftx0x) & (shiftx1x) & (!ax31x) & (!ax30x) & (!ax29x) & (ax28x)) + ((shiftx0x) & (shiftx1x) & (!ax31x) & (!ax30x) & (ax29x) & (ax28x)) + ((shiftx0x) & (shiftx1x) & (!ax31x) & (ax30x) & (!ax29x) & (ax28x)) + ((shiftx0x) & (shiftx1x) & (!ax31x) & (ax30x) & (ax29x) & (ax28x)) + ((shiftx0x) & (shiftx1x) & (ax31x) & (!ax30x) & (!ax29x) & (ax28x)) + ((shiftx0x) & (shiftx1x) & (ax31x) & (!ax30x) & (ax29x) & (ax28x)) + ((shiftx0x) & (shiftx1x) & (ax31x) & (ax30x) & (!ax29x) & (ax28x)) + ((shiftx0x) & (shiftx1x) & (ax31x) & (ax30x) & (ax29x) & (ax28x)));
	assign g147 = (((!shiftx0x) & (!shiftx1x) & (!ax20x) & (ax23x) & (!ax22x) & (!ax21x)) + ((!shiftx0x) & (!shiftx1x) & (!ax20x) & (ax23x) & (!ax22x) & (ax21x)) + ((!shiftx0x) & (!shiftx1x) & (!ax20x) & (ax23x) & (ax22x) & (!ax21x)) + ((!shiftx0x) & (!shiftx1x) & (!ax20x) & (ax23x) & (ax22x) & (ax21x)) + ((!shiftx0x) & (!shiftx1x) & (ax20x) & (ax23x) & (!ax22x) & (!ax21x)) + ((!shiftx0x) & (!shiftx1x) & (ax20x) & (ax23x) & (!ax22x) & (ax21x)) + ((!shiftx0x) & (!shiftx1x) & (ax20x) & (ax23x) & (ax22x) & (!ax21x)) + ((!shiftx0x) & (!shiftx1x) & (ax20x) & (ax23x) & (ax22x) & (ax21x)) + ((!shiftx0x) & (shiftx1x) & (!ax20x) & (!ax23x) & (!ax22x) & (ax21x)) + ((!shiftx0x) & (shiftx1x) & (!ax20x) & (!ax23x) & (ax22x) & (ax21x)) + ((!shiftx0x) & (shiftx1x) & (!ax20x) & (ax23x) & (!ax22x) & (ax21x)) + ((!shiftx0x) & (shiftx1x) & (!ax20x) & (ax23x) & (ax22x) & (ax21x)) + ((!shiftx0x) & (shiftx1x) & (ax20x) & (!ax23x) & (!ax22x) & (ax21x)) + ((!shiftx0x) & (shiftx1x) & (ax20x) & (!ax23x) & (ax22x) & (ax21x)) + ((!shiftx0x) & (shiftx1x) & (ax20x) & (ax23x) & (!ax22x) & (ax21x)) + ((!shiftx0x) & (shiftx1x) & (ax20x) & (ax23x) & (ax22x) & (ax21x)) + ((shiftx0x) & (!shiftx1x) & (!ax20x) & (!ax23x) & (ax22x) & (!ax21x)) + ((shiftx0x) & (!shiftx1x) & (!ax20x) & (!ax23x) & (ax22x) & (ax21x)) + ((shiftx0x) & (!shiftx1x) & (!ax20x) & (ax23x) & (ax22x) & (!ax21x)) + ((shiftx0x) & (!shiftx1x) & (!ax20x) & (ax23x) & (ax22x) & (ax21x)) + ((shiftx0x) & (!shiftx1x) & (ax20x) & (!ax23x) & (ax22x) & (!ax21x)) + ((shiftx0x) & (!shiftx1x) & (ax20x) & (!ax23x) & (ax22x) & (ax21x)) + ((shiftx0x) & (!shiftx1x) & (ax20x) & (ax23x) & (ax22x) & (!ax21x)) + ((shiftx0x) & (!shiftx1x) & (ax20x) & (ax23x) & (ax22x) & (ax21x)) + ((shiftx0x) & (shiftx1x) & (ax20x) & (!ax23x) & (!ax22x) & (!ax21x)) + ((shiftx0x) & (shiftx1x) & (ax20x) & (!ax23x) & (!ax22x) & (ax21x)) + ((shiftx0x) & (shiftx1x) & (ax20x) & (!ax23x) & (ax22x) & (!ax21x)) + ((shiftx0x) & (shiftx1x) & (ax20x) & (!ax23x) & (ax22x) & (ax21x)) + ((shiftx0x) & (shiftx1x) & (ax20x) & (ax23x) & (!ax22x) & (!ax21x)) + ((shiftx0x) & (shiftx1x) & (ax20x) & (ax23x) & (!ax22x) & (ax21x)) + ((shiftx0x) & (shiftx1x) & (ax20x) & (ax23x) & (ax22x) & (!ax21x)) + ((shiftx0x) & (shiftx1x) & (ax20x) & (ax23x) & (ax22x) & (ax21x)));
	assign g148 = (((!shiftx0x) & (!shiftx1x) & (ax27x) & (!ax26x) & (!ax25x) & (!ax24x)) + ((!shiftx0x) & (!shiftx1x) & (ax27x) & (!ax26x) & (!ax25x) & (ax24x)) + ((!shiftx0x) & (!shiftx1x) & (ax27x) & (!ax26x) & (ax25x) & (!ax24x)) + ((!shiftx0x) & (!shiftx1x) & (ax27x) & (!ax26x) & (ax25x) & (ax24x)) + ((!shiftx0x) & (!shiftx1x) & (ax27x) & (ax26x) & (!ax25x) & (!ax24x)) + ((!shiftx0x) & (!shiftx1x) & (ax27x) & (ax26x) & (!ax25x) & (ax24x)) + ((!shiftx0x) & (!shiftx1x) & (ax27x) & (ax26x) & (ax25x) & (!ax24x)) + ((!shiftx0x) & (!shiftx1x) & (ax27x) & (ax26x) & (ax25x) & (ax24x)) + ((!shiftx0x) & (shiftx1x) & (!ax27x) & (!ax26x) & (ax25x) & (!ax24x)) + ((!shiftx0x) & (shiftx1x) & (!ax27x) & (!ax26x) & (ax25x) & (ax24x)) + ((!shiftx0x) & (shiftx1x) & (!ax27x) & (ax26x) & (ax25x) & (!ax24x)) + ((!shiftx0x) & (shiftx1x) & (!ax27x) & (ax26x) & (ax25x) & (ax24x)) + ((!shiftx0x) & (shiftx1x) & (ax27x) & (!ax26x) & (ax25x) & (!ax24x)) + ((!shiftx0x) & (shiftx1x) & (ax27x) & (!ax26x) & (ax25x) & (ax24x)) + ((!shiftx0x) & (shiftx1x) & (ax27x) & (ax26x) & (ax25x) & (!ax24x)) + ((!shiftx0x) & (shiftx1x) & (ax27x) & (ax26x) & (ax25x) & (ax24x)) + ((shiftx0x) & (!shiftx1x) & (!ax27x) & (ax26x) & (!ax25x) & (!ax24x)) + ((shiftx0x) & (!shiftx1x) & (!ax27x) & (ax26x) & (!ax25x) & (ax24x)) + ((shiftx0x) & (!shiftx1x) & (!ax27x) & (ax26x) & (ax25x) & (!ax24x)) + ((shiftx0x) & (!shiftx1x) & (!ax27x) & (ax26x) & (ax25x) & (ax24x)) + ((shiftx0x) & (!shiftx1x) & (ax27x) & (ax26x) & (!ax25x) & (!ax24x)) + ((shiftx0x) & (!shiftx1x) & (ax27x) & (ax26x) & (!ax25x) & (ax24x)) + ((shiftx0x) & (!shiftx1x) & (ax27x) & (ax26x) & (ax25x) & (!ax24x)) + ((shiftx0x) & (!shiftx1x) & (ax27x) & (ax26x) & (ax25x) & (ax24x)) + ((shiftx0x) & (shiftx1x) & (!ax27x) & (!ax26x) & (!ax25x) & (ax24x)) + ((shiftx0x) & (shiftx1x) & (!ax27x) & (!ax26x) & (ax25x) & (ax24x)) + ((shiftx0x) & (shiftx1x) & (!ax27x) & (ax26x) & (!ax25x) & (ax24x)) + ((shiftx0x) & (shiftx1x) & (!ax27x) & (ax26x) & (ax25x) & (ax24x)) + ((shiftx0x) & (shiftx1x) & (ax27x) & (!ax26x) & (!ax25x) & (ax24x)) + ((shiftx0x) & (shiftx1x) & (ax27x) & (!ax26x) & (ax25x) & (ax24x)) + ((shiftx0x) & (shiftx1x) & (ax27x) & (ax26x) & (!ax25x) & (ax24x)) + ((shiftx0x) & (shiftx1x) & (ax27x) & (ax26x) & (ax25x) & (ax24x)));
	assign g149 = (((!shiftx2x) & (!shiftx3x) & (g145) & (!g146) & (!g147) & (!g148)) + ((!shiftx2x) & (!shiftx3x) & (g145) & (!g146) & (!g147) & (g148)) + ((!shiftx2x) & (!shiftx3x) & (g145) & (!g146) & (g147) & (!g148)) + ((!shiftx2x) & (!shiftx3x) & (g145) & (!g146) & (g147) & (g148)) + ((!shiftx2x) & (!shiftx3x) & (g145) & (g146) & (!g147) & (!g148)) + ((!shiftx2x) & (!shiftx3x) & (g145) & (g146) & (!g147) & (g148)) + ((!shiftx2x) & (!shiftx3x) & (g145) & (g146) & (g147) & (!g148)) + ((!shiftx2x) & (!shiftx3x) & (g145) & (g146) & (g147) & (g148)) + ((!shiftx2x) & (shiftx3x) & (!g145) & (!g146) & (!g147) & (g148)) + ((!shiftx2x) & (shiftx3x) & (!g145) & (!g146) & (g147) & (g148)) + ((!shiftx2x) & (shiftx3x) & (!g145) & (g146) & (!g147) & (g148)) + ((!shiftx2x) & (shiftx3x) & (!g145) & (g146) & (g147) & (g148)) + ((!shiftx2x) & (shiftx3x) & (g145) & (!g146) & (!g147) & (g148)) + ((!shiftx2x) & (shiftx3x) & (g145) & (!g146) & (g147) & (g148)) + ((!shiftx2x) & (shiftx3x) & (g145) & (g146) & (!g147) & (g148)) + ((!shiftx2x) & (shiftx3x) & (g145) & (g146) & (g147) & (g148)) + ((shiftx2x) & (!shiftx3x) & (!g145) & (g146) & (!g147) & (!g148)) + ((shiftx2x) & (!shiftx3x) & (!g145) & (g146) & (!g147) & (g148)) + ((shiftx2x) & (!shiftx3x) & (!g145) & (g146) & (g147) & (!g148)) + ((shiftx2x) & (!shiftx3x) & (!g145) & (g146) & (g147) & (g148)) + ((shiftx2x) & (!shiftx3x) & (g145) & (g146) & (!g147) & (!g148)) + ((shiftx2x) & (!shiftx3x) & (g145) & (g146) & (!g147) & (g148)) + ((shiftx2x) & (!shiftx3x) & (g145) & (g146) & (g147) & (!g148)) + ((shiftx2x) & (!shiftx3x) & (g145) & (g146) & (g147) & (g148)) + ((shiftx2x) & (shiftx3x) & (!g145) & (!g146) & (g147) & (!g148)) + ((shiftx2x) & (shiftx3x) & (!g145) & (!g146) & (g147) & (g148)) + ((shiftx2x) & (shiftx3x) & (!g145) & (g146) & (g147) & (!g148)) + ((shiftx2x) & (shiftx3x) & (!g145) & (g146) & (g147) & (g148)) + ((shiftx2x) & (shiftx3x) & (g145) & (!g146) & (g147) & (!g148)) + ((shiftx2x) & (shiftx3x) & (g145) & (!g146) & (g147) & (g148)) + ((shiftx2x) & (shiftx3x) & (g145) & (g146) & (g147) & (!g148)) + ((shiftx2x) & (shiftx3x) & (g145) & (g146) & (g147) & (g148)));
	assign g150 = (((!shiftx4x) & (!shiftx5x) & (g134) & (!g139) & (!g144) & (!g149)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (!g139) & (!g144) & (g149)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (!g139) & (g144) & (!g149)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (!g139) & (g144) & (g149)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (g139) & (!g144) & (!g149)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (g139) & (!g144) & (g149)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (g139) & (g144) & (!g149)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (g139) & (g144) & (g149)) + ((!shiftx4x) & (shiftx5x) & (!g134) & (!g139) & (!g144) & (g149)) + ((!shiftx4x) & (shiftx5x) & (!g134) & (!g139) & (g144) & (g149)) + ((!shiftx4x) & (shiftx5x) & (!g134) & (g139) & (!g144) & (g149)) + ((!shiftx4x) & (shiftx5x) & (!g134) & (g139) & (g144) & (g149)) + ((!shiftx4x) & (shiftx5x) & (g134) & (!g139) & (!g144) & (g149)) + ((!shiftx4x) & (shiftx5x) & (g134) & (!g139) & (g144) & (g149)) + ((!shiftx4x) & (shiftx5x) & (g134) & (g139) & (!g144) & (g149)) + ((!shiftx4x) & (shiftx5x) & (g134) & (g139) & (g144) & (g149)) + ((shiftx4x) & (!shiftx5x) & (!g134) & (g139) & (!g144) & (!g149)) + ((shiftx4x) & (!shiftx5x) & (!g134) & (g139) & (!g144) & (g149)) + ((shiftx4x) & (!shiftx5x) & (!g134) & (g139) & (g144) & (!g149)) + ((shiftx4x) & (!shiftx5x) & (!g134) & (g139) & (g144) & (g149)) + ((shiftx4x) & (!shiftx5x) & (g134) & (g139) & (!g144) & (!g149)) + ((shiftx4x) & (!shiftx5x) & (g134) & (g139) & (!g144) & (g149)) + ((shiftx4x) & (!shiftx5x) & (g134) & (g139) & (g144) & (!g149)) + ((shiftx4x) & (!shiftx5x) & (g134) & (g139) & (g144) & (g149)) + ((shiftx4x) & (shiftx5x) & (!g134) & (!g139) & (g144) & (!g149)) + ((shiftx4x) & (shiftx5x) & (!g134) & (!g139) & (g144) & (g149)) + ((shiftx4x) & (shiftx5x) & (!g134) & (g139) & (g144) & (!g149)) + ((shiftx4x) & (shiftx5x) & (!g134) & (g139) & (g144) & (g149)) + ((shiftx4x) & (shiftx5x) & (g134) & (!g139) & (g144) & (!g149)) + ((shiftx4x) & (shiftx5x) & (g134) & (!g139) & (g144) & (g149)) + ((shiftx4x) & (shiftx5x) & (g134) & (g139) & (g144) & (!g149)) + ((shiftx4x) & (shiftx5x) & (g134) & (g139) & (g144) & (g149)));
	assign g151 = (((!shiftx0x) & (!shiftx1x) & (ax115x) & (!ax114x) & (!ax113x) & (!ax112x)) + ((!shiftx0x) & (!shiftx1x) & (ax115x) & (!ax114x) & (!ax113x) & (ax112x)) + ((!shiftx0x) & (!shiftx1x) & (ax115x) & (!ax114x) & (ax113x) & (!ax112x)) + ((!shiftx0x) & (!shiftx1x) & (ax115x) & (!ax114x) & (ax113x) & (ax112x)) + ((!shiftx0x) & (!shiftx1x) & (ax115x) & (ax114x) & (!ax113x) & (!ax112x)) + ((!shiftx0x) & (!shiftx1x) & (ax115x) & (ax114x) & (!ax113x) & (ax112x)) + ((!shiftx0x) & (!shiftx1x) & (ax115x) & (ax114x) & (ax113x) & (!ax112x)) + ((!shiftx0x) & (!shiftx1x) & (ax115x) & (ax114x) & (ax113x) & (ax112x)) + ((!shiftx0x) & (shiftx1x) & (!ax115x) & (!ax114x) & (ax113x) & (!ax112x)) + ((!shiftx0x) & (shiftx1x) & (!ax115x) & (!ax114x) & (ax113x) & (ax112x)) + ((!shiftx0x) & (shiftx1x) & (!ax115x) & (ax114x) & (ax113x) & (!ax112x)) + ((!shiftx0x) & (shiftx1x) & (!ax115x) & (ax114x) & (ax113x) & (ax112x)) + ((!shiftx0x) & (shiftx1x) & (ax115x) & (!ax114x) & (ax113x) & (!ax112x)) + ((!shiftx0x) & (shiftx1x) & (ax115x) & (!ax114x) & (ax113x) & (ax112x)) + ((!shiftx0x) & (shiftx1x) & (ax115x) & (ax114x) & (ax113x) & (!ax112x)) + ((!shiftx0x) & (shiftx1x) & (ax115x) & (ax114x) & (ax113x) & (ax112x)) + ((shiftx0x) & (!shiftx1x) & (!ax115x) & (ax114x) & (!ax113x) & (!ax112x)) + ((shiftx0x) & (!shiftx1x) & (!ax115x) & (ax114x) & (!ax113x) & (ax112x)) + ((shiftx0x) & (!shiftx1x) & (!ax115x) & (ax114x) & (ax113x) & (!ax112x)) + ((shiftx0x) & (!shiftx1x) & (!ax115x) & (ax114x) & (ax113x) & (ax112x)) + ((shiftx0x) & (!shiftx1x) & (ax115x) & (ax114x) & (!ax113x) & (!ax112x)) + ((shiftx0x) & (!shiftx1x) & (ax115x) & (ax114x) & (!ax113x) & (ax112x)) + ((shiftx0x) & (!shiftx1x) & (ax115x) & (ax114x) & (ax113x) & (!ax112x)) + ((shiftx0x) & (!shiftx1x) & (ax115x) & (ax114x) & (ax113x) & (ax112x)) + ((shiftx0x) & (shiftx1x) & (!ax115x) & (!ax114x) & (!ax113x) & (ax112x)) + ((shiftx0x) & (shiftx1x) & (!ax115x) & (!ax114x) & (ax113x) & (ax112x)) + ((shiftx0x) & (shiftx1x) & (!ax115x) & (ax114x) & (!ax113x) & (ax112x)) + ((shiftx0x) & (shiftx1x) & (!ax115x) & (ax114x) & (ax113x) & (ax112x)) + ((shiftx0x) & (shiftx1x) & (ax115x) & (!ax114x) & (!ax113x) & (ax112x)) + ((shiftx0x) & (shiftx1x) & (ax115x) & (!ax114x) & (ax113x) & (ax112x)) + ((shiftx0x) & (shiftx1x) & (ax115x) & (ax114x) & (!ax113x) & (ax112x)) + ((shiftx0x) & (shiftx1x) & (ax115x) & (ax114x) & (ax113x) & (ax112x)));
	assign g152 = (((!shiftx0x) & (!shiftx1x) & (ax111x) & (!ax110x) & (!ax109x) & (!ax108x)) + ((!shiftx0x) & (!shiftx1x) & (ax111x) & (!ax110x) & (!ax109x) & (ax108x)) + ((!shiftx0x) & (!shiftx1x) & (ax111x) & (!ax110x) & (ax109x) & (!ax108x)) + ((!shiftx0x) & (!shiftx1x) & (ax111x) & (!ax110x) & (ax109x) & (ax108x)) + ((!shiftx0x) & (!shiftx1x) & (ax111x) & (ax110x) & (!ax109x) & (!ax108x)) + ((!shiftx0x) & (!shiftx1x) & (ax111x) & (ax110x) & (!ax109x) & (ax108x)) + ((!shiftx0x) & (!shiftx1x) & (ax111x) & (ax110x) & (ax109x) & (!ax108x)) + ((!shiftx0x) & (!shiftx1x) & (ax111x) & (ax110x) & (ax109x) & (ax108x)) + ((!shiftx0x) & (shiftx1x) & (!ax111x) & (!ax110x) & (ax109x) & (!ax108x)) + ((!shiftx0x) & (shiftx1x) & (!ax111x) & (!ax110x) & (ax109x) & (ax108x)) + ((!shiftx0x) & (shiftx1x) & (!ax111x) & (ax110x) & (ax109x) & (!ax108x)) + ((!shiftx0x) & (shiftx1x) & (!ax111x) & (ax110x) & (ax109x) & (ax108x)) + ((!shiftx0x) & (shiftx1x) & (ax111x) & (!ax110x) & (ax109x) & (!ax108x)) + ((!shiftx0x) & (shiftx1x) & (ax111x) & (!ax110x) & (ax109x) & (ax108x)) + ((!shiftx0x) & (shiftx1x) & (ax111x) & (ax110x) & (ax109x) & (!ax108x)) + ((!shiftx0x) & (shiftx1x) & (ax111x) & (ax110x) & (ax109x) & (ax108x)) + ((shiftx0x) & (!shiftx1x) & (!ax111x) & (ax110x) & (!ax109x) & (!ax108x)) + ((shiftx0x) & (!shiftx1x) & (!ax111x) & (ax110x) & (!ax109x) & (ax108x)) + ((shiftx0x) & (!shiftx1x) & (!ax111x) & (ax110x) & (ax109x) & (!ax108x)) + ((shiftx0x) & (!shiftx1x) & (!ax111x) & (ax110x) & (ax109x) & (ax108x)) + ((shiftx0x) & (!shiftx1x) & (ax111x) & (ax110x) & (!ax109x) & (!ax108x)) + ((shiftx0x) & (!shiftx1x) & (ax111x) & (ax110x) & (!ax109x) & (ax108x)) + ((shiftx0x) & (!shiftx1x) & (ax111x) & (ax110x) & (ax109x) & (!ax108x)) + ((shiftx0x) & (!shiftx1x) & (ax111x) & (ax110x) & (ax109x) & (ax108x)) + ((shiftx0x) & (shiftx1x) & (!ax111x) & (!ax110x) & (!ax109x) & (ax108x)) + ((shiftx0x) & (shiftx1x) & (!ax111x) & (!ax110x) & (ax109x) & (ax108x)) + ((shiftx0x) & (shiftx1x) & (!ax111x) & (ax110x) & (!ax109x) & (ax108x)) + ((shiftx0x) & (shiftx1x) & (!ax111x) & (ax110x) & (ax109x) & (ax108x)) + ((shiftx0x) & (shiftx1x) & (ax111x) & (!ax110x) & (!ax109x) & (ax108x)) + ((shiftx0x) & (shiftx1x) & (ax111x) & (!ax110x) & (ax109x) & (ax108x)) + ((shiftx0x) & (shiftx1x) & (ax111x) & (ax110x) & (!ax109x) & (ax108x)) + ((shiftx0x) & (shiftx1x) & (ax111x) & (ax110x) & (ax109x) & (ax108x)));
	assign g153 = (((!shiftx0x) & (!shiftx1x) & (!ax100x) & (ax103x) & (!ax102x) & (!ax101x)) + ((!shiftx0x) & (!shiftx1x) & (!ax100x) & (ax103x) & (!ax102x) & (ax101x)) + ((!shiftx0x) & (!shiftx1x) & (!ax100x) & (ax103x) & (ax102x) & (!ax101x)) + ((!shiftx0x) & (!shiftx1x) & (!ax100x) & (ax103x) & (ax102x) & (ax101x)) + ((!shiftx0x) & (!shiftx1x) & (ax100x) & (ax103x) & (!ax102x) & (!ax101x)) + ((!shiftx0x) & (!shiftx1x) & (ax100x) & (ax103x) & (!ax102x) & (ax101x)) + ((!shiftx0x) & (!shiftx1x) & (ax100x) & (ax103x) & (ax102x) & (!ax101x)) + ((!shiftx0x) & (!shiftx1x) & (ax100x) & (ax103x) & (ax102x) & (ax101x)) + ((!shiftx0x) & (shiftx1x) & (!ax100x) & (!ax103x) & (!ax102x) & (ax101x)) + ((!shiftx0x) & (shiftx1x) & (!ax100x) & (!ax103x) & (ax102x) & (ax101x)) + ((!shiftx0x) & (shiftx1x) & (!ax100x) & (ax103x) & (!ax102x) & (ax101x)) + ((!shiftx0x) & (shiftx1x) & (!ax100x) & (ax103x) & (ax102x) & (ax101x)) + ((!shiftx0x) & (shiftx1x) & (ax100x) & (!ax103x) & (!ax102x) & (ax101x)) + ((!shiftx0x) & (shiftx1x) & (ax100x) & (!ax103x) & (ax102x) & (ax101x)) + ((!shiftx0x) & (shiftx1x) & (ax100x) & (ax103x) & (!ax102x) & (ax101x)) + ((!shiftx0x) & (shiftx1x) & (ax100x) & (ax103x) & (ax102x) & (ax101x)) + ((shiftx0x) & (!shiftx1x) & (!ax100x) & (!ax103x) & (ax102x) & (!ax101x)) + ((shiftx0x) & (!shiftx1x) & (!ax100x) & (!ax103x) & (ax102x) & (ax101x)) + ((shiftx0x) & (!shiftx1x) & (!ax100x) & (ax103x) & (ax102x) & (!ax101x)) + ((shiftx0x) & (!shiftx1x) & (!ax100x) & (ax103x) & (ax102x) & (ax101x)) + ((shiftx0x) & (!shiftx1x) & (ax100x) & (!ax103x) & (ax102x) & (!ax101x)) + ((shiftx0x) & (!shiftx1x) & (ax100x) & (!ax103x) & (ax102x) & (ax101x)) + ((shiftx0x) & (!shiftx1x) & (ax100x) & (ax103x) & (ax102x) & (!ax101x)) + ((shiftx0x) & (!shiftx1x) & (ax100x) & (ax103x) & (ax102x) & (ax101x)) + ((shiftx0x) & (shiftx1x) & (ax100x) & (!ax103x) & (!ax102x) & (!ax101x)) + ((shiftx0x) & (shiftx1x) & (ax100x) & (!ax103x) & (!ax102x) & (ax101x)) + ((shiftx0x) & (shiftx1x) & (ax100x) & (!ax103x) & (ax102x) & (!ax101x)) + ((shiftx0x) & (shiftx1x) & (ax100x) & (!ax103x) & (ax102x) & (ax101x)) + ((shiftx0x) & (shiftx1x) & (ax100x) & (ax103x) & (!ax102x) & (!ax101x)) + ((shiftx0x) & (shiftx1x) & (ax100x) & (ax103x) & (!ax102x) & (ax101x)) + ((shiftx0x) & (shiftx1x) & (ax100x) & (ax103x) & (ax102x) & (!ax101x)) + ((shiftx0x) & (shiftx1x) & (ax100x) & (ax103x) & (ax102x) & (ax101x)));
	assign g154 = (((!shiftx0x) & (!shiftx1x) & (ax107x) & (!ax106x) & (!ax105x) & (!ax104x)) + ((!shiftx0x) & (!shiftx1x) & (ax107x) & (!ax106x) & (!ax105x) & (ax104x)) + ((!shiftx0x) & (!shiftx1x) & (ax107x) & (!ax106x) & (ax105x) & (!ax104x)) + ((!shiftx0x) & (!shiftx1x) & (ax107x) & (!ax106x) & (ax105x) & (ax104x)) + ((!shiftx0x) & (!shiftx1x) & (ax107x) & (ax106x) & (!ax105x) & (!ax104x)) + ((!shiftx0x) & (!shiftx1x) & (ax107x) & (ax106x) & (!ax105x) & (ax104x)) + ((!shiftx0x) & (!shiftx1x) & (ax107x) & (ax106x) & (ax105x) & (!ax104x)) + ((!shiftx0x) & (!shiftx1x) & (ax107x) & (ax106x) & (ax105x) & (ax104x)) + ((!shiftx0x) & (shiftx1x) & (!ax107x) & (!ax106x) & (ax105x) & (!ax104x)) + ((!shiftx0x) & (shiftx1x) & (!ax107x) & (!ax106x) & (ax105x) & (ax104x)) + ((!shiftx0x) & (shiftx1x) & (!ax107x) & (ax106x) & (ax105x) & (!ax104x)) + ((!shiftx0x) & (shiftx1x) & (!ax107x) & (ax106x) & (ax105x) & (ax104x)) + ((!shiftx0x) & (shiftx1x) & (ax107x) & (!ax106x) & (ax105x) & (!ax104x)) + ((!shiftx0x) & (shiftx1x) & (ax107x) & (!ax106x) & (ax105x) & (ax104x)) + ((!shiftx0x) & (shiftx1x) & (ax107x) & (ax106x) & (ax105x) & (!ax104x)) + ((!shiftx0x) & (shiftx1x) & (ax107x) & (ax106x) & (ax105x) & (ax104x)) + ((shiftx0x) & (!shiftx1x) & (!ax107x) & (ax106x) & (!ax105x) & (!ax104x)) + ((shiftx0x) & (!shiftx1x) & (!ax107x) & (ax106x) & (!ax105x) & (ax104x)) + ((shiftx0x) & (!shiftx1x) & (!ax107x) & (ax106x) & (ax105x) & (!ax104x)) + ((shiftx0x) & (!shiftx1x) & (!ax107x) & (ax106x) & (ax105x) & (ax104x)) + ((shiftx0x) & (!shiftx1x) & (ax107x) & (ax106x) & (!ax105x) & (!ax104x)) + ((shiftx0x) & (!shiftx1x) & (ax107x) & (ax106x) & (!ax105x) & (ax104x)) + ((shiftx0x) & (!shiftx1x) & (ax107x) & (ax106x) & (ax105x) & (!ax104x)) + ((shiftx0x) & (!shiftx1x) & (ax107x) & (ax106x) & (ax105x) & (ax104x)) + ((shiftx0x) & (shiftx1x) & (!ax107x) & (!ax106x) & (!ax105x) & (ax104x)) + ((shiftx0x) & (shiftx1x) & (!ax107x) & (!ax106x) & (ax105x) & (ax104x)) + ((shiftx0x) & (shiftx1x) & (!ax107x) & (ax106x) & (!ax105x) & (ax104x)) + ((shiftx0x) & (shiftx1x) & (!ax107x) & (ax106x) & (ax105x) & (ax104x)) + ((shiftx0x) & (shiftx1x) & (ax107x) & (!ax106x) & (!ax105x) & (ax104x)) + ((shiftx0x) & (shiftx1x) & (ax107x) & (!ax106x) & (ax105x) & (ax104x)) + ((shiftx0x) & (shiftx1x) & (ax107x) & (ax106x) & (!ax105x) & (ax104x)) + ((shiftx0x) & (shiftx1x) & (ax107x) & (ax106x) & (ax105x) & (ax104x)));
	assign g155 = (((!shiftx2x) & (!shiftx3x) & (g151) & (!g152) & (!g153) & (!g154)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (!g152) & (!g153) & (g154)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (!g152) & (g153) & (!g154)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (!g152) & (g153) & (g154)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (g152) & (!g153) & (!g154)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (g152) & (!g153) & (g154)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (g152) & (g153) & (!g154)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (g152) & (g153) & (g154)) + ((!shiftx2x) & (shiftx3x) & (!g151) & (!g152) & (!g153) & (g154)) + ((!shiftx2x) & (shiftx3x) & (!g151) & (!g152) & (g153) & (g154)) + ((!shiftx2x) & (shiftx3x) & (!g151) & (g152) & (!g153) & (g154)) + ((!shiftx2x) & (shiftx3x) & (!g151) & (g152) & (g153) & (g154)) + ((!shiftx2x) & (shiftx3x) & (g151) & (!g152) & (!g153) & (g154)) + ((!shiftx2x) & (shiftx3x) & (g151) & (!g152) & (g153) & (g154)) + ((!shiftx2x) & (shiftx3x) & (g151) & (g152) & (!g153) & (g154)) + ((!shiftx2x) & (shiftx3x) & (g151) & (g152) & (g153) & (g154)) + ((shiftx2x) & (!shiftx3x) & (!g151) & (g152) & (!g153) & (!g154)) + ((shiftx2x) & (!shiftx3x) & (!g151) & (g152) & (!g153) & (g154)) + ((shiftx2x) & (!shiftx3x) & (!g151) & (g152) & (g153) & (!g154)) + ((shiftx2x) & (!shiftx3x) & (!g151) & (g152) & (g153) & (g154)) + ((shiftx2x) & (!shiftx3x) & (g151) & (g152) & (!g153) & (!g154)) + ((shiftx2x) & (!shiftx3x) & (g151) & (g152) & (!g153) & (g154)) + ((shiftx2x) & (!shiftx3x) & (g151) & (g152) & (g153) & (!g154)) + ((shiftx2x) & (!shiftx3x) & (g151) & (g152) & (g153) & (g154)) + ((shiftx2x) & (shiftx3x) & (!g151) & (!g152) & (g153) & (!g154)) + ((shiftx2x) & (shiftx3x) & (!g151) & (!g152) & (g153) & (g154)) + ((shiftx2x) & (shiftx3x) & (!g151) & (g152) & (g153) & (!g154)) + ((shiftx2x) & (shiftx3x) & (!g151) & (g152) & (g153) & (g154)) + ((shiftx2x) & (shiftx3x) & (g151) & (!g152) & (g153) & (!g154)) + ((shiftx2x) & (shiftx3x) & (g151) & (!g152) & (g153) & (g154)) + ((shiftx2x) & (shiftx3x) & (g151) & (g152) & (g153) & (!g154)) + ((shiftx2x) & (shiftx3x) & (g151) & (g152) & (g153) & (g154)));
	assign g156 = (((!shiftx0x) & (!shiftx1x) & (!ax96x) & (ax99x) & (!ax98x) & (!ax97x)) + ((!shiftx0x) & (!shiftx1x) & (!ax96x) & (ax99x) & (!ax98x) & (ax97x)) + ((!shiftx0x) & (!shiftx1x) & (!ax96x) & (ax99x) & (ax98x) & (!ax97x)) + ((!shiftx0x) & (!shiftx1x) & (!ax96x) & (ax99x) & (ax98x) & (ax97x)) + ((!shiftx0x) & (!shiftx1x) & (ax96x) & (ax99x) & (!ax98x) & (!ax97x)) + ((!shiftx0x) & (!shiftx1x) & (ax96x) & (ax99x) & (!ax98x) & (ax97x)) + ((!shiftx0x) & (!shiftx1x) & (ax96x) & (ax99x) & (ax98x) & (!ax97x)) + ((!shiftx0x) & (!shiftx1x) & (ax96x) & (ax99x) & (ax98x) & (ax97x)) + ((!shiftx0x) & (shiftx1x) & (!ax96x) & (!ax99x) & (!ax98x) & (ax97x)) + ((!shiftx0x) & (shiftx1x) & (!ax96x) & (!ax99x) & (ax98x) & (ax97x)) + ((!shiftx0x) & (shiftx1x) & (!ax96x) & (ax99x) & (!ax98x) & (ax97x)) + ((!shiftx0x) & (shiftx1x) & (!ax96x) & (ax99x) & (ax98x) & (ax97x)) + ((!shiftx0x) & (shiftx1x) & (ax96x) & (!ax99x) & (!ax98x) & (ax97x)) + ((!shiftx0x) & (shiftx1x) & (ax96x) & (!ax99x) & (ax98x) & (ax97x)) + ((!shiftx0x) & (shiftx1x) & (ax96x) & (ax99x) & (!ax98x) & (ax97x)) + ((!shiftx0x) & (shiftx1x) & (ax96x) & (ax99x) & (ax98x) & (ax97x)) + ((shiftx0x) & (!shiftx1x) & (!ax96x) & (!ax99x) & (ax98x) & (!ax97x)) + ((shiftx0x) & (!shiftx1x) & (!ax96x) & (!ax99x) & (ax98x) & (ax97x)) + ((shiftx0x) & (!shiftx1x) & (!ax96x) & (ax99x) & (ax98x) & (!ax97x)) + ((shiftx0x) & (!shiftx1x) & (!ax96x) & (ax99x) & (ax98x) & (ax97x)) + ((shiftx0x) & (!shiftx1x) & (ax96x) & (!ax99x) & (ax98x) & (!ax97x)) + ((shiftx0x) & (!shiftx1x) & (ax96x) & (!ax99x) & (ax98x) & (ax97x)) + ((shiftx0x) & (!shiftx1x) & (ax96x) & (ax99x) & (ax98x) & (!ax97x)) + ((shiftx0x) & (!shiftx1x) & (ax96x) & (ax99x) & (ax98x) & (ax97x)) + ((shiftx0x) & (shiftx1x) & (ax96x) & (!ax99x) & (!ax98x) & (!ax97x)) + ((shiftx0x) & (shiftx1x) & (ax96x) & (!ax99x) & (!ax98x) & (ax97x)) + ((shiftx0x) & (shiftx1x) & (ax96x) & (!ax99x) & (ax98x) & (!ax97x)) + ((shiftx0x) & (shiftx1x) & (ax96x) & (!ax99x) & (ax98x) & (ax97x)) + ((shiftx0x) & (shiftx1x) & (ax96x) & (ax99x) & (!ax98x) & (!ax97x)) + ((shiftx0x) & (shiftx1x) & (ax96x) & (ax99x) & (!ax98x) & (ax97x)) + ((shiftx0x) & (shiftx1x) & (ax96x) & (ax99x) & (ax98x) & (!ax97x)) + ((shiftx0x) & (shiftx1x) & (ax96x) & (ax99x) & (ax98x) & (ax97x)));
	assign g157 = (((!shiftx0x) & (!shiftx1x) & (ax95x) & (!ax94x) & (!ax93x) & (!ax92x)) + ((!shiftx0x) & (!shiftx1x) & (ax95x) & (!ax94x) & (!ax93x) & (ax92x)) + ((!shiftx0x) & (!shiftx1x) & (ax95x) & (!ax94x) & (ax93x) & (!ax92x)) + ((!shiftx0x) & (!shiftx1x) & (ax95x) & (!ax94x) & (ax93x) & (ax92x)) + ((!shiftx0x) & (!shiftx1x) & (ax95x) & (ax94x) & (!ax93x) & (!ax92x)) + ((!shiftx0x) & (!shiftx1x) & (ax95x) & (ax94x) & (!ax93x) & (ax92x)) + ((!shiftx0x) & (!shiftx1x) & (ax95x) & (ax94x) & (ax93x) & (!ax92x)) + ((!shiftx0x) & (!shiftx1x) & (ax95x) & (ax94x) & (ax93x) & (ax92x)) + ((!shiftx0x) & (shiftx1x) & (!ax95x) & (!ax94x) & (ax93x) & (!ax92x)) + ((!shiftx0x) & (shiftx1x) & (!ax95x) & (!ax94x) & (ax93x) & (ax92x)) + ((!shiftx0x) & (shiftx1x) & (!ax95x) & (ax94x) & (ax93x) & (!ax92x)) + ((!shiftx0x) & (shiftx1x) & (!ax95x) & (ax94x) & (ax93x) & (ax92x)) + ((!shiftx0x) & (shiftx1x) & (ax95x) & (!ax94x) & (ax93x) & (!ax92x)) + ((!shiftx0x) & (shiftx1x) & (ax95x) & (!ax94x) & (ax93x) & (ax92x)) + ((!shiftx0x) & (shiftx1x) & (ax95x) & (ax94x) & (ax93x) & (!ax92x)) + ((!shiftx0x) & (shiftx1x) & (ax95x) & (ax94x) & (ax93x) & (ax92x)) + ((shiftx0x) & (!shiftx1x) & (!ax95x) & (ax94x) & (!ax93x) & (!ax92x)) + ((shiftx0x) & (!shiftx1x) & (!ax95x) & (ax94x) & (!ax93x) & (ax92x)) + ((shiftx0x) & (!shiftx1x) & (!ax95x) & (ax94x) & (ax93x) & (!ax92x)) + ((shiftx0x) & (!shiftx1x) & (!ax95x) & (ax94x) & (ax93x) & (ax92x)) + ((shiftx0x) & (!shiftx1x) & (ax95x) & (ax94x) & (!ax93x) & (!ax92x)) + ((shiftx0x) & (!shiftx1x) & (ax95x) & (ax94x) & (!ax93x) & (ax92x)) + ((shiftx0x) & (!shiftx1x) & (ax95x) & (ax94x) & (ax93x) & (!ax92x)) + ((shiftx0x) & (!shiftx1x) & (ax95x) & (ax94x) & (ax93x) & (ax92x)) + ((shiftx0x) & (shiftx1x) & (!ax95x) & (!ax94x) & (!ax93x) & (ax92x)) + ((shiftx0x) & (shiftx1x) & (!ax95x) & (!ax94x) & (ax93x) & (ax92x)) + ((shiftx0x) & (shiftx1x) & (!ax95x) & (ax94x) & (!ax93x) & (ax92x)) + ((shiftx0x) & (shiftx1x) & (!ax95x) & (ax94x) & (ax93x) & (ax92x)) + ((shiftx0x) & (shiftx1x) & (ax95x) & (!ax94x) & (!ax93x) & (ax92x)) + ((shiftx0x) & (shiftx1x) & (ax95x) & (!ax94x) & (ax93x) & (ax92x)) + ((shiftx0x) & (shiftx1x) & (ax95x) & (ax94x) & (!ax93x) & (ax92x)) + ((shiftx0x) & (shiftx1x) & (ax95x) & (ax94x) & (ax93x) & (ax92x)));
	assign g158 = (((!shiftx0x) & (!shiftx1x) & (!ax84x) & (ax87x) & (!ax86x) & (!ax85x)) + ((!shiftx0x) & (!shiftx1x) & (!ax84x) & (ax87x) & (!ax86x) & (ax85x)) + ((!shiftx0x) & (!shiftx1x) & (!ax84x) & (ax87x) & (ax86x) & (!ax85x)) + ((!shiftx0x) & (!shiftx1x) & (!ax84x) & (ax87x) & (ax86x) & (ax85x)) + ((!shiftx0x) & (!shiftx1x) & (ax84x) & (ax87x) & (!ax86x) & (!ax85x)) + ((!shiftx0x) & (!shiftx1x) & (ax84x) & (ax87x) & (!ax86x) & (ax85x)) + ((!shiftx0x) & (!shiftx1x) & (ax84x) & (ax87x) & (ax86x) & (!ax85x)) + ((!shiftx0x) & (!shiftx1x) & (ax84x) & (ax87x) & (ax86x) & (ax85x)) + ((!shiftx0x) & (shiftx1x) & (!ax84x) & (!ax87x) & (!ax86x) & (ax85x)) + ((!shiftx0x) & (shiftx1x) & (!ax84x) & (!ax87x) & (ax86x) & (ax85x)) + ((!shiftx0x) & (shiftx1x) & (!ax84x) & (ax87x) & (!ax86x) & (ax85x)) + ((!shiftx0x) & (shiftx1x) & (!ax84x) & (ax87x) & (ax86x) & (ax85x)) + ((!shiftx0x) & (shiftx1x) & (ax84x) & (!ax87x) & (!ax86x) & (ax85x)) + ((!shiftx0x) & (shiftx1x) & (ax84x) & (!ax87x) & (ax86x) & (ax85x)) + ((!shiftx0x) & (shiftx1x) & (ax84x) & (ax87x) & (!ax86x) & (ax85x)) + ((!shiftx0x) & (shiftx1x) & (ax84x) & (ax87x) & (ax86x) & (ax85x)) + ((shiftx0x) & (!shiftx1x) & (!ax84x) & (!ax87x) & (ax86x) & (!ax85x)) + ((shiftx0x) & (!shiftx1x) & (!ax84x) & (!ax87x) & (ax86x) & (ax85x)) + ((shiftx0x) & (!shiftx1x) & (!ax84x) & (ax87x) & (ax86x) & (!ax85x)) + ((shiftx0x) & (!shiftx1x) & (!ax84x) & (ax87x) & (ax86x) & (ax85x)) + ((shiftx0x) & (!shiftx1x) & (ax84x) & (!ax87x) & (ax86x) & (!ax85x)) + ((shiftx0x) & (!shiftx1x) & (ax84x) & (!ax87x) & (ax86x) & (ax85x)) + ((shiftx0x) & (!shiftx1x) & (ax84x) & (ax87x) & (ax86x) & (!ax85x)) + ((shiftx0x) & (!shiftx1x) & (ax84x) & (ax87x) & (ax86x) & (ax85x)) + ((shiftx0x) & (shiftx1x) & (ax84x) & (!ax87x) & (!ax86x) & (!ax85x)) + ((shiftx0x) & (shiftx1x) & (ax84x) & (!ax87x) & (!ax86x) & (ax85x)) + ((shiftx0x) & (shiftx1x) & (ax84x) & (!ax87x) & (ax86x) & (!ax85x)) + ((shiftx0x) & (shiftx1x) & (ax84x) & (!ax87x) & (ax86x) & (ax85x)) + ((shiftx0x) & (shiftx1x) & (ax84x) & (ax87x) & (!ax86x) & (!ax85x)) + ((shiftx0x) & (shiftx1x) & (ax84x) & (ax87x) & (!ax86x) & (ax85x)) + ((shiftx0x) & (shiftx1x) & (ax84x) & (ax87x) & (ax86x) & (!ax85x)) + ((shiftx0x) & (shiftx1x) & (ax84x) & (ax87x) & (ax86x) & (ax85x)));
	assign g159 = (((!shiftx0x) & (!shiftx1x) & (ax91x) & (!ax90x) & (!ax89x) & (!ax88x)) + ((!shiftx0x) & (!shiftx1x) & (ax91x) & (!ax90x) & (!ax89x) & (ax88x)) + ((!shiftx0x) & (!shiftx1x) & (ax91x) & (!ax90x) & (ax89x) & (!ax88x)) + ((!shiftx0x) & (!shiftx1x) & (ax91x) & (!ax90x) & (ax89x) & (ax88x)) + ((!shiftx0x) & (!shiftx1x) & (ax91x) & (ax90x) & (!ax89x) & (!ax88x)) + ((!shiftx0x) & (!shiftx1x) & (ax91x) & (ax90x) & (!ax89x) & (ax88x)) + ((!shiftx0x) & (!shiftx1x) & (ax91x) & (ax90x) & (ax89x) & (!ax88x)) + ((!shiftx0x) & (!shiftx1x) & (ax91x) & (ax90x) & (ax89x) & (ax88x)) + ((!shiftx0x) & (shiftx1x) & (!ax91x) & (!ax90x) & (ax89x) & (!ax88x)) + ((!shiftx0x) & (shiftx1x) & (!ax91x) & (!ax90x) & (ax89x) & (ax88x)) + ((!shiftx0x) & (shiftx1x) & (!ax91x) & (ax90x) & (ax89x) & (!ax88x)) + ((!shiftx0x) & (shiftx1x) & (!ax91x) & (ax90x) & (ax89x) & (ax88x)) + ((!shiftx0x) & (shiftx1x) & (ax91x) & (!ax90x) & (ax89x) & (!ax88x)) + ((!shiftx0x) & (shiftx1x) & (ax91x) & (!ax90x) & (ax89x) & (ax88x)) + ((!shiftx0x) & (shiftx1x) & (ax91x) & (ax90x) & (ax89x) & (!ax88x)) + ((!shiftx0x) & (shiftx1x) & (ax91x) & (ax90x) & (ax89x) & (ax88x)) + ((shiftx0x) & (!shiftx1x) & (!ax91x) & (ax90x) & (!ax89x) & (!ax88x)) + ((shiftx0x) & (!shiftx1x) & (!ax91x) & (ax90x) & (!ax89x) & (ax88x)) + ((shiftx0x) & (!shiftx1x) & (!ax91x) & (ax90x) & (ax89x) & (!ax88x)) + ((shiftx0x) & (!shiftx1x) & (!ax91x) & (ax90x) & (ax89x) & (ax88x)) + ((shiftx0x) & (!shiftx1x) & (ax91x) & (ax90x) & (!ax89x) & (!ax88x)) + ((shiftx0x) & (!shiftx1x) & (ax91x) & (ax90x) & (!ax89x) & (ax88x)) + ((shiftx0x) & (!shiftx1x) & (ax91x) & (ax90x) & (ax89x) & (!ax88x)) + ((shiftx0x) & (!shiftx1x) & (ax91x) & (ax90x) & (ax89x) & (ax88x)) + ((shiftx0x) & (shiftx1x) & (!ax91x) & (!ax90x) & (!ax89x) & (ax88x)) + ((shiftx0x) & (shiftx1x) & (!ax91x) & (!ax90x) & (ax89x) & (ax88x)) + ((shiftx0x) & (shiftx1x) & (!ax91x) & (ax90x) & (!ax89x) & (ax88x)) + ((shiftx0x) & (shiftx1x) & (!ax91x) & (ax90x) & (ax89x) & (ax88x)) + ((shiftx0x) & (shiftx1x) & (ax91x) & (!ax90x) & (!ax89x) & (ax88x)) + ((shiftx0x) & (shiftx1x) & (ax91x) & (!ax90x) & (ax89x) & (ax88x)) + ((shiftx0x) & (shiftx1x) & (ax91x) & (ax90x) & (!ax89x) & (ax88x)) + ((shiftx0x) & (shiftx1x) & (ax91x) & (ax90x) & (ax89x) & (ax88x)));
	assign g160 = (((!shiftx2x) & (!shiftx3x) & (g156) & (!g157) & (!g158) & (!g159)) + ((!shiftx2x) & (!shiftx3x) & (g156) & (!g157) & (!g158) & (g159)) + ((!shiftx2x) & (!shiftx3x) & (g156) & (!g157) & (g158) & (!g159)) + ((!shiftx2x) & (!shiftx3x) & (g156) & (!g157) & (g158) & (g159)) + ((!shiftx2x) & (!shiftx3x) & (g156) & (g157) & (!g158) & (!g159)) + ((!shiftx2x) & (!shiftx3x) & (g156) & (g157) & (!g158) & (g159)) + ((!shiftx2x) & (!shiftx3x) & (g156) & (g157) & (g158) & (!g159)) + ((!shiftx2x) & (!shiftx3x) & (g156) & (g157) & (g158) & (g159)) + ((!shiftx2x) & (shiftx3x) & (!g156) & (!g157) & (!g158) & (g159)) + ((!shiftx2x) & (shiftx3x) & (!g156) & (!g157) & (g158) & (g159)) + ((!shiftx2x) & (shiftx3x) & (!g156) & (g157) & (!g158) & (g159)) + ((!shiftx2x) & (shiftx3x) & (!g156) & (g157) & (g158) & (g159)) + ((!shiftx2x) & (shiftx3x) & (g156) & (!g157) & (!g158) & (g159)) + ((!shiftx2x) & (shiftx3x) & (g156) & (!g157) & (g158) & (g159)) + ((!shiftx2x) & (shiftx3x) & (g156) & (g157) & (!g158) & (g159)) + ((!shiftx2x) & (shiftx3x) & (g156) & (g157) & (g158) & (g159)) + ((shiftx2x) & (!shiftx3x) & (!g156) & (g157) & (!g158) & (!g159)) + ((shiftx2x) & (!shiftx3x) & (!g156) & (g157) & (!g158) & (g159)) + ((shiftx2x) & (!shiftx3x) & (!g156) & (g157) & (g158) & (!g159)) + ((shiftx2x) & (!shiftx3x) & (!g156) & (g157) & (g158) & (g159)) + ((shiftx2x) & (!shiftx3x) & (g156) & (g157) & (!g158) & (!g159)) + ((shiftx2x) & (!shiftx3x) & (g156) & (g157) & (!g158) & (g159)) + ((shiftx2x) & (!shiftx3x) & (g156) & (g157) & (g158) & (!g159)) + ((shiftx2x) & (!shiftx3x) & (g156) & (g157) & (g158) & (g159)) + ((shiftx2x) & (shiftx3x) & (!g156) & (!g157) & (g158) & (!g159)) + ((shiftx2x) & (shiftx3x) & (!g156) & (!g157) & (g158) & (g159)) + ((shiftx2x) & (shiftx3x) & (!g156) & (g157) & (g158) & (!g159)) + ((shiftx2x) & (shiftx3x) & (!g156) & (g157) & (g158) & (g159)) + ((shiftx2x) & (shiftx3x) & (g156) & (!g157) & (g158) & (!g159)) + ((shiftx2x) & (shiftx3x) & (g156) & (!g157) & (g158) & (g159)) + ((shiftx2x) & (shiftx3x) & (g156) & (g157) & (g158) & (!g159)) + ((shiftx2x) & (shiftx3x) & (g156) & (g157) & (g158) & (g159)));
	assign g161 = (((!shiftx0x) & (!shiftx1x) & (ax3x) & (!ax2x) & (!ax1x) & (!ax0x)) + ((!shiftx0x) & (!shiftx1x) & (ax3x) & (!ax2x) & (!ax1x) & (ax0x)) + ((!shiftx0x) & (!shiftx1x) & (ax3x) & (!ax2x) & (ax1x) & (!ax0x)) + ((!shiftx0x) & (!shiftx1x) & (ax3x) & (!ax2x) & (ax1x) & (ax0x)) + ((!shiftx0x) & (!shiftx1x) & (ax3x) & (ax2x) & (!ax1x) & (!ax0x)) + ((!shiftx0x) & (!shiftx1x) & (ax3x) & (ax2x) & (!ax1x) & (ax0x)) + ((!shiftx0x) & (!shiftx1x) & (ax3x) & (ax2x) & (ax1x) & (!ax0x)) + ((!shiftx0x) & (!shiftx1x) & (ax3x) & (ax2x) & (ax1x) & (ax0x)) + ((!shiftx0x) & (shiftx1x) & (!ax3x) & (!ax2x) & (ax1x) & (!ax0x)) + ((!shiftx0x) & (shiftx1x) & (!ax3x) & (!ax2x) & (ax1x) & (ax0x)) + ((!shiftx0x) & (shiftx1x) & (!ax3x) & (ax2x) & (ax1x) & (!ax0x)) + ((!shiftx0x) & (shiftx1x) & (!ax3x) & (ax2x) & (ax1x) & (ax0x)) + ((!shiftx0x) & (shiftx1x) & (ax3x) & (!ax2x) & (ax1x) & (!ax0x)) + ((!shiftx0x) & (shiftx1x) & (ax3x) & (!ax2x) & (ax1x) & (ax0x)) + ((!shiftx0x) & (shiftx1x) & (ax3x) & (ax2x) & (ax1x) & (!ax0x)) + ((!shiftx0x) & (shiftx1x) & (ax3x) & (ax2x) & (ax1x) & (ax0x)) + ((shiftx0x) & (!shiftx1x) & (!ax3x) & (ax2x) & (!ax1x) & (!ax0x)) + ((shiftx0x) & (!shiftx1x) & (!ax3x) & (ax2x) & (!ax1x) & (ax0x)) + ((shiftx0x) & (!shiftx1x) & (!ax3x) & (ax2x) & (ax1x) & (!ax0x)) + ((shiftx0x) & (!shiftx1x) & (!ax3x) & (ax2x) & (ax1x) & (ax0x)) + ((shiftx0x) & (!shiftx1x) & (ax3x) & (ax2x) & (!ax1x) & (!ax0x)) + ((shiftx0x) & (!shiftx1x) & (ax3x) & (ax2x) & (!ax1x) & (ax0x)) + ((shiftx0x) & (!shiftx1x) & (ax3x) & (ax2x) & (ax1x) & (!ax0x)) + ((shiftx0x) & (!shiftx1x) & (ax3x) & (ax2x) & (ax1x) & (ax0x)) + ((shiftx0x) & (shiftx1x) & (!ax3x) & (!ax2x) & (!ax1x) & (ax0x)) + ((shiftx0x) & (shiftx1x) & (!ax3x) & (!ax2x) & (ax1x) & (ax0x)) + ((shiftx0x) & (shiftx1x) & (!ax3x) & (ax2x) & (!ax1x) & (ax0x)) + ((shiftx0x) & (shiftx1x) & (!ax3x) & (ax2x) & (ax1x) & (ax0x)) + ((shiftx0x) & (shiftx1x) & (ax3x) & (!ax2x) & (!ax1x) & (ax0x)) + ((shiftx0x) & (shiftx1x) & (ax3x) & (!ax2x) & (ax1x) & (ax0x)) + ((shiftx0x) & (shiftx1x) & (ax3x) & (ax2x) & (!ax1x) & (ax0x)) + ((shiftx0x) & (shiftx1x) & (ax3x) & (ax2x) & (ax1x) & (ax0x)));
	assign g162 = (((!shiftx0x) & (!shiftx1x) & (ax127x) & (!ax126x) & (!ax125x) & (!ax124x)) + ((!shiftx0x) & (!shiftx1x) & (ax127x) & (!ax126x) & (!ax125x) & (ax124x)) + ((!shiftx0x) & (!shiftx1x) & (ax127x) & (!ax126x) & (ax125x) & (!ax124x)) + ((!shiftx0x) & (!shiftx1x) & (ax127x) & (!ax126x) & (ax125x) & (ax124x)) + ((!shiftx0x) & (!shiftx1x) & (ax127x) & (ax126x) & (!ax125x) & (!ax124x)) + ((!shiftx0x) & (!shiftx1x) & (ax127x) & (ax126x) & (!ax125x) & (ax124x)) + ((!shiftx0x) & (!shiftx1x) & (ax127x) & (ax126x) & (ax125x) & (!ax124x)) + ((!shiftx0x) & (!shiftx1x) & (ax127x) & (ax126x) & (ax125x) & (ax124x)) + ((!shiftx0x) & (shiftx1x) & (!ax127x) & (!ax126x) & (ax125x) & (!ax124x)) + ((!shiftx0x) & (shiftx1x) & (!ax127x) & (!ax126x) & (ax125x) & (ax124x)) + ((!shiftx0x) & (shiftx1x) & (!ax127x) & (ax126x) & (ax125x) & (!ax124x)) + ((!shiftx0x) & (shiftx1x) & (!ax127x) & (ax126x) & (ax125x) & (ax124x)) + ((!shiftx0x) & (shiftx1x) & (ax127x) & (!ax126x) & (ax125x) & (!ax124x)) + ((!shiftx0x) & (shiftx1x) & (ax127x) & (!ax126x) & (ax125x) & (ax124x)) + ((!shiftx0x) & (shiftx1x) & (ax127x) & (ax126x) & (ax125x) & (!ax124x)) + ((!shiftx0x) & (shiftx1x) & (ax127x) & (ax126x) & (ax125x) & (ax124x)) + ((shiftx0x) & (!shiftx1x) & (!ax127x) & (ax126x) & (!ax125x) & (!ax124x)) + ((shiftx0x) & (!shiftx1x) & (!ax127x) & (ax126x) & (!ax125x) & (ax124x)) + ((shiftx0x) & (!shiftx1x) & (!ax127x) & (ax126x) & (ax125x) & (!ax124x)) + ((shiftx0x) & (!shiftx1x) & (!ax127x) & (ax126x) & (ax125x) & (ax124x)) + ((shiftx0x) & (!shiftx1x) & (ax127x) & (ax126x) & (!ax125x) & (!ax124x)) + ((shiftx0x) & (!shiftx1x) & (ax127x) & (ax126x) & (!ax125x) & (ax124x)) + ((shiftx0x) & (!shiftx1x) & (ax127x) & (ax126x) & (ax125x) & (!ax124x)) + ((shiftx0x) & (!shiftx1x) & (ax127x) & (ax126x) & (ax125x) & (ax124x)) + ((shiftx0x) & (shiftx1x) & (!ax127x) & (!ax126x) & (!ax125x) & (ax124x)) + ((shiftx0x) & (shiftx1x) & (!ax127x) & (!ax126x) & (ax125x) & (ax124x)) + ((shiftx0x) & (shiftx1x) & (!ax127x) & (ax126x) & (!ax125x) & (ax124x)) + ((shiftx0x) & (shiftx1x) & (!ax127x) & (ax126x) & (ax125x) & (ax124x)) + ((shiftx0x) & (shiftx1x) & (ax127x) & (!ax126x) & (!ax125x) & (ax124x)) + ((shiftx0x) & (shiftx1x) & (ax127x) & (!ax126x) & (ax125x) & (ax124x)) + ((shiftx0x) & (shiftx1x) & (ax127x) & (ax126x) & (!ax125x) & (ax124x)) + ((shiftx0x) & (shiftx1x) & (ax127x) & (ax126x) & (ax125x) & (ax124x)));
	assign g163 = (((!shiftx0x) & (!shiftx1x) & (!ax116x) & (ax119x) & (!ax118x) & (!ax117x)) + ((!shiftx0x) & (!shiftx1x) & (!ax116x) & (ax119x) & (!ax118x) & (ax117x)) + ((!shiftx0x) & (!shiftx1x) & (!ax116x) & (ax119x) & (ax118x) & (!ax117x)) + ((!shiftx0x) & (!shiftx1x) & (!ax116x) & (ax119x) & (ax118x) & (ax117x)) + ((!shiftx0x) & (!shiftx1x) & (ax116x) & (ax119x) & (!ax118x) & (!ax117x)) + ((!shiftx0x) & (!shiftx1x) & (ax116x) & (ax119x) & (!ax118x) & (ax117x)) + ((!shiftx0x) & (!shiftx1x) & (ax116x) & (ax119x) & (ax118x) & (!ax117x)) + ((!shiftx0x) & (!shiftx1x) & (ax116x) & (ax119x) & (ax118x) & (ax117x)) + ((!shiftx0x) & (shiftx1x) & (!ax116x) & (!ax119x) & (!ax118x) & (ax117x)) + ((!shiftx0x) & (shiftx1x) & (!ax116x) & (!ax119x) & (ax118x) & (ax117x)) + ((!shiftx0x) & (shiftx1x) & (!ax116x) & (ax119x) & (!ax118x) & (ax117x)) + ((!shiftx0x) & (shiftx1x) & (!ax116x) & (ax119x) & (ax118x) & (ax117x)) + ((!shiftx0x) & (shiftx1x) & (ax116x) & (!ax119x) & (!ax118x) & (ax117x)) + ((!shiftx0x) & (shiftx1x) & (ax116x) & (!ax119x) & (ax118x) & (ax117x)) + ((!shiftx0x) & (shiftx1x) & (ax116x) & (ax119x) & (!ax118x) & (ax117x)) + ((!shiftx0x) & (shiftx1x) & (ax116x) & (ax119x) & (ax118x) & (ax117x)) + ((shiftx0x) & (!shiftx1x) & (!ax116x) & (!ax119x) & (ax118x) & (!ax117x)) + ((shiftx0x) & (!shiftx1x) & (!ax116x) & (!ax119x) & (ax118x) & (ax117x)) + ((shiftx0x) & (!shiftx1x) & (!ax116x) & (ax119x) & (ax118x) & (!ax117x)) + ((shiftx0x) & (!shiftx1x) & (!ax116x) & (ax119x) & (ax118x) & (ax117x)) + ((shiftx0x) & (!shiftx1x) & (ax116x) & (!ax119x) & (ax118x) & (!ax117x)) + ((shiftx0x) & (!shiftx1x) & (ax116x) & (!ax119x) & (ax118x) & (ax117x)) + ((shiftx0x) & (!shiftx1x) & (ax116x) & (ax119x) & (ax118x) & (!ax117x)) + ((shiftx0x) & (!shiftx1x) & (ax116x) & (ax119x) & (ax118x) & (ax117x)) + ((shiftx0x) & (shiftx1x) & (ax116x) & (!ax119x) & (!ax118x) & (!ax117x)) + ((shiftx0x) & (shiftx1x) & (ax116x) & (!ax119x) & (!ax118x) & (ax117x)) + ((shiftx0x) & (shiftx1x) & (ax116x) & (!ax119x) & (ax118x) & (!ax117x)) + ((shiftx0x) & (shiftx1x) & (ax116x) & (!ax119x) & (ax118x) & (ax117x)) + ((shiftx0x) & (shiftx1x) & (ax116x) & (ax119x) & (!ax118x) & (!ax117x)) + ((shiftx0x) & (shiftx1x) & (ax116x) & (ax119x) & (!ax118x) & (ax117x)) + ((shiftx0x) & (shiftx1x) & (ax116x) & (ax119x) & (ax118x) & (!ax117x)) + ((shiftx0x) & (shiftx1x) & (ax116x) & (ax119x) & (ax118x) & (ax117x)));
	assign g164 = (((!shiftx0x) & (!shiftx1x) & (ax123x) & (!ax122x) & (!ax121x) & (!ax120x)) + ((!shiftx0x) & (!shiftx1x) & (ax123x) & (!ax122x) & (!ax121x) & (ax120x)) + ((!shiftx0x) & (!shiftx1x) & (ax123x) & (!ax122x) & (ax121x) & (!ax120x)) + ((!shiftx0x) & (!shiftx1x) & (ax123x) & (!ax122x) & (ax121x) & (ax120x)) + ((!shiftx0x) & (!shiftx1x) & (ax123x) & (ax122x) & (!ax121x) & (!ax120x)) + ((!shiftx0x) & (!shiftx1x) & (ax123x) & (ax122x) & (!ax121x) & (ax120x)) + ((!shiftx0x) & (!shiftx1x) & (ax123x) & (ax122x) & (ax121x) & (!ax120x)) + ((!shiftx0x) & (!shiftx1x) & (ax123x) & (ax122x) & (ax121x) & (ax120x)) + ((!shiftx0x) & (shiftx1x) & (!ax123x) & (!ax122x) & (ax121x) & (!ax120x)) + ((!shiftx0x) & (shiftx1x) & (!ax123x) & (!ax122x) & (ax121x) & (ax120x)) + ((!shiftx0x) & (shiftx1x) & (!ax123x) & (ax122x) & (ax121x) & (!ax120x)) + ((!shiftx0x) & (shiftx1x) & (!ax123x) & (ax122x) & (ax121x) & (ax120x)) + ((!shiftx0x) & (shiftx1x) & (ax123x) & (!ax122x) & (ax121x) & (!ax120x)) + ((!shiftx0x) & (shiftx1x) & (ax123x) & (!ax122x) & (ax121x) & (ax120x)) + ((!shiftx0x) & (shiftx1x) & (ax123x) & (ax122x) & (ax121x) & (!ax120x)) + ((!shiftx0x) & (shiftx1x) & (ax123x) & (ax122x) & (ax121x) & (ax120x)) + ((shiftx0x) & (!shiftx1x) & (!ax123x) & (ax122x) & (!ax121x) & (!ax120x)) + ((shiftx0x) & (!shiftx1x) & (!ax123x) & (ax122x) & (!ax121x) & (ax120x)) + ((shiftx0x) & (!shiftx1x) & (!ax123x) & (ax122x) & (ax121x) & (!ax120x)) + ((shiftx0x) & (!shiftx1x) & (!ax123x) & (ax122x) & (ax121x) & (ax120x)) + ((shiftx0x) & (!shiftx1x) & (ax123x) & (ax122x) & (!ax121x) & (!ax120x)) + ((shiftx0x) & (!shiftx1x) & (ax123x) & (ax122x) & (!ax121x) & (ax120x)) + ((shiftx0x) & (!shiftx1x) & (ax123x) & (ax122x) & (ax121x) & (!ax120x)) + ((shiftx0x) & (!shiftx1x) & (ax123x) & (ax122x) & (ax121x) & (ax120x)) + ((shiftx0x) & (shiftx1x) & (!ax123x) & (!ax122x) & (!ax121x) & (ax120x)) + ((shiftx0x) & (shiftx1x) & (!ax123x) & (!ax122x) & (ax121x) & (ax120x)) + ((shiftx0x) & (shiftx1x) & (!ax123x) & (ax122x) & (!ax121x) & (ax120x)) + ((shiftx0x) & (shiftx1x) & (!ax123x) & (ax122x) & (ax121x) & (ax120x)) + ((shiftx0x) & (shiftx1x) & (ax123x) & (!ax122x) & (!ax121x) & (ax120x)) + ((shiftx0x) & (shiftx1x) & (ax123x) & (!ax122x) & (ax121x) & (ax120x)) + ((shiftx0x) & (shiftx1x) & (ax123x) & (ax122x) & (!ax121x) & (ax120x)) + ((shiftx0x) & (shiftx1x) & (ax123x) & (ax122x) & (ax121x) & (ax120x)));
	assign g165 = (((!shiftx2x) & (!shiftx3x) & (g161) & (!g162) & (!g163) & (!g164)) + ((!shiftx2x) & (!shiftx3x) & (g161) & (!g162) & (!g163) & (g164)) + ((!shiftx2x) & (!shiftx3x) & (g161) & (!g162) & (g163) & (!g164)) + ((!shiftx2x) & (!shiftx3x) & (g161) & (!g162) & (g163) & (g164)) + ((!shiftx2x) & (!shiftx3x) & (g161) & (g162) & (!g163) & (!g164)) + ((!shiftx2x) & (!shiftx3x) & (g161) & (g162) & (!g163) & (g164)) + ((!shiftx2x) & (!shiftx3x) & (g161) & (g162) & (g163) & (!g164)) + ((!shiftx2x) & (!shiftx3x) & (g161) & (g162) & (g163) & (g164)) + ((!shiftx2x) & (shiftx3x) & (!g161) & (!g162) & (!g163) & (g164)) + ((!shiftx2x) & (shiftx3x) & (!g161) & (!g162) & (g163) & (g164)) + ((!shiftx2x) & (shiftx3x) & (!g161) & (g162) & (!g163) & (g164)) + ((!shiftx2x) & (shiftx3x) & (!g161) & (g162) & (g163) & (g164)) + ((!shiftx2x) & (shiftx3x) & (g161) & (!g162) & (!g163) & (g164)) + ((!shiftx2x) & (shiftx3x) & (g161) & (!g162) & (g163) & (g164)) + ((!shiftx2x) & (shiftx3x) & (g161) & (g162) & (!g163) & (g164)) + ((!shiftx2x) & (shiftx3x) & (g161) & (g162) & (g163) & (g164)) + ((shiftx2x) & (!shiftx3x) & (!g161) & (g162) & (!g163) & (!g164)) + ((shiftx2x) & (!shiftx3x) & (!g161) & (g162) & (!g163) & (g164)) + ((shiftx2x) & (!shiftx3x) & (!g161) & (g162) & (g163) & (!g164)) + ((shiftx2x) & (!shiftx3x) & (!g161) & (g162) & (g163) & (g164)) + ((shiftx2x) & (!shiftx3x) & (g161) & (g162) & (!g163) & (!g164)) + ((shiftx2x) & (!shiftx3x) & (g161) & (g162) & (!g163) & (g164)) + ((shiftx2x) & (!shiftx3x) & (g161) & (g162) & (g163) & (!g164)) + ((shiftx2x) & (!shiftx3x) & (g161) & (g162) & (g163) & (g164)) + ((shiftx2x) & (shiftx3x) & (!g161) & (!g162) & (g163) & (!g164)) + ((shiftx2x) & (shiftx3x) & (!g161) & (!g162) & (g163) & (g164)) + ((shiftx2x) & (shiftx3x) & (!g161) & (g162) & (g163) & (!g164)) + ((shiftx2x) & (shiftx3x) & (!g161) & (g162) & (g163) & (g164)) + ((shiftx2x) & (shiftx3x) & (g161) & (!g162) & (g163) & (!g164)) + ((shiftx2x) & (shiftx3x) & (g161) & (!g162) & (g163) & (g164)) + ((shiftx2x) & (shiftx3x) & (g161) & (g162) & (g163) & (!g164)) + ((shiftx2x) & (shiftx3x) & (g161) & (g162) & (g163) & (g164)));
	assign g166 = (((!shiftx0x) & (!shiftx1x) & (!ax80x) & (ax83x) & (!ax82x) & (!ax81x)) + ((!shiftx0x) & (!shiftx1x) & (!ax80x) & (ax83x) & (!ax82x) & (ax81x)) + ((!shiftx0x) & (!shiftx1x) & (!ax80x) & (ax83x) & (ax82x) & (!ax81x)) + ((!shiftx0x) & (!shiftx1x) & (!ax80x) & (ax83x) & (ax82x) & (ax81x)) + ((!shiftx0x) & (!shiftx1x) & (ax80x) & (ax83x) & (!ax82x) & (!ax81x)) + ((!shiftx0x) & (!shiftx1x) & (ax80x) & (ax83x) & (!ax82x) & (ax81x)) + ((!shiftx0x) & (!shiftx1x) & (ax80x) & (ax83x) & (ax82x) & (!ax81x)) + ((!shiftx0x) & (!shiftx1x) & (ax80x) & (ax83x) & (ax82x) & (ax81x)) + ((!shiftx0x) & (shiftx1x) & (!ax80x) & (!ax83x) & (!ax82x) & (ax81x)) + ((!shiftx0x) & (shiftx1x) & (!ax80x) & (!ax83x) & (ax82x) & (ax81x)) + ((!shiftx0x) & (shiftx1x) & (!ax80x) & (ax83x) & (!ax82x) & (ax81x)) + ((!shiftx0x) & (shiftx1x) & (!ax80x) & (ax83x) & (ax82x) & (ax81x)) + ((!shiftx0x) & (shiftx1x) & (ax80x) & (!ax83x) & (!ax82x) & (ax81x)) + ((!shiftx0x) & (shiftx1x) & (ax80x) & (!ax83x) & (ax82x) & (ax81x)) + ((!shiftx0x) & (shiftx1x) & (ax80x) & (ax83x) & (!ax82x) & (ax81x)) + ((!shiftx0x) & (shiftx1x) & (ax80x) & (ax83x) & (ax82x) & (ax81x)) + ((shiftx0x) & (!shiftx1x) & (!ax80x) & (!ax83x) & (ax82x) & (!ax81x)) + ((shiftx0x) & (!shiftx1x) & (!ax80x) & (!ax83x) & (ax82x) & (ax81x)) + ((shiftx0x) & (!shiftx1x) & (!ax80x) & (ax83x) & (ax82x) & (!ax81x)) + ((shiftx0x) & (!shiftx1x) & (!ax80x) & (ax83x) & (ax82x) & (ax81x)) + ((shiftx0x) & (!shiftx1x) & (ax80x) & (!ax83x) & (ax82x) & (!ax81x)) + ((shiftx0x) & (!shiftx1x) & (ax80x) & (!ax83x) & (ax82x) & (ax81x)) + ((shiftx0x) & (!shiftx1x) & (ax80x) & (ax83x) & (ax82x) & (!ax81x)) + ((shiftx0x) & (!shiftx1x) & (ax80x) & (ax83x) & (ax82x) & (ax81x)) + ((shiftx0x) & (shiftx1x) & (ax80x) & (!ax83x) & (!ax82x) & (!ax81x)) + ((shiftx0x) & (shiftx1x) & (ax80x) & (!ax83x) & (!ax82x) & (ax81x)) + ((shiftx0x) & (shiftx1x) & (ax80x) & (!ax83x) & (ax82x) & (!ax81x)) + ((shiftx0x) & (shiftx1x) & (ax80x) & (!ax83x) & (ax82x) & (ax81x)) + ((shiftx0x) & (shiftx1x) & (ax80x) & (ax83x) & (!ax82x) & (!ax81x)) + ((shiftx0x) & (shiftx1x) & (ax80x) & (ax83x) & (!ax82x) & (ax81x)) + ((shiftx0x) & (shiftx1x) & (ax80x) & (ax83x) & (ax82x) & (!ax81x)) + ((shiftx0x) & (shiftx1x) & (ax80x) & (ax83x) & (ax82x) & (ax81x)));
	assign g167 = (((!shiftx0x) & (!shiftx1x) & (ax79x) & (!ax78x) & (!ax77x) & (!ax76x)) + ((!shiftx0x) & (!shiftx1x) & (ax79x) & (!ax78x) & (!ax77x) & (ax76x)) + ((!shiftx0x) & (!shiftx1x) & (ax79x) & (!ax78x) & (ax77x) & (!ax76x)) + ((!shiftx0x) & (!shiftx1x) & (ax79x) & (!ax78x) & (ax77x) & (ax76x)) + ((!shiftx0x) & (!shiftx1x) & (ax79x) & (ax78x) & (!ax77x) & (!ax76x)) + ((!shiftx0x) & (!shiftx1x) & (ax79x) & (ax78x) & (!ax77x) & (ax76x)) + ((!shiftx0x) & (!shiftx1x) & (ax79x) & (ax78x) & (ax77x) & (!ax76x)) + ((!shiftx0x) & (!shiftx1x) & (ax79x) & (ax78x) & (ax77x) & (ax76x)) + ((!shiftx0x) & (shiftx1x) & (!ax79x) & (!ax78x) & (ax77x) & (!ax76x)) + ((!shiftx0x) & (shiftx1x) & (!ax79x) & (!ax78x) & (ax77x) & (ax76x)) + ((!shiftx0x) & (shiftx1x) & (!ax79x) & (ax78x) & (ax77x) & (!ax76x)) + ((!shiftx0x) & (shiftx1x) & (!ax79x) & (ax78x) & (ax77x) & (ax76x)) + ((!shiftx0x) & (shiftx1x) & (ax79x) & (!ax78x) & (ax77x) & (!ax76x)) + ((!shiftx0x) & (shiftx1x) & (ax79x) & (!ax78x) & (ax77x) & (ax76x)) + ((!shiftx0x) & (shiftx1x) & (ax79x) & (ax78x) & (ax77x) & (!ax76x)) + ((!shiftx0x) & (shiftx1x) & (ax79x) & (ax78x) & (ax77x) & (ax76x)) + ((shiftx0x) & (!shiftx1x) & (!ax79x) & (ax78x) & (!ax77x) & (!ax76x)) + ((shiftx0x) & (!shiftx1x) & (!ax79x) & (ax78x) & (!ax77x) & (ax76x)) + ((shiftx0x) & (!shiftx1x) & (!ax79x) & (ax78x) & (ax77x) & (!ax76x)) + ((shiftx0x) & (!shiftx1x) & (!ax79x) & (ax78x) & (ax77x) & (ax76x)) + ((shiftx0x) & (!shiftx1x) & (ax79x) & (ax78x) & (!ax77x) & (!ax76x)) + ((shiftx0x) & (!shiftx1x) & (ax79x) & (ax78x) & (!ax77x) & (ax76x)) + ((shiftx0x) & (!shiftx1x) & (ax79x) & (ax78x) & (ax77x) & (!ax76x)) + ((shiftx0x) & (!shiftx1x) & (ax79x) & (ax78x) & (ax77x) & (ax76x)) + ((shiftx0x) & (shiftx1x) & (!ax79x) & (!ax78x) & (!ax77x) & (ax76x)) + ((shiftx0x) & (shiftx1x) & (!ax79x) & (!ax78x) & (ax77x) & (ax76x)) + ((shiftx0x) & (shiftx1x) & (!ax79x) & (ax78x) & (!ax77x) & (ax76x)) + ((shiftx0x) & (shiftx1x) & (!ax79x) & (ax78x) & (ax77x) & (ax76x)) + ((shiftx0x) & (shiftx1x) & (ax79x) & (!ax78x) & (!ax77x) & (ax76x)) + ((shiftx0x) & (shiftx1x) & (ax79x) & (!ax78x) & (ax77x) & (ax76x)) + ((shiftx0x) & (shiftx1x) & (ax79x) & (ax78x) & (!ax77x) & (ax76x)) + ((shiftx0x) & (shiftx1x) & (ax79x) & (ax78x) & (ax77x) & (ax76x)));
	assign g168 = (((!shiftx0x) & (!shiftx1x) & (!ax68x) & (ax71x) & (!ax70x) & (!ax69x)) + ((!shiftx0x) & (!shiftx1x) & (!ax68x) & (ax71x) & (!ax70x) & (ax69x)) + ((!shiftx0x) & (!shiftx1x) & (!ax68x) & (ax71x) & (ax70x) & (!ax69x)) + ((!shiftx0x) & (!shiftx1x) & (!ax68x) & (ax71x) & (ax70x) & (ax69x)) + ((!shiftx0x) & (!shiftx1x) & (ax68x) & (ax71x) & (!ax70x) & (!ax69x)) + ((!shiftx0x) & (!shiftx1x) & (ax68x) & (ax71x) & (!ax70x) & (ax69x)) + ((!shiftx0x) & (!shiftx1x) & (ax68x) & (ax71x) & (ax70x) & (!ax69x)) + ((!shiftx0x) & (!shiftx1x) & (ax68x) & (ax71x) & (ax70x) & (ax69x)) + ((!shiftx0x) & (shiftx1x) & (!ax68x) & (!ax71x) & (!ax70x) & (ax69x)) + ((!shiftx0x) & (shiftx1x) & (!ax68x) & (!ax71x) & (ax70x) & (ax69x)) + ((!shiftx0x) & (shiftx1x) & (!ax68x) & (ax71x) & (!ax70x) & (ax69x)) + ((!shiftx0x) & (shiftx1x) & (!ax68x) & (ax71x) & (ax70x) & (ax69x)) + ((!shiftx0x) & (shiftx1x) & (ax68x) & (!ax71x) & (!ax70x) & (ax69x)) + ((!shiftx0x) & (shiftx1x) & (ax68x) & (!ax71x) & (ax70x) & (ax69x)) + ((!shiftx0x) & (shiftx1x) & (ax68x) & (ax71x) & (!ax70x) & (ax69x)) + ((!shiftx0x) & (shiftx1x) & (ax68x) & (ax71x) & (ax70x) & (ax69x)) + ((shiftx0x) & (!shiftx1x) & (!ax68x) & (!ax71x) & (ax70x) & (!ax69x)) + ((shiftx0x) & (!shiftx1x) & (!ax68x) & (!ax71x) & (ax70x) & (ax69x)) + ((shiftx0x) & (!shiftx1x) & (!ax68x) & (ax71x) & (ax70x) & (!ax69x)) + ((shiftx0x) & (!shiftx1x) & (!ax68x) & (ax71x) & (ax70x) & (ax69x)) + ((shiftx0x) & (!shiftx1x) & (ax68x) & (!ax71x) & (ax70x) & (!ax69x)) + ((shiftx0x) & (!shiftx1x) & (ax68x) & (!ax71x) & (ax70x) & (ax69x)) + ((shiftx0x) & (!shiftx1x) & (ax68x) & (ax71x) & (ax70x) & (!ax69x)) + ((shiftx0x) & (!shiftx1x) & (ax68x) & (ax71x) & (ax70x) & (ax69x)) + ((shiftx0x) & (shiftx1x) & (ax68x) & (!ax71x) & (!ax70x) & (!ax69x)) + ((shiftx0x) & (shiftx1x) & (ax68x) & (!ax71x) & (!ax70x) & (ax69x)) + ((shiftx0x) & (shiftx1x) & (ax68x) & (!ax71x) & (ax70x) & (!ax69x)) + ((shiftx0x) & (shiftx1x) & (ax68x) & (!ax71x) & (ax70x) & (ax69x)) + ((shiftx0x) & (shiftx1x) & (ax68x) & (ax71x) & (!ax70x) & (!ax69x)) + ((shiftx0x) & (shiftx1x) & (ax68x) & (ax71x) & (!ax70x) & (ax69x)) + ((shiftx0x) & (shiftx1x) & (ax68x) & (ax71x) & (ax70x) & (!ax69x)) + ((shiftx0x) & (shiftx1x) & (ax68x) & (ax71x) & (ax70x) & (ax69x)));
	assign g169 = (((!shiftx0x) & (!shiftx1x) & (ax75x) & (!ax74x) & (!ax73x) & (!ax72x)) + ((!shiftx0x) & (!shiftx1x) & (ax75x) & (!ax74x) & (!ax73x) & (ax72x)) + ((!shiftx0x) & (!shiftx1x) & (ax75x) & (!ax74x) & (ax73x) & (!ax72x)) + ((!shiftx0x) & (!shiftx1x) & (ax75x) & (!ax74x) & (ax73x) & (ax72x)) + ((!shiftx0x) & (!shiftx1x) & (ax75x) & (ax74x) & (!ax73x) & (!ax72x)) + ((!shiftx0x) & (!shiftx1x) & (ax75x) & (ax74x) & (!ax73x) & (ax72x)) + ((!shiftx0x) & (!shiftx1x) & (ax75x) & (ax74x) & (ax73x) & (!ax72x)) + ((!shiftx0x) & (!shiftx1x) & (ax75x) & (ax74x) & (ax73x) & (ax72x)) + ((!shiftx0x) & (shiftx1x) & (!ax75x) & (!ax74x) & (ax73x) & (!ax72x)) + ((!shiftx0x) & (shiftx1x) & (!ax75x) & (!ax74x) & (ax73x) & (ax72x)) + ((!shiftx0x) & (shiftx1x) & (!ax75x) & (ax74x) & (ax73x) & (!ax72x)) + ((!shiftx0x) & (shiftx1x) & (!ax75x) & (ax74x) & (ax73x) & (ax72x)) + ((!shiftx0x) & (shiftx1x) & (ax75x) & (!ax74x) & (ax73x) & (!ax72x)) + ((!shiftx0x) & (shiftx1x) & (ax75x) & (!ax74x) & (ax73x) & (ax72x)) + ((!shiftx0x) & (shiftx1x) & (ax75x) & (ax74x) & (ax73x) & (!ax72x)) + ((!shiftx0x) & (shiftx1x) & (ax75x) & (ax74x) & (ax73x) & (ax72x)) + ((shiftx0x) & (!shiftx1x) & (!ax75x) & (ax74x) & (!ax73x) & (!ax72x)) + ((shiftx0x) & (!shiftx1x) & (!ax75x) & (ax74x) & (!ax73x) & (ax72x)) + ((shiftx0x) & (!shiftx1x) & (!ax75x) & (ax74x) & (ax73x) & (!ax72x)) + ((shiftx0x) & (!shiftx1x) & (!ax75x) & (ax74x) & (ax73x) & (ax72x)) + ((shiftx0x) & (!shiftx1x) & (ax75x) & (ax74x) & (!ax73x) & (!ax72x)) + ((shiftx0x) & (!shiftx1x) & (ax75x) & (ax74x) & (!ax73x) & (ax72x)) + ((shiftx0x) & (!shiftx1x) & (ax75x) & (ax74x) & (ax73x) & (!ax72x)) + ((shiftx0x) & (!shiftx1x) & (ax75x) & (ax74x) & (ax73x) & (ax72x)) + ((shiftx0x) & (shiftx1x) & (!ax75x) & (!ax74x) & (!ax73x) & (ax72x)) + ((shiftx0x) & (shiftx1x) & (!ax75x) & (!ax74x) & (ax73x) & (ax72x)) + ((shiftx0x) & (shiftx1x) & (!ax75x) & (ax74x) & (!ax73x) & (ax72x)) + ((shiftx0x) & (shiftx1x) & (!ax75x) & (ax74x) & (ax73x) & (ax72x)) + ((shiftx0x) & (shiftx1x) & (ax75x) & (!ax74x) & (!ax73x) & (ax72x)) + ((shiftx0x) & (shiftx1x) & (ax75x) & (!ax74x) & (ax73x) & (ax72x)) + ((shiftx0x) & (shiftx1x) & (ax75x) & (ax74x) & (!ax73x) & (ax72x)) + ((shiftx0x) & (shiftx1x) & (ax75x) & (ax74x) & (ax73x) & (ax72x)));
	assign g170 = (((!shiftx2x) & (!shiftx3x) & (g166) & (!g167) & (!g168) & (!g169)) + ((!shiftx2x) & (!shiftx3x) & (g166) & (!g167) & (!g168) & (g169)) + ((!shiftx2x) & (!shiftx3x) & (g166) & (!g167) & (g168) & (!g169)) + ((!shiftx2x) & (!shiftx3x) & (g166) & (!g167) & (g168) & (g169)) + ((!shiftx2x) & (!shiftx3x) & (g166) & (g167) & (!g168) & (!g169)) + ((!shiftx2x) & (!shiftx3x) & (g166) & (g167) & (!g168) & (g169)) + ((!shiftx2x) & (!shiftx3x) & (g166) & (g167) & (g168) & (!g169)) + ((!shiftx2x) & (!shiftx3x) & (g166) & (g167) & (g168) & (g169)) + ((!shiftx2x) & (shiftx3x) & (!g166) & (!g167) & (!g168) & (g169)) + ((!shiftx2x) & (shiftx3x) & (!g166) & (!g167) & (g168) & (g169)) + ((!shiftx2x) & (shiftx3x) & (!g166) & (g167) & (!g168) & (g169)) + ((!shiftx2x) & (shiftx3x) & (!g166) & (g167) & (g168) & (g169)) + ((!shiftx2x) & (shiftx3x) & (g166) & (!g167) & (!g168) & (g169)) + ((!shiftx2x) & (shiftx3x) & (g166) & (!g167) & (g168) & (g169)) + ((!shiftx2x) & (shiftx3x) & (g166) & (g167) & (!g168) & (g169)) + ((!shiftx2x) & (shiftx3x) & (g166) & (g167) & (g168) & (g169)) + ((shiftx2x) & (!shiftx3x) & (!g166) & (g167) & (!g168) & (!g169)) + ((shiftx2x) & (!shiftx3x) & (!g166) & (g167) & (!g168) & (g169)) + ((shiftx2x) & (!shiftx3x) & (!g166) & (g167) & (g168) & (!g169)) + ((shiftx2x) & (!shiftx3x) & (!g166) & (g167) & (g168) & (g169)) + ((shiftx2x) & (!shiftx3x) & (g166) & (g167) & (!g168) & (!g169)) + ((shiftx2x) & (!shiftx3x) & (g166) & (g167) & (!g168) & (g169)) + ((shiftx2x) & (!shiftx3x) & (g166) & (g167) & (g168) & (!g169)) + ((shiftx2x) & (!shiftx3x) & (g166) & (g167) & (g168) & (g169)) + ((shiftx2x) & (shiftx3x) & (!g166) & (!g167) & (g168) & (!g169)) + ((shiftx2x) & (shiftx3x) & (!g166) & (!g167) & (g168) & (g169)) + ((shiftx2x) & (shiftx3x) & (!g166) & (g167) & (g168) & (!g169)) + ((shiftx2x) & (shiftx3x) & (!g166) & (g167) & (g168) & (g169)) + ((shiftx2x) & (shiftx3x) & (g166) & (!g167) & (g168) & (!g169)) + ((shiftx2x) & (shiftx3x) & (g166) & (!g167) & (g168) & (g169)) + ((shiftx2x) & (shiftx3x) & (g166) & (g167) & (g168) & (!g169)) + ((shiftx2x) & (shiftx3x) & (g166) & (g167) & (g168) & (g169)));
	assign g171 = (((!shiftx4x) & (!shiftx5x) & (!g155) & (!g160) & (g165) & (!g170)) + ((!shiftx4x) & (!shiftx5x) & (!g155) & (!g160) & (g165) & (g170)) + ((!shiftx4x) & (!shiftx5x) & (!g155) & (g160) & (g165) & (!g170)) + ((!shiftx4x) & (!shiftx5x) & (!g155) & (g160) & (g165) & (g170)) + ((!shiftx4x) & (!shiftx5x) & (g155) & (!g160) & (g165) & (!g170)) + ((!shiftx4x) & (!shiftx5x) & (g155) & (!g160) & (g165) & (g170)) + ((!shiftx4x) & (!shiftx5x) & (g155) & (g160) & (g165) & (!g170)) + ((!shiftx4x) & (!shiftx5x) & (g155) & (g160) & (g165) & (g170)) + ((!shiftx4x) & (shiftx5x) & (!g155) & (g160) & (!g165) & (!g170)) + ((!shiftx4x) & (shiftx5x) & (!g155) & (g160) & (!g165) & (g170)) + ((!shiftx4x) & (shiftx5x) & (!g155) & (g160) & (g165) & (!g170)) + ((!shiftx4x) & (shiftx5x) & (!g155) & (g160) & (g165) & (g170)) + ((!shiftx4x) & (shiftx5x) & (g155) & (g160) & (!g165) & (!g170)) + ((!shiftx4x) & (shiftx5x) & (g155) & (g160) & (!g165) & (g170)) + ((!shiftx4x) & (shiftx5x) & (g155) & (g160) & (g165) & (!g170)) + ((!shiftx4x) & (shiftx5x) & (g155) & (g160) & (g165) & (g170)) + ((shiftx4x) & (!shiftx5x) & (g155) & (!g160) & (!g165) & (!g170)) + ((shiftx4x) & (!shiftx5x) & (g155) & (!g160) & (!g165) & (g170)) + ((shiftx4x) & (!shiftx5x) & (g155) & (!g160) & (g165) & (!g170)) + ((shiftx4x) & (!shiftx5x) & (g155) & (!g160) & (g165) & (g170)) + ((shiftx4x) & (!shiftx5x) & (g155) & (g160) & (!g165) & (!g170)) + ((shiftx4x) & (!shiftx5x) & (g155) & (g160) & (!g165) & (g170)) + ((shiftx4x) & (!shiftx5x) & (g155) & (g160) & (g165) & (!g170)) + ((shiftx4x) & (!shiftx5x) & (g155) & (g160) & (g165) & (g170)) + ((shiftx4x) & (shiftx5x) & (!g155) & (!g160) & (!g165) & (g170)) + ((shiftx4x) & (shiftx5x) & (!g155) & (!g160) & (g165) & (g170)) + ((shiftx4x) & (shiftx5x) & (!g155) & (g160) & (!g165) & (g170)) + ((shiftx4x) & (shiftx5x) & (!g155) & (g160) & (g165) & (g170)) + ((shiftx4x) & (shiftx5x) & (g155) & (!g160) & (!g165) & (g170)) + ((shiftx4x) & (shiftx5x) & (g155) & (!g160) & (g165) & (g170)) + ((shiftx4x) & (shiftx5x) & (g155) & (g160) & (!g165) & (g170)) + ((shiftx4x) & (shiftx5x) & (g155) & (g160) & (g165) & (g170)));
	assign resultx3x = (((!sk[43]) & (shiftx6x) & (!g150) & (!g171)) + ((!sk[43]) & (shiftx6x) & (!g150) & (g171)) + ((!sk[43]) & (shiftx6x) & (g150) & (!g171)) + ((!sk[43]) & (shiftx6x) & (g150) & (g171)) + ((sk[43]) & (!shiftx6x) & (!g150) & (g171)) + ((sk[43]) & (!shiftx6x) & (g150) & (g171)) + ((sk[43]) & (shiftx6x) & (g150) & (!g171)) + ((sk[43]) & (shiftx6x) & (g150) & (g171)));
	assign g173 = (((!shiftx2x) & (!shiftx3x) & (g13) & (!g16) & (!g17) & (!g19)) + ((!shiftx2x) & (!shiftx3x) & (g13) & (!g16) & (!g17) & (g19)) + ((!shiftx2x) & (!shiftx3x) & (g13) & (!g16) & (g17) & (!g19)) + ((!shiftx2x) & (!shiftx3x) & (g13) & (!g16) & (g17) & (g19)) + ((!shiftx2x) & (!shiftx3x) & (g13) & (g16) & (!g17) & (!g19)) + ((!shiftx2x) & (!shiftx3x) & (g13) & (g16) & (!g17) & (g19)) + ((!shiftx2x) & (!shiftx3x) & (g13) & (g16) & (g17) & (!g19)) + ((!shiftx2x) & (!shiftx3x) & (g13) & (g16) & (g17) & (g19)) + ((!shiftx2x) & (shiftx3x) & (!g13) & (!g16) & (g17) & (!g19)) + ((!shiftx2x) & (shiftx3x) & (!g13) & (!g16) & (g17) & (g19)) + ((!shiftx2x) & (shiftx3x) & (!g13) & (g16) & (g17) & (!g19)) + ((!shiftx2x) & (shiftx3x) & (!g13) & (g16) & (g17) & (g19)) + ((!shiftx2x) & (shiftx3x) & (g13) & (!g16) & (g17) & (!g19)) + ((!shiftx2x) & (shiftx3x) & (g13) & (!g16) & (g17) & (g19)) + ((!shiftx2x) & (shiftx3x) & (g13) & (g16) & (g17) & (!g19)) + ((!shiftx2x) & (shiftx3x) & (g13) & (g16) & (g17) & (g19)) + ((shiftx2x) & (!shiftx3x) & (!g13) & (g16) & (!g17) & (!g19)) + ((shiftx2x) & (!shiftx3x) & (!g13) & (g16) & (!g17) & (g19)) + ((shiftx2x) & (!shiftx3x) & (!g13) & (g16) & (g17) & (!g19)) + ((shiftx2x) & (!shiftx3x) & (!g13) & (g16) & (g17) & (g19)) + ((shiftx2x) & (!shiftx3x) & (g13) & (g16) & (!g17) & (!g19)) + ((shiftx2x) & (!shiftx3x) & (g13) & (g16) & (!g17) & (g19)) + ((shiftx2x) & (!shiftx3x) & (g13) & (g16) & (g17) & (!g19)) + ((shiftx2x) & (!shiftx3x) & (g13) & (g16) & (g17) & (g19)) + ((shiftx2x) & (shiftx3x) & (!g13) & (!g16) & (!g17) & (g19)) + ((shiftx2x) & (shiftx3x) & (!g13) & (!g16) & (g17) & (g19)) + ((shiftx2x) & (shiftx3x) & (!g13) & (g16) & (!g17) & (g19)) + ((shiftx2x) & (shiftx3x) & (!g13) & (g16) & (g17) & (g19)) + ((shiftx2x) & (shiftx3x) & (g13) & (!g16) & (!g17) & (g19)) + ((shiftx2x) & (shiftx3x) & (g13) & (!g16) & (g17) & (g19)) + ((shiftx2x) & (shiftx3x) & (g13) & (g16) & (!g17) & (g19)) + ((shiftx2x) & (shiftx3x) & (g13) & (g16) & (g17) & (g19)));
	assign g174 = (((!shiftx2x) & (!shiftx3x) & (!g11) & (!g12) & (!g14) & (g24)) + ((!shiftx2x) & (!shiftx3x) & (!g11) & (!g12) & (g14) & (g24)) + ((!shiftx2x) & (!shiftx3x) & (!g11) & (g12) & (!g14) & (g24)) + ((!shiftx2x) & (!shiftx3x) & (!g11) & (g12) & (g14) & (g24)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (!g12) & (!g14) & (g24)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (!g12) & (g14) & (g24)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (g12) & (!g14) & (g24)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (g12) & (g14) & (g24)) + ((!shiftx2x) & (shiftx3x) & (!g11) & (g12) & (!g14) & (!g24)) + ((!shiftx2x) & (shiftx3x) & (!g11) & (g12) & (!g14) & (g24)) + ((!shiftx2x) & (shiftx3x) & (!g11) & (g12) & (g14) & (!g24)) + ((!shiftx2x) & (shiftx3x) & (!g11) & (g12) & (g14) & (g24)) + ((!shiftx2x) & (shiftx3x) & (g11) & (g12) & (!g14) & (!g24)) + ((!shiftx2x) & (shiftx3x) & (g11) & (g12) & (!g14) & (g24)) + ((!shiftx2x) & (shiftx3x) & (g11) & (g12) & (g14) & (!g24)) + ((!shiftx2x) & (shiftx3x) & (g11) & (g12) & (g14) & (g24)) + ((shiftx2x) & (!shiftx3x) & (g11) & (!g12) & (!g14) & (!g24)) + ((shiftx2x) & (!shiftx3x) & (g11) & (!g12) & (!g14) & (g24)) + ((shiftx2x) & (!shiftx3x) & (g11) & (!g12) & (g14) & (!g24)) + ((shiftx2x) & (!shiftx3x) & (g11) & (!g12) & (g14) & (g24)) + ((shiftx2x) & (!shiftx3x) & (g11) & (g12) & (!g14) & (!g24)) + ((shiftx2x) & (!shiftx3x) & (g11) & (g12) & (!g14) & (g24)) + ((shiftx2x) & (!shiftx3x) & (g11) & (g12) & (g14) & (!g24)) + ((shiftx2x) & (!shiftx3x) & (g11) & (g12) & (g14) & (g24)) + ((shiftx2x) & (shiftx3x) & (!g11) & (!g12) & (g14) & (!g24)) + ((shiftx2x) & (shiftx3x) & (!g11) & (!g12) & (g14) & (g24)) + ((shiftx2x) & (shiftx3x) & (!g11) & (g12) & (g14) & (!g24)) + ((shiftx2x) & (shiftx3x) & (!g11) & (g12) & (g14) & (g24)) + ((shiftx2x) & (shiftx3x) & (g11) & (!g12) & (g14) & (!g24)) + ((shiftx2x) & (shiftx3x) & (g11) & (!g12) & (g14) & (g24)) + ((shiftx2x) & (shiftx3x) & (g11) & (g12) & (g14) & (!g24)) + ((shiftx2x) & (shiftx3x) & (g11) & (g12) & (g14) & (g24)));
	assign g175 = (((!shiftx2x) & (!shiftx3x) & (!g6) & (!g7) & (!g9) & (g18)) + ((!shiftx2x) & (!shiftx3x) & (!g6) & (!g7) & (g9) & (g18)) + ((!shiftx2x) & (!shiftx3x) & (!g6) & (g7) & (!g9) & (g18)) + ((!shiftx2x) & (!shiftx3x) & (!g6) & (g7) & (g9) & (g18)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (!g7) & (!g9) & (g18)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (!g7) & (g9) & (g18)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (g7) & (!g9) & (g18)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (g7) & (g9) & (g18)) + ((!shiftx2x) & (shiftx3x) & (!g6) & (g7) & (!g9) & (!g18)) + ((!shiftx2x) & (shiftx3x) & (!g6) & (g7) & (!g9) & (g18)) + ((!shiftx2x) & (shiftx3x) & (!g6) & (g7) & (g9) & (!g18)) + ((!shiftx2x) & (shiftx3x) & (!g6) & (g7) & (g9) & (g18)) + ((!shiftx2x) & (shiftx3x) & (g6) & (g7) & (!g9) & (!g18)) + ((!shiftx2x) & (shiftx3x) & (g6) & (g7) & (!g9) & (g18)) + ((!shiftx2x) & (shiftx3x) & (g6) & (g7) & (g9) & (!g18)) + ((!shiftx2x) & (shiftx3x) & (g6) & (g7) & (g9) & (g18)) + ((shiftx2x) & (!shiftx3x) & (g6) & (!g7) & (!g9) & (!g18)) + ((shiftx2x) & (!shiftx3x) & (g6) & (!g7) & (!g9) & (g18)) + ((shiftx2x) & (!shiftx3x) & (g6) & (!g7) & (g9) & (!g18)) + ((shiftx2x) & (!shiftx3x) & (g6) & (!g7) & (g9) & (g18)) + ((shiftx2x) & (!shiftx3x) & (g6) & (g7) & (!g9) & (!g18)) + ((shiftx2x) & (!shiftx3x) & (g6) & (g7) & (!g9) & (g18)) + ((shiftx2x) & (!shiftx3x) & (g6) & (g7) & (g9) & (!g18)) + ((shiftx2x) & (!shiftx3x) & (g6) & (g7) & (g9) & (g18)) + ((shiftx2x) & (shiftx3x) & (!g6) & (!g7) & (g9) & (!g18)) + ((shiftx2x) & (shiftx3x) & (!g6) & (!g7) & (g9) & (g18)) + ((shiftx2x) & (shiftx3x) & (!g6) & (g7) & (g9) & (!g18)) + ((shiftx2x) & (shiftx3x) & (!g6) & (g7) & (g9) & (g18)) + ((shiftx2x) & (shiftx3x) & (g6) & (!g7) & (g9) & (!g18)) + ((shiftx2x) & (shiftx3x) & (g6) & (!g7) & (g9) & (g18)) + ((shiftx2x) & (shiftx3x) & (g6) & (g7) & (g9) & (!g18)) + ((shiftx2x) & (shiftx3x) & (g6) & (g7) & (g9) & (g18)));
	assign g176 = (((!shiftx2x) & (!shiftx3x) & (!g1) & (!g2) & (!g4) & (g8)) + ((!shiftx2x) & (!shiftx3x) & (!g1) & (!g2) & (g4) & (g8)) + ((!shiftx2x) & (!shiftx3x) & (!g1) & (g2) & (!g4) & (g8)) + ((!shiftx2x) & (!shiftx3x) & (!g1) & (g2) & (g4) & (g8)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (!g2) & (!g4) & (g8)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (!g2) & (g4) & (g8)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (g2) & (!g4) & (g8)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (g2) & (g4) & (g8)) + ((!shiftx2x) & (shiftx3x) & (!g1) & (g2) & (!g4) & (!g8)) + ((!shiftx2x) & (shiftx3x) & (!g1) & (g2) & (!g4) & (g8)) + ((!shiftx2x) & (shiftx3x) & (!g1) & (g2) & (g4) & (!g8)) + ((!shiftx2x) & (shiftx3x) & (!g1) & (g2) & (g4) & (g8)) + ((!shiftx2x) & (shiftx3x) & (g1) & (g2) & (!g4) & (!g8)) + ((!shiftx2x) & (shiftx3x) & (g1) & (g2) & (!g4) & (g8)) + ((!shiftx2x) & (shiftx3x) & (g1) & (g2) & (g4) & (!g8)) + ((!shiftx2x) & (shiftx3x) & (g1) & (g2) & (g4) & (g8)) + ((shiftx2x) & (!shiftx3x) & (g1) & (!g2) & (!g4) & (!g8)) + ((shiftx2x) & (!shiftx3x) & (g1) & (!g2) & (!g4) & (g8)) + ((shiftx2x) & (!shiftx3x) & (g1) & (!g2) & (g4) & (!g8)) + ((shiftx2x) & (!shiftx3x) & (g1) & (!g2) & (g4) & (g8)) + ((shiftx2x) & (!shiftx3x) & (g1) & (g2) & (!g4) & (!g8)) + ((shiftx2x) & (!shiftx3x) & (g1) & (g2) & (!g4) & (g8)) + ((shiftx2x) & (!shiftx3x) & (g1) & (g2) & (g4) & (!g8)) + ((shiftx2x) & (!shiftx3x) & (g1) & (g2) & (g4) & (g8)) + ((shiftx2x) & (shiftx3x) & (!g1) & (!g2) & (g4) & (!g8)) + ((shiftx2x) & (shiftx3x) & (!g1) & (!g2) & (g4) & (g8)) + ((shiftx2x) & (shiftx3x) & (!g1) & (g2) & (g4) & (!g8)) + ((shiftx2x) & (shiftx3x) & (!g1) & (g2) & (g4) & (g8)) + ((shiftx2x) & (shiftx3x) & (g1) & (!g2) & (g4) & (!g8)) + ((shiftx2x) & (shiftx3x) & (g1) & (!g2) & (g4) & (g8)) + ((shiftx2x) & (shiftx3x) & (g1) & (g2) & (g4) & (!g8)) + ((shiftx2x) & (shiftx3x) & (g1) & (g2) & (g4) & (g8)));
	assign g177 = (((!shiftx4x) & (!shiftx5x) & (!g173) & (g174) & (!g175) & (!g176)) + ((!shiftx4x) & (!shiftx5x) & (!g173) & (g174) & (!g175) & (g176)) + ((!shiftx4x) & (!shiftx5x) & (!g173) & (g174) & (g175) & (!g176)) + ((!shiftx4x) & (!shiftx5x) & (!g173) & (g174) & (g175) & (g176)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (g174) & (!g175) & (!g176)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (g174) & (!g175) & (g176)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (g174) & (g175) & (!g176)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (g174) & (g175) & (g176)) + ((!shiftx4x) & (shiftx5x) & (!g173) & (!g174) & (g175) & (!g176)) + ((!shiftx4x) & (shiftx5x) & (!g173) & (!g174) & (g175) & (g176)) + ((!shiftx4x) & (shiftx5x) & (!g173) & (g174) & (g175) & (!g176)) + ((!shiftx4x) & (shiftx5x) & (!g173) & (g174) & (g175) & (g176)) + ((!shiftx4x) & (shiftx5x) & (g173) & (!g174) & (g175) & (!g176)) + ((!shiftx4x) & (shiftx5x) & (g173) & (!g174) & (g175) & (g176)) + ((!shiftx4x) & (shiftx5x) & (g173) & (g174) & (g175) & (!g176)) + ((!shiftx4x) & (shiftx5x) & (g173) & (g174) & (g175) & (g176)) + ((shiftx4x) & (!shiftx5x) & (g173) & (!g174) & (!g175) & (!g176)) + ((shiftx4x) & (!shiftx5x) & (g173) & (!g174) & (!g175) & (g176)) + ((shiftx4x) & (!shiftx5x) & (g173) & (!g174) & (g175) & (!g176)) + ((shiftx4x) & (!shiftx5x) & (g173) & (!g174) & (g175) & (g176)) + ((shiftx4x) & (!shiftx5x) & (g173) & (g174) & (!g175) & (!g176)) + ((shiftx4x) & (!shiftx5x) & (g173) & (g174) & (!g175) & (g176)) + ((shiftx4x) & (!shiftx5x) & (g173) & (g174) & (g175) & (!g176)) + ((shiftx4x) & (!shiftx5x) & (g173) & (g174) & (g175) & (g176)) + ((shiftx4x) & (shiftx5x) & (!g173) & (!g174) & (!g175) & (g176)) + ((shiftx4x) & (shiftx5x) & (!g173) & (!g174) & (g175) & (g176)) + ((shiftx4x) & (shiftx5x) & (!g173) & (g174) & (!g175) & (g176)) + ((shiftx4x) & (shiftx5x) & (!g173) & (g174) & (g175) & (g176)) + ((shiftx4x) & (shiftx5x) & (g173) & (!g174) & (!g175) & (g176)) + ((shiftx4x) & (shiftx5x) & (g173) & (!g174) & (g175) & (g176)) + ((shiftx4x) & (shiftx5x) & (g173) & (g174) & (!g175) & (g176)) + ((shiftx4x) & (shiftx5x) & (g173) & (g174) & (g175) & (g176)));
	assign g178 = (((!shiftx2x) & (!shiftx3x) & (!g22) & (!g23) & (!g25) & (g29)) + ((!shiftx2x) & (!shiftx3x) & (!g22) & (!g23) & (g25) & (g29)) + ((!shiftx2x) & (!shiftx3x) & (!g22) & (g23) & (!g25) & (g29)) + ((!shiftx2x) & (!shiftx3x) & (!g22) & (g23) & (g25) & (g29)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (!g23) & (!g25) & (g29)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (!g23) & (g25) & (g29)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (g23) & (!g25) & (g29)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (g23) & (g25) & (g29)) + ((!shiftx2x) & (shiftx3x) & (!g22) & (g23) & (!g25) & (!g29)) + ((!shiftx2x) & (shiftx3x) & (!g22) & (g23) & (!g25) & (g29)) + ((!shiftx2x) & (shiftx3x) & (!g22) & (g23) & (g25) & (!g29)) + ((!shiftx2x) & (shiftx3x) & (!g22) & (g23) & (g25) & (g29)) + ((!shiftx2x) & (shiftx3x) & (g22) & (g23) & (!g25) & (!g29)) + ((!shiftx2x) & (shiftx3x) & (g22) & (g23) & (!g25) & (g29)) + ((!shiftx2x) & (shiftx3x) & (g22) & (g23) & (g25) & (!g29)) + ((!shiftx2x) & (shiftx3x) & (g22) & (g23) & (g25) & (g29)) + ((shiftx2x) & (!shiftx3x) & (g22) & (!g23) & (!g25) & (!g29)) + ((shiftx2x) & (!shiftx3x) & (g22) & (!g23) & (!g25) & (g29)) + ((shiftx2x) & (!shiftx3x) & (g22) & (!g23) & (g25) & (!g29)) + ((shiftx2x) & (!shiftx3x) & (g22) & (!g23) & (g25) & (g29)) + ((shiftx2x) & (!shiftx3x) & (g22) & (g23) & (!g25) & (!g29)) + ((shiftx2x) & (!shiftx3x) & (g22) & (g23) & (!g25) & (g29)) + ((shiftx2x) & (!shiftx3x) & (g22) & (g23) & (g25) & (!g29)) + ((shiftx2x) & (!shiftx3x) & (g22) & (g23) & (g25) & (g29)) + ((shiftx2x) & (shiftx3x) & (!g22) & (!g23) & (g25) & (!g29)) + ((shiftx2x) & (shiftx3x) & (!g22) & (!g23) & (g25) & (g29)) + ((shiftx2x) & (shiftx3x) & (!g22) & (g23) & (g25) & (!g29)) + ((shiftx2x) & (shiftx3x) & (!g22) & (g23) & (g25) & (g29)) + ((shiftx2x) & (shiftx3x) & (g22) & (!g23) & (g25) & (!g29)) + ((shiftx2x) & (shiftx3x) & (g22) & (!g23) & (g25) & (g29)) + ((shiftx2x) & (shiftx3x) & (g22) & (g23) & (g25) & (!g29)) + ((shiftx2x) & (shiftx3x) & (g22) & (g23) & (g25) & (g29)));
	assign g179 = (((!shiftx2x) & (!shiftx3x) & (!g27) & (!g28) & (!g30) & (g39)) + ((!shiftx2x) & (!shiftx3x) & (!g27) & (!g28) & (g30) & (g39)) + ((!shiftx2x) & (!shiftx3x) & (!g27) & (g28) & (!g30) & (g39)) + ((!shiftx2x) & (!shiftx3x) & (!g27) & (g28) & (g30) & (g39)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (!g28) & (!g30) & (g39)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (!g28) & (g30) & (g39)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (g28) & (!g30) & (g39)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (g28) & (g30) & (g39)) + ((!shiftx2x) & (shiftx3x) & (!g27) & (g28) & (!g30) & (!g39)) + ((!shiftx2x) & (shiftx3x) & (!g27) & (g28) & (!g30) & (g39)) + ((!shiftx2x) & (shiftx3x) & (!g27) & (g28) & (g30) & (!g39)) + ((!shiftx2x) & (shiftx3x) & (!g27) & (g28) & (g30) & (g39)) + ((!shiftx2x) & (shiftx3x) & (g27) & (g28) & (!g30) & (!g39)) + ((!shiftx2x) & (shiftx3x) & (g27) & (g28) & (!g30) & (g39)) + ((!shiftx2x) & (shiftx3x) & (g27) & (g28) & (g30) & (!g39)) + ((!shiftx2x) & (shiftx3x) & (g27) & (g28) & (g30) & (g39)) + ((shiftx2x) & (!shiftx3x) & (g27) & (!g28) & (!g30) & (!g39)) + ((shiftx2x) & (!shiftx3x) & (g27) & (!g28) & (!g30) & (g39)) + ((shiftx2x) & (!shiftx3x) & (g27) & (!g28) & (g30) & (!g39)) + ((shiftx2x) & (!shiftx3x) & (g27) & (!g28) & (g30) & (g39)) + ((shiftx2x) & (!shiftx3x) & (g27) & (g28) & (!g30) & (!g39)) + ((shiftx2x) & (!shiftx3x) & (g27) & (g28) & (!g30) & (g39)) + ((shiftx2x) & (!shiftx3x) & (g27) & (g28) & (g30) & (!g39)) + ((shiftx2x) & (!shiftx3x) & (g27) & (g28) & (g30) & (g39)) + ((shiftx2x) & (shiftx3x) & (!g27) & (!g28) & (g30) & (!g39)) + ((shiftx2x) & (shiftx3x) & (!g27) & (!g28) & (g30) & (g39)) + ((shiftx2x) & (shiftx3x) & (!g27) & (g28) & (g30) & (!g39)) + ((shiftx2x) & (shiftx3x) & (!g27) & (g28) & (g30) & (g39)) + ((shiftx2x) & (shiftx3x) & (g27) & (!g28) & (g30) & (!g39)) + ((shiftx2x) & (shiftx3x) & (g27) & (!g28) & (g30) & (g39)) + ((shiftx2x) & (shiftx3x) & (g27) & (g28) & (g30) & (!g39)) + ((shiftx2x) & (shiftx3x) & (g27) & (g28) & (g30) & (g39)));
	assign g180 = (((!shiftx2x) & (!shiftx3x) & (g3) & (!g32) & (!g33) & (!g35)) + ((!shiftx2x) & (!shiftx3x) & (g3) & (!g32) & (!g33) & (g35)) + ((!shiftx2x) & (!shiftx3x) & (g3) & (!g32) & (g33) & (!g35)) + ((!shiftx2x) & (!shiftx3x) & (g3) & (!g32) & (g33) & (g35)) + ((!shiftx2x) & (!shiftx3x) & (g3) & (g32) & (!g33) & (!g35)) + ((!shiftx2x) & (!shiftx3x) & (g3) & (g32) & (!g33) & (g35)) + ((!shiftx2x) & (!shiftx3x) & (g3) & (g32) & (g33) & (!g35)) + ((!shiftx2x) & (!shiftx3x) & (g3) & (g32) & (g33) & (g35)) + ((!shiftx2x) & (shiftx3x) & (!g3) & (!g32) & (g33) & (!g35)) + ((!shiftx2x) & (shiftx3x) & (!g3) & (!g32) & (g33) & (g35)) + ((!shiftx2x) & (shiftx3x) & (!g3) & (g32) & (g33) & (!g35)) + ((!shiftx2x) & (shiftx3x) & (!g3) & (g32) & (g33) & (g35)) + ((!shiftx2x) & (shiftx3x) & (g3) & (!g32) & (g33) & (!g35)) + ((!shiftx2x) & (shiftx3x) & (g3) & (!g32) & (g33) & (g35)) + ((!shiftx2x) & (shiftx3x) & (g3) & (g32) & (g33) & (!g35)) + ((!shiftx2x) & (shiftx3x) & (g3) & (g32) & (g33) & (g35)) + ((shiftx2x) & (!shiftx3x) & (!g3) & (g32) & (!g33) & (!g35)) + ((shiftx2x) & (!shiftx3x) & (!g3) & (g32) & (!g33) & (g35)) + ((shiftx2x) & (!shiftx3x) & (!g3) & (g32) & (g33) & (!g35)) + ((shiftx2x) & (!shiftx3x) & (!g3) & (g32) & (g33) & (g35)) + ((shiftx2x) & (!shiftx3x) & (g3) & (g32) & (!g33) & (!g35)) + ((shiftx2x) & (!shiftx3x) & (g3) & (g32) & (!g33) & (g35)) + ((shiftx2x) & (!shiftx3x) & (g3) & (g32) & (g33) & (!g35)) + ((shiftx2x) & (!shiftx3x) & (g3) & (g32) & (g33) & (g35)) + ((shiftx2x) & (shiftx3x) & (!g3) & (!g32) & (!g33) & (g35)) + ((shiftx2x) & (shiftx3x) & (!g3) & (!g32) & (g33) & (g35)) + ((shiftx2x) & (shiftx3x) & (!g3) & (g32) & (!g33) & (g35)) + ((shiftx2x) & (shiftx3x) & (!g3) & (g32) & (g33) & (g35)) + ((shiftx2x) & (shiftx3x) & (g3) & (!g32) & (!g33) & (g35)) + ((shiftx2x) & (shiftx3x) & (g3) & (!g32) & (g33) & (g35)) + ((shiftx2x) & (shiftx3x) & (g3) & (g32) & (!g33) & (g35)) + ((shiftx2x) & (shiftx3x) & (g3) & (g32) & (g33) & (g35)));
	assign g181 = (((!shiftx2x) & (!shiftx3x) & (g34) & (!g37) & (!g38) & (!g40)) + ((!shiftx2x) & (!shiftx3x) & (g34) & (!g37) & (!g38) & (g40)) + ((!shiftx2x) & (!shiftx3x) & (g34) & (!g37) & (g38) & (!g40)) + ((!shiftx2x) & (!shiftx3x) & (g34) & (!g37) & (g38) & (g40)) + ((!shiftx2x) & (!shiftx3x) & (g34) & (g37) & (!g38) & (!g40)) + ((!shiftx2x) & (!shiftx3x) & (g34) & (g37) & (!g38) & (g40)) + ((!shiftx2x) & (!shiftx3x) & (g34) & (g37) & (g38) & (!g40)) + ((!shiftx2x) & (!shiftx3x) & (g34) & (g37) & (g38) & (g40)) + ((!shiftx2x) & (shiftx3x) & (!g34) & (!g37) & (g38) & (!g40)) + ((!shiftx2x) & (shiftx3x) & (!g34) & (!g37) & (g38) & (g40)) + ((!shiftx2x) & (shiftx3x) & (!g34) & (g37) & (g38) & (!g40)) + ((!shiftx2x) & (shiftx3x) & (!g34) & (g37) & (g38) & (g40)) + ((!shiftx2x) & (shiftx3x) & (g34) & (!g37) & (g38) & (!g40)) + ((!shiftx2x) & (shiftx3x) & (g34) & (!g37) & (g38) & (g40)) + ((!shiftx2x) & (shiftx3x) & (g34) & (g37) & (g38) & (!g40)) + ((!shiftx2x) & (shiftx3x) & (g34) & (g37) & (g38) & (g40)) + ((shiftx2x) & (!shiftx3x) & (!g34) & (g37) & (!g38) & (!g40)) + ((shiftx2x) & (!shiftx3x) & (!g34) & (g37) & (!g38) & (g40)) + ((shiftx2x) & (!shiftx3x) & (!g34) & (g37) & (g38) & (!g40)) + ((shiftx2x) & (!shiftx3x) & (!g34) & (g37) & (g38) & (g40)) + ((shiftx2x) & (!shiftx3x) & (g34) & (g37) & (!g38) & (!g40)) + ((shiftx2x) & (!shiftx3x) & (g34) & (g37) & (!g38) & (g40)) + ((shiftx2x) & (!shiftx3x) & (g34) & (g37) & (g38) & (!g40)) + ((shiftx2x) & (!shiftx3x) & (g34) & (g37) & (g38) & (g40)) + ((shiftx2x) & (shiftx3x) & (!g34) & (!g37) & (!g38) & (g40)) + ((shiftx2x) & (shiftx3x) & (!g34) & (!g37) & (g38) & (g40)) + ((shiftx2x) & (shiftx3x) & (!g34) & (g37) & (!g38) & (g40)) + ((shiftx2x) & (shiftx3x) & (!g34) & (g37) & (g38) & (g40)) + ((shiftx2x) & (shiftx3x) & (g34) & (!g37) & (!g38) & (g40)) + ((shiftx2x) & (shiftx3x) & (g34) & (!g37) & (g38) & (g40)) + ((shiftx2x) & (shiftx3x) & (g34) & (g37) & (!g38) & (g40)) + ((shiftx2x) & (shiftx3x) & (g34) & (g37) & (g38) & (g40)));
	assign g182 = (((!shiftx4x) & (!shiftx5x) & (!g178) & (!g179) & (g180) & (!g181)) + ((!shiftx4x) & (!shiftx5x) & (!g178) & (!g179) & (g180) & (g181)) + ((!shiftx4x) & (!shiftx5x) & (!g178) & (g179) & (g180) & (!g181)) + ((!shiftx4x) & (!shiftx5x) & (!g178) & (g179) & (g180) & (g181)) + ((!shiftx4x) & (!shiftx5x) & (g178) & (!g179) & (g180) & (!g181)) + ((!shiftx4x) & (!shiftx5x) & (g178) & (!g179) & (g180) & (g181)) + ((!shiftx4x) & (!shiftx5x) & (g178) & (g179) & (g180) & (!g181)) + ((!shiftx4x) & (!shiftx5x) & (g178) & (g179) & (g180) & (g181)) + ((!shiftx4x) & (shiftx5x) & (!g178) & (g179) & (!g180) & (!g181)) + ((!shiftx4x) & (shiftx5x) & (!g178) & (g179) & (!g180) & (g181)) + ((!shiftx4x) & (shiftx5x) & (!g178) & (g179) & (g180) & (!g181)) + ((!shiftx4x) & (shiftx5x) & (!g178) & (g179) & (g180) & (g181)) + ((!shiftx4x) & (shiftx5x) & (g178) & (g179) & (!g180) & (!g181)) + ((!shiftx4x) & (shiftx5x) & (g178) & (g179) & (!g180) & (g181)) + ((!shiftx4x) & (shiftx5x) & (g178) & (g179) & (g180) & (!g181)) + ((!shiftx4x) & (shiftx5x) & (g178) & (g179) & (g180) & (g181)) + ((shiftx4x) & (!shiftx5x) & (!g178) & (!g179) & (!g180) & (g181)) + ((shiftx4x) & (!shiftx5x) & (!g178) & (!g179) & (g180) & (g181)) + ((shiftx4x) & (!shiftx5x) & (!g178) & (g179) & (!g180) & (g181)) + ((shiftx4x) & (!shiftx5x) & (!g178) & (g179) & (g180) & (g181)) + ((shiftx4x) & (!shiftx5x) & (g178) & (!g179) & (!g180) & (g181)) + ((shiftx4x) & (!shiftx5x) & (g178) & (!g179) & (g180) & (g181)) + ((shiftx4x) & (!shiftx5x) & (g178) & (g179) & (!g180) & (g181)) + ((shiftx4x) & (!shiftx5x) & (g178) & (g179) & (g180) & (g181)) + ((shiftx4x) & (shiftx5x) & (g178) & (!g179) & (!g180) & (!g181)) + ((shiftx4x) & (shiftx5x) & (g178) & (!g179) & (!g180) & (g181)) + ((shiftx4x) & (shiftx5x) & (g178) & (!g179) & (g180) & (!g181)) + ((shiftx4x) & (shiftx5x) & (g178) & (!g179) & (g180) & (g181)) + ((shiftx4x) & (shiftx5x) & (g178) & (g179) & (!g180) & (!g181)) + ((shiftx4x) & (shiftx5x) & (g178) & (g179) & (!g180) & (g181)) + ((shiftx4x) & (shiftx5x) & (g178) & (g179) & (g180) & (!g181)) + ((shiftx4x) & (shiftx5x) & (g178) & (g179) & (g180) & (g181)));
	assign resultx4x = (((!sk[54]) & (shiftx6x) & (!g177) & (!g182)) + ((!sk[54]) & (shiftx6x) & (!g177) & (g182)) + ((!sk[54]) & (shiftx6x) & (g177) & (!g182)) + ((!sk[54]) & (shiftx6x) & (g177) & (g182)) + ((sk[54]) & (!shiftx6x) & (!g177) & (g182)) + ((sk[54]) & (!shiftx6x) & (g177) & (g182)) + ((sk[54]) & (shiftx6x) & (g177) & (!g182)) + ((sk[54]) & (shiftx6x) & (g177) & (g182)));
	assign g184 = (((!shiftx2x) & (!shiftx3x) & (g46) & (!g54) & (!g55) & (!g57)) + ((!shiftx2x) & (!shiftx3x) & (g46) & (!g54) & (!g55) & (g57)) + ((!shiftx2x) & (!shiftx3x) & (g46) & (!g54) & (g55) & (!g57)) + ((!shiftx2x) & (!shiftx3x) & (g46) & (!g54) & (g55) & (g57)) + ((!shiftx2x) & (!shiftx3x) & (g46) & (g54) & (!g55) & (!g57)) + ((!shiftx2x) & (!shiftx3x) & (g46) & (g54) & (!g55) & (g57)) + ((!shiftx2x) & (!shiftx3x) & (g46) & (g54) & (g55) & (!g57)) + ((!shiftx2x) & (!shiftx3x) & (g46) & (g54) & (g55) & (g57)) + ((!shiftx2x) & (shiftx3x) & (!g46) & (!g54) & (g55) & (!g57)) + ((!shiftx2x) & (shiftx3x) & (!g46) & (!g54) & (g55) & (g57)) + ((!shiftx2x) & (shiftx3x) & (!g46) & (g54) & (g55) & (!g57)) + ((!shiftx2x) & (shiftx3x) & (!g46) & (g54) & (g55) & (g57)) + ((!shiftx2x) & (shiftx3x) & (g46) & (!g54) & (g55) & (!g57)) + ((!shiftx2x) & (shiftx3x) & (g46) & (!g54) & (g55) & (g57)) + ((!shiftx2x) & (shiftx3x) & (g46) & (g54) & (g55) & (!g57)) + ((!shiftx2x) & (shiftx3x) & (g46) & (g54) & (g55) & (g57)) + ((shiftx2x) & (!shiftx3x) & (!g46) & (g54) & (!g55) & (!g57)) + ((shiftx2x) & (!shiftx3x) & (!g46) & (g54) & (!g55) & (g57)) + ((shiftx2x) & (!shiftx3x) & (!g46) & (g54) & (g55) & (!g57)) + ((shiftx2x) & (!shiftx3x) & (!g46) & (g54) & (g55) & (g57)) + ((shiftx2x) & (!shiftx3x) & (g46) & (g54) & (!g55) & (!g57)) + ((shiftx2x) & (!shiftx3x) & (g46) & (g54) & (!g55) & (g57)) + ((shiftx2x) & (!shiftx3x) & (g46) & (g54) & (g55) & (!g57)) + ((shiftx2x) & (!shiftx3x) & (g46) & (g54) & (g55) & (g57)) + ((shiftx2x) & (shiftx3x) & (!g46) & (!g54) & (!g55) & (g57)) + ((shiftx2x) & (shiftx3x) & (!g46) & (!g54) & (g55) & (g57)) + ((shiftx2x) & (shiftx3x) & (!g46) & (g54) & (!g55) & (g57)) + ((shiftx2x) & (shiftx3x) & (!g46) & (g54) & (g55) & (g57)) + ((shiftx2x) & (shiftx3x) & (g46) & (!g54) & (!g55) & (g57)) + ((shiftx2x) & (shiftx3x) & (g46) & (!g54) & (g55) & (g57)) + ((shiftx2x) & (shiftx3x) & (g46) & (g54) & (!g55) & (g57)) + ((shiftx2x) & (shiftx3x) & (g46) & (g54) & (g55) & (g57)));
	assign g185 = (((!shiftx2x) & (!shiftx3x) & (!g44) & (!g45) & (!g47) & (g67)) + ((!shiftx2x) & (!shiftx3x) & (!g44) & (!g45) & (g47) & (g67)) + ((!shiftx2x) & (!shiftx3x) & (!g44) & (g45) & (!g47) & (g67)) + ((!shiftx2x) & (!shiftx3x) & (!g44) & (g45) & (g47) & (g67)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (!g45) & (!g47) & (g67)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (!g45) & (g47) & (g67)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (g45) & (!g47) & (g67)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (g45) & (g47) & (g67)) + ((!shiftx2x) & (shiftx3x) & (!g44) & (g45) & (!g47) & (!g67)) + ((!shiftx2x) & (shiftx3x) & (!g44) & (g45) & (!g47) & (g67)) + ((!shiftx2x) & (shiftx3x) & (!g44) & (g45) & (g47) & (!g67)) + ((!shiftx2x) & (shiftx3x) & (!g44) & (g45) & (g47) & (g67)) + ((!shiftx2x) & (shiftx3x) & (g44) & (g45) & (!g47) & (!g67)) + ((!shiftx2x) & (shiftx3x) & (g44) & (g45) & (!g47) & (g67)) + ((!shiftx2x) & (shiftx3x) & (g44) & (g45) & (g47) & (!g67)) + ((!shiftx2x) & (shiftx3x) & (g44) & (g45) & (g47) & (g67)) + ((shiftx2x) & (!shiftx3x) & (g44) & (!g45) & (!g47) & (!g67)) + ((shiftx2x) & (!shiftx3x) & (g44) & (!g45) & (!g47) & (g67)) + ((shiftx2x) & (!shiftx3x) & (g44) & (!g45) & (g47) & (!g67)) + ((shiftx2x) & (!shiftx3x) & (g44) & (!g45) & (g47) & (g67)) + ((shiftx2x) & (!shiftx3x) & (g44) & (g45) & (!g47) & (!g67)) + ((shiftx2x) & (!shiftx3x) & (g44) & (g45) & (!g47) & (g67)) + ((shiftx2x) & (!shiftx3x) & (g44) & (g45) & (g47) & (!g67)) + ((shiftx2x) & (!shiftx3x) & (g44) & (g45) & (g47) & (g67)) + ((shiftx2x) & (shiftx3x) & (!g44) & (!g45) & (g47) & (!g67)) + ((shiftx2x) & (shiftx3x) & (!g44) & (!g45) & (g47) & (g67)) + ((shiftx2x) & (shiftx3x) & (!g44) & (g45) & (g47) & (!g67)) + ((shiftx2x) & (shiftx3x) & (!g44) & (g45) & (g47) & (g67)) + ((shiftx2x) & (shiftx3x) & (g44) & (!g45) & (g47) & (!g67)) + ((shiftx2x) & (shiftx3x) & (g44) & (!g45) & (g47) & (g67)) + ((shiftx2x) & (shiftx3x) & (g44) & (g45) & (g47) & (!g67)) + ((shiftx2x) & (shiftx3x) & (g44) & (g45) & (g47) & (g67)));
	assign g186 = (((!shiftx2x) & (!shiftx3x) & (g56) & (!g59) & (!g60) & (!g62)) + ((!shiftx2x) & (!shiftx3x) & (g56) & (!g59) & (!g60) & (g62)) + ((!shiftx2x) & (!shiftx3x) & (g56) & (!g59) & (g60) & (!g62)) + ((!shiftx2x) & (!shiftx3x) & (g56) & (!g59) & (g60) & (g62)) + ((!shiftx2x) & (!shiftx3x) & (g56) & (g59) & (!g60) & (!g62)) + ((!shiftx2x) & (!shiftx3x) & (g56) & (g59) & (!g60) & (g62)) + ((!shiftx2x) & (!shiftx3x) & (g56) & (g59) & (g60) & (!g62)) + ((!shiftx2x) & (!shiftx3x) & (g56) & (g59) & (g60) & (g62)) + ((!shiftx2x) & (shiftx3x) & (!g56) & (!g59) & (g60) & (!g62)) + ((!shiftx2x) & (shiftx3x) & (!g56) & (!g59) & (g60) & (g62)) + ((!shiftx2x) & (shiftx3x) & (!g56) & (g59) & (g60) & (!g62)) + ((!shiftx2x) & (shiftx3x) & (!g56) & (g59) & (g60) & (g62)) + ((!shiftx2x) & (shiftx3x) & (g56) & (!g59) & (g60) & (!g62)) + ((!shiftx2x) & (shiftx3x) & (g56) & (!g59) & (g60) & (g62)) + ((!shiftx2x) & (shiftx3x) & (g56) & (g59) & (g60) & (!g62)) + ((!shiftx2x) & (shiftx3x) & (g56) & (g59) & (g60) & (g62)) + ((shiftx2x) & (!shiftx3x) & (!g56) & (g59) & (!g60) & (!g62)) + ((shiftx2x) & (!shiftx3x) & (!g56) & (g59) & (!g60) & (g62)) + ((shiftx2x) & (!shiftx3x) & (!g56) & (g59) & (g60) & (!g62)) + ((shiftx2x) & (!shiftx3x) & (!g56) & (g59) & (g60) & (g62)) + ((shiftx2x) & (!shiftx3x) & (g56) & (g59) & (!g60) & (!g62)) + ((shiftx2x) & (!shiftx3x) & (g56) & (g59) & (!g60) & (g62)) + ((shiftx2x) & (!shiftx3x) & (g56) & (g59) & (g60) & (!g62)) + ((shiftx2x) & (!shiftx3x) & (g56) & (g59) & (g60) & (g62)) + ((shiftx2x) & (shiftx3x) & (!g56) & (!g59) & (!g60) & (g62)) + ((shiftx2x) & (shiftx3x) & (!g56) & (!g59) & (g60) & (g62)) + ((shiftx2x) & (shiftx3x) & (!g56) & (g59) & (!g60) & (g62)) + ((shiftx2x) & (shiftx3x) & (!g56) & (g59) & (g60) & (g62)) + ((shiftx2x) & (shiftx3x) & (g56) & (!g59) & (!g60) & (g62)) + ((shiftx2x) & (shiftx3x) & (g56) & (!g59) & (g60) & (g62)) + ((shiftx2x) & (shiftx3x) & (g56) & (g59) & (!g60) & (g62)) + ((shiftx2x) & (shiftx3x) & (g56) & (g59) & (g60) & (g62)));
	assign g187 = (((!shiftx2x) & (!shiftx3x) & (!g49) & (!g50) & (!g52) & (g61)) + ((!shiftx2x) & (!shiftx3x) & (!g49) & (!g50) & (g52) & (g61)) + ((!shiftx2x) & (!shiftx3x) & (!g49) & (g50) & (!g52) & (g61)) + ((!shiftx2x) & (!shiftx3x) & (!g49) & (g50) & (g52) & (g61)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (!g50) & (!g52) & (g61)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (!g50) & (g52) & (g61)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (g50) & (!g52) & (g61)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (g50) & (g52) & (g61)) + ((!shiftx2x) & (shiftx3x) & (!g49) & (g50) & (!g52) & (!g61)) + ((!shiftx2x) & (shiftx3x) & (!g49) & (g50) & (!g52) & (g61)) + ((!shiftx2x) & (shiftx3x) & (!g49) & (g50) & (g52) & (!g61)) + ((!shiftx2x) & (shiftx3x) & (!g49) & (g50) & (g52) & (g61)) + ((!shiftx2x) & (shiftx3x) & (g49) & (g50) & (!g52) & (!g61)) + ((!shiftx2x) & (shiftx3x) & (g49) & (g50) & (!g52) & (g61)) + ((!shiftx2x) & (shiftx3x) & (g49) & (g50) & (g52) & (!g61)) + ((!shiftx2x) & (shiftx3x) & (g49) & (g50) & (g52) & (g61)) + ((shiftx2x) & (!shiftx3x) & (g49) & (!g50) & (!g52) & (!g61)) + ((shiftx2x) & (!shiftx3x) & (g49) & (!g50) & (!g52) & (g61)) + ((shiftx2x) & (!shiftx3x) & (g49) & (!g50) & (g52) & (!g61)) + ((shiftx2x) & (!shiftx3x) & (g49) & (!g50) & (g52) & (g61)) + ((shiftx2x) & (!shiftx3x) & (g49) & (g50) & (!g52) & (!g61)) + ((shiftx2x) & (!shiftx3x) & (g49) & (g50) & (!g52) & (g61)) + ((shiftx2x) & (!shiftx3x) & (g49) & (g50) & (g52) & (!g61)) + ((shiftx2x) & (!shiftx3x) & (g49) & (g50) & (g52) & (g61)) + ((shiftx2x) & (shiftx3x) & (!g49) & (!g50) & (g52) & (!g61)) + ((shiftx2x) & (shiftx3x) & (!g49) & (!g50) & (g52) & (g61)) + ((shiftx2x) & (shiftx3x) & (!g49) & (g50) & (g52) & (!g61)) + ((shiftx2x) & (shiftx3x) & (!g49) & (g50) & (g52) & (g61)) + ((shiftx2x) & (shiftx3x) & (g49) & (!g50) & (g52) & (!g61)) + ((shiftx2x) & (shiftx3x) & (g49) & (!g50) & (g52) & (g61)) + ((shiftx2x) & (shiftx3x) & (g49) & (g50) & (g52) & (!g61)) + ((shiftx2x) & (shiftx3x) & (g49) & (g50) & (g52) & (g61)));
	assign g188 = (((!shiftx4x) & (!shiftx5x) & (!g184) & (g185) & (!g186) & (!g187)) + ((!shiftx4x) & (!shiftx5x) & (!g184) & (g185) & (!g186) & (g187)) + ((!shiftx4x) & (!shiftx5x) & (!g184) & (g185) & (g186) & (!g187)) + ((!shiftx4x) & (!shiftx5x) & (!g184) & (g185) & (g186) & (g187)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (g185) & (!g186) & (!g187)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (g185) & (!g186) & (g187)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (g185) & (g186) & (!g187)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (g185) & (g186) & (g187)) + ((!shiftx4x) & (shiftx5x) & (!g184) & (!g185) & (g186) & (!g187)) + ((!shiftx4x) & (shiftx5x) & (!g184) & (!g185) & (g186) & (g187)) + ((!shiftx4x) & (shiftx5x) & (!g184) & (g185) & (g186) & (!g187)) + ((!shiftx4x) & (shiftx5x) & (!g184) & (g185) & (g186) & (g187)) + ((!shiftx4x) & (shiftx5x) & (g184) & (!g185) & (g186) & (!g187)) + ((!shiftx4x) & (shiftx5x) & (g184) & (!g185) & (g186) & (g187)) + ((!shiftx4x) & (shiftx5x) & (g184) & (g185) & (g186) & (!g187)) + ((!shiftx4x) & (shiftx5x) & (g184) & (g185) & (g186) & (g187)) + ((shiftx4x) & (!shiftx5x) & (g184) & (!g185) & (!g186) & (!g187)) + ((shiftx4x) & (!shiftx5x) & (g184) & (!g185) & (!g186) & (g187)) + ((shiftx4x) & (!shiftx5x) & (g184) & (!g185) & (g186) & (!g187)) + ((shiftx4x) & (!shiftx5x) & (g184) & (!g185) & (g186) & (g187)) + ((shiftx4x) & (!shiftx5x) & (g184) & (g185) & (!g186) & (!g187)) + ((shiftx4x) & (!shiftx5x) & (g184) & (g185) & (!g186) & (g187)) + ((shiftx4x) & (!shiftx5x) & (g184) & (g185) & (g186) & (!g187)) + ((shiftx4x) & (!shiftx5x) & (g184) & (g185) & (g186) & (g187)) + ((shiftx4x) & (shiftx5x) & (!g184) & (!g185) & (!g186) & (g187)) + ((shiftx4x) & (shiftx5x) & (!g184) & (!g185) & (g186) & (g187)) + ((shiftx4x) & (shiftx5x) & (!g184) & (g185) & (!g186) & (g187)) + ((shiftx4x) & (shiftx5x) & (!g184) & (g185) & (g186) & (g187)) + ((shiftx4x) & (shiftx5x) & (g184) & (!g185) & (!g186) & (g187)) + ((shiftx4x) & (shiftx5x) & (g184) & (!g185) & (g186) & (g187)) + ((shiftx4x) & (shiftx5x) & (g184) & (g185) & (!g186) & (g187)) + ((shiftx4x) & (shiftx5x) & (g184) & (g185) & (g186) & (g187)));
	assign g189 = (((!shiftx2x) & (!shiftx3x) & (!g65) & (!g66) & (!g68) & (g72)) + ((!shiftx2x) & (!shiftx3x) & (!g65) & (!g66) & (g68) & (g72)) + ((!shiftx2x) & (!shiftx3x) & (!g65) & (g66) & (!g68) & (g72)) + ((!shiftx2x) & (!shiftx3x) & (!g65) & (g66) & (g68) & (g72)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (!g66) & (!g68) & (g72)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (!g66) & (g68) & (g72)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (g66) & (!g68) & (g72)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (g66) & (g68) & (g72)) + ((!shiftx2x) & (shiftx3x) & (!g65) & (g66) & (!g68) & (!g72)) + ((!shiftx2x) & (shiftx3x) & (!g65) & (g66) & (!g68) & (g72)) + ((!shiftx2x) & (shiftx3x) & (!g65) & (g66) & (g68) & (!g72)) + ((!shiftx2x) & (shiftx3x) & (!g65) & (g66) & (g68) & (g72)) + ((!shiftx2x) & (shiftx3x) & (g65) & (g66) & (!g68) & (!g72)) + ((!shiftx2x) & (shiftx3x) & (g65) & (g66) & (!g68) & (g72)) + ((!shiftx2x) & (shiftx3x) & (g65) & (g66) & (g68) & (!g72)) + ((!shiftx2x) & (shiftx3x) & (g65) & (g66) & (g68) & (g72)) + ((shiftx2x) & (!shiftx3x) & (g65) & (!g66) & (!g68) & (!g72)) + ((shiftx2x) & (!shiftx3x) & (g65) & (!g66) & (!g68) & (g72)) + ((shiftx2x) & (!shiftx3x) & (g65) & (!g66) & (g68) & (!g72)) + ((shiftx2x) & (!shiftx3x) & (g65) & (!g66) & (g68) & (g72)) + ((shiftx2x) & (!shiftx3x) & (g65) & (g66) & (!g68) & (!g72)) + ((shiftx2x) & (!shiftx3x) & (g65) & (g66) & (!g68) & (g72)) + ((shiftx2x) & (!shiftx3x) & (g65) & (g66) & (g68) & (!g72)) + ((shiftx2x) & (!shiftx3x) & (g65) & (g66) & (g68) & (g72)) + ((shiftx2x) & (shiftx3x) & (!g65) & (!g66) & (g68) & (!g72)) + ((shiftx2x) & (shiftx3x) & (!g65) & (!g66) & (g68) & (g72)) + ((shiftx2x) & (shiftx3x) & (!g65) & (g66) & (g68) & (!g72)) + ((shiftx2x) & (shiftx3x) & (!g65) & (g66) & (g68) & (g72)) + ((shiftx2x) & (shiftx3x) & (g65) & (!g66) & (g68) & (!g72)) + ((shiftx2x) & (shiftx3x) & (g65) & (!g66) & (g68) & (g72)) + ((shiftx2x) & (shiftx3x) & (g65) & (g66) & (g68) & (!g72)) + ((shiftx2x) & (shiftx3x) & (g65) & (g66) & (g68) & (g72)));
	assign g190 = (((!shiftx2x) & (!shiftx3x) & (!g70) & (!g71) & (!g73) & (g82)) + ((!shiftx2x) & (!shiftx3x) & (!g70) & (!g71) & (g73) & (g82)) + ((!shiftx2x) & (!shiftx3x) & (!g70) & (g71) & (!g73) & (g82)) + ((!shiftx2x) & (!shiftx3x) & (!g70) & (g71) & (g73) & (g82)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (!g71) & (!g73) & (g82)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (!g71) & (g73) & (g82)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (g71) & (!g73) & (g82)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (g71) & (g73) & (g82)) + ((!shiftx2x) & (shiftx3x) & (!g70) & (g71) & (!g73) & (!g82)) + ((!shiftx2x) & (shiftx3x) & (!g70) & (g71) & (!g73) & (g82)) + ((!shiftx2x) & (shiftx3x) & (!g70) & (g71) & (g73) & (!g82)) + ((!shiftx2x) & (shiftx3x) & (!g70) & (g71) & (g73) & (g82)) + ((!shiftx2x) & (shiftx3x) & (g70) & (g71) & (!g73) & (!g82)) + ((!shiftx2x) & (shiftx3x) & (g70) & (g71) & (!g73) & (g82)) + ((!shiftx2x) & (shiftx3x) & (g70) & (g71) & (g73) & (!g82)) + ((!shiftx2x) & (shiftx3x) & (g70) & (g71) & (g73) & (g82)) + ((shiftx2x) & (!shiftx3x) & (g70) & (!g71) & (!g73) & (!g82)) + ((shiftx2x) & (!shiftx3x) & (g70) & (!g71) & (!g73) & (g82)) + ((shiftx2x) & (!shiftx3x) & (g70) & (!g71) & (g73) & (!g82)) + ((shiftx2x) & (!shiftx3x) & (g70) & (!g71) & (g73) & (g82)) + ((shiftx2x) & (!shiftx3x) & (g70) & (g71) & (!g73) & (!g82)) + ((shiftx2x) & (!shiftx3x) & (g70) & (g71) & (!g73) & (g82)) + ((shiftx2x) & (!shiftx3x) & (g70) & (g71) & (g73) & (!g82)) + ((shiftx2x) & (!shiftx3x) & (g70) & (g71) & (g73) & (g82)) + ((shiftx2x) & (shiftx3x) & (!g70) & (!g71) & (g73) & (!g82)) + ((shiftx2x) & (shiftx3x) & (!g70) & (!g71) & (g73) & (g82)) + ((shiftx2x) & (shiftx3x) & (!g70) & (g71) & (g73) & (!g82)) + ((shiftx2x) & (shiftx3x) & (!g70) & (g71) & (g73) & (g82)) + ((shiftx2x) & (shiftx3x) & (g70) & (!g71) & (g73) & (!g82)) + ((shiftx2x) & (shiftx3x) & (g70) & (!g71) & (g73) & (g82)) + ((shiftx2x) & (shiftx3x) & (g70) & (g71) & (g73) & (!g82)) + ((shiftx2x) & (shiftx3x) & (g70) & (g71) & (g73) & (g82)));
	assign g191 = (((!shiftx2x) & (!shiftx3x) & (g51) & (!g75) & (!g76) & (!g78)) + ((!shiftx2x) & (!shiftx3x) & (g51) & (!g75) & (!g76) & (g78)) + ((!shiftx2x) & (!shiftx3x) & (g51) & (!g75) & (g76) & (!g78)) + ((!shiftx2x) & (!shiftx3x) & (g51) & (!g75) & (g76) & (g78)) + ((!shiftx2x) & (!shiftx3x) & (g51) & (g75) & (!g76) & (!g78)) + ((!shiftx2x) & (!shiftx3x) & (g51) & (g75) & (!g76) & (g78)) + ((!shiftx2x) & (!shiftx3x) & (g51) & (g75) & (g76) & (!g78)) + ((!shiftx2x) & (!shiftx3x) & (g51) & (g75) & (g76) & (g78)) + ((!shiftx2x) & (shiftx3x) & (!g51) & (!g75) & (g76) & (!g78)) + ((!shiftx2x) & (shiftx3x) & (!g51) & (!g75) & (g76) & (g78)) + ((!shiftx2x) & (shiftx3x) & (!g51) & (g75) & (g76) & (!g78)) + ((!shiftx2x) & (shiftx3x) & (!g51) & (g75) & (g76) & (g78)) + ((!shiftx2x) & (shiftx3x) & (g51) & (!g75) & (g76) & (!g78)) + ((!shiftx2x) & (shiftx3x) & (g51) & (!g75) & (g76) & (g78)) + ((!shiftx2x) & (shiftx3x) & (g51) & (g75) & (g76) & (!g78)) + ((!shiftx2x) & (shiftx3x) & (g51) & (g75) & (g76) & (g78)) + ((shiftx2x) & (!shiftx3x) & (!g51) & (g75) & (!g76) & (!g78)) + ((shiftx2x) & (!shiftx3x) & (!g51) & (g75) & (!g76) & (g78)) + ((shiftx2x) & (!shiftx3x) & (!g51) & (g75) & (g76) & (!g78)) + ((shiftx2x) & (!shiftx3x) & (!g51) & (g75) & (g76) & (g78)) + ((shiftx2x) & (!shiftx3x) & (g51) & (g75) & (!g76) & (!g78)) + ((shiftx2x) & (!shiftx3x) & (g51) & (g75) & (!g76) & (g78)) + ((shiftx2x) & (!shiftx3x) & (g51) & (g75) & (g76) & (!g78)) + ((shiftx2x) & (!shiftx3x) & (g51) & (g75) & (g76) & (g78)) + ((shiftx2x) & (shiftx3x) & (!g51) & (!g75) & (!g76) & (g78)) + ((shiftx2x) & (shiftx3x) & (!g51) & (!g75) & (g76) & (g78)) + ((shiftx2x) & (shiftx3x) & (!g51) & (g75) & (!g76) & (g78)) + ((shiftx2x) & (shiftx3x) & (!g51) & (g75) & (g76) & (g78)) + ((shiftx2x) & (shiftx3x) & (g51) & (!g75) & (!g76) & (g78)) + ((shiftx2x) & (shiftx3x) & (g51) & (!g75) & (g76) & (g78)) + ((shiftx2x) & (shiftx3x) & (g51) & (g75) & (!g76) & (g78)) + ((shiftx2x) & (shiftx3x) & (g51) & (g75) & (g76) & (g78)));
	assign g192 = (((!shiftx2x) & (!shiftx3x) & (g77) & (!g80) & (!g81) & (!g83)) + ((!shiftx2x) & (!shiftx3x) & (g77) & (!g80) & (!g81) & (g83)) + ((!shiftx2x) & (!shiftx3x) & (g77) & (!g80) & (g81) & (!g83)) + ((!shiftx2x) & (!shiftx3x) & (g77) & (!g80) & (g81) & (g83)) + ((!shiftx2x) & (!shiftx3x) & (g77) & (g80) & (!g81) & (!g83)) + ((!shiftx2x) & (!shiftx3x) & (g77) & (g80) & (!g81) & (g83)) + ((!shiftx2x) & (!shiftx3x) & (g77) & (g80) & (g81) & (!g83)) + ((!shiftx2x) & (!shiftx3x) & (g77) & (g80) & (g81) & (g83)) + ((!shiftx2x) & (shiftx3x) & (!g77) & (!g80) & (g81) & (!g83)) + ((!shiftx2x) & (shiftx3x) & (!g77) & (!g80) & (g81) & (g83)) + ((!shiftx2x) & (shiftx3x) & (!g77) & (g80) & (g81) & (!g83)) + ((!shiftx2x) & (shiftx3x) & (!g77) & (g80) & (g81) & (g83)) + ((!shiftx2x) & (shiftx3x) & (g77) & (!g80) & (g81) & (!g83)) + ((!shiftx2x) & (shiftx3x) & (g77) & (!g80) & (g81) & (g83)) + ((!shiftx2x) & (shiftx3x) & (g77) & (g80) & (g81) & (!g83)) + ((!shiftx2x) & (shiftx3x) & (g77) & (g80) & (g81) & (g83)) + ((shiftx2x) & (!shiftx3x) & (!g77) & (g80) & (!g81) & (!g83)) + ((shiftx2x) & (!shiftx3x) & (!g77) & (g80) & (!g81) & (g83)) + ((shiftx2x) & (!shiftx3x) & (!g77) & (g80) & (g81) & (!g83)) + ((shiftx2x) & (!shiftx3x) & (!g77) & (g80) & (g81) & (g83)) + ((shiftx2x) & (!shiftx3x) & (g77) & (g80) & (!g81) & (!g83)) + ((shiftx2x) & (!shiftx3x) & (g77) & (g80) & (!g81) & (g83)) + ((shiftx2x) & (!shiftx3x) & (g77) & (g80) & (g81) & (!g83)) + ((shiftx2x) & (!shiftx3x) & (g77) & (g80) & (g81) & (g83)) + ((shiftx2x) & (shiftx3x) & (!g77) & (!g80) & (!g81) & (g83)) + ((shiftx2x) & (shiftx3x) & (!g77) & (!g80) & (g81) & (g83)) + ((shiftx2x) & (shiftx3x) & (!g77) & (g80) & (!g81) & (g83)) + ((shiftx2x) & (shiftx3x) & (!g77) & (g80) & (g81) & (g83)) + ((shiftx2x) & (shiftx3x) & (g77) & (!g80) & (!g81) & (g83)) + ((shiftx2x) & (shiftx3x) & (g77) & (!g80) & (g81) & (g83)) + ((shiftx2x) & (shiftx3x) & (g77) & (g80) & (!g81) & (g83)) + ((shiftx2x) & (shiftx3x) & (g77) & (g80) & (g81) & (g83)));
	assign g193 = (((!shiftx4x) & (!shiftx5x) & (!g189) & (!g190) & (g191) & (!g192)) + ((!shiftx4x) & (!shiftx5x) & (!g189) & (!g190) & (g191) & (g192)) + ((!shiftx4x) & (!shiftx5x) & (!g189) & (g190) & (g191) & (!g192)) + ((!shiftx4x) & (!shiftx5x) & (!g189) & (g190) & (g191) & (g192)) + ((!shiftx4x) & (!shiftx5x) & (g189) & (!g190) & (g191) & (!g192)) + ((!shiftx4x) & (!shiftx5x) & (g189) & (!g190) & (g191) & (g192)) + ((!shiftx4x) & (!shiftx5x) & (g189) & (g190) & (g191) & (!g192)) + ((!shiftx4x) & (!shiftx5x) & (g189) & (g190) & (g191) & (g192)) + ((!shiftx4x) & (shiftx5x) & (!g189) & (g190) & (!g191) & (!g192)) + ((!shiftx4x) & (shiftx5x) & (!g189) & (g190) & (!g191) & (g192)) + ((!shiftx4x) & (shiftx5x) & (!g189) & (g190) & (g191) & (!g192)) + ((!shiftx4x) & (shiftx5x) & (!g189) & (g190) & (g191) & (g192)) + ((!shiftx4x) & (shiftx5x) & (g189) & (g190) & (!g191) & (!g192)) + ((!shiftx4x) & (shiftx5x) & (g189) & (g190) & (!g191) & (g192)) + ((!shiftx4x) & (shiftx5x) & (g189) & (g190) & (g191) & (!g192)) + ((!shiftx4x) & (shiftx5x) & (g189) & (g190) & (g191) & (g192)) + ((shiftx4x) & (!shiftx5x) & (!g189) & (!g190) & (!g191) & (g192)) + ((shiftx4x) & (!shiftx5x) & (!g189) & (!g190) & (g191) & (g192)) + ((shiftx4x) & (!shiftx5x) & (!g189) & (g190) & (!g191) & (g192)) + ((shiftx4x) & (!shiftx5x) & (!g189) & (g190) & (g191) & (g192)) + ((shiftx4x) & (!shiftx5x) & (g189) & (!g190) & (!g191) & (g192)) + ((shiftx4x) & (!shiftx5x) & (g189) & (!g190) & (g191) & (g192)) + ((shiftx4x) & (!shiftx5x) & (g189) & (g190) & (!g191) & (g192)) + ((shiftx4x) & (!shiftx5x) & (g189) & (g190) & (g191) & (g192)) + ((shiftx4x) & (shiftx5x) & (g189) & (!g190) & (!g191) & (!g192)) + ((shiftx4x) & (shiftx5x) & (g189) & (!g190) & (!g191) & (g192)) + ((shiftx4x) & (shiftx5x) & (g189) & (!g190) & (g191) & (!g192)) + ((shiftx4x) & (shiftx5x) & (g189) & (!g190) & (g191) & (g192)) + ((shiftx4x) & (shiftx5x) & (g189) & (g190) & (!g191) & (!g192)) + ((shiftx4x) & (shiftx5x) & (g189) & (g190) & (!g191) & (g192)) + ((shiftx4x) & (shiftx5x) & (g189) & (g190) & (g191) & (!g192)) + ((shiftx4x) & (shiftx5x) & (g189) & (g190) & (g191) & (g192)));
	assign resultx5x = (((!shiftx6x) & (!g188) & (sk[65]) & (g193)) + ((!shiftx6x) & (g188) & (sk[65]) & (g193)) + ((shiftx6x) & (!g188) & (!sk[65]) & (!g193)) + ((shiftx6x) & (!g188) & (!sk[65]) & (g193)) + ((shiftx6x) & (g188) & (!sk[65]) & (!g193)) + ((shiftx6x) & (g188) & (!sk[65]) & (g193)) + ((shiftx6x) & (g188) & (sk[65]) & (!g193)) + ((shiftx6x) & (g188) & (sk[65]) & (g193)));
	assign g195 = (((!shiftx2x) & (!shiftx3x) & (g89) & (!g97) & (!g98) & (!g100)) + ((!shiftx2x) & (!shiftx3x) & (g89) & (!g97) & (!g98) & (g100)) + ((!shiftx2x) & (!shiftx3x) & (g89) & (!g97) & (g98) & (!g100)) + ((!shiftx2x) & (!shiftx3x) & (g89) & (!g97) & (g98) & (g100)) + ((!shiftx2x) & (!shiftx3x) & (g89) & (g97) & (!g98) & (!g100)) + ((!shiftx2x) & (!shiftx3x) & (g89) & (g97) & (!g98) & (g100)) + ((!shiftx2x) & (!shiftx3x) & (g89) & (g97) & (g98) & (!g100)) + ((!shiftx2x) & (!shiftx3x) & (g89) & (g97) & (g98) & (g100)) + ((!shiftx2x) & (shiftx3x) & (!g89) & (!g97) & (g98) & (!g100)) + ((!shiftx2x) & (shiftx3x) & (!g89) & (!g97) & (g98) & (g100)) + ((!shiftx2x) & (shiftx3x) & (!g89) & (g97) & (g98) & (!g100)) + ((!shiftx2x) & (shiftx3x) & (!g89) & (g97) & (g98) & (g100)) + ((!shiftx2x) & (shiftx3x) & (g89) & (!g97) & (g98) & (!g100)) + ((!shiftx2x) & (shiftx3x) & (g89) & (!g97) & (g98) & (g100)) + ((!shiftx2x) & (shiftx3x) & (g89) & (g97) & (g98) & (!g100)) + ((!shiftx2x) & (shiftx3x) & (g89) & (g97) & (g98) & (g100)) + ((shiftx2x) & (!shiftx3x) & (!g89) & (g97) & (!g98) & (!g100)) + ((shiftx2x) & (!shiftx3x) & (!g89) & (g97) & (!g98) & (g100)) + ((shiftx2x) & (!shiftx3x) & (!g89) & (g97) & (g98) & (!g100)) + ((shiftx2x) & (!shiftx3x) & (!g89) & (g97) & (g98) & (g100)) + ((shiftx2x) & (!shiftx3x) & (g89) & (g97) & (!g98) & (!g100)) + ((shiftx2x) & (!shiftx3x) & (g89) & (g97) & (!g98) & (g100)) + ((shiftx2x) & (!shiftx3x) & (g89) & (g97) & (g98) & (!g100)) + ((shiftx2x) & (!shiftx3x) & (g89) & (g97) & (g98) & (g100)) + ((shiftx2x) & (shiftx3x) & (!g89) & (!g97) & (!g98) & (g100)) + ((shiftx2x) & (shiftx3x) & (!g89) & (!g97) & (g98) & (g100)) + ((shiftx2x) & (shiftx3x) & (!g89) & (g97) & (!g98) & (g100)) + ((shiftx2x) & (shiftx3x) & (!g89) & (g97) & (g98) & (g100)) + ((shiftx2x) & (shiftx3x) & (g89) & (!g97) & (!g98) & (g100)) + ((shiftx2x) & (shiftx3x) & (g89) & (!g97) & (g98) & (g100)) + ((shiftx2x) & (shiftx3x) & (g89) & (g97) & (!g98) & (g100)) + ((shiftx2x) & (shiftx3x) & (g89) & (g97) & (g98) & (g100)));
	assign g196 = (((!shiftx2x) & (!shiftx3x) & (!g87) & (!g88) & (!g90) & (g110)) + ((!shiftx2x) & (!shiftx3x) & (!g87) & (!g88) & (g90) & (g110)) + ((!shiftx2x) & (!shiftx3x) & (!g87) & (g88) & (!g90) & (g110)) + ((!shiftx2x) & (!shiftx3x) & (!g87) & (g88) & (g90) & (g110)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (!g88) & (!g90) & (g110)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (!g88) & (g90) & (g110)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (g88) & (!g90) & (g110)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (g88) & (g90) & (g110)) + ((!shiftx2x) & (shiftx3x) & (!g87) & (g88) & (!g90) & (!g110)) + ((!shiftx2x) & (shiftx3x) & (!g87) & (g88) & (!g90) & (g110)) + ((!shiftx2x) & (shiftx3x) & (!g87) & (g88) & (g90) & (!g110)) + ((!shiftx2x) & (shiftx3x) & (!g87) & (g88) & (g90) & (g110)) + ((!shiftx2x) & (shiftx3x) & (g87) & (g88) & (!g90) & (!g110)) + ((!shiftx2x) & (shiftx3x) & (g87) & (g88) & (!g90) & (g110)) + ((!shiftx2x) & (shiftx3x) & (g87) & (g88) & (g90) & (!g110)) + ((!shiftx2x) & (shiftx3x) & (g87) & (g88) & (g90) & (g110)) + ((shiftx2x) & (!shiftx3x) & (g87) & (!g88) & (!g90) & (!g110)) + ((shiftx2x) & (!shiftx3x) & (g87) & (!g88) & (!g90) & (g110)) + ((shiftx2x) & (!shiftx3x) & (g87) & (!g88) & (g90) & (!g110)) + ((shiftx2x) & (!shiftx3x) & (g87) & (!g88) & (g90) & (g110)) + ((shiftx2x) & (!shiftx3x) & (g87) & (g88) & (!g90) & (!g110)) + ((shiftx2x) & (!shiftx3x) & (g87) & (g88) & (!g90) & (g110)) + ((shiftx2x) & (!shiftx3x) & (g87) & (g88) & (g90) & (!g110)) + ((shiftx2x) & (!shiftx3x) & (g87) & (g88) & (g90) & (g110)) + ((shiftx2x) & (shiftx3x) & (!g87) & (!g88) & (g90) & (!g110)) + ((shiftx2x) & (shiftx3x) & (!g87) & (!g88) & (g90) & (g110)) + ((shiftx2x) & (shiftx3x) & (!g87) & (g88) & (g90) & (!g110)) + ((shiftx2x) & (shiftx3x) & (!g87) & (g88) & (g90) & (g110)) + ((shiftx2x) & (shiftx3x) & (g87) & (!g88) & (g90) & (!g110)) + ((shiftx2x) & (shiftx3x) & (g87) & (!g88) & (g90) & (g110)) + ((shiftx2x) & (shiftx3x) & (g87) & (g88) & (g90) & (!g110)) + ((shiftx2x) & (shiftx3x) & (g87) & (g88) & (g90) & (g110)));
	assign g197 = (((!shiftx2x) & (!shiftx3x) & (g99) & (!g102) & (!g103) & (!g105)) + ((!shiftx2x) & (!shiftx3x) & (g99) & (!g102) & (!g103) & (g105)) + ((!shiftx2x) & (!shiftx3x) & (g99) & (!g102) & (g103) & (!g105)) + ((!shiftx2x) & (!shiftx3x) & (g99) & (!g102) & (g103) & (g105)) + ((!shiftx2x) & (!shiftx3x) & (g99) & (g102) & (!g103) & (!g105)) + ((!shiftx2x) & (!shiftx3x) & (g99) & (g102) & (!g103) & (g105)) + ((!shiftx2x) & (!shiftx3x) & (g99) & (g102) & (g103) & (!g105)) + ((!shiftx2x) & (!shiftx3x) & (g99) & (g102) & (g103) & (g105)) + ((!shiftx2x) & (shiftx3x) & (!g99) & (!g102) & (g103) & (!g105)) + ((!shiftx2x) & (shiftx3x) & (!g99) & (!g102) & (g103) & (g105)) + ((!shiftx2x) & (shiftx3x) & (!g99) & (g102) & (g103) & (!g105)) + ((!shiftx2x) & (shiftx3x) & (!g99) & (g102) & (g103) & (g105)) + ((!shiftx2x) & (shiftx3x) & (g99) & (!g102) & (g103) & (!g105)) + ((!shiftx2x) & (shiftx3x) & (g99) & (!g102) & (g103) & (g105)) + ((!shiftx2x) & (shiftx3x) & (g99) & (g102) & (g103) & (!g105)) + ((!shiftx2x) & (shiftx3x) & (g99) & (g102) & (g103) & (g105)) + ((shiftx2x) & (!shiftx3x) & (!g99) & (g102) & (!g103) & (!g105)) + ((shiftx2x) & (!shiftx3x) & (!g99) & (g102) & (!g103) & (g105)) + ((shiftx2x) & (!shiftx3x) & (!g99) & (g102) & (g103) & (!g105)) + ((shiftx2x) & (!shiftx3x) & (!g99) & (g102) & (g103) & (g105)) + ((shiftx2x) & (!shiftx3x) & (g99) & (g102) & (!g103) & (!g105)) + ((shiftx2x) & (!shiftx3x) & (g99) & (g102) & (!g103) & (g105)) + ((shiftx2x) & (!shiftx3x) & (g99) & (g102) & (g103) & (!g105)) + ((shiftx2x) & (!shiftx3x) & (g99) & (g102) & (g103) & (g105)) + ((shiftx2x) & (shiftx3x) & (!g99) & (!g102) & (!g103) & (g105)) + ((shiftx2x) & (shiftx3x) & (!g99) & (!g102) & (g103) & (g105)) + ((shiftx2x) & (shiftx3x) & (!g99) & (g102) & (!g103) & (g105)) + ((shiftx2x) & (shiftx3x) & (!g99) & (g102) & (g103) & (g105)) + ((shiftx2x) & (shiftx3x) & (g99) & (!g102) & (!g103) & (g105)) + ((shiftx2x) & (shiftx3x) & (g99) & (!g102) & (g103) & (g105)) + ((shiftx2x) & (shiftx3x) & (g99) & (g102) & (!g103) & (g105)) + ((shiftx2x) & (shiftx3x) & (g99) & (g102) & (g103) & (g105)));
	assign g198 = (((!shiftx2x) & (!shiftx3x) & (!g92) & (!g93) & (!g95) & (g104)) + ((!shiftx2x) & (!shiftx3x) & (!g92) & (!g93) & (g95) & (g104)) + ((!shiftx2x) & (!shiftx3x) & (!g92) & (g93) & (!g95) & (g104)) + ((!shiftx2x) & (!shiftx3x) & (!g92) & (g93) & (g95) & (g104)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (!g93) & (!g95) & (g104)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (!g93) & (g95) & (g104)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (g93) & (!g95) & (g104)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (g93) & (g95) & (g104)) + ((!shiftx2x) & (shiftx3x) & (!g92) & (g93) & (!g95) & (!g104)) + ((!shiftx2x) & (shiftx3x) & (!g92) & (g93) & (!g95) & (g104)) + ((!shiftx2x) & (shiftx3x) & (!g92) & (g93) & (g95) & (!g104)) + ((!shiftx2x) & (shiftx3x) & (!g92) & (g93) & (g95) & (g104)) + ((!shiftx2x) & (shiftx3x) & (g92) & (g93) & (!g95) & (!g104)) + ((!shiftx2x) & (shiftx3x) & (g92) & (g93) & (!g95) & (g104)) + ((!shiftx2x) & (shiftx3x) & (g92) & (g93) & (g95) & (!g104)) + ((!shiftx2x) & (shiftx3x) & (g92) & (g93) & (g95) & (g104)) + ((shiftx2x) & (!shiftx3x) & (g92) & (!g93) & (!g95) & (!g104)) + ((shiftx2x) & (!shiftx3x) & (g92) & (!g93) & (!g95) & (g104)) + ((shiftx2x) & (!shiftx3x) & (g92) & (!g93) & (g95) & (!g104)) + ((shiftx2x) & (!shiftx3x) & (g92) & (!g93) & (g95) & (g104)) + ((shiftx2x) & (!shiftx3x) & (g92) & (g93) & (!g95) & (!g104)) + ((shiftx2x) & (!shiftx3x) & (g92) & (g93) & (!g95) & (g104)) + ((shiftx2x) & (!shiftx3x) & (g92) & (g93) & (g95) & (!g104)) + ((shiftx2x) & (!shiftx3x) & (g92) & (g93) & (g95) & (g104)) + ((shiftx2x) & (shiftx3x) & (!g92) & (!g93) & (g95) & (!g104)) + ((shiftx2x) & (shiftx3x) & (!g92) & (!g93) & (g95) & (g104)) + ((shiftx2x) & (shiftx3x) & (!g92) & (g93) & (g95) & (!g104)) + ((shiftx2x) & (shiftx3x) & (!g92) & (g93) & (g95) & (g104)) + ((shiftx2x) & (shiftx3x) & (g92) & (!g93) & (g95) & (!g104)) + ((shiftx2x) & (shiftx3x) & (g92) & (!g93) & (g95) & (g104)) + ((shiftx2x) & (shiftx3x) & (g92) & (g93) & (g95) & (!g104)) + ((shiftx2x) & (shiftx3x) & (g92) & (g93) & (g95) & (g104)));
	assign g199 = (((!shiftx4x) & (!shiftx5x) & (!g195) & (g196) & (!g197) & (!g198)) + ((!shiftx4x) & (!shiftx5x) & (!g195) & (g196) & (!g197) & (g198)) + ((!shiftx4x) & (!shiftx5x) & (!g195) & (g196) & (g197) & (!g198)) + ((!shiftx4x) & (!shiftx5x) & (!g195) & (g196) & (g197) & (g198)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (g196) & (!g197) & (!g198)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (g196) & (!g197) & (g198)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (g196) & (g197) & (!g198)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (g196) & (g197) & (g198)) + ((!shiftx4x) & (shiftx5x) & (!g195) & (!g196) & (g197) & (!g198)) + ((!shiftx4x) & (shiftx5x) & (!g195) & (!g196) & (g197) & (g198)) + ((!shiftx4x) & (shiftx5x) & (!g195) & (g196) & (g197) & (!g198)) + ((!shiftx4x) & (shiftx5x) & (!g195) & (g196) & (g197) & (g198)) + ((!shiftx4x) & (shiftx5x) & (g195) & (!g196) & (g197) & (!g198)) + ((!shiftx4x) & (shiftx5x) & (g195) & (!g196) & (g197) & (g198)) + ((!shiftx4x) & (shiftx5x) & (g195) & (g196) & (g197) & (!g198)) + ((!shiftx4x) & (shiftx5x) & (g195) & (g196) & (g197) & (g198)) + ((shiftx4x) & (!shiftx5x) & (g195) & (!g196) & (!g197) & (!g198)) + ((shiftx4x) & (!shiftx5x) & (g195) & (!g196) & (!g197) & (g198)) + ((shiftx4x) & (!shiftx5x) & (g195) & (!g196) & (g197) & (!g198)) + ((shiftx4x) & (!shiftx5x) & (g195) & (!g196) & (g197) & (g198)) + ((shiftx4x) & (!shiftx5x) & (g195) & (g196) & (!g197) & (!g198)) + ((shiftx4x) & (!shiftx5x) & (g195) & (g196) & (!g197) & (g198)) + ((shiftx4x) & (!shiftx5x) & (g195) & (g196) & (g197) & (!g198)) + ((shiftx4x) & (!shiftx5x) & (g195) & (g196) & (g197) & (g198)) + ((shiftx4x) & (shiftx5x) & (!g195) & (!g196) & (!g197) & (g198)) + ((shiftx4x) & (shiftx5x) & (!g195) & (!g196) & (g197) & (g198)) + ((shiftx4x) & (shiftx5x) & (!g195) & (g196) & (!g197) & (g198)) + ((shiftx4x) & (shiftx5x) & (!g195) & (g196) & (g197) & (g198)) + ((shiftx4x) & (shiftx5x) & (g195) & (!g196) & (!g197) & (g198)) + ((shiftx4x) & (shiftx5x) & (g195) & (!g196) & (g197) & (g198)) + ((shiftx4x) & (shiftx5x) & (g195) & (g196) & (!g197) & (g198)) + ((shiftx4x) & (shiftx5x) & (g195) & (g196) & (g197) & (g198)));
	assign g200 = (((!shiftx2x) & (!shiftx3x) & (!g108) & (!g109) & (!g111) & (g115)) + ((!shiftx2x) & (!shiftx3x) & (!g108) & (!g109) & (g111) & (g115)) + ((!shiftx2x) & (!shiftx3x) & (!g108) & (g109) & (!g111) & (g115)) + ((!shiftx2x) & (!shiftx3x) & (!g108) & (g109) & (g111) & (g115)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (!g109) & (!g111) & (g115)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (!g109) & (g111) & (g115)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (g109) & (!g111) & (g115)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (g109) & (g111) & (g115)) + ((!shiftx2x) & (shiftx3x) & (!g108) & (g109) & (!g111) & (!g115)) + ((!shiftx2x) & (shiftx3x) & (!g108) & (g109) & (!g111) & (g115)) + ((!shiftx2x) & (shiftx3x) & (!g108) & (g109) & (g111) & (!g115)) + ((!shiftx2x) & (shiftx3x) & (!g108) & (g109) & (g111) & (g115)) + ((!shiftx2x) & (shiftx3x) & (g108) & (g109) & (!g111) & (!g115)) + ((!shiftx2x) & (shiftx3x) & (g108) & (g109) & (!g111) & (g115)) + ((!shiftx2x) & (shiftx3x) & (g108) & (g109) & (g111) & (!g115)) + ((!shiftx2x) & (shiftx3x) & (g108) & (g109) & (g111) & (g115)) + ((shiftx2x) & (!shiftx3x) & (g108) & (!g109) & (!g111) & (!g115)) + ((shiftx2x) & (!shiftx3x) & (g108) & (!g109) & (!g111) & (g115)) + ((shiftx2x) & (!shiftx3x) & (g108) & (!g109) & (g111) & (!g115)) + ((shiftx2x) & (!shiftx3x) & (g108) & (!g109) & (g111) & (g115)) + ((shiftx2x) & (!shiftx3x) & (g108) & (g109) & (!g111) & (!g115)) + ((shiftx2x) & (!shiftx3x) & (g108) & (g109) & (!g111) & (g115)) + ((shiftx2x) & (!shiftx3x) & (g108) & (g109) & (g111) & (!g115)) + ((shiftx2x) & (!shiftx3x) & (g108) & (g109) & (g111) & (g115)) + ((shiftx2x) & (shiftx3x) & (!g108) & (!g109) & (g111) & (!g115)) + ((shiftx2x) & (shiftx3x) & (!g108) & (!g109) & (g111) & (g115)) + ((shiftx2x) & (shiftx3x) & (!g108) & (g109) & (g111) & (!g115)) + ((shiftx2x) & (shiftx3x) & (!g108) & (g109) & (g111) & (g115)) + ((shiftx2x) & (shiftx3x) & (g108) & (!g109) & (g111) & (!g115)) + ((shiftx2x) & (shiftx3x) & (g108) & (!g109) & (g111) & (g115)) + ((shiftx2x) & (shiftx3x) & (g108) & (g109) & (g111) & (!g115)) + ((shiftx2x) & (shiftx3x) & (g108) & (g109) & (g111) & (g115)));
	assign g201 = (((!shiftx2x) & (!shiftx3x) & (!g113) & (!g114) & (!g116) & (g125)) + ((!shiftx2x) & (!shiftx3x) & (!g113) & (!g114) & (g116) & (g125)) + ((!shiftx2x) & (!shiftx3x) & (!g113) & (g114) & (!g116) & (g125)) + ((!shiftx2x) & (!shiftx3x) & (!g113) & (g114) & (g116) & (g125)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (!g114) & (!g116) & (g125)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (!g114) & (g116) & (g125)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (g114) & (!g116) & (g125)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (g114) & (g116) & (g125)) + ((!shiftx2x) & (shiftx3x) & (!g113) & (g114) & (!g116) & (!g125)) + ((!shiftx2x) & (shiftx3x) & (!g113) & (g114) & (!g116) & (g125)) + ((!shiftx2x) & (shiftx3x) & (!g113) & (g114) & (g116) & (!g125)) + ((!shiftx2x) & (shiftx3x) & (!g113) & (g114) & (g116) & (g125)) + ((!shiftx2x) & (shiftx3x) & (g113) & (g114) & (!g116) & (!g125)) + ((!shiftx2x) & (shiftx3x) & (g113) & (g114) & (!g116) & (g125)) + ((!shiftx2x) & (shiftx3x) & (g113) & (g114) & (g116) & (!g125)) + ((!shiftx2x) & (shiftx3x) & (g113) & (g114) & (g116) & (g125)) + ((shiftx2x) & (!shiftx3x) & (g113) & (!g114) & (!g116) & (!g125)) + ((shiftx2x) & (!shiftx3x) & (g113) & (!g114) & (!g116) & (g125)) + ((shiftx2x) & (!shiftx3x) & (g113) & (!g114) & (g116) & (!g125)) + ((shiftx2x) & (!shiftx3x) & (g113) & (!g114) & (g116) & (g125)) + ((shiftx2x) & (!shiftx3x) & (g113) & (g114) & (!g116) & (!g125)) + ((shiftx2x) & (!shiftx3x) & (g113) & (g114) & (!g116) & (g125)) + ((shiftx2x) & (!shiftx3x) & (g113) & (g114) & (g116) & (!g125)) + ((shiftx2x) & (!shiftx3x) & (g113) & (g114) & (g116) & (g125)) + ((shiftx2x) & (shiftx3x) & (!g113) & (!g114) & (g116) & (!g125)) + ((shiftx2x) & (shiftx3x) & (!g113) & (!g114) & (g116) & (g125)) + ((shiftx2x) & (shiftx3x) & (!g113) & (g114) & (g116) & (!g125)) + ((shiftx2x) & (shiftx3x) & (!g113) & (g114) & (g116) & (g125)) + ((shiftx2x) & (shiftx3x) & (g113) & (!g114) & (g116) & (!g125)) + ((shiftx2x) & (shiftx3x) & (g113) & (!g114) & (g116) & (g125)) + ((shiftx2x) & (shiftx3x) & (g113) & (g114) & (g116) & (!g125)) + ((shiftx2x) & (shiftx3x) & (g113) & (g114) & (g116) & (g125)));
	assign g202 = (((!shiftx2x) & (!shiftx3x) & (g94) & (!g118) & (!g119) & (!g121)) + ((!shiftx2x) & (!shiftx3x) & (g94) & (!g118) & (!g119) & (g121)) + ((!shiftx2x) & (!shiftx3x) & (g94) & (!g118) & (g119) & (!g121)) + ((!shiftx2x) & (!shiftx3x) & (g94) & (!g118) & (g119) & (g121)) + ((!shiftx2x) & (!shiftx3x) & (g94) & (g118) & (!g119) & (!g121)) + ((!shiftx2x) & (!shiftx3x) & (g94) & (g118) & (!g119) & (g121)) + ((!shiftx2x) & (!shiftx3x) & (g94) & (g118) & (g119) & (!g121)) + ((!shiftx2x) & (!shiftx3x) & (g94) & (g118) & (g119) & (g121)) + ((!shiftx2x) & (shiftx3x) & (!g94) & (!g118) & (g119) & (!g121)) + ((!shiftx2x) & (shiftx3x) & (!g94) & (!g118) & (g119) & (g121)) + ((!shiftx2x) & (shiftx3x) & (!g94) & (g118) & (g119) & (!g121)) + ((!shiftx2x) & (shiftx3x) & (!g94) & (g118) & (g119) & (g121)) + ((!shiftx2x) & (shiftx3x) & (g94) & (!g118) & (g119) & (!g121)) + ((!shiftx2x) & (shiftx3x) & (g94) & (!g118) & (g119) & (g121)) + ((!shiftx2x) & (shiftx3x) & (g94) & (g118) & (g119) & (!g121)) + ((!shiftx2x) & (shiftx3x) & (g94) & (g118) & (g119) & (g121)) + ((shiftx2x) & (!shiftx3x) & (!g94) & (g118) & (!g119) & (!g121)) + ((shiftx2x) & (!shiftx3x) & (!g94) & (g118) & (!g119) & (g121)) + ((shiftx2x) & (!shiftx3x) & (!g94) & (g118) & (g119) & (!g121)) + ((shiftx2x) & (!shiftx3x) & (!g94) & (g118) & (g119) & (g121)) + ((shiftx2x) & (!shiftx3x) & (g94) & (g118) & (!g119) & (!g121)) + ((shiftx2x) & (!shiftx3x) & (g94) & (g118) & (!g119) & (g121)) + ((shiftx2x) & (!shiftx3x) & (g94) & (g118) & (g119) & (!g121)) + ((shiftx2x) & (!shiftx3x) & (g94) & (g118) & (g119) & (g121)) + ((shiftx2x) & (shiftx3x) & (!g94) & (!g118) & (!g119) & (g121)) + ((shiftx2x) & (shiftx3x) & (!g94) & (!g118) & (g119) & (g121)) + ((shiftx2x) & (shiftx3x) & (!g94) & (g118) & (!g119) & (g121)) + ((shiftx2x) & (shiftx3x) & (!g94) & (g118) & (g119) & (g121)) + ((shiftx2x) & (shiftx3x) & (g94) & (!g118) & (!g119) & (g121)) + ((shiftx2x) & (shiftx3x) & (g94) & (!g118) & (g119) & (g121)) + ((shiftx2x) & (shiftx3x) & (g94) & (g118) & (!g119) & (g121)) + ((shiftx2x) & (shiftx3x) & (g94) & (g118) & (g119) & (g121)));
	assign g203 = (((!shiftx2x) & (!shiftx3x) & (g120) & (!g123) & (!g124) & (!g126)) + ((!shiftx2x) & (!shiftx3x) & (g120) & (!g123) & (!g124) & (g126)) + ((!shiftx2x) & (!shiftx3x) & (g120) & (!g123) & (g124) & (!g126)) + ((!shiftx2x) & (!shiftx3x) & (g120) & (!g123) & (g124) & (g126)) + ((!shiftx2x) & (!shiftx3x) & (g120) & (g123) & (!g124) & (!g126)) + ((!shiftx2x) & (!shiftx3x) & (g120) & (g123) & (!g124) & (g126)) + ((!shiftx2x) & (!shiftx3x) & (g120) & (g123) & (g124) & (!g126)) + ((!shiftx2x) & (!shiftx3x) & (g120) & (g123) & (g124) & (g126)) + ((!shiftx2x) & (shiftx3x) & (!g120) & (!g123) & (g124) & (!g126)) + ((!shiftx2x) & (shiftx3x) & (!g120) & (!g123) & (g124) & (g126)) + ((!shiftx2x) & (shiftx3x) & (!g120) & (g123) & (g124) & (!g126)) + ((!shiftx2x) & (shiftx3x) & (!g120) & (g123) & (g124) & (g126)) + ((!shiftx2x) & (shiftx3x) & (g120) & (!g123) & (g124) & (!g126)) + ((!shiftx2x) & (shiftx3x) & (g120) & (!g123) & (g124) & (g126)) + ((!shiftx2x) & (shiftx3x) & (g120) & (g123) & (g124) & (!g126)) + ((!shiftx2x) & (shiftx3x) & (g120) & (g123) & (g124) & (g126)) + ((shiftx2x) & (!shiftx3x) & (!g120) & (g123) & (!g124) & (!g126)) + ((shiftx2x) & (!shiftx3x) & (!g120) & (g123) & (!g124) & (g126)) + ((shiftx2x) & (!shiftx3x) & (!g120) & (g123) & (g124) & (!g126)) + ((shiftx2x) & (!shiftx3x) & (!g120) & (g123) & (g124) & (g126)) + ((shiftx2x) & (!shiftx3x) & (g120) & (g123) & (!g124) & (!g126)) + ((shiftx2x) & (!shiftx3x) & (g120) & (g123) & (!g124) & (g126)) + ((shiftx2x) & (!shiftx3x) & (g120) & (g123) & (g124) & (!g126)) + ((shiftx2x) & (!shiftx3x) & (g120) & (g123) & (g124) & (g126)) + ((shiftx2x) & (shiftx3x) & (!g120) & (!g123) & (!g124) & (g126)) + ((shiftx2x) & (shiftx3x) & (!g120) & (!g123) & (g124) & (g126)) + ((shiftx2x) & (shiftx3x) & (!g120) & (g123) & (!g124) & (g126)) + ((shiftx2x) & (shiftx3x) & (!g120) & (g123) & (g124) & (g126)) + ((shiftx2x) & (shiftx3x) & (g120) & (!g123) & (!g124) & (g126)) + ((shiftx2x) & (shiftx3x) & (g120) & (!g123) & (g124) & (g126)) + ((shiftx2x) & (shiftx3x) & (g120) & (g123) & (!g124) & (g126)) + ((shiftx2x) & (shiftx3x) & (g120) & (g123) & (g124) & (g126)));
	assign g204 = (((!shiftx4x) & (!shiftx5x) & (!g200) & (!g201) & (g202) & (!g203)) + ((!shiftx4x) & (!shiftx5x) & (!g200) & (!g201) & (g202) & (g203)) + ((!shiftx4x) & (!shiftx5x) & (!g200) & (g201) & (g202) & (!g203)) + ((!shiftx4x) & (!shiftx5x) & (!g200) & (g201) & (g202) & (g203)) + ((!shiftx4x) & (!shiftx5x) & (g200) & (!g201) & (g202) & (!g203)) + ((!shiftx4x) & (!shiftx5x) & (g200) & (!g201) & (g202) & (g203)) + ((!shiftx4x) & (!shiftx5x) & (g200) & (g201) & (g202) & (!g203)) + ((!shiftx4x) & (!shiftx5x) & (g200) & (g201) & (g202) & (g203)) + ((!shiftx4x) & (shiftx5x) & (!g200) & (g201) & (!g202) & (!g203)) + ((!shiftx4x) & (shiftx5x) & (!g200) & (g201) & (!g202) & (g203)) + ((!shiftx4x) & (shiftx5x) & (!g200) & (g201) & (g202) & (!g203)) + ((!shiftx4x) & (shiftx5x) & (!g200) & (g201) & (g202) & (g203)) + ((!shiftx4x) & (shiftx5x) & (g200) & (g201) & (!g202) & (!g203)) + ((!shiftx4x) & (shiftx5x) & (g200) & (g201) & (!g202) & (g203)) + ((!shiftx4x) & (shiftx5x) & (g200) & (g201) & (g202) & (!g203)) + ((!shiftx4x) & (shiftx5x) & (g200) & (g201) & (g202) & (g203)) + ((shiftx4x) & (!shiftx5x) & (!g200) & (!g201) & (!g202) & (g203)) + ((shiftx4x) & (!shiftx5x) & (!g200) & (!g201) & (g202) & (g203)) + ((shiftx4x) & (!shiftx5x) & (!g200) & (g201) & (!g202) & (g203)) + ((shiftx4x) & (!shiftx5x) & (!g200) & (g201) & (g202) & (g203)) + ((shiftx4x) & (!shiftx5x) & (g200) & (!g201) & (!g202) & (g203)) + ((shiftx4x) & (!shiftx5x) & (g200) & (!g201) & (g202) & (g203)) + ((shiftx4x) & (!shiftx5x) & (g200) & (g201) & (!g202) & (g203)) + ((shiftx4x) & (!shiftx5x) & (g200) & (g201) & (g202) & (g203)) + ((shiftx4x) & (shiftx5x) & (g200) & (!g201) & (!g202) & (!g203)) + ((shiftx4x) & (shiftx5x) & (g200) & (!g201) & (!g202) & (g203)) + ((shiftx4x) & (shiftx5x) & (g200) & (!g201) & (g202) & (!g203)) + ((shiftx4x) & (shiftx5x) & (g200) & (!g201) & (g202) & (g203)) + ((shiftx4x) & (shiftx5x) & (g200) & (g201) & (!g202) & (!g203)) + ((shiftx4x) & (shiftx5x) & (g200) & (g201) & (!g202) & (g203)) + ((shiftx4x) & (shiftx5x) & (g200) & (g201) & (g202) & (!g203)) + ((shiftx4x) & (shiftx5x) & (g200) & (g201) & (g202) & (g203)));
	assign resultx6x = (((!shiftx6x) & (sk[76]) & (!g199) & (g204)) + ((!shiftx6x) & (sk[76]) & (g199) & (g204)) + ((shiftx6x) & (!sk[76]) & (!g199) & (!g204)) + ((shiftx6x) & (!sk[76]) & (!g199) & (g204)) + ((shiftx6x) & (!sk[76]) & (g199) & (!g204)) + ((shiftx6x) & (!sk[76]) & (g199) & (g204)) + ((shiftx6x) & (sk[76]) & (g199) & (!g204)) + ((shiftx6x) & (sk[76]) & (g199) & (g204)));
	assign g206 = (((!shiftx2x) & (!shiftx3x) & (g132) & (!g135) & (!g136) & (!g138)) + ((!shiftx2x) & (!shiftx3x) & (g132) & (!g135) & (!g136) & (g138)) + ((!shiftx2x) & (!shiftx3x) & (g132) & (!g135) & (g136) & (!g138)) + ((!shiftx2x) & (!shiftx3x) & (g132) & (!g135) & (g136) & (g138)) + ((!shiftx2x) & (!shiftx3x) & (g132) & (g135) & (!g136) & (!g138)) + ((!shiftx2x) & (!shiftx3x) & (g132) & (g135) & (!g136) & (g138)) + ((!shiftx2x) & (!shiftx3x) & (g132) & (g135) & (g136) & (!g138)) + ((!shiftx2x) & (!shiftx3x) & (g132) & (g135) & (g136) & (g138)) + ((!shiftx2x) & (shiftx3x) & (!g132) & (!g135) & (g136) & (!g138)) + ((!shiftx2x) & (shiftx3x) & (!g132) & (!g135) & (g136) & (g138)) + ((!shiftx2x) & (shiftx3x) & (!g132) & (g135) & (g136) & (!g138)) + ((!shiftx2x) & (shiftx3x) & (!g132) & (g135) & (g136) & (g138)) + ((!shiftx2x) & (shiftx3x) & (g132) & (!g135) & (g136) & (!g138)) + ((!shiftx2x) & (shiftx3x) & (g132) & (!g135) & (g136) & (g138)) + ((!shiftx2x) & (shiftx3x) & (g132) & (g135) & (g136) & (!g138)) + ((!shiftx2x) & (shiftx3x) & (g132) & (g135) & (g136) & (g138)) + ((shiftx2x) & (!shiftx3x) & (!g132) & (g135) & (!g136) & (!g138)) + ((shiftx2x) & (!shiftx3x) & (!g132) & (g135) & (!g136) & (g138)) + ((shiftx2x) & (!shiftx3x) & (!g132) & (g135) & (g136) & (!g138)) + ((shiftx2x) & (!shiftx3x) & (!g132) & (g135) & (g136) & (g138)) + ((shiftx2x) & (!shiftx3x) & (g132) & (g135) & (!g136) & (!g138)) + ((shiftx2x) & (!shiftx3x) & (g132) & (g135) & (!g136) & (g138)) + ((shiftx2x) & (!shiftx3x) & (g132) & (g135) & (g136) & (!g138)) + ((shiftx2x) & (!shiftx3x) & (g132) & (g135) & (g136) & (g138)) + ((shiftx2x) & (shiftx3x) & (!g132) & (!g135) & (!g136) & (g138)) + ((shiftx2x) & (shiftx3x) & (!g132) & (!g135) & (g136) & (g138)) + ((shiftx2x) & (shiftx3x) & (!g132) & (g135) & (!g136) & (g138)) + ((shiftx2x) & (shiftx3x) & (!g132) & (g135) & (g136) & (g138)) + ((shiftx2x) & (shiftx3x) & (g132) & (!g135) & (!g136) & (g138)) + ((shiftx2x) & (shiftx3x) & (g132) & (!g135) & (g136) & (g138)) + ((shiftx2x) & (shiftx3x) & (g132) & (g135) & (!g136) & (g138)) + ((shiftx2x) & (shiftx3x) & (g132) & (g135) & (g136) & (g138)));
	assign g207 = (((!shiftx2x) & (!shiftx3x) & (!g130) & (!g131) & (!g133) & (g168)) + ((!shiftx2x) & (!shiftx3x) & (!g130) & (!g131) & (g133) & (g168)) + ((!shiftx2x) & (!shiftx3x) & (!g130) & (g131) & (!g133) & (g168)) + ((!shiftx2x) & (!shiftx3x) & (!g130) & (g131) & (g133) & (g168)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (!g131) & (!g133) & (g168)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (!g131) & (g133) & (g168)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (g131) & (!g133) & (g168)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (g131) & (g133) & (g168)) + ((!shiftx2x) & (shiftx3x) & (!g130) & (g131) & (!g133) & (!g168)) + ((!shiftx2x) & (shiftx3x) & (!g130) & (g131) & (!g133) & (g168)) + ((!shiftx2x) & (shiftx3x) & (!g130) & (g131) & (g133) & (!g168)) + ((!shiftx2x) & (shiftx3x) & (!g130) & (g131) & (g133) & (g168)) + ((!shiftx2x) & (shiftx3x) & (g130) & (g131) & (!g133) & (!g168)) + ((!shiftx2x) & (shiftx3x) & (g130) & (g131) & (!g133) & (g168)) + ((!shiftx2x) & (shiftx3x) & (g130) & (g131) & (g133) & (!g168)) + ((!shiftx2x) & (shiftx3x) & (g130) & (g131) & (g133) & (g168)) + ((shiftx2x) & (!shiftx3x) & (g130) & (!g131) & (!g133) & (!g168)) + ((shiftx2x) & (!shiftx3x) & (g130) & (!g131) & (!g133) & (g168)) + ((shiftx2x) & (!shiftx3x) & (g130) & (!g131) & (g133) & (!g168)) + ((shiftx2x) & (!shiftx3x) & (g130) & (!g131) & (g133) & (g168)) + ((shiftx2x) & (!shiftx3x) & (g130) & (g131) & (!g133) & (!g168)) + ((shiftx2x) & (!shiftx3x) & (g130) & (g131) & (!g133) & (g168)) + ((shiftx2x) & (!shiftx3x) & (g130) & (g131) & (g133) & (!g168)) + ((shiftx2x) & (!shiftx3x) & (g130) & (g131) & (g133) & (g168)) + ((shiftx2x) & (shiftx3x) & (!g130) & (!g131) & (g133) & (!g168)) + ((shiftx2x) & (shiftx3x) & (!g130) & (!g131) & (g133) & (g168)) + ((shiftx2x) & (shiftx3x) & (!g130) & (g131) & (g133) & (!g168)) + ((shiftx2x) & (shiftx3x) & (!g130) & (g131) & (g133) & (g168)) + ((shiftx2x) & (shiftx3x) & (g130) & (!g131) & (g133) & (!g168)) + ((shiftx2x) & (shiftx3x) & (g130) & (!g131) & (g133) & (g168)) + ((shiftx2x) & (shiftx3x) & (g130) & (g131) & (g133) & (!g168)) + ((shiftx2x) & (shiftx3x) & (g130) & (g131) & (g133) & (g168)));
	assign g208 = (((!shiftx2x) & (!shiftx3x) & (g137) & (!g145) & (!g146) & (!g148)) + ((!shiftx2x) & (!shiftx3x) & (g137) & (!g145) & (!g146) & (g148)) + ((!shiftx2x) & (!shiftx3x) & (g137) & (!g145) & (g146) & (!g148)) + ((!shiftx2x) & (!shiftx3x) & (g137) & (!g145) & (g146) & (g148)) + ((!shiftx2x) & (!shiftx3x) & (g137) & (g145) & (!g146) & (!g148)) + ((!shiftx2x) & (!shiftx3x) & (g137) & (g145) & (!g146) & (g148)) + ((!shiftx2x) & (!shiftx3x) & (g137) & (g145) & (g146) & (!g148)) + ((!shiftx2x) & (!shiftx3x) & (g137) & (g145) & (g146) & (g148)) + ((!shiftx2x) & (shiftx3x) & (!g137) & (!g145) & (g146) & (!g148)) + ((!shiftx2x) & (shiftx3x) & (!g137) & (!g145) & (g146) & (g148)) + ((!shiftx2x) & (shiftx3x) & (!g137) & (g145) & (g146) & (!g148)) + ((!shiftx2x) & (shiftx3x) & (!g137) & (g145) & (g146) & (g148)) + ((!shiftx2x) & (shiftx3x) & (g137) & (!g145) & (g146) & (!g148)) + ((!shiftx2x) & (shiftx3x) & (g137) & (!g145) & (g146) & (g148)) + ((!shiftx2x) & (shiftx3x) & (g137) & (g145) & (g146) & (!g148)) + ((!shiftx2x) & (shiftx3x) & (g137) & (g145) & (g146) & (g148)) + ((shiftx2x) & (!shiftx3x) & (!g137) & (g145) & (!g146) & (!g148)) + ((shiftx2x) & (!shiftx3x) & (!g137) & (g145) & (!g146) & (g148)) + ((shiftx2x) & (!shiftx3x) & (!g137) & (g145) & (g146) & (!g148)) + ((shiftx2x) & (!shiftx3x) & (!g137) & (g145) & (g146) & (g148)) + ((shiftx2x) & (!shiftx3x) & (g137) & (g145) & (!g146) & (!g148)) + ((shiftx2x) & (!shiftx3x) & (g137) & (g145) & (!g146) & (g148)) + ((shiftx2x) & (!shiftx3x) & (g137) & (g145) & (g146) & (!g148)) + ((shiftx2x) & (!shiftx3x) & (g137) & (g145) & (g146) & (g148)) + ((shiftx2x) & (shiftx3x) & (!g137) & (!g145) & (!g146) & (g148)) + ((shiftx2x) & (shiftx3x) & (!g137) & (!g145) & (g146) & (g148)) + ((shiftx2x) & (shiftx3x) & (!g137) & (g145) & (!g146) & (g148)) + ((shiftx2x) & (shiftx3x) & (!g137) & (g145) & (g146) & (g148)) + ((shiftx2x) & (shiftx3x) & (g137) & (!g145) & (!g146) & (g148)) + ((shiftx2x) & (shiftx3x) & (g137) & (!g145) & (g146) & (g148)) + ((shiftx2x) & (shiftx3x) & (g137) & (g145) & (!g146) & (g148)) + ((shiftx2x) & (shiftx3x) & (g137) & (g145) & (g146) & (g148)));
	assign g209 = (((!shiftx2x) & (!shiftx3x) & (!g140) & (!g141) & (!g143) & (g147)) + ((!shiftx2x) & (!shiftx3x) & (!g140) & (!g141) & (g143) & (g147)) + ((!shiftx2x) & (!shiftx3x) & (!g140) & (g141) & (!g143) & (g147)) + ((!shiftx2x) & (!shiftx3x) & (!g140) & (g141) & (g143) & (g147)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (!g141) & (!g143) & (g147)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (!g141) & (g143) & (g147)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (g141) & (!g143) & (g147)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (g141) & (g143) & (g147)) + ((!shiftx2x) & (shiftx3x) & (!g140) & (g141) & (!g143) & (!g147)) + ((!shiftx2x) & (shiftx3x) & (!g140) & (g141) & (!g143) & (g147)) + ((!shiftx2x) & (shiftx3x) & (!g140) & (g141) & (g143) & (!g147)) + ((!shiftx2x) & (shiftx3x) & (!g140) & (g141) & (g143) & (g147)) + ((!shiftx2x) & (shiftx3x) & (g140) & (g141) & (!g143) & (!g147)) + ((!shiftx2x) & (shiftx3x) & (g140) & (g141) & (!g143) & (g147)) + ((!shiftx2x) & (shiftx3x) & (g140) & (g141) & (g143) & (!g147)) + ((!shiftx2x) & (shiftx3x) & (g140) & (g141) & (g143) & (g147)) + ((shiftx2x) & (!shiftx3x) & (g140) & (!g141) & (!g143) & (!g147)) + ((shiftx2x) & (!shiftx3x) & (g140) & (!g141) & (!g143) & (g147)) + ((shiftx2x) & (!shiftx3x) & (g140) & (!g141) & (g143) & (!g147)) + ((shiftx2x) & (!shiftx3x) & (g140) & (!g141) & (g143) & (g147)) + ((shiftx2x) & (!shiftx3x) & (g140) & (g141) & (!g143) & (!g147)) + ((shiftx2x) & (!shiftx3x) & (g140) & (g141) & (!g143) & (g147)) + ((shiftx2x) & (!shiftx3x) & (g140) & (g141) & (g143) & (!g147)) + ((shiftx2x) & (!shiftx3x) & (g140) & (g141) & (g143) & (g147)) + ((shiftx2x) & (shiftx3x) & (!g140) & (!g141) & (g143) & (!g147)) + ((shiftx2x) & (shiftx3x) & (!g140) & (!g141) & (g143) & (g147)) + ((shiftx2x) & (shiftx3x) & (!g140) & (g141) & (g143) & (!g147)) + ((shiftx2x) & (shiftx3x) & (!g140) & (g141) & (g143) & (g147)) + ((shiftx2x) & (shiftx3x) & (g140) & (!g141) & (g143) & (!g147)) + ((shiftx2x) & (shiftx3x) & (g140) & (!g141) & (g143) & (g147)) + ((shiftx2x) & (shiftx3x) & (g140) & (g141) & (g143) & (!g147)) + ((shiftx2x) & (shiftx3x) & (g140) & (g141) & (g143) & (g147)));
	assign g210 = (((!shiftx4x) & (!shiftx5x) & (!g206) & (g207) & (!g208) & (!g209)) + ((!shiftx4x) & (!shiftx5x) & (!g206) & (g207) & (!g208) & (g209)) + ((!shiftx4x) & (!shiftx5x) & (!g206) & (g207) & (g208) & (!g209)) + ((!shiftx4x) & (!shiftx5x) & (!g206) & (g207) & (g208) & (g209)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (g207) & (!g208) & (!g209)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (g207) & (!g208) & (g209)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (g207) & (g208) & (!g209)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (g207) & (g208) & (g209)) + ((!shiftx4x) & (shiftx5x) & (!g206) & (!g207) & (g208) & (!g209)) + ((!shiftx4x) & (shiftx5x) & (!g206) & (!g207) & (g208) & (g209)) + ((!shiftx4x) & (shiftx5x) & (!g206) & (g207) & (g208) & (!g209)) + ((!shiftx4x) & (shiftx5x) & (!g206) & (g207) & (g208) & (g209)) + ((!shiftx4x) & (shiftx5x) & (g206) & (!g207) & (g208) & (!g209)) + ((!shiftx4x) & (shiftx5x) & (g206) & (!g207) & (g208) & (g209)) + ((!shiftx4x) & (shiftx5x) & (g206) & (g207) & (g208) & (!g209)) + ((!shiftx4x) & (shiftx5x) & (g206) & (g207) & (g208) & (g209)) + ((shiftx4x) & (!shiftx5x) & (g206) & (!g207) & (!g208) & (!g209)) + ((shiftx4x) & (!shiftx5x) & (g206) & (!g207) & (!g208) & (g209)) + ((shiftx4x) & (!shiftx5x) & (g206) & (!g207) & (g208) & (!g209)) + ((shiftx4x) & (!shiftx5x) & (g206) & (!g207) & (g208) & (g209)) + ((shiftx4x) & (!shiftx5x) & (g206) & (g207) & (!g208) & (!g209)) + ((shiftx4x) & (!shiftx5x) & (g206) & (g207) & (!g208) & (g209)) + ((shiftx4x) & (!shiftx5x) & (g206) & (g207) & (g208) & (!g209)) + ((shiftx4x) & (!shiftx5x) & (g206) & (g207) & (g208) & (g209)) + ((shiftx4x) & (shiftx5x) & (!g206) & (!g207) & (!g208) & (g209)) + ((shiftx4x) & (shiftx5x) & (!g206) & (!g207) & (g208) & (g209)) + ((shiftx4x) & (shiftx5x) & (!g206) & (g207) & (!g208) & (g209)) + ((shiftx4x) & (shiftx5x) & (!g206) & (g207) & (g208) & (g209)) + ((shiftx4x) & (shiftx5x) & (g206) & (!g207) & (!g208) & (g209)) + ((shiftx4x) & (shiftx5x) & (g206) & (!g207) & (g208) & (g209)) + ((shiftx4x) & (shiftx5x) & (g206) & (g207) & (!g208) & (g209)) + ((shiftx4x) & (shiftx5x) & (g206) & (g207) & (g208) & (g209)));
	assign g211 = (((!shiftx2x) & (!shiftx3x) & (g158) & (!g166) & (!g167) & (!g169)) + ((!shiftx2x) & (!shiftx3x) & (g158) & (!g166) & (!g167) & (g169)) + ((!shiftx2x) & (!shiftx3x) & (g158) & (!g166) & (g167) & (!g169)) + ((!shiftx2x) & (!shiftx3x) & (g158) & (!g166) & (g167) & (g169)) + ((!shiftx2x) & (!shiftx3x) & (g158) & (g166) & (!g167) & (!g169)) + ((!shiftx2x) & (!shiftx3x) & (g158) & (g166) & (!g167) & (g169)) + ((!shiftx2x) & (!shiftx3x) & (g158) & (g166) & (g167) & (!g169)) + ((!shiftx2x) & (!shiftx3x) & (g158) & (g166) & (g167) & (g169)) + ((!shiftx2x) & (shiftx3x) & (!g158) & (!g166) & (g167) & (!g169)) + ((!shiftx2x) & (shiftx3x) & (!g158) & (!g166) & (g167) & (g169)) + ((!shiftx2x) & (shiftx3x) & (!g158) & (g166) & (g167) & (!g169)) + ((!shiftx2x) & (shiftx3x) & (!g158) & (g166) & (g167) & (g169)) + ((!shiftx2x) & (shiftx3x) & (g158) & (!g166) & (g167) & (!g169)) + ((!shiftx2x) & (shiftx3x) & (g158) & (!g166) & (g167) & (g169)) + ((!shiftx2x) & (shiftx3x) & (g158) & (g166) & (g167) & (!g169)) + ((!shiftx2x) & (shiftx3x) & (g158) & (g166) & (g167) & (g169)) + ((shiftx2x) & (!shiftx3x) & (!g158) & (g166) & (!g167) & (!g169)) + ((shiftx2x) & (!shiftx3x) & (!g158) & (g166) & (!g167) & (g169)) + ((shiftx2x) & (!shiftx3x) & (!g158) & (g166) & (g167) & (!g169)) + ((shiftx2x) & (!shiftx3x) & (!g158) & (g166) & (g167) & (g169)) + ((shiftx2x) & (!shiftx3x) & (g158) & (g166) & (!g167) & (!g169)) + ((shiftx2x) & (!shiftx3x) & (g158) & (g166) & (!g167) & (g169)) + ((shiftx2x) & (!shiftx3x) & (g158) & (g166) & (g167) & (!g169)) + ((shiftx2x) & (!shiftx3x) & (g158) & (g166) & (g167) & (g169)) + ((shiftx2x) & (shiftx3x) & (!g158) & (!g166) & (!g167) & (g169)) + ((shiftx2x) & (shiftx3x) & (!g158) & (!g166) & (g167) & (g169)) + ((shiftx2x) & (shiftx3x) & (!g158) & (g166) & (!g167) & (g169)) + ((shiftx2x) & (shiftx3x) & (!g158) & (g166) & (g167) & (g169)) + ((shiftx2x) & (shiftx3x) & (g158) & (!g166) & (!g167) & (g169)) + ((shiftx2x) & (shiftx3x) & (g158) & (!g166) & (g167) & (g169)) + ((shiftx2x) & (shiftx3x) & (g158) & (g166) & (!g167) & (g169)) + ((shiftx2x) & (shiftx3x) & (g158) & (g166) & (g167) & (g169)));
	assign g212 = (((!shiftx2x) & (!shiftx3x) & (g153) & (!g156) & (!g157) & (!g159)) + ((!shiftx2x) & (!shiftx3x) & (g153) & (!g156) & (!g157) & (g159)) + ((!shiftx2x) & (!shiftx3x) & (g153) & (!g156) & (g157) & (!g159)) + ((!shiftx2x) & (!shiftx3x) & (g153) & (!g156) & (g157) & (g159)) + ((!shiftx2x) & (!shiftx3x) & (g153) & (g156) & (!g157) & (!g159)) + ((!shiftx2x) & (!shiftx3x) & (g153) & (g156) & (!g157) & (g159)) + ((!shiftx2x) & (!shiftx3x) & (g153) & (g156) & (g157) & (!g159)) + ((!shiftx2x) & (!shiftx3x) & (g153) & (g156) & (g157) & (g159)) + ((!shiftx2x) & (shiftx3x) & (!g153) & (!g156) & (g157) & (!g159)) + ((!shiftx2x) & (shiftx3x) & (!g153) & (!g156) & (g157) & (g159)) + ((!shiftx2x) & (shiftx3x) & (!g153) & (g156) & (g157) & (!g159)) + ((!shiftx2x) & (shiftx3x) & (!g153) & (g156) & (g157) & (g159)) + ((!shiftx2x) & (shiftx3x) & (g153) & (!g156) & (g157) & (!g159)) + ((!shiftx2x) & (shiftx3x) & (g153) & (!g156) & (g157) & (g159)) + ((!shiftx2x) & (shiftx3x) & (g153) & (g156) & (g157) & (!g159)) + ((!shiftx2x) & (shiftx3x) & (g153) & (g156) & (g157) & (g159)) + ((shiftx2x) & (!shiftx3x) & (!g153) & (g156) & (!g157) & (!g159)) + ((shiftx2x) & (!shiftx3x) & (!g153) & (g156) & (!g157) & (g159)) + ((shiftx2x) & (!shiftx3x) & (!g153) & (g156) & (g157) & (!g159)) + ((shiftx2x) & (!shiftx3x) & (!g153) & (g156) & (g157) & (g159)) + ((shiftx2x) & (!shiftx3x) & (g153) & (g156) & (!g157) & (!g159)) + ((shiftx2x) & (!shiftx3x) & (g153) & (g156) & (!g157) & (g159)) + ((shiftx2x) & (!shiftx3x) & (g153) & (g156) & (g157) & (!g159)) + ((shiftx2x) & (!shiftx3x) & (g153) & (g156) & (g157) & (g159)) + ((shiftx2x) & (shiftx3x) & (!g153) & (!g156) & (!g157) & (g159)) + ((shiftx2x) & (shiftx3x) & (!g153) & (!g156) & (g157) & (g159)) + ((shiftx2x) & (shiftx3x) & (!g153) & (g156) & (!g157) & (g159)) + ((shiftx2x) & (shiftx3x) & (!g153) & (g156) & (g157) & (g159)) + ((shiftx2x) & (shiftx3x) & (g153) & (!g156) & (!g157) & (g159)) + ((shiftx2x) & (shiftx3x) & (g153) & (!g156) & (g157) & (g159)) + ((shiftx2x) & (shiftx3x) & (g153) & (g156) & (!g157) & (g159)) + ((shiftx2x) & (shiftx3x) & (g153) & (g156) & (g157) & (g159)));
	assign g213 = (((!shiftx2x) & (!shiftx3x) & (g142) & (!g161) & (!g162) & (!g164)) + ((!shiftx2x) & (!shiftx3x) & (g142) & (!g161) & (!g162) & (g164)) + ((!shiftx2x) & (!shiftx3x) & (g142) & (!g161) & (g162) & (!g164)) + ((!shiftx2x) & (!shiftx3x) & (g142) & (!g161) & (g162) & (g164)) + ((!shiftx2x) & (!shiftx3x) & (g142) & (g161) & (!g162) & (!g164)) + ((!shiftx2x) & (!shiftx3x) & (g142) & (g161) & (!g162) & (g164)) + ((!shiftx2x) & (!shiftx3x) & (g142) & (g161) & (g162) & (!g164)) + ((!shiftx2x) & (!shiftx3x) & (g142) & (g161) & (g162) & (g164)) + ((!shiftx2x) & (shiftx3x) & (!g142) & (!g161) & (g162) & (!g164)) + ((!shiftx2x) & (shiftx3x) & (!g142) & (!g161) & (g162) & (g164)) + ((!shiftx2x) & (shiftx3x) & (!g142) & (g161) & (g162) & (!g164)) + ((!shiftx2x) & (shiftx3x) & (!g142) & (g161) & (g162) & (g164)) + ((!shiftx2x) & (shiftx3x) & (g142) & (!g161) & (g162) & (!g164)) + ((!shiftx2x) & (shiftx3x) & (g142) & (!g161) & (g162) & (g164)) + ((!shiftx2x) & (shiftx3x) & (g142) & (g161) & (g162) & (!g164)) + ((!shiftx2x) & (shiftx3x) & (g142) & (g161) & (g162) & (g164)) + ((shiftx2x) & (!shiftx3x) & (!g142) & (g161) & (!g162) & (!g164)) + ((shiftx2x) & (!shiftx3x) & (!g142) & (g161) & (!g162) & (g164)) + ((shiftx2x) & (!shiftx3x) & (!g142) & (g161) & (g162) & (!g164)) + ((shiftx2x) & (!shiftx3x) & (!g142) & (g161) & (g162) & (g164)) + ((shiftx2x) & (!shiftx3x) & (g142) & (g161) & (!g162) & (!g164)) + ((shiftx2x) & (!shiftx3x) & (g142) & (g161) & (!g162) & (g164)) + ((shiftx2x) & (!shiftx3x) & (g142) & (g161) & (g162) & (!g164)) + ((shiftx2x) & (!shiftx3x) & (g142) & (g161) & (g162) & (g164)) + ((shiftx2x) & (shiftx3x) & (!g142) & (!g161) & (!g162) & (g164)) + ((shiftx2x) & (shiftx3x) & (!g142) & (!g161) & (g162) & (g164)) + ((shiftx2x) & (shiftx3x) & (!g142) & (g161) & (!g162) & (g164)) + ((shiftx2x) & (shiftx3x) & (!g142) & (g161) & (g162) & (g164)) + ((shiftx2x) & (shiftx3x) & (g142) & (!g161) & (!g162) & (g164)) + ((shiftx2x) & (shiftx3x) & (g142) & (!g161) & (g162) & (g164)) + ((shiftx2x) & (shiftx3x) & (g142) & (g161) & (!g162) & (g164)) + ((shiftx2x) & (shiftx3x) & (g142) & (g161) & (g162) & (g164)));
	assign g214 = (((!shiftx2x) & (!shiftx3x) & (!g151) & (!g152) & (!g154) & (g163)) + ((!shiftx2x) & (!shiftx3x) & (!g151) & (!g152) & (g154) & (g163)) + ((!shiftx2x) & (!shiftx3x) & (!g151) & (g152) & (!g154) & (g163)) + ((!shiftx2x) & (!shiftx3x) & (!g151) & (g152) & (g154) & (g163)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (!g152) & (!g154) & (g163)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (!g152) & (g154) & (g163)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (g152) & (!g154) & (g163)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (g152) & (g154) & (g163)) + ((!shiftx2x) & (shiftx3x) & (!g151) & (g152) & (!g154) & (!g163)) + ((!shiftx2x) & (shiftx3x) & (!g151) & (g152) & (!g154) & (g163)) + ((!shiftx2x) & (shiftx3x) & (!g151) & (g152) & (g154) & (!g163)) + ((!shiftx2x) & (shiftx3x) & (!g151) & (g152) & (g154) & (g163)) + ((!shiftx2x) & (shiftx3x) & (g151) & (g152) & (!g154) & (!g163)) + ((!shiftx2x) & (shiftx3x) & (g151) & (g152) & (!g154) & (g163)) + ((!shiftx2x) & (shiftx3x) & (g151) & (g152) & (g154) & (!g163)) + ((!shiftx2x) & (shiftx3x) & (g151) & (g152) & (g154) & (g163)) + ((shiftx2x) & (!shiftx3x) & (g151) & (!g152) & (!g154) & (!g163)) + ((shiftx2x) & (!shiftx3x) & (g151) & (!g152) & (!g154) & (g163)) + ((shiftx2x) & (!shiftx3x) & (g151) & (!g152) & (g154) & (!g163)) + ((shiftx2x) & (!shiftx3x) & (g151) & (!g152) & (g154) & (g163)) + ((shiftx2x) & (!shiftx3x) & (g151) & (g152) & (!g154) & (!g163)) + ((shiftx2x) & (!shiftx3x) & (g151) & (g152) & (!g154) & (g163)) + ((shiftx2x) & (!shiftx3x) & (g151) & (g152) & (g154) & (!g163)) + ((shiftx2x) & (!shiftx3x) & (g151) & (g152) & (g154) & (g163)) + ((shiftx2x) & (shiftx3x) & (!g151) & (!g152) & (g154) & (!g163)) + ((shiftx2x) & (shiftx3x) & (!g151) & (!g152) & (g154) & (g163)) + ((shiftx2x) & (shiftx3x) & (!g151) & (g152) & (g154) & (!g163)) + ((shiftx2x) & (shiftx3x) & (!g151) & (g152) & (g154) & (g163)) + ((shiftx2x) & (shiftx3x) & (g151) & (!g152) & (g154) & (!g163)) + ((shiftx2x) & (shiftx3x) & (g151) & (!g152) & (g154) & (g163)) + ((shiftx2x) & (shiftx3x) & (g151) & (g152) & (g154) & (!g163)) + ((shiftx2x) & (shiftx3x) & (g151) & (g152) & (g154) & (g163)));
	assign g215 = (((!shiftx4x) & (!shiftx5x) & (!g211) & (!g212) & (g213) & (!g214)) + ((!shiftx4x) & (!shiftx5x) & (!g211) & (!g212) & (g213) & (g214)) + ((!shiftx4x) & (!shiftx5x) & (!g211) & (g212) & (g213) & (!g214)) + ((!shiftx4x) & (!shiftx5x) & (!g211) & (g212) & (g213) & (g214)) + ((!shiftx4x) & (!shiftx5x) & (g211) & (!g212) & (g213) & (!g214)) + ((!shiftx4x) & (!shiftx5x) & (g211) & (!g212) & (g213) & (g214)) + ((!shiftx4x) & (!shiftx5x) & (g211) & (g212) & (g213) & (!g214)) + ((!shiftx4x) & (!shiftx5x) & (g211) & (g212) & (g213) & (g214)) + ((!shiftx4x) & (shiftx5x) & (!g211) & (g212) & (!g213) & (!g214)) + ((!shiftx4x) & (shiftx5x) & (!g211) & (g212) & (!g213) & (g214)) + ((!shiftx4x) & (shiftx5x) & (!g211) & (g212) & (g213) & (!g214)) + ((!shiftx4x) & (shiftx5x) & (!g211) & (g212) & (g213) & (g214)) + ((!shiftx4x) & (shiftx5x) & (g211) & (g212) & (!g213) & (!g214)) + ((!shiftx4x) & (shiftx5x) & (g211) & (g212) & (!g213) & (g214)) + ((!shiftx4x) & (shiftx5x) & (g211) & (g212) & (g213) & (!g214)) + ((!shiftx4x) & (shiftx5x) & (g211) & (g212) & (g213) & (g214)) + ((shiftx4x) & (!shiftx5x) & (!g211) & (!g212) & (!g213) & (g214)) + ((shiftx4x) & (!shiftx5x) & (!g211) & (!g212) & (g213) & (g214)) + ((shiftx4x) & (!shiftx5x) & (!g211) & (g212) & (!g213) & (g214)) + ((shiftx4x) & (!shiftx5x) & (!g211) & (g212) & (g213) & (g214)) + ((shiftx4x) & (!shiftx5x) & (g211) & (!g212) & (!g213) & (g214)) + ((shiftx4x) & (!shiftx5x) & (g211) & (!g212) & (g213) & (g214)) + ((shiftx4x) & (!shiftx5x) & (g211) & (g212) & (!g213) & (g214)) + ((shiftx4x) & (!shiftx5x) & (g211) & (g212) & (g213) & (g214)) + ((shiftx4x) & (shiftx5x) & (g211) & (!g212) & (!g213) & (!g214)) + ((shiftx4x) & (shiftx5x) & (g211) & (!g212) & (!g213) & (g214)) + ((shiftx4x) & (shiftx5x) & (g211) & (!g212) & (g213) & (!g214)) + ((shiftx4x) & (shiftx5x) & (g211) & (!g212) & (g213) & (g214)) + ((shiftx4x) & (shiftx5x) & (g211) & (g212) & (!g213) & (!g214)) + ((shiftx4x) & (shiftx5x) & (g211) & (g212) & (!g213) & (g214)) + ((shiftx4x) & (shiftx5x) & (g211) & (g212) & (g213) & (!g214)) + ((shiftx4x) & (shiftx5x) & (g211) & (g212) & (g213) & (g214)));
	assign resultx7x = (((!shiftx6x) & (sk[87]) & (!g210) & (g215)) + ((!shiftx6x) & (sk[87]) & (g210) & (g215)) + ((shiftx6x) & (!sk[87]) & (!g210) & (!g215)) + ((shiftx6x) & (!sk[87]) & (!g210) & (g215)) + ((shiftx6x) & (!sk[87]) & (g210) & (!g215)) + ((shiftx6x) & (!sk[87]) & (g210) & (g215)) + ((shiftx6x) & (sk[87]) & (g210) & (!g215)) + ((shiftx6x) & (sk[87]) & (g210) & (g215)));
	assign g217 = (((!shiftx2x) & (!shiftx3x) & (!g13) & (g14) & (!g16) & (!g17)) + ((!shiftx2x) & (!shiftx3x) & (!g13) & (g14) & (!g16) & (g17)) + ((!shiftx2x) & (!shiftx3x) & (!g13) & (g14) & (g16) & (!g17)) + ((!shiftx2x) & (!shiftx3x) & (!g13) & (g14) & (g16) & (g17)) + ((!shiftx2x) & (!shiftx3x) & (g13) & (g14) & (!g16) & (!g17)) + ((!shiftx2x) & (!shiftx3x) & (g13) & (g14) & (!g16) & (g17)) + ((!shiftx2x) & (!shiftx3x) & (g13) & (g14) & (g16) & (!g17)) + ((!shiftx2x) & (!shiftx3x) & (g13) & (g14) & (g16) & (g17)) + ((!shiftx2x) & (shiftx3x) & (!g13) & (!g14) & (g16) & (!g17)) + ((!shiftx2x) & (shiftx3x) & (!g13) & (!g14) & (g16) & (g17)) + ((!shiftx2x) & (shiftx3x) & (!g13) & (g14) & (g16) & (!g17)) + ((!shiftx2x) & (shiftx3x) & (!g13) & (g14) & (g16) & (g17)) + ((!shiftx2x) & (shiftx3x) & (g13) & (!g14) & (g16) & (!g17)) + ((!shiftx2x) & (shiftx3x) & (g13) & (!g14) & (g16) & (g17)) + ((!shiftx2x) & (shiftx3x) & (g13) & (g14) & (g16) & (!g17)) + ((!shiftx2x) & (shiftx3x) & (g13) & (g14) & (g16) & (g17)) + ((shiftx2x) & (!shiftx3x) & (g13) & (!g14) & (!g16) & (!g17)) + ((shiftx2x) & (!shiftx3x) & (g13) & (!g14) & (!g16) & (g17)) + ((shiftx2x) & (!shiftx3x) & (g13) & (!g14) & (g16) & (!g17)) + ((shiftx2x) & (!shiftx3x) & (g13) & (!g14) & (g16) & (g17)) + ((shiftx2x) & (!shiftx3x) & (g13) & (g14) & (!g16) & (!g17)) + ((shiftx2x) & (!shiftx3x) & (g13) & (g14) & (!g16) & (g17)) + ((shiftx2x) & (!shiftx3x) & (g13) & (g14) & (g16) & (!g17)) + ((shiftx2x) & (!shiftx3x) & (g13) & (g14) & (g16) & (g17)) + ((shiftx2x) & (shiftx3x) & (!g13) & (!g14) & (!g16) & (g17)) + ((shiftx2x) & (shiftx3x) & (!g13) & (!g14) & (g16) & (g17)) + ((shiftx2x) & (shiftx3x) & (!g13) & (g14) & (!g16) & (g17)) + ((shiftx2x) & (shiftx3x) & (!g13) & (g14) & (g16) & (g17)) + ((shiftx2x) & (shiftx3x) & (g13) & (!g14) & (!g16) & (g17)) + ((shiftx2x) & (shiftx3x) & (g13) & (!g14) & (g16) & (g17)) + ((shiftx2x) & (shiftx3x) & (g13) & (g14) & (!g16) & (g17)) + ((shiftx2x) & (shiftx3x) & (g13) & (g14) & (g16) & (g17)));
	assign g218 = (((!shiftx2x) & (!shiftx3x) & (!g11) & (!g12) & (!g24) & (g25)) + ((!shiftx2x) & (!shiftx3x) & (!g11) & (!g12) & (g24) & (g25)) + ((!shiftx2x) & (!shiftx3x) & (!g11) & (g12) & (!g24) & (g25)) + ((!shiftx2x) & (!shiftx3x) & (!g11) & (g12) & (g24) & (g25)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (!g12) & (!g24) & (g25)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (!g12) & (g24) & (g25)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (g12) & (!g24) & (g25)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (g12) & (g24) & (g25)) + ((!shiftx2x) & (shiftx3x) & (g11) & (!g12) & (!g24) & (!g25)) + ((!shiftx2x) & (shiftx3x) & (g11) & (!g12) & (!g24) & (g25)) + ((!shiftx2x) & (shiftx3x) & (g11) & (!g12) & (g24) & (!g25)) + ((!shiftx2x) & (shiftx3x) & (g11) & (!g12) & (g24) & (g25)) + ((!shiftx2x) & (shiftx3x) & (g11) & (g12) & (!g24) & (!g25)) + ((!shiftx2x) & (shiftx3x) & (g11) & (g12) & (!g24) & (g25)) + ((!shiftx2x) & (shiftx3x) & (g11) & (g12) & (g24) & (!g25)) + ((!shiftx2x) & (shiftx3x) & (g11) & (g12) & (g24) & (g25)) + ((shiftx2x) & (!shiftx3x) & (!g11) & (!g12) & (g24) & (!g25)) + ((shiftx2x) & (!shiftx3x) & (!g11) & (!g12) & (g24) & (g25)) + ((shiftx2x) & (!shiftx3x) & (!g11) & (g12) & (g24) & (!g25)) + ((shiftx2x) & (!shiftx3x) & (!g11) & (g12) & (g24) & (g25)) + ((shiftx2x) & (!shiftx3x) & (g11) & (!g12) & (g24) & (!g25)) + ((shiftx2x) & (!shiftx3x) & (g11) & (!g12) & (g24) & (g25)) + ((shiftx2x) & (!shiftx3x) & (g11) & (g12) & (g24) & (!g25)) + ((shiftx2x) & (!shiftx3x) & (g11) & (g12) & (g24) & (g25)) + ((shiftx2x) & (shiftx3x) & (!g11) & (g12) & (!g24) & (!g25)) + ((shiftx2x) & (shiftx3x) & (!g11) & (g12) & (!g24) & (g25)) + ((shiftx2x) & (shiftx3x) & (!g11) & (g12) & (g24) & (!g25)) + ((shiftx2x) & (shiftx3x) & (!g11) & (g12) & (g24) & (g25)) + ((shiftx2x) & (shiftx3x) & (g11) & (g12) & (!g24) & (!g25)) + ((shiftx2x) & (shiftx3x) & (g11) & (g12) & (!g24) & (g25)) + ((shiftx2x) & (shiftx3x) & (g11) & (g12) & (g24) & (!g25)) + ((shiftx2x) & (shiftx3x) & (g11) & (g12) & (g24) & (g25)));
	assign g219 = (((!shiftx2x) & (!shiftx3x) & (!g6) & (!g7) & (!g18) & (g19)) + ((!shiftx2x) & (!shiftx3x) & (!g6) & (!g7) & (g18) & (g19)) + ((!shiftx2x) & (!shiftx3x) & (!g6) & (g7) & (!g18) & (g19)) + ((!shiftx2x) & (!shiftx3x) & (!g6) & (g7) & (g18) & (g19)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (!g7) & (!g18) & (g19)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (!g7) & (g18) & (g19)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (g7) & (!g18) & (g19)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (g7) & (g18) & (g19)) + ((!shiftx2x) & (shiftx3x) & (g6) & (!g7) & (!g18) & (!g19)) + ((!shiftx2x) & (shiftx3x) & (g6) & (!g7) & (!g18) & (g19)) + ((!shiftx2x) & (shiftx3x) & (g6) & (!g7) & (g18) & (!g19)) + ((!shiftx2x) & (shiftx3x) & (g6) & (!g7) & (g18) & (g19)) + ((!shiftx2x) & (shiftx3x) & (g6) & (g7) & (!g18) & (!g19)) + ((!shiftx2x) & (shiftx3x) & (g6) & (g7) & (!g18) & (g19)) + ((!shiftx2x) & (shiftx3x) & (g6) & (g7) & (g18) & (!g19)) + ((!shiftx2x) & (shiftx3x) & (g6) & (g7) & (g18) & (g19)) + ((shiftx2x) & (!shiftx3x) & (!g6) & (!g7) & (g18) & (!g19)) + ((shiftx2x) & (!shiftx3x) & (!g6) & (!g7) & (g18) & (g19)) + ((shiftx2x) & (!shiftx3x) & (!g6) & (g7) & (g18) & (!g19)) + ((shiftx2x) & (!shiftx3x) & (!g6) & (g7) & (g18) & (g19)) + ((shiftx2x) & (!shiftx3x) & (g6) & (!g7) & (g18) & (!g19)) + ((shiftx2x) & (!shiftx3x) & (g6) & (!g7) & (g18) & (g19)) + ((shiftx2x) & (!shiftx3x) & (g6) & (g7) & (g18) & (!g19)) + ((shiftx2x) & (!shiftx3x) & (g6) & (g7) & (g18) & (g19)) + ((shiftx2x) & (shiftx3x) & (!g6) & (g7) & (!g18) & (!g19)) + ((shiftx2x) & (shiftx3x) & (!g6) & (g7) & (!g18) & (g19)) + ((shiftx2x) & (shiftx3x) & (!g6) & (g7) & (g18) & (!g19)) + ((shiftx2x) & (shiftx3x) & (!g6) & (g7) & (g18) & (g19)) + ((shiftx2x) & (shiftx3x) & (g6) & (g7) & (!g18) & (!g19)) + ((shiftx2x) & (shiftx3x) & (g6) & (g7) & (!g18) & (g19)) + ((shiftx2x) & (shiftx3x) & (g6) & (g7) & (g18) & (!g19)) + ((shiftx2x) & (shiftx3x) & (g6) & (g7) & (g18) & (g19)));
	assign g220 = (((!shiftx2x) & (!shiftx3x) & (!g1) & (!g2) & (!g8) & (g9)) + ((!shiftx2x) & (!shiftx3x) & (!g1) & (!g2) & (g8) & (g9)) + ((!shiftx2x) & (!shiftx3x) & (!g1) & (g2) & (!g8) & (g9)) + ((!shiftx2x) & (!shiftx3x) & (!g1) & (g2) & (g8) & (g9)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (!g2) & (!g8) & (g9)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (!g2) & (g8) & (g9)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (g2) & (!g8) & (g9)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (g2) & (g8) & (g9)) + ((!shiftx2x) & (shiftx3x) & (g1) & (!g2) & (!g8) & (!g9)) + ((!shiftx2x) & (shiftx3x) & (g1) & (!g2) & (!g8) & (g9)) + ((!shiftx2x) & (shiftx3x) & (g1) & (!g2) & (g8) & (!g9)) + ((!shiftx2x) & (shiftx3x) & (g1) & (!g2) & (g8) & (g9)) + ((!shiftx2x) & (shiftx3x) & (g1) & (g2) & (!g8) & (!g9)) + ((!shiftx2x) & (shiftx3x) & (g1) & (g2) & (!g8) & (g9)) + ((!shiftx2x) & (shiftx3x) & (g1) & (g2) & (g8) & (!g9)) + ((!shiftx2x) & (shiftx3x) & (g1) & (g2) & (g8) & (g9)) + ((shiftx2x) & (!shiftx3x) & (!g1) & (!g2) & (g8) & (!g9)) + ((shiftx2x) & (!shiftx3x) & (!g1) & (!g2) & (g8) & (g9)) + ((shiftx2x) & (!shiftx3x) & (!g1) & (g2) & (g8) & (!g9)) + ((shiftx2x) & (!shiftx3x) & (!g1) & (g2) & (g8) & (g9)) + ((shiftx2x) & (!shiftx3x) & (g1) & (!g2) & (g8) & (!g9)) + ((shiftx2x) & (!shiftx3x) & (g1) & (!g2) & (g8) & (g9)) + ((shiftx2x) & (!shiftx3x) & (g1) & (g2) & (g8) & (!g9)) + ((shiftx2x) & (!shiftx3x) & (g1) & (g2) & (g8) & (g9)) + ((shiftx2x) & (shiftx3x) & (!g1) & (g2) & (!g8) & (!g9)) + ((shiftx2x) & (shiftx3x) & (!g1) & (g2) & (!g8) & (g9)) + ((shiftx2x) & (shiftx3x) & (!g1) & (g2) & (g8) & (!g9)) + ((shiftx2x) & (shiftx3x) & (!g1) & (g2) & (g8) & (g9)) + ((shiftx2x) & (shiftx3x) & (g1) & (g2) & (!g8) & (!g9)) + ((shiftx2x) & (shiftx3x) & (g1) & (g2) & (!g8) & (g9)) + ((shiftx2x) & (shiftx3x) & (g1) & (g2) & (g8) & (!g9)) + ((shiftx2x) & (shiftx3x) & (g1) & (g2) & (g8) & (g9)));
	assign g221 = (((!shiftx4x) & (!shiftx5x) & (!g217) & (g218) & (!g219) & (!g220)) + ((!shiftx4x) & (!shiftx5x) & (!g217) & (g218) & (!g219) & (g220)) + ((!shiftx4x) & (!shiftx5x) & (!g217) & (g218) & (g219) & (!g220)) + ((!shiftx4x) & (!shiftx5x) & (!g217) & (g218) & (g219) & (g220)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (g218) & (!g219) & (!g220)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (g218) & (!g219) & (g220)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (g218) & (g219) & (!g220)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (g218) & (g219) & (g220)) + ((!shiftx4x) & (shiftx5x) & (!g217) & (!g218) & (g219) & (!g220)) + ((!shiftx4x) & (shiftx5x) & (!g217) & (!g218) & (g219) & (g220)) + ((!shiftx4x) & (shiftx5x) & (!g217) & (g218) & (g219) & (!g220)) + ((!shiftx4x) & (shiftx5x) & (!g217) & (g218) & (g219) & (g220)) + ((!shiftx4x) & (shiftx5x) & (g217) & (!g218) & (g219) & (!g220)) + ((!shiftx4x) & (shiftx5x) & (g217) & (!g218) & (g219) & (g220)) + ((!shiftx4x) & (shiftx5x) & (g217) & (g218) & (g219) & (!g220)) + ((!shiftx4x) & (shiftx5x) & (g217) & (g218) & (g219) & (g220)) + ((shiftx4x) & (!shiftx5x) & (g217) & (!g218) & (!g219) & (!g220)) + ((shiftx4x) & (!shiftx5x) & (g217) & (!g218) & (!g219) & (g220)) + ((shiftx4x) & (!shiftx5x) & (g217) & (!g218) & (g219) & (!g220)) + ((shiftx4x) & (!shiftx5x) & (g217) & (!g218) & (g219) & (g220)) + ((shiftx4x) & (!shiftx5x) & (g217) & (g218) & (!g219) & (!g220)) + ((shiftx4x) & (!shiftx5x) & (g217) & (g218) & (!g219) & (g220)) + ((shiftx4x) & (!shiftx5x) & (g217) & (g218) & (g219) & (!g220)) + ((shiftx4x) & (!shiftx5x) & (g217) & (g218) & (g219) & (g220)) + ((shiftx4x) & (shiftx5x) & (!g217) & (!g218) & (!g219) & (g220)) + ((shiftx4x) & (shiftx5x) & (!g217) & (!g218) & (g219) & (g220)) + ((shiftx4x) & (shiftx5x) & (!g217) & (g218) & (!g219) & (g220)) + ((shiftx4x) & (shiftx5x) & (!g217) & (g218) & (g219) & (g220)) + ((shiftx4x) & (shiftx5x) & (g217) & (!g218) & (!g219) & (g220)) + ((shiftx4x) & (shiftx5x) & (g217) & (!g218) & (g219) & (g220)) + ((shiftx4x) & (shiftx5x) & (g217) & (g218) & (!g219) & (g220)) + ((shiftx4x) & (shiftx5x) & (g217) & (g218) & (g219) & (g220)));
	assign g222 = (((!shiftx2x) & (!shiftx3x) & (!g22) & (!g23) & (!g29) & (g30)) + ((!shiftx2x) & (!shiftx3x) & (!g22) & (!g23) & (g29) & (g30)) + ((!shiftx2x) & (!shiftx3x) & (!g22) & (g23) & (!g29) & (g30)) + ((!shiftx2x) & (!shiftx3x) & (!g22) & (g23) & (g29) & (g30)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (!g23) & (!g29) & (g30)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (!g23) & (g29) & (g30)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (g23) & (!g29) & (g30)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (g23) & (g29) & (g30)) + ((!shiftx2x) & (shiftx3x) & (g22) & (!g23) & (!g29) & (!g30)) + ((!shiftx2x) & (shiftx3x) & (g22) & (!g23) & (!g29) & (g30)) + ((!shiftx2x) & (shiftx3x) & (g22) & (!g23) & (g29) & (!g30)) + ((!shiftx2x) & (shiftx3x) & (g22) & (!g23) & (g29) & (g30)) + ((!shiftx2x) & (shiftx3x) & (g22) & (g23) & (!g29) & (!g30)) + ((!shiftx2x) & (shiftx3x) & (g22) & (g23) & (!g29) & (g30)) + ((!shiftx2x) & (shiftx3x) & (g22) & (g23) & (g29) & (!g30)) + ((!shiftx2x) & (shiftx3x) & (g22) & (g23) & (g29) & (g30)) + ((shiftx2x) & (!shiftx3x) & (!g22) & (!g23) & (g29) & (!g30)) + ((shiftx2x) & (!shiftx3x) & (!g22) & (!g23) & (g29) & (g30)) + ((shiftx2x) & (!shiftx3x) & (!g22) & (g23) & (g29) & (!g30)) + ((shiftx2x) & (!shiftx3x) & (!g22) & (g23) & (g29) & (g30)) + ((shiftx2x) & (!shiftx3x) & (g22) & (!g23) & (g29) & (!g30)) + ((shiftx2x) & (!shiftx3x) & (g22) & (!g23) & (g29) & (g30)) + ((shiftx2x) & (!shiftx3x) & (g22) & (g23) & (g29) & (!g30)) + ((shiftx2x) & (!shiftx3x) & (g22) & (g23) & (g29) & (g30)) + ((shiftx2x) & (shiftx3x) & (!g22) & (g23) & (!g29) & (!g30)) + ((shiftx2x) & (shiftx3x) & (!g22) & (g23) & (!g29) & (g30)) + ((shiftx2x) & (shiftx3x) & (!g22) & (g23) & (g29) & (!g30)) + ((shiftx2x) & (shiftx3x) & (!g22) & (g23) & (g29) & (g30)) + ((shiftx2x) & (shiftx3x) & (g22) & (g23) & (!g29) & (!g30)) + ((shiftx2x) & (shiftx3x) & (g22) & (g23) & (!g29) & (g30)) + ((shiftx2x) & (shiftx3x) & (g22) & (g23) & (g29) & (!g30)) + ((shiftx2x) & (shiftx3x) & (g22) & (g23) & (g29) & (g30)));
	assign g223 = (((!shiftx2x) & (!shiftx3x) & (!g27) & (!g28) & (!g39) & (g40)) + ((!shiftx2x) & (!shiftx3x) & (!g27) & (!g28) & (g39) & (g40)) + ((!shiftx2x) & (!shiftx3x) & (!g27) & (g28) & (!g39) & (g40)) + ((!shiftx2x) & (!shiftx3x) & (!g27) & (g28) & (g39) & (g40)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (!g28) & (!g39) & (g40)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (!g28) & (g39) & (g40)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (g28) & (!g39) & (g40)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (g28) & (g39) & (g40)) + ((!shiftx2x) & (shiftx3x) & (g27) & (!g28) & (!g39) & (!g40)) + ((!shiftx2x) & (shiftx3x) & (g27) & (!g28) & (!g39) & (g40)) + ((!shiftx2x) & (shiftx3x) & (g27) & (!g28) & (g39) & (!g40)) + ((!shiftx2x) & (shiftx3x) & (g27) & (!g28) & (g39) & (g40)) + ((!shiftx2x) & (shiftx3x) & (g27) & (g28) & (!g39) & (!g40)) + ((!shiftx2x) & (shiftx3x) & (g27) & (g28) & (!g39) & (g40)) + ((!shiftx2x) & (shiftx3x) & (g27) & (g28) & (g39) & (!g40)) + ((!shiftx2x) & (shiftx3x) & (g27) & (g28) & (g39) & (g40)) + ((shiftx2x) & (!shiftx3x) & (!g27) & (!g28) & (g39) & (!g40)) + ((shiftx2x) & (!shiftx3x) & (!g27) & (!g28) & (g39) & (g40)) + ((shiftx2x) & (!shiftx3x) & (!g27) & (g28) & (g39) & (!g40)) + ((shiftx2x) & (!shiftx3x) & (!g27) & (g28) & (g39) & (g40)) + ((shiftx2x) & (!shiftx3x) & (g27) & (!g28) & (g39) & (!g40)) + ((shiftx2x) & (!shiftx3x) & (g27) & (!g28) & (g39) & (g40)) + ((shiftx2x) & (!shiftx3x) & (g27) & (g28) & (g39) & (!g40)) + ((shiftx2x) & (!shiftx3x) & (g27) & (g28) & (g39) & (g40)) + ((shiftx2x) & (shiftx3x) & (!g27) & (g28) & (!g39) & (!g40)) + ((shiftx2x) & (shiftx3x) & (!g27) & (g28) & (!g39) & (g40)) + ((shiftx2x) & (shiftx3x) & (!g27) & (g28) & (g39) & (!g40)) + ((shiftx2x) & (shiftx3x) & (!g27) & (g28) & (g39) & (g40)) + ((shiftx2x) & (shiftx3x) & (g27) & (g28) & (!g39) & (!g40)) + ((shiftx2x) & (shiftx3x) & (g27) & (g28) & (!g39) & (g40)) + ((shiftx2x) & (shiftx3x) & (g27) & (g28) & (g39) & (!g40)) + ((shiftx2x) & (shiftx3x) & (g27) & (g28) & (g39) & (g40)));
	assign g224 = (((!shiftx2x) & (!shiftx3x) & (!g3) & (g4) & (!g32) & (!g33)) + ((!shiftx2x) & (!shiftx3x) & (!g3) & (g4) & (!g32) & (g33)) + ((!shiftx2x) & (!shiftx3x) & (!g3) & (g4) & (g32) & (!g33)) + ((!shiftx2x) & (!shiftx3x) & (!g3) & (g4) & (g32) & (g33)) + ((!shiftx2x) & (!shiftx3x) & (g3) & (g4) & (!g32) & (!g33)) + ((!shiftx2x) & (!shiftx3x) & (g3) & (g4) & (!g32) & (g33)) + ((!shiftx2x) & (!shiftx3x) & (g3) & (g4) & (g32) & (!g33)) + ((!shiftx2x) & (!shiftx3x) & (g3) & (g4) & (g32) & (g33)) + ((!shiftx2x) & (shiftx3x) & (!g3) & (!g4) & (g32) & (!g33)) + ((!shiftx2x) & (shiftx3x) & (!g3) & (!g4) & (g32) & (g33)) + ((!shiftx2x) & (shiftx3x) & (!g3) & (g4) & (g32) & (!g33)) + ((!shiftx2x) & (shiftx3x) & (!g3) & (g4) & (g32) & (g33)) + ((!shiftx2x) & (shiftx3x) & (g3) & (!g4) & (g32) & (!g33)) + ((!shiftx2x) & (shiftx3x) & (g3) & (!g4) & (g32) & (g33)) + ((!shiftx2x) & (shiftx3x) & (g3) & (g4) & (g32) & (!g33)) + ((!shiftx2x) & (shiftx3x) & (g3) & (g4) & (g32) & (g33)) + ((shiftx2x) & (!shiftx3x) & (g3) & (!g4) & (!g32) & (!g33)) + ((shiftx2x) & (!shiftx3x) & (g3) & (!g4) & (!g32) & (g33)) + ((shiftx2x) & (!shiftx3x) & (g3) & (!g4) & (g32) & (!g33)) + ((shiftx2x) & (!shiftx3x) & (g3) & (!g4) & (g32) & (g33)) + ((shiftx2x) & (!shiftx3x) & (g3) & (g4) & (!g32) & (!g33)) + ((shiftx2x) & (!shiftx3x) & (g3) & (g4) & (!g32) & (g33)) + ((shiftx2x) & (!shiftx3x) & (g3) & (g4) & (g32) & (!g33)) + ((shiftx2x) & (!shiftx3x) & (g3) & (g4) & (g32) & (g33)) + ((shiftx2x) & (shiftx3x) & (!g3) & (!g4) & (!g32) & (g33)) + ((shiftx2x) & (shiftx3x) & (!g3) & (!g4) & (g32) & (g33)) + ((shiftx2x) & (shiftx3x) & (!g3) & (g4) & (!g32) & (g33)) + ((shiftx2x) & (shiftx3x) & (!g3) & (g4) & (g32) & (g33)) + ((shiftx2x) & (shiftx3x) & (g3) & (!g4) & (!g32) & (g33)) + ((shiftx2x) & (shiftx3x) & (g3) & (!g4) & (g32) & (g33)) + ((shiftx2x) & (shiftx3x) & (g3) & (g4) & (!g32) & (g33)) + ((shiftx2x) & (shiftx3x) & (g3) & (g4) & (g32) & (g33)));
	assign g225 = (((!shiftx2x) & (!shiftx3x) & (!g34) & (g35) & (!g37) & (!g38)) + ((!shiftx2x) & (!shiftx3x) & (!g34) & (g35) & (!g37) & (g38)) + ((!shiftx2x) & (!shiftx3x) & (!g34) & (g35) & (g37) & (!g38)) + ((!shiftx2x) & (!shiftx3x) & (!g34) & (g35) & (g37) & (g38)) + ((!shiftx2x) & (!shiftx3x) & (g34) & (g35) & (!g37) & (!g38)) + ((!shiftx2x) & (!shiftx3x) & (g34) & (g35) & (!g37) & (g38)) + ((!shiftx2x) & (!shiftx3x) & (g34) & (g35) & (g37) & (!g38)) + ((!shiftx2x) & (!shiftx3x) & (g34) & (g35) & (g37) & (g38)) + ((!shiftx2x) & (shiftx3x) & (!g34) & (!g35) & (g37) & (!g38)) + ((!shiftx2x) & (shiftx3x) & (!g34) & (!g35) & (g37) & (g38)) + ((!shiftx2x) & (shiftx3x) & (!g34) & (g35) & (g37) & (!g38)) + ((!shiftx2x) & (shiftx3x) & (!g34) & (g35) & (g37) & (g38)) + ((!shiftx2x) & (shiftx3x) & (g34) & (!g35) & (g37) & (!g38)) + ((!shiftx2x) & (shiftx3x) & (g34) & (!g35) & (g37) & (g38)) + ((!shiftx2x) & (shiftx3x) & (g34) & (g35) & (g37) & (!g38)) + ((!shiftx2x) & (shiftx3x) & (g34) & (g35) & (g37) & (g38)) + ((shiftx2x) & (!shiftx3x) & (g34) & (!g35) & (!g37) & (!g38)) + ((shiftx2x) & (!shiftx3x) & (g34) & (!g35) & (!g37) & (g38)) + ((shiftx2x) & (!shiftx3x) & (g34) & (!g35) & (g37) & (!g38)) + ((shiftx2x) & (!shiftx3x) & (g34) & (!g35) & (g37) & (g38)) + ((shiftx2x) & (!shiftx3x) & (g34) & (g35) & (!g37) & (!g38)) + ((shiftx2x) & (!shiftx3x) & (g34) & (g35) & (!g37) & (g38)) + ((shiftx2x) & (!shiftx3x) & (g34) & (g35) & (g37) & (!g38)) + ((shiftx2x) & (!shiftx3x) & (g34) & (g35) & (g37) & (g38)) + ((shiftx2x) & (shiftx3x) & (!g34) & (!g35) & (!g37) & (g38)) + ((shiftx2x) & (shiftx3x) & (!g34) & (!g35) & (g37) & (g38)) + ((shiftx2x) & (shiftx3x) & (!g34) & (g35) & (!g37) & (g38)) + ((shiftx2x) & (shiftx3x) & (!g34) & (g35) & (g37) & (g38)) + ((shiftx2x) & (shiftx3x) & (g34) & (!g35) & (!g37) & (g38)) + ((shiftx2x) & (shiftx3x) & (g34) & (!g35) & (g37) & (g38)) + ((shiftx2x) & (shiftx3x) & (g34) & (g35) & (!g37) & (g38)) + ((shiftx2x) & (shiftx3x) & (g34) & (g35) & (g37) & (g38)));
	assign g226 = (((!shiftx4x) & (!shiftx5x) & (!g222) & (!g223) & (g224) & (!g225)) + ((!shiftx4x) & (!shiftx5x) & (!g222) & (!g223) & (g224) & (g225)) + ((!shiftx4x) & (!shiftx5x) & (!g222) & (g223) & (g224) & (!g225)) + ((!shiftx4x) & (!shiftx5x) & (!g222) & (g223) & (g224) & (g225)) + ((!shiftx4x) & (!shiftx5x) & (g222) & (!g223) & (g224) & (!g225)) + ((!shiftx4x) & (!shiftx5x) & (g222) & (!g223) & (g224) & (g225)) + ((!shiftx4x) & (!shiftx5x) & (g222) & (g223) & (g224) & (!g225)) + ((!shiftx4x) & (!shiftx5x) & (g222) & (g223) & (g224) & (g225)) + ((!shiftx4x) & (shiftx5x) & (!g222) & (g223) & (!g224) & (!g225)) + ((!shiftx4x) & (shiftx5x) & (!g222) & (g223) & (!g224) & (g225)) + ((!shiftx4x) & (shiftx5x) & (!g222) & (g223) & (g224) & (!g225)) + ((!shiftx4x) & (shiftx5x) & (!g222) & (g223) & (g224) & (g225)) + ((!shiftx4x) & (shiftx5x) & (g222) & (g223) & (!g224) & (!g225)) + ((!shiftx4x) & (shiftx5x) & (g222) & (g223) & (!g224) & (g225)) + ((!shiftx4x) & (shiftx5x) & (g222) & (g223) & (g224) & (!g225)) + ((!shiftx4x) & (shiftx5x) & (g222) & (g223) & (g224) & (g225)) + ((shiftx4x) & (!shiftx5x) & (!g222) & (!g223) & (!g224) & (g225)) + ((shiftx4x) & (!shiftx5x) & (!g222) & (!g223) & (g224) & (g225)) + ((shiftx4x) & (!shiftx5x) & (!g222) & (g223) & (!g224) & (g225)) + ((shiftx4x) & (!shiftx5x) & (!g222) & (g223) & (g224) & (g225)) + ((shiftx4x) & (!shiftx5x) & (g222) & (!g223) & (!g224) & (g225)) + ((shiftx4x) & (!shiftx5x) & (g222) & (!g223) & (g224) & (g225)) + ((shiftx4x) & (!shiftx5x) & (g222) & (g223) & (!g224) & (g225)) + ((shiftx4x) & (!shiftx5x) & (g222) & (g223) & (g224) & (g225)) + ((shiftx4x) & (shiftx5x) & (g222) & (!g223) & (!g224) & (!g225)) + ((shiftx4x) & (shiftx5x) & (g222) & (!g223) & (!g224) & (g225)) + ((shiftx4x) & (shiftx5x) & (g222) & (!g223) & (g224) & (!g225)) + ((shiftx4x) & (shiftx5x) & (g222) & (!g223) & (g224) & (g225)) + ((shiftx4x) & (shiftx5x) & (g222) & (g223) & (!g224) & (!g225)) + ((shiftx4x) & (shiftx5x) & (g222) & (g223) & (!g224) & (g225)) + ((shiftx4x) & (shiftx5x) & (g222) & (g223) & (g224) & (!g225)) + ((shiftx4x) & (shiftx5x) & (g222) & (g223) & (g224) & (g225)));
	assign resultx8x = (((!shiftx6x) & (sk[98]) & (!g221) & (g226)) + ((!shiftx6x) & (sk[98]) & (g221) & (g226)) + ((shiftx6x) & (!sk[98]) & (!g221) & (!g226)) + ((shiftx6x) & (!sk[98]) & (!g221) & (g226)) + ((shiftx6x) & (!sk[98]) & (g221) & (!g226)) + ((shiftx6x) & (!sk[98]) & (g221) & (g226)) + ((shiftx6x) & (sk[98]) & (g221) & (!g226)) + ((shiftx6x) & (sk[98]) & (g221) & (g226)));
	assign g228 = (((!shiftx2x) & (!shiftx3x) & (!g46) & (g47) & (!g54) & (!g55)) + ((!shiftx2x) & (!shiftx3x) & (!g46) & (g47) & (!g54) & (g55)) + ((!shiftx2x) & (!shiftx3x) & (!g46) & (g47) & (g54) & (!g55)) + ((!shiftx2x) & (!shiftx3x) & (!g46) & (g47) & (g54) & (g55)) + ((!shiftx2x) & (!shiftx3x) & (g46) & (g47) & (!g54) & (!g55)) + ((!shiftx2x) & (!shiftx3x) & (g46) & (g47) & (!g54) & (g55)) + ((!shiftx2x) & (!shiftx3x) & (g46) & (g47) & (g54) & (!g55)) + ((!shiftx2x) & (!shiftx3x) & (g46) & (g47) & (g54) & (g55)) + ((!shiftx2x) & (shiftx3x) & (!g46) & (!g47) & (g54) & (!g55)) + ((!shiftx2x) & (shiftx3x) & (!g46) & (!g47) & (g54) & (g55)) + ((!shiftx2x) & (shiftx3x) & (!g46) & (g47) & (g54) & (!g55)) + ((!shiftx2x) & (shiftx3x) & (!g46) & (g47) & (g54) & (g55)) + ((!shiftx2x) & (shiftx3x) & (g46) & (!g47) & (g54) & (!g55)) + ((!shiftx2x) & (shiftx3x) & (g46) & (!g47) & (g54) & (g55)) + ((!shiftx2x) & (shiftx3x) & (g46) & (g47) & (g54) & (!g55)) + ((!shiftx2x) & (shiftx3x) & (g46) & (g47) & (g54) & (g55)) + ((shiftx2x) & (!shiftx3x) & (g46) & (!g47) & (!g54) & (!g55)) + ((shiftx2x) & (!shiftx3x) & (g46) & (!g47) & (!g54) & (g55)) + ((shiftx2x) & (!shiftx3x) & (g46) & (!g47) & (g54) & (!g55)) + ((shiftx2x) & (!shiftx3x) & (g46) & (!g47) & (g54) & (g55)) + ((shiftx2x) & (!shiftx3x) & (g46) & (g47) & (!g54) & (!g55)) + ((shiftx2x) & (!shiftx3x) & (g46) & (g47) & (!g54) & (g55)) + ((shiftx2x) & (!shiftx3x) & (g46) & (g47) & (g54) & (!g55)) + ((shiftx2x) & (!shiftx3x) & (g46) & (g47) & (g54) & (g55)) + ((shiftx2x) & (shiftx3x) & (!g46) & (!g47) & (!g54) & (g55)) + ((shiftx2x) & (shiftx3x) & (!g46) & (!g47) & (g54) & (g55)) + ((shiftx2x) & (shiftx3x) & (!g46) & (g47) & (!g54) & (g55)) + ((shiftx2x) & (shiftx3x) & (!g46) & (g47) & (g54) & (g55)) + ((shiftx2x) & (shiftx3x) & (g46) & (!g47) & (!g54) & (g55)) + ((shiftx2x) & (shiftx3x) & (g46) & (!g47) & (g54) & (g55)) + ((shiftx2x) & (shiftx3x) & (g46) & (g47) & (!g54) & (g55)) + ((shiftx2x) & (shiftx3x) & (g46) & (g47) & (g54) & (g55)));
	assign g229 = (((!shiftx2x) & (!shiftx3x) & (!g44) & (!g45) & (!g67) & (g68)) + ((!shiftx2x) & (!shiftx3x) & (!g44) & (!g45) & (g67) & (g68)) + ((!shiftx2x) & (!shiftx3x) & (!g44) & (g45) & (!g67) & (g68)) + ((!shiftx2x) & (!shiftx3x) & (!g44) & (g45) & (g67) & (g68)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (!g45) & (!g67) & (g68)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (!g45) & (g67) & (g68)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (g45) & (!g67) & (g68)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (g45) & (g67) & (g68)) + ((!shiftx2x) & (shiftx3x) & (g44) & (!g45) & (!g67) & (!g68)) + ((!shiftx2x) & (shiftx3x) & (g44) & (!g45) & (!g67) & (g68)) + ((!shiftx2x) & (shiftx3x) & (g44) & (!g45) & (g67) & (!g68)) + ((!shiftx2x) & (shiftx3x) & (g44) & (!g45) & (g67) & (g68)) + ((!shiftx2x) & (shiftx3x) & (g44) & (g45) & (!g67) & (!g68)) + ((!shiftx2x) & (shiftx3x) & (g44) & (g45) & (!g67) & (g68)) + ((!shiftx2x) & (shiftx3x) & (g44) & (g45) & (g67) & (!g68)) + ((!shiftx2x) & (shiftx3x) & (g44) & (g45) & (g67) & (g68)) + ((shiftx2x) & (!shiftx3x) & (!g44) & (!g45) & (g67) & (!g68)) + ((shiftx2x) & (!shiftx3x) & (!g44) & (!g45) & (g67) & (g68)) + ((shiftx2x) & (!shiftx3x) & (!g44) & (g45) & (g67) & (!g68)) + ((shiftx2x) & (!shiftx3x) & (!g44) & (g45) & (g67) & (g68)) + ((shiftx2x) & (!shiftx3x) & (g44) & (!g45) & (g67) & (!g68)) + ((shiftx2x) & (!shiftx3x) & (g44) & (!g45) & (g67) & (g68)) + ((shiftx2x) & (!shiftx3x) & (g44) & (g45) & (g67) & (!g68)) + ((shiftx2x) & (!shiftx3x) & (g44) & (g45) & (g67) & (g68)) + ((shiftx2x) & (shiftx3x) & (!g44) & (g45) & (!g67) & (!g68)) + ((shiftx2x) & (shiftx3x) & (!g44) & (g45) & (!g67) & (g68)) + ((shiftx2x) & (shiftx3x) & (!g44) & (g45) & (g67) & (!g68)) + ((shiftx2x) & (shiftx3x) & (!g44) & (g45) & (g67) & (g68)) + ((shiftx2x) & (shiftx3x) & (g44) & (g45) & (!g67) & (!g68)) + ((shiftx2x) & (shiftx3x) & (g44) & (g45) & (!g67) & (g68)) + ((shiftx2x) & (shiftx3x) & (g44) & (g45) & (g67) & (!g68)) + ((shiftx2x) & (shiftx3x) & (g44) & (g45) & (g67) & (g68)));
	assign g230 = (((!shiftx2x) & (!shiftx3x) & (!g56) & (g57) & (!g59) & (!g60)) + ((!shiftx2x) & (!shiftx3x) & (!g56) & (g57) & (!g59) & (g60)) + ((!shiftx2x) & (!shiftx3x) & (!g56) & (g57) & (g59) & (!g60)) + ((!shiftx2x) & (!shiftx3x) & (!g56) & (g57) & (g59) & (g60)) + ((!shiftx2x) & (!shiftx3x) & (g56) & (g57) & (!g59) & (!g60)) + ((!shiftx2x) & (!shiftx3x) & (g56) & (g57) & (!g59) & (g60)) + ((!shiftx2x) & (!shiftx3x) & (g56) & (g57) & (g59) & (!g60)) + ((!shiftx2x) & (!shiftx3x) & (g56) & (g57) & (g59) & (g60)) + ((!shiftx2x) & (shiftx3x) & (!g56) & (!g57) & (g59) & (!g60)) + ((!shiftx2x) & (shiftx3x) & (!g56) & (!g57) & (g59) & (g60)) + ((!shiftx2x) & (shiftx3x) & (!g56) & (g57) & (g59) & (!g60)) + ((!shiftx2x) & (shiftx3x) & (!g56) & (g57) & (g59) & (g60)) + ((!shiftx2x) & (shiftx3x) & (g56) & (!g57) & (g59) & (!g60)) + ((!shiftx2x) & (shiftx3x) & (g56) & (!g57) & (g59) & (g60)) + ((!shiftx2x) & (shiftx3x) & (g56) & (g57) & (g59) & (!g60)) + ((!shiftx2x) & (shiftx3x) & (g56) & (g57) & (g59) & (g60)) + ((shiftx2x) & (!shiftx3x) & (g56) & (!g57) & (!g59) & (!g60)) + ((shiftx2x) & (!shiftx3x) & (g56) & (!g57) & (!g59) & (g60)) + ((shiftx2x) & (!shiftx3x) & (g56) & (!g57) & (g59) & (!g60)) + ((shiftx2x) & (!shiftx3x) & (g56) & (!g57) & (g59) & (g60)) + ((shiftx2x) & (!shiftx3x) & (g56) & (g57) & (!g59) & (!g60)) + ((shiftx2x) & (!shiftx3x) & (g56) & (g57) & (!g59) & (g60)) + ((shiftx2x) & (!shiftx3x) & (g56) & (g57) & (g59) & (!g60)) + ((shiftx2x) & (!shiftx3x) & (g56) & (g57) & (g59) & (g60)) + ((shiftx2x) & (shiftx3x) & (!g56) & (!g57) & (!g59) & (g60)) + ((shiftx2x) & (shiftx3x) & (!g56) & (!g57) & (g59) & (g60)) + ((shiftx2x) & (shiftx3x) & (!g56) & (g57) & (!g59) & (g60)) + ((shiftx2x) & (shiftx3x) & (!g56) & (g57) & (g59) & (g60)) + ((shiftx2x) & (shiftx3x) & (g56) & (!g57) & (!g59) & (g60)) + ((shiftx2x) & (shiftx3x) & (g56) & (!g57) & (g59) & (g60)) + ((shiftx2x) & (shiftx3x) & (g56) & (g57) & (!g59) & (g60)) + ((shiftx2x) & (shiftx3x) & (g56) & (g57) & (g59) & (g60)));
	assign g231 = (((!shiftx2x) & (!shiftx3x) & (!g49) & (!g50) & (!g61) & (g62)) + ((!shiftx2x) & (!shiftx3x) & (!g49) & (!g50) & (g61) & (g62)) + ((!shiftx2x) & (!shiftx3x) & (!g49) & (g50) & (!g61) & (g62)) + ((!shiftx2x) & (!shiftx3x) & (!g49) & (g50) & (g61) & (g62)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (!g50) & (!g61) & (g62)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (!g50) & (g61) & (g62)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (g50) & (!g61) & (g62)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (g50) & (g61) & (g62)) + ((!shiftx2x) & (shiftx3x) & (g49) & (!g50) & (!g61) & (!g62)) + ((!shiftx2x) & (shiftx3x) & (g49) & (!g50) & (!g61) & (g62)) + ((!shiftx2x) & (shiftx3x) & (g49) & (!g50) & (g61) & (!g62)) + ((!shiftx2x) & (shiftx3x) & (g49) & (!g50) & (g61) & (g62)) + ((!shiftx2x) & (shiftx3x) & (g49) & (g50) & (!g61) & (!g62)) + ((!shiftx2x) & (shiftx3x) & (g49) & (g50) & (!g61) & (g62)) + ((!shiftx2x) & (shiftx3x) & (g49) & (g50) & (g61) & (!g62)) + ((!shiftx2x) & (shiftx3x) & (g49) & (g50) & (g61) & (g62)) + ((shiftx2x) & (!shiftx3x) & (!g49) & (!g50) & (g61) & (!g62)) + ((shiftx2x) & (!shiftx3x) & (!g49) & (!g50) & (g61) & (g62)) + ((shiftx2x) & (!shiftx3x) & (!g49) & (g50) & (g61) & (!g62)) + ((shiftx2x) & (!shiftx3x) & (!g49) & (g50) & (g61) & (g62)) + ((shiftx2x) & (!shiftx3x) & (g49) & (!g50) & (g61) & (!g62)) + ((shiftx2x) & (!shiftx3x) & (g49) & (!g50) & (g61) & (g62)) + ((shiftx2x) & (!shiftx3x) & (g49) & (g50) & (g61) & (!g62)) + ((shiftx2x) & (!shiftx3x) & (g49) & (g50) & (g61) & (g62)) + ((shiftx2x) & (shiftx3x) & (!g49) & (g50) & (!g61) & (!g62)) + ((shiftx2x) & (shiftx3x) & (!g49) & (g50) & (!g61) & (g62)) + ((shiftx2x) & (shiftx3x) & (!g49) & (g50) & (g61) & (!g62)) + ((shiftx2x) & (shiftx3x) & (!g49) & (g50) & (g61) & (g62)) + ((shiftx2x) & (shiftx3x) & (g49) & (g50) & (!g61) & (!g62)) + ((shiftx2x) & (shiftx3x) & (g49) & (g50) & (!g61) & (g62)) + ((shiftx2x) & (shiftx3x) & (g49) & (g50) & (g61) & (!g62)) + ((shiftx2x) & (shiftx3x) & (g49) & (g50) & (g61) & (g62)));
	assign g232 = (((!shiftx4x) & (!shiftx5x) & (!g228) & (g229) & (!g230) & (!g231)) + ((!shiftx4x) & (!shiftx5x) & (!g228) & (g229) & (!g230) & (g231)) + ((!shiftx4x) & (!shiftx5x) & (!g228) & (g229) & (g230) & (!g231)) + ((!shiftx4x) & (!shiftx5x) & (!g228) & (g229) & (g230) & (g231)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (g229) & (!g230) & (!g231)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (g229) & (!g230) & (g231)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (g229) & (g230) & (!g231)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (g229) & (g230) & (g231)) + ((!shiftx4x) & (shiftx5x) & (!g228) & (!g229) & (g230) & (!g231)) + ((!shiftx4x) & (shiftx5x) & (!g228) & (!g229) & (g230) & (g231)) + ((!shiftx4x) & (shiftx5x) & (!g228) & (g229) & (g230) & (!g231)) + ((!shiftx4x) & (shiftx5x) & (!g228) & (g229) & (g230) & (g231)) + ((!shiftx4x) & (shiftx5x) & (g228) & (!g229) & (g230) & (!g231)) + ((!shiftx4x) & (shiftx5x) & (g228) & (!g229) & (g230) & (g231)) + ((!shiftx4x) & (shiftx5x) & (g228) & (g229) & (g230) & (!g231)) + ((!shiftx4x) & (shiftx5x) & (g228) & (g229) & (g230) & (g231)) + ((shiftx4x) & (!shiftx5x) & (g228) & (!g229) & (!g230) & (!g231)) + ((shiftx4x) & (!shiftx5x) & (g228) & (!g229) & (!g230) & (g231)) + ((shiftx4x) & (!shiftx5x) & (g228) & (!g229) & (g230) & (!g231)) + ((shiftx4x) & (!shiftx5x) & (g228) & (!g229) & (g230) & (g231)) + ((shiftx4x) & (!shiftx5x) & (g228) & (g229) & (!g230) & (!g231)) + ((shiftx4x) & (!shiftx5x) & (g228) & (g229) & (!g230) & (g231)) + ((shiftx4x) & (!shiftx5x) & (g228) & (g229) & (g230) & (!g231)) + ((shiftx4x) & (!shiftx5x) & (g228) & (g229) & (g230) & (g231)) + ((shiftx4x) & (shiftx5x) & (!g228) & (!g229) & (!g230) & (g231)) + ((shiftx4x) & (shiftx5x) & (!g228) & (!g229) & (g230) & (g231)) + ((shiftx4x) & (shiftx5x) & (!g228) & (g229) & (!g230) & (g231)) + ((shiftx4x) & (shiftx5x) & (!g228) & (g229) & (g230) & (g231)) + ((shiftx4x) & (shiftx5x) & (g228) & (!g229) & (!g230) & (g231)) + ((shiftx4x) & (shiftx5x) & (g228) & (!g229) & (g230) & (g231)) + ((shiftx4x) & (shiftx5x) & (g228) & (g229) & (!g230) & (g231)) + ((shiftx4x) & (shiftx5x) & (g228) & (g229) & (g230) & (g231)));
	assign g233 = (((!shiftx2x) & (!shiftx3x) & (!g65) & (!g66) & (!g72) & (g73)) + ((!shiftx2x) & (!shiftx3x) & (!g65) & (!g66) & (g72) & (g73)) + ((!shiftx2x) & (!shiftx3x) & (!g65) & (g66) & (!g72) & (g73)) + ((!shiftx2x) & (!shiftx3x) & (!g65) & (g66) & (g72) & (g73)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (!g66) & (!g72) & (g73)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (!g66) & (g72) & (g73)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (g66) & (!g72) & (g73)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (g66) & (g72) & (g73)) + ((!shiftx2x) & (shiftx3x) & (g65) & (!g66) & (!g72) & (!g73)) + ((!shiftx2x) & (shiftx3x) & (g65) & (!g66) & (!g72) & (g73)) + ((!shiftx2x) & (shiftx3x) & (g65) & (!g66) & (g72) & (!g73)) + ((!shiftx2x) & (shiftx3x) & (g65) & (!g66) & (g72) & (g73)) + ((!shiftx2x) & (shiftx3x) & (g65) & (g66) & (!g72) & (!g73)) + ((!shiftx2x) & (shiftx3x) & (g65) & (g66) & (!g72) & (g73)) + ((!shiftx2x) & (shiftx3x) & (g65) & (g66) & (g72) & (!g73)) + ((!shiftx2x) & (shiftx3x) & (g65) & (g66) & (g72) & (g73)) + ((shiftx2x) & (!shiftx3x) & (!g65) & (!g66) & (g72) & (!g73)) + ((shiftx2x) & (!shiftx3x) & (!g65) & (!g66) & (g72) & (g73)) + ((shiftx2x) & (!shiftx3x) & (!g65) & (g66) & (g72) & (!g73)) + ((shiftx2x) & (!shiftx3x) & (!g65) & (g66) & (g72) & (g73)) + ((shiftx2x) & (!shiftx3x) & (g65) & (!g66) & (g72) & (!g73)) + ((shiftx2x) & (!shiftx3x) & (g65) & (!g66) & (g72) & (g73)) + ((shiftx2x) & (!shiftx3x) & (g65) & (g66) & (g72) & (!g73)) + ((shiftx2x) & (!shiftx3x) & (g65) & (g66) & (g72) & (g73)) + ((shiftx2x) & (shiftx3x) & (!g65) & (g66) & (!g72) & (!g73)) + ((shiftx2x) & (shiftx3x) & (!g65) & (g66) & (!g72) & (g73)) + ((shiftx2x) & (shiftx3x) & (!g65) & (g66) & (g72) & (!g73)) + ((shiftx2x) & (shiftx3x) & (!g65) & (g66) & (g72) & (g73)) + ((shiftx2x) & (shiftx3x) & (g65) & (g66) & (!g72) & (!g73)) + ((shiftx2x) & (shiftx3x) & (g65) & (g66) & (!g72) & (g73)) + ((shiftx2x) & (shiftx3x) & (g65) & (g66) & (g72) & (!g73)) + ((shiftx2x) & (shiftx3x) & (g65) & (g66) & (g72) & (g73)));
	assign g234 = (((!shiftx2x) & (!shiftx3x) & (!g70) & (!g71) & (!g82) & (g83)) + ((!shiftx2x) & (!shiftx3x) & (!g70) & (!g71) & (g82) & (g83)) + ((!shiftx2x) & (!shiftx3x) & (!g70) & (g71) & (!g82) & (g83)) + ((!shiftx2x) & (!shiftx3x) & (!g70) & (g71) & (g82) & (g83)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (!g71) & (!g82) & (g83)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (!g71) & (g82) & (g83)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (g71) & (!g82) & (g83)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (g71) & (g82) & (g83)) + ((!shiftx2x) & (shiftx3x) & (g70) & (!g71) & (!g82) & (!g83)) + ((!shiftx2x) & (shiftx3x) & (g70) & (!g71) & (!g82) & (g83)) + ((!shiftx2x) & (shiftx3x) & (g70) & (!g71) & (g82) & (!g83)) + ((!shiftx2x) & (shiftx3x) & (g70) & (!g71) & (g82) & (g83)) + ((!shiftx2x) & (shiftx3x) & (g70) & (g71) & (!g82) & (!g83)) + ((!shiftx2x) & (shiftx3x) & (g70) & (g71) & (!g82) & (g83)) + ((!shiftx2x) & (shiftx3x) & (g70) & (g71) & (g82) & (!g83)) + ((!shiftx2x) & (shiftx3x) & (g70) & (g71) & (g82) & (g83)) + ((shiftx2x) & (!shiftx3x) & (!g70) & (!g71) & (g82) & (!g83)) + ((shiftx2x) & (!shiftx3x) & (!g70) & (!g71) & (g82) & (g83)) + ((shiftx2x) & (!shiftx3x) & (!g70) & (g71) & (g82) & (!g83)) + ((shiftx2x) & (!shiftx3x) & (!g70) & (g71) & (g82) & (g83)) + ((shiftx2x) & (!shiftx3x) & (g70) & (!g71) & (g82) & (!g83)) + ((shiftx2x) & (!shiftx3x) & (g70) & (!g71) & (g82) & (g83)) + ((shiftx2x) & (!shiftx3x) & (g70) & (g71) & (g82) & (!g83)) + ((shiftx2x) & (!shiftx3x) & (g70) & (g71) & (g82) & (g83)) + ((shiftx2x) & (shiftx3x) & (!g70) & (g71) & (!g82) & (!g83)) + ((shiftx2x) & (shiftx3x) & (!g70) & (g71) & (!g82) & (g83)) + ((shiftx2x) & (shiftx3x) & (!g70) & (g71) & (g82) & (!g83)) + ((shiftx2x) & (shiftx3x) & (!g70) & (g71) & (g82) & (g83)) + ((shiftx2x) & (shiftx3x) & (g70) & (g71) & (!g82) & (!g83)) + ((shiftx2x) & (shiftx3x) & (g70) & (g71) & (!g82) & (g83)) + ((shiftx2x) & (shiftx3x) & (g70) & (g71) & (g82) & (!g83)) + ((shiftx2x) & (shiftx3x) & (g70) & (g71) & (g82) & (g83)));
	assign g235 = (((!shiftx2x) & (!shiftx3x) & (!g51) & (g52) & (!g75) & (!g76)) + ((!shiftx2x) & (!shiftx3x) & (!g51) & (g52) & (!g75) & (g76)) + ((!shiftx2x) & (!shiftx3x) & (!g51) & (g52) & (g75) & (!g76)) + ((!shiftx2x) & (!shiftx3x) & (!g51) & (g52) & (g75) & (g76)) + ((!shiftx2x) & (!shiftx3x) & (g51) & (g52) & (!g75) & (!g76)) + ((!shiftx2x) & (!shiftx3x) & (g51) & (g52) & (!g75) & (g76)) + ((!shiftx2x) & (!shiftx3x) & (g51) & (g52) & (g75) & (!g76)) + ((!shiftx2x) & (!shiftx3x) & (g51) & (g52) & (g75) & (g76)) + ((!shiftx2x) & (shiftx3x) & (!g51) & (!g52) & (g75) & (!g76)) + ((!shiftx2x) & (shiftx3x) & (!g51) & (!g52) & (g75) & (g76)) + ((!shiftx2x) & (shiftx3x) & (!g51) & (g52) & (g75) & (!g76)) + ((!shiftx2x) & (shiftx3x) & (!g51) & (g52) & (g75) & (g76)) + ((!shiftx2x) & (shiftx3x) & (g51) & (!g52) & (g75) & (!g76)) + ((!shiftx2x) & (shiftx3x) & (g51) & (!g52) & (g75) & (g76)) + ((!shiftx2x) & (shiftx3x) & (g51) & (g52) & (g75) & (!g76)) + ((!shiftx2x) & (shiftx3x) & (g51) & (g52) & (g75) & (g76)) + ((shiftx2x) & (!shiftx3x) & (g51) & (!g52) & (!g75) & (!g76)) + ((shiftx2x) & (!shiftx3x) & (g51) & (!g52) & (!g75) & (g76)) + ((shiftx2x) & (!shiftx3x) & (g51) & (!g52) & (g75) & (!g76)) + ((shiftx2x) & (!shiftx3x) & (g51) & (!g52) & (g75) & (g76)) + ((shiftx2x) & (!shiftx3x) & (g51) & (g52) & (!g75) & (!g76)) + ((shiftx2x) & (!shiftx3x) & (g51) & (g52) & (!g75) & (g76)) + ((shiftx2x) & (!shiftx3x) & (g51) & (g52) & (g75) & (!g76)) + ((shiftx2x) & (!shiftx3x) & (g51) & (g52) & (g75) & (g76)) + ((shiftx2x) & (shiftx3x) & (!g51) & (!g52) & (!g75) & (g76)) + ((shiftx2x) & (shiftx3x) & (!g51) & (!g52) & (g75) & (g76)) + ((shiftx2x) & (shiftx3x) & (!g51) & (g52) & (!g75) & (g76)) + ((shiftx2x) & (shiftx3x) & (!g51) & (g52) & (g75) & (g76)) + ((shiftx2x) & (shiftx3x) & (g51) & (!g52) & (!g75) & (g76)) + ((shiftx2x) & (shiftx3x) & (g51) & (!g52) & (g75) & (g76)) + ((shiftx2x) & (shiftx3x) & (g51) & (g52) & (!g75) & (g76)) + ((shiftx2x) & (shiftx3x) & (g51) & (g52) & (g75) & (g76)));
	assign g236 = (((!shiftx2x) & (!shiftx3x) & (!g77) & (g78) & (!g80) & (!g81)) + ((!shiftx2x) & (!shiftx3x) & (!g77) & (g78) & (!g80) & (g81)) + ((!shiftx2x) & (!shiftx3x) & (!g77) & (g78) & (g80) & (!g81)) + ((!shiftx2x) & (!shiftx3x) & (!g77) & (g78) & (g80) & (g81)) + ((!shiftx2x) & (!shiftx3x) & (g77) & (g78) & (!g80) & (!g81)) + ((!shiftx2x) & (!shiftx3x) & (g77) & (g78) & (!g80) & (g81)) + ((!shiftx2x) & (!shiftx3x) & (g77) & (g78) & (g80) & (!g81)) + ((!shiftx2x) & (!shiftx3x) & (g77) & (g78) & (g80) & (g81)) + ((!shiftx2x) & (shiftx3x) & (!g77) & (!g78) & (g80) & (!g81)) + ((!shiftx2x) & (shiftx3x) & (!g77) & (!g78) & (g80) & (g81)) + ((!shiftx2x) & (shiftx3x) & (!g77) & (g78) & (g80) & (!g81)) + ((!shiftx2x) & (shiftx3x) & (!g77) & (g78) & (g80) & (g81)) + ((!shiftx2x) & (shiftx3x) & (g77) & (!g78) & (g80) & (!g81)) + ((!shiftx2x) & (shiftx3x) & (g77) & (!g78) & (g80) & (g81)) + ((!shiftx2x) & (shiftx3x) & (g77) & (g78) & (g80) & (!g81)) + ((!shiftx2x) & (shiftx3x) & (g77) & (g78) & (g80) & (g81)) + ((shiftx2x) & (!shiftx3x) & (g77) & (!g78) & (!g80) & (!g81)) + ((shiftx2x) & (!shiftx3x) & (g77) & (!g78) & (!g80) & (g81)) + ((shiftx2x) & (!shiftx3x) & (g77) & (!g78) & (g80) & (!g81)) + ((shiftx2x) & (!shiftx3x) & (g77) & (!g78) & (g80) & (g81)) + ((shiftx2x) & (!shiftx3x) & (g77) & (g78) & (!g80) & (!g81)) + ((shiftx2x) & (!shiftx3x) & (g77) & (g78) & (!g80) & (g81)) + ((shiftx2x) & (!shiftx3x) & (g77) & (g78) & (g80) & (!g81)) + ((shiftx2x) & (!shiftx3x) & (g77) & (g78) & (g80) & (g81)) + ((shiftx2x) & (shiftx3x) & (!g77) & (!g78) & (!g80) & (g81)) + ((shiftx2x) & (shiftx3x) & (!g77) & (!g78) & (g80) & (g81)) + ((shiftx2x) & (shiftx3x) & (!g77) & (g78) & (!g80) & (g81)) + ((shiftx2x) & (shiftx3x) & (!g77) & (g78) & (g80) & (g81)) + ((shiftx2x) & (shiftx3x) & (g77) & (!g78) & (!g80) & (g81)) + ((shiftx2x) & (shiftx3x) & (g77) & (!g78) & (g80) & (g81)) + ((shiftx2x) & (shiftx3x) & (g77) & (g78) & (!g80) & (g81)) + ((shiftx2x) & (shiftx3x) & (g77) & (g78) & (g80) & (g81)));
	assign g237 = (((!shiftx4x) & (!shiftx5x) & (!g233) & (!g234) & (g235) & (!g236)) + ((!shiftx4x) & (!shiftx5x) & (!g233) & (!g234) & (g235) & (g236)) + ((!shiftx4x) & (!shiftx5x) & (!g233) & (g234) & (g235) & (!g236)) + ((!shiftx4x) & (!shiftx5x) & (!g233) & (g234) & (g235) & (g236)) + ((!shiftx4x) & (!shiftx5x) & (g233) & (!g234) & (g235) & (!g236)) + ((!shiftx4x) & (!shiftx5x) & (g233) & (!g234) & (g235) & (g236)) + ((!shiftx4x) & (!shiftx5x) & (g233) & (g234) & (g235) & (!g236)) + ((!shiftx4x) & (!shiftx5x) & (g233) & (g234) & (g235) & (g236)) + ((!shiftx4x) & (shiftx5x) & (!g233) & (g234) & (!g235) & (!g236)) + ((!shiftx4x) & (shiftx5x) & (!g233) & (g234) & (!g235) & (g236)) + ((!shiftx4x) & (shiftx5x) & (!g233) & (g234) & (g235) & (!g236)) + ((!shiftx4x) & (shiftx5x) & (!g233) & (g234) & (g235) & (g236)) + ((!shiftx4x) & (shiftx5x) & (g233) & (g234) & (!g235) & (!g236)) + ((!shiftx4x) & (shiftx5x) & (g233) & (g234) & (!g235) & (g236)) + ((!shiftx4x) & (shiftx5x) & (g233) & (g234) & (g235) & (!g236)) + ((!shiftx4x) & (shiftx5x) & (g233) & (g234) & (g235) & (g236)) + ((shiftx4x) & (!shiftx5x) & (!g233) & (!g234) & (!g235) & (g236)) + ((shiftx4x) & (!shiftx5x) & (!g233) & (!g234) & (g235) & (g236)) + ((shiftx4x) & (!shiftx5x) & (!g233) & (g234) & (!g235) & (g236)) + ((shiftx4x) & (!shiftx5x) & (!g233) & (g234) & (g235) & (g236)) + ((shiftx4x) & (!shiftx5x) & (g233) & (!g234) & (!g235) & (g236)) + ((shiftx4x) & (!shiftx5x) & (g233) & (!g234) & (g235) & (g236)) + ((shiftx4x) & (!shiftx5x) & (g233) & (g234) & (!g235) & (g236)) + ((shiftx4x) & (!shiftx5x) & (g233) & (g234) & (g235) & (g236)) + ((shiftx4x) & (shiftx5x) & (g233) & (!g234) & (!g235) & (!g236)) + ((shiftx4x) & (shiftx5x) & (g233) & (!g234) & (!g235) & (g236)) + ((shiftx4x) & (shiftx5x) & (g233) & (!g234) & (g235) & (!g236)) + ((shiftx4x) & (shiftx5x) & (g233) & (!g234) & (g235) & (g236)) + ((shiftx4x) & (shiftx5x) & (g233) & (g234) & (!g235) & (!g236)) + ((shiftx4x) & (shiftx5x) & (g233) & (g234) & (!g235) & (g236)) + ((shiftx4x) & (shiftx5x) & (g233) & (g234) & (g235) & (!g236)) + ((shiftx4x) & (shiftx5x) & (g233) & (g234) & (g235) & (g236)));
	assign resultx9x = (((!shiftx6x) & (sk[109]) & (!g232) & (g237)) + ((!shiftx6x) & (sk[109]) & (g232) & (g237)) + ((shiftx6x) & (!sk[109]) & (!g232) & (!g237)) + ((shiftx6x) & (!sk[109]) & (!g232) & (g237)) + ((shiftx6x) & (!sk[109]) & (g232) & (!g237)) + ((shiftx6x) & (!sk[109]) & (g232) & (g237)) + ((shiftx6x) & (sk[109]) & (g232) & (!g237)) + ((shiftx6x) & (sk[109]) & (g232) & (g237)));
	assign g239 = (((!shiftx2x) & (!shiftx3x) & (!g89) & (g90) & (!g97) & (!g98)) + ((!shiftx2x) & (!shiftx3x) & (!g89) & (g90) & (!g97) & (g98)) + ((!shiftx2x) & (!shiftx3x) & (!g89) & (g90) & (g97) & (!g98)) + ((!shiftx2x) & (!shiftx3x) & (!g89) & (g90) & (g97) & (g98)) + ((!shiftx2x) & (!shiftx3x) & (g89) & (g90) & (!g97) & (!g98)) + ((!shiftx2x) & (!shiftx3x) & (g89) & (g90) & (!g97) & (g98)) + ((!shiftx2x) & (!shiftx3x) & (g89) & (g90) & (g97) & (!g98)) + ((!shiftx2x) & (!shiftx3x) & (g89) & (g90) & (g97) & (g98)) + ((!shiftx2x) & (shiftx3x) & (!g89) & (!g90) & (g97) & (!g98)) + ((!shiftx2x) & (shiftx3x) & (!g89) & (!g90) & (g97) & (g98)) + ((!shiftx2x) & (shiftx3x) & (!g89) & (g90) & (g97) & (!g98)) + ((!shiftx2x) & (shiftx3x) & (!g89) & (g90) & (g97) & (g98)) + ((!shiftx2x) & (shiftx3x) & (g89) & (!g90) & (g97) & (!g98)) + ((!shiftx2x) & (shiftx3x) & (g89) & (!g90) & (g97) & (g98)) + ((!shiftx2x) & (shiftx3x) & (g89) & (g90) & (g97) & (!g98)) + ((!shiftx2x) & (shiftx3x) & (g89) & (g90) & (g97) & (g98)) + ((shiftx2x) & (!shiftx3x) & (g89) & (!g90) & (!g97) & (!g98)) + ((shiftx2x) & (!shiftx3x) & (g89) & (!g90) & (!g97) & (g98)) + ((shiftx2x) & (!shiftx3x) & (g89) & (!g90) & (g97) & (!g98)) + ((shiftx2x) & (!shiftx3x) & (g89) & (!g90) & (g97) & (g98)) + ((shiftx2x) & (!shiftx3x) & (g89) & (g90) & (!g97) & (!g98)) + ((shiftx2x) & (!shiftx3x) & (g89) & (g90) & (!g97) & (g98)) + ((shiftx2x) & (!shiftx3x) & (g89) & (g90) & (g97) & (!g98)) + ((shiftx2x) & (!shiftx3x) & (g89) & (g90) & (g97) & (g98)) + ((shiftx2x) & (shiftx3x) & (!g89) & (!g90) & (!g97) & (g98)) + ((shiftx2x) & (shiftx3x) & (!g89) & (!g90) & (g97) & (g98)) + ((shiftx2x) & (shiftx3x) & (!g89) & (g90) & (!g97) & (g98)) + ((shiftx2x) & (shiftx3x) & (!g89) & (g90) & (g97) & (g98)) + ((shiftx2x) & (shiftx3x) & (g89) & (!g90) & (!g97) & (g98)) + ((shiftx2x) & (shiftx3x) & (g89) & (!g90) & (g97) & (g98)) + ((shiftx2x) & (shiftx3x) & (g89) & (g90) & (!g97) & (g98)) + ((shiftx2x) & (shiftx3x) & (g89) & (g90) & (g97) & (g98)));
	assign g240 = (((!shiftx2x) & (!shiftx3x) & (!g87) & (!g88) & (!g110) & (g111)) + ((!shiftx2x) & (!shiftx3x) & (!g87) & (!g88) & (g110) & (g111)) + ((!shiftx2x) & (!shiftx3x) & (!g87) & (g88) & (!g110) & (g111)) + ((!shiftx2x) & (!shiftx3x) & (!g87) & (g88) & (g110) & (g111)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (!g88) & (!g110) & (g111)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (!g88) & (g110) & (g111)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (g88) & (!g110) & (g111)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (g88) & (g110) & (g111)) + ((!shiftx2x) & (shiftx3x) & (g87) & (!g88) & (!g110) & (!g111)) + ((!shiftx2x) & (shiftx3x) & (g87) & (!g88) & (!g110) & (g111)) + ((!shiftx2x) & (shiftx3x) & (g87) & (!g88) & (g110) & (!g111)) + ((!shiftx2x) & (shiftx3x) & (g87) & (!g88) & (g110) & (g111)) + ((!shiftx2x) & (shiftx3x) & (g87) & (g88) & (!g110) & (!g111)) + ((!shiftx2x) & (shiftx3x) & (g87) & (g88) & (!g110) & (g111)) + ((!shiftx2x) & (shiftx3x) & (g87) & (g88) & (g110) & (!g111)) + ((!shiftx2x) & (shiftx3x) & (g87) & (g88) & (g110) & (g111)) + ((shiftx2x) & (!shiftx3x) & (!g87) & (!g88) & (g110) & (!g111)) + ((shiftx2x) & (!shiftx3x) & (!g87) & (!g88) & (g110) & (g111)) + ((shiftx2x) & (!shiftx3x) & (!g87) & (g88) & (g110) & (!g111)) + ((shiftx2x) & (!shiftx3x) & (!g87) & (g88) & (g110) & (g111)) + ((shiftx2x) & (!shiftx3x) & (g87) & (!g88) & (g110) & (!g111)) + ((shiftx2x) & (!shiftx3x) & (g87) & (!g88) & (g110) & (g111)) + ((shiftx2x) & (!shiftx3x) & (g87) & (g88) & (g110) & (!g111)) + ((shiftx2x) & (!shiftx3x) & (g87) & (g88) & (g110) & (g111)) + ((shiftx2x) & (shiftx3x) & (!g87) & (g88) & (!g110) & (!g111)) + ((shiftx2x) & (shiftx3x) & (!g87) & (g88) & (!g110) & (g111)) + ((shiftx2x) & (shiftx3x) & (!g87) & (g88) & (g110) & (!g111)) + ((shiftx2x) & (shiftx3x) & (!g87) & (g88) & (g110) & (g111)) + ((shiftx2x) & (shiftx3x) & (g87) & (g88) & (!g110) & (!g111)) + ((shiftx2x) & (shiftx3x) & (g87) & (g88) & (!g110) & (g111)) + ((shiftx2x) & (shiftx3x) & (g87) & (g88) & (g110) & (!g111)) + ((shiftx2x) & (shiftx3x) & (g87) & (g88) & (g110) & (g111)));
	assign g241 = (((!shiftx2x) & (!shiftx3x) & (!g99) & (g100) & (!g102) & (!g103)) + ((!shiftx2x) & (!shiftx3x) & (!g99) & (g100) & (!g102) & (g103)) + ((!shiftx2x) & (!shiftx3x) & (!g99) & (g100) & (g102) & (!g103)) + ((!shiftx2x) & (!shiftx3x) & (!g99) & (g100) & (g102) & (g103)) + ((!shiftx2x) & (!shiftx3x) & (g99) & (g100) & (!g102) & (!g103)) + ((!shiftx2x) & (!shiftx3x) & (g99) & (g100) & (!g102) & (g103)) + ((!shiftx2x) & (!shiftx3x) & (g99) & (g100) & (g102) & (!g103)) + ((!shiftx2x) & (!shiftx3x) & (g99) & (g100) & (g102) & (g103)) + ((!shiftx2x) & (shiftx3x) & (!g99) & (!g100) & (g102) & (!g103)) + ((!shiftx2x) & (shiftx3x) & (!g99) & (!g100) & (g102) & (g103)) + ((!shiftx2x) & (shiftx3x) & (!g99) & (g100) & (g102) & (!g103)) + ((!shiftx2x) & (shiftx3x) & (!g99) & (g100) & (g102) & (g103)) + ((!shiftx2x) & (shiftx3x) & (g99) & (!g100) & (g102) & (!g103)) + ((!shiftx2x) & (shiftx3x) & (g99) & (!g100) & (g102) & (g103)) + ((!shiftx2x) & (shiftx3x) & (g99) & (g100) & (g102) & (!g103)) + ((!shiftx2x) & (shiftx3x) & (g99) & (g100) & (g102) & (g103)) + ((shiftx2x) & (!shiftx3x) & (g99) & (!g100) & (!g102) & (!g103)) + ((shiftx2x) & (!shiftx3x) & (g99) & (!g100) & (!g102) & (g103)) + ((shiftx2x) & (!shiftx3x) & (g99) & (!g100) & (g102) & (!g103)) + ((shiftx2x) & (!shiftx3x) & (g99) & (!g100) & (g102) & (g103)) + ((shiftx2x) & (!shiftx3x) & (g99) & (g100) & (!g102) & (!g103)) + ((shiftx2x) & (!shiftx3x) & (g99) & (g100) & (!g102) & (g103)) + ((shiftx2x) & (!shiftx3x) & (g99) & (g100) & (g102) & (!g103)) + ((shiftx2x) & (!shiftx3x) & (g99) & (g100) & (g102) & (g103)) + ((shiftx2x) & (shiftx3x) & (!g99) & (!g100) & (!g102) & (g103)) + ((shiftx2x) & (shiftx3x) & (!g99) & (!g100) & (g102) & (g103)) + ((shiftx2x) & (shiftx3x) & (!g99) & (g100) & (!g102) & (g103)) + ((shiftx2x) & (shiftx3x) & (!g99) & (g100) & (g102) & (g103)) + ((shiftx2x) & (shiftx3x) & (g99) & (!g100) & (!g102) & (g103)) + ((shiftx2x) & (shiftx3x) & (g99) & (!g100) & (g102) & (g103)) + ((shiftx2x) & (shiftx3x) & (g99) & (g100) & (!g102) & (g103)) + ((shiftx2x) & (shiftx3x) & (g99) & (g100) & (g102) & (g103)));
	assign g242 = (((!shiftx2x) & (!shiftx3x) & (!g92) & (!g93) & (!g104) & (g105)) + ((!shiftx2x) & (!shiftx3x) & (!g92) & (!g93) & (g104) & (g105)) + ((!shiftx2x) & (!shiftx3x) & (!g92) & (g93) & (!g104) & (g105)) + ((!shiftx2x) & (!shiftx3x) & (!g92) & (g93) & (g104) & (g105)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (!g93) & (!g104) & (g105)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (!g93) & (g104) & (g105)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (g93) & (!g104) & (g105)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (g93) & (g104) & (g105)) + ((!shiftx2x) & (shiftx3x) & (g92) & (!g93) & (!g104) & (!g105)) + ((!shiftx2x) & (shiftx3x) & (g92) & (!g93) & (!g104) & (g105)) + ((!shiftx2x) & (shiftx3x) & (g92) & (!g93) & (g104) & (!g105)) + ((!shiftx2x) & (shiftx3x) & (g92) & (!g93) & (g104) & (g105)) + ((!shiftx2x) & (shiftx3x) & (g92) & (g93) & (!g104) & (!g105)) + ((!shiftx2x) & (shiftx3x) & (g92) & (g93) & (!g104) & (g105)) + ((!shiftx2x) & (shiftx3x) & (g92) & (g93) & (g104) & (!g105)) + ((!shiftx2x) & (shiftx3x) & (g92) & (g93) & (g104) & (g105)) + ((shiftx2x) & (!shiftx3x) & (!g92) & (!g93) & (g104) & (!g105)) + ((shiftx2x) & (!shiftx3x) & (!g92) & (!g93) & (g104) & (g105)) + ((shiftx2x) & (!shiftx3x) & (!g92) & (g93) & (g104) & (!g105)) + ((shiftx2x) & (!shiftx3x) & (!g92) & (g93) & (g104) & (g105)) + ((shiftx2x) & (!shiftx3x) & (g92) & (!g93) & (g104) & (!g105)) + ((shiftx2x) & (!shiftx3x) & (g92) & (!g93) & (g104) & (g105)) + ((shiftx2x) & (!shiftx3x) & (g92) & (g93) & (g104) & (!g105)) + ((shiftx2x) & (!shiftx3x) & (g92) & (g93) & (g104) & (g105)) + ((shiftx2x) & (shiftx3x) & (!g92) & (g93) & (!g104) & (!g105)) + ((shiftx2x) & (shiftx3x) & (!g92) & (g93) & (!g104) & (g105)) + ((shiftx2x) & (shiftx3x) & (!g92) & (g93) & (g104) & (!g105)) + ((shiftx2x) & (shiftx3x) & (!g92) & (g93) & (g104) & (g105)) + ((shiftx2x) & (shiftx3x) & (g92) & (g93) & (!g104) & (!g105)) + ((shiftx2x) & (shiftx3x) & (g92) & (g93) & (!g104) & (g105)) + ((shiftx2x) & (shiftx3x) & (g92) & (g93) & (g104) & (!g105)) + ((shiftx2x) & (shiftx3x) & (g92) & (g93) & (g104) & (g105)));
	assign g243 = (((!shiftx4x) & (!shiftx5x) & (!g239) & (g240) & (!g241) & (!g242)) + ((!shiftx4x) & (!shiftx5x) & (!g239) & (g240) & (!g241) & (g242)) + ((!shiftx4x) & (!shiftx5x) & (!g239) & (g240) & (g241) & (!g242)) + ((!shiftx4x) & (!shiftx5x) & (!g239) & (g240) & (g241) & (g242)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (g240) & (!g241) & (!g242)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (g240) & (!g241) & (g242)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (g240) & (g241) & (!g242)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (g240) & (g241) & (g242)) + ((!shiftx4x) & (shiftx5x) & (!g239) & (!g240) & (g241) & (!g242)) + ((!shiftx4x) & (shiftx5x) & (!g239) & (!g240) & (g241) & (g242)) + ((!shiftx4x) & (shiftx5x) & (!g239) & (g240) & (g241) & (!g242)) + ((!shiftx4x) & (shiftx5x) & (!g239) & (g240) & (g241) & (g242)) + ((!shiftx4x) & (shiftx5x) & (g239) & (!g240) & (g241) & (!g242)) + ((!shiftx4x) & (shiftx5x) & (g239) & (!g240) & (g241) & (g242)) + ((!shiftx4x) & (shiftx5x) & (g239) & (g240) & (g241) & (!g242)) + ((!shiftx4x) & (shiftx5x) & (g239) & (g240) & (g241) & (g242)) + ((shiftx4x) & (!shiftx5x) & (g239) & (!g240) & (!g241) & (!g242)) + ((shiftx4x) & (!shiftx5x) & (g239) & (!g240) & (!g241) & (g242)) + ((shiftx4x) & (!shiftx5x) & (g239) & (!g240) & (g241) & (!g242)) + ((shiftx4x) & (!shiftx5x) & (g239) & (!g240) & (g241) & (g242)) + ((shiftx4x) & (!shiftx5x) & (g239) & (g240) & (!g241) & (!g242)) + ((shiftx4x) & (!shiftx5x) & (g239) & (g240) & (!g241) & (g242)) + ((shiftx4x) & (!shiftx5x) & (g239) & (g240) & (g241) & (!g242)) + ((shiftx4x) & (!shiftx5x) & (g239) & (g240) & (g241) & (g242)) + ((shiftx4x) & (shiftx5x) & (!g239) & (!g240) & (!g241) & (g242)) + ((shiftx4x) & (shiftx5x) & (!g239) & (!g240) & (g241) & (g242)) + ((shiftx4x) & (shiftx5x) & (!g239) & (g240) & (!g241) & (g242)) + ((shiftx4x) & (shiftx5x) & (!g239) & (g240) & (g241) & (g242)) + ((shiftx4x) & (shiftx5x) & (g239) & (!g240) & (!g241) & (g242)) + ((shiftx4x) & (shiftx5x) & (g239) & (!g240) & (g241) & (g242)) + ((shiftx4x) & (shiftx5x) & (g239) & (g240) & (!g241) & (g242)) + ((shiftx4x) & (shiftx5x) & (g239) & (g240) & (g241) & (g242)));
	assign g244 = (((!shiftx2x) & (!shiftx3x) & (!g108) & (!g109) & (!g115) & (g116)) + ((!shiftx2x) & (!shiftx3x) & (!g108) & (!g109) & (g115) & (g116)) + ((!shiftx2x) & (!shiftx3x) & (!g108) & (g109) & (!g115) & (g116)) + ((!shiftx2x) & (!shiftx3x) & (!g108) & (g109) & (g115) & (g116)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (!g109) & (!g115) & (g116)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (!g109) & (g115) & (g116)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (g109) & (!g115) & (g116)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (g109) & (g115) & (g116)) + ((!shiftx2x) & (shiftx3x) & (g108) & (!g109) & (!g115) & (!g116)) + ((!shiftx2x) & (shiftx3x) & (g108) & (!g109) & (!g115) & (g116)) + ((!shiftx2x) & (shiftx3x) & (g108) & (!g109) & (g115) & (!g116)) + ((!shiftx2x) & (shiftx3x) & (g108) & (!g109) & (g115) & (g116)) + ((!shiftx2x) & (shiftx3x) & (g108) & (g109) & (!g115) & (!g116)) + ((!shiftx2x) & (shiftx3x) & (g108) & (g109) & (!g115) & (g116)) + ((!shiftx2x) & (shiftx3x) & (g108) & (g109) & (g115) & (!g116)) + ((!shiftx2x) & (shiftx3x) & (g108) & (g109) & (g115) & (g116)) + ((shiftx2x) & (!shiftx3x) & (!g108) & (!g109) & (g115) & (!g116)) + ((shiftx2x) & (!shiftx3x) & (!g108) & (!g109) & (g115) & (g116)) + ((shiftx2x) & (!shiftx3x) & (!g108) & (g109) & (g115) & (!g116)) + ((shiftx2x) & (!shiftx3x) & (!g108) & (g109) & (g115) & (g116)) + ((shiftx2x) & (!shiftx3x) & (g108) & (!g109) & (g115) & (!g116)) + ((shiftx2x) & (!shiftx3x) & (g108) & (!g109) & (g115) & (g116)) + ((shiftx2x) & (!shiftx3x) & (g108) & (g109) & (g115) & (!g116)) + ((shiftx2x) & (!shiftx3x) & (g108) & (g109) & (g115) & (g116)) + ((shiftx2x) & (shiftx3x) & (!g108) & (g109) & (!g115) & (!g116)) + ((shiftx2x) & (shiftx3x) & (!g108) & (g109) & (!g115) & (g116)) + ((shiftx2x) & (shiftx3x) & (!g108) & (g109) & (g115) & (!g116)) + ((shiftx2x) & (shiftx3x) & (!g108) & (g109) & (g115) & (g116)) + ((shiftx2x) & (shiftx3x) & (g108) & (g109) & (!g115) & (!g116)) + ((shiftx2x) & (shiftx3x) & (g108) & (g109) & (!g115) & (g116)) + ((shiftx2x) & (shiftx3x) & (g108) & (g109) & (g115) & (!g116)) + ((shiftx2x) & (shiftx3x) & (g108) & (g109) & (g115) & (g116)));
	assign g245 = (((!shiftx2x) & (!shiftx3x) & (!g113) & (!g114) & (!g125) & (g126)) + ((!shiftx2x) & (!shiftx3x) & (!g113) & (!g114) & (g125) & (g126)) + ((!shiftx2x) & (!shiftx3x) & (!g113) & (g114) & (!g125) & (g126)) + ((!shiftx2x) & (!shiftx3x) & (!g113) & (g114) & (g125) & (g126)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (!g114) & (!g125) & (g126)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (!g114) & (g125) & (g126)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (g114) & (!g125) & (g126)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (g114) & (g125) & (g126)) + ((!shiftx2x) & (shiftx3x) & (g113) & (!g114) & (!g125) & (!g126)) + ((!shiftx2x) & (shiftx3x) & (g113) & (!g114) & (!g125) & (g126)) + ((!shiftx2x) & (shiftx3x) & (g113) & (!g114) & (g125) & (!g126)) + ((!shiftx2x) & (shiftx3x) & (g113) & (!g114) & (g125) & (g126)) + ((!shiftx2x) & (shiftx3x) & (g113) & (g114) & (!g125) & (!g126)) + ((!shiftx2x) & (shiftx3x) & (g113) & (g114) & (!g125) & (g126)) + ((!shiftx2x) & (shiftx3x) & (g113) & (g114) & (g125) & (!g126)) + ((!shiftx2x) & (shiftx3x) & (g113) & (g114) & (g125) & (g126)) + ((shiftx2x) & (!shiftx3x) & (!g113) & (!g114) & (g125) & (!g126)) + ((shiftx2x) & (!shiftx3x) & (!g113) & (!g114) & (g125) & (g126)) + ((shiftx2x) & (!shiftx3x) & (!g113) & (g114) & (g125) & (!g126)) + ((shiftx2x) & (!shiftx3x) & (!g113) & (g114) & (g125) & (g126)) + ((shiftx2x) & (!shiftx3x) & (g113) & (!g114) & (g125) & (!g126)) + ((shiftx2x) & (!shiftx3x) & (g113) & (!g114) & (g125) & (g126)) + ((shiftx2x) & (!shiftx3x) & (g113) & (g114) & (g125) & (!g126)) + ((shiftx2x) & (!shiftx3x) & (g113) & (g114) & (g125) & (g126)) + ((shiftx2x) & (shiftx3x) & (!g113) & (g114) & (!g125) & (!g126)) + ((shiftx2x) & (shiftx3x) & (!g113) & (g114) & (!g125) & (g126)) + ((shiftx2x) & (shiftx3x) & (!g113) & (g114) & (g125) & (!g126)) + ((shiftx2x) & (shiftx3x) & (!g113) & (g114) & (g125) & (g126)) + ((shiftx2x) & (shiftx3x) & (g113) & (g114) & (!g125) & (!g126)) + ((shiftx2x) & (shiftx3x) & (g113) & (g114) & (!g125) & (g126)) + ((shiftx2x) & (shiftx3x) & (g113) & (g114) & (g125) & (!g126)) + ((shiftx2x) & (shiftx3x) & (g113) & (g114) & (g125) & (g126)));
	assign g246 = (((!shiftx2x) & (!shiftx3x) & (!g94) & (g95) & (!g118) & (!g119)) + ((!shiftx2x) & (!shiftx3x) & (!g94) & (g95) & (!g118) & (g119)) + ((!shiftx2x) & (!shiftx3x) & (!g94) & (g95) & (g118) & (!g119)) + ((!shiftx2x) & (!shiftx3x) & (!g94) & (g95) & (g118) & (g119)) + ((!shiftx2x) & (!shiftx3x) & (g94) & (g95) & (!g118) & (!g119)) + ((!shiftx2x) & (!shiftx3x) & (g94) & (g95) & (!g118) & (g119)) + ((!shiftx2x) & (!shiftx3x) & (g94) & (g95) & (g118) & (!g119)) + ((!shiftx2x) & (!shiftx3x) & (g94) & (g95) & (g118) & (g119)) + ((!shiftx2x) & (shiftx3x) & (!g94) & (!g95) & (g118) & (!g119)) + ((!shiftx2x) & (shiftx3x) & (!g94) & (!g95) & (g118) & (g119)) + ((!shiftx2x) & (shiftx3x) & (!g94) & (g95) & (g118) & (!g119)) + ((!shiftx2x) & (shiftx3x) & (!g94) & (g95) & (g118) & (g119)) + ((!shiftx2x) & (shiftx3x) & (g94) & (!g95) & (g118) & (!g119)) + ((!shiftx2x) & (shiftx3x) & (g94) & (!g95) & (g118) & (g119)) + ((!shiftx2x) & (shiftx3x) & (g94) & (g95) & (g118) & (!g119)) + ((!shiftx2x) & (shiftx3x) & (g94) & (g95) & (g118) & (g119)) + ((shiftx2x) & (!shiftx3x) & (g94) & (!g95) & (!g118) & (!g119)) + ((shiftx2x) & (!shiftx3x) & (g94) & (!g95) & (!g118) & (g119)) + ((shiftx2x) & (!shiftx3x) & (g94) & (!g95) & (g118) & (!g119)) + ((shiftx2x) & (!shiftx3x) & (g94) & (!g95) & (g118) & (g119)) + ((shiftx2x) & (!shiftx3x) & (g94) & (g95) & (!g118) & (!g119)) + ((shiftx2x) & (!shiftx3x) & (g94) & (g95) & (!g118) & (g119)) + ((shiftx2x) & (!shiftx3x) & (g94) & (g95) & (g118) & (!g119)) + ((shiftx2x) & (!shiftx3x) & (g94) & (g95) & (g118) & (g119)) + ((shiftx2x) & (shiftx3x) & (!g94) & (!g95) & (!g118) & (g119)) + ((shiftx2x) & (shiftx3x) & (!g94) & (!g95) & (g118) & (g119)) + ((shiftx2x) & (shiftx3x) & (!g94) & (g95) & (!g118) & (g119)) + ((shiftx2x) & (shiftx3x) & (!g94) & (g95) & (g118) & (g119)) + ((shiftx2x) & (shiftx3x) & (g94) & (!g95) & (!g118) & (g119)) + ((shiftx2x) & (shiftx3x) & (g94) & (!g95) & (g118) & (g119)) + ((shiftx2x) & (shiftx3x) & (g94) & (g95) & (!g118) & (g119)) + ((shiftx2x) & (shiftx3x) & (g94) & (g95) & (g118) & (g119)));
	assign g247 = (((!shiftx2x) & (!shiftx3x) & (!g120) & (g121) & (!g123) & (!g124)) + ((!shiftx2x) & (!shiftx3x) & (!g120) & (g121) & (!g123) & (g124)) + ((!shiftx2x) & (!shiftx3x) & (!g120) & (g121) & (g123) & (!g124)) + ((!shiftx2x) & (!shiftx3x) & (!g120) & (g121) & (g123) & (g124)) + ((!shiftx2x) & (!shiftx3x) & (g120) & (g121) & (!g123) & (!g124)) + ((!shiftx2x) & (!shiftx3x) & (g120) & (g121) & (!g123) & (g124)) + ((!shiftx2x) & (!shiftx3x) & (g120) & (g121) & (g123) & (!g124)) + ((!shiftx2x) & (!shiftx3x) & (g120) & (g121) & (g123) & (g124)) + ((!shiftx2x) & (shiftx3x) & (!g120) & (!g121) & (g123) & (!g124)) + ((!shiftx2x) & (shiftx3x) & (!g120) & (!g121) & (g123) & (g124)) + ((!shiftx2x) & (shiftx3x) & (!g120) & (g121) & (g123) & (!g124)) + ((!shiftx2x) & (shiftx3x) & (!g120) & (g121) & (g123) & (g124)) + ((!shiftx2x) & (shiftx3x) & (g120) & (!g121) & (g123) & (!g124)) + ((!shiftx2x) & (shiftx3x) & (g120) & (!g121) & (g123) & (g124)) + ((!shiftx2x) & (shiftx3x) & (g120) & (g121) & (g123) & (!g124)) + ((!shiftx2x) & (shiftx3x) & (g120) & (g121) & (g123) & (g124)) + ((shiftx2x) & (!shiftx3x) & (g120) & (!g121) & (!g123) & (!g124)) + ((shiftx2x) & (!shiftx3x) & (g120) & (!g121) & (!g123) & (g124)) + ((shiftx2x) & (!shiftx3x) & (g120) & (!g121) & (g123) & (!g124)) + ((shiftx2x) & (!shiftx3x) & (g120) & (!g121) & (g123) & (g124)) + ((shiftx2x) & (!shiftx3x) & (g120) & (g121) & (!g123) & (!g124)) + ((shiftx2x) & (!shiftx3x) & (g120) & (g121) & (!g123) & (g124)) + ((shiftx2x) & (!shiftx3x) & (g120) & (g121) & (g123) & (!g124)) + ((shiftx2x) & (!shiftx3x) & (g120) & (g121) & (g123) & (g124)) + ((shiftx2x) & (shiftx3x) & (!g120) & (!g121) & (!g123) & (g124)) + ((shiftx2x) & (shiftx3x) & (!g120) & (!g121) & (g123) & (g124)) + ((shiftx2x) & (shiftx3x) & (!g120) & (g121) & (!g123) & (g124)) + ((shiftx2x) & (shiftx3x) & (!g120) & (g121) & (g123) & (g124)) + ((shiftx2x) & (shiftx3x) & (g120) & (!g121) & (!g123) & (g124)) + ((shiftx2x) & (shiftx3x) & (g120) & (!g121) & (g123) & (g124)) + ((shiftx2x) & (shiftx3x) & (g120) & (g121) & (!g123) & (g124)) + ((shiftx2x) & (shiftx3x) & (g120) & (g121) & (g123) & (g124)));
	assign g248 = (((!shiftx4x) & (!shiftx5x) & (!g244) & (!g245) & (g246) & (!g247)) + ((!shiftx4x) & (!shiftx5x) & (!g244) & (!g245) & (g246) & (g247)) + ((!shiftx4x) & (!shiftx5x) & (!g244) & (g245) & (g246) & (!g247)) + ((!shiftx4x) & (!shiftx5x) & (!g244) & (g245) & (g246) & (g247)) + ((!shiftx4x) & (!shiftx5x) & (g244) & (!g245) & (g246) & (!g247)) + ((!shiftx4x) & (!shiftx5x) & (g244) & (!g245) & (g246) & (g247)) + ((!shiftx4x) & (!shiftx5x) & (g244) & (g245) & (g246) & (!g247)) + ((!shiftx4x) & (!shiftx5x) & (g244) & (g245) & (g246) & (g247)) + ((!shiftx4x) & (shiftx5x) & (!g244) & (g245) & (!g246) & (!g247)) + ((!shiftx4x) & (shiftx5x) & (!g244) & (g245) & (!g246) & (g247)) + ((!shiftx4x) & (shiftx5x) & (!g244) & (g245) & (g246) & (!g247)) + ((!shiftx4x) & (shiftx5x) & (!g244) & (g245) & (g246) & (g247)) + ((!shiftx4x) & (shiftx5x) & (g244) & (g245) & (!g246) & (!g247)) + ((!shiftx4x) & (shiftx5x) & (g244) & (g245) & (!g246) & (g247)) + ((!shiftx4x) & (shiftx5x) & (g244) & (g245) & (g246) & (!g247)) + ((!shiftx4x) & (shiftx5x) & (g244) & (g245) & (g246) & (g247)) + ((shiftx4x) & (!shiftx5x) & (!g244) & (!g245) & (!g246) & (g247)) + ((shiftx4x) & (!shiftx5x) & (!g244) & (!g245) & (g246) & (g247)) + ((shiftx4x) & (!shiftx5x) & (!g244) & (g245) & (!g246) & (g247)) + ((shiftx4x) & (!shiftx5x) & (!g244) & (g245) & (g246) & (g247)) + ((shiftx4x) & (!shiftx5x) & (g244) & (!g245) & (!g246) & (g247)) + ((shiftx4x) & (!shiftx5x) & (g244) & (!g245) & (g246) & (g247)) + ((shiftx4x) & (!shiftx5x) & (g244) & (g245) & (!g246) & (g247)) + ((shiftx4x) & (!shiftx5x) & (g244) & (g245) & (g246) & (g247)) + ((shiftx4x) & (shiftx5x) & (g244) & (!g245) & (!g246) & (!g247)) + ((shiftx4x) & (shiftx5x) & (g244) & (!g245) & (!g246) & (g247)) + ((shiftx4x) & (shiftx5x) & (g244) & (!g245) & (g246) & (!g247)) + ((shiftx4x) & (shiftx5x) & (g244) & (!g245) & (g246) & (g247)) + ((shiftx4x) & (shiftx5x) & (g244) & (g245) & (!g246) & (!g247)) + ((shiftx4x) & (shiftx5x) & (g244) & (g245) & (!g246) & (g247)) + ((shiftx4x) & (shiftx5x) & (g244) & (g245) & (g246) & (!g247)) + ((shiftx4x) & (shiftx5x) & (g244) & (g245) & (g246) & (g247)));
	assign resultx10x = (((!sk[120]) & (shiftx6x) & (!g243) & (!g248)) + ((!sk[120]) & (shiftx6x) & (!g243) & (g248)) + ((!sk[120]) & (shiftx6x) & (g243) & (!g248)) + ((!sk[120]) & (shiftx6x) & (g243) & (g248)) + ((sk[120]) & (!shiftx6x) & (!g243) & (g248)) + ((sk[120]) & (!shiftx6x) & (g243) & (g248)) + ((sk[120]) & (shiftx6x) & (g243) & (!g248)) + ((sk[120]) & (shiftx6x) & (g243) & (g248)));
	assign g250 = (((!shiftx2x) & (!shiftx3x) & (!g132) & (g133) & (!g135) & (!g136)) + ((!shiftx2x) & (!shiftx3x) & (!g132) & (g133) & (!g135) & (g136)) + ((!shiftx2x) & (!shiftx3x) & (!g132) & (g133) & (g135) & (!g136)) + ((!shiftx2x) & (!shiftx3x) & (!g132) & (g133) & (g135) & (g136)) + ((!shiftx2x) & (!shiftx3x) & (g132) & (g133) & (!g135) & (!g136)) + ((!shiftx2x) & (!shiftx3x) & (g132) & (g133) & (!g135) & (g136)) + ((!shiftx2x) & (!shiftx3x) & (g132) & (g133) & (g135) & (!g136)) + ((!shiftx2x) & (!shiftx3x) & (g132) & (g133) & (g135) & (g136)) + ((!shiftx2x) & (shiftx3x) & (!g132) & (!g133) & (g135) & (!g136)) + ((!shiftx2x) & (shiftx3x) & (!g132) & (!g133) & (g135) & (g136)) + ((!shiftx2x) & (shiftx3x) & (!g132) & (g133) & (g135) & (!g136)) + ((!shiftx2x) & (shiftx3x) & (!g132) & (g133) & (g135) & (g136)) + ((!shiftx2x) & (shiftx3x) & (g132) & (!g133) & (g135) & (!g136)) + ((!shiftx2x) & (shiftx3x) & (g132) & (!g133) & (g135) & (g136)) + ((!shiftx2x) & (shiftx3x) & (g132) & (g133) & (g135) & (!g136)) + ((!shiftx2x) & (shiftx3x) & (g132) & (g133) & (g135) & (g136)) + ((shiftx2x) & (!shiftx3x) & (g132) & (!g133) & (!g135) & (!g136)) + ((shiftx2x) & (!shiftx3x) & (g132) & (!g133) & (!g135) & (g136)) + ((shiftx2x) & (!shiftx3x) & (g132) & (!g133) & (g135) & (!g136)) + ((shiftx2x) & (!shiftx3x) & (g132) & (!g133) & (g135) & (g136)) + ((shiftx2x) & (!shiftx3x) & (g132) & (g133) & (!g135) & (!g136)) + ((shiftx2x) & (!shiftx3x) & (g132) & (g133) & (!g135) & (g136)) + ((shiftx2x) & (!shiftx3x) & (g132) & (g133) & (g135) & (!g136)) + ((shiftx2x) & (!shiftx3x) & (g132) & (g133) & (g135) & (g136)) + ((shiftx2x) & (shiftx3x) & (!g132) & (!g133) & (!g135) & (g136)) + ((shiftx2x) & (shiftx3x) & (!g132) & (!g133) & (g135) & (g136)) + ((shiftx2x) & (shiftx3x) & (!g132) & (g133) & (!g135) & (g136)) + ((shiftx2x) & (shiftx3x) & (!g132) & (g133) & (g135) & (g136)) + ((shiftx2x) & (shiftx3x) & (g132) & (!g133) & (!g135) & (g136)) + ((shiftx2x) & (shiftx3x) & (g132) & (!g133) & (g135) & (g136)) + ((shiftx2x) & (shiftx3x) & (g132) & (g133) & (!g135) & (g136)) + ((shiftx2x) & (shiftx3x) & (g132) & (g133) & (g135) & (g136)));
	assign g251 = (((!shiftx2x) & (!shiftx3x) & (!g130) & (!g131) & (!g168) & (g169)) + ((!shiftx2x) & (!shiftx3x) & (!g130) & (!g131) & (g168) & (g169)) + ((!shiftx2x) & (!shiftx3x) & (!g130) & (g131) & (!g168) & (g169)) + ((!shiftx2x) & (!shiftx3x) & (!g130) & (g131) & (g168) & (g169)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (!g131) & (!g168) & (g169)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (!g131) & (g168) & (g169)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (g131) & (!g168) & (g169)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (g131) & (g168) & (g169)) + ((!shiftx2x) & (shiftx3x) & (g130) & (!g131) & (!g168) & (!g169)) + ((!shiftx2x) & (shiftx3x) & (g130) & (!g131) & (!g168) & (g169)) + ((!shiftx2x) & (shiftx3x) & (g130) & (!g131) & (g168) & (!g169)) + ((!shiftx2x) & (shiftx3x) & (g130) & (!g131) & (g168) & (g169)) + ((!shiftx2x) & (shiftx3x) & (g130) & (g131) & (!g168) & (!g169)) + ((!shiftx2x) & (shiftx3x) & (g130) & (g131) & (!g168) & (g169)) + ((!shiftx2x) & (shiftx3x) & (g130) & (g131) & (g168) & (!g169)) + ((!shiftx2x) & (shiftx3x) & (g130) & (g131) & (g168) & (g169)) + ((shiftx2x) & (!shiftx3x) & (!g130) & (!g131) & (g168) & (!g169)) + ((shiftx2x) & (!shiftx3x) & (!g130) & (!g131) & (g168) & (g169)) + ((shiftx2x) & (!shiftx3x) & (!g130) & (g131) & (g168) & (!g169)) + ((shiftx2x) & (!shiftx3x) & (!g130) & (g131) & (g168) & (g169)) + ((shiftx2x) & (!shiftx3x) & (g130) & (!g131) & (g168) & (!g169)) + ((shiftx2x) & (!shiftx3x) & (g130) & (!g131) & (g168) & (g169)) + ((shiftx2x) & (!shiftx3x) & (g130) & (g131) & (g168) & (!g169)) + ((shiftx2x) & (!shiftx3x) & (g130) & (g131) & (g168) & (g169)) + ((shiftx2x) & (shiftx3x) & (!g130) & (g131) & (!g168) & (!g169)) + ((shiftx2x) & (shiftx3x) & (!g130) & (g131) & (!g168) & (g169)) + ((shiftx2x) & (shiftx3x) & (!g130) & (g131) & (g168) & (!g169)) + ((shiftx2x) & (shiftx3x) & (!g130) & (g131) & (g168) & (g169)) + ((shiftx2x) & (shiftx3x) & (g130) & (g131) & (!g168) & (!g169)) + ((shiftx2x) & (shiftx3x) & (g130) & (g131) & (!g168) & (g169)) + ((shiftx2x) & (shiftx3x) & (g130) & (g131) & (g168) & (!g169)) + ((shiftx2x) & (shiftx3x) & (g130) & (g131) & (g168) & (g169)));
	assign g252 = (((!shiftx2x) & (!shiftx3x) & (!g137) & (g138) & (!g145) & (!g146)) + ((!shiftx2x) & (!shiftx3x) & (!g137) & (g138) & (!g145) & (g146)) + ((!shiftx2x) & (!shiftx3x) & (!g137) & (g138) & (g145) & (!g146)) + ((!shiftx2x) & (!shiftx3x) & (!g137) & (g138) & (g145) & (g146)) + ((!shiftx2x) & (!shiftx3x) & (g137) & (g138) & (!g145) & (!g146)) + ((!shiftx2x) & (!shiftx3x) & (g137) & (g138) & (!g145) & (g146)) + ((!shiftx2x) & (!shiftx3x) & (g137) & (g138) & (g145) & (!g146)) + ((!shiftx2x) & (!shiftx3x) & (g137) & (g138) & (g145) & (g146)) + ((!shiftx2x) & (shiftx3x) & (!g137) & (!g138) & (g145) & (!g146)) + ((!shiftx2x) & (shiftx3x) & (!g137) & (!g138) & (g145) & (g146)) + ((!shiftx2x) & (shiftx3x) & (!g137) & (g138) & (g145) & (!g146)) + ((!shiftx2x) & (shiftx3x) & (!g137) & (g138) & (g145) & (g146)) + ((!shiftx2x) & (shiftx3x) & (g137) & (!g138) & (g145) & (!g146)) + ((!shiftx2x) & (shiftx3x) & (g137) & (!g138) & (g145) & (g146)) + ((!shiftx2x) & (shiftx3x) & (g137) & (g138) & (g145) & (!g146)) + ((!shiftx2x) & (shiftx3x) & (g137) & (g138) & (g145) & (g146)) + ((shiftx2x) & (!shiftx3x) & (g137) & (!g138) & (!g145) & (!g146)) + ((shiftx2x) & (!shiftx3x) & (g137) & (!g138) & (!g145) & (g146)) + ((shiftx2x) & (!shiftx3x) & (g137) & (!g138) & (g145) & (!g146)) + ((shiftx2x) & (!shiftx3x) & (g137) & (!g138) & (g145) & (g146)) + ((shiftx2x) & (!shiftx3x) & (g137) & (g138) & (!g145) & (!g146)) + ((shiftx2x) & (!shiftx3x) & (g137) & (g138) & (!g145) & (g146)) + ((shiftx2x) & (!shiftx3x) & (g137) & (g138) & (g145) & (!g146)) + ((shiftx2x) & (!shiftx3x) & (g137) & (g138) & (g145) & (g146)) + ((shiftx2x) & (shiftx3x) & (!g137) & (!g138) & (!g145) & (g146)) + ((shiftx2x) & (shiftx3x) & (!g137) & (!g138) & (g145) & (g146)) + ((shiftx2x) & (shiftx3x) & (!g137) & (g138) & (!g145) & (g146)) + ((shiftx2x) & (shiftx3x) & (!g137) & (g138) & (g145) & (g146)) + ((shiftx2x) & (shiftx3x) & (g137) & (!g138) & (!g145) & (g146)) + ((shiftx2x) & (shiftx3x) & (g137) & (!g138) & (g145) & (g146)) + ((shiftx2x) & (shiftx3x) & (g137) & (g138) & (!g145) & (g146)) + ((shiftx2x) & (shiftx3x) & (g137) & (g138) & (g145) & (g146)));
	assign g253 = (((!shiftx2x) & (!shiftx3x) & (!g140) & (!g141) & (!g147) & (g148)) + ((!shiftx2x) & (!shiftx3x) & (!g140) & (!g141) & (g147) & (g148)) + ((!shiftx2x) & (!shiftx3x) & (!g140) & (g141) & (!g147) & (g148)) + ((!shiftx2x) & (!shiftx3x) & (!g140) & (g141) & (g147) & (g148)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (!g141) & (!g147) & (g148)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (!g141) & (g147) & (g148)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (g141) & (!g147) & (g148)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (g141) & (g147) & (g148)) + ((!shiftx2x) & (shiftx3x) & (g140) & (!g141) & (!g147) & (!g148)) + ((!shiftx2x) & (shiftx3x) & (g140) & (!g141) & (!g147) & (g148)) + ((!shiftx2x) & (shiftx3x) & (g140) & (!g141) & (g147) & (!g148)) + ((!shiftx2x) & (shiftx3x) & (g140) & (!g141) & (g147) & (g148)) + ((!shiftx2x) & (shiftx3x) & (g140) & (g141) & (!g147) & (!g148)) + ((!shiftx2x) & (shiftx3x) & (g140) & (g141) & (!g147) & (g148)) + ((!shiftx2x) & (shiftx3x) & (g140) & (g141) & (g147) & (!g148)) + ((!shiftx2x) & (shiftx3x) & (g140) & (g141) & (g147) & (g148)) + ((shiftx2x) & (!shiftx3x) & (!g140) & (!g141) & (g147) & (!g148)) + ((shiftx2x) & (!shiftx3x) & (!g140) & (!g141) & (g147) & (g148)) + ((shiftx2x) & (!shiftx3x) & (!g140) & (g141) & (g147) & (!g148)) + ((shiftx2x) & (!shiftx3x) & (!g140) & (g141) & (g147) & (g148)) + ((shiftx2x) & (!shiftx3x) & (g140) & (!g141) & (g147) & (!g148)) + ((shiftx2x) & (!shiftx3x) & (g140) & (!g141) & (g147) & (g148)) + ((shiftx2x) & (!shiftx3x) & (g140) & (g141) & (g147) & (!g148)) + ((shiftx2x) & (!shiftx3x) & (g140) & (g141) & (g147) & (g148)) + ((shiftx2x) & (shiftx3x) & (!g140) & (g141) & (!g147) & (!g148)) + ((shiftx2x) & (shiftx3x) & (!g140) & (g141) & (!g147) & (g148)) + ((shiftx2x) & (shiftx3x) & (!g140) & (g141) & (g147) & (!g148)) + ((shiftx2x) & (shiftx3x) & (!g140) & (g141) & (g147) & (g148)) + ((shiftx2x) & (shiftx3x) & (g140) & (g141) & (!g147) & (!g148)) + ((shiftx2x) & (shiftx3x) & (g140) & (g141) & (!g147) & (g148)) + ((shiftx2x) & (shiftx3x) & (g140) & (g141) & (g147) & (!g148)) + ((shiftx2x) & (shiftx3x) & (g140) & (g141) & (g147) & (g148)));
	assign g254 = (((!shiftx4x) & (!shiftx5x) & (!g250) & (g251) & (!g252) & (!g253)) + ((!shiftx4x) & (!shiftx5x) & (!g250) & (g251) & (!g252) & (g253)) + ((!shiftx4x) & (!shiftx5x) & (!g250) & (g251) & (g252) & (!g253)) + ((!shiftx4x) & (!shiftx5x) & (!g250) & (g251) & (g252) & (g253)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (g251) & (!g252) & (!g253)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (g251) & (!g252) & (g253)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (g251) & (g252) & (!g253)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (g251) & (g252) & (g253)) + ((!shiftx4x) & (shiftx5x) & (!g250) & (!g251) & (g252) & (!g253)) + ((!shiftx4x) & (shiftx5x) & (!g250) & (!g251) & (g252) & (g253)) + ((!shiftx4x) & (shiftx5x) & (!g250) & (g251) & (g252) & (!g253)) + ((!shiftx4x) & (shiftx5x) & (!g250) & (g251) & (g252) & (g253)) + ((!shiftx4x) & (shiftx5x) & (g250) & (!g251) & (g252) & (!g253)) + ((!shiftx4x) & (shiftx5x) & (g250) & (!g251) & (g252) & (g253)) + ((!shiftx4x) & (shiftx5x) & (g250) & (g251) & (g252) & (!g253)) + ((!shiftx4x) & (shiftx5x) & (g250) & (g251) & (g252) & (g253)) + ((shiftx4x) & (!shiftx5x) & (g250) & (!g251) & (!g252) & (!g253)) + ((shiftx4x) & (!shiftx5x) & (g250) & (!g251) & (!g252) & (g253)) + ((shiftx4x) & (!shiftx5x) & (g250) & (!g251) & (g252) & (!g253)) + ((shiftx4x) & (!shiftx5x) & (g250) & (!g251) & (g252) & (g253)) + ((shiftx4x) & (!shiftx5x) & (g250) & (g251) & (!g252) & (!g253)) + ((shiftx4x) & (!shiftx5x) & (g250) & (g251) & (!g252) & (g253)) + ((shiftx4x) & (!shiftx5x) & (g250) & (g251) & (g252) & (!g253)) + ((shiftx4x) & (!shiftx5x) & (g250) & (g251) & (g252) & (g253)) + ((shiftx4x) & (shiftx5x) & (!g250) & (!g251) & (!g252) & (g253)) + ((shiftx4x) & (shiftx5x) & (!g250) & (!g251) & (g252) & (g253)) + ((shiftx4x) & (shiftx5x) & (!g250) & (g251) & (!g252) & (g253)) + ((shiftx4x) & (shiftx5x) & (!g250) & (g251) & (g252) & (g253)) + ((shiftx4x) & (shiftx5x) & (g250) & (!g251) & (!g252) & (g253)) + ((shiftx4x) & (shiftx5x) & (g250) & (!g251) & (g252) & (g253)) + ((shiftx4x) & (shiftx5x) & (g250) & (g251) & (!g252) & (g253)) + ((shiftx4x) & (shiftx5x) & (g250) & (g251) & (g252) & (g253)));
	assign g255 = (((!shiftx2x) & (!shiftx3x) & (!g158) & (g159) & (!g166) & (!g167)) + ((!shiftx2x) & (!shiftx3x) & (!g158) & (g159) & (!g166) & (g167)) + ((!shiftx2x) & (!shiftx3x) & (!g158) & (g159) & (g166) & (!g167)) + ((!shiftx2x) & (!shiftx3x) & (!g158) & (g159) & (g166) & (g167)) + ((!shiftx2x) & (!shiftx3x) & (g158) & (g159) & (!g166) & (!g167)) + ((!shiftx2x) & (!shiftx3x) & (g158) & (g159) & (!g166) & (g167)) + ((!shiftx2x) & (!shiftx3x) & (g158) & (g159) & (g166) & (!g167)) + ((!shiftx2x) & (!shiftx3x) & (g158) & (g159) & (g166) & (g167)) + ((!shiftx2x) & (shiftx3x) & (!g158) & (!g159) & (g166) & (!g167)) + ((!shiftx2x) & (shiftx3x) & (!g158) & (!g159) & (g166) & (g167)) + ((!shiftx2x) & (shiftx3x) & (!g158) & (g159) & (g166) & (!g167)) + ((!shiftx2x) & (shiftx3x) & (!g158) & (g159) & (g166) & (g167)) + ((!shiftx2x) & (shiftx3x) & (g158) & (!g159) & (g166) & (!g167)) + ((!shiftx2x) & (shiftx3x) & (g158) & (!g159) & (g166) & (g167)) + ((!shiftx2x) & (shiftx3x) & (g158) & (g159) & (g166) & (!g167)) + ((!shiftx2x) & (shiftx3x) & (g158) & (g159) & (g166) & (g167)) + ((shiftx2x) & (!shiftx3x) & (g158) & (!g159) & (!g166) & (!g167)) + ((shiftx2x) & (!shiftx3x) & (g158) & (!g159) & (!g166) & (g167)) + ((shiftx2x) & (!shiftx3x) & (g158) & (!g159) & (g166) & (!g167)) + ((shiftx2x) & (!shiftx3x) & (g158) & (!g159) & (g166) & (g167)) + ((shiftx2x) & (!shiftx3x) & (g158) & (g159) & (!g166) & (!g167)) + ((shiftx2x) & (!shiftx3x) & (g158) & (g159) & (!g166) & (g167)) + ((shiftx2x) & (!shiftx3x) & (g158) & (g159) & (g166) & (!g167)) + ((shiftx2x) & (!shiftx3x) & (g158) & (g159) & (g166) & (g167)) + ((shiftx2x) & (shiftx3x) & (!g158) & (!g159) & (!g166) & (g167)) + ((shiftx2x) & (shiftx3x) & (!g158) & (!g159) & (g166) & (g167)) + ((shiftx2x) & (shiftx3x) & (!g158) & (g159) & (!g166) & (g167)) + ((shiftx2x) & (shiftx3x) & (!g158) & (g159) & (g166) & (g167)) + ((shiftx2x) & (shiftx3x) & (g158) & (!g159) & (!g166) & (g167)) + ((shiftx2x) & (shiftx3x) & (g158) & (!g159) & (g166) & (g167)) + ((shiftx2x) & (shiftx3x) & (g158) & (g159) & (!g166) & (g167)) + ((shiftx2x) & (shiftx3x) & (g158) & (g159) & (g166) & (g167)));
	assign g256 = (((!shiftx2x) & (!shiftx3x) & (!g153) & (g154) & (!g156) & (!g157)) + ((!shiftx2x) & (!shiftx3x) & (!g153) & (g154) & (!g156) & (g157)) + ((!shiftx2x) & (!shiftx3x) & (!g153) & (g154) & (g156) & (!g157)) + ((!shiftx2x) & (!shiftx3x) & (!g153) & (g154) & (g156) & (g157)) + ((!shiftx2x) & (!shiftx3x) & (g153) & (g154) & (!g156) & (!g157)) + ((!shiftx2x) & (!shiftx3x) & (g153) & (g154) & (!g156) & (g157)) + ((!shiftx2x) & (!shiftx3x) & (g153) & (g154) & (g156) & (!g157)) + ((!shiftx2x) & (!shiftx3x) & (g153) & (g154) & (g156) & (g157)) + ((!shiftx2x) & (shiftx3x) & (!g153) & (!g154) & (g156) & (!g157)) + ((!shiftx2x) & (shiftx3x) & (!g153) & (!g154) & (g156) & (g157)) + ((!shiftx2x) & (shiftx3x) & (!g153) & (g154) & (g156) & (!g157)) + ((!shiftx2x) & (shiftx3x) & (!g153) & (g154) & (g156) & (g157)) + ((!shiftx2x) & (shiftx3x) & (g153) & (!g154) & (g156) & (!g157)) + ((!shiftx2x) & (shiftx3x) & (g153) & (!g154) & (g156) & (g157)) + ((!shiftx2x) & (shiftx3x) & (g153) & (g154) & (g156) & (!g157)) + ((!shiftx2x) & (shiftx3x) & (g153) & (g154) & (g156) & (g157)) + ((shiftx2x) & (!shiftx3x) & (g153) & (!g154) & (!g156) & (!g157)) + ((shiftx2x) & (!shiftx3x) & (g153) & (!g154) & (!g156) & (g157)) + ((shiftx2x) & (!shiftx3x) & (g153) & (!g154) & (g156) & (!g157)) + ((shiftx2x) & (!shiftx3x) & (g153) & (!g154) & (g156) & (g157)) + ((shiftx2x) & (!shiftx3x) & (g153) & (g154) & (!g156) & (!g157)) + ((shiftx2x) & (!shiftx3x) & (g153) & (g154) & (!g156) & (g157)) + ((shiftx2x) & (!shiftx3x) & (g153) & (g154) & (g156) & (!g157)) + ((shiftx2x) & (!shiftx3x) & (g153) & (g154) & (g156) & (g157)) + ((shiftx2x) & (shiftx3x) & (!g153) & (!g154) & (!g156) & (g157)) + ((shiftx2x) & (shiftx3x) & (!g153) & (!g154) & (g156) & (g157)) + ((shiftx2x) & (shiftx3x) & (!g153) & (g154) & (!g156) & (g157)) + ((shiftx2x) & (shiftx3x) & (!g153) & (g154) & (g156) & (g157)) + ((shiftx2x) & (shiftx3x) & (g153) & (!g154) & (!g156) & (g157)) + ((shiftx2x) & (shiftx3x) & (g153) & (!g154) & (g156) & (g157)) + ((shiftx2x) & (shiftx3x) & (g153) & (g154) & (!g156) & (g157)) + ((shiftx2x) & (shiftx3x) & (g153) & (g154) & (g156) & (g157)));
	assign g257 = (((!shiftx2x) & (!shiftx3x) & (!g142) & (g143) & (!g161) & (!g162)) + ((!shiftx2x) & (!shiftx3x) & (!g142) & (g143) & (!g161) & (g162)) + ((!shiftx2x) & (!shiftx3x) & (!g142) & (g143) & (g161) & (!g162)) + ((!shiftx2x) & (!shiftx3x) & (!g142) & (g143) & (g161) & (g162)) + ((!shiftx2x) & (!shiftx3x) & (g142) & (g143) & (!g161) & (!g162)) + ((!shiftx2x) & (!shiftx3x) & (g142) & (g143) & (!g161) & (g162)) + ((!shiftx2x) & (!shiftx3x) & (g142) & (g143) & (g161) & (!g162)) + ((!shiftx2x) & (!shiftx3x) & (g142) & (g143) & (g161) & (g162)) + ((!shiftx2x) & (shiftx3x) & (!g142) & (!g143) & (g161) & (!g162)) + ((!shiftx2x) & (shiftx3x) & (!g142) & (!g143) & (g161) & (g162)) + ((!shiftx2x) & (shiftx3x) & (!g142) & (g143) & (g161) & (!g162)) + ((!shiftx2x) & (shiftx3x) & (!g142) & (g143) & (g161) & (g162)) + ((!shiftx2x) & (shiftx3x) & (g142) & (!g143) & (g161) & (!g162)) + ((!shiftx2x) & (shiftx3x) & (g142) & (!g143) & (g161) & (g162)) + ((!shiftx2x) & (shiftx3x) & (g142) & (g143) & (g161) & (!g162)) + ((!shiftx2x) & (shiftx3x) & (g142) & (g143) & (g161) & (g162)) + ((shiftx2x) & (!shiftx3x) & (g142) & (!g143) & (!g161) & (!g162)) + ((shiftx2x) & (!shiftx3x) & (g142) & (!g143) & (!g161) & (g162)) + ((shiftx2x) & (!shiftx3x) & (g142) & (!g143) & (g161) & (!g162)) + ((shiftx2x) & (!shiftx3x) & (g142) & (!g143) & (g161) & (g162)) + ((shiftx2x) & (!shiftx3x) & (g142) & (g143) & (!g161) & (!g162)) + ((shiftx2x) & (!shiftx3x) & (g142) & (g143) & (!g161) & (g162)) + ((shiftx2x) & (!shiftx3x) & (g142) & (g143) & (g161) & (!g162)) + ((shiftx2x) & (!shiftx3x) & (g142) & (g143) & (g161) & (g162)) + ((shiftx2x) & (shiftx3x) & (!g142) & (!g143) & (!g161) & (g162)) + ((shiftx2x) & (shiftx3x) & (!g142) & (!g143) & (g161) & (g162)) + ((shiftx2x) & (shiftx3x) & (!g142) & (g143) & (!g161) & (g162)) + ((shiftx2x) & (shiftx3x) & (!g142) & (g143) & (g161) & (g162)) + ((shiftx2x) & (shiftx3x) & (g142) & (!g143) & (!g161) & (g162)) + ((shiftx2x) & (shiftx3x) & (g142) & (!g143) & (g161) & (g162)) + ((shiftx2x) & (shiftx3x) & (g142) & (g143) & (!g161) & (g162)) + ((shiftx2x) & (shiftx3x) & (g142) & (g143) & (g161) & (g162)));
	assign g258 = (((!shiftx2x) & (!shiftx3x) & (!g151) & (!g152) & (!g163) & (g164)) + ((!shiftx2x) & (!shiftx3x) & (!g151) & (!g152) & (g163) & (g164)) + ((!shiftx2x) & (!shiftx3x) & (!g151) & (g152) & (!g163) & (g164)) + ((!shiftx2x) & (!shiftx3x) & (!g151) & (g152) & (g163) & (g164)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (!g152) & (!g163) & (g164)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (!g152) & (g163) & (g164)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (g152) & (!g163) & (g164)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (g152) & (g163) & (g164)) + ((!shiftx2x) & (shiftx3x) & (g151) & (!g152) & (!g163) & (!g164)) + ((!shiftx2x) & (shiftx3x) & (g151) & (!g152) & (!g163) & (g164)) + ((!shiftx2x) & (shiftx3x) & (g151) & (!g152) & (g163) & (!g164)) + ((!shiftx2x) & (shiftx3x) & (g151) & (!g152) & (g163) & (g164)) + ((!shiftx2x) & (shiftx3x) & (g151) & (g152) & (!g163) & (!g164)) + ((!shiftx2x) & (shiftx3x) & (g151) & (g152) & (!g163) & (g164)) + ((!shiftx2x) & (shiftx3x) & (g151) & (g152) & (g163) & (!g164)) + ((!shiftx2x) & (shiftx3x) & (g151) & (g152) & (g163) & (g164)) + ((shiftx2x) & (!shiftx3x) & (!g151) & (!g152) & (g163) & (!g164)) + ((shiftx2x) & (!shiftx3x) & (!g151) & (!g152) & (g163) & (g164)) + ((shiftx2x) & (!shiftx3x) & (!g151) & (g152) & (g163) & (!g164)) + ((shiftx2x) & (!shiftx3x) & (!g151) & (g152) & (g163) & (g164)) + ((shiftx2x) & (!shiftx3x) & (g151) & (!g152) & (g163) & (!g164)) + ((shiftx2x) & (!shiftx3x) & (g151) & (!g152) & (g163) & (g164)) + ((shiftx2x) & (!shiftx3x) & (g151) & (g152) & (g163) & (!g164)) + ((shiftx2x) & (!shiftx3x) & (g151) & (g152) & (g163) & (g164)) + ((shiftx2x) & (shiftx3x) & (!g151) & (g152) & (!g163) & (!g164)) + ((shiftx2x) & (shiftx3x) & (!g151) & (g152) & (!g163) & (g164)) + ((shiftx2x) & (shiftx3x) & (!g151) & (g152) & (g163) & (!g164)) + ((shiftx2x) & (shiftx3x) & (!g151) & (g152) & (g163) & (g164)) + ((shiftx2x) & (shiftx3x) & (g151) & (g152) & (!g163) & (!g164)) + ((shiftx2x) & (shiftx3x) & (g151) & (g152) & (!g163) & (g164)) + ((shiftx2x) & (shiftx3x) & (g151) & (g152) & (g163) & (!g164)) + ((shiftx2x) & (shiftx3x) & (g151) & (g152) & (g163) & (g164)));
	assign g259 = (((!shiftx4x) & (!shiftx5x) & (!g255) & (!g256) & (g257) & (!g258)) + ((!shiftx4x) & (!shiftx5x) & (!g255) & (!g256) & (g257) & (g258)) + ((!shiftx4x) & (!shiftx5x) & (!g255) & (g256) & (g257) & (!g258)) + ((!shiftx4x) & (!shiftx5x) & (!g255) & (g256) & (g257) & (g258)) + ((!shiftx4x) & (!shiftx5x) & (g255) & (!g256) & (g257) & (!g258)) + ((!shiftx4x) & (!shiftx5x) & (g255) & (!g256) & (g257) & (g258)) + ((!shiftx4x) & (!shiftx5x) & (g255) & (g256) & (g257) & (!g258)) + ((!shiftx4x) & (!shiftx5x) & (g255) & (g256) & (g257) & (g258)) + ((!shiftx4x) & (shiftx5x) & (!g255) & (g256) & (!g257) & (!g258)) + ((!shiftx4x) & (shiftx5x) & (!g255) & (g256) & (!g257) & (g258)) + ((!shiftx4x) & (shiftx5x) & (!g255) & (g256) & (g257) & (!g258)) + ((!shiftx4x) & (shiftx5x) & (!g255) & (g256) & (g257) & (g258)) + ((!shiftx4x) & (shiftx5x) & (g255) & (g256) & (!g257) & (!g258)) + ((!shiftx4x) & (shiftx5x) & (g255) & (g256) & (!g257) & (g258)) + ((!shiftx4x) & (shiftx5x) & (g255) & (g256) & (g257) & (!g258)) + ((!shiftx4x) & (shiftx5x) & (g255) & (g256) & (g257) & (g258)) + ((shiftx4x) & (!shiftx5x) & (!g255) & (!g256) & (!g257) & (g258)) + ((shiftx4x) & (!shiftx5x) & (!g255) & (!g256) & (g257) & (g258)) + ((shiftx4x) & (!shiftx5x) & (!g255) & (g256) & (!g257) & (g258)) + ((shiftx4x) & (!shiftx5x) & (!g255) & (g256) & (g257) & (g258)) + ((shiftx4x) & (!shiftx5x) & (g255) & (!g256) & (!g257) & (g258)) + ((shiftx4x) & (!shiftx5x) & (g255) & (!g256) & (g257) & (g258)) + ((shiftx4x) & (!shiftx5x) & (g255) & (g256) & (!g257) & (g258)) + ((shiftx4x) & (!shiftx5x) & (g255) & (g256) & (g257) & (g258)) + ((shiftx4x) & (shiftx5x) & (g255) & (!g256) & (!g257) & (!g258)) + ((shiftx4x) & (shiftx5x) & (g255) & (!g256) & (!g257) & (g258)) + ((shiftx4x) & (shiftx5x) & (g255) & (!g256) & (g257) & (!g258)) + ((shiftx4x) & (shiftx5x) & (g255) & (!g256) & (g257) & (g258)) + ((shiftx4x) & (shiftx5x) & (g255) & (g256) & (!g257) & (!g258)) + ((shiftx4x) & (shiftx5x) & (g255) & (g256) & (!g257) & (g258)) + ((shiftx4x) & (shiftx5x) & (g255) & (g256) & (g257) & (!g258)) + ((shiftx4x) & (shiftx5x) & (g255) & (g256) & (g257) & (g258)));
	assign resultx11x = (((!shiftx6x) & (sk[3]) & (!g254) & (g259)) + ((!shiftx6x) & (sk[3]) & (g254) & (g259)) + ((shiftx6x) & (!sk[3]) & (!g254) & (!g259)) + ((shiftx6x) & (!sk[3]) & (!g254) & (g259)) + ((shiftx6x) & (!sk[3]) & (g254) & (!g259)) + ((shiftx6x) & (!sk[3]) & (g254) & (g259)) + ((shiftx6x) & (sk[3]) & (g254) & (!g259)) + ((shiftx6x) & (sk[3]) & (g254) & (g259)));
	assign g261 = (((!shiftx2x) & (!shiftx3x) & (g12) & (!g13) & (!g14) & (!g16)) + ((!shiftx2x) & (!shiftx3x) & (g12) & (!g13) & (!g14) & (g16)) + ((!shiftx2x) & (!shiftx3x) & (g12) & (!g13) & (g14) & (!g16)) + ((!shiftx2x) & (!shiftx3x) & (g12) & (!g13) & (g14) & (g16)) + ((!shiftx2x) & (!shiftx3x) & (g12) & (g13) & (!g14) & (!g16)) + ((!shiftx2x) & (!shiftx3x) & (g12) & (g13) & (!g14) & (g16)) + ((!shiftx2x) & (!shiftx3x) & (g12) & (g13) & (g14) & (!g16)) + ((!shiftx2x) & (!shiftx3x) & (g12) & (g13) & (g14) & (g16)) + ((!shiftx2x) & (shiftx3x) & (!g12) & (g13) & (!g14) & (!g16)) + ((!shiftx2x) & (shiftx3x) & (!g12) & (g13) & (!g14) & (g16)) + ((!shiftx2x) & (shiftx3x) & (!g12) & (g13) & (g14) & (!g16)) + ((!shiftx2x) & (shiftx3x) & (!g12) & (g13) & (g14) & (g16)) + ((!shiftx2x) & (shiftx3x) & (g12) & (g13) & (!g14) & (!g16)) + ((!shiftx2x) & (shiftx3x) & (g12) & (g13) & (!g14) & (g16)) + ((!shiftx2x) & (shiftx3x) & (g12) & (g13) & (g14) & (!g16)) + ((!shiftx2x) & (shiftx3x) & (g12) & (g13) & (g14) & (g16)) + ((shiftx2x) & (!shiftx3x) & (!g12) & (!g13) & (g14) & (!g16)) + ((shiftx2x) & (!shiftx3x) & (!g12) & (!g13) & (g14) & (g16)) + ((shiftx2x) & (!shiftx3x) & (!g12) & (g13) & (g14) & (!g16)) + ((shiftx2x) & (!shiftx3x) & (!g12) & (g13) & (g14) & (g16)) + ((shiftx2x) & (!shiftx3x) & (g12) & (!g13) & (g14) & (!g16)) + ((shiftx2x) & (!shiftx3x) & (g12) & (!g13) & (g14) & (g16)) + ((shiftx2x) & (!shiftx3x) & (g12) & (g13) & (g14) & (!g16)) + ((shiftx2x) & (!shiftx3x) & (g12) & (g13) & (g14) & (g16)) + ((shiftx2x) & (shiftx3x) & (!g12) & (!g13) & (!g14) & (g16)) + ((shiftx2x) & (shiftx3x) & (!g12) & (!g13) & (g14) & (g16)) + ((shiftx2x) & (shiftx3x) & (!g12) & (g13) & (!g14) & (g16)) + ((shiftx2x) & (shiftx3x) & (!g12) & (g13) & (g14) & (g16)) + ((shiftx2x) & (shiftx3x) & (g12) & (!g13) & (!g14) & (g16)) + ((shiftx2x) & (shiftx3x) & (g12) & (!g13) & (g14) & (g16)) + ((shiftx2x) & (shiftx3x) & (g12) & (g13) & (!g14) & (g16)) + ((shiftx2x) & (shiftx3x) & (g12) & (g13) & (g14) & (g16)));
	assign g262 = (((!shiftx2x) & (!shiftx3x) & (!g11) & (g23) & (!g24) & (!g25)) + ((!shiftx2x) & (!shiftx3x) & (!g11) & (g23) & (!g24) & (g25)) + ((!shiftx2x) & (!shiftx3x) & (!g11) & (g23) & (g24) & (!g25)) + ((!shiftx2x) & (!shiftx3x) & (!g11) & (g23) & (g24) & (g25)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (g23) & (!g24) & (!g25)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (g23) & (!g24) & (g25)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (g23) & (g24) & (!g25)) + ((!shiftx2x) & (!shiftx3x) & (g11) & (g23) & (g24) & (g25)) + ((!shiftx2x) & (shiftx3x) & (!g11) & (!g23) & (g24) & (!g25)) + ((!shiftx2x) & (shiftx3x) & (!g11) & (!g23) & (g24) & (g25)) + ((!shiftx2x) & (shiftx3x) & (!g11) & (g23) & (g24) & (!g25)) + ((!shiftx2x) & (shiftx3x) & (!g11) & (g23) & (g24) & (g25)) + ((!shiftx2x) & (shiftx3x) & (g11) & (!g23) & (g24) & (!g25)) + ((!shiftx2x) & (shiftx3x) & (g11) & (!g23) & (g24) & (g25)) + ((!shiftx2x) & (shiftx3x) & (g11) & (g23) & (g24) & (!g25)) + ((!shiftx2x) & (shiftx3x) & (g11) & (g23) & (g24) & (g25)) + ((shiftx2x) & (!shiftx3x) & (!g11) & (!g23) & (!g24) & (g25)) + ((shiftx2x) & (!shiftx3x) & (!g11) & (!g23) & (g24) & (g25)) + ((shiftx2x) & (!shiftx3x) & (!g11) & (g23) & (!g24) & (g25)) + ((shiftx2x) & (!shiftx3x) & (!g11) & (g23) & (g24) & (g25)) + ((shiftx2x) & (!shiftx3x) & (g11) & (!g23) & (!g24) & (g25)) + ((shiftx2x) & (!shiftx3x) & (g11) & (!g23) & (g24) & (g25)) + ((shiftx2x) & (!shiftx3x) & (g11) & (g23) & (!g24) & (g25)) + ((shiftx2x) & (!shiftx3x) & (g11) & (g23) & (g24) & (g25)) + ((shiftx2x) & (shiftx3x) & (g11) & (!g23) & (!g24) & (!g25)) + ((shiftx2x) & (shiftx3x) & (g11) & (!g23) & (!g24) & (g25)) + ((shiftx2x) & (shiftx3x) & (g11) & (!g23) & (g24) & (!g25)) + ((shiftx2x) & (shiftx3x) & (g11) & (!g23) & (g24) & (g25)) + ((shiftx2x) & (shiftx3x) & (g11) & (g23) & (!g24) & (!g25)) + ((shiftx2x) & (shiftx3x) & (g11) & (g23) & (!g24) & (g25)) + ((shiftx2x) & (shiftx3x) & (g11) & (g23) & (g24) & (!g25)) + ((shiftx2x) & (shiftx3x) & (g11) & (g23) & (g24) & (g25)));
	assign g263 = (((!shiftx2x) & (!shiftx3x) & (!g6) & (g17) & (!g18) & (!g19)) + ((!shiftx2x) & (!shiftx3x) & (!g6) & (g17) & (!g18) & (g19)) + ((!shiftx2x) & (!shiftx3x) & (!g6) & (g17) & (g18) & (!g19)) + ((!shiftx2x) & (!shiftx3x) & (!g6) & (g17) & (g18) & (g19)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (g17) & (!g18) & (!g19)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (g17) & (!g18) & (g19)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (g17) & (g18) & (!g19)) + ((!shiftx2x) & (!shiftx3x) & (g6) & (g17) & (g18) & (g19)) + ((!shiftx2x) & (shiftx3x) & (!g6) & (!g17) & (g18) & (!g19)) + ((!shiftx2x) & (shiftx3x) & (!g6) & (!g17) & (g18) & (g19)) + ((!shiftx2x) & (shiftx3x) & (!g6) & (g17) & (g18) & (!g19)) + ((!shiftx2x) & (shiftx3x) & (!g6) & (g17) & (g18) & (g19)) + ((!shiftx2x) & (shiftx3x) & (g6) & (!g17) & (g18) & (!g19)) + ((!shiftx2x) & (shiftx3x) & (g6) & (!g17) & (g18) & (g19)) + ((!shiftx2x) & (shiftx3x) & (g6) & (g17) & (g18) & (!g19)) + ((!shiftx2x) & (shiftx3x) & (g6) & (g17) & (g18) & (g19)) + ((shiftx2x) & (!shiftx3x) & (!g6) & (!g17) & (!g18) & (g19)) + ((shiftx2x) & (!shiftx3x) & (!g6) & (!g17) & (g18) & (g19)) + ((shiftx2x) & (!shiftx3x) & (!g6) & (g17) & (!g18) & (g19)) + ((shiftx2x) & (!shiftx3x) & (!g6) & (g17) & (g18) & (g19)) + ((shiftx2x) & (!shiftx3x) & (g6) & (!g17) & (!g18) & (g19)) + ((shiftx2x) & (!shiftx3x) & (g6) & (!g17) & (g18) & (g19)) + ((shiftx2x) & (!shiftx3x) & (g6) & (g17) & (!g18) & (g19)) + ((shiftx2x) & (!shiftx3x) & (g6) & (g17) & (g18) & (g19)) + ((shiftx2x) & (shiftx3x) & (g6) & (!g17) & (!g18) & (!g19)) + ((shiftx2x) & (shiftx3x) & (g6) & (!g17) & (!g18) & (g19)) + ((shiftx2x) & (shiftx3x) & (g6) & (!g17) & (g18) & (!g19)) + ((shiftx2x) & (shiftx3x) & (g6) & (!g17) & (g18) & (g19)) + ((shiftx2x) & (shiftx3x) & (g6) & (g17) & (!g18) & (!g19)) + ((shiftx2x) & (shiftx3x) & (g6) & (g17) & (!g18) & (g19)) + ((shiftx2x) & (shiftx3x) & (g6) & (g17) & (g18) & (!g19)) + ((shiftx2x) & (shiftx3x) & (g6) & (g17) & (g18) & (g19)));
	assign g264 = (((!shiftx2x) & (!shiftx3x) & (!g1) & (g7) & (!g8) & (!g9)) + ((!shiftx2x) & (!shiftx3x) & (!g1) & (g7) & (!g8) & (g9)) + ((!shiftx2x) & (!shiftx3x) & (!g1) & (g7) & (g8) & (!g9)) + ((!shiftx2x) & (!shiftx3x) & (!g1) & (g7) & (g8) & (g9)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (g7) & (!g8) & (!g9)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (g7) & (!g8) & (g9)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (g7) & (g8) & (!g9)) + ((!shiftx2x) & (!shiftx3x) & (g1) & (g7) & (g8) & (g9)) + ((!shiftx2x) & (shiftx3x) & (!g1) & (!g7) & (g8) & (!g9)) + ((!shiftx2x) & (shiftx3x) & (!g1) & (!g7) & (g8) & (g9)) + ((!shiftx2x) & (shiftx3x) & (!g1) & (g7) & (g8) & (!g9)) + ((!shiftx2x) & (shiftx3x) & (!g1) & (g7) & (g8) & (g9)) + ((!shiftx2x) & (shiftx3x) & (g1) & (!g7) & (g8) & (!g9)) + ((!shiftx2x) & (shiftx3x) & (g1) & (!g7) & (g8) & (g9)) + ((!shiftx2x) & (shiftx3x) & (g1) & (g7) & (g8) & (!g9)) + ((!shiftx2x) & (shiftx3x) & (g1) & (g7) & (g8) & (g9)) + ((shiftx2x) & (!shiftx3x) & (!g1) & (!g7) & (!g8) & (g9)) + ((shiftx2x) & (!shiftx3x) & (!g1) & (!g7) & (g8) & (g9)) + ((shiftx2x) & (!shiftx3x) & (!g1) & (g7) & (!g8) & (g9)) + ((shiftx2x) & (!shiftx3x) & (!g1) & (g7) & (g8) & (g9)) + ((shiftx2x) & (!shiftx3x) & (g1) & (!g7) & (!g8) & (g9)) + ((shiftx2x) & (!shiftx3x) & (g1) & (!g7) & (g8) & (g9)) + ((shiftx2x) & (!shiftx3x) & (g1) & (g7) & (!g8) & (g9)) + ((shiftx2x) & (!shiftx3x) & (g1) & (g7) & (g8) & (g9)) + ((shiftx2x) & (shiftx3x) & (g1) & (!g7) & (!g8) & (!g9)) + ((shiftx2x) & (shiftx3x) & (g1) & (!g7) & (!g8) & (g9)) + ((shiftx2x) & (shiftx3x) & (g1) & (!g7) & (g8) & (!g9)) + ((shiftx2x) & (shiftx3x) & (g1) & (!g7) & (g8) & (g9)) + ((shiftx2x) & (shiftx3x) & (g1) & (g7) & (!g8) & (!g9)) + ((shiftx2x) & (shiftx3x) & (g1) & (g7) & (!g8) & (g9)) + ((shiftx2x) & (shiftx3x) & (g1) & (g7) & (g8) & (!g9)) + ((shiftx2x) & (shiftx3x) & (g1) & (g7) & (g8) & (g9)));
	assign g265 = (((!shiftx4x) & (!shiftx5x) & (!g261) & (g262) & (!g263) & (!g264)) + ((!shiftx4x) & (!shiftx5x) & (!g261) & (g262) & (!g263) & (g264)) + ((!shiftx4x) & (!shiftx5x) & (!g261) & (g262) & (g263) & (!g264)) + ((!shiftx4x) & (!shiftx5x) & (!g261) & (g262) & (g263) & (g264)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (g262) & (!g263) & (!g264)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (g262) & (!g263) & (g264)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (g262) & (g263) & (!g264)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (g262) & (g263) & (g264)) + ((!shiftx4x) & (shiftx5x) & (!g261) & (!g262) & (g263) & (!g264)) + ((!shiftx4x) & (shiftx5x) & (!g261) & (!g262) & (g263) & (g264)) + ((!shiftx4x) & (shiftx5x) & (!g261) & (g262) & (g263) & (!g264)) + ((!shiftx4x) & (shiftx5x) & (!g261) & (g262) & (g263) & (g264)) + ((!shiftx4x) & (shiftx5x) & (g261) & (!g262) & (g263) & (!g264)) + ((!shiftx4x) & (shiftx5x) & (g261) & (!g262) & (g263) & (g264)) + ((!shiftx4x) & (shiftx5x) & (g261) & (g262) & (g263) & (!g264)) + ((!shiftx4x) & (shiftx5x) & (g261) & (g262) & (g263) & (g264)) + ((shiftx4x) & (!shiftx5x) & (g261) & (!g262) & (!g263) & (!g264)) + ((shiftx4x) & (!shiftx5x) & (g261) & (!g262) & (!g263) & (g264)) + ((shiftx4x) & (!shiftx5x) & (g261) & (!g262) & (g263) & (!g264)) + ((shiftx4x) & (!shiftx5x) & (g261) & (!g262) & (g263) & (g264)) + ((shiftx4x) & (!shiftx5x) & (g261) & (g262) & (!g263) & (!g264)) + ((shiftx4x) & (!shiftx5x) & (g261) & (g262) & (!g263) & (g264)) + ((shiftx4x) & (!shiftx5x) & (g261) & (g262) & (g263) & (!g264)) + ((shiftx4x) & (!shiftx5x) & (g261) & (g262) & (g263) & (g264)) + ((shiftx4x) & (shiftx5x) & (!g261) & (!g262) & (!g263) & (g264)) + ((shiftx4x) & (shiftx5x) & (!g261) & (!g262) & (g263) & (g264)) + ((shiftx4x) & (shiftx5x) & (!g261) & (g262) & (!g263) & (g264)) + ((shiftx4x) & (shiftx5x) & (!g261) & (g262) & (g263) & (g264)) + ((shiftx4x) & (shiftx5x) & (g261) & (!g262) & (!g263) & (g264)) + ((shiftx4x) & (shiftx5x) & (g261) & (!g262) & (g263) & (g264)) + ((shiftx4x) & (shiftx5x) & (g261) & (g262) & (!g263) & (g264)) + ((shiftx4x) & (shiftx5x) & (g261) & (g262) & (g263) & (g264)));
	assign g266 = (((!shiftx2x) & (!shiftx3x) & (!g22) & (g28) & (!g29) & (!g30)) + ((!shiftx2x) & (!shiftx3x) & (!g22) & (g28) & (!g29) & (g30)) + ((!shiftx2x) & (!shiftx3x) & (!g22) & (g28) & (g29) & (!g30)) + ((!shiftx2x) & (!shiftx3x) & (!g22) & (g28) & (g29) & (g30)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (g28) & (!g29) & (!g30)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (g28) & (!g29) & (g30)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (g28) & (g29) & (!g30)) + ((!shiftx2x) & (!shiftx3x) & (g22) & (g28) & (g29) & (g30)) + ((!shiftx2x) & (shiftx3x) & (!g22) & (!g28) & (g29) & (!g30)) + ((!shiftx2x) & (shiftx3x) & (!g22) & (!g28) & (g29) & (g30)) + ((!shiftx2x) & (shiftx3x) & (!g22) & (g28) & (g29) & (!g30)) + ((!shiftx2x) & (shiftx3x) & (!g22) & (g28) & (g29) & (g30)) + ((!shiftx2x) & (shiftx3x) & (g22) & (!g28) & (g29) & (!g30)) + ((!shiftx2x) & (shiftx3x) & (g22) & (!g28) & (g29) & (g30)) + ((!shiftx2x) & (shiftx3x) & (g22) & (g28) & (g29) & (!g30)) + ((!shiftx2x) & (shiftx3x) & (g22) & (g28) & (g29) & (g30)) + ((shiftx2x) & (!shiftx3x) & (!g22) & (!g28) & (!g29) & (g30)) + ((shiftx2x) & (!shiftx3x) & (!g22) & (!g28) & (g29) & (g30)) + ((shiftx2x) & (!shiftx3x) & (!g22) & (g28) & (!g29) & (g30)) + ((shiftx2x) & (!shiftx3x) & (!g22) & (g28) & (g29) & (g30)) + ((shiftx2x) & (!shiftx3x) & (g22) & (!g28) & (!g29) & (g30)) + ((shiftx2x) & (!shiftx3x) & (g22) & (!g28) & (g29) & (g30)) + ((shiftx2x) & (!shiftx3x) & (g22) & (g28) & (!g29) & (g30)) + ((shiftx2x) & (!shiftx3x) & (g22) & (g28) & (g29) & (g30)) + ((shiftx2x) & (shiftx3x) & (g22) & (!g28) & (!g29) & (!g30)) + ((shiftx2x) & (shiftx3x) & (g22) & (!g28) & (!g29) & (g30)) + ((shiftx2x) & (shiftx3x) & (g22) & (!g28) & (g29) & (!g30)) + ((shiftx2x) & (shiftx3x) & (g22) & (!g28) & (g29) & (g30)) + ((shiftx2x) & (shiftx3x) & (g22) & (g28) & (!g29) & (!g30)) + ((shiftx2x) & (shiftx3x) & (g22) & (g28) & (!g29) & (g30)) + ((shiftx2x) & (shiftx3x) & (g22) & (g28) & (g29) & (!g30)) + ((shiftx2x) & (shiftx3x) & (g22) & (g28) & (g29) & (g30)));
	assign g267 = (((!shiftx2x) & (!shiftx3x) & (!g27) & (g38) & (!g39) & (!g40)) + ((!shiftx2x) & (!shiftx3x) & (!g27) & (g38) & (!g39) & (g40)) + ((!shiftx2x) & (!shiftx3x) & (!g27) & (g38) & (g39) & (!g40)) + ((!shiftx2x) & (!shiftx3x) & (!g27) & (g38) & (g39) & (g40)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (g38) & (!g39) & (!g40)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (g38) & (!g39) & (g40)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (g38) & (g39) & (!g40)) + ((!shiftx2x) & (!shiftx3x) & (g27) & (g38) & (g39) & (g40)) + ((!shiftx2x) & (shiftx3x) & (!g27) & (!g38) & (g39) & (!g40)) + ((!shiftx2x) & (shiftx3x) & (!g27) & (!g38) & (g39) & (g40)) + ((!shiftx2x) & (shiftx3x) & (!g27) & (g38) & (g39) & (!g40)) + ((!shiftx2x) & (shiftx3x) & (!g27) & (g38) & (g39) & (g40)) + ((!shiftx2x) & (shiftx3x) & (g27) & (!g38) & (g39) & (!g40)) + ((!shiftx2x) & (shiftx3x) & (g27) & (!g38) & (g39) & (g40)) + ((!shiftx2x) & (shiftx3x) & (g27) & (g38) & (g39) & (!g40)) + ((!shiftx2x) & (shiftx3x) & (g27) & (g38) & (g39) & (g40)) + ((shiftx2x) & (!shiftx3x) & (!g27) & (!g38) & (!g39) & (g40)) + ((shiftx2x) & (!shiftx3x) & (!g27) & (!g38) & (g39) & (g40)) + ((shiftx2x) & (!shiftx3x) & (!g27) & (g38) & (!g39) & (g40)) + ((shiftx2x) & (!shiftx3x) & (!g27) & (g38) & (g39) & (g40)) + ((shiftx2x) & (!shiftx3x) & (g27) & (!g38) & (!g39) & (g40)) + ((shiftx2x) & (!shiftx3x) & (g27) & (!g38) & (g39) & (g40)) + ((shiftx2x) & (!shiftx3x) & (g27) & (g38) & (!g39) & (g40)) + ((shiftx2x) & (!shiftx3x) & (g27) & (g38) & (g39) & (g40)) + ((shiftx2x) & (shiftx3x) & (g27) & (!g38) & (!g39) & (!g40)) + ((shiftx2x) & (shiftx3x) & (g27) & (!g38) & (!g39) & (g40)) + ((shiftx2x) & (shiftx3x) & (g27) & (!g38) & (g39) & (!g40)) + ((shiftx2x) & (shiftx3x) & (g27) & (!g38) & (g39) & (g40)) + ((shiftx2x) & (shiftx3x) & (g27) & (g38) & (!g39) & (!g40)) + ((shiftx2x) & (shiftx3x) & (g27) & (g38) & (!g39) & (g40)) + ((shiftx2x) & (shiftx3x) & (g27) & (g38) & (g39) & (!g40)) + ((shiftx2x) & (shiftx3x) & (g27) & (g38) & (g39) & (g40)));
	assign g268 = (((!shiftx2x) & (!shiftx3x) & (g2) & (!g3) & (!g4) & (!g32)) + ((!shiftx2x) & (!shiftx3x) & (g2) & (!g3) & (!g4) & (g32)) + ((!shiftx2x) & (!shiftx3x) & (g2) & (!g3) & (g4) & (!g32)) + ((!shiftx2x) & (!shiftx3x) & (g2) & (!g3) & (g4) & (g32)) + ((!shiftx2x) & (!shiftx3x) & (g2) & (g3) & (!g4) & (!g32)) + ((!shiftx2x) & (!shiftx3x) & (g2) & (g3) & (!g4) & (g32)) + ((!shiftx2x) & (!shiftx3x) & (g2) & (g3) & (g4) & (!g32)) + ((!shiftx2x) & (!shiftx3x) & (g2) & (g3) & (g4) & (g32)) + ((!shiftx2x) & (shiftx3x) & (!g2) & (g3) & (!g4) & (!g32)) + ((!shiftx2x) & (shiftx3x) & (!g2) & (g3) & (!g4) & (g32)) + ((!shiftx2x) & (shiftx3x) & (!g2) & (g3) & (g4) & (!g32)) + ((!shiftx2x) & (shiftx3x) & (!g2) & (g3) & (g4) & (g32)) + ((!shiftx2x) & (shiftx3x) & (g2) & (g3) & (!g4) & (!g32)) + ((!shiftx2x) & (shiftx3x) & (g2) & (g3) & (!g4) & (g32)) + ((!shiftx2x) & (shiftx3x) & (g2) & (g3) & (g4) & (!g32)) + ((!shiftx2x) & (shiftx3x) & (g2) & (g3) & (g4) & (g32)) + ((shiftx2x) & (!shiftx3x) & (!g2) & (!g3) & (g4) & (!g32)) + ((shiftx2x) & (!shiftx3x) & (!g2) & (!g3) & (g4) & (g32)) + ((shiftx2x) & (!shiftx3x) & (!g2) & (g3) & (g4) & (!g32)) + ((shiftx2x) & (!shiftx3x) & (!g2) & (g3) & (g4) & (g32)) + ((shiftx2x) & (!shiftx3x) & (g2) & (!g3) & (g4) & (!g32)) + ((shiftx2x) & (!shiftx3x) & (g2) & (!g3) & (g4) & (g32)) + ((shiftx2x) & (!shiftx3x) & (g2) & (g3) & (g4) & (!g32)) + ((shiftx2x) & (!shiftx3x) & (g2) & (g3) & (g4) & (g32)) + ((shiftx2x) & (shiftx3x) & (!g2) & (!g3) & (!g4) & (g32)) + ((shiftx2x) & (shiftx3x) & (!g2) & (!g3) & (g4) & (g32)) + ((shiftx2x) & (shiftx3x) & (!g2) & (g3) & (!g4) & (g32)) + ((shiftx2x) & (shiftx3x) & (!g2) & (g3) & (g4) & (g32)) + ((shiftx2x) & (shiftx3x) & (g2) & (!g3) & (!g4) & (g32)) + ((shiftx2x) & (shiftx3x) & (g2) & (!g3) & (g4) & (g32)) + ((shiftx2x) & (shiftx3x) & (g2) & (g3) & (!g4) & (g32)) + ((shiftx2x) & (shiftx3x) & (g2) & (g3) & (g4) & (g32)));
	assign g269 = (((!shiftx2x) & (!shiftx3x) & (g33) & (!g34) & (!g35) & (!g37)) + ((!shiftx2x) & (!shiftx3x) & (g33) & (!g34) & (!g35) & (g37)) + ((!shiftx2x) & (!shiftx3x) & (g33) & (!g34) & (g35) & (!g37)) + ((!shiftx2x) & (!shiftx3x) & (g33) & (!g34) & (g35) & (g37)) + ((!shiftx2x) & (!shiftx3x) & (g33) & (g34) & (!g35) & (!g37)) + ((!shiftx2x) & (!shiftx3x) & (g33) & (g34) & (!g35) & (g37)) + ((!shiftx2x) & (!shiftx3x) & (g33) & (g34) & (g35) & (!g37)) + ((!shiftx2x) & (!shiftx3x) & (g33) & (g34) & (g35) & (g37)) + ((!shiftx2x) & (shiftx3x) & (!g33) & (g34) & (!g35) & (!g37)) + ((!shiftx2x) & (shiftx3x) & (!g33) & (g34) & (!g35) & (g37)) + ((!shiftx2x) & (shiftx3x) & (!g33) & (g34) & (g35) & (!g37)) + ((!shiftx2x) & (shiftx3x) & (!g33) & (g34) & (g35) & (g37)) + ((!shiftx2x) & (shiftx3x) & (g33) & (g34) & (!g35) & (!g37)) + ((!shiftx2x) & (shiftx3x) & (g33) & (g34) & (!g35) & (g37)) + ((!shiftx2x) & (shiftx3x) & (g33) & (g34) & (g35) & (!g37)) + ((!shiftx2x) & (shiftx3x) & (g33) & (g34) & (g35) & (g37)) + ((shiftx2x) & (!shiftx3x) & (!g33) & (!g34) & (g35) & (!g37)) + ((shiftx2x) & (!shiftx3x) & (!g33) & (!g34) & (g35) & (g37)) + ((shiftx2x) & (!shiftx3x) & (!g33) & (g34) & (g35) & (!g37)) + ((shiftx2x) & (!shiftx3x) & (!g33) & (g34) & (g35) & (g37)) + ((shiftx2x) & (!shiftx3x) & (g33) & (!g34) & (g35) & (!g37)) + ((shiftx2x) & (!shiftx3x) & (g33) & (!g34) & (g35) & (g37)) + ((shiftx2x) & (!shiftx3x) & (g33) & (g34) & (g35) & (!g37)) + ((shiftx2x) & (!shiftx3x) & (g33) & (g34) & (g35) & (g37)) + ((shiftx2x) & (shiftx3x) & (!g33) & (!g34) & (!g35) & (g37)) + ((shiftx2x) & (shiftx3x) & (!g33) & (!g34) & (g35) & (g37)) + ((shiftx2x) & (shiftx3x) & (!g33) & (g34) & (!g35) & (g37)) + ((shiftx2x) & (shiftx3x) & (!g33) & (g34) & (g35) & (g37)) + ((shiftx2x) & (shiftx3x) & (g33) & (!g34) & (!g35) & (g37)) + ((shiftx2x) & (shiftx3x) & (g33) & (!g34) & (g35) & (g37)) + ((shiftx2x) & (shiftx3x) & (g33) & (g34) & (!g35) & (g37)) + ((shiftx2x) & (shiftx3x) & (g33) & (g34) & (g35) & (g37)));
	assign g270 = (((!shiftx4x) & (!shiftx5x) & (!g266) & (!g267) & (g268) & (!g269)) + ((!shiftx4x) & (!shiftx5x) & (!g266) & (!g267) & (g268) & (g269)) + ((!shiftx4x) & (!shiftx5x) & (!g266) & (g267) & (g268) & (!g269)) + ((!shiftx4x) & (!shiftx5x) & (!g266) & (g267) & (g268) & (g269)) + ((!shiftx4x) & (!shiftx5x) & (g266) & (!g267) & (g268) & (!g269)) + ((!shiftx4x) & (!shiftx5x) & (g266) & (!g267) & (g268) & (g269)) + ((!shiftx4x) & (!shiftx5x) & (g266) & (g267) & (g268) & (!g269)) + ((!shiftx4x) & (!shiftx5x) & (g266) & (g267) & (g268) & (g269)) + ((!shiftx4x) & (shiftx5x) & (!g266) & (g267) & (!g268) & (!g269)) + ((!shiftx4x) & (shiftx5x) & (!g266) & (g267) & (!g268) & (g269)) + ((!shiftx4x) & (shiftx5x) & (!g266) & (g267) & (g268) & (!g269)) + ((!shiftx4x) & (shiftx5x) & (!g266) & (g267) & (g268) & (g269)) + ((!shiftx4x) & (shiftx5x) & (g266) & (g267) & (!g268) & (!g269)) + ((!shiftx4x) & (shiftx5x) & (g266) & (g267) & (!g268) & (g269)) + ((!shiftx4x) & (shiftx5x) & (g266) & (g267) & (g268) & (!g269)) + ((!shiftx4x) & (shiftx5x) & (g266) & (g267) & (g268) & (g269)) + ((shiftx4x) & (!shiftx5x) & (!g266) & (!g267) & (!g268) & (g269)) + ((shiftx4x) & (!shiftx5x) & (!g266) & (!g267) & (g268) & (g269)) + ((shiftx4x) & (!shiftx5x) & (!g266) & (g267) & (!g268) & (g269)) + ((shiftx4x) & (!shiftx5x) & (!g266) & (g267) & (g268) & (g269)) + ((shiftx4x) & (!shiftx5x) & (g266) & (!g267) & (!g268) & (g269)) + ((shiftx4x) & (!shiftx5x) & (g266) & (!g267) & (g268) & (g269)) + ((shiftx4x) & (!shiftx5x) & (g266) & (g267) & (!g268) & (g269)) + ((shiftx4x) & (!shiftx5x) & (g266) & (g267) & (g268) & (g269)) + ((shiftx4x) & (shiftx5x) & (g266) & (!g267) & (!g268) & (!g269)) + ((shiftx4x) & (shiftx5x) & (g266) & (!g267) & (!g268) & (g269)) + ((shiftx4x) & (shiftx5x) & (g266) & (!g267) & (g268) & (!g269)) + ((shiftx4x) & (shiftx5x) & (g266) & (!g267) & (g268) & (g269)) + ((shiftx4x) & (shiftx5x) & (g266) & (g267) & (!g268) & (!g269)) + ((shiftx4x) & (shiftx5x) & (g266) & (g267) & (!g268) & (g269)) + ((shiftx4x) & (shiftx5x) & (g266) & (g267) & (g268) & (!g269)) + ((shiftx4x) & (shiftx5x) & (g266) & (g267) & (g268) & (g269)));
	assign resultx12x = (((!shiftx6x) & (!g265) & (sk[14]) & (g270)) + ((!shiftx6x) & (g265) & (sk[14]) & (g270)) + ((shiftx6x) & (!g265) & (!sk[14]) & (!g270)) + ((shiftx6x) & (!g265) & (!sk[14]) & (g270)) + ((shiftx6x) & (g265) & (!sk[14]) & (!g270)) + ((shiftx6x) & (g265) & (!sk[14]) & (g270)) + ((shiftx6x) & (g265) & (sk[14]) & (!g270)) + ((shiftx6x) & (g265) & (sk[14]) & (g270)));
	assign g272 = (((!shiftx2x) & (!shiftx3x) & (g45) & (!g46) & (!g47) & (!g54)) + ((!shiftx2x) & (!shiftx3x) & (g45) & (!g46) & (!g47) & (g54)) + ((!shiftx2x) & (!shiftx3x) & (g45) & (!g46) & (g47) & (!g54)) + ((!shiftx2x) & (!shiftx3x) & (g45) & (!g46) & (g47) & (g54)) + ((!shiftx2x) & (!shiftx3x) & (g45) & (g46) & (!g47) & (!g54)) + ((!shiftx2x) & (!shiftx3x) & (g45) & (g46) & (!g47) & (g54)) + ((!shiftx2x) & (!shiftx3x) & (g45) & (g46) & (g47) & (!g54)) + ((!shiftx2x) & (!shiftx3x) & (g45) & (g46) & (g47) & (g54)) + ((!shiftx2x) & (shiftx3x) & (!g45) & (g46) & (!g47) & (!g54)) + ((!shiftx2x) & (shiftx3x) & (!g45) & (g46) & (!g47) & (g54)) + ((!shiftx2x) & (shiftx3x) & (!g45) & (g46) & (g47) & (!g54)) + ((!shiftx2x) & (shiftx3x) & (!g45) & (g46) & (g47) & (g54)) + ((!shiftx2x) & (shiftx3x) & (g45) & (g46) & (!g47) & (!g54)) + ((!shiftx2x) & (shiftx3x) & (g45) & (g46) & (!g47) & (g54)) + ((!shiftx2x) & (shiftx3x) & (g45) & (g46) & (g47) & (!g54)) + ((!shiftx2x) & (shiftx3x) & (g45) & (g46) & (g47) & (g54)) + ((shiftx2x) & (!shiftx3x) & (!g45) & (!g46) & (g47) & (!g54)) + ((shiftx2x) & (!shiftx3x) & (!g45) & (!g46) & (g47) & (g54)) + ((shiftx2x) & (!shiftx3x) & (!g45) & (g46) & (g47) & (!g54)) + ((shiftx2x) & (!shiftx3x) & (!g45) & (g46) & (g47) & (g54)) + ((shiftx2x) & (!shiftx3x) & (g45) & (!g46) & (g47) & (!g54)) + ((shiftx2x) & (!shiftx3x) & (g45) & (!g46) & (g47) & (g54)) + ((shiftx2x) & (!shiftx3x) & (g45) & (g46) & (g47) & (!g54)) + ((shiftx2x) & (!shiftx3x) & (g45) & (g46) & (g47) & (g54)) + ((shiftx2x) & (shiftx3x) & (!g45) & (!g46) & (!g47) & (g54)) + ((shiftx2x) & (shiftx3x) & (!g45) & (!g46) & (g47) & (g54)) + ((shiftx2x) & (shiftx3x) & (!g45) & (g46) & (!g47) & (g54)) + ((shiftx2x) & (shiftx3x) & (!g45) & (g46) & (g47) & (g54)) + ((shiftx2x) & (shiftx3x) & (g45) & (!g46) & (!g47) & (g54)) + ((shiftx2x) & (shiftx3x) & (g45) & (!g46) & (g47) & (g54)) + ((shiftx2x) & (shiftx3x) & (g45) & (g46) & (!g47) & (g54)) + ((shiftx2x) & (shiftx3x) & (g45) & (g46) & (g47) & (g54)));
	assign g273 = (((!shiftx2x) & (!shiftx3x) & (!g44) & (g66) & (!g67) & (!g68)) + ((!shiftx2x) & (!shiftx3x) & (!g44) & (g66) & (!g67) & (g68)) + ((!shiftx2x) & (!shiftx3x) & (!g44) & (g66) & (g67) & (!g68)) + ((!shiftx2x) & (!shiftx3x) & (!g44) & (g66) & (g67) & (g68)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (g66) & (!g67) & (!g68)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (g66) & (!g67) & (g68)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (g66) & (g67) & (!g68)) + ((!shiftx2x) & (!shiftx3x) & (g44) & (g66) & (g67) & (g68)) + ((!shiftx2x) & (shiftx3x) & (!g44) & (!g66) & (g67) & (!g68)) + ((!shiftx2x) & (shiftx3x) & (!g44) & (!g66) & (g67) & (g68)) + ((!shiftx2x) & (shiftx3x) & (!g44) & (g66) & (g67) & (!g68)) + ((!shiftx2x) & (shiftx3x) & (!g44) & (g66) & (g67) & (g68)) + ((!shiftx2x) & (shiftx3x) & (g44) & (!g66) & (g67) & (!g68)) + ((!shiftx2x) & (shiftx3x) & (g44) & (!g66) & (g67) & (g68)) + ((!shiftx2x) & (shiftx3x) & (g44) & (g66) & (g67) & (!g68)) + ((!shiftx2x) & (shiftx3x) & (g44) & (g66) & (g67) & (g68)) + ((shiftx2x) & (!shiftx3x) & (!g44) & (!g66) & (!g67) & (g68)) + ((shiftx2x) & (!shiftx3x) & (!g44) & (!g66) & (g67) & (g68)) + ((shiftx2x) & (!shiftx3x) & (!g44) & (g66) & (!g67) & (g68)) + ((shiftx2x) & (!shiftx3x) & (!g44) & (g66) & (g67) & (g68)) + ((shiftx2x) & (!shiftx3x) & (g44) & (!g66) & (!g67) & (g68)) + ((shiftx2x) & (!shiftx3x) & (g44) & (!g66) & (g67) & (g68)) + ((shiftx2x) & (!shiftx3x) & (g44) & (g66) & (!g67) & (g68)) + ((shiftx2x) & (!shiftx3x) & (g44) & (g66) & (g67) & (g68)) + ((shiftx2x) & (shiftx3x) & (g44) & (!g66) & (!g67) & (!g68)) + ((shiftx2x) & (shiftx3x) & (g44) & (!g66) & (!g67) & (g68)) + ((shiftx2x) & (shiftx3x) & (g44) & (!g66) & (g67) & (!g68)) + ((shiftx2x) & (shiftx3x) & (g44) & (!g66) & (g67) & (g68)) + ((shiftx2x) & (shiftx3x) & (g44) & (g66) & (!g67) & (!g68)) + ((shiftx2x) & (shiftx3x) & (g44) & (g66) & (!g67) & (g68)) + ((shiftx2x) & (shiftx3x) & (g44) & (g66) & (g67) & (!g68)) + ((shiftx2x) & (shiftx3x) & (g44) & (g66) & (g67) & (g68)));
	assign g274 = (((!shiftx2x) & (!shiftx3x) & (g55) & (!g56) & (!g57) & (!g59)) + ((!shiftx2x) & (!shiftx3x) & (g55) & (!g56) & (!g57) & (g59)) + ((!shiftx2x) & (!shiftx3x) & (g55) & (!g56) & (g57) & (!g59)) + ((!shiftx2x) & (!shiftx3x) & (g55) & (!g56) & (g57) & (g59)) + ((!shiftx2x) & (!shiftx3x) & (g55) & (g56) & (!g57) & (!g59)) + ((!shiftx2x) & (!shiftx3x) & (g55) & (g56) & (!g57) & (g59)) + ((!shiftx2x) & (!shiftx3x) & (g55) & (g56) & (g57) & (!g59)) + ((!shiftx2x) & (!shiftx3x) & (g55) & (g56) & (g57) & (g59)) + ((!shiftx2x) & (shiftx3x) & (!g55) & (g56) & (!g57) & (!g59)) + ((!shiftx2x) & (shiftx3x) & (!g55) & (g56) & (!g57) & (g59)) + ((!shiftx2x) & (shiftx3x) & (!g55) & (g56) & (g57) & (!g59)) + ((!shiftx2x) & (shiftx3x) & (!g55) & (g56) & (g57) & (g59)) + ((!shiftx2x) & (shiftx3x) & (g55) & (g56) & (!g57) & (!g59)) + ((!shiftx2x) & (shiftx3x) & (g55) & (g56) & (!g57) & (g59)) + ((!shiftx2x) & (shiftx3x) & (g55) & (g56) & (g57) & (!g59)) + ((!shiftx2x) & (shiftx3x) & (g55) & (g56) & (g57) & (g59)) + ((shiftx2x) & (!shiftx3x) & (!g55) & (!g56) & (g57) & (!g59)) + ((shiftx2x) & (!shiftx3x) & (!g55) & (!g56) & (g57) & (g59)) + ((shiftx2x) & (!shiftx3x) & (!g55) & (g56) & (g57) & (!g59)) + ((shiftx2x) & (!shiftx3x) & (!g55) & (g56) & (g57) & (g59)) + ((shiftx2x) & (!shiftx3x) & (g55) & (!g56) & (g57) & (!g59)) + ((shiftx2x) & (!shiftx3x) & (g55) & (!g56) & (g57) & (g59)) + ((shiftx2x) & (!shiftx3x) & (g55) & (g56) & (g57) & (!g59)) + ((shiftx2x) & (!shiftx3x) & (g55) & (g56) & (g57) & (g59)) + ((shiftx2x) & (shiftx3x) & (!g55) & (!g56) & (!g57) & (g59)) + ((shiftx2x) & (shiftx3x) & (!g55) & (!g56) & (g57) & (g59)) + ((shiftx2x) & (shiftx3x) & (!g55) & (g56) & (!g57) & (g59)) + ((shiftx2x) & (shiftx3x) & (!g55) & (g56) & (g57) & (g59)) + ((shiftx2x) & (shiftx3x) & (g55) & (!g56) & (!g57) & (g59)) + ((shiftx2x) & (shiftx3x) & (g55) & (!g56) & (g57) & (g59)) + ((shiftx2x) & (shiftx3x) & (g55) & (g56) & (!g57) & (g59)) + ((shiftx2x) & (shiftx3x) & (g55) & (g56) & (g57) & (g59)));
	assign g275 = (((!shiftx2x) & (!shiftx3x) & (!g49) & (g60) & (!g61) & (!g62)) + ((!shiftx2x) & (!shiftx3x) & (!g49) & (g60) & (!g61) & (g62)) + ((!shiftx2x) & (!shiftx3x) & (!g49) & (g60) & (g61) & (!g62)) + ((!shiftx2x) & (!shiftx3x) & (!g49) & (g60) & (g61) & (g62)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (g60) & (!g61) & (!g62)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (g60) & (!g61) & (g62)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (g60) & (g61) & (!g62)) + ((!shiftx2x) & (!shiftx3x) & (g49) & (g60) & (g61) & (g62)) + ((!shiftx2x) & (shiftx3x) & (!g49) & (!g60) & (g61) & (!g62)) + ((!shiftx2x) & (shiftx3x) & (!g49) & (!g60) & (g61) & (g62)) + ((!shiftx2x) & (shiftx3x) & (!g49) & (g60) & (g61) & (!g62)) + ((!shiftx2x) & (shiftx3x) & (!g49) & (g60) & (g61) & (g62)) + ((!shiftx2x) & (shiftx3x) & (g49) & (!g60) & (g61) & (!g62)) + ((!shiftx2x) & (shiftx3x) & (g49) & (!g60) & (g61) & (g62)) + ((!shiftx2x) & (shiftx3x) & (g49) & (g60) & (g61) & (!g62)) + ((!shiftx2x) & (shiftx3x) & (g49) & (g60) & (g61) & (g62)) + ((shiftx2x) & (!shiftx3x) & (!g49) & (!g60) & (!g61) & (g62)) + ((shiftx2x) & (!shiftx3x) & (!g49) & (!g60) & (g61) & (g62)) + ((shiftx2x) & (!shiftx3x) & (!g49) & (g60) & (!g61) & (g62)) + ((shiftx2x) & (!shiftx3x) & (!g49) & (g60) & (g61) & (g62)) + ((shiftx2x) & (!shiftx3x) & (g49) & (!g60) & (!g61) & (g62)) + ((shiftx2x) & (!shiftx3x) & (g49) & (!g60) & (g61) & (g62)) + ((shiftx2x) & (!shiftx3x) & (g49) & (g60) & (!g61) & (g62)) + ((shiftx2x) & (!shiftx3x) & (g49) & (g60) & (g61) & (g62)) + ((shiftx2x) & (shiftx3x) & (g49) & (!g60) & (!g61) & (!g62)) + ((shiftx2x) & (shiftx3x) & (g49) & (!g60) & (!g61) & (g62)) + ((shiftx2x) & (shiftx3x) & (g49) & (!g60) & (g61) & (!g62)) + ((shiftx2x) & (shiftx3x) & (g49) & (!g60) & (g61) & (g62)) + ((shiftx2x) & (shiftx3x) & (g49) & (g60) & (!g61) & (!g62)) + ((shiftx2x) & (shiftx3x) & (g49) & (g60) & (!g61) & (g62)) + ((shiftx2x) & (shiftx3x) & (g49) & (g60) & (g61) & (!g62)) + ((shiftx2x) & (shiftx3x) & (g49) & (g60) & (g61) & (g62)));
	assign g276 = (((!shiftx4x) & (!shiftx5x) & (!g272) & (g273) & (!g274) & (!g275)) + ((!shiftx4x) & (!shiftx5x) & (!g272) & (g273) & (!g274) & (g275)) + ((!shiftx4x) & (!shiftx5x) & (!g272) & (g273) & (g274) & (!g275)) + ((!shiftx4x) & (!shiftx5x) & (!g272) & (g273) & (g274) & (g275)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (g273) & (!g274) & (!g275)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (g273) & (!g274) & (g275)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (g273) & (g274) & (!g275)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (g273) & (g274) & (g275)) + ((!shiftx4x) & (shiftx5x) & (!g272) & (!g273) & (g274) & (!g275)) + ((!shiftx4x) & (shiftx5x) & (!g272) & (!g273) & (g274) & (g275)) + ((!shiftx4x) & (shiftx5x) & (!g272) & (g273) & (g274) & (!g275)) + ((!shiftx4x) & (shiftx5x) & (!g272) & (g273) & (g274) & (g275)) + ((!shiftx4x) & (shiftx5x) & (g272) & (!g273) & (g274) & (!g275)) + ((!shiftx4x) & (shiftx5x) & (g272) & (!g273) & (g274) & (g275)) + ((!shiftx4x) & (shiftx5x) & (g272) & (g273) & (g274) & (!g275)) + ((!shiftx4x) & (shiftx5x) & (g272) & (g273) & (g274) & (g275)) + ((shiftx4x) & (!shiftx5x) & (g272) & (!g273) & (!g274) & (!g275)) + ((shiftx4x) & (!shiftx5x) & (g272) & (!g273) & (!g274) & (g275)) + ((shiftx4x) & (!shiftx5x) & (g272) & (!g273) & (g274) & (!g275)) + ((shiftx4x) & (!shiftx5x) & (g272) & (!g273) & (g274) & (g275)) + ((shiftx4x) & (!shiftx5x) & (g272) & (g273) & (!g274) & (!g275)) + ((shiftx4x) & (!shiftx5x) & (g272) & (g273) & (!g274) & (g275)) + ((shiftx4x) & (!shiftx5x) & (g272) & (g273) & (g274) & (!g275)) + ((shiftx4x) & (!shiftx5x) & (g272) & (g273) & (g274) & (g275)) + ((shiftx4x) & (shiftx5x) & (!g272) & (!g273) & (!g274) & (g275)) + ((shiftx4x) & (shiftx5x) & (!g272) & (!g273) & (g274) & (g275)) + ((shiftx4x) & (shiftx5x) & (!g272) & (g273) & (!g274) & (g275)) + ((shiftx4x) & (shiftx5x) & (!g272) & (g273) & (g274) & (g275)) + ((shiftx4x) & (shiftx5x) & (g272) & (!g273) & (!g274) & (g275)) + ((shiftx4x) & (shiftx5x) & (g272) & (!g273) & (g274) & (g275)) + ((shiftx4x) & (shiftx5x) & (g272) & (g273) & (!g274) & (g275)) + ((shiftx4x) & (shiftx5x) & (g272) & (g273) & (g274) & (g275)));
	assign g277 = (((!shiftx2x) & (!shiftx3x) & (!g65) & (g71) & (!g72) & (!g73)) + ((!shiftx2x) & (!shiftx3x) & (!g65) & (g71) & (!g72) & (g73)) + ((!shiftx2x) & (!shiftx3x) & (!g65) & (g71) & (g72) & (!g73)) + ((!shiftx2x) & (!shiftx3x) & (!g65) & (g71) & (g72) & (g73)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (g71) & (!g72) & (!g73)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (g71) & (!g72) & (g73)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (g71) & (g72) & (!g73)) + ((!shiftx2x) & (!shiftx3x) & (g65) & (g71) & (g72) & (g73)) + ((!shiftx2x) & (shiftx3x) & (!g65) & (!g71) & (g72) & (!g73)) + ((!shiftx2x) & (shiftx3x) & (!g65) & (!g71) & (g72) & (g73)) + ((!shiftx2x) & (shiftx3x) & (!g65) & (g71) & (g72) & (!g73)) + ((!shiftx2x) & (shiftx3x) & (!g65) & (g71) & (g72) & (g73)) + ((!shiftx2x) & (shiftx3x) & (g65) & (!g71) & (g72) & (!g73)) + ((!shiftx2x) & (shiftx3x) & (g65) & (!g71) & (g72) & (g73)) + ((!shiftx2x) & (shiftx3x) & (g65) & (g71) & (g72) & (!g73)) + ((!shiftx2x) & (shiftx3x) & (g65) & (g71) & (g72) & (g73)) + ((shiftx2x) & (!shiftx3x) & (!g65) & (!g71) & (!g72) & (g73)) + ((shiftx2x) & (!shiftx3x) & (!g65) & (!g71) & (g72) & (g73)) + ((shiftx2x) & (!shiftx3x) & (!g65) & (g71) & (!g72) & (g73)) + ((shiftx2x) & (!shiftx3x) & (!g65) & (g71) & (g72) & (g73)) + ((shiftx2x) & (!shiftx3x) & (g65) & (!g71) & (!g72) & (g73)) + ((shiftx2x) & (!shiftx3x) & (g65) & (!g71) & (g72) & (g73)) + ((shiftx2x) & (!shiftx3x) & (g65) & (g71) & (!g72) & (g73)) + ((shiftx2x) & (!shiftx3x) & (g65) & (g71) & (g72) & (g73)) + ((shiftx2x) & (shiftx3x) & (g65) & (!g71) & (!g72) & (!g73)) + ((shiftx2x) & (shiftx3x) & (g65) & (!g71) & (!g72) & (g73)) + ((shiftx2x) & (shiftx3x) & (g65) & (!g71) & (g72) & (!g73)) + ((shiftx2x) & (shiftx3x) & (g65) & (!g71) & (g72) & (g73)) + ((shiftx2x) & (shiftx3x) & (g65) & (g71) & (!g72) & (!g73)) + ((shiftx2x) & (shiftx3x) & (g65) & (g71) & (!g72) & (g73)) + ((shiftx2x) & (shiftx3x) & (g65) & (g71) & (g72) & (!g73)) + ((shiftx2x) & (shiftx3x) & (g65) & (g71) & (g72) & (g73)));
	assign g278 = (((!shiftx2x) & (!shiftx3x) & (!g70) & (g81) & (!g82) & (!g83)) + ((!shiftx2x) & (!shiftx3x) & (!g70) & (g81) & (!g82) & (g83)) + ((!shiftx2x) & (!shiftx3x) & (!g70) & (g81) & (g82) & (!g83)) + ((!shiftx2x) & (!shiftx3x) & (!g70) & (g81) & (g82) & (g83)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (g81) & (!g82) & (!g83)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (g81) & (!g82) & (g83)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (g81) & (g82) & (!g83)) + ((!shiftx2x) & (!shiftx3x) & (g70) & (g81) & (g82) & (g83)) + ((!shiftx2x) & (shiftx3x) & (!g70) & (!g81) & (g82) & (!g83)) + ((!shiftx2x) & (shiftx3x) & (!g70) & (!g81) & (g82) & (g83)) + ((!shiftx2x) & (shiftx3x) & (!g70) & (g81) & (g82) & (!g83)) + ((!shiftx2x) & (shiftx3x) & (!g70) & (g81) & (g82) & (g83)) + ((!shiftx2x) & (shiftx3x) & (g70) & (!g81) & (g82) & (!g83)) + ((!shiftx2x) & (shiftx3x) & (g70) & (!g81) & (g82) & (g83)) + ((!shiftx2x) & (shiftx3x) & (g70) & (g81) & (g82) & (!g83)) + ((!shiftx2x) & (shiftx3x) & (g70) & (g81) & (g82) & (g83)) + ((shiftx2x) & (!shiftx3x) & (!g70) & (!g81) & (!g82) & (g83)) + ((shiftx2x) & (!shiftx3x) & (!g70) & (!g81) & (g82) & (g83)) + ((shiftx2x) & (!shiftx3x) & (!g70) & (g81) & (!g82) & (g83)) + ((shiftx2x) & (!shiftx3x) & (!g70) & (g81) & (g82) & (g83)) + ((shiftx2x) & (!shiftx3x) & (g70) & (!g81) & (!g82) & (g83)) + ((shiftx2x) & (!shiftx3x) & (g70) & (!g81) & (g82) & (g83)) + ((shiftx2x) & (!shiftx3x) & (g70) & (g81) & (!g82) & (g83)) + ((shiftx2x) & (!shiftx3x) & (g70) & (g81) & (g82) & (g83)) + ((shiftx2x) & (shiftx3x) & (g70) & (!g81) & (!g82) & (!g83)) + ((shiftx2x) & (shiftx3x) & (g70) & (!g81) & (!g82) & (g83)) + ((shiftx2x) & (shiftx3x) & (g70) & (!g81) & (g82) & (!g83)) + ((shiftx2x) & (shiftx3x) & (g70) & (!g81) & (g82) & (g83)) + ((shiftx2x) & (shiftx3x) & (g70) & (g81) & (!g82) & (!g83)) + ((shiftx2x) & (shiftx3x) & (g70) & (g81) & (!g82) & (g83)) + ((shiftx2x) & (shiftx3x) & (g70) & (g81) & (g82) & (!g83)) + ((shiftx2x) & (shiftx3x) & (g70) & (g81) & (g82) & (g83)));
	assign g279 = (((!shiftx2x) & (!shiftx3x) & (g50) & (!g51) & (!g52) & (!g75)) + ((!shiftx2x) & (!shiftx3x) & (g50) & (!g51) & (!g52) & (g75)) + ((!shiftx2x) & (!shiftx3x) & (g50) & (!g51) & (g52) & (!g75)) + ((!shiftx2x) & (!shiftx3x) & (g50) & (!g51) & (g52) & (g75)) + ((!shiftx2x) & (!shiftx3x) & (g50) & (g51) & (!g52) & (!g75)) + ((!shiftx2x) & (!shiftx3x) & (g50) & (g51) & (!g52) & (g75)) + ((!shiftx2x) & (!shiftx3x) & (g50) & (g51) & (g52) & (!g75)) + ((!shiftx2x) & (!shiftx3x) & (g50) & (g51) & (g52) & (g75)) + ((!shiftx2x) & (shiftx3x) & (!g50) & (g51) & (!g52) & (!g75)) + ((!shiftx2x) & (shiftx3x) & (!g50) & (g51) & (!g52) & (g75)) + ((!shiftx2x) & (shiftx3x) & (!g50) & (g51) & (g52) & (!g75)) + ((!shiftx2x) & (shiftx3x) & (!g50) & (g51) & (g52) & (g75)) + ((!shiftx2x) & (shiftx3x) & (g50) & (g51) & (!g52) & (!g75)) + ((!shiftx2x) & (shiftx3x) & (g50) & (g51) & (!g52) & (g75)) + ((!shiftx2x) & (shiftx3x) & (g50) & (g51) & (g52) & (!g75)) + ((!shiftx2x) & (shiftx3x) & (g50) & (g51) & (g52) & (g75)) + ((shiftx2x) & (!shiftx3x) & (!g50) & (!g51) & (g52) & (!g75)) + ((shiftx2x) & (!shiftx3x) & (!g50) & (!g51) & (g52) & (g75)) + ((shiftx2x) & (!shiftx3x) & (!g50) & (g51) & (g52) & (!g75)) + ((shiftx2x) & (!shiftx3x) & (!g50) & (g51) & (g52) & (g75)) + ((shiftx2x) & (!shiftx3x) & (g50) & (!g51) & (g52) & (!g75)) + ((shiftx2x) & (!shiftx3x) & (g50) & (!g51) & (g52) & (g75)) + ((shiftx2x) & (!shiftx3x) & (g50) & (g51) & (g52) & (!g75)) + ((shiftx2x) & (!shiftx3x) & (g50) & (g51) & (g52) & (g75)) + ((shiftx2x) & (shiftx3x) & (!g50) & (!g51) & (!g52) & (g75)) + ((shiftx2x) & (shiftx3x) & (!g50) & (!g51) & (g52) & (g75)) + ((shiftx2x) & (shiftx3x) & (!g50) & (g51) & (!g52) & (g75)) + ((shiftx2x) & (shiftx3x) & (!g50) & (g51) & (g52) & (g75)) + ((shiftx2x) & (shiftx3x) & (g50) & (!g51) & (!g52) & (g75)) + ((shiftx2x) & (shiftx3x) & (g50) & (!g51) & (g52) & (g75)) + ((shiftx2x) & (shiftx3x) & (g50) & (g51) & (!g52) & (g75)) + ((shiftx2x) & (shiftx3x) & (g50) & (g51) & (g52) & (g75)));
	assign g280 = (((!shiftx2x) & (!shiftx3x) & (g76) & (!g77) & (!g78) & (!g80)) + ((!shiftx2x) & (!shiftx3x) & (g76) & (!g77) & (!g78) & (g80)) + ((!shiftx2x) & (!shiftx3x) & (g76) & (!g77) & (g78) & (!g80)) + ((!shiftx2x) & (!shiftx3x) & (g76) & (!g77) & (g78) & (g80)) + ((!shiftx2x) & (!shiftx3x) & (g76) & (g77) & (!g78) & (!g80)) + ((!shiftx2x) & (!shiftx3x) & (g76) & (g77) & (!g78) & (g80)) + ((!shiftx2x) & (!shiftx3x) & (g76) & (g77) & (g78) & (!g80)) + ((!shiftx2x) & (!shiftx3x) & (g76) & (g77) & (g78) & (g80)) + ((!shiftx2x) & (shiftx3x) & (!g76) & (g77) & (!g78) & (!g80)) + ((!shiftx2x) & (shiftx3x) & (!g76) & (g77) & (!g78) & (g80)) + ((!shiftx2x) & (shiftx3x) & (!g76) & (g77) & (g78) & (!g80)) + ((!shiftx2x) & (shiftx3x) & (!g76) & (g77) & (g78) & (g80)) + ((!shiftx2x) & (shiftx3x) & (g76) & (g77) & (!g78) & (!g80)) + ((!shiftx2x) & (shiftx3x) & (g76) & (g77) & (!g78) & (g80)) + ((!shiftx2x) & (shiftx3x) & (g76) & (g77) & (g78) & (!g80)) + ((!shiftx2x) & (shiftx3x) & (g76) & (g77) & (g78) & (g80)) + ((shiftx2x) & (!shiftx3x) & (!g76) & (!g77) & (g78) & (!g80)) + ((shiftx2x) & (!shiftx3x) & (!g76) & (!g77) & (g78) & (g80)) + ((shiftx2x) & (!shiftx3x) & (!g76) & (g77) & (g78) & (!g80)) + ((shiftx2x) & (!shiftx3x) & (!g76) & (g77) & (g78) & (g80)) + ((shiftx2x) & (!shiftx3x) & (g76) & (!g77) & (g78) & (!g80)) + ((shiftx2x) & (!shiftx3x) & (g76) & (!g77) & (g78) & (g80)) + ((shiftx2x) & (!shiftx3x) & (g76) & (g77) & (g78) & (!g80)) + ((shiftx2x) & (!shiftx3x) & (g76) & (g77) & (g78) & (g80)) + ((shiftx2x) & (shiftx3x) & (!g76) & (!g77) & (!g78) & (g80)) + ((shiftx2x) & (shiftx3x) & (!g76) & (!g77) & (g78) & (g80)) + ((shiftx2x) & (shiftx3x) & (!g76) & (g77) & (!g78) & (g80)) + ((shiftx2x) & (shiftx3x) & (!g76) & (g77) & (g78) & (g80)) + ((shiftx2x) & (shiftx3x) & (g76) & (!g77) & (!g78) & (g80)) + ((shiftx2x) & (shiftx3x) & (g76) & (!g77) & (g78) & (g80)) + ((shiftx2x) & (shiftx3x) & (g76) & (g77) & (!g78) & (g80)) + ((shiftx2x) & (shiftx3x) & (g76) & (g77) & (g78) & (g80)));
	assign g281 = (((!shiftx4x) & (!shiftx5x) & (!g277) & (!g278) & (g279) & (!g280)) + ((!shiftx4x) & (!shiftx5x) & (!g277) & (!g278) & (g279) & (g280)) + ((!shiftx4x) & (!shiftx5x) & (!g277) & (g278) & (g279) & (!g280)) + ((!shiftx4x) & (!shiftx5x) & (!g277) & (g278) & (g279) & (g280)) + ((!shiftx4x) & (!shiftx5x) & (g277) & (!g278) & (g279) & (!g280)) + ((!shiftx4x) & (!shiftx5x) & (g277) & (!g278) & (g279) & (g280)) + ((!shiftx4x) & (!shiftx5x) & (g277) & (g278) & (g279) & (!g280)) + ((!shiftx4x) & (!shiftx5x) & (g277) & (g278) & (g279) & (g280)) + ((!shiftx4x) & (shiftx5x) & (!g277) & (g278) & (!g279) & (!g280)) + ((!shiftx4x) & (shiftx5x) & (!g277) & (g278) & (!g279) & (g280)) + ((!shiftx4x) & (shiftx5x) & (!g277) & (g278) & (g279) & (!g280)) + ((!shiftx4x) & (shiftx5x) & (!g277) & (g278) & (g279) & (g280)) + ((!shiftx4x) & (shiftx5x) & (g277) & (g278) & (!g279) & (!g280)) + ((!shiftx4x) & (shiftx5x) & (g277) & (g278) & (!g279) & (g280)) + ((!shiftx4x) & (shiftx5x) & (g277) & (g278) & (g279) & (!g280)) + ((!shiftx4x) & (shiftx5x) & (g277) & (g278) & (g279) & (g280)) + ((shiftx4x) & (!shiftx5x) & (!g277) & (!g278) & (!g279) & (g280)) + ((shiftx4x) & (!shiftx5x) & (!g277) & (!g278) & (g279) & (g280)) + ((shiftx4x) & (!shiftx5x) & (!g277) & (g278) & (!g279) & (g280)) + ((shiftx4x) & (!shiftx5x) & (!g277) & (g278) & (g279) & (g280)) + ((shiftx4x) & (!shiftx5x) & (g277) & (!g278) & (!g279) & (g280)) + ((shiftx4x) & (!shiftx5x) & (g277) & (!g278) & (g279) & (g280)) + ((shiftx4x) & (!shiftx5x) & (g277) & (g278) & (!g279) & (g280)) + ((shiftx4x) & (!shiftx5x) & (g277) & (g278) & (g279) & (g280)) + ((shiftx4x) & (shiftx5x) & (g277) & (!g278) & (!g279) & (!g280)) + ((shiftx4x) & (shiftx5x) & (g277) & (!g278) & (!g279) & (g280)) + ((shiftx4x) & (shiftx5x) & (g277) & (!g278) & (g279) & (!g280)) + ((shiftx4x) & (shiftx5x) & (g277) & (!g278) & (g279) & (g280)) + ((shiftx4x) & (shiftx5x) & (g277) & (g278) & (!g279) & (!g280)) + ((shiftx4x) & (shiftx5x) & (g277) & (g278) & (!g279) & (g280)) + ((shiftx4x) & (shiftx5x) & (g277) & (g278) & (g279) & (!g280)) + ((shiftx4x) & (shiftx5x) & (g277) & (g278) & (g279) & (g280)));
	assign resultx13x = (((!shiftx6x) & (!g276) & (sk[25]) & (g281)) + ((!shiftx6x) & (g276) & (sk[25]) & (g281)) + ((shiftx6x) & (!g276) & (!sk[25]) & (!g281)) + ((shiftx6x) & (!g276) & (!sk[25]) & (g281)) + ((shiftx6x) & (g276) & (!sk[25]) & (!g281)) + ((shiftx6x) & (g276) & (!sk[25]) & (g281)) + ((shiftx6x) & (g276) & (sk[25]) & (!g281)) + ((shiftx6x) & (g276) & (sk[25]) & (g281)));
	assign g283 = (((!shiftx2x) & (!shiftx3x) & (g88) & (!g89) & (!g90) & (!g97)) + ((!shiftx2x) & (!shiftx3x) & (g88) & (!g89) & (!g90) & (g97)) + ((!shiftx2x) & (!shiftx3x) & (g88) & (!g89) & (g90) & (!g97)) + ((!shiftx2x) & (!shiftx3x) & (g88) & (!g89) & (g90) & (g97)) + ((!shiftx2x) & (!shiftx3x) & (g88) & (g89) & (!g90) & (!g97)) + ((!shiftx2x) & (!shiftx3x) & (g88) & (g89) & (!g90) & (g97)) + ((!shiftx2x) & (!shiftx3x) & (g88) & (g89) & (g90) & (!g97)) + ((!shiftx2x) & (!shiftx3x) & (g88) & (g89) & (g90) & (g97)) + ((!shiftx2x) & (shiftx3x) & (!g88) & (g89) & (!g90) & (!g97)) + ((!shiftx2x) & (shiftx3x) & (!g88) & (g89) & (!g90) & (g97)) + ((!shiftx2x) & (shiftx3x) & (!g88) & (g89) & (g90) & (!g97)) + ((!shiftx2x) & (shiftx3x) & (!g88) & (g89) & (g90) & (g97)) + ((!shiftx2x) & (shiftx3x) & (g88) & (g89) & (!g90) & (!g97)) + ((!shiftx2x) & (shiftx3x) & (g88) & (g89) & (!g90) & (g97)) + ((!shiftx2x) & (shiftx3x) & (g88) & (g89) & (g90) & (!g97)) + ((!shiftx2x) & (shiftx3x) & (g88) & (g89) & (g90) & (g97)) + ((shiftx2x) & (!shiftx3x) & (!g88) & (!g89) & (g90) & (!g97)) + ((shiftx2x) & (!shiftx3x) & (!g88) & (!g89) & (g90) & (g97)) + ((shiftx2x) & (!shiftx3x) & (!g88) & (g89) & (g90) & (!g97)) + ((shiftx2x) & (!shiftx3x) & (!g88) & (g89) & (g90) & (g97)) + ((shiftx2x) & (!shiftx3x) & (g88) & (!g89) & (g90) & (!g97)) + ((shiftx2x) & (!shiftx3x) & (g88) & (!g89) & (g90) & (g97)) + ((shiftx2x) & (!shiftx3x) & (g88) & (g89) & (g90) & (!g97)) + ((shiftx2x) & (!shiftx3x) & (g88) & (g89) & (g90) & (g97)) + ((shiftx2x) & (shiftx3x) & (!g88) & (!g89) & (!g90) & (g97)) + ((shiftx2x) & (shiftx3x) & (!g88) & (!g89) & (g90) & (g97)) + ((shiftx2x) & (shiftx3x) & (!g88) & (g89) & (!g90) & (g97)) + ((shiftx2x) & (shiftx3x) & (!g88) & (g89) & (g90) & (g97)) + ((shiftx2x) & (shiftx3x) & (g88) & (!g89) & (!g90) & (g97)) + ((shiftx2x) & (shiftx3x) & (g88) & (!g89) & (g90) & (g97)) + ((shiftx2x) & (shiftx3x) & (g88) & (g89) & (!g90) & (g97)) + ((shiftx2x) & (shiftx3x) & (g88) & (g89) & (g90) & (g97)));
	assign g284 = (((!shiftx2x) & (!shiftx3x) & (!g87) & (g109) & (!g110) & (!g111)) + ((!shiftx2x) & (!shiftx3x) & (!g87) & (g109) & (!g110) & (g111)) + ((!shiftx2x) & (!shiftx3x) & (!g87) & (g109) & (g110) & (!g111)) + ((!shiftx2x) & (!shiftx3x) & (!g87) & (g109) & (g110) & (g111)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (g109) & (!g110) & (!g111)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (g109) & (!g110) & (g111)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (g109) & (g110) & (!g111)) + ((!shiftx2x) & (!shiftx3x) & (g87) & (g109) & (g110) & (g111)) + ((!shiftx2x) & (shiftx3x) & (!g87) & (!g109) & (g110) & (!g111)) + ((!shiftx2x) & (shiftx3x) & (!g87) & (!g109) & (g110) & (g111)) + ((!shiftx2x) & (shiftx3x) & (!g87) & (g109) & (g110) & (!g111)) + ((!shiftx2x) & (shiftx3x) & (!g87) & (g109) & (g110) & (g111)) + ((!shiftx2x) & (shiftx3x) & (g87) & (!g109) & (g110) & (!g111)) + ((!shiftx2x) & (shiftx3x) & (g87) & (!g109) & (g110) & (g111)) + ((!shiftx2x) & (shiftx3x) & (g87) & (g109) & (g110) & (!g111)) + ((!shiftx2x) & (shiftx3x) & (g87) & (g109) & (g110) & (g111)) + ((shiftx2x) & (!shiftx3x) & (!g87) & (!g109) & (!g110) & (g111)) + ((shiftx2x) & (!shiftx3x) & (!g87) & (!g109) & (g110) & (g111)) + ((shiftx2x) & (!shiftx3x) & (!g87) & (g109) & (!g110) & (g111)) + ((shiftx2x) & (!shiftx3x) & (!g87) & (g109) & (g110) & (g111)) + ((shiftx2x) & (!shiftx3x) & (g87) & (!g109) & (!g110) & (g111)) + ((shiftx2x) & (!shiftx3x) & (g87) & (!g109) & (g110) & (g111)) + ((shiftx2x) & (!shiftx3x) & (g87) & (g109) & (!g110) & (g111)) + ((shiftx2x) & (!shiftx3x) & (g87) & (g109) & (g110) & (g111)) + ((shiftx2x) & (shiftx3x) & (g87) & (!g109) & (!g110) & (!g111)) + ((shiftx2x) & (shiftx3x) & (g87) & (!g109) & (!g110) & (g111)) + ((shiftx2x) & (shiftx3x) & (g87) & (!g109) & (g110) & (!g111)) + ((shiftx2x) & (shiftx3x) & (g87) & (!g109) & (g110) & (g111)) + ((shiftx2x) & (shiftx3x) & (g87) & (g109) & (!g110) & (!g111)) + ((shiftx2x) & (shiftx3x) & (g87) & (g109) & (!g110) & (g111)) + ((shiftx2x) & (shiftx3x) & (g87) & (g109) & (g110) & (!g111)) + ((shiftx2x) & (shiftx3x) & (g87) & (g109) & (g110) & (g111)));
	assign g285 = (((!shiftx2x) & (!shiftx3x) & (g98) & (!g99) & (!g100) & (!g102)) + ((!shiftx2x) & (!shiftx3x) & (g98) & (!g99) & (!g100) & (g102)) + ((!shiftx2x) & (!shiftx3x) & (g98) & (!g99) & (g100) & (!g102)) + ((!shiftx2x) & (!shiftx3x) & (g98) & (!g99) & (g100) & (g102)) + ((!shiftx2x) & (!shiftx3x) & (g98) & (g99) & (!g100) & (!g102)) + ((!shiftx2x) & (!shiftx3x) & (g98) & (g99) & (!g100) & (g102)) + ((!shiftx2x) & (!shiftx3x) & (g98) & (g99) & (g100) & (!g102)) + ((!shiftx2x) & (!shiftx3x) & (g98) & (g99) & (g100) & (g102)) + ((!shiftx2x) & (shiftx3x) & (!g98) & (g99) & (!g100) & (!g102)) + ((!shiftx2x) & (shiftx3x) & (!g98) & (g99) & (!g100) & (g102)) + ((!shiftx2x) & (shiftx3x) & (!g98) & (g99) & (g100) & (!g102)) + ((!shiftx2x) & (shiftx3x) & (!g98) & (g99) & (g100) & (g102)) + ((!shiftx2x) & (shiftx3x) & (g98) & (g99) & (!g100) & (!g102)) + ((!shiftx2x) & (shiftx3x) & (g98) & (g99) & (!g100) & (g102)) + ((!shiftx2x) & (shiftx3x) & (g98) & (g99) & (g100) & (!g102)) + ((!shiftx2x) & (shiftx3x) & (g98) & (g99) & (g100) & (g102)) + ((shiftx2x) & (!shiftx3x) & (!g98) & (!g99) & (g100) & (!g102)) + ((shiftx2x) & (!shiftx3x) & (!g98) & (!g99) & (g100) & (g102)) + ((shiftx2x) & (!shiftx3x) & (!g98) & (g99) & (g100) & (!g102)) + ((shiftx2x) & (!shiftx3x) & (!g98) & (g99) & (g100) & (g102)) + ((shiftx2x) & (!shiftx3x) & (g98) & (!g99) & (g100) & (!g102)) + ((shiftx2x) & (!shiftx3x) & (g98) & (!g99) & (g100) & (g102)) + ((shiftx2x) & (!shiftx3x) & (g98) & (g99) & (g100) & (!g102)) + ((shiftx2x) & (!shiftx3x) & (g98) & (g99) & (g100) & (g102)) + ((shiftx2x) & (shiftx3x) & (!g98) & (!g99) & (!g100) & (g102)) + ((shiftx2x) & (shiftx3x) & (!g98) & (!g99) & (g100) & (g102)) + ((shiftx2x) & (shiftx3x) & (!g98) & (g99) & (!g100) & (g102)) + ((shiftx2x) & (shiftx3x) & (!g98) & (g99) & (g100) & (g102)) + ((shiftx2x) & (shiftx3x) & (g98) & (!g99) & (!g100) & (g102)) + ((shiftx2x) & (shiftx3x) & (g98) & (!g99) & (g100) & (g102)) + ((shiftx2x) & (shiftx3x) & (g98) & (g99) & (!g100) & (g102)) + ((shiftx2x) & (shiftx3x) & (g98) & (g99) & (g100) & (g102)));
	assign g286 = (((!shiftx2x) & (!shiftx3x) & (!g92) & (g103) & (!g104) & (!g105)) + ((!shiftx2x) & (!shiftx3x) & (!g92) & (g103) & (!g104) & (g105)) + ((!shiftx2x) & (!shiftx3x) & (!g92) & (g103) & (g104) & (!g105)) + ((!shiftx2x) & (!shiftx3x) & (!g92) & (g103) & (g104) & (g105)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (g103) & (!g104) & (!g105)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (g103) & (!g104) & (g105)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (g103) & (g104) & (!g105)) + ((!shiftx2x) & (!shiftx3x) & (g92) & (g103) & (g104) & (g105)) + ((!shiftx2x) & (shiftx3x) & (!g92) & (!g103) & (g104) & (!g105)) + ((!shiftx2x) & (shiftx3x) & (!g92) & (!g103) & (g104) & (g105)) + ((!shiftx2x) & (shiftx3x) & (!g92) & (g103) & (g104) & (!g105)) + ((!shiftx2x) & (shiftx3x) & (!g92) & (g103) & (g104) & (g105)) + ((!shiftx2x) & (shiftx3x) & (g92) & (!g103) & (g104) & (!g105)) + ((!shiftx2x) & (shiftx3x) & (g92) & (!g103) & (g104) & (g105)) + ((!shiftx2x) & (shiftx3x) & (g92) & (g103) & (g104) & (!g105)) + ((!shiftx2x) & (shiftx3x) & (g92) & (g103) & (g104) & (g105)) + ((shiftx2x) & (!shiftx3x) & (!g92) & (!g103) & (!g104) & (g105)) + ((shiftx2x) & (!shiftx3x) & (!g92) & (!g103) & (g104) & (g105)) + ((shiftx2x) & (!shiftx3x) & (!g92) & (g103) & (!g104) & (g105)) + ((shiftx2x) & (!shiftx3x) & (!g92) & (g103) & (g104) & (g105)) + ((shiftx2x) & (!shiftx3x) & (g92) & (!g103) & (!g104) & (g105)) + ((shiftx2x) & (!shiftx3x) & (g92) & (!g103) & (g104) & (g105)) + ((shiftx2x) & (!shiftx3x) & (g92) & (g103) & (!g104) & (g105)) + ((shiftx2x) & (!shiftx3x) & (g92) & (g103) & (g104) & (g105)) + ((shiftx2x) & (shiftx3x) & (g92) & (!g103) & (!g104) & (!g105)) + ((shiftx2x) & (shiftx3x) & (g92) & (!g103) & (!g104) & (g105)) + ((shiftx2x) & (shiftx3x) & (g92) & (!g103) & (g104) & (!g105)) + ((shiftx2x) & (shiftx3x) & (g92) & (!g103) & (g104) & (g105)) + ((shiftx2x) & (shiftx3x) & (g92) & (g103) & (!g104) & (!g105)) + ((shiftx2x) & (shiftx3x) & (g92) & (g103) & (!g104) & (g105)) + ((shiftx2x) & (shiftx3x) & (g92) & (g103) & (g104) & (!g105)) + ((shiftx2x) & (shiftx3x) & (g92) & (g103) & (g104) & (g105)));
	assign g287 = (((!shiftx4x) & (!shiftx5x) & (!g283) & (g284) & (!g285) & (!g286)) + ((!shiftx4x) & (!shiftx5x) & (!g283) & (g284) & (!g285) & (g286)) + ((!shiftx4x) & (!shiftx5x) & (!g283) & (g284) & (g285) & (!g286)) + ((!shiftx4x) & (!shiftx5x) & (!g283) & (g284) & (g285) & (g286)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (g284) & (!g285) & (!g286)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (g284) & (!g285) & (g286)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (g284) & (g285) & (!g286)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (g284) & (g285) & (g286)) + ((!shiftx4x) & (shiftx5x) & (!g283) & (!g284) & (g285) & (!g286)) + ((!shiftx4x) & (shiftx5x) & (!g283) & (!g284) & (g285) & (g286)) + ((!shiftx4x) & (shiftx5x) & (!g283) & (g284) & (g285) & (!g286)) + ((!shiftx4x) & (shiftx5x) & (!g283) & (g284) & (g285) & (g286)) + ((!shiftx4x) & (shiftx5x) & (g283) & (!g284) & (g285) & (!g286)) + ((!shiftx4x) & (shiftx5x) & (g283) & (!g284) & (g285) & (g286)) + ((!shiftx4x) & (shiftx5x) & (g283) & (g284) & (g285) & (!g286)) + ((!shiftx4x) & (shiftx5x) & (g283) & (g284) & (g285) & (g286)) + ((shiftx4x) & (!shiftx5x) & (g283) & (!g284) & (!g285) & (!g286)) + ((shiftx4x) & (!shiftx5x) & (g283) & (!g284) & (!g285) & (g286)) + ((shiftx4x) & (!shiftx5x) & (g283) & (!g284) & (g285) & (!g286)) + ((shiftx4x) & (!shiftx5x) & (g283) & (!g284) & (g285) & (g286)) + ((shiftx4x) & (!shiftx5x) & (g283) & (g284) & (!g285) & (!g286)) + ((shiftx4x) & (!shiftx5x) & (g283) & (g284) & (!g285) & (g286)) + ((shiftx4x) & (!shiftx5x) & (g283) & (g284) & (g285) & (!g286)) + ((shiftx4x) & (!shiftx5x) & (g283) & (g284) & (g285) & (g286)) + ((shiftx4x) & (shiftx5x) & (!g283) & (!g284) & (!g285) & (g286)) + ((shiftx4x) & (shiftx5x) & (!g283) & (!g284) & (g285) & (g286)) + ((shiftx4x) & (shiftx5x) & (!g283) & (g284) & (!g285) & (g286)) + ((shiftx4x) & (shiftx5x) & (!g283) & (g284) & (g285) & (g286)) + ((shiftx4x) & (shiftx5x) & (g283) & (!g284) & (!g285) & (g286)) + ((shiftx4x) & (shiftx5x) & (g283) & (!g284) & (g285) & (g286)) + ((shiftx4x) & (shiftx5x) & (g283) & (g284) & (!g285) & (g286)) + ((shiftx4x) & (shiftx5x) & (g283) & (g284) & (g285) & (g286)));
	assign g288 = (((!shiftx2x) & (!shiftx3x) & (!g108) & (g114) & (!g115) & (!g116)) + ((!shiftx2x) & (!shiftx3x) & (!g108) & (g114) & (!g115) & (g116)) + ((!shiftx2x) & (!shiftx3x) & (!g108) & (g114) & (g115) & (!g116)) + ((!shiftx2x) & (!shiftx3x) & (!g108) & (g114) & (g115) & (g116)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (g114) & (!g115) & (!g116)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (g114) & (!g115) & (g116)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (g114) & (g115) & (!g116)) + ((!shiftx2x) & (!shiftx3x) & (g108) & (g114) & (g115) & (g116)) + ((!shiftx2x) & (shiftx3x) & (!g108) & (!g114) & (g115) & (!g116)) + ((!shiftx2x) & (shiftx3x) & (!g108) & (!g114) & (g115) & (g116)) + ((!shiftx2x) & (shiftx3x) & (!g108) & (g114) & (g115) & (!g116)) + ((!shiftx2x) & (shiftx3x) & (!g108) & (g114) & (g115) & (g116)) + ((!shiftx2x) & (shiftx3x) & (g108) & (!g114) & (g115) & (!g116)) + ((!shiftx2x) & (shiftx3x) & (g108) & (!g114) & (g115) & (g116)) + ((!shiftx2x) & (shiftx3x) & (g108) & (g114) & (g115) & (!g116)) + ((!shiftx2x) & (shiftx3x) & (g108) & (g114) & (g115) & (g116)) + ((shiftx2x) & (!shiftx3x) & (!g108) & (!g114) & (!g115) & (g116)) + ((shiftx2x) & (!shiftx3x) & (!g108) & (!g114) & (g115) & (g116)) + ((shiftx2x) & (!shiftx3x) & (!g108) & (g114) & (!g115) & (g116)) + ((shiftx2x) & (!shiftx3x) & (!g108) & (g114) & (g115) & (g116)) + ((shiftx2x) & (!shiftx3x) & (g108) & (!g114) & (!g115) & (g116)) + ((shiftx2x) & (!shiftx3x) & (g108) & (!g114) & (g115) & (g116)) + ((shiftx2x) & (!shiftx3x) & (g108) & (g114) & (!g115) & (g116)) + ((shiftx2x) & (!shiftx3x) & (g108) & (g114) & (g115) & (g116)) + ((shiftx2x) & (shiftx3x) & (g108) & (!g114) & (!g115) & (!g116)) + ((shiftx2x) & (shiftx3x) & (g108) & (!g114) & (!g115) & (g116)) + ((shiftx2x) & (shiftx3x) & (g108) & (!g114) & (g115) & (!g116)) + ((shiftx2x) & (shiftx3x) & (g108) & (!g114) & (g115) & (g116)) + ((shiftx2x) & (shiftx3x) & (g108) & (g114) & (!g115) & (!g116)) + ((shiftx2x) & (shiftx3x) & (g108) & (g114) & (!g115) & (g116)) + ((shiftx2x) & (shiftx3x) & (g108) & (g114) & (g115) & (!g116)) + ((shiftx2x) & (shiftx3x) & (g108) & (g114) & (g115) & (g116)));
	assign g289 = (((!shiftx2x) & (!shiftx3x) & (!g113) & (g124) & (!g125) & (!g126)) + ((!shiftx2x) & (!shiftx3x) & (!g113) & (g124) & (!g125) & (g126)) + ((!shiftx2x) & (!shiftx3x) & (!g113) & (g124) & (g125) & (!g126)) + ((!shiftx2x) & (!shiftx3x) & (!g113) & (g124) & (g125) & (g126)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (g124) & (!g125) & (!g126)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (g124) & (!g125) & (g126)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (g124) & (g125) & (!g126)) + ((!shiftx2x) & (!shiftx3x) & (g113) & (g124) & (g125) & (g126)) + ((!shiftx2x) & (shiftx3x) & (!g113) & (!g124) & (g125) & (!g126)) + ((!shiftx2x) & (shiftx3x) & (!g113) & (!g124) & (g125) & (g126)) + ((!shiftx2x) & (shiftx3x) & (!g113) & (g124) & (g125) & (!g126)) + ((!shiftx2x) & (shiftx3x) & (!g113) & (g124) & (g125) & (g126)) + ((!shiftx2x) & (shiftx3x) & (g113) & (!g124) & (g125) & (!g126)) + ((!shiftx2x) & (shiftx3x) & (g113) & (!g124) & (g125) & (g126)) + ((!shiftx2x) & (shiftx3x) & (g113) & (g124) & (g125) & (!g126)) + ((!shiftx2x) & (shiftx3x) & (g113) & (g124) & (g125) & (g126)) + ((shiftx2x) & (!shiftx3x) & (!g113) & (!g124) & (!g125) & (g126)) + ((shiftx2x) & (!shiftx3x) & (!g113) & (!g124) & (g125) & (g126)) + ((shiftx2x) & (!shiftx3x) & (!g113) & (g124) & (!g125) & (g126)) + ((shiftx2x) & (!shiftx3x) & (!g113) & (g124) & (g125) & (g126)) + ((shiftx2x) & (!shiftx3x) & (g113) & (!g124) & (!g125) & (g126)) + ((shiftx2x) & (!shiftx3x) & (g113) & (!g124) & (g125) & (g126)) + ((shiftx2x) & (!shiftx3x) & (g113) & (g124) & (!g125) & (g126)) + ((shiftx2x) & (!shiftx3x) & (g113) & (g124) & (g125) & (g126)) + ((shiftx2x) & (shiftx3x) & (g113) & (!g124) & (!g125) & (!g126)) + ((shiftx2x) & (shiftx3x) & (g113) & (!g124) & (!g125) & (g126)) + ((shiftx2x) & (shiftx3x) & (g113) & (!g124) & (g125) & (!g126)) + ((shiftx2x) & (shiftx3x) & (g113) & (!g124) & (g125) & (g126)) + ((shiftx2x) & (shiftx3x) & (g113) & (g124) & (!g125) & (!g126)) + ((shiftx2x) & (shiftx3x) & (g113) & (g124) & (!g125) & (g126)) + ((shiftx2x) & (shiftx3x) & (g113) & (g124) & (g125) & (!g126)) + ((shiftx2x) & (shiftx3x) & (g113) & (g124) & (g125) & (g126)));
	assign g290 = (((!shiftx2x) & (!shiftx3x) & (g93) & (!g94) & (!g95) & (!g118)) + ((!shiftx2x) & (!shiftx3x) & (g93) & (!g94) & (!g95) & (g118)) + ((!shiftx2x) & (!shiftx3x) & (g93) & (!g94) & (g95) & (!g118)) + ((!shiftx2x) & (!shiftx3x) & (g93) & (!g94) & (g95) & (g118)) + ((!shiftx2x) & (!shiftx3x) & (g93) & (g94) & (!g95) & (!g118)) + ((!shiftx2x) & (!shiftx3x) & (g93) & (g94) & (!g95) & (g118)) + ((!shiftx2x) & (!shiftx3x) & (g93) & (g94) & (g95) & (!g118)) + ((!shiftx2x) & (!shiftx3x) & (g93) & (g94) & (g95) & (g118)) + ((!shiftx2x) & (shiftx3x) & (!g93) & (g94) & (!g95) & (!g118)) + ((!shiftx2x) & (shiftx3x) & (!g93) & (g94) & (!g95) & (g118)) + ((!shiftx2x) & (shiftx3x) & (!g93) & (g94) & (g95) & (!g118)) + ((!shiftx2x) & (shiftx3x) & (!g93) & (g94) & (g95) & (g118)) + ((!shiftx2x) & (shiftx3x) & (g93) & (g94) & (!g95) & (!g118)) + ((!shiftx2x) & (shiftx3x) & (g93) & (g94) & (!g95) & (g118)) + ((!shiftx2x) & (shiftx3x) & (g93) & (g94) & (g95) & (!g118)) + ((!shiftx2x) & (shiftx3x) & (g93) & (g94) & (g95) & (g118)) + ((shiftx2x) & (!shiftx3x) & (!g93) & (!g94) & (g95) & (!g118)) + ((shiftx2x) & (!shiftx3x) & (!g93) & (!g94) & (g95) & (g118)) + ((shiftx2x) & (!shiftx3x) & (!g93) & (g94) & (g95) & (!g118)) + ((shiftx2x) & (!shiftx3x) & (!g93) & (g94) & (g95) & (g118)) + ((shiftx2x) & (!shiftx3x) & (g93) & (!g94) & (g95) & (!g118)) + ((shiftx2x) & (!shiftx3x) & (g93) & (!g94) & (g95) & (g118)) + ((shiftx2x) & (!shiftx3x) & (g93) & (g94) & (g95) & (!g118)) + ((shiftx2x) & (!shiftx3x) & (g93) & (g94) & (g95) & (g118)) + ((shiftx2x) & (shiftx3x) & (!g93) & (!g94) & (!g95) & (g118)) + ((shiftx2x) & (shiftx3x) & (!g93) & (!g94) & (g95) & (g118)) + ((shiftx2x) & (shiftx3x) & (!g93) & (g94) & (!g95) & (g118)) + ((shiftx2x) & (shiftx3x) & (!g93) & (g94) & (g95) & (g118)) + ((shiftx2x) & (shiftx3x) & (g93) & (!g94) & (!g95) & (g118)) + ((shiftx2x) & (shiftx3x) & (g93) & (!g94) & (g95) & (g118)) + ((shiftx2x) & (shiftx3x) & (g93) & (g94) & (!g95) & (g118)) + ((shiftx2x) & (shiftx3x) & (g93) & (g94) & (g95) & (g118)));
	assign g291 = (((!shiftx2x) & (!shiftx3x) & (g119) & (!g120) & (!g121) & (!g123)) + ((!shiftx2x) & (!shiftx3x) & (g119) & (!g120) & (!g121) & (g123)) + ((!shiftx2x) & (!shiftx3x) & (g119) & (!g120) & (g121) & (!g123)) + ((!shiftx2x) & (!shiftx3x) & (g119) & (!g120) & (g121) & (g123)) + ((!shiftx2x) & (!shiftx3x) & (g119) & (g120) & (!g121) & (!g123)) + ((!shiftx2x) & (!shiftx3x) & (g119) & (g120) & (!g121) & (g123)) + ((!shiftx2x) & (!shiftx3x) & (g119) & (g120) & (g121) & (!g123)) + ((!shiftx2x) & (!shiftx3x) & (g119) & (g120) & (g121) & (g123)) + ((!shiftx2x) & (shiftx3x) & (!g119) & (g120) & (!g121) & (!g123)) + ((!shiftx2x) & (shiftx3x) & (!g119) & (g120) & (!g121) & (g123)) + ((!shiftx2x) & (shiftx3x) & (!g119) & (g120) & (g121) & (!g123)) + ((!shiftx2x) & (shiftx3x) & (!g119) & (g120) & (g121) & (g123)) + ((!shiftx2x) & (shiftx3x) & (g119) & (g120) & (!g121) & (!g123)) + ((!shiftx2x) & (shiftx3x) & (g119) & (g120) & (!g121) & (g123)) + ((!shiftx2x) & (shiftx3x) & (g119) & (g120) & (g121) & (!g123)) + ((!shiftx2x) & (shiftx3x) & (g119) & (g120) & (g121) & (g123)) + ((shiftx2x) & (!shiftx3x) & (!g119) & (!g120) & (g121) & (!g123)) + ((shiftx2x) & (!shiftx3x) & (!g119) & (!g120) & (g121) & (g123)) + ((shiftx2x) & (!shiftx3x) & (!g119) & (g120) & (g121) & (!g123)) + ((shiftx2x) & (!shiftx3x) & (!g119) & (g120) & (g121) & (g123)) + ((shiftx2x) & (!shiftx3x) & (g119) & (!g120) & (g121) & (!g123)) + ((shiftx2x) & (!shiftx3x) & (g119) & (!g120) & (g121) & (g123)) + ((shiftx2x) & (!shiftx3x) & (g119) & (g120) & (g121) & (!g123)) + ((shiftx2x) & (!shiftx3x) & (g119) & (g120) & (g121) & (g123)) + ((shiftx2x) & (shiftx3x) & (!g119) & (!g120) & (!g121) & (g123)) + ((shiftx2x) & (shiftx3x) & (!g119) & (!g120) & (g121) & (g123)) + ((shiftx2x) & (shiftx3x) & (!g119) & (g120) & (!g121) & (g123)) + ((shiftx2x) & (shiftx3x) & (!g119) & (g120) & (g121) & (g123)) + ((shiftx2x) & (shiftx3x) & (g119) & (!g120) & (!g121) & (g123)) + ((shiftx2x) & (shiftx3x) & (g119) & (!g120) & (g121) & (g123)) + ((shiftx2x) & (shiftx3x) & (g119) & (g120) & (!g121) & (g123)) + ((shiftx2x) & (shiftx3x) & (g119) & (g120) & (g121) & (g123)));
	assign g292 = (((!shiftx4x) & (!shiftx5x) & (!g288) & (!g289) & (g290) & (!g291)) + ((!shiftx4x) & (!shiftx5x) & (!g288) & (!g289) & (g290) & (g291)) + ((!shiftx4x) & (!shiftx5x) & (!g288) & (g289) & (g290) & (!g291)) + ((!shiftx4x) & (!shiftx5x) & (!g288) & (g289) & (g290) & (g291)) + ((!shiftx4x) & (!shiftx5x) & (g288) & (!g289) & (g290) & (!g291)) + ((!shiftx4x) & (!shiftx5x) & (g288) & (!g289) & (g290) & (g291)) + ((!shiftx4x) & (!shiftx5x) & (g288) & (g289) & (g290) & (!g291)) + ((!shiftx4x) & (!shiftx5x) & (g288) & (g289) & (g290) & (g291)) + ((!shiftx4x) & (shiftx5x) & (!g288) & (g289) & (!g290) & (!g291)) + ((!shiftx4x) & (shiftx5x) & (!g288) & (g289) & (!g290) & (g291)) + ((!shiftx4x) & (shiftx5x) & (!g288) & (g289) & (g290) & (!g291)) + ((!shiftx4x) & (shiftx5x) & (!g288) & (g289) & (g290) & (g291)) + ((!shiftx4x) & (shiftx5x) & (g288) & (g289) & (!g290) & (!g291)) + ((!shiftx4x) & (shiftx5x) & (g288) & (g289) & (!g290) & (g291)) + ((!shiftx4x) & (shiftx5x) & (g288) & (g289) & (g290) & (!g291)) + ((!shiftx4x) & (shiftx5x) & (g288) & (g289) & (g290) & (g291)) + ((shiftx4x) & (!shiftx5x) & (!g288) & (!g289) & (!g290) & (g291)) + ((shiftx4x) & (!shiftx5x) & (!g288) & (!g289) & (g290) & (g291)) + ((shiftx4x) & (!shiftx5x) & (!g288) & (g289) & (!g290) & (g291)) + ((shiftx4x) & (!shiftx5x) & (!g288) & (g289) & (g290) & (g291)) + ((shiftx4x) & (!shiftx5x) & (g288) & (!g289) & (!g290) & (g291)) + ((shiftx4x) & (!shiftx5x) & (g288) & (!g289) & (g290) & (g291)) + ((shiftx4x) & (!shiftx5x) & (g288) & (g289) & (!g290) & (g291)) + ((shiftx4x) & (!shiftx5x) & (g288) & (g289) & (g290) & (g291)) + ((shiftx4x) & (shiftx5x) & (g288) & (!g289) & (!g290) & (!g291)) + ((shiftx4x) & (shiftx5x) & (g288) & (!g289) & (!g290) & (g291)) + ((shiftx4x) & (shiftx5x) & (g288) & (!g289) & (g290) & (!g291)) + ((shiftx4x) & (shiftx5x) & (g288) & (!g289) & (g290) & (g291)) + ((shiftx4x) & (shiftx5x) & (g288) & (g289) & (!g290) & (!g291)) + ((shiftx4x) & (shiftx5x) & (g288) & (g289) & (!g290) & (g291)) + ((shiftx4x) & (shiftx5x) & (g288) & (g289) & (g290) & (!g291)) + ((shiftx4x) & (shiftx5x) & (g288) & (g289) & (g290) & (g291)));
	assign resultx14x = (((!sk[36]) & (shiftx6x) & (!g287) & (!g292)) + ((!sk[36]) & (shiftx6x) & (!g287) & (g292)) + ((!sk[36]) & (shiftx6x) & (g287) & (!g292)) + ((!sk[36]) & (shiftx6x) & (g287) & (g292)) + ((sk[36]) & (!shiftx6x) & (!g287) & (g292)) + ((sk[36]) & (!shiftx6x) & (g287) & (g292)) + ((sk[36]) & (shiftx6x) & (g287) & (!g292)) + ((sk[36]) & (shiftx6x) & (g287) & (g292)));
	assign g294 = (((!shiftx2x) & (!shiftx3x) & (g131) & (!g132) & (!g133) & (!g135)) + ((!shiftx2x) & (!shiftx3x) & (g131) & (!g132) & (!g133) & (g135)) + ((!shiftx2x) & (!shiftx3x) & (g131) & (!g132) & (g133) & (!g135)) + ((!shiftx2x) & (!shiftx3x) & (g131) & (!g132) & (g133) & (g135)) + ((!shiftx2x) & (!shiftx3x) & (g131) & (g132) & (!g133) & (!g135)) + ((!shiftx2x) & (!shiftx3x) & (g131) & (g132) & (!g133) & (g135)) + ((!shiftx2x) & (!shiftx3x) & (g131) & (g132) & (g133) & (!g135)) + ((!shiftx2x) & (!shiftx3x) & (g131) & (g132) & (g133) & (g135)) + ((!shiftx2x) & (shiftx3x) & (!g131) & (g132) & (!g133) & (!g135)) + ((!shiftx2x) & (shiftx3x) & (!g131) & (g132) & (!g133) & (g135)) + ((!shiftx2x) & (shiftx3x) & (!g131) & (g132) & (g133) & (!g135)) + ((!shiftx2x) & (shiftx3x) & (!g131) & (g132) & (g133) & (g135)) + ((!shiftx2x) & (shiftx3x) & (g131) & (g132) & (!g133) & (!g135)) + ((!shiftx2x) & (shiftx3x) & (g131) & (g132) & (!g133) & (g135)) + ((!shiftx2x) & (shiftx3x) & (g131) & (g132) & (g133) & (!g135)) + ((!shiftx2x) & (shiftx3x) & (g131) & (g132) & (g133) & (g135)) + ((shiftx2x) & (!shiftx3x) & (!g131) & (!g132) & (g133) & (!g135)) + ((shiftx2x) & (!shiftx3x) & (!g131) & (!g132) & (g133) & (g135)) + ((shiftx2x) & (!shiftx3x) & (!g131) & (g132) & (g133) & (!g135)) + ((shiftx2x) & (!shiftx3x) & (!g131) & (g132) & (g133) & (g135)) + ((shiftx2x) & (!shiftx3x) & (g131) & (!g132) & (g133) & (!g135)) + ((shiftx2x) & (!shiftx3x) & (g131) & (!g132) & (g133) & (g135)) + ((shiftx2x) & (!shiftx3x) & (g131) & (g132) & (g133) & (!g135)) + ((shiftx2x) & (!shiftx3x) & (g131) & (g132) & (g133) & (g135)) + ((shiftx2x) & (shiftx3x) & (!g131) & (!g132) & (!g133) & (g135)) + ((shiftx2x) & (shiftx3x) & (!g131) & (!g132) & (g133) & (g135)) + ((shiftx2x) & (shiftx3x) & (!g131) & (g132) & (!g133) & (g135)) + ((shiftx2x) & (shiftx3x) & (!g131) & (g132) & (g133) & (g135)) + ((shiftx2x) & (shiftx3x) & (g131) & (!g132) & (!g133) & (g135)) + ((shiftx2x) & (shiftx3x) & (g131) & (!g132) & (g133) & (g135)) + ((shiftx2x) & (shiftx3x) & (g131) & (g132) & (!g133) & (g135)) + ((shiftx2x) & (shiftx3x) & (g131) & (g132) & (g133) & (g135)));
	assign g295 = (((!shiftx2x) & (!shiftx3x) & (!g130) & (g167) & (!g168) & (!g169)) + ((!shiftx2x) & (!shiftx3x) & (!g130) & (g167) & (!g168) & (g169)) + ((!shiftx2x) & (!shiftx3x) & (!g130) & (g167) & (g168) & (!g169)) + ((!shiftx2x) & (!shiftx3x) & (!g130) & (g167) & (g168) & (g169)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (g167) & (!g168) & (!g169)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (g167) & (!g168) & (g169)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (g167) & (g168) & (!g169)) + ((!shiftx2x) & (!shiftx3x) & (g130) & (g167) & (g168) & (g169)) + ((!shiftx2x) & (shiftx3x) & (!g130) & (!g167) & (g168) & (!g169)) + ((!shiftx2x) & (shiftx3x) & (!g130) & (!g167) & (g168) & (g169)) + ((!shiftx2x) & (shiftx3x) & (!g130) & (g167) & (g168) & (!g169)) + ((!shiftx2x) & (shiftx3x) & (!g130) & (g167) & (g168) & (g169)) + ((!shiftx2x) & (shiftx3x) & (g130) & (!g167) & (g168) & (!g169)) + ((!shiftx2x) & (shiftx3x) & (g130) & (!g167) & (g168) & (g169)) + ((!shiftx2x) & (shiftx3x) & (g130) & (g167) & (g168) & (!g169)) + ((!shiftx2x) & (shiftx3x) & (g130) & (g167) & (g168) & (g169)) + ((shiftx2x) & (!shiftx3x) & (!g130) & (!g167) & (!g168) & (g169)) + ((shiftx2x) & (!shiftx3x) & (!g130) & (!g167) & (g168) & (g169)) + ((shiftx2x) & (!shiftx3x) & (!g130) & (g167) & (!g168) & (g169)) + ((shiftx2x) & (!shiftx3x) & (!g130) & (g167) & (g168) & (g169)) + ((shiftx2x) & (!shiftx3x) & (g130) & (!g167) & (!g168) & (g169)) + ((shiftx2x) & (!shiftx3x) & (g130) & (!g167) & (g168) & (g169)) + ((shiftx2x) & (!shiftx3x) & (g130) & (g167) & (!g168) & (g169)) + ((shiftx2x) & (!shiftx3x) & (g130) & (g167) & (g168) & (g169)) + ((shiftx2x) & (shiftx3x) & (g130) & (!g167) & (!g168) & (!g169)) + ((shiftx2x) & (shiftx3x) & (g130) & (!g167) & (!g168) & (g169)) + ((shiftx2x) & (shiftx3x) & (g130) & (!g167) & (g168) & (!g169)) + ((shiftx2x) & (shiftx3x) & (g130) & (!g167) & (g168) & (g169)) + ((shiftx2x) & (shiftx3x) & (g130) & (g167) & (!g168) & (!g169)) + ((shiftx2x) & (shiftx3x) & (g130) & (g167) & (!g168) & (g169)) + ((shiftx2x) & (shiftx3x) & (g130) & (g167) & (g168) & (!g169)) + ((shiftx2x) & (shiftx3x) & (g130) & (g167) & (g168) & (g169)));
	assign g296 = (((!shiftx2x) & (!shiftx3x) & (g136) & (!g137) & (!g138) & (!g145)) + ((!shiftx2x) & (!shiftx3x) & (g136) & (!g137) & (!g138) & (g145)) + ((!shiftx2x) & (!shiftx3x) & (g136) & (!g137) & (g138) & (!g145)) + ((!shiftx2x) & (!shiftx3x) & (g136) & (!g137) & (g138) & (g145)) + ((!shiftx2x) & (!shiftx3x) & (g136) & (g137) & (!g138) & (!g145)) + ((!shiftx2x) & (!shiftx3x) & (g136) & (g137) & (!g138) & (g145)) + ((!shiftx2x) & (!shiftx3x) & (g136) & (g137) & (g138) & (!g145)) + ((!shiftx2x) & (!shiftx3x) & (g136) & (g137) & (g138) & (g145)) + ((!shiftx2x) & (shiftx3x) & (!g136) & (g137) & (!g138) & (!g145)) + ((!shiftx2x) & (shiftx3x) & (!g136) & (g137) & (!g138) & (g145)) + ((!shiftx2x) & (shiftx3x) & (!g136) & (g137) & (g138) & (!g145)) + ((!shiftx2x) & (shiftx3x) & (!g136) & (g137) & (g138) & (g145)) + ((!shiftx2x) & (shiftx3x) & (g136) & (g137) & (!g138) & (!g145)) + ((!shiftx2x) & (shiftx3x) & (g136) & (g137) & (!g138) & (g145)) + ((!shiftx2x) & (shiftx3x) & (g136) & (g137) & (g138) & (!g145)) + ((!shiftx2x) & (shiftx3x) & (g136) & (g137) & (g138) & (g145)) + ((shiftx2x) & (!shiftx3x) & (!g136) & (!g137) & (g138) & (!g145)) + ((shiftx2x) & (!shiftx3x) & (!g136) & (!g137) & (g138) & (g145)) + ((shiftx2x) & (!shiftx3x) & (!g136) & (g137) & (g138) & (!g145)) + ((shiftx2x) & (!shiftx3x) & (!g136) & (g137) & (g138) & (g145)) + ((shiftx2x) & (!shiftx3x) & (g136) & (!g137) & (g138) & (!g145)) + ((shiftx2x) & (!shiftx3x) & (g136) & (!g137) & (g138) & (g145)) + ((shiftx2x) & (!shiftx3x) & (g136) & (g137) & (g138) & (!g145)) + ((shiftx2x) & (!shiftx3x) & (g136) & (g137) & (g138) & (g145)) + ((shiftx2x) & (shiftx3x) & (!g136) & (!g137) & (!g138) & (g145)) + ((shiftx2x) & (shiftx3x) & (!g136) & (!g137) & (g138) & (g145)) + ((shiftx2x) & (shiftx3x) & (!g136) & (g137) & (!g138) & (g145)) + ((shiftx2x) & (shiftx3x) & (!g136) & (g137) & (g138) & (g145)) + ((shiftx2x) & (shiftx3x) & (g136) & (!g137) & (!g138) & (g145)) + ((shiftx2x) & (shiftx3x) & (g136) & (!g137) & (g138) & (g145)) + ((shiftx2x) & (shiftx3x) & (g136) & (g137) & (!g138) & (g145)) + ((shiftx2x) & (shiftx3x) & (g136) & (g137) & (g138) & (g145)));
	assign g297 = (((!shiftx2x) & (!shiftx3x) & (!g140) & (g146) & (!g147) & (!g148)) + ((!shiftx2x) & (!shiftx3x) & (!g140) & (g146) & (!g147) & (g148)) + ((!shiftx2x) & (!shiftx3x) & (!g140) & (g146) & (g147) & (!g148)) + ((!shiftx2x) & (!shiftx3x) & (!g140) & (g146) & (g147) & (g148)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (g146) & (!g147) & (!g148)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (g146) & (!g147) & (g148)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (g146) & (g147) & (!g148)) + ((!shiftx2x) & (!shiftx3x) & (g140) & (g146) & (g147) & (g148)) + ((!shiftx2x) & (shiftx3x) & (!g140) & (!g146) & (g147) & (!g148)) + ((!shiftx2x) & (shiftx3x) & (!g140) & (!g146) & (g147) & (g148)) + ((!shiftx2x) & (shiftx3x) & (!g140) & (g146) & (g147) & (!g148)) + ((!shiftx2x) & (shiftx3x) & (!g140) & (g146) & (g147) & (g148)) + ((!shiftx2x) & (shiftx3x) & (g140) & (!g146) & (g147) & (!g148)) + ((!shiftx2x) & (shiftx3x) & (g140) & (!g146) & (g147) & (g148)) + ((!shiftx2x) & (shiftx3x) & (g140) & (g146) & (g147) & (!g148)) + ((!shiftx2x) & (shiftx3x) & (g140) & (g146) & (g147) & (g148)) + ((shiftx2x) & (!shiftx3x) & (!g140) & (!g146) & (!g147) & (g148)) + ((shiftx2x) & (!shiftx3x) & (!g140) & (!g146) & (g147) & (g148)) + ((shiftx2x) & (!shiftx3x) & (!g140) & (g146) & (!g147) & (g148)) + ((shiftx2x) & (!shiftx3x) & (!g140) & (g146) & (g147) & (g148)) + ((shiftx2x) & (!shiftx3x) & (g140) & (!g146) & (!g147) & (g148)) + ((shiftx2x) & (!shiftx3x) & (g140) & (!g146) & (g147) & (g148)) + ((shiftx2x) & (!shiftx3x) & (g140) & (g146) & (!g147) & (g148)) + ((shiftx2x) & (!shiftx3x) & (g140) & (g146) & (g147) & (g148)) + ((shiftx2x) & (shiftx3x) & (g140) & (!g146) & (!g147) & (!g148)) + ((shiftx2x) & (shiftx3x) & (g140) & (!g146) & (!g147) & (g148)) + ((shiftx2x) & (shiftx3x) & (g140) & (!g146) & (g147) & (!g148)) + ((shiftx2x) & (shiftx3x) & (g140) & (!g146) & (g147) & (g148)) + ((shiftx2x) & (shiftx3x) & (g140) & (g146) & (!g147) & (!g148)) + ((shiftx2x) & (shiftx3x) & (g140) & (g146) & (!g147) & (g148)) + ((shiftx2x) & (shiftx3x) & (g140) & (g146) & (g147) & (!g148)) + ((shiftx2x) & (shiftx3x) & (g140) & (g146) & (g147) & (g148)));
	assign g298 = (((!shiftx4x) & (!shiftx5x) & (!g294) & (g295) & (!g296) & (!g297)) + ((!shiftx4x) & (!shiftx5x) & (!g294) & (g295) & (!g296) & (g297)) + ((!shiftx4x) & (!shiftx5x) & (!g294) & (g295) & (g296) & (!g297)) + ((!shiftx4x) & (!shiftx5x) & (!g294) & (g295) & (g296) & (g297)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (g295) & (!g296) & (!g297)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (g295) & (!g296) & (g297)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (g295) & (g296) & (!g297)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (g295) & (g296) & (g297)) + ((!shiftx4x) & (shiftx5x) & (!g294) & (!g295) & (g296) & (!g297)) + ((!shiftx4x) & (shiftx5x) & (!g294) & (!g295) & (g296) & (g297)) + ((!shiftx4x) & (shiftx5x) & (!g294) & (g295) & (g296) & (!g297)) + ((!shiftx4x) & (shiftx5x) & (!g294) & (g295) & (g296) & (g297)) + ((!shiftx4x) & (shiftx5x) & (g294) & (!g295) & (g296) & (!g297)) + ((!shiftx4x) & (shiftx5x) & (g294) & (!g295) & (g296) & (g297)) + ((!shiftx4x) & (shiftx5x) & (g294) & (g295) & (g296) & (!g297)) + ((!shiftx4x) & (shiftx5x) & (g294) & (g295) & (g296) & (g297)) + ((shiftx4x) & (!shiftx5x) & (g294) & (!g295) & (!g296) & (!g297)) + ((shiftx4x) & (!shiftx5x) & (g294) & (!g295) & (!g296) & (g297)) + ((shiftx4x) & (!shiftx5x) & (g294) & (!g295) & (g296) & (!g297)) + ((shiftx4x) & (!shiftx5x) & (g294) & (!g295) & (g296) & (g297)) + ((shiftx4x) & (!shiftx5x) & (g294) & (g295) & (!g296) & (!g297)) + ((shiftx4x) & (!shiftx5x) & (g294) & (g295) & (!g296) & (g297)) + ((shiftx4x) & (!shiftx5x) & (g294) & (g295) & (g296) & (!g297)) + ((shiftx4x) & (!shiftx5x) & (g294) & (g295) & (g296) & (g297)) + ((shiftx4x) & (shiftx5x) & (!g294) & (!g295) & (!g296) & (g297)) + ((shiftx4x) & (shiftx5x) & (!g294) & (!g295) & (g296) & (g297)) + ((shiftx4x) & (shiftx5x) & (!g294) & (g295) & (!g296) & (g297)) + ((shiftx4x) & (shiftx5x) & (!g294) & (g295) & (g296) & (g297)) + ((shiftx4x) & (shiftx5x) & (g294) & (!g295) & (!g296) & (g297)) + ((shiftx4x) & (shiftx5x) & (g294) & (!g295) & (g296) & (g297)) + ((shiftx4x) & (shiftx5x) & (g294) & (g295) & (!g296) & (g297)) + ((shiftx4x) & (shiftx5x) & (g294) & (g295) & (g296) & (g297)));
	assign g299 = (((!shiftx2x) & (!shiftx3x) & (g157) & (!g158) & (!g159) & (!g166)) + ((!shiftx2x) & (!shiftx3x) & (g157) & (!g158) & (!g159) & (g166)) + ((!shiftx2x) & (!shiftx3x) & (g157) & (!g158) & (g159) & (!g166)) + ((!shiftx2x) & (!shiftx3x) & (g157) & (!g158) & (g159) & (g166)) + ((!shiftx2x) & (!shiftx3x) & (g157) & (g158) & (!g159) & (!g166)) + ((!shiftx2x) & (!shiftx3x) & (g157) & (g158) & (!g159) & (g166)) + ((!shiftx2x) & (!shiftx3x) & (g157) & (g158) & (g159) & (!g166)) + ((!shiftx2x) & (!shiftx3x) & (g157) & (g158) & (g159) & (g166)) + ((!shiftx2x) & (shiftx3x) & (!g157) & (g158) & (!g159) & (!g166)) + ((!shiftx2x) & (shiftx3x) & (!g157) & (g158) & (!g159) & (g166)) + ((!shiftx2x) & (shiftx3x) & (!g157) & (g158) & (g159) & (!g166)) + ((!shiftx2x) & (shiftx3x) & (!g157) & (g158) & (g159) & (g166)) + ((!shiftx2x) & (shiftx3x) & (g157) & (g158) & (!g159) & (!g166)) + ((!shiftx2x) & (shiftx3x) & (g157) & (g158) & (!g159) & (g166)) + ((!shiftx2x) & (shiftx3x) & (g157) & (g158) & (g159) & (!g166)) + ((!shiftx2x) & (shiftx3x) & (g157) & (g158) & (g159) & (g166)) + ((shiftx2x) & (!shiftx3x) & (!g157) & (!g158) & (g159) & (!g166)) + ((shiftx2x) & (!shiftx3x) & (!g157) & (!g158) & (g159) & (g166)) + ((shiftx2x) & (!shiftx3x) & (!g157) & (g158) & (g159) & (!g166)) + ((shiftx2x) & (!shiftx3x) & (!g157) & (g158) & (g159) & (g166)) + ((shiftx2x) & (!shiftx3x) & (g157) & (!g158) & (g159) & (!g166)) + ((shiftx2x) & (!shiftx3x) & (g157) & (!g158) & (g159) & (g166)) + ((shiftx2x) & (!shiftx3x) & (g157) & (g158) & (g159) & (!g166)) + ((shiftx2x) & (!shiftx3x) & (g157) & (g158) & (g159) & (g166)) + ((shiftx2x) & (shiftx3x) & (!g157) & (!g158) & (!g159) & (g166)) + ((shiftx2x) & (shiftx3x) & (!g157) & (!g158) & (g159) & (g166)) + ((shiftx2x) & (shiftx3x) & (!g157) & (g158) & (!g159) & (g166)) + ((shiftx2x) & (shiftx3x) & (!g157) & (g158) & (g159) & (g166)) + ((shiftx2x) & (shiftx3x) & (g157) & (!g158) & (!g159) & (g166)) + ((shiftx2x) & (shiftx3x) & (g157) & (!g158) & (g159) & (g166)) + ((shiftx2x) & (shiftx3x) & (g157) & (g158) & (!g159) & (g166)) + ((shiftx2x) & (shiftx3x) & (g157) & (g158) & (g159) & (g166)));
	assign g300 = (((!shiftx2x) & (!shiftx3x) & (g152) & (!g153) & (!g154) & (!g156)) + ((!shiftx2x) & (!shiftx3x) & (g152) & (!g153) & (!g154) & (g156)) + ((!shiftx2x) & (!shiftx3x) & (g152) & (!g153) & (g154) & (!g156)) + ((!shiftx2x) & (!shiftx3x) & (g152) & (!g153) & (g154) & (g156)) + ((!shiftx2x) & (!shiftx3x) & (g152) & (g153) & (!g154) & (!g156)) + ((!shiftx2x) & (!shiftx3x) & (g152) & (g153) & (!g154) & (g156)) + ((!shiftx2x) & (!shiftx3x) & (g152) & (g153) & (g154) & (!g156)) + ((!shiftx2x) & (!shiftx3x) & (g152) & (g153) & (g154) & (g156)) + ((!shiftx2x) & (shiftx3x) & (!g152) & (g153) & (!g154) & (!g156)) + ((!shiftx2x) & (shiftx3x) & (!g152) & (g153) & (!g154) & (g156)) + ((!shiftx2x) & (shiftx3x) & (!g152) & (g153) & (g154) & (!g156)) + ((!shiftx2x) & (shiftx3x) & (!g152) & (g153) & (g154) & (g156)) + ((!shiftx2x) & (shiftx3x) & (g152) & (g153) & (!g154) & (!g156)) + ((!shiftx2x) & (shiftx3x) & (g152) & (g153) & (!g154) & (g156)) + ((!shiftx2x) & (shiftx3x) & (g152) & (g153) & (g154) & (!g156)) + ((!shiftx2x) & (shiftx3x) & (g152) & (g153) & (g154) & (g156)) + ((shiftx2x) & (!shiftx3x) & (!g152) & (!g153) & (g154) & (!g156)) + ((shiftx2x) & (!shiftx3x) & (!g152) & (!g153) & (g154) & (g156)) + ((shiftx2x) & (!shiftx3x) & (!g152) & (g153) & (g154) & (!g156)) + ((shiftx2x) & (!shiftx3x) & (!g152) & (g153) & (g154) & (g156)) + ((shiftx2x) & (!shiftx3x) & (g152) & (!g153) & (g154) & (!g156)) + ((shiftx2x) & (!shiftx3x) & (g152) & (!g153) & (g154) & (g156)) + ((shiftx2x) & (!shiftx3x) & (g152) & (g153) & (g154) & (!g156)) + ((shiftx2x) & (!shiftx3x) & (g152) & (g153) & (g154) & (g156)) + ((shiftx2x) & (shiftx3x) & (!g152) & (!g153) & (!g154) & (g156)) + ((shiftx2x) & (shiftx3x) & (!g152) & (!g153) & (g154) & (g156)) + ((shiftx2x) & (shiftx3x) & (!g152) & (g153) & (!g154) & (g156)) + ((shiftx2x) & (shiftx3x) & (!g152) & (g153) & (g154) & (g156)) + ((shiftx2x) & (shiftx3x) & (g152) & (!g153) & (!g154) & (g156)) + ((shiftx2x) & (shiftx3x) & (g152) & (!g153) & (g154) & (g156)) + ((shiftx2x) & (shiftx3x) & (g152) & (g153) & (!g154) & (g156)) + ((shiftx2x) & (shiftx3x) & (g152) & (g153) & (g154) & (g156)));
	assign g301 = (((!shiftx2x) & (!shiftx3x) & (g141) & (!g142) & (!g143) & (!g161)) + ((!shiftx2x) & (!shiftx3x) & (g141) & (!g142) & (!g143) & (g161)) + ((!shiftx2x) & (!shiftx3x) & (g141) & (!g142) & (g143) & (!g161)) + ((!shiftx2x) & (!shiftx3x) & (g141) & (!g142) & (g143) & (g161)) + ((!shiftx2x) & (!shiftx3x) & (g141) & (g142) & (!g143) & (!g161)) + ((!shiftx2x) & (!shiftx3x) & (g141) & (g142) & (!g143) & (g161)) + ((!shiftx2x) & (!shiftx3x) & (g141) & (g142) & (g143) & (!g161)) + ((!shiftx2x) & (!shiftx3x) & (g141) & (g142) & (g143) & (g161)) + ((!shiftx2x) & (shiftx3x) & (!g141) & (g142) & (!g143) & (!g161)) + ((!shiftx2x) & (shiftx3x) & (!g141) & (g142) & (!g143) & (g161)) + ((!shiftx2x) & (shiftx3x) & (!g141) & (g142) & (g143) & (!g161)) + ((!shiftx2x) & (shiftx3x) & (!g141) & (g142) & (g143) & (g161)) + ((!shiftx2x) & (shiftx3x) & (g141) & (g142) & (!g143) & (!g161)) + ((!shiftx2x) & (shiftx3x) & (g141) & (g142) & (!g143) & (g161)) + ((!shiftx2x) & (shiftx3x) & (g141) & (g142) & (g143) & (!g161)) + ((!shiftx2x) & (shiftx3x) & (g141) & (g142) & (g143) & (g161)) + ((shiftx2x) & (!shiftx3x) & (!g141) & (!g142) & (g143) & (!g161)) + ((shiftx2x) & (!shiftx3x) & (!g141) & (!g142) & (g143) & (g161)) + ((shiftx2x) & (!shiftx3x) & (!g141) & (g142) & (g143) & (!g161)) + ((shiftx2x) & (!shiftx3x) & (!g141) & (g142) & (g143) & (g161)) + ((shiftx2x) & (!shiftx3x) & (g141) & (!g142) & (g143) & (!g161)) + ((shiftx2x) & (!shiftx3x) & (g141) & (!g142) & (g143) & (g161)) + ((shiftx2x) & (!shiftx3x) & (g141) & (g142) & (g143) & (!g161)) + ((shiftx2x) & (!shiftx3x) & (g141) & (g142) & (g143) & (g161)) + ((shiftx2x) & (shiftx3x) & (!g141) & (!g142) & (!g143) & (g161)) + ((shiftx2x) & (shiftx3x) & (!g141) & (!g142) & (g143) & (g161)) + ((shiftx2x) & (shiftx3x) & (!g141) & (g142) & (!g143) & (g161)) + ((shiftx2x) & (shiftx3x) & (!g141) & (g142) & (g143) & (g161)) + ((shiftx2x) & (shiftx3x) & (g141) & (!g142) & (!g143) & (g161)) + ((shiftx2x) & (shiftx3x) & (g141) & (!g142) & (g143) & (g161)) + ((shiftx2x) & (shiftx3x) & (g141) & (g142) & (!g143) & (g161)) + ((shiftx2x) & (shiftx3x) & (g141) & (g142) & (g143) & (g161)));
	assign g302 = (((!shiftx2x) & (!shiftx3x) & (!g151) & (g162) & (!g163) & (!g164)) + ((!shiftx2x) & (!shiftx3x) & (!g151) & (g162) & (!g163) & (g164)) + ((!shiftx2x) & (!shiftx3x) & (!g151) & (g162) & (g163) & (!g164)) + ((!shiftx2x) & (!shiftx3x) & (!g151) & (g162) & (g163) & (g164)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (g162) & (!g163) & (!g164)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (g162) & (!g163) & (g164)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (g162) & (g163) & (!g164)) + ((!shiftx2x) & (!shiftx3x) & (g151) & (g162) & (g163) & (g164)) + ((!shiftx2x) & (shiftx3x) & (!g151) & (!g162) & (g163) & (!g164)) + ((!shiftx2x) & (shiftx3x) & (!g151) & (!g162) & (g163) & (g164)) + ((!shiftx2x) & (shiftx3x) & (!g151) & (g162) & (g163) & (!g164)) + ((!shiftx2x) & (shiftx3x) & (!g151) & (g162) & (g163) & (g164)) + ((!shiftx2x) & (shiftx3x) & (g151) & (!g162) & (g163) & (!g164)) + ((!shiftx2x) & (shiftx3x) & (g151) & (!g162) & (g163) & (g164)) + ((!shiftx2x) & (shiftx3x) & (g151) & (g162) & (g163) & (!g164)) + ((!shiftx2x) & (shiftx3x) & (g151) & (g162) & (g163) & (g164)) + ((shiftx2x) & (!shiftx3x) & (!g151) & (!g162) & (!g163) & (g164)) + ((shiftx2x) & (!shiftx3x) & (!g151) & (!g162) & (g163) & (g164)) + ((shiftx2x) & (!shiftx3x) & (!g151) & (g162) & (!g163) & (g164)) + ((shiftx2x) & (!shiftx3x) & (!g151) & (g162) & (g163) & (g164)) + ((shiftx2x) & (!shiftx3x) & (g151) & (!g162) & (!g163) & (g164)) + ((shiftx2x) & (!shiftx3x) & (g151) & (!g162) & (g163) & (g164)) + ((shiftx2x) & (!shiftx3x) & (g151) & (g162) & (!g163) & (g164)) + ((shiftx2x) & (!shiftx3x) & (g151) & (g162) & (g163) & (g164)) + ((shiftx2x) & (shiftx3x) & (g151) & (!g162) & (!g163) & (!g164)) + ((shiftx2x) & (shiftx3x) & (g151) & (!g162) & (!g163) & (g164)) + ((shiftx2x) & (shiftx3x) & (g151) & (!g162) & (g163) & (!g164)) + ((shiftx2x) & (shiftx3x) & (g151) & (!g162) & (g163) & (g164)) + ((shiftx2x) & (shiftx3x) & (g151) & (g162) & (!g163) & (!g164)) + ((shiftx2x) & (shiftx3x) & (g151) & (g162) & (!g163) & (g164)) + ((shiftx2x) & (shiftx3x) & (g151) & (g162) & (g163) & (!g164)) + ((shiftx2x) & (shiftx3x) & (g151) & (g162) & (g163) & (g164)));
	assign g303 = (((!shiftx4x) & (!shiftx5x) & (!g299) & (!g300) & (g301) & (!g302)) + ((!shiftx4x) & (!shiftx5x) & (!g299) & (!g300) & (g301) & (g302)) + ((!shiftx4x) & (!shiftx5x) & (!g299) & (g300) & (g301) & (!g302)) + ((!shiftx4x) & (!shiftx5x) & (!g299) & (g300) & (g301) & (g302)) + ((!shiftx4x) & (!shiftx5x) & (g299) & (!g300) & (g301) & (!g302)) + ((!shiftx4x) & (!shiftx5x) & (g299) & (!g300) & (g301) & (g302)) + ((!shiftx4x) & (!shiftx5x) & (g299) & (g300) & (g301) & (!g302)) + ((!shiftx4x) & (!shiftx5x) & (g299) & (g300) & (g301) & (g302)) + ((!shiftx4x) & (shiftx5x) & (!g299) & (g300) & (!g301) & (!g302)) + ((!shiftx4x) & (shiftx5x) & (!g299) & (g300) & (!g301) & (g302)) + ((!shiftx4x) & (shiftx5x) & (!g299) & (g300) & (g301) & (!g302)) + ((!shiftx4x) & (shiftx5x) & (!g299) & (g300) & (g301) & (g302)) + ((!shiftx4x) & (shiftx5x) & (g299) & (g300) & (!g301) & (!g302)) + ((!shiftx4x) & (shiftx5x) & (g299) & (g300) & (!g301) & (g302)) + ((!shiftx4x) & (shiftx5x) & (g299) & (g300) & (g301) & (!g302)) + ((!shiftx4x) & (shiftx5x) & (g299) & (g300) & (g301) & (g302)) + ((shiftx4x) & (!shiftx5x) & (!g299) & (!g300) & (!g301) & (g302)) + ((shiftx4x) & (!shiftx5x) & (!g299) & (!g300) & (g301) & (g302)) + ((shiftx4x) & (!shiftx5x) & (!g299) & (g300) & (!g301) & (g302)) + ((shiftx4x) & (!shiftx5x) & (!g299) & (g300) & (g301) & (g302)) + ((shiftx4x) & (!shiftx5x) & (g299) & (!g300) & (!g301) & (g302)) + ((shiftx4x) & (!shiftx5x) & (g299) & (!g300) & (g301) & (g302)) + ((shiftx4x) & (!shiftx5x) & (g299) & (g300) & (!g301) & (g302)) + ((shiftx4x) & (!shiftx5x) & (g299) & (g300) & (g301) & (g302)) + ((shiftx4x) & (shiftx5x) & (g299) & (!g300) & (!g301) & (!g302)) + ((shiftx4x) & (shiftx5x) & (g299) & (!g300) & (!g301) & (g302)) + ((shiftx4x) & (shiftx5x) & (g299) & (!g300) & (g301) & (!g302)) + ((shiftx4x) & (shiftx5x) & (g299) & (!g300) & (g301) & (g302)) + ((shiftx4x) & (shiftx5x) & (g299) & (g300) & (!g301) & (!g302)) + ((shiftx4x) & (shiftx5x) & (g299) & (g300) & (!g301) & (g302)) + ((shiftx4x) & (shiftx5x) & (g299) & (g300) & (g301) & (!g302)) + ((shiftx4x) & (shiftx5x) & (g299) & (g300) & (g301) & (g302)));
	assign resultx15x = (((!sk[47]) & (shiftx6x) & (!g298) & (!g303)) + ((!sk[47]) & (shiftx6x) & (!g298) & (g303)) + ((!sk[47]) & (shiftx6x) & (g298) & (!g303)) + ((!sk[47]) & (shiftx6x) & (g298) & (g303)) + ((sk[47]) & (!shiftx6x) & (!g298) & (g303)) + ((sk[47]) & (!shiftx6x) & (g298) & (g303)) + ((sk[47]) & (shiftx6x) & (g298) & (!g303)) + ((sk[47]) & (shiftx6x) & (g298) & (g303)));
	assign g305 = (((!shiftx4x) & (!shiftx5x) & (!g10) & (!g15) & (!g20) & (g26)) + ((!shiftx4x) & (!shiftx5x) & (!g10) & (!g15) & (g20) & (g26)) + ((!shiftx4x) & (!shiftx5x) & (!g10) & (g15) & (!g20) & (g26)) + ((!shiftx4x) & (!shiftx5x) & (!g10) & (g15) & (g20) & (g26)) + ((!shiftx4x) & (!shiftx5x) & (g10) & (!g15) & (!g20) & (g26)) + ((!shiftx4x) & (!shiftx5x) & (g10) & (!g15) & (g20) & (g26)) + ((!shiftx4x) & (!shiftx5x) & (g10) & (g15) & (!g20) & (g26)) + ((!shiftx4x) & (!shiftx5x) & (g10) & (g15) & (g20) & (g26)) + ((!shiftx4x) & (shiftx5x) & (!g10) & (!g15) & (g20) & (!g26)) + ((!shiftx4x) & (shiftx5x) & (!g10) & (!g15) & (g20) & (g26)) + ((!shiftx4x) & (shiftx5x) & (!g10) & (g15) & (g20) & (!g26)) + ((!shiftx4x) & (shiftx5x) & (!g10) & (g15) & (g20) & (g26)) + ((!shiftx4x) & (shiftx5x) & (g10) & (!g15) & (g20) & (!g26)) + ((!shiftx4x) & (shiftx5x) & (g10) & (!g15) & (g20) & (g26)) + ((!shiftx4x) & (shiftx5x) & (g10) & (g15) & (g20) & (!g26)) + ((!shiftx4x) & (shiftx5x) & (g10) & (g15) & (g20) & (g26)) + ((shiftx4x) & (!shiftx5x) & (!g10) & (g15) & (!g20) & (!g26)) + ((shiftx4x) & (!shiftx5x) & (!g10) & (g15) & (!g20) & (g26)) + ((shiftx4x) & (!shiftx5x) & (!g10) & (g15) & (g20) & (!g26)) + ((shiftx4x) & (!shiftx5x) & (!g10) & (g15) & (g20) & (g26)) + ((shiftx4x) & (!shiftx5x) & (g10) & (g15) & (!g20) & (!g26)) + ((shiftx4x) & (!shiftx5x) & (g10) & (g15) & (!g20) & (g26)) + ((shiftx4x) & (!shiftx5x) & (g10) & (g15) & (g20) & (!g26)) + ((shiftx4x) & (!shiftx5x) & (g10) & (g15) & (g20) & (g26)) + ((shiftx4x) & (shiftx5x) & (g10) & (!g15) & (!g20) & (!g26)) + ((shiftx4x) & (shiftx5x) & (g10) & (!g15) & (!g20) & (g26)) + ((shiftx4x) & (shiftx5x) & (g10) & (!g15) & (g20) & (!g26)) + ((shiftx4x) & (shiftx5x) & (g10) & (!g15) & (g20) & (g26)) + ((shiftx4x) & (shiftx5x) & (g10) & (g15) & (!g20) & (!g26)) + ((shiftx4x) & (shiftx5x) & (g10) & (g15) & (!g20) & (g26)) + ((shiftx4x) & (shiftx5x) & (g10) & (g15) & (g20) & (!g26)) + ((shiftx4x) & (shiftx5x) & (g10) & (g15) & (g20) & (g26)));
	assign g306 = (((!shiftx4x) & (!shiftx5x) & (g5) & (!g31) & (!g36) & (!g41)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (!g31) & (!g36) & (g41)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (!g31) & (g36) & (!g41)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (!g31) & (g36) & (g41)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (g31) & (!g36) & (!g41)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (g31) & (!g36) & (g41)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (g31) & (g36) & (!g41)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (g31) & (g36) & (g41)) + ((!shiftx4x) & (shiftx5x) & (!g5) & (!g31) & (!g36) & (g41)) + ((!shiftx4x) & (shiftx5x) & (!g5) & (!g31) & (g36) & (g41)) + ((!shiftx4x) & (shiftx5x) & (!g5) & (g31) & (!g36) & (g41)) + ((!shiftx4x) & (shiftx5x) & (!g5) & (g31) & (g36) & (g41)) + ((!shiftx4x) & (shiftx5x) & (g5) & (!g31) & (!g36) & (g41)) + ((!shiftx4x) & (shiftx5x) & (g5) & (!g31) & (g36) & (g41)) + ((!shiftx4x) & (shiftx5x) & (g5) & (g31) & (!g36) & (g41)) + ((!shiftx4x) & (shiftx5x) & (g5) & (g31) & (g36) & (g41)) + ((shiftx4x) & (!shiftx5x) & (!g5) & (!g31) & (g36) & (!g41)) + ((shiftx4x) & (!shiftx5x) & (!g5) & (!g31) & (g36) & (g41)) + ((shiftx4x) & (!shiftx5x) & (!g5) & (g31) & (g36) & (!g41)) + ((shiftx4x) & (!shiftx5x) & (!g5) & (g31) & (g36) & (g41)) + ((shiftx4x) & (!shiftx5x) & (g5) & (!g31) & (g36) & (!g41)) + ((shiftx4x) & (!shiftx5x) & (g5) & (!g31) & (g36) & (g41)) + ((shiftx4x) & (!shiftx5x) & (g5) & (g31) & (g36) & (!g41)) + ((shiftx4x) & (!shiftx5x) & (g5) & (g31) & (g36) & (g41)) + ((shiftx4x) & (shiftx5x) & (!g5) & (g31) & (!g36) & (!g41)) + ((shiftx4x) & (shiftx5x) & (!g5) & (g31) & (!g36) & (g41)) + ((shiftx4x) & (shiftx5x) & (!g5) & (g31) & (g36) & (!g41)) + ((shiftx4x) & (shiftx5x) & (!g5) & (g31) & (g36) & (g41)) + ((shiftx4x) & (shiftx5x) & (g5) & (g31) & (!g36) & (!g41)) + ((shiftx4x) & (shiftx5x) & (g5) & (g31) & (!g36) & (g41)) + ((shiftx4x) & (shiftx5x) & (g5) & (g31) & (g36) & (!g41)) + ((shiftx4x) & (shiftx5x) & (g5) & (g31) & (g36) & (g41)));
	assign resultx16x = (((!shiftx6x) & (!g305) & (sk[50]) & (g306)) + ((!shiftx6x) & (g305) & (sk[50]) & (g306)) + ((shiftx6x) & (!g305) & (!sk[50]) & (!g306)) + ((shiftx6x) & (!g305) & (!sk[50]) & (g306)) + ((shiftx6x) & (g305) & (!sk[50]) & (!g306)) + ((shiftx6x) & (g305) & (!sk[50]) & (g306)) + ((shiftx6x) & (g305) & (sk[50]) & (!g306)) + ((shiftx6x) & (g305) & (sk[50]) & (g306)));
	assign g308 = (((!shiftx4x) & (!shiftx5x) & (!g48) & (!g58) & (!g63) & (g69)) + ((!shiftx4x) & (!shiftx5x) & (!g48) & (!g58) & (g63) & (g69)) + ((!shiftx4x) & (!shiftx5x) & (!g48) & (g58) & (!g63) & (g69)) + ((!shiftx4x) & (!shiftx5x) & (!g48) & (g58) & (g63) & (g69)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (!g58) & (!g63) & (g69)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (!g58) & (g63) & (g69)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (g58) & (!g63) & (g69)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (g58) & (g63) & (g69)) + ((!shiftx4x) & (shiftx5x) & (!g48) & (g58) & (!g63) & (!g69)) + ((!shiftx4x) & (shiftx5x) & (!g48) & (g58) & (!g63) & (g69)) + ((!shiftx4x) & (shiftx5x) & (!g48) & (g58) & (g63) & (!g69)) + ((!shiftx4x) & (shiftx5x) & (!g48) & (g58) & (g63) & (g69)) + ((!shiftx4x) & (shiftx5x) & (g48) & (g58) & (!g63) & (!g69)) + ((!shiftx4x) & (shiftx5x) & (g48) & (g58) & (!g63) & (g69)) + ((!shiftx4x) & (shiftx5x) & (g48) & (g58) & (g63) & (!g69)) + ((!shiftx4x) & (shiftx5x) & (g48) & (g58) & (g63) & (g69)) + ((shiftx4x) & (!shiftx5x) & (g48) & (!g58) & (!g63) & (!g69)) + ((shiftx4x) & (!shiftx5x) & (g48) & (!g58) & (!g63) & (g69)) + ((shiftx4x) & (!shiftx5x) & (g48) & (!g58) & (g63) & (!g69)) + ((shiftx4x) & (!shiftx5x) & (g48) & (!g58) & (g63) & (g69)) + ((shiftx4x) & (!shiftx5x) & (g48) & (g58) & (!g63) & (!g69)) + ((shiftx4x) & (!shiftx5x) & (g48) & (g58) & (!g63) & (g69)) + ((shiftx4x) & (!shiftx5x) & (g48) & (g58) & (g63) & (!g69)) + ((shiftx4x) & (!shiftx5x) & (g48) & (g58) & (g63) & (g69)) + ((shiftx4x) & (shiftx5x) & (!g48) & (!g58) & (g63) & (!g69)) + ((shiftx4x) & (shiftx5x) & (!g48) & (!g58) & (g63) & (g69)) + ((shiftx4x) & (shiftx5x) & (!g48) & (g58) & (g63) & (!g69)) + ((shiftx4x) & (shiftx5x) & (!g48) & (g58) & (g63) & (g69)) + ((shiftx4x) & (shiftx5x) & (g48) & (!g58) & (g63) & (!g69)) + ((shiftx4x) & (shiftx5x) & (g48) & (!g58) & (g63) & (g69)) + ((shiftx4x) & (shiftx5x) & (g48) & (g58) & (g63) & (!g69)) + ((shiftx4x) & (shiftx5x) & (g48) & (g58) & (g63) & (g69)));
	assign g309 = (((!shiftx4x) & (!shiftx5x) & (g53) & (!g74) & (!g79) & (!g84)) + ((!shiftx4x) & (!shiftx5x) & (g53) & (!g74) & (!g79) & (g84)) + ((!shiftx4x) & (!shiftx5x) & (g53) & (!g74) & (g79) & (!g84)) + ((!shiftx4x) & (!shiftx5x) & (g53) & (!g74) & (g79) & (g84)) + ((!shiftx4x) & (!shiftx5x) & (g53) & (g74) & (!g79) & (!g84)) + ((!shiftx4x) & (!shiftx5x) & (g53) & (g74) & (!g79) & (g84)) + ((!shiftx4x) & (!shiftx5x) & (g53) & (g74) & (g79) & (!g84)) + ((!shiftx4x) & (!shiftx5x) & (g53) & (g74) & (g79) & (g84)) + ((!shiftx4x) & (shiftx5x) & (!g53) & (!g74) & (!g79) & (g84)) + ((!shiftx4x) & (shiftx5x) & (!g53) & (!g74) & (g79) & (g84)) + ((!shiftx4x) & (shiftx5x) & (!g53) & (g74) & (!g79) & (g84)) + ((!shiftx4x) & (shiftx5x) & (!g53) & (g74) & (g79) & (g84)) + ((!shiftx4x) & (shiftx5x) & (g53) & (!g74) & (!g79) & (g84)) + ((!shiftx4x) & (shiftx5x) & (g53) & (!g74) & (g79) & (g84)) + ((!shiftx4x) & (shiftx5x) & (g53) & (g74) & (!g79) & (g84)) + ((!shiftx4x) & (shiftx5x) & (g53) & (g74) & (g79) & (g84)) + ((shiftx4x) & (!shiftx5x) & (!g53) & (!g74) & (g79) & (!g84)) + ((shiftx4x) & (!shiftx5x) & (!g53) & (!g74) & (g79) & (g84)) + ((shiftx4x) & (!shiftx5x) & (!g53) & (g74) & (g79) & (!g84)) + ((shiftx4x) & (!shiftx5x) & (!g53) & (g74) & (g79) & (g84)) + ((shiftx4x) & (!shiftx5x) & (g53) & (!g74) & (g79) & (!g84)) + ((shiftx4x) & (!shiftx5x) & (g53) & (!g74) & (g79) & (g84)) + ((shiftx4x) & (!shiftx5x) & (g53) & (g74) & (g79) & (!g84)) + ((shiftx4x) & (!shiftx5x) & (g53) & (g74) & (g79) & (g84)) + ((shiftx4x) & (shiftx5x) & (!g53) & (g74) & (!g79) & (!g84)) + ((shiftx4x) & (shiftx5x) & (!g53) & (g74) & (!g79) & (g84)) + ((shiftx4x) & (shiftx5x) & (!g53) & (g74) & (g79) & (!g84)) + ((shiftx4x) & (shiftx5x) & (!g53) & (g74) & (g79) & (g84)) + ((shiftx4x) & (shiftx5x) & (g53) & (g74) & (!g79) & (!g84)) + ((shiftx4x) & (shiftx5x) & (g53) & (g74) & (!g79) & (g84)) + ((shiftx4x) & (shiftx5x) & (g53) & (g74) & (g79) & (!g84)) + ((shiftx4x) & (shiftx5x) & (g53) & (g74) & (g79) & (g84)));
	assign resultx17x = (((!shiftx6x) & (sk[53]) & (!g308) & (g309)) + ((!shiftx6x) & (sk[53]) & (g308) & (g309)) + ((shiftx6x) & (!sk[53]) & (!g308) & (!g309)) + ((shiftx6x) & (!sk[53]) & (!g308) & (g309)) + ((shiftx6x) & (!sk[53]) & (g308) & (!g309)) + ((shiftx6x) & (!sk[53]) & (g308) & (g309)) + ((shiftx6x) & (sk[53]) & (g308) & (!g309)) + ((shiftx6x) & (sk[53]) & (g308) & (g309)));
	assign g311 = (((!shiftx4x) & (!shiftx5x) & (!g91) & (!g101) & (!g106) & (g112)) + ((!shiftx4x) & (!shiftx5x) & (!g91) & (!g101) & (g106) & (g112)) + ((!shiftx4x) & (!shiftx5x) & (!g91) & (g101) & (!g106) & (g112)) + ((!shiftx4x) & (!shiftx5x) & (!g91) & (g101) & (g106) & (g112)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (!g101) & (!g106) & (g112)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (!g101) & (g106) & (g112)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (g101) & (!g106) & (g112)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (g101) & (g106) & (g112)) + ((!shiftx4x) & (shiftx5x) & (!g91) & (g101) & (!g106) & (!g112)) + ((!shiftx4x) & (shiftx5x) & (!g91) & (g101) & (!g106) & (g112)) + ((!shiftx4x) & (shiftx5x) & (!g91) & (g101) & (g106) & (!g112)) + ((!shiftx4x) & (shiftx5x) & (!g91) & (g101) & (g106) & (g112)) + ((!shiftx4x) & (shiftx5x) & (g91) & (g101) & (!g106) & (!g112)) + ((!shiftx4x) & (shiftx5x) & (g91) & (g101) & (!g106) & (g112)) + ((!shiftx4x) & (shiftx5x) & (g91) & (g101) & (g106) & (!g112)) + ((!shiftx4x) & (shiftx5x) & (g91) & (g101) & (g106) & (g112)) + ((shiftx4x) & (!shiftx5x) & (g91) & (!g101) & (!g106) & (!g112)) + ((shiftx4x) & (!shiftx5x) & (g91) & (!g101) & (!g106) & (g112)) + ((shiftx4x) & (!shiftx5x) & (g91) & (!g101) & (g106) & (!g112)) + ((shiftx4x) & (!shiftx5x) & (g91) & (!g101) & (g106) & (g112)) + ((shiftx4x) & (!shiftx5x) & (g91) & (g101) & (!g106) & (!g112)) + ((shiftx4x) & (!shiftx5x) & (g91) & (g101) & (!g106) & (g112)) + ((shiftx4x) & (!shiftx5x) & (g91) & (g101) & (g106) & (!g112)) + ((shiftx4x) & (!shiftx5x) & (g91) & (g101) & (g106) & (g112)) + ((shiftx4x) & (shiftx5x) & (!g91) & (!g101) & (g106) & (!g112)) + ((shiftx4x) & (shiftx5x) & (!g91) & (!g101) & (g106) & (g112)) + ((shiftx4x) & (shiftx5x) & (!g91) & (g101) & (g106) & (!g112)) + ((shiftx4x) & (shiftx5x) & (!g91) & (g101) & (g106) & (g112)) + ((shiftx4x) & (shiftx5x) & (g91) & (!g101) & (g106) & (!g112)) + ((shiftx4x) & (shiftx5x) & (g91) & (!g101) & (g106) & (g112)) + ((shiftx4x) & (shiftx5x) & (g91) & (g101) & (g106) & (!g112)) + ((shiftx4x) & (shiftx5x) & (g91) & (g101) & (g106) & (g112)));
	assign g312 = (((!shiftx4x) & (!shiftx5x) & (g96) & (!g117) & (!g122) & (!g127)) + ((!shiftx4x) & (!shiftx5x) & (g96) & (!g117) & (!g122) & (g127)) + ((!shiftx4x) & (!shiftx5x) & (g96) & (!g117) & (g122) & (!g127)) + ((!shiftx4x) & (!shiftx5x) & (g96) & (!g117) & (g122) & (g127)) + ((!shiftx4x) & (!shiftx5x) & (g96) & (g117) & (!g122) & (!g127)) + ((!shiftx4x) & (!shiftx5x) & (g96) & (g117) & (!g122) & (g127)) + ((!shiftx4x) & (!shiftx5x) & (g96) & (g117) & (g122) & (!g127)) + ((!shiftx4x) & (!shiftx5x) & (g96) & (g117) & (g122) & (g127)) + ((!shiftx4x) & (shiftx5x) & (!g96) & (!g117) & (!g122) & (g127)) + ((!shiftx4x) & (shiftx5x) & (!g96) & (!g117) & (g122) & (g127)) + ((!shiftx4x) & (shiftx5x) & (!g96) & (g117) & (!g122) & (g127)) + ((!shiftx4x) & (shiftx5x) & (!g96) & (g117) & (g122) & (g127)) + ((!shiftx4x) & (shiftx5x) & (g96) & (!g117) & (!g122) & (g127)) + ((!shiftx4x) & (shiftx5x) & (g96) & (!g117) & (g122) & (g127)) + ((!shiftx4x) & (shiftx5x) & (g96) & (g117) & (!g122) & (g127)) + ((!shiftx4x) & (shiftx5x) & (g96) & (g117) & (g122) & (g127)) + ((shiftx4x) & (!shiftx5x) & (!g96) & (!g117) & (g122) & (!g127)) + ((shiftx4x) & (!shiftx5x) & (!g96) & (!g117) & (g122) & (g127)) + ((shiftx4x) & (!shiftx5x) & (!g96) & (g117) & (g122) & (!g127)) + ((shiftx4x) & (!shiftx5x) & (!g96) & (g117) & (g122) & (g127)) + ((shiftx4x) & (!shiftx5x) & (g96) & (!g117) & (g122) & (!g127)) + ((shiftx4x) & (!shiftx5x) & (g96) & (!g117) & (g122) & (g127)) + ((shiftx4x) & (!shiftx5x) & (g96) & (g117) & (g122) & (!g127)) + ((shiftx4x) & (!shiftx5x) & (g96) & (g117) & (g122) & (g127)) + ((shiftx4x) & (shiftx5x) & (!g96) & (g117) & (!g122) & (!g127)) + ((shiftx4x) & (shiftx5x) & (!g96) & (g117) & (!g122) & (g127)) + ((shiftx4x) & (shiftx5x) & (!g96) & (g117) & (g122) & (!g127)) + ((shiftx4x) & (shiftx5x) & (!g96) & (g117) & (g122) & (g127)) + ((shiftx4x) & (shiftx5x) & (g96) & (g117) & (!g122) & (!g127)) + ((shiftx4x) & (shiftx5x) & (g96) & (g117) & (!g122) & (g127)) + ((shiftx4x) & (shiftx5x) & (g96) & (g117) & (g122) & (!g127)) + ((shiftx4x) & (shiftx5x) & (g96) & (g117) & (g122) & (g127)));
	assign resultx18x = (((!shiftx6x) & (!g311) & (sk[56]) & (g312)) + ((!shiftx6x) & (g311) & (sk[56]) & (g312)) + ((shiftx6x) & (!g311) & (!sk[56]) & (!g312)) + ((shiftx6x) & (!g311) & (!sk[56]) & (g312)) + ((shiftx6x) & (g311) & (!sk[56]) & (!g312)) + ((shiftx6x) & (g311) & (!sk[56]) & (g312)) + ((shiftx6x) & (g311) & (sk[56]) & (!g312)) + ((shiftx6x) & (g311) & (sk[56]) & (g312)));
	assign g314 = (((!shiftx4x) & (!shiftx5x) & (!g134) & (!g139) & (!g149) & (g170)) + ((!shiftx4x) & (!shiftx5x) & (!g134) & (!g139) & (g149) & (g170)) + ((!shiftx4x) & (!shiftx5x) & (!g134) & (g139) & (!g149) & (g170)) + ((!shiftx4x) & (!shiftx5x) & (!g134) & (g139) & (g149) & (g170)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (!g139) & (!g149) & (g170)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (!g139) & (g149) & (g170)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (g139) & (!g149) & (g170)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (g139) & (g149) & (g170)) + ((!shiftx4x) & (shiftx5x) & (!g134) & (g139) & (!g149) & (!g170)) + ((!shiftx4x) & (shiftx5x) & (!g134) & (g139) & (!g149) & (g170)) + ((!shiftx4x) & (shiftx5x) & (!g134) & (g139) & (g149) & (!g170)) + ((!shiftx4x) & (shiftx5x) & (!g134) & (g139) & (g149) & (g170)) + ((!shiftx4x) & (shiftx5x) & (g134) & (g139) & (!g149) & (!g170)) + ((!shiftx4x) & (shiftx5x) & (g134) & (g139) & (!g149) & (g170)) + ((!shiftx4x) & (shiftx5x) & (g134) & (g139) & (g149) & (!g170)) + ((!shiftx4x) & (shiftx5x) & (g134) & (g139) & (g149) & (g170)) + ((shiftx4x) & (!shiftx5x) & (g134) & (!g139) & (!g149) & (!g170)) + ((shiftx4x) & (!shiftx5x) & (g134) & (!g139) & (!g149) & (g170)) + ((shiftx4x) & (!shiftx5x) & (g134) & (!g139) & (g149) & (!g170)) + ((shiftx4x) & (!shiftx5x) & (g134) & (!g139) & (g149) & (g170)) + ((shiftx4x) & (!shiftx5x) & (g134) & (g139) & (!g149) & (!g170)) + ((shiftx4x) & (!shiftx5x) & (g134) & (g139) & (!g149) & (g170)) + ((shiftx4x) & (!shiftx5x) & (g134) & (g139) & (g149) & (!g170)) + ((shiftx4x) & (!shiftx5x) & (g134) & (g139) & (g149) & (g170)) + ((shiftx4x) & (shiftx5x) & (!g134) & (!g139) & (g149) & (!g170)) + ((shiftx4x) & (shiftx5x) & (!g134) & (!g139) & (g149) & (g170)) + ((shiftx4x) & (shiftx5x) & (!g134) & (g139) & (g149) & (!g170)) + ((shiftx4x) & (shiftx5x) & (!g134) & (g139) & (g149) & (g170)) + ((shiftx4x) & (shiftx5x) & (g134) & (!g139) & (g149) & (!g170)) + ((shiftx4x) & (shiftx5x) & (g134) & (!g139) & (g149) & (g170)) + ((shiftx4x) & (shiftx5x) & (g134) & (g139) & (g149) & (!g170)) + ((shiftx4x) & (shiftx5x) & (g134) & (g139) & (g149) & (g170)));
	assign g315 = (((!shiftx4x) & (!shiftx5x) & (g144) & (!g155) & (!g160) & (!g165)) + ((!shiftx4x) & (!shiftx5x) & (g144) & (!g155) & (!g160) & (g165)) + ((!shiftx4x) & (!shiftx5x) & (g144) & (!g155) & (g160) & (!g165)) + ((!shiftx4x) & (!shiftx5x) & (g144) & (!g155) & (g160) & (g165)) + ((!shiftx4x) & (!shiftx5x) & (g144) & (g155) & (!g160) & (!g165)) + ((!shiftx4x) & (!shiftx5x) & (g144) & (g155) & (!g160) & (g165)) + ((!shiftx4x) & (!shiftx5x) & (g144) & (g155) & (g160) & (!g165)) + ((!shiftx4x) & (!shiftx5x) & (g144) & (g155) & (g160) & (g165)) + ((!shiftx4x) & (shiftx5x) & (!g144) & (g155) & (!g160) & (!g165)) + ((!shiftx4x) & (shiftx5x) & (!g144) & (g155) & (!g160) & (g165)) + ((!shiftx4x) & (shiftx5x) & (!g144) & (g155) & (g160) & (!g165)) + ((!shiftx4x) & (shiftx5x) & (!g144) & (g155) & (g160) & (g165)) + ((!shiftx4x) & (shiftx5x) & (g144) & (g155) & (!g160) & (!g165)) + ((!shiftx4x) & (shiftx5x) & (g144) & (g155) & (!g160) & (g165)) + ((!shiftx4x) & (shiftx5x) & (g144) & (g155) & (g160) & (!g165)) + ((!shiftx4x) & (shiftx5x) & (g144) & (g155) & (g160) & (g165)) + ((shiftx4x) & (!shiftx5x) & (!g144) & (!g155) & (!g160) & (g165)) + ((shiftx4x) & (!shiftx5x) & (!g144) & (!g155) & (g160) & (g165)) + ((shiftx4x) & (!shiftx5x) & (!g144) & (g155) & (!g160) & (g165)) + ((shiftx4x) & (!shiftx5x) & (!g144) & (g155) & (g160) & (g165)) + ((shiftx4x) & (!shiftx5x) & (g144) & (!g155) & (!g160) & (g165)) + ((shiftx4x) & (!shiftx5x) & (g144) & (!g155) & (g160) & (g165)) + ((shiftx4x) & (!shiftx5x) & (g144) & (g155) & (!g160) & (g165)) + ((shiftx4x) & (!shiftx5x) & (g144) & (g155) & (g160) & (g165)) + ((shiftx4x) & (shiftx5x) & (!g144) & (!g155) & (g160) & (!g165)) + ((shiftx4x) & (shiftx5x) & (!g144) & (!g155) & (g160) & (g165)) + ((shiftx4x) & (shiftx5x) & (!g144) & (g155) & (g160) & (!g165)) + ((shiftx4x) & (shiftx5x) & (!g144) & (g155) & (g160) & (g165)) + ((shiftx4x) & (shiftx5x) & (g144) & (!g155) & (g160) & (!g165)) + ((shiftx4x) & (shiftx5x) & (g144) & (!g155) & (g160) & (g165)) + ((shiftx4x) & (shiftx5x) & (g144) & (g155) & (g160) & (!g165)) + ((shiftx4x) & (shiftx5x) & (g144) & (g155) & (g160) & (g165)));
	assign resultx19x = (((!sk[59]) & (shiftx6x) & (!g314) & (!g315)) + ((!sk[59]) & (shiftx6x) & (!g314) & (g315)) + ((!sk[59]) & (shiftx6x) & (g314) & (!g315)) + ((!sk[59]) & (shiftx6x) & (g314) & (g315)) + ((sk[59]) & (!shiftx6x) & (!g314) & (g315)) + ((sk[59]) & (!shiftx6x) & (g314) & (g315)) + ((sk[59]) & (shiftx6x) & (g314) & (!g315)) + ((sk[59]) & (shiftx6x) & (g314) & (g315)));
	assign g317 = (((!shiftx4x) & (!shiftx5x) & (!g173) & (!g174) & (!g175) & (g178)) + ((!shiftx4x) & (!shiftx5x) & (!g173) & (!g174) & (g175) & (g178)) + ((!shiftx4x) & (!shiftx5x) & (!g173) & (g174) & (!g175) & (g178)) + ((!shiftx4x) & (!shiftx5x) & (!g173) & (g174) & (g175) & (g178)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (!g174) & (!g175) & (g178)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (!g174) & (g175) & (g178)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (g174) & (!g175) & (g178)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (g174) & (g175) & (g178)) + ((!shiftx4x) & (shiftx5x) & (g173) & (!g174) & (!g175) & (!g178)) + ((!shiftx4x) & (shiftx5x) & (g173) & (!g174) & (!g175) & (g178)) + ((!shiftx4x) & (shiftx5x) & (g173) & (!g174) & (g175) & (!g178)) + ((!shiftx4x) & (shiftx5x) & (g173) & (!g174) & (g175) & (g178)) + ((!shiftx4x) & (shiftx5x) & (g173) & (g174) & (!g175) & (!g178)) + ((!shiftx4x) & (shiftx5x) & (g173) & (g174) & (!g175) & (g178)) + ((!shiftx4x) & (shiftx5x) & (g173) & (g174) & (g175) & (!g178)) + ((!shiftx4x) & (shiftx5x) & (g173) & (g174) & (g175) & (g178)) + ((shiftx4x) & (!shiftx5x) & (!g173) & (g174) & (!g175) & (!g178)) + ((shiftx4x) & (!shiftx5x) & (!g173) & (g174) & (!g175) & (g178)) + ((shiftx4x) & (!shiftx5x) & (!g173) & (g174) & (g175) & (!g178)) + ((shiftx4x) & (!shiftx5x) & (!g173) & (g174) & (g175) & (g178)) + ((shiftx4x) & (!shiftx5x) & (g173) & (g174) & (!g175) & (!g178)) + ((shiftx4x) & (!shiftx5x) & (g173) & (g174) & (!g175) & (g178)) + ((shiftx4x) & (!shiftx5x) & (g173) & (g174) & (g175) & (!g178)) + ((shiftx4x) & (!shiftx5x) & (g173) & (g174) & (g175) & (g178)) + ((shiftx4x) & (shiftx5x) & (!g173) & (!g174) & (g175) & (!g178)) + ((shiftx4x) & (shiftx5x) & (!g173) & (!g174) & (g175) & (g178)) + ((shiftx4x) & (shiftx5x) & (!g173) & (g174) & (g175) & (!g178)) + ((shiftx4x) & (shiftx5x) & (!g173) & (g174) & (g175) & (g178)) + ((shiftx4x) & (shiftx5x) & (g173) & (!g174) & (g175) & (!g178)) + ((shiftx4x) & (shiftx5x) & (g173) & (!g174) & (g175) & (g178)) + ((shiftx4x) & (shiftx5x) & (g173) & (g174) & (g175) & (!g178)) + ((shiftx4x) & (shiftx5x) & (g173) & (g174) & (g175) & (g178)));
	assign g318 = (((!shiftx4x) & (!shiftx5x) & (g176) & (!g179) & (!g180) & (!g181)) + ((!shiftx4x) & (!shiftx5x) & (g176) & (!g179) & (!g180) & (g181)) + ((!shiftx4x) & (!shiftx5x) & (g176) & (!g179) & (g180) & (!g181)) + ((!shiftx4x) & (!shiftx5x) & (g176) & (!g179) & (g180) & (g181)) + ((!shiftx4x) & (!shiftx5x) & (g176) & (g179) & (!g180) & (!g181)) + ((!shiftx4x) & (!shiftx5x) & (g176) & (g179) & (!g180) & (g181)) + ((!shiftx4x) & (!shiftx5x) & (g176) & (g179) & (g180) & (!g181)) + ((!shiftx4x) & (!shiftx5x) & (g176) & (g179) & (g180) & (g181)) + ((!shiftx4x) & (shiftx5x) & (!g176) & (!g179) & (!g180) & (g181)) + ((!shiftx4x) & (shiftx5x) & (!g176) & (!g179) & (g180) & (g181)) + ((!shiftx4x) & (shiftx5x) & (!g176) & (g179) & (!g180) & (g181)) + ((!shiftx4x) & (shiftx5x) & (!g176) & (g179) & (g180) & (g181)) + ((!shiftx4x) & (shiftx5x) & (g176) & (!g179) & (!g180) & (g181)) + ((!shiftx4x) & (shiftx5x) & (g176) & (!g179) & (g180) & (g181)) + ((!shiftx4x) & (shiftx5x) & (g176) & (g179) & (!g180) & (g181)) + ((!shiftx4x) & (shiftx5x) & (g176) & (g179) & (g180) & (g181)) + ((shiftx4x) & (!shiftx5x) & (!g176) & (!g179) & (g180) & (!g181)) + ((shiftx4x) & (!shiftx5x) & (!g176) & (!g179) & (g180) & (g181)) + ((shiftx4x) & (!shiftx5x) & (!g176) & (g179) & (g180) & (!g181)) + ((shiftx4x) & (!shiftx5x) & (!g176) & (g179) & (g180) & (g181)) + ((shiftx4x) & (!shiftx5x) & (g176) & (!g179) & (g180) & (!g181)) + ((shiftx4x) & (!shiftx5x) & (g176) & (!g179) & (g180) & (g181)) + ((shiftx4x) & (!shiftx5x) & (g176) & (g179) & (g180) & (!g181)) + ((shiftx4x) & (!shiftx5x) & (g176) & (g179) & (g180) & (g181)) + ((shiftx4x) & (shiftx5x) & (!g176) & (g179) & (!g180) & (!g181)) + ((shiftx4x) & (shiftx5x) & (!g176) & (g179) & (!g180) & (g181)) + ((shiftx4x) & (shiftx5x) & (!g176) & (g179) & (g180) & (!g181)) + ((shiftx4x) & (shiftx5x) & (!g176) & (g179) & (g180) & (g181)) + ((shiftx4x) & (shiftx5x) & (g176) & (g179) & (!g180) & (!g181)) + ((shiftx4x) & (shiftx5x) & (g176) & (g179) & (!g180) & (g181)) + ((shiftx4x) & (shiftx5x) & (g176) & (g179) & (g180) & (!g181)) + ((shiftx4x) & (shiftx5x) & (g176) & (g179) & (g180) & (g181)));
	assign resultx20x = (((!shiftx6x) & (!g317) & (sk[62]) & (g318)) + ((!shiftx6x) & (g317) & (sk[62]) & (g318)) + ((shiftx6x) & (!g317) & (!sk[62]) & (!g318)) + ((shiftx6x) & (!g317) & (!sk[62]) & (g318)) + ((shiftx6x) & (g317) & (!sk[62]) & (!g318)) + ((shiftx6x) & (g317) & (!sk[62]) & (g318)) + ((shiftx6x) & (g317) & (sk[62]) & (!g318)) + ((shiftx6x) & (g317) & (sk[62]) & (g318)));
	assign g320 = (((!shiftx4x) & (!shiftx5x) & (!g184) & (!g185) & (!g186) & (g189)) + ((!shiftx4x) & (!shiftx5x) & (!g184) & (!g185) & (g186) & (g189)) + ((!shiftx4x) & (!shiftx5x) & (!g184) & (g185) & (!g186) & (g189)) + ((!shiftx4x) & (!shiftx5x) & (!g184) & (g185) & (g186) & (g189)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (!g185) & (!g186) & (g189)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (!g185) & (g186) & (g189)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (g185) & (!g186) & (g189)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (g185) & (g186) & (g189)) + ((!shiftx4x) & (shiftx5x) & (g184) & (!g185) & (!g186) & (!g189)) + ((!shiftx4x) & (shiftx5x) & (g184) & (!g185) & (!g186) & (g189)) + ((!shiftx4x) & (shiftx5x) & (g184) & (!g185) & (g186) & (!g189)) + ((!shiftx4x) & (shiftx5x) & (g184) & (!g185) & (g186) & (g189)) + ((!shiftx4x) & (shiftx5x) & (g184) & (g185) & (!g186) & (!g189)) + ((!shiftx4x) & (shiftx5x) & (g184) & (g185) & (!g186) & (g189)) + ((!shiftx4x) & (shiftx5x) & (g184) & (g185) & (g186) & (!g189)) + ((!shiftx4x) & (shiftx5x) & (g184) & (g185) & (g186) & (g189)) + ((shiftx4x) & (!shiftx5x) & (!g184) & (g185) & (!g186) & (!g189)) + ((shiftx4x) & (!shiftx5x) & (!g184) & (g185) & (!g186) & (g189)) + ((shiftx4x) & (!shiftx5x) & (!g184) & (g185) & (g186) & (!g189)) + ((shiftx4x) & (!shiftx5x) & (!g184) & (g185) & (g186) & (g189)) + ((shiftx4x) & (!shiftx5x) & (g184) & (g185) & (!g186) & (!g189)) + ((shiftx4x) & (!shiftx5x) & (g184) & (g185) & (!g186) & (g189)) + ((shiftx4x) & (!shiftx5x) & (g184) & (g185) & (g186) & (!g189)) + ((shiftx4x) & (!shiftx5x) & (g184) & (g185) & (g186) & (g189)) + ((shiftx4x) & (shiftx5x) & (!g184) & (!g185) & (g186) & (!g189)) + ((shiftx4x) & (shiftx5x) & (!g184) & (!g185) & (g186) & (g189)) + ((shiftx4x) & (shiftx5x) & (!g184) & (g185) & (g186) & (!g189)) + ((shiftx4x) & (shiftx5x) & (!g184) & (g185) & (g186) & (g189)) + ((shiftx4x) & (shiftx5x) & (g184) & (!g185) & (g186) & (!g189)) + ((shiftx4x) & (shiftx5x) & (g184) & (!g185) & (g186) & (g189)) + ((shiftx4x) & (shiftx5x) & (g184) & (g185) & (g186) & (!g189)) + ((shiftx4x) & (shiftx5x) & (g184) & (g185) & (g186) & (g189)));
	assign g321 = (((!shiftx4x) & (!shiftx5x) & (g187) & (!g190) & (!g191) & (!g192)) + ((!shiftx4x) & (!shiftx5x) & (g187) & (!g190) & (!g191) & (g192)) + ((!shiftx4x) & (!shiftx5x) & (g187) & (!g190) & (g191) & (!g192)) + ((!shiftx4x) & (!shiftx5x) & (g187) & (!g190) & (g191) & (g192)) + ((!shiftx4x) & (!shiftx5x) & (g187) & (g190) & (!g191) & (!g192)) + ((!shiftx4x) & (!shiftx5x) & (g187) & (g190) & (!g191) & (g192)) + ((!shiftx4x) & (!shiftx5x) & (g187) & (g190) & (g191) & (!g192)) + ((!shiftx4x) & (!shiftx5x) & (g187) & (g190) & (g191) & (g192)) + ((!shiftx4x) & (shiftx5x) & (!g187) & (!g190) & (!g191) & (g192)) + ((!shiftx4x) & (shiftx5x) & (!g187) & (!g190) & (g191) & (g192)) + ((!shiftx4x) & (shiftx5x) & (!g187) & (g190) & (!g191) & (g192)) + ((!shiftx4x) & (shiftx5x) & (!g187) & (g190) & (g191) & (g192)) + ((!shiftx4x) & (shiftx5x) & (g187) & (!g190) & (!g191) & (g192)) + ((!shiftx4x) & (shiftx5x) & (g187) & (!g190) & (g191) & (g192)) + ((!shiftx4x) & (shiftx5x) & (g187) & (g190) & (!g191) & (g192)) + ((!shiftx4x) & (shiftx5x) & (g187) & (g190) & (g191) & (g192)) + ((shiftx4x) & (!shiftx5x) & (!g187) & (!g190) & (g191) & (!g192)) + ((shiftx4x) & (!shiftx5x) & (!g187) & (!g190) & (g191) & (g192)) + ((shiftx4x) & (!shiftx5x) & (!g187) & (g190) & (g191) & (!g192)) + ((shiftx4x) & (!shiftx5x) & (!g187) & (g190) & (g191) & (g192)) + ((shiftx4x) & (!shiftx5x) & (g187) & (!g190) & (g191) & (!g192)) + ((shiftx4x) & (!shiftx5x) & (g187) & (!g190) & (g191) & (g192)) + ((shiftx4x) & (!shiftx5x) & (g187) & (g190) & (g191) & (!g192)) + ((shiftx4x) & (!shiftx5x) & (g187) & (g190) & (g191) & (g192)) + ((shiftx4x) & (shiftx5x) & (!g187) & (g190) & (!g191) & (!g192)) + ((shiftx4x) & (shiftx5x) & (!g187) & (g190) & (!g191) & (g192)) + ((shiftx4x) & (shiftx5x) & (!g187) & (g190) & (g191) & (!g192)) + ((shiftx4x) & (shiftx5x) & (!g187) & (g190) & (g191) & (g192)) + ((shiftx4x) & (shiftx5x) & (g187) & (g190) & (!g191) & (!g192)) + ((shiftx4x) & (shiftx5x) & (g187) & (g190) & (!g191) & (g192)) + ((shiftx4x) & (shiftx5x) & (g187) & (g190) & (g191) & (!g192)) + ((shiftx4x) & (shiftx5x) & (g187) & (g190) & (g191) & (g192)));
	assign resultx21x = (((!shiftx6x) & (!g320) & (sk[65]) & (g321)) + ((!shiftx6x) & (g320) & (sk[65]) & (g321)) + ((shiftx6x) & (!g320) & (!sk[65]) & (!g321)) + ((shiftx6x) & (!g320) & (!sk[65]) & (g321)) + ((shiftx6x) & (g320) & (!sk[65]) & (!g321)) + ((shiftx6x) & (g320) & (!sk[65]) & (g321)) + ((shiftx6x) & (g320) & (sk[65]) & (!g321)) + ((shiftx6x) & (g320) & (sk[65]) & (g321)));
	assign g323 = (((!shiftx4x) & (!shiftx5x) & (!g195) & (!g196) & (!g197) & (g200)) + ((!shiftx4x) & (!shiftx5x) & (!g195) & (!g196) & (g197) & (g200)) + ((!shiftx4x) & (!shiftx5x) & (!g195) & (g196) & (!g197) & (g200)) + ((!shiftx4x) & (!shiftx5x) & (!g195) & (g196) & (g197) & (g200)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (!g196) & (!g197) & (g200)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (!g196) & (g197) & (g200)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (g196) & (!g197) & (g200)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (g196) & (g197) & (g200)) + ((!shiftx4x) & (shiftx5x) & (g195) & (!g196) & (!g197) & (!g200)) + ((!shiftx4x) & (shiftx5x) & (g195) & (!g196) & (!g197) & (g200)) + ((!shiftx4x) & (shiftx5x) & (g195) & (!g196) & (g197) & (!g200)) + ((!shiftx4x) & (shiftx5x) & (g195) & (!g196) & (g197) & (g200)) + ((!shiftx4x) & (shiftx5x) & (g195) & (g196) & (!g197) & (!g200)) + ((!shiftx4x) & (shiftx5x) & (g195) & (g196) & (!g197) & (g200)) + ((!shiftx4x) & (shiftx5x) & (g195) & (g196) & (g197) & (!g200)) + ((!shiftx4x) & (shiftx5x) & (g195) & (g196) & (g197) & (g200)) + ((shiftx4x) & (!shiftx5x) & (!g195) & (g196) & (!g197) & (!g200)) + ((shiftx4x) & (!shiftx5x) & (!g195) & (g196) & (!g197) & (g200)) + ((shiftx4x) & (!shiftx5x) & (!g195) & (g196) & (g197) & (!g200)) + ((shiftx4x) & (!shiftx5x) & (!g195) & (g196) & (g197) & (g200)) + ((shiftx4x) & (!shiftx5x) & (g195) & (g196) & (!g197) & (!g200)) + ((shiftx4x) & (!shiftx5x) & (g195) & (g196) & (!g197) & (g200)) + ((shiftx4x) & (!shiftx5x) & (g195) & (g196) & (g197) & (!g200)) + ((shiftx4x) & (!shiftx5x) & (g195) & (g196) & (g197) & (g200)) + ((shiftx4x) & (shiftx5x) & (!g195) & (!g196) & (g197) & (!g200)) + ((shiftx4x) & (shiftx5x) & (!g195) & (!g196) & (g197) & (g200)) + ((shiftx4x) & (shiftx5x) & (!g195) & (g196) & (g197) & (!g200)) + ((shiftx4x) & (shiftx5x) & (!g195) & (g196) & (g197) & (g200)) + ((shiftx4x) & (shiftx5x) & (g195) & (!g196) & (g197) & (!g200)) + ((shiftx4x) & (shiftx5x) & (g195) & (!g196) & (g197) & (g200)) + ((shiftx4x) & (shiftx5x) & (g195) & (g196) & (g197) & (!g200)) + ((shiftx4x) & (shiftx5x) & (g195) & (g196) & (g197) & (g200)));
	assign g324 = (((!shiftx4x) & (!shiftx5x) & (g198) & (!g201) & (!g202) & (!g203)) + ((!shiftx4x) & (!shiftx5x) & (g198) & (!g201) & (!g202) & (g203)) + ((!shiftx4x) & (!shiftx5x) & (g198) & (!g201) & (g202) & (!g203)) + ((!shiftx4x) & (!shiftx5x) & (g198) & (!g201) & (g202) & (g203)) + ((!shiftx4x) & (!shiftx5x) & (g198) & (g201) & (!g202) & (!g203)) + ((!shiftx4x) & (!shiftx5x) & (g198) & (g201) & (!g202) & (g203)) + ((!shiftx4x) & (!shiftx5x) & (g198) & (g201) & (g202) & (!g203)) + ((!shiftx4x) & (!shiftx5x) & (g198) & (g201) & (g202) & (g203)) + ((!shiftx4x) & (shiftx5x) & (!g198) & (!g201) & (!g202) & (g203)) + ((!shiftx4x) & (shiftx5x) & (!g198) & (!g201) & (g202) & (g203)) + ((!shiftx4x) & (shiftx5x) & (!g198) & (g201) & (!g202) & (g203)) + ((!shiftx4x) & (shiftx5x) & (!g198) & (g201) & (g202) & (g203)) + ((!shiftx4x) & (shiftx5x) & (g198) & (!g201) & (!g202) & (g203)) + ((!shiftx4x) & (shiftx5x) & (g198) & (!g201) & (g202) & (g203)) + ((!shiftx4x) & (shiftx5x) & (g198) & (g201) & (!g202) & (g203)) + ((!shiftx4x) & (shiftx5x) & (g198) & (g201) & (g202) & (g203)) + ((shiftx4x) & (!shiftx5x) & (!g198) & (!g201) & (g202) & (!g203)) + ((shiftx4x) & (!shiftx5x) & (!g198) & (!g201) & (g202) & (g203)) + ((shiftx4x) & (!shiftx5x) & (!g198) & (g201) & (g202) & (!g203)) + ((shiftx4x) & (!shiftx5x) & (!g198) & (g201) & (g202) & (g203)) + ((shiftx4x) & (!shiftx5x) & (g198) & (!g201) & (g202) & (!g203)) + ((shiftx4x) & (!shiftx5x) & (g198) & (!g201) & (g202) & (g203)) + ((shiftx4x) & (!shiftx5x) & (g198) & (g201) & (g202) & (!g203)) + ((shiftx4x) & (!shiftx5x) & (g198) & (g201) & (g202) & (g203)) + ((shiftx4x) & (shiftx5x) & (!g198) & (g201) & (!g202) & (!g203)) + ((shiftx4x) & (shiftx5x) & (!g198) & (g201) & (!g202) & (g203)) + ((shiftx4x) & (shiftx5x) & (!g198) & (g201) & (g202) & (!g203)) + ((shiftx4x) & (shiftx5x) & (!g198) & (g201) & (g202) & (g203)) + ((shiftx4x) & (shiftx5x) & (g198) & (g201) & (!g202) & (!g203)) + ((shiftx4x) & (shiftx5x) & (g198) & (g201) & (!g202) & (g203)) + ((shiftx4x) & (shiftx5x) & (g198) & (g201) & (g202) & (!g203)) + ((shiftx4x) & (shiftx5x) & (g198) & (g201) & (g202) & (g203)));
	assign resultx22x = (((!shiftx6x) & (!g323) & (sk[68]) & (g324)) + ((!shiftx6x) & (g323) & (sk[68]) & (g324)) + ((shiftx6x) & (!g323) & (!sk[68]) & (!g324)) + ((shiftx6x) & (!g323) & (!sk[68]) & (g324)) + ((shiftx6x) & (g323) & (!sk[68]) & (!g324)) + ((shiftx6x) & (g323) & (!sk[68]) & (g324)) + ((shiftx6x) & (g323) & (sk[68]) & (!g324)) + ((shiftx6x) & (g323) & (sk[68]) & (g324)));
	assign g326 = (((!shiftx4x) & (!shiftx5x) & (!g206) & (!g207) & (!g208) & (g211)) + ((!shiftx4x) & (!shiftx5x) & (!g206) & (!g207) & (g208) & (g211)) + ((!shiftx4x) & (!shiftx5x) & (!g206) & (g207) & (!g208) & (g211)) + ((!shiftx4x) & (!shiftx5x) & (!g206) & (g207) & (g208) & (g211)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (!g207) & (!g208) & (g211)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (!g207) & (g208) & (g211)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (g207) & (!g208) & (g211)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (g207) & (g208) & (g211)) + ((!shiftx4x) & (shiftx5x) & (g206) & (!g207) & (!g208) & (!g211)) + ((!shiftx4x) & (shiftx5x) & (g206) & (!g207) & (!g208) & (g211)) + ((!shiftx4x) & (shiftx5x) & (g206) & (!g207) & (g208) & (!g211)) + ((!shiftx4x) & (shiftx5x) & (g206) & (!g207) & (g208) & (g211)) + ((!shiftx4x) & (shiftx5x) & (g206) & (g207) & (!g208) & (!g211)) + ((!shiftx4x) & (shiftx5x) & (g206) & (g207) & (!g208) & (g211)) + ((!shiftx4x) & (shiftx5x) & (g206) & (g207) & (g208) & (!g211)) + ((!shiftx4x) & (shiftx5x) & (g206) & (g207) & (g208) & (g211)) + ((shiftx4x) & (!shiftx5x) & (!g206) & (g207) & (!g208) & (!g211)) + ((shiftx4x) & (!shiftx5x) & (!g206) & (g207) & (!g208) & (g211)) + ((shiftx4x) & (!shiftx5x) & (!g206) & (g207) & (g208) & (!g211)) + ((shiftx4x) & (!shiftx5x) & (!g206) & (g207) & (g208) & (g211)) + ((shiftx4x) & (!shiftx5x) & (g206) & (g207) & (!g208) & (!g211)) + ((shiftx4x) & (!shiftx5x) & (g206) & (g207) & (!g208) & (g211)) + ((shiftx4x) & (!shiftx5x) & (g206) & (g207) & (g208) & (!g211)) + ((shiftx4x) & (!shiftx5x) & (g206) & (g207) & (g208) & (g211)) + ((shiftx4x) & (shiftx5x) & (!g206) & (!g207) & (g208) & (!g211)) + ((shiftx4x) & (shiftx5x) & (!g206) & (!g207) & (g208) & (g211)) + ((shiftx4x) & (shiftx5x) & (!g206) & (g207) & (g208) & (!g211)) + ((shiftx4x) & (shiftx5x) & (!g206) & (g207) & (g208) & (g211)) + ((shiftx4x) & (shiftx5x) & (g206) & (!g207) & (g208) & (!g211)) + ((shiftx4x) & (shiftx5x) & (g206) & (!g207) & (g208) & (g211)) + ((shiftx4x) & (shiftx5x) & (g206) & (g207) & (g208) & (!g211)) + ((shiftx4x) & (shiftx5x) & (g206) & (g207) & (g208) & (g211)));
	assign g327 = (((!shiftx4x) & (!shiftx5x) & (g209) & (!g212) & (!g213) & (!g214)) + ((!shiftx4x) & (!shiftx5x) & (g209) & (!g212) & (!g213) & (g214)) + ((!shiftx4x) & (!shiftx5x) & (g209) & (!g212) & (g213) & (!g214)) + ((!shiftx4x) & (!shiftx5x) & (g209) & (!g212) & (g213) & (g214)) + ((!shiftx4x) & (!shiftx5x) & (g209) & (g212) & (!g213) & (!g214)) + ((!shiftx4x) & (!shiftx5x) & (g209) & (g212) & (!g213) & (g214)) + ((!shiftx4x) & (!shiftx5x) & (g209) & (g212) & (g213) & (!g214)) + ((!shiftx4x) & (!shiftx5x) & (g209) & (g212) & (g213) & (g214)) + ((!shiftx4x) & (shiftx5x) & (!g209) & (!g212) & (!g213) & (g214)) + ((!shiftx4x) & (shiftx5x) & (!g209) & (!g212) & (g213) & (g214)) + ((!shiftx4x) & (shiftx5x) & (!g209) & (g212) & (!g213) & (g214)) + ((!shiftx4x) & (shiftx5x) & (!g209) & (g212) & (g213) & (g214)) + ((!shiftx4x) & (shiftx5x) & (g209) & (!g212) & (!g213) & (g214)) + ((!shiftx4x) & (shiftx5x) & (g209) & (!g212) & (g213) & (g214)) + ((!shiftx4x) & (shiftx5x) & (g209) & (g212) & (!g213) & (g214)) + ((!shiftx4x) & (shiftx5x) & (g209) & (g212) & (g213) & (g214)) + ((shiftx4x) & (!shiftx5x) & (!g209) & (!g212) & (g213) & (!g214)) + ((shiftx4x) & (!shiftx5x) & (!g209) & (!g212) & (g213) & (g214)) + ((shiftx4x) & (!shiftx5x) & (!g209) & (g212) & (g213) & (!g214)) + ((shiftx4x) & (!shiftx5x) & (!g209) & (g212) & (g213) & (g214)) + ((shiftx4x) & (!shiftx5x) & (g209) & (!g212) & (g213) & (!g214)) + ((shiftx4x) & (!shiftx5x) & (g209) & (!g212) & (g213) & (g214)) + ((shiftx4x) & (!shiftx5x) & (g209) & (g212) & (g213) & (!g214)) + ((shiftx4x) & (!shiftx5x) & (g209) & (g212) & (g213) & (g214)) + ((shiftx4x) & (shiftx5x) & (!g209) & (g212) & (!g213) & (!g214)) + ((shiftx4x) & (shiftx5x) & (!g209) & (g212) & (!g213) & (g214)) + ((shiftx4x) & (shiftx5x) & (!g209) & (g212) & (g213) & (!g214)) + ((shiftx4x) & (shiftx5x) & (!g209) & (g212) & (g213) & (g214)) + ((shiftx4x) & (shiftx5x) & (g209) & (g212) & (!g213) & (!g214)) + ((shiftx4x) & (shiftx5x) & (g209) & (g212) & (!g213) & (g214)) + ((shiftx4x) & (shiftx5x) & (g209) & (g212) & (g213) & (!g214)) + ((shiftx4x) & (shiftx5x) & (g209) & (g212) & (g213) & (g214)));
	assign resultx23x = (((!shiftx6x) & (!g326) & (sk[71]) & (g327)) + ((!shiftx6x) & (g326) & (sk[71]) & (g327)) + ((shiftx6x) & (!g326) & (!sk[71]) & (!g327)) + ((shiftx6x) & (!g326) & (!sk[71]) & (g327)) + ((shiftx6x) & (g326) & (!sk[71]) & (!g327)) + ((shiftx6x) & (g326) & (!sk[71]) & (g327)) + ((shiftx6x) & (g326) & (sk[71]) & (!g327)) + ((shiftx6x) & (g326) & (sk[71]) & (g327)));
	assign g329 = (((!shiftx4x) & (!shiftx5x) & (!g217) & (!g218) & (!g219) & (g222)) + ((!shiftx4x) & (!shiftx5x) & (!g217) & (!g218) & (g219) & (g222)) + ((!shiftx4x) & (!shiftx5x) & (!g217) & (g218) & (!g219) & (g222)) + ((!shiftx4x) & (!shiftx5x) & (!g217) & (g218) & (g219) & (g222)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (!g218) & (!g219) & (g222)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (!g218) & (g219) & (g222)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (g218) & (!g219) & (g222)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (g218) & (g219) & (g222)) + ((!shiftx4x) & (shiftx5x) & (g217) & (!g218) & (!g219) & (!g222)) + ((!shiftx4x) & (shiftx5x) & (g217) & (!g218) & (!g219) & (g222)) + ((!shiftx4x) & (shiftx5x) & (g217) & (!g218) & (g219) & (!g222)) + ((!shiftx4x) & (shiftx5x) & (g217) & (!g218) & (g219) & (g222)) + ((!shiftx4x) & (shiftx5x) & (g217) & (g218) & (!g219) & (!g222)) + ((!shiftx4x) & (shiftx5x) & (g217) & (g218) & (!g219) & (g222)) + ((!shiftx4x) & (shiftx5x) & (g217) & (g218) & (g219) & (!g222)) + ((!shiftx4x) & (shiftx5x) & (g217) & (g218) & (g219) & (g222)) + ((shiftx4x) & (!shiftx5x) & (!g217) & (g218) & (!g219) & (!g222)) + ((shiftx4x) & (!shiftx5x) & (!g217) & (g218) & (!g219) & (g222)) + ((shiftx4x) & (!shiftx5x) & (!g217) & (g218) & (g219) & (!g222)) + ((shiftx4x) & (!shiftx5x) & (!g217) & (g218) & (g219) & (g222)) + ((shiftx4x) & (!shiftx5x) & (g217) & (g218) & (!g219) & (!g222)) + ((shiftx4x) & (!shiftx5x) & (g217) & (g218) & (!g219) & (g222)) + ((shiftx4x) & (!shiftx5x) & (g217) & (g218) & (g219) & (!g222)) + ((shiftx4x) & (!shiftx5x) & (g217) & (g218) & (g219) & (g222)) + ((shiftx4x) & (shiftx5x) & (!g217) & (!g218) & (g219) & (!g222)) + ((shiftx4x) & (shiftx5x) & (!g217) & (!g218) & (g219) & (g222)) + ((shiftx4x) & (shiftx5x) & (!g217) & (g218) & (g219) & (!g222)) + ((shiftx4x) & (shiftx5x) & (!g217) & (g218) & (g219) & (g222)) + ((shiftx4x) & (shiftx5x) & (g217) & (!g218) & (g219) & (!g222)) + ((shiftx4x) & (shiftx5x) & (g217) & (!g218) & (g219) & (g222)) + ((shiftx4x) & (shiftx5x) & (g217) & (g218) & (g219) & (!g222)) + ((shiftx4x) & (shiftx5x) & (g217) & (g218) & (g219) & (g222)));
	assign g330 = (((!shiftx4x) & (!shiftx5x) & (g220) & (!g223) & (!g224) & (!g225)) + ((!shiftx4x) & (!shiftx5x) & (g220) & (!g223) & (!g224) & (g225)) + ((!shiftx4x) & (!shiftx5x) & (g220) & (!g223) & (g224) & (!g225)) + ((!shiftx4x) & (!shiftx5x) & (g220) & (!g223) & (g224) & (g225)) + ((!shiftx4x) & (!shiftx5x) & (g220) & (g223) & (!g224) & (!g225)) + ((!shiftx4x) & (!shiftx5x) & (g220) & (g223) & (!g224) & (g225)) + ((!shiftx4x) & (!shiftx5x) & (g220) & (g223) & (g224) & (!g225)) + ((!shiftx4x) & (!shiftx5x) & (g220) & (g223) & (g224) & (g225)) + ((!shiftx4x) & (shiftx5x) & (!g220) & (!g223) & (!g224) & (g225)) + ((!shiftx4x) & (shiftx5x) & (!g220) & (!g223) & (g224) & (g225)) + ((!shiftx4x) & (shiftx5x) & (!g220) & (g223) & (!g224) & (g225)) + ((!shiftx4x) & (shiftx5x) & (!g220) & (g223) & (g224) & (g225)) + ((!shiftx4x) & (shiftx5x) & (g220) & (!g223) & (!g224) & (g225)) + ((!shiftx4x) & (shiftx5x) & (g220) & (!g223) & (g224) & (g225)) + ((!shiftx4x) & (shiftx5x) & (g220) & (g223) & (!g224) & (g225)) + ((!shiftx4x) & (shiftx5x) & (g220) & (g223) & (g224) & (g225)) + ((shiftx4x) & (!shiftx5x) & (!g220) & (!g223) & (g224) & (!g225)) + ((shiftx4x) & (!shiftx5x) & (!g220) & (!g223) & (g224) & (g225)) + ((shiftx4x) & (!shiftx5x) & (!g220) & (g223) & (g224) & (!g225)) + ((shiftx4x) & (!shiftx5x) & (!g220) & (g223) & (g224) & (g225)) + ((shiftx4x) & (!shiftx5x) & (g220) & (!g223) & (g224) & (!g225)) + ((shiftx4x) & (!shiftx5x) & (g220) & (!g223) & (g224) & (g225)) + ((shiftx4x) & (!shiftx5x) & (g220) & (g223) & (g224) & (!g225)) + ((shiftx4x) & (!shiftx5x) & (g220) & (g223) & (g224) & (g225)) + ((shiftx4x) & (shiftx5x) & (!g220) & (g223) & (!g224) & (!g225)) + ((shiftx4x) & (shiftx5x) & (!g220) & (g223) & (!g224) & (g225)) + ((shiftx4x) & (shiftx5x) & (!g220) & (g223) & (g224) & (!g225)) + ((shiftx4x) & (shiftx5x) & (!g220) & (g223) & (g224) & (g225)) + ((shiftx4x) & (shiftx5x) & (g220) & (g223) & (!g224) & (!g225)) + ((shiftx4x) & (shiftx5x) & (g220) & (g223) & (!g224) & (g225)) + ((shiftx4x) & (shiftx5x) & (g220) & (g223) & (g224) & (!g225)) + ((shiftx4x) & (shiftx5x) & (g220) & (g223) & (g224) & (g225)));
	assign resultx24x = (((!shiftx6x) & (sk[74]) & (!g329) & (g330)) + ((!shiftx6x) & (sk[74]) & (g329) & (g330)) + ((shiftx6x) & (!sk[74]) & (!g329) & (!g330)) + ((shiftx6x) & (!sk[74]) & (!g329) & (g330)) + ((shiftx6x) & (!sk[74]) & (g329) & (!g330)) + ((shiftx6x) & (!sk[74]) & (g329) & (g330)) + ((shiftx6x) & (sk[74]) & (g329) & (!g330)) + ((shiftx6x) & (sk[74]) & (g329) & (g330)));
	assign g332 = (((!shiftx4x) & (!shiftx5x) & (!g228) & (!g229) & (!g230) & (g233)) + ((!shiftx4x) & (!shiftx5x) & (!g228) & (!g229) & (g230) & (g233)) + ((!shiftx4x) & (!shiftx5x) & (!g228) & (g229) & (!g230) & (g233)) + ((!shiftx4x) & (!shiftx5x) & (!g228) & (g229) & (g230) & (g233)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (!g229) & (!g230) & (g233)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (!g229) & (g230) & (g233)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (g229) & (!g230) & (g233)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (g229) & (g230) & (g233)) + ((!shiftx4x) & (shiftx5x) & (g228) & (!g229) & (!g230) & (!g233)) + ((!shiftx4x) & (shiftx5x) & (g228) & (!g229) & (!g230) & (g233)) + ((!shiftx4x) & (shiftx5x) & (g228) & (!g229) & (g230) & (!g233)) + ((!shiftx4x) & (shiftx5x) & (g228) & (!g229) & (g230) & (g233)) + ((!shiftx4x) & (shiftx5x) & (g228) & (g229) & (!g230) & (!g233)) + ((!shiftx4x) & (shiftx5x) & (g228) & (g229) & (!g230) & (g233)) + ((!shiftx4x) & (shiftx5x) & (g228) & (g229) & (g230) & (!g233)) + ((!shiftx4x) & (shiftx5x) & (g228) & (g229) & (g230) & (g233)) + ((shiftx4x) & (!shiftx5x) & (!g228) & (g229) & (!g230) & (!g233)) + ((shiftx4x) & (!shiftx5x) & (!g228) & (g229) & (!g230) & (g233)) + ((shiftx4x) & (!shiftx5x) & (!g228) & (g229) & (g230) & (!g233)) + ((shiftx4x) & (!shiftx5x) & (!g228) & (g229) & (g230) & (g233)) + ((shiftx4x) & (!shiftx5x) & (g228) & (g229) & (!g230) & (!g233)) + ((shiftx4x) & (!shiftx5x) & (g228) & (g229) & (!g230) & (g233)) + ((shiftx4x) & (!shiftx5x) & (g228) & (g229) & (g230) & (!g233)) + ((shiftx4x) & (!shiftx5x) & (g228) & (g229) & (g230) & (g233)) + ((shiftx4x) & (shiftx5x) & (!g228) & (!g229) & (g230) & (!g233)) + ((shiftx4x) & (shiftx5x) & (!g228) & (!g229) & (g230) & (g233)) + ((shiftx4x) & (shiftx5x) & (!g228) & (g229) & (g230) & (!g233)) + ((shiftx4x) & (shiftx5x) & (!g228) & (g229) & (g230) & (g233)) + ((shiftx4x) & (shiftx5x) & (g228) & (!g229) & (g230) & (!g233)) + ((shiftx4x) & (shiftx5x) & (g228) & (!g229) & (g230) & (g233)) + ((shiftx4x) & (shiftx5x) & (g228) & (g229) & (g230) & (!g233)) + ((shiftx4x) & (shiftx5x) & (g228) & (g229) & (g230) & (g233)));
	assign g333 = (((!shiftx4x) & (!shiftx5x) & (g231) & (!g234) & (!g235) & (!g236)) + ((!shiftx4x) & (!shiftx5x) & (g231) & (!g234) & (!g235) & (g236)) + ((!shiftx4x) & (!shiftx5x) & (g231) & (!g234) & (g235) & (!g236)) + ((!shiftx4x) & (!shiftx5x) & (g231) & (!g234) & (g235) & (g236)) + ((!shiftx4x) & (!shiftx5x) & (g231) & (g234) & (!g235) & (!g236)) + ((!shiftx4x) & (!shiftx5x) & (g231) & (g234) & (!g235) & (g236)) + ((!shiftx4x) & (!shiftx5x) & (g231) & (g234) & (g235) & (!g236)) + ((!shiftx4x) & (!shiftx5x) & (g231) & (g234) & (g235) & (g236)) + ((!shiftx4x) & (shiftx5x) & (!g231) & (!g234) & (!g235) & (g236)) + ((!shiftx4x) & (shiftx5x) & (!g231) & (!g234) & (g235) & (g236)) + ((!shiftx4x) & (shiftx5x) & (!g231) & (g234) & (!g235) & (g236)) + ((!shiftx4x) & (shiftx5x) & (!g231) & (g234) & (g235) & (g236)) + ((!shiftx4x) & (shiftx5x) & (g231) & (!g234) & (!g235) & (g236)) + ((!shiftx4x) & (shiftx5x) & (g231) & (!g234) & (g235) & (g236)) + ((!shiftx4x) & (shiftx5x) & (g231) & (g234) & (!g235) & (g236)) + ((!shiftx4x) & (shiftx5x) & (g231) & (g234) & (g235) & (g236)) + ((shiftx4x) & (!shiftx5x) & (!g231) & (!g234) & (g235) & (!g236)) + ((shiftx4x) & (!shiftx5x) & (!g231) & (!g234) & (g235) & (g236)) + ((shiftx4x) & (!shiftx5x) & (!g231) & (g234) & (g235) & (!g236)) + ((shiftx4x) & (!shiftx5x) & (!g231) & (g234) & (g235) & (g236)) + ((shiftx4x) & (!shiftx5x) & (g231) & (!g234) & (g235) & (!g236)) + ((shiftx4x) & (!shiftx5x) & (g231) & (!g234) & (g235) & (g236)) + ((shiftx4x) & (!shiftx5x) & (g231) & (g234) & (g235) & (!g236)) + ((shiftx4x) & (!shiftx5x) & (g231) & (g234) & (g235) & (g236)) + ((shiftx4x) & (shiftx5x) & (!g231) & (g234) & (!g235) & (!g236)) + ((shiftx4x) & (shiftx5x) & (!g231) & (g234) & (!g235) & (g236)) + ((shiftx4x) & (shiftx5x) & (!g231) & (g234) & (g235) & (!g236)) + ((shiftx4x) & (shiftx5x) & (!g231) & (g234) & (g235) & (g236)) + ((shiftx4x) & (shiftx5x) & (g231) & (g234) & (!g235) & (!g236)) + ((shiftx4x) & (shiftx5x) & (g231) & (g234) & (!g235) & (g236)) + ((shiftx4x) & (shiftx5x) & (g231) & (g234) & (g235) & (!g236)) + ((shiftx4x) & (shiftx5x) & (g231) & (g234) & (g235) & (g236)));
	assign resultx25x = (((!sk[77]) & (shiftx6x) & (!g332) & (!g333)) + ((!sk[77]) & (shiftx6x) & (!g332) & (g333)) + ((!sk[77]) & (shiftx6x) & (g332) & (!g333)) + ((!sk[77]) & (shiftx6x) & (g332) & (g333)) + ((sk[77]) & (!shiftx6x) & (!g332) & (g333)) + ((sk[77]) & (!shiftx6x) & (g332) & (g333)) + ((sk[77]) & (shiftx6x) & (g332) & (!g333)) + ((sk[77]) & (shiftx6x) & (g332) & (g333)));
	assign g335 = (((!shiftx4x) & (!shiftx5x) & (!g239) & (!g240) & (!g241) & (g244)) + ((!shiftx4x) & (!shiftx5x) & (!g239) & (!g240) & (g241) & (g244)) + ((!shiftx4x) & (!shiftx5x) & (!g239) & (g240) & (!g241) & (g244)) + ((!shiftx4x) & (!shiftx5x) & (!g239) & (g240) & (g241) & (g244)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (!g240) & (!g241) & (g244)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (!g240) & (g241) & (g244)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (g240) & (!g241) & (g244)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (g240) & (g241) & (g244)) + ((!shiftx4x) & (shiftx5x) & (g239) & (!g240) & (!g241) & (!g244)) + ((!shiftx4x) & (shiftx5x) & (g239) & (!g240) & (!g241) & (g244)) + ((!shiftx4x) & (shiftx5x) & (g239) & (!g240) & (g241) & (!g244)) + ((!shiftx4x) & (shiftx5x) & (g239) & (!g240) & (g241) & (g244)) + ((!shiftx4x) & (shiftx5x) & (g239) & (g240) & (!g241) & (!g244)) + ((!shiftx4x) & (shiftx5x) & (g239) & (g240) & (!g241) & (g244)) + ((!shiftx4x) & (shiftx5x) & (g239) & (g240) & (g241) & (!g244)) + ((!shiftx4x) & (shiftx5x) & (g239) & (g240) & (g241) & (g244)) + ((shiftx4x) & (!shiftx5x) & (!g239) & (g240) & (!g241) & (!g244)) + ((shiftx4x) & (!shiftx5x) & (!g239) & (g240) & (!g241) & (g244)) + ((shiftx4x) & (!shiftx5x) & (!g239) & (g240) & (g241) & (!g244)) + ((shiftx4x) & (!shiftx5x) & (!g239) & (g240) & (g241) & (g244)) + ((shiftx4x) & (!shiftx5x) & (g239) & (g240) & (!g241) & (!g244)) + ((shiftx4x) & (!shiftx5x) & (g239) & (g240) & (!g241) & (g244)) + ((shiftx4x) & (!shiftx5x) & (g239) & (g240) & (g241) & (!g244)) + ((shiftx4x) & (!shiftx5x) & (g239) & (g240) & (g241) & (g244)) + ((shiftx4x) & (shiftx5x) & (!g239) & (!g240) & (g241) & (!g244)) + ((shiftx4x) & (shiftx5x) & (!g239) & (!g240) & (g241) & (g244)) + ((shiftx4x) & (shiftx5x) & (!g239) & (g240) & (g241) & (!g244)) + ((shiftx4x) & (shiftx5x) & (!g239) & (g240) & (g241) & (g244)) + ((shiftx4x) & (shiftx5x) & (g239) & (!g240) & (g241) & (!g244)) + ((shiftx4x) & (shiftx5x) & (g239) & (!g240) & (g241) & (g244)) + ((shiftx4x) & (shiftx5x) & (g239) & (g240) & (g241) & (!g244)) + ((shiftx4x) & (shiftx5x) & (g239) & (g240) & (g241) & (g244)));
	assign g336 = (((!shiftx4x) & (!shiftx5x) & (g242) & (!g245) & (!g246) & (!g247)) + ((!shiftx4x) & (!shiftx5x) & (g242) & (!g245) & (!g246) & (g247)) + ((!shiftx4x) & (!shiftx5x) & (g242) & (!g245) & (g246) & (!g247)) + ((!shiftx4x) & (!shiftx5x) & (g242) & (!g245) & (g246) & (g247)) + ((!shiftx4x) & (!shiftx5x) & (g242) & (g245) & (!g246) & (!g247)) + ((!shiftx4x) & (!shiftx5x) & (g242) & (g245) & (!g246) & (g247)) + ((!shiftx4x) & (!shiftx5x) & (g242) & (g245) & (g246) & (!g247)) + ((!shiftx4x) & (!shiftx5x) & (g242) & (g245) & (g246) & (g247)) + ((!shiftx4x) & (shiftx5x) & (!g242) & (!g245) & (!g246) & (g247)) + ((!shiftx4x) & (shiftx5x) & (!g242) & (!g245) & (g246) & (g247)) + ((!shiftx4x) & (shiftx5x) & (!g242) & (g245) & (!g246) & (g247)) + ((!shiftx4x) & (shiftx5x) & (!g242) & (g245) & (g246) & (g247)) + ((!shiftx4x) & (shiftx5x) & (g242) & (!g245) & (!g246) & (g247)) + ((!shiftx4x) & (shiftx5x) & (g242) & (!g245) & (g246) & (g247)) + ((!shiftx4x) & (shiftx5x) & (g242) & (g245) & (!g246) & (g247)) + ((!shiftx4x) & (shiftx5x) & (g242) & (g245) & (g246) & (g247)) + ((shiftx4x) & (!shiftx5x) & (!g242) & (!g245) & (g246) & (!g247)) + ((shiftx4x) & (!shiftx5x) & (!g242) & (!g245) & (g246) & (g247)) + ((shiftx4x) & (!shiftx5x) & (!g242) & (g245) & (g246) & (!g247)) + ((shiftx4x) & (!shiftx5x) & (!g242) & (g245) & (g246) & (g247)) + ((shiftx4x) & (!shiftx5x) & (g242) & (!g245) & (g246) & (!g247)) + ((shiftx4x) & (!shiftx5x) & (g242) & (!g245) & (g246) & (g247)) + ((shiftx4x) & (!shiftx5x) & (g242) & (g245) & (g246) & (!g247)) + ((shiftx4x) & (!shiftx5x) & (g242) & (g245) & (g246) & (g247)) + ((shiftx4x) & (shiftx5x) & (!g242) & (g245) & (!g246) & (!g247)) + ((shiftx4x) & (shiftx5x) & (!g242) & (g245) & (!g246) & (g247)) + ((shiftx4x) & (shiftx5x) & (!g242) & (g245) & (g246) & (!g247)) + ((shiftx4x) & (shiftx5x) & (!g242) & (g245) & (g246) & (g247)) + ((shiftx4x) & (shiftx5x) & (g242) & (g245) & (!g246) & (!g247)) + ((shiftx4x) & (shiftx5x) & (g242) & (g245) & (!g246) & (g247)) + ((shiftx4x) & (shiftx5x) & (g242) & (g245) & (g246) & (!g247)) + ((shiftx4x) & (shiftx5x) & (g242) & (g245) & (g246) & (g247)));
	assign resultx26x = (((!sk[80]) & (shiftx6x) & (!g335) & (!g336)) + ((!sk[80]) & (shiftx6x) & (!g335) & (g336)) + ((!sk[80]) & (shiftx6x) & (g335) & (!g336)) + ((!sk[80]) & (shiftx6x) & (g335) & (g336)) + ((sk[80]) & (!shiftx6x) & (!g335) & (g336)) + ((sk[80]) & (!shiftx6x) & (g335) & (g336)) + ((sk[80]) & (shiftx6x) & (g335) & (!g336)) + ((sk[80]) & (shiftx6x) & (g335) & (g336)));
	assign g338 = (((!shiftx4x) & (!shiftx5x) & (!g250) & (!g251) & (!g252) & (g255)) + ((!shiftx4x) & (!shiftx5x) & (!g250) & (!g251) & (g252) & (g255)) + ((!shiftx4x) & (!shiftx5x) & (!g250) & (g251) & (!g252) & (g255)) + ((!shiftx4x) & (!shiftx5x) & (!g250) & (g251) & (g252) & (g255)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (!g251) & (!g252) & (g255)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (!g251) & (g252) & (g255)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (g251) & (!g252) & (g255)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (g251) & (g252) & (g255)) + ((!shiftx4x) & (shiftx5x) & (g250) & (!g251) & (!g252) & (!g255)) + ((!shiftx4x) & (shiftx5x) & (g250) & (!g251) & (!g252) & (g255)) + ((!shiftx4x) & (shiftx5x) & (g250) & (!g251) & (g252) & (!g255)) + ((!shiftx4x) & (shiftx5x) & (g250) & (!g251) & (g252) & (g255)) + ((!shiftx4x) & (shiftx5x) & (g250) & (g251) & (!g252) & (!g255)) + ((!shiftx4x) & (shiftx5x) & (g250) & (g251) & (!g252) & (g255)) + ((!shiftx4x) & (shiftx5x) & (g250) & (g251) & (g252) & (!g255)) + ((!shiftx4x) & (shiftx5x) & (g250) & (g251) & (g252) & (g255)) + ((shiftx4x) & (!shiftx5x) & (!g250) & (g251) & (!g252) & (!g255)) + ((shiftx4x) & (!shiftx5x) & (!g250) & (g251) & (!g252) & (g255)) + ((shiftx4x) & (!shiftx5x) & (!g250) & (g251) & (g252) & (!g255)) + ((shiftx4x) & (!shiftx5x) & (!g250) & (g251) & (g252) & (g255)) + ((shiftx4x) & (!shiftx5x) & (g250) & (g251) & (!g252) & (!g255)) + ((shiftx4x) & (!shiftx5x) & (g250) & (g251) & (!g252) & (g255)) + ((shiftx4x) & (!shiftx5x) & (g250) & (g251) & (g252) & (!g255)) + ((shiftx4x) & (!shiftx5x) & (g250) & (g251) & (g252) & (g255)) + ((shiftx4x) & (shiftx5x) & (!g250) & (!g251) & (g252) & (!g255)) + ((shiftx4x) & (shiftx5x) & (!g250) & (!g251) & (g252) & (g255)) + ((shiftx4x) & (shiftx5x) & (!g250) & (g251) & (g252) & (!g255)) + ((shiftx4x) & (shiftx5x) & (!g250) & (g251) & (g252) & (g255)) + ((shiftx4x) & (shiftx5x) & (g250) & (!g251) & (g252) & (!g255)) + ((shiftx4x) & (shiftx5x) & (g250) & (!g251) & (g252) & (g255)) + ((shiftx4x) & (shiftx5x) & (g250) & (g251) & (g252) & (!g255)) + ((shiftx4x) & (shiftx5x) & (g250) & (g251) & (g252) & (g255)));
	assign g339 = (((!shiftx4x) & (!shiftx5x) & (g253) & (!g256) & (!g257) & (!g258)) + ((!shiftx4x) & (!shiftx5x) & (g253) & (!g256) & (!g257) & (g258)) + ((!shiftx4x) & (!shiftx5x) & (g253) & (!g256) & (g257) & (!g258)) + ((!shiftx4x) & (!shiftx5x) & (g253) & (!g256) & (g257) & (g258)) + ((!shiftx4x) & (!shiftx5x) & (g253) & (g256) & (!g257) & (!g258)) + ((!shiftx4x) & (!shiftx5x) & (g253) & (g256) & (!g257) & (g258)) + ((!shiftx4x) & (!shiftx5x) & (g253) & (g256) & (g257) & (!g258)) + ((!shiftx4x) & (!shiftx5x) & (g253) & (g256) & (g257) & (g258)) + ((!shiftx4x) & (shiftx5x) & (!g253) & (!g256) & (!g257) & (g258)) + ((!shiftx4x) & (shiftx5x) & (!g253) & (!g256) & (g257) & (g258)) + ((!shiftx4x) & (shiftx5x) & (!g253) & (g256) & (!g257) & (g258)) + ((!shiftx4x) & (shiftx5x) & (!g253) & (g256) & (g257) & (g258)) + ((!shiftx4x) & (shiftx5x) & (g253) & (!g256) & (!g257) & (g258)) + ((!shiftx4x) & (shiftx5x) & (g253) & (!g256) & (g257) & (g258)) + ((!shiftx4x) & (shiftx5x) & (g253) & (g256) & (!g257) & (g258)) + ((!shiftx4x) & (shiftx5x) & (g253) & (g256) & (g257) & (g258)) + ((shiftx4x) & (!shiftx5x) & (!g253) & (!g256) & (g257) & (!g258)) + ((shiftx4x) & (!shiftx5x) & (!g253) & (!g256) & (g257) & (g258)) + ((shiftx4x) & (!shiftx5x) & (!g253) & (g256) & (g257) & (!g258)) + ((shiftx4x) & (!shiftx5x) & (!g253) & (g256) & (g257) & (g258)) + ((shiftx4x) & (!shiftx5x) & (g253) & (!g256) & (g257) & (!g258)) + ((shiftx4x) & (!shiftx5x) & (g253) & (!g256) & (g257) & (g258)) + ((shiftx4x) & (!shiftx5x) & (g253) & (g256) & (g257) & (!g258)) + ((shiftx4x) & (!shiftx5x) & (g253) & (g256) & (g257) & (g258)) + ((shiftx4x) & (shiftx5x) & (!g253) & (g256) & (!g257) & (!g258)) + ((shiftx4x) & (shiftx5x) & (!g253) & (g256) & (!g257) & (g258)) + ((shiftx4x) & (shiftx5x) & (!g253) & (g256) & (g257) & (!g258)) + ((shiftx4x) & (shiftx5x) & (!g253) & (g256) & (g257) & (g258)) + ((shiftx4x) & (shiftx5x) & (g253) & (g256) & (!g257) & (!g258)) + ((shiftx4x) & (shiftx5x) & (g253) & (g256) & (!g257) & (g258)) + ((shiftx4x) & (shiftx5x) & (g253) & (g256) & (g257) & (!g258)) + ((shiftx4x) & (shiftx5x) & (g253) & (g256) & (g257) & (g258)));
	assign resultx27x = (((!sk[83]) & (shiftx6x) & (!g338) & (!g339)) + ((!sk[83]) & (shiftx6x) & (!g338) & (g339)) + ((!sk[83]) & (shiftx6x) & (g338) & (!g339)) + ((!sk[83]) & (shiftx6x) & (g338) & (g339)) + ((sk[83]) & (!shiftx6x) & (!g338) & (g339)) + ((sk[83]) & (!shiftx6x) & (g338) & (g339)) + ((sk[83]) & (shiftx6x) & (g338) & (!g339)) + ((sk[83]) & (shiftx6x) & (g338) & (g339)));
	assign g341 = (((!shiftx4x) & (!shiftx5x) & (!g261) & (!g262) & (!g263) & (g266)) + ((!shiftx4x) & (!shiftx5x) & (!g261) & (!g262) & (g263) & (g266)) + ((!shiftx4x) & (!shiftx5x) & (!g261) & (g262) & (!g263) & (g266)) + ((!shiftx4x) & (!shiftx5x) & (!g261) & (g262) & (g263) & (g266)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (!g262) & (!g263) & (g266)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (!g262) & (g263) & (g266)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (g262) & (!g263) & (g266)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (g262) & (g263) & (g266)) + ((!shiftx4x) & (shiftx5x) & (g261) & (!g262) & (!g263) & (!g266)) + ((!shiftx4x) & (shiftx5x) & (g261) & (!g262) & (!g263) & (g266)) + ((!shiftx4x) & (shiftx5x) & (g261) & (!g262) & (g263) & (!g266)) + ((!shiftx4x) & (shiftx5x) & (g261) & (!g262) & (g263) & (g266)) + ((!shiftx4x) & (shiftx5x) & (g261) & (g262) & (!g263) & (!g266)) + ((!shiftx4x) & (shiftx5x) & (g261) & (g262) & (!g263) & (g266)) + ((!shiftx4x) & (shiftx5x) & (g261) & (g262) & (g263) & (!g266)) + ((!shiftx4x) & (shiftx5x) & (g261) & (g262) & (g263) & (g266)) + ((shiftx4x) & (!shiftx5x) & (!g261) & (g262) & (!g263) & (!g266)) + ((shiftx4x) & (!shiftx5x) & (!g261) & (g262) & (!g263) & (g266)) + ((shiftx4x) & (!shiftx5x) & (!g261) & (g262) & (g263) & (!g266)) + ((shiftx4x) & (!shiftx5x) & (!g261) & (g262) & (g263) & (g266)) + ((shiftx4x) & (!shiftx5x) & (g261) & (g262) & (!g263) & (!g266)) + ((shiftx4x) & (!shiftx5x) & (g261) & (g262) & (!g263) & (g266)) + ((shiftx4x) & (!shiftx5x) & (g261) & (g262) & (g263) & (!g266)) + ((shiftx4x) & (!shiftx5x) & (g261) & (g262) & (g263) & (g266)) + ((shiftx4x) & (shiftx5x) & (!g261) & (!g262) & (g263) & (!g266)) + ((shiftx4x) & (shiftx5x) & (!g261) & (!g262) & (g263) & (g266)) + ((shiftx4x) & (shiftx5x) & (!g261) & (g262) & (g263) & (!g266)) + ((shiftx4x) & (shiftx5x) & (!g261) & (g262) & (g263) & (g266)) + ((shiftx4x) & (shiftx5x) & (g261) & (!g262) & (g263) & (!g266)) + ((shiftx4x) & (shiftx5x) & (g261) & (!g262) & (g263) & (g266)) + ((shiftx4x) & (shiftx5x) & (g261) & (g262) & (g263) & (!g266)) + ((shiftx4x) & (shiftx5x) & (g261) & (g262) & (g263) & (g266)));
	assign g342 = (((!shiftx4x) & (!shiftx5x) & (g264) & (!g267) & (!g268) & (!g269)) + ((!shiftx4x) & (!shiftx5x) & (g264) & (!g267) & (!g268) & (g269)) + ((!shiftx4x) & (!shiftx5x) & (g264) & (!g267) & (g268) & (!g269)) + ((!shiftx4x) & (!shiftx5x) & (g264) & (!g267) & (g268) & (g269)) + ((!shiftx4x) & (!shiftx5x) & (g264) & (g267) & (!g268) & (!g269)) + ((!shiftx4x) & (!shiftx5x) & (g264) & (g267) & (!g268) & (g269)) + ((!shiftx4x) & (!shiftx5x) & (g264) & (g267) & (g268) & (!g269)) + ((!shiftx4x) & (!shiftx5x) & (g264) & (g267) & (g268) & (g269)) + ((!shiftx4x) & (shiftx5x) & (!g264) & (!g267) & (!g268) & (g269)) + ((!shiftx4x) & (shiftx5x) & (!g264) & (!g267) & (g268) & (g269)) + ((!shiftx4x) & (shiftx5x) & (!g264) & (g267) & (!g268) & (g269)) + ((!shiftx4x) & (shiftx5x) & (!g264) & (g267) & (g268) & (g269)) + ((!shiftx4x) & (shiftx5x) & (g264) & (!g267) & (!g268) & (g269)) + ((!shiftx4x) & (shiftx5x) & (g264) & (!g267) & (g268) & (g269)) + ((!shiftx4x) & (shiftx5x) & (g264) & (g267) & (!g268) & (g269)) + ((!shiftx4x) & (shiftx5x) & (g264) & (g267) & (g268) & (g269)) + ((shiftx4x) & (!shiftx5x) & (!g264) & (!g267) & (g268) & (!g269)) + ((shiftx4x) & (!shiftx5x) & (!g264) & (!g267) & (g268) & (g269)) + ((shiftx4x) & (!shiftx5x) & (!g264) & (g267) & (g268) & (!g269)) + ((shiftx4x) & (!shiftx5x) & (!g264) & (g267) & (g268) & (g269)) + ((shiftx4x) & (!shiftx5x) & (g264) & (!g267) & (g268) & (!g269)) + ((shiftx4x) & (!shiftx5x) & (g264) & (!g267) & (g268) & (g269)) + ((shiftx4x) & (!shiftx5x) & (g264) & (g267) & (g268) & (!g269)) + ((shiftx4x) & (!shiftx5x) & (g264) & (g267) & (g268) & (g269)) + ((shiftx4x) & (shiftx5x) & (!g264) & (g267) & (!g268) & (!g269)) + ((shiftx4x) & (shiftx5x) & (!g264) & (g267) & (!g268) & (g269)) + ((shiftx4x) & (shiftx5x) & (!g264) & (g267) & (g268) & (!g269)) + ((shiftx4x) & (shiftx5x) & (!g264) & (g267) & (g268) & (g269)) + ((shiftx4x) & (shiftx5x) & (g264) & (g267) & (!g268) & (!g269)) + ((shiftx4x) & (shiftx5x) & (g264) & (g267) & (!g268) & (g269)) + ((shiftx4x) & (shiftx5x) & (g264) & (g267) & (g268) & (!g269)) + ((shiftx4x) & (shiftx5x) & (g264) & (g267) & (g268) & (g269)));
	assign resultx28x = (((!sk[86]) & (shiftx6x) & (!g341) & (!g342)) + ((!sk[86]) & (shiftx6x) & (!g341) & (g342)) + ((!sk[86]) & (shiftx6x) & (g341) & (!g342)) + ((!sk[86]) & (shiftx6x) & (g341) & (g342)) + ((sk[86]) & (!shiftx6x) & (!g341) & (g342)) + ((sk[86]) & (!shiftx6x) & (g341) & (g342)) + ((sk[86]) & (shiftx6x) & (g341) & (!g342)) + ((sk[86]) & (shiftx6x) & (g341) & (g342)));
	assign g344 = (((!shiftx4x) & (!shiftx5x) & (!g272) & (!g273) & (!g274) & (g277)) + ((!shiftx4x) & (!shiftx5x) & (!g272) & (!g273) & (g274) & (g277)) + ((!shiftx4x) & (!shiftx5x) & (!g272) & (g273) & (!g274) & (g277)) + ((!shiftx4x) & (!shiftx5x) & (!g272) & (g273) & (g274) & (g277)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (!g273) & (!g274) & (g277)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (!g273) & (g274) & (g277)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (g273) & (!g274) & (g277)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (g273) & (g274) & (g277)) + ((!shiftx4x) & (shiftx5x) & (g272) & (!g273) & (!g274) & (!g277)) + ((!shiftx4x) & (shiftx5x) & (g272) & (!g273) & (!g274) & (g277)) + ((!shiftx4x) & (shiftx5x) & (g272) & (!g273) & (g274) & (!g277)) + ((!shiftx4x) & (shiftx5x) & (g272) & (!g273) & (g274) & (g277)) + ((!shiftx4x) & (shiftx5x) & (g272) & (g273) & (!g274) & (!g277)) + ((!shiftx4x) & (shiftx5x) & (g272) & (g273) & (!g274) & (g277)) + ((!shiftx4x) & (shiftx5x) & (g272) & (g273) & (g274) & (!g277)) + ((!shiftx4x) & (shiftx5x) & (g272) & (g273) & (g274) & (g277)) + ((shiftx4x) & (!shiftx5x) & (!g272) & (g273) & (!g274) & (!g277)) + ((shiftx4x) & (!shiftx5x) & (!g272) & (g273) & (!g274) & (g277)) + ((shiftx4x) & (!shiftx5x) & (!g272) & (g273) & (g274) & (!g277)) + ((shiftx4x) & (!shiftx5x) & (!g272) & (g273) & (g274) & (g277)) + ((shiftx4x) & (!shiftx5x) & (g272) & (g273) & (!g274) & (!g277)) + ((shiftx4x) & (!shiftx5x) & (g272) & (g273) & (!g274) & (g277)) + ((shiftx4x) & (!shiftx5x) & (g272) & (g273) & (g274) & (!g277)) + ((shiftx4x) & (!shiftx5x) & (g272) & (g273) & (g274) & (g277)) + ((shiftx4x) & (shiftx5x) & (!g272) & (!g273) & (g274) & (!g277)) + ((shiftx4x) & (shiftx5x) & (!g272) & (!g273) & (g274) & (g277)) + ((shiftx4x) & (shiftx5x) & (!g272) & (g273) & (g274) & (!g277)) + ((shiftx4x) & (shiftx5x) & (!g272) & (g273) & (g274) & (g277)) + ((shiftx4x) & (shiftx5x) & (g272) & (!g273) & (g274) & (!g277)) + ((shiftx4x) & (shiftx5x) & (g272) & (!g273) & (g274) & (g277)) + ((shiftx4x) & (shiftx5x) & (g272) & (g273) & (g274) & (!g277)) + ((shiftx4x) & (shiftx5x) & (g272) & (g273) & (g274) & (g277)));
	assign g345 = (((!shiftx4x) & (!shiftx5x) & (g275) & (!g278) & (!g279) & (!g280)) + ((!shiftx4x) & (!shiftx5x) & (g275) & (!g278) & (!g279) & (g280)) + ((!shiftx4x) & (!shiftx5x) & (g275) & (!g278) & (g279) & (!g280)) + ((!shiftx4x) & (!shiftx5x) & (g275) & (!g278) & (g279) & (g280)) + ((!shiftx4x) & (!shiftx5x) & (g275) & (g278) & (!g279) & (!g280)) + ((!shiftx4x) & (!shiftx5x) & (g275) & (g278) & (!g279) & (g280)) + ((!shiftx4x) & (!shiftx5x) & (g275) & (g278) & (g279) & (!g280)) + ((!shiftx4x) & (!shiftx5x) & (g275) & (g278) & (g279) & (g280)) + ((!shiftx4x) & (shiftx5x) & (!g275) & (!g278) & (!g279) & (g280)) + ((!shiftx4x) & (shiftx5x) & (!g275) & (!g278) & (g279) & (g280)) + ((!shiftx4x) & (shiftx5x) & (!g275) & (g278) & (!g279) & (g280)) + ((!shiftx4x) & (shiftx5x) & (!g275) & (g278) & (g279) & (g280)) + ((!shiftx4x) & (shiftx5x) & (g275) & (!g278) & (!g279) & (g280)) + ((!shiftx4x) & (shiftx5x) & (g275) & (!g278) & (g279) & (g280)) + ((!shiftx4x) & (shiftx5x) & (g275) & (g278) & (!g279) & (g280)) + ((!shiftx4x) & (shiftx5x) & (g275) & (g278) & (g279) & (g280)) + ((shiftx4x) & (!shiftx5x) & (!g275) & (!g278) & (g279) & (!g280)) + ((shiftx4x) & (!shiftx5x) & (!g275) & (!g278) & (g279) & (g280)) + ((shiftx4x) & (!shiftx5x) & (!g275) & (g278) & (g279) & (!g280)) + ((shiftx4x) & (!shiftx5x) & (!g275) & (g278) & (g279) & (g280)) + ((shiftx4x) & (!shiftx5x) & (g275) & (!g278) & (g279) & (!g280)) + ((shiftx4x) & (!shiftx5x) & (g275) & (!g278) & (g279) & (g280)) + ((shiftx4x) & (!shiftx5x) & (g275) & (g278) & (g279) & (!g280)) + ((shiftx4x) & (!shiftx5x) & (g275) & (g278) & (g279) & (g280)) + ((shiftx4x) & (shiftx5x) & (!g275) & (g278) & (!g279) & (!g280)) + ((shiftx4x) & (shiftx5x) & (!g275) & (g278) & (!g279) & (g280)) + ((shiftx4x) & (shiftx5x) & (!g275) & (g278) & (g279) & (!g280)) + ((shiftx4x) & (shiftx5x) & (!g275) & (g278) & (g279) & (g280)) + ((shiftx4x) & (shiftx5x) & (g275) & (g278) & (!g279) & (!g280)) + ((shiftx4x) & (shiftx5x) & (g275) & (g278) & (!g279) & (g280)) + ((shiftx4x) & (shiftx5x) & (g275) & (g278) & (g279) & (!g280)) + ((shiftx4x) & (shiftx5x) & (g275) & (g278) & (g279) & (g280)));
	assign resultx29x = (((!sk[89]) & (shiftx6x) & (!g344) & (!g345)) + ((!sk[89]) & (shiftx6x) & (!g344) & (g345)) + ((!sk[89]) & (shiftx6x) & (g344) & (!g345)) + ((!sk[89]) & (shiftx6x) & (g344) & (g345)) + ((sk[89]) & (!shiftx6x) & (!g344) & (g345)) + ((sk[89]) & (!shiftx6x) & (g344) & (g345)) + ((sk[89]) & (shiftx6x) & (g344) & (!g345)) + ((sk[89]) & (shiftx6x) & (g344) & (g345)));
	assign g347 = (((!shiftx4x) & (!shiftx5x) & (!g283) & (!g284) & (!g285) & (g288)) + ((!shiftx4x) & (!shiftx5x) & (!g283) & (!g284) & (g285) & (g288)) + ((!shiftx4x) & (!shiftx5x) & (!g283) & (g284) & (!g285) & (g288)) + ((!shiftx4x) & (!shiftx5x) & (!g283) & (g284) & (g285) & (g288)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (!g284) & (!g285) & (g288)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (!g284) & (g285) & (g288)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (g284) & (!g285) & (g288)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (g284) & (g285) & (g288)) + ((!shiftx4x) & (shiftx5x) & (g283) & (!g284) & (!g285) & (!g288)) + ((!shiftx4x) & (shiftx5x) & (g283) & (!g284) & (!g285) & (g288)) + ((!shiftx4x) & (shiftx5x) & (g283) & (!g284) & (g285) & (!g288)) + ((!shiftx4x) & (shiftx5x) & (g283) & (!g284) & (g285) & (g288)) + ((!shiftx4x) & (shiftx5x) & (g283) & (g284) & (!g285) & (!g288)) + ((!shiftx4x) & (shiftx5x) & (g283) & (g284) & (!g285) & (g288)) + ((!shiftx4x) & (shiftx5x) & (g283) & (g284) & (g285) & (!g288)) + ((!shiftx4x) & (shiftx5x) & (g283) & (g284) & (g285) & (g288)) + ((shiftx4x) & (!shiftx5x) & (!g283) & (g284) & (!g285) & (!g288)) + ((shiftx4x) & (!shiftx5x) & (!g283) & (g284) & (!g285) & (g288)) + ((shiftx4x) & (!shiftx5x) & (!g283) & (g284) & (g285) & (!g288)) + ((shiftx4x) & (!shiftx5x) & (!g283) & (g284) & (g285) & (g288)) + ((shiftx4x) & (!shiftx5x) & (g283) & (g284) & (!g285) & (!g288)) + ((shiftx4x) & (!shiftx5x) & (g283) & (g284) & (!g285) & (g288)) + ((shiftx4x) & (!shiftx5x) & (g283) & (g284) & (g285) & (!g288)) + ((shiftx4x) & (!shiftx5x) & (g283) & (g284) & (g285) & (g288)) + ((shiftx4x) & (shiftx5x) & (!g283) & (!g284) & (g285) & (!g288)) + ((shiftx4x) & (shiftx5x) & (!g283) & (!g284) & (g285) & (g288)) + ((shiftx4x) & (shiftx5x) & (!g283) & (g284) & (g285) & (!g288)) + ((shiftx4x) & (shiftx5x) & (!g283) & (g284) & (g285) & (g288)) + ((shiftx4x) & (shiftx5x) & (g283) & (!g284) & (g285) & (!g288)) + ((shiftx4x) & (shiftx5x) & (g283) & (!g284) & (g285) & (g288)) + ((shiftx4x) & (shiftx5x) & (g283) & (g284) & (g285) & (!g288)) + ((shiftx4x) & (shiftx5x) & (g283) & (g284) & (g285) & (g288)));
	assign g348 = (((!shiftx4x) & (!shiftx5x) & (g286) & (!g289) & (!g290) & (!g291)) + ((!shiftx4x) & (!shiftx5x) & (g286) & (!g289) & (!g290) & (g291)) + ((!shiftx4x) & (!shiftx5x) & (g286) & (!g289) & (g290) & (!g291)) + ((!shiftx4x) & (!shiftx5x) & (g286) & (!g289) & (g290) & (g291)) + ((!shiftx4x) & (!shiftx5x) & (g286) & (g289) & (!g290) & (!g291)) + ((!shiftx4x) & (!shiftx5x) & (g286) & (g289) & (!g290) & (g291)) + ((!shiftx4x) & (!shiftx5x) & (g286) & (g289) & (g290) & (!g291)) + ((!shiftx4x) & (!shiftx5x) & (g286) & (g289) & (g290) & (g291)) + ((!shiftx4x) & (shiftx5x) & (!g286) & (!g289) & (!g290) & (g291)) + ((!shiftx4x) & (shiftx5x) & (!g286) & (!g289) & (g290) & (g291)) + ((!shiftx4x) & (shiftx5x) & (!g286) & (g289) & (!g290) & (g291)) + ((!shiftx4x) & (shiftx5x) & (!g286) & (g289) & (g290) & (g291)) + ((!shiftx4x) & (shiftx5x) & (g286) & (!g289) & (!g290) & (g291)) + ((!shiftx4x) & (shiftx5x) & (g286) & (!g289) & (g290) & (g291)) + ((!shiftx4x) & (shiftx5x) & (g286) & (g289) & (!g290) & (g291)) + ((!shiftx4x) & (shiftx5x) & (g286) & (g289) & (g290) & (g291)) + ((shiftx4x) & (!shiftx5x) & (!g286) & (!g289) & (g290) & (!g291)) + ((shiftx4x) & (!shiftx5x) & (!g286) & (!g289) & (g290) & (g291)) + ((shiftx4x) & (!shiftx5x) & (!g286) & (g289) & (g290) & (!g291)) + ((shiftx4x) & (!shiftx5x) & (!g286) & (g289) & (g290) & (g291)) + ((shiftx4x) & (!shiftx5x) & (g286) & (!g289) & (g290) & (!g291)) + ((shiftx4x) & (!shiftx5x) & (g286) & (!g289) & (g290) & (g291)) + ((shiftx4x) & (!shiftx5x) & (g286) & (g289) & (g290) & (!g291)) + ((shiftx4x) & (!shiftx5x) & (g286) & (g289) & (g290) & (g291)) + ((shiftx4x) & (shiftx5x) & (!g286) & (g289) & (!g290) & (!g291)) + ((shiftx4x) & (shiftx5x) & (!g286) & (g289) & (!g290) & (g291)) + ((shiftx4x) & (shiftx5x) & (!g286) & (g289) & (g290) & (!g291)) + ((shiftx4x) & (shiftx5x) & (!g286) & (g289) & (g290) & (g291)) + ((shiftx4x) & (shiftx5x) & (g286) & (g289) & (!g290) & (!g291)) + ((shiftx4x) & (shiftx5x) & (g286) & (g289) & (!g290) & (g291)) + ((shiftx4x) & (shiftx5x) & (g286) & (g289) & (g290) & (!g291)) + ((shiftx4x) & (shiftx5x) & (g286) & (g289) & (g290) & (g291)));
	assign resultx30x = (((!sk[92]) & (shiftx6x) & (!g347) & (!g348)) + ((!sk[92]) & (shiftx6x) & (!g347) & (g348)) + ((!sk[92]) & (shiftx6x) & (g347) & (!g348)) + ((!sk[92]) & (shiftx6x) & (g347) & (g348)) + ((sk[92]) & (!shiftx6x) & (!g347) & (g348)) + ((sk[92]) & (!shiftx6x) & (g347) & (g348)) + ((sk[92]) & (shiftx6x) & (g347) & (!g348)) + ((sk[92]) & (shiftx6x) & (g347) & (g348)));
	assign g350 = (((!shiftx4x) & (!shiftx5x) & (!g294) & (!g295) & (!g296) & (g299)) + ((!shiftx4x) & (!shiftx5x) & (!g294) & (!g295) & (g296) & (g299)) + ((!shiftx4x) & (!shiftx5x) & (!g294) & (g295) & (!g296) & (g299)) + ((!shiftx4x) & (!shiftx5x) & (!g294) & (g295) & (g296) & (g299)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (!g295) & (!g296) & (g299)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (!g295) & (g296) & (g299)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (g295) & (!g296) & (g299)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (g295) & (g296) & (g299)) + ((!shiftx4x) & (shiftx5x) & (g294) & (!g295) & (!g296) & (!g299)) + ((!shiftx4x) & (shiftx5x) & (g294) & (!g295) & (!g296) & (g299)) + ((!shiftx4x) & (shiftx5x) & (g294) & (!g295) & (g296) & (!g299)) + ((!shiftx4x) & (shiftx5x) & (g294) & (!g295) & (g296) & (g299)) + ((!shiftx4x) & (shiftx5x) & (g294) & (g295) & (!g296) & (!g299)) + ((!shiftx4x) & (shiftx5x) & (g294) & (g295) & (!g296) & (g299)) + ((!shiftx4x) & (shiftx5x) & (g294) & (g295) & (g296) & (!g299)) + ((!shiftx4x) & (shiftx5x) & (g294) & (g295) & (g296) & (g299)) + ((shiftx4x) & (!shiftx5x) & (!g294) & (g295) & (!g296) & (!g299)) + ((shiftx4x) & (!shiftx5x) & (!g294) & (g295) & (!g296) & (g299)) + ((shiftx4x) & (!shiftx5x) & (!g294) & (g295) & (g296) & (!g299)) + ((shiftx4x) & (!shiftx5x) & (!g294) & (g295) & (g296) & (g299)) + ((shiftx4x) & (!shiftx5x) & (g294) & (g295) & (!g296) & (!g299)) + ((shiftx4x) & (!shiftx5x) & (g294) & (g295) & (!g296) & (g299)) + ((shiftx4x) & (!shiftx5x) & (g294) & (g295) & (g296) & (!g299)) + ((shiftx4x) & (!shiftx5x) & (g294) & (g295) & (g296) & (g299)) + ((shiftx4x) & (shiftx5x) & (!g294) & (!g295) & (g296) & (!g299)) + ((shiftx4x) & (shiftx5x) & (!g294) & (!g295) & (g296) & (g299)) + ((shiftx4x) & (shiftx5x) & (!g294) & (g295) & (g296) & (!g299)) + ((shiftx4x) & (shiftx5x) & (!g294) & (g295) & (g296) & (g299)) + ((shiftx4x) & (shiftx5x) & (g294) & (!g295) & (g296) & (!g299)) + ((shiftx4x) & (shiftx5x) & (g294) & (!g295) & (g296) & (g299)) + ((shiftx4x) & (shiftx5x) & (g294) & (g295) & (g296) & (!g299)) + ((shiftx4x) & (shiftx5x) & (g294) & (g295) & (g296) & (g299)));
	assign g351 = (((!shiftx4x) & (!shiftx5x) & (g297) & (!g300) & (!g301) & (!g302)) + ((!shiftx4x) & (!shiftx5x) & (g297) & (!g300) & (!g301) & (g302)) + ((!shiftx4x) & (!shiftx5x) & (g297) & (!g300) & (g301) & (!g302)) + ((!shiftx4x) & (!shiftx5x) & (g297) & (!g300) & (g301) & (g302)) + ((!shiftx4x) & (!shiftx5x) & (g297) & (g300) & (!g301) & (!g302)) + ((!shiftx4x) & (!shiftx5x) & (g297) & (g300) & (!g301) & (g302)) + ((!shiftx4x) & (!shiftx5x) & (g297) & (g300) & (g301) & (!g302)) + ((!shiftx4x) & (!shiftx5x) & (g297) & (g300) & (g301) & (g302)) + ((!shiftx4x) & (shiftx5x) & (!g297) & (!g300) & (!g301) & (g302)) + ((!shiftx4x) & (shiftx5x) & (!g297) & (!g300) & (g301) & (g302)) + ((!shiftx4x) & (shiftx5x) & (!g297) & (g300) & (!g301) & (g302)) + ((!shiftx4x) & (shiftx5x) & (!g297) & (g300) & (g301) & (g302)) + ((!shiftx4x) & (shiftx5x) & (g297) & (!g300) & (!g301) & (g302)) + ((!shiftx4x) & (shiftx5x) & (g297) & (!g300) & (g301) & (g302)) + ((!shiftx4x) & (shiftx5x) & (g297) & (g300) & (!g301) & (g302)) + ((!shiftx4x) & (shiftx5x) & (g297) & (g300) & (g301) & (g302)) + ((shiftx4x) & (!shiftx5x) & (!g297) & (!g300) & (g301) & (!g302)) + ((shiftx4x) & (!shiftx5x) & (!g297) & (!g300) & (g301) & (g302)) + ((shiftx4x) & (!shiftx5x) & (!g297) & (g300) & (g301) & (!g302)) + ((shiftx4x) & (!shiftx5x) & (!g297) & (g300) & (g301) & (g302)) + ((shiftx4x) & (!shiftx5x) & (g297) & (!g300) & (g301) & (!g302)) + ((shiftx4x) & (!shiftx5x) & (g297) & (!g300) & (g301) & (g302)) + ((shiftx4x) & (!shiftx5x) & (g297) & (g300) & (g301) & (!g302)) + ((shiftx4x) & (!shiftx5x) & (g297) & (g300) & (g301) & (g302)) + ((shiftx4x) & (shiftx5x) & (!g297) & (g300) & (!g301) & (!g302)) + ((shiftx4x) & (shiftx5x) & (!g297) & (g300) & (!g301) & (g302)) + ((shiftx4x) & (shiftx5x) & (!g297) & (g300) & (g301) & (!g302)) + ((shiftx4x) & (shiftx5x) & (!g297) & (g300) & (g301) & (g302)) + ((shiftx4x) & (shiftx5x) & (g297) & (g300) & (!g301) & (!g302)) + ((shiftx4x) & (shiftx5x) & (g297) & (g300) & (!g301) & (g302)) + ((shiftx4x) & (shiftx5x) & (g297) & (g300) & (g301) & (!g302)) + ((shiftx4x) & (shiftx5x) & (g297) & (g300) & (g301) & (g302)));
	assign resultx31x = (((!shiftx6x) & (!g350) & (sk[95]) & (g351)) + ((!shiftx6x) & (g350) & (sk[95]) & (g351)) + ((shiftx6x) & (!g350) & (!sk[95]) & (!g351)) + ((shiftx6x) & (!g350) & (!sk[95]) & (g351)) + ((shiftx6x) & (g350) & (!sk[95]) & (!g351)) + ((shiftx6x) & (g350) & (!sk[95]) & (g351)) + ((shiftx6x) & (g350) & (sk[95]) & (!g351)) + ((shiftx6x) & (g350) & (sk[95]) & (g351)));
	assign g353 = (((!shiftx4x) & (!shiftx5x) & (!g15) & (!g20) & (!g26) & (g31)) + ((!shiftx4x) & (!shiftx5x) & (!g15) & (!g20) & (g26) & (g31)) + ((!shiftx4x) & (!shiftx5x) & (!g15) & (g20) & (!g26) & (g31)) + ((!shiftx4x) & (!shiftx5x) & (!g15) & (g20) & (g26) & (g31)) + ((!shiftx4x) & (!shiftx5x) & (g15) & (!g20) & (!g26) & (g31)) + ((!shiftx4x) & (!shiftx5x) & (g15) & (!g20) & (g26) & (g31)) + ((!shiftx4x) & (!shiftx5x) & (g15) & (g20) & (!g26) & (g31)) + ((!shiftx4x) & (!shiftx5x) & (g15) & (g20) & (g26) & (g31)) + ((!shiftx4x) & (shiftx5x) & (g15) & (!g20) & (!g26) & (!g31)) + ((!shiftx4x) & (shiftx5x) & (g15) & (!g20) & (!g26) & (g31)) + ((!shiftx4x) & (shiftx5x) & (g15) & (!g20) & (g26) & (!g31)) + ((!shiftx4x) & (shiftx5x) & (g15) & (!g20) & (g26) & (g31)) + ((!shiftx4x) & (shiftx5x) & (g15) & (g20) & (!g26) & (!g31)) + ((!shiftx4x) & (shiftx5x) & (g15) & (g20) & (!g26) & (g31)) + ((!shiftx4x) & (shiftx5x) & (g15) & (g20) & (g26) & (!g31)) + ((!shiftx4x) & (shiftx5x) & (g15) & (g20) & (g26) & (g31)) + ((shiftx4x) & (!shiftx5x) & (!g15) & (!g20) & (g26) & (!g31)) + ((shiftx4x) & (!shiftx5x) & (!g15) & (!g20) & (g26) & (g31)) + ((shiftx4x) & (!shiftx5x) & (!g15) & (g20) & (g26) & (!g31)) + ((shiftx4x) & (!shiftx5x) & (!g15) & (g20) & (g26) & (g31)) + ((shiftx4x) & (!shiftx5x) & (g15) & (!g20) & (g26) & (!g31)) + ((shiftx4x) & (!shiftx5x) & (g15) & (!g20) & (g26) & (g31)) + ((shiftx4x) & (!shiftx5x) & (g15) & (g20) & (g26) & (!g31)) + ((shiftx4x) & (!shiftx5x) & (g15) & (g20) & (g26) & (g31)) + ((shiftx4x) & (shiftx5x) & (!g15) & (g20) & (!g26) & (!g31)) + ((shiftx4x) & (shiftx5x) & (!g15) & (g20) & (!g26) & (g31)) + ((shiftx4x) & (shiftx5x) & (!g15) & (g20) & (g26) & (!g31)) + ((shiftx4x) & (shiftx5x) & (!g15) & (g20) & (g26) & (g31)) + ((shiftx4x) & (shiftx5x) & (g15) & (g20) & (!g26) & (!g31)) + ((shiftx4x) & (shiftx5x) & (g15) & (g20) & (!g26) & (g31)) + ((shiftx4x) & (shiftx5x) & (g15) & (g20) & (g26) & (!g31)) + ((shiftx4x) & (shiftx5x) & (g15) & (g20) & (g26) & (g31)));
	assign g354 = (((!shiftx4x) & (!shiftx5x) & (!g5) & (g10) & (!g36) & (!g41)) + ((!shiftx4x) & (!shiftx5x) & (!g5) & (g10) & (!g36) & (g41)) + ((!shiftx4x) & (!shiftx5x) & (!g5) & (g10) & (g36) & (!g41)) + ((!shiftx4x) & (!shiftx5x) & (!g5) & (g10) & (g36) & (g41)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (g10) & (!g36) & (!g41)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (g10) & (!g36) & (g41)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (g10) & (g36) & (!g41)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (g10) & (g36) & (g41)) + ((!shiftx4x) & (shiftx5x) & (!g5) & (!g10) & (g36) & (!g41)) + ((!shiftx4x) & (shiftx5x) & (!g5) & (!g10) & (g36) & (g41)) + ((!shiftx4x) & (shiftx5x) & (!g5) & (g10) & (g36) & (!g41)) + ((!shiftx4x) & (shiftx5x) & (!g5) & (g10) & (g36) & (g41)) + ((!shiftx4x) & (shiftx5x) & (g5) & (!g10) & (g36) & (!g41)) + ((!shiftx4x) & (shiftx5x) & (g5) & (!g10) & (g36) & (g41)) + ((!shiftx4x) & (shiftx5x) & (g5) & (g10) & (g36) & (!g41)) + ((!shiftx4x) & (shiftx5x) & (g5) & (g10) & (g36) & (g41)) + ((shiftx4x) & (!shiftx5x) & (g5) & (!g10) & (!g36) & (!g41)) + ((shiftx4x) & (!shiftx5x) & (g5) & (!g10) & (!g36) & (g41)) + ((shiftx4x) & (!shiftx5x) & (g5) & (!g10) & (g36) & (!g41)) + ((shiftx4x) & (!shiftx5x) & (g5) & (!g10) & (g36) & (g41)) + ((shiftx4x) & (!shiftx5x) & (g5) & (g10) & (!g36) & (!g41)) + ((shiftx4x) & (!shiftx5x) & (g5) & (g10) & (!g36) & (g41)) + ((shiftx4x) & (!shiftx5x) & (g5) & (g10) & (g36) & (!g41)) + ((shiftx4x) & (!shiftx5x) & (g5) & (g10) & (g36) & (g41)) + ((shiftx4x) & (shiftx5x) & (!g5) & (!g10) & (!g36) & (g41)) + ((shiftx4x) & (shiftx5x) & (!g5) & (!g10) & (g36) & (g41)) + ((shiftx4x) & (shiftx5x) & (!g5) & (g10) & (!g36) & (g41)) + ((shiftx4x) & (shiftx5x) & (!g5) & (g10) & (g36) & (g41)) + ((shiftx4x) & (shiftx5x) & (g5) & (!g10) & (!g36) & (g41)) + ((shiftx4x) & (shiftx5x) & (g5) & (!g10) & (g36) & (g41)) + ((shiftx4x) & (shiftx5x) & (g5) & (g10) & (!g36) & (g41)) + ((shiftx4x) & (shiftx5x) & (g5) & (g10) & (g36) & (g41)));
	assign resultx32x = (((!shiftx6x) & (sk[98]) & (!g353) & (g354)) + ((!shiftx6x) & (sk[98]) & (g353) & (g354)) + ((shiftx6x) & (!sk[98]) & (!g353) & (!g354)) + ((shiftx6x) & (!sk[98]) & (!g353) & (g354)) + ((shiftx6x) & (!sk[98]) & (g353) & (!g354)) + ((shiftx6x) & (!sk[98]) & (g353) & (g354)) + ((shiftx6x) & (sk[98]) & (g353) & (!g354)) + ((shiftx6x) & (sk[98]) & (g353) & (g354)));
	assign g356 = (((!shiftx4x) & (!shiftx5x) & (!g48) & (!g58) & (!g69) & (g74)) + ((!shiftx4x) & (!shiftx5x) & (!g48) & (!g58) & (g69) & (g74)) + ((!shiftx4x) & (!shiftx5x) & (!g48) & (g58) & (!g69) & (g74)) + ((!shiftx4x) & (!shiftx5x) & (!g48) & (g58) & (g69) & (g74)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (!g58) & (!g69) & (g74)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (!g58) & (g69) & (g74)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (g58) & (!g69) & (g74)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (g58) & (g69) & (g74)) + ((!shiftx4x) & (shiftx5x) & (g48) & (!g58) & (!g69) & (!g74)) + ((!shiftx4x) & (shiftx5x) & (g48) & (!g58) & (!g69) & (g74)) + ((!shiftx4x) & (shiftx5x) & (g48) & (!g58) & (g69) & (!g74)) + ((!shiftx4x) & (shiftx5x) & (g48) & (!g58) & (g69) & (g74)) + ((!shiftx4x) & (shiftx5x) & (g48) & (g58) & (!g69) & (!g74)) + ((!shiftx4x) & (shiftx5x) & (g48) & (g58) & (!g69) & (g74)) + ((!shiftx4x) & (shiftx5x) & (g48) & (g58) & (g69) & (!g74)) + ((!shiftx4x) & (shiftx5x) & (g48) & (g58) & (g69) & (g74)) + ((shiftx4x) & (!shiftx5x) & (!g48) & (!g58) & (g69) & (!g74)) + ((shiftx4x) & (!shiftx5x) & (!g48) & (!g58) & (g69) & (g74)) + ((shiftx4x) & (!shiftx5x) & (!g48) & (g58) & (g69) & (!g74)) + ((shiftx4x) & (!shiftx5x) & (!g48) & (g58) & (g69) & (g74)) + ((shiftx4x) & (!shiftx5x) & (g48) & (!g58) & (g69) & (!g74)) + ((shiftx4x) & (!shiftx5x) & (g48) & (!g58) & (g69) & (g74)) + ((shiftx4x) & (!shiftx5x) & (g48) & (g58) & (g69) & (!g74)) + ((shiftx4x) & (!shiftx5x) & (g48) & (g58) & (g69) & (g74)) + ((shiftx4x) & (shiftx5x) & (!g48) & (g58) & (!g69) & (!g74)) + ((shiftx4x) & (shiftx5x) & (!g48) & (g58) & (!g69) & (g74)) + ((shiftx4x) & (shiftx5x) & (!g48) & (g58) & (g69) & (!g74)) + ((shiftx4x) & (shiftx5x) & (!g48) & (g58) & (g69) & (g74)) + ((shiftx4x) & (shiftx5x) & (g48) & (g58) & (!g69) & (!g74)) + ((shiftx4x) & (shiftx5x) & (g48) & (g58) & (!g69) & (g74)) + ((shiftx4x) & (shiftx5x) & (g48) & (g58) & (g69) & (!g74)) + ((shiftx4x) & (shiftx5x) & (g48) & (g58) & (g69) & (g74)));
	assign g357 = (((!shiftx4x) & (!shiftx5x) & (!g53) & (g63) & (!g79) & (!g84)) + ((!shiftx4x) & (!shiftx5x) & (!g53) & (g63) & (!g79) & (g84)) + ((!shiftx4x) & (!shiftx5x) & (!g53) & (g63) & (g79) & (!g84)) + ((!shiftx4x) & (!shiftx5x) & (!g53) & (g63) & (g79) & (g84)) + ((!shiftx4x) & (!shiftx5x) & (g53) & (g63) & (!g79) & (!g84)) + ((!shiftx4x) & (!shiftx5x) & (g53) & (g63) & (!g79) & (g84)) + ((!shiftx4x) & (!shiftx5x) & (g53) & (g63) & (g79) & (!g84)) + ((!shiftx4x) & (!shiftx5x) & (g53) & (g63) & (g79) & (g84)) + ((!shiftx4x) & (shiftx5x) & (!g53) & (!g63) & (g79) & (!g84)) + ((!shiftx4x) & (shiftx5x) & (!g53) & (!g63) & (g79) & (g84)) + ((!shiftx4x) & (shiftx5x) & (!g53) & (g63) & (g79) & (!g84)) + ((!shiftx4x) & (shiftx5x) & (!g53) & (g63) & (g79) & (g84)) + ((!shiftx4x) & (shiftx5x) & (g53) & (!g63) & (g79) & (!g84)) + ((!shiftx4x) & (shiftx5x) & (g53) & (!g63) & (g79) & (g84)) + ((!shiftx4x) & (shiftx5x) & (g53) & (g63) & (g79) & (!g84)) + ((!shiftx4x) & (shiftx5x) & (g53) & (g63) & (g79) & (g84)) + ((shiftx4x) & (!shiftx5x) & (g53) & (!g63) & (!g79) & (!g84)) + ((shiftx4x) & (!shiftx5x) & (g53) & (!g63) & (!g79) & (g84)) + ((shiftx4x) & (!shiftx5x) & (g53) & (!g63) & (g79) & (!g84)) + ((shiftx4x) & (!shiftx5x) & (g53) & (!g63) & (g79) & (g84)) + ((shiftx4x) & (!shiftx5x) & (g53) & (g63) & (!g79) & (!g84)) + ((shiftx4x) & (!shiftx5x) & (g53) & (g63) & (!g79) & (g84)) + ((shiftx4x) & (!shiftx5x) & (g53) & (g63) & (g79) & (!g84)) + ((shiftx4x) & (!shiftx5x) & (g53) & (g63) & (g79) & (g84)) + ((shiftx4x) & (shiftx5x) & (!g53) & (!g63) & (!g79) & (g84)) + ((shiftx4x) & (shiftx5x) & (!g53) & (!g63) & (g79) & (g84)) + ((shiftx4x) & (shiftx5x) & (!g53) & (g63) & (!g79) & (g84)) + ((shiftx4x) & (shiftx5x) & (!g53) & (g63) & (g79) & (g84)) + ((shiftx4x) & (shiftx5x) & (g53) & (!g63) & (!g79) & (g84)) + ((shiftx4x) & (shiftx5x) & (g53) & (!g63) & (g79) & (g84)) + ((shiftx4x) & (shiftx5x) & (g53) & (g63) & (!g79) & (g84)) + ((shiftx4x) & (shiftx5x) & (g53) & (g63) & (g79) & (g84)));
	assign resultx33x = (((!shiftx6x) & (sk[101]) & (!g356) & (g357)) + ((!shiftx6x) & (sk[101]) & (g356) & (g357)) + ((shiftx6x) & (!sk[101]) & (!g356) & (!g357)) + ((shiftx6x) & (!sk[101]) & (!g356) & (g357)) + ((shiftx6x) & (!sk[101]) & (g356) & (!g357)) + ((shiftx6x) & (!sk[101]) & (g356) & (g357)) + ((shiftx6x) & (sk[101]) & (g356) & (!g357)) + ((shiftx6x) & (sk[101]) & (g356) & (g357)));
	assign g359 = (((!shiftx4x) & (!shiftx5x) & (!g91) & (!g101) & (!g112) & (g117)) + ((!shiftx4x) & (!shiftx5x) & (!g91) & (!g101) & (g112) & (g117)) + ((!shiftx4x) & (!shiftx5x) & (!g91) & (g101) & (!g112) & (g117)) + ((!shiftx4x) & (!shiftx5x) & (!g91) & (g101) & (g112) & (g117)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (!g101) & (!g112) & (g117)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (!g101) & (g112) & (g117)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (g101) & (!g112) & (g117)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (g101) & (g112) & (g117)) + ((!shiftx4x) & (shiftx5x) & (g91) & (!g101) & (!g112) & (!g117)) + ((!shiftx4x) & (shiftx5x) & (g91) & (!g101) & (!g112) & (g117)) + ((!shiftx4x) & (shiftx5x) & (g91) & (!g101) & (g112) & (!g117)) + ((!shiftx4x) & (shiftx5x) & (g91) & (!g101) & (g112) & (g117)) + ((!shiftx4x) & (shiftx5x) & (g91) & (g101) & (!g112) & (!g117)) + ((!shiftx4x) & (shiftx5x) & (g91) & (g101) & (!g112) & (g117)) + ((!shiftx4x) & (shiftx5x) & (g91) & (g101) & (g112) & (!g117)) + ((!shiftx4x) & (shiftx5x) & (g91) & (g101) & (g112) & (g117)) + ((shiftx4x) & (!shiftx5x) & (!g91) & (!g101) & (g112) & (!g117)) + ((shiftx4x) & (!shiftx5x) & (!g91) & (!g101) & (g112) & (g117)) + ((shiftx4x) & (!shiftx5x) & (!g91) & (g101) & (g112) & (!g117)) + ((shiftx4x) & (!shiftx5x) & (!g91) & (g101) & (g112) & (g117)) + ((shiftx4x) & (!shiftx5x) & (g91) & (!g101) & (g112) & (!g117)) + ((shiftx4x) & (!shiftx5x) & (g91) & (!g101) & (g112) & (g117)) + ((shiftx4x) & (!shiftx5x) & (g91) & (g101) & (g112) & (!g117)) + ((shiftx4x) & (!shiftx5x) & (g91) & (g101) & (g112) & (g117)) + ((shiftx4x) & (shiftx5x) & (!g91) & (g101) & (!g112) & (!g117)) + ((shiftx4x) & (shiftx5x) & (!g91) & (g101) & (!g112) & (g117)) + ((shiftx4x) & (shiftx5x) & (!g91) & (g101) & (g112) & (!g117)) + ((shiftx4x) & (shiftx5x) & (!g91) & (g101) & (g112) & (g117)) + ((shiftx4x) & (shiftx5x) & (g91) & (g101) & (!g112) & (!g117)) + ((shiftx4x) & (shiftx5x) & (g91) & (g101) & (!g112) & (g117)) + ((shiftx4x) & (shiftx5x) & (g91) & (g101) & (g112) & (!g117)) + ((shiftx4x) & (shiftx5x) & (g91) & (g101) & (g112) & (g117)));
	assign g360 = (((!shiftx4x) & (!shiftx5x) & (!g96) & (g106) & (!g122) & (!g127)) + ((!shiftx4x) & (!shiftx5x) & (!g96) & (g106) & (!g122) & (g127)) + ((!shiftx4x) & (!shiftx5x) & (!g96) & (g106) & (g122) & (!g127)) + ((!shiftx4x) & (!shiftx5x) & (!g96) & (g106) & (g122) & (g127)) + ((!shiftx4x) & (!shiftx5x) & (g96) & (g106) & (!g122) & (!g127)) + ((!shiftx4x) & (!shiftx5x) & (g96) & (g106) & (!g122) & (g127)) + ((!shiftx4x) & (!shiftx5x) & (g96) & (g106) & (g122) & (!g127)) + ((!shiftx4x) & (!shiftx5x) & (g96) & (g106) & (g122) & (g127)) + ((!shiftx4x) & (shiftx5x) & (!g96) & (!g106) & (g122) & (!g127)) + ((!shiftx4x) & (shiftx5x) & (!g96) & (!g106) & (g122) & (g127)) + ((!shiftx4x) & (shiftx5x) & (!g96) & (g106) & (g122) & (!g127)) + ((!shiftx4x) & (shiftx5x) & (!g96) & (g106) & (g122) & (g127)) + ((!shiftx4x) & (shiftx5x) & (g96) & (!g106) & (g122) & (!g127)) + ((!shiftx4x) & (shiftx5x) & (g96) & (!g106) & (g122) & (g127)) + ((!shiftx4x) & (shiftx5x) & (g96) & (g106) & (g122) & (!g127)) + ((!shiftx4x) & (shiftx5x) & (g96) & (g106) & (g122) & (g127)) + ((shiftx4x) & (!shiftx5x) & (g96) & (!g106) & (!g122) & (!g127)) + ((shiftx4x) & (!shiftx5x) & (g96) & (!g106) & (!g122) & (g127)) + ((shiftx4x) & (!shiftx5x) & (g96) & (!g106) & (g122) & (!g127)) + ((shiftx4x) & (!shiftx5x) & (g96) & (!g106) & (g122) & (g127)) + ((shiftx4x) & (!shiftx5x) & (g96) & (g106) & (!g122) & (!g127)) + ((shiftx4x) & (!shiftx5x) & (g96) & (g106) & (!g122) & (g127)) + ((shiftx4x) & (!shiftx5x) & (g96) & (g106) & (g122) & (!g127)) + ((shiftx4x) & (!shiftx5x) & (g96) & (g106) & (g122) & (g127)) + ((shiftx4x) & (shiftx5x) & (!g96) & (!g106) & (!g122) & (g127)) + ((shiftx4x) & (shiftx5x) & (!g96) & (!g106) & (g122) & (g127)) + ((shiftx4x) & (shiftx5x) & (!g96) & (g106) & (!g122) & (g127)) + ((shiftx4x) & (shiftx5x) & (!g96) & (g106) & (g122) & (g127)) + ((shiftx4x) & (shiftx5x) & (g96) & (!g106) & (!g122) & (g127)) + ((shiftx4x) & (shiftx5x) & (g96) & (!g106) & (g122) & (g127)) + ((shiftx4x) & (shiftx5x) & (g96) & (g106) & (!g122) & (g127)) + ((shiftx4x) & (shiftx5x) & (g96) & (g106) & (g122) & (g127)));
	assign resultx34x = (((!shiftx6x) & (sk[104]) & (!g359) & (g360)) + ((!shiftx6x) & (sk[104]) & (g359) & (g360)) + ((shiftx6x) & (!sk[104]) & (!g359) & (!g360)) + ((shiftx6x) & (!sk[104]) & (!g359) & (g360)) + ((shiftx6x) & (!sk[104]) & (g359) & (!g360)) + ((shiftx6x) & (!sk[104]) & (g359) & (g360)) + ((shiftx6x) & (sk[104]) & (g359) & (!g360)) + ((shiftx6x) & (sk[104]) & (g359) & (g360)));
	assign g362 = (((!shiftx4x) & (!shiftx5x) & (!g134) & (!g139) & (g160) & (!g170)) + ((!shiftx4x) & (!shiftx5x) & (!g134) & (!g139) & (g160) & (g170)) + ((!shiftx4x) & (!shiftx5x) & (!g134) & (g139) & (g160) & (!g170)) + ((!shiftx4x) & (!shiftx5x) & (!g134) & (g139) & (g160) & (g170)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (!g139) & (g160) & (!g170)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (!g139) & (g160) & (g170)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (g139) & (g160) & (!g170)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (g139) & (g160) & (g170)) + ((!shiftx4x) & (shiftx5x) & (g134) & (!g139) & (!g160) & (!g170)) + ((!shiftx4x) & (shiftx5x) & (g134) & (!g139) & (!g160) & (g170)) + ((!shiftx4x) & (shiftx5x) & (g134) & (!g139) & (g160) & (!g170)) + ((!shiftx4x) & (shiftx5x) & (g134) & (!g139) & (g160) & (g170)) + ((!shiftx4x) & (shiftx5x) & (g134) & (g139) & (!g160) & (!g170)) + ((!shiftx4x) & (shiftx5x) & (g134) & (g139) & (!g160) & (g170)) + ((!shiftx4x) & (shiftx5x) & (g134) & (g139) & (g160) & (!g170)) + ((!shiftx4x) & (shiftx5x) & (g134) & (g139) & (g160) & (g170)) + ((shiftx4x) & (!shiftx5x) & (!g134) & (!g139) & (!g160) & (g170)) + ((shiftx4x) & (!shiftx5x) & (!g134) & (!g139) & (g160) & (g170)) + ((shiftx4x) & (!shiftx5x) & (!g134) & (g139) & (!g160) & (g170)) + ((shiftx4x) & (!shiftx5x) & (!g134) & (g139) & (g160) & (g170)) + ((shiftx4x) & (!shiftx5x) & (g134) & (!g139) & (!g160) & (g170)) + ((shiftx4x) & (!shiftx5x) & (g134) & (!g139) & (g160) & (g170)) + ((shiftx4x) & (!shiftx5x) & (g134) & (g139) & (!g160) & (g170)) + ((shiftx4x) & (!shiftx5x) & (g134) & (g139) & (g160) & (g170)) + ((shiftx4x) & (shiftx5x) & (!g134) & (g139) & (!g160) & (!g170)) + ((shiftx4x) & (shiftx5x) & (!g134) & (g139) & (!g160) & (g170)) + ((shiftx4x) & (shiftx5x) & (!g134) & (g139) & (g160) & (!g170)) + ((shiftx4x) & (shiftx5x) & (!g134) & (g139) & (g160) & (g170)) + ((shiftx4x) & (shiftx5x) & (g134) & (g139) & (!g160) & (!g170)) + ((shiftx4x) & (shiftx5x) & (g134) & (g139) & (!g160) & (g170)) + ((shiftx4x) & (shiftx5x) & (g134) & (g139) & (g160) & (!g170)) + ((shiftx4x) & (shiftx5x) & (g134) & (g139) & (g160) & (g170)));
	assign g363 = (((!shiftx4x) & (!shiftx5x) & (!g144) & (g149) & (!g155) & (!g165)) + ((!shiftx4x) & (!shiftx5x) & (!g144) & (g149) & (!g155) & (g165)) + ((!shiftx4x) & (!shiftx5x) & (!g144) & (g149) & (g155) & (!g165)) + ((!shiftx4x) & (!shiftx5x) & (!g144) & (g149) & (g155) & (g165)) + ((!shiftx4x) & (!shiftx5x) & (g144) & (g149) & (!g155) & (!g165)) + ((!shiftx4x) & (!shiftx5x) & (g144) & (g149) & (!g155) & (g165)) + ((!shiftx4x) & (!shiftx5x) & (g144) & (g149) & (g155) & (!g165)) + ((!shiftx4x) & (!shiftx5x) & (g144) & (g149) & (g155) & (g165)) + ((!shiftx4x) & (shiftx5x) & (!g144) & (!g149) & (!g155) & (g165)) + ((!shiftx4x) & (shiftx5x) & (!g144) & (!g149) & (g155) & (g165)) + ((!shiftx4x) & (shiftx5x) & (!g144) & (g149) & (!g155) & (g165)) + ((!shiftx4x) & (shiftx5x) & (!g144) & (g149) & (g155) & (g165)) + ((!shiftx4x) & (shiftx5x) & (g144) & (!g149) & (!g155) & (g165)) + ((!shiftx4x) & (shiftx5x) & (g144) & (!g149) & (g155) & (g165)) + ((!shiftx4x) & (shiftx5x) & (g144) & (g149) & (!g155) & (g165)) + ((!shiftx4x) & (shiftx5x) & (g144) & (g149) & (g155) & (g165)) + ((shiftx4x) & (!shiftx5x) & (g144) & (!g149) & (!g155) & (!g165)) + ((shiftx4x) & (!shiftx5x) & (g144) & (!g149) & (!g155) & (g165)) + ((shiftx4x) & (!shiftx5x) & (g144) & (!g149) & (g155) & (!g165)) + ((shiftx4x) & (!shiftx5x) & (g144) & (!g149) & (g155) & (g165)) + ((shiftx4x) & (!shiftx5x) & (g144) & (g149) & (!g155) & (!g165)) + ((shiftx4x) & (!shiftx5x) & (g144) & (g149) & (!g155) & (g165)) + ((shiftx4x) & (!shiftx5x) & (g144) & (g149) & (g155) & (!g165)) + ((shiftx4x) & (!shiftx5x) & (g144) & (g149) & (g155) & (g165)) + ((shiftx4x) & (shiftx5x) & (!g144) & (!g149) & (g155) & (!g165)) + ((shiftx4x) & (shiftx5x) & (!g144) & (!g149) & (g155) & (g165)) + ((shiftx4x) & (shiftx5x) & (!g144) & (g149) & (g155) & (!g165)) + ((shiftx4x) & (shiftx5x) & (!g144) & (g149) & (g155) & (g165)) + ((shiftx4x) & (shiftx5x) & (g144) & (!g149) & (g155) & (!g165)) + ((shiftx4x) & (shiftx5x) & (g144) & (!g149) & (g155) & (g165)) + ((shiftx4x) & (shiftx5x) & (g144) & (g149) & (g155) & (!g165)) + ((shiftx4x) & (shiftx5x) & (g144) & (g149) & (g155) & (g165)));
	assign resultx35x = (((!shiftx6x) & (!g362) & (sk[107]) & (g363)) + ((!shiftx6x) & (g362) & (sk[107]) & (g363)) + ((shiftx6x) & (!g362) & (!sk[107]) & (!g363)) + ((shiftx6x) & (!g362) & (!sk[107]) & (g363)) + ((shiftx6x) & (g362) & (!sk[107]) & (!g363)) + ((shiftx6x) & (g362) & (!sk[107]) & (g363)) + ((shiftx6x) & (g362) & (sk[107]) & (!g363)) + ((shiftx6x) & (g362) & (sk[107]) & (g363)));
	assign g365 = (((!shiftx4x) & (!shiftx5x) & (!g173) & (!g174) & (!g178) & (g179)) + ((!shiftx4x) & (!shiftx5x) & (!g173) & (!g174) & (g178) & (g179)) + ((!shiftx4x) & (!shiftx5x) & (!g173) & (g174) & (!g178) & (g179)) + ((!shiftx4x) & (!shiftx5x) & (!g173) & (g174) & (g178) & (g179)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (!g174) & (!g178) & (g179)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (!g174) & (g178) & (g179)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (g174) & (!g178) & (g179)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (g174) & (g178) & (g179)) + ((!shiftx4x) & (shiftx5x) & (!g173) & (g174) & (!g178) & (!g179)) + ((!shiftx4x) & (shiftx5x) & (!g173) & (g174) & (!g178) & (g179)) + ((!shiftx4x) & (shiftx5x) & (!g173) & (g174) & (g178) & (!g179)) + ((!shiftx4x) & (shiftx5x) & (!g173) & (g174) & (g178) & (g179)) + ((!shiftx4x) & (shiftx5x) & (g173) & (g174) & (!g178) & (!g179)) + ((!shiftx4x) & (shiftx5x) & (g173) & (g174) & (!g178) & (g179)) + ((!shiftx4x) & (shiftx5x) & (g173) & (g174) & (g178) & (!g179)) + ((!shiftx4x) & (shiftx5x) & (g173) & (g174) & (g178) & (g179)) + ((shiftx4x) & (!shiftx5x) & (!g173) & (!g174) & (g178) & (!g179)) + ((shiftx4x) & (!shiftx5x) & (!g173) & (!g174) & (g178) & (g179)) + ((shiftx4x) & (!shiftx5x) & (!g173) & (g174) & (g178) & (!g179)) + ((shiftx4x) & (!shiftx5x) & (!g173) & (g174) & (g178) & (g179)) + ((shiftx4x) & (!shiftx5x) & (g173) & (!g174) & (g178) & (!g179)) + ((shiftx4x) & (!shiftx5x) & (g173) & (!g174) & (g178) & (g179)) + ((shiftx4x) & (!shiftx5x) & (g173) & (g174) & (g178) & (!g179)) + ((shiftx4x) & (!shiftx5x) & (g173) & (g174) & (g178) & (g179)) + ((shiftx4x) & (shiftx5x) & (g173) & (!g174) & (!g178) & (!g179)) + ((shiftx4x) & (shiftx5x) & (g173) & (!g174) & (!g178) & (g179)) + ((shiftx4x) & (shiftx5x) & (g173) & (!g174) & (g178) & (!g179)) + ((shiftx4x) & (shiftx5x) & (g173) & (!g174) & (g178) & (g179)) + ((shiftx4x) & (shiftx5x) & (g173) & (g174) & (!g178) & (!g179)) + ((shiftx4x) & (shiftx5x) & (g173) & (g174) & (!g178) & (g179)) + ((shiftx4x) & (shiftx5x) & (g173) & (g174) & (g178) & (!g179)) + ((shiftx4x) & (shiftx5x) & (g173) & (g174) & (g178) & (g179)));
	assign g366 = (((!shiftx4x) & (!shiftx5x) & (g175) & (!g176) & (!g180) & (!g181)) + ((!shiftx4x) & (!shiftx5x) & (g175) & (!g176) & (!g180) & (g181)) + ((!shiftx4x) & (!shiftx5x) & (g175) & (!g176) & (g180) & (!g181)) + ((!shiftx4x) & (!shiftx5x) & (g175) & (!g176) & (g180) & (g181)) + ((!shiftx4x) & (!shiftx5x) & (g175) & (g176) & (!g180) & (!g181)) + ((!shiftx4x) & (!shiftx5x) & (g175) & (g176) & (!g180) & (g181)) + ((!shiftx4x) & (!shiftx5x) & (g175) & (g176) & (g180) & (!g181)) + ((!shiftx4x) & (!shiftx5x) & (g175) & (g176) & (g180) & (g181)) + ((!shiftx4x) & (shiftx5x) & (!g175) & (!g176) & (g180) & (!g181)) + ((!shiftx4x) & (shiftx5x) & (!g175) & (!g176) & (g180) & (g181)) + ((!shiftx4x) & (shiftx5x) & (!g175) & (g176) & (g180) & (!g181)) + ((!shiftx4x) & (shiftx5x) & (!g175) & (g176) & (g180) & (g181)) + ((!shiftx4x) & (shiftx5x) & (g175) & (!g176) & (g180) & (!g181)) + ((!shiftx4x) & (shiftx5x) & (g175) & (!g176) & (g180) & (g181)) + ((!shiftx4x) & (shiftx5x) & (g175) & (g176) & (g180) & (!g181)) + ((!shiftx4x) & (shiftx5x) & (g175) & (g176) & (g180) & (g181)) + ((shiftx4x) & (!shiftx5x) & (!g175) & (g176) & (!g180) & (!g181)) + ((shiftx4x) & (!shiftx5x) & (!g175) & (g176) & (!g180) & (g181)) + ((shiftx4x) & (!shiftx5x) & (!g175) & (g176) & (g180) & (!g181)) + ((shiftx4x) & (!shiftx5x) & (!g175) & (g176) & (g180) & (g181)) + ((shiftx4x) & (!shiftx5x) & (g175) & (g176) & (!g180) & (!g181)) + ((shiftx4x) & (!shiftx5x) & (g175) & (g176) & (!g180) & (g181)) + ((shiftx4x) & (!shiftx5x) & (g175) & (g176) & (g180) & (!g181)) + ((shiftx4x) & (!shiftx5x) & (g175) & (g176) & (g180) & (g181)) + ((shiftx4x) & (shiftx5x) & (!g175) & (!g176) & (!g180) & (g181)) + ((shiftx4x) & (shiftx5x) & (!g175) & (!g176) & (g180) & (g181)) + ((shiftx4x) & (shiftx5x) & (!g175) & (g176) & (!g180) & (g181)) + ((shiftx4x) & (shiftx5x) & (!g175) & (g176) & (g180) & (g181)) + ((shiftx4x) & (shiftx5x) & (g175) & (!g176) & (!g180) & (g181)) + ((shiftx4x) & (shiftx5x) & (g175) & (!g176) & (g180) & (g181)) + ((shiftx4x) & (shiftx5x) & (g175) & (g176) & (!g180) & (g181)) + ((shiftx4x) & (shiftx5x) & (g175) & (g176) & (g180) & (g181)));
	assign resultx36x = (((!sk[110]) & (shiftx6x) & (!g365) & (!g366)) + ((!sk[110]) & (shiftx6x) & (!g365) & (g366)) + ((!sk[110]) & (shiftx6x) & (g365) & (!g366)) + ((!sk[110]) & (shiftx6x) & (g365) & (g366)) + ((sk[110]) & (!shiftx6x) & (!g365) & (g366)) + ((sk[110]) & (!shiftx6x) & (g365) & (g366)) + ((sk[110]) & (shiftx6x) & (g365) & (!g366)) + ((sk[110]) & (shiftx6x) & (g365) & (g366)));
	assign g368 = (((!shiftx4x) & (!shiftx5x) & (!g184) & (!g185) & (!g189) & (g190)) + ((!shiftx4x) & (!shiftx5x) & (!g184) & (!g185) & (g189) & (g190)) + ((!shiftx4x) & (!shiftx5x) & (!g184) & (g185) & (!g189) & (g190)) + ((!shiftx4x) & (!shiftx5x) & (!g184) & (g185) & (g189) & (g190)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (!g185) & (!g189) & (g190)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (!g185) & (g189) & (g190)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (g185) & (!g189) & (g190)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (g185) & (g189) & (g190)) + ((!shiftx4x) & (shiftx5x) & (!g184) & (g185) & (!g189) & (!g190)) + ((!shiftx4x) & (shiftx5x) & (!g184) & (g185) & (!g189) & (g190)) + ((!shiftx4x) & (shiftx5x) & (!g184) & (g185) & (g189) & (!g190)) + ((!shiftx4x) & (shiftx5x) & (!g184) & (g185) & (g189) & (g190)) + ((!shiftx4x) & (shiftx5x) & (g184) & (g185) & (!g189) & (!g190)) + ((!shiftx4x) & (shiftx5x) & (g184) & (g185) & (!g189) & (g190)) + ((!shiftx4x) & (shiftx5x) & (g184) & (g185) & (g189) & (!g190)) + ((!shiftx4x) & (shiftx5x) & (g184) & (g185) & (g189) & (g190)) + ((shiftx4x) & (!shiftx5x) & (!g184) & (!g185) & (g189) & (!g190)) + ((shiftx4x) & (!shiftx5x) & (!g184) & (!g185) & (g189) & (g190)) + ((shiftx4x) & (!shiftx5x) & (!g184) & (g185) & (g189) & (!g190)) + ((shiftx4x) & (!shiftx5x) & (!g184) & (g185) & (g189) & (g190)) + ((shiftx4x) & (!shiftx5x) & (g184) & (!g185) & (g189) & (!g190)) + ((shiftx4x) & (!shiftx5x) & (g184) & (!g185) & (g189) & (g190)) + ((shiftx4x) & (!shiftx5x) & (g184) & (g185) & (g189) & (!g190)) + ((shiftx4x) & (!shiftx5x) & (g184) & (g185) & (g189) & (g190)) + ((shiftx4x) & (shiftx5x) & (g184) & (!g185) & (!g189) & (!g190)) + ((shiftx4x) & (shiftx5x) & (g184) & (!g185) & (!g189) & (g190)) + ((shiftx4x) & (shiftx5x) & (g184) & (!g185) & (g189) & (!g190)) + ((shiftx4x) & (shiftx5x) & (g184) & (!g185) & (g189) & (g190)) + ((shiftx4x) & (shiftx5x) & (g184) & (g185) & (!g189) & (!g190)) + ((shiftx4x) & (shiftx5x) & (g184) & (g185) & (!g189) & (g190)) + ((shiftx4x) & (shiftx5x) & (g184) & (g185) & (g189) & (!g190)) + ((shiftx4x) & (shiftx5x) & (g184) & (g185) & (g189) & (g190)));
	assign g369 = (((!shiftx4x) & (!shiftx5x) & (g186) & (!g187) & (!g191) & (!g192)) + ((!shiftx4x) & (!shiftx5x) & (g186) & (!g187) & (!g191) & (g192)) + ((!shiftx4x) & (!shiftx5x) & (g186) & (!g187) & (g191) & (!g192)) + ((!shiftx4x) & (!shiftx5x) & (g186) & (!g187) & (g191) & (g192)) + ((!shiftx4x) & (!shiftx5x) & (g186) & (g187) & (!g191) & (!g192)) + ((!shiftx4x) & (!shiftx5x) & (g186) & (g187) & (!g191) & (g192)) + ((!shiftx4x) & (!shiftx5x) & (g186) & (g187) & (g191) & (!g192)) + ((!shiftx4x) & (!shiftx5x) & (g186) & (g187) & (g191) & (g192)) + ((!shiftx4x) & (shiftx5x) & (!g186) & (!g187) & (g191) & (!g192)) + ((!shiftx4x) & (shiftx5x) & (!g186) & (!g187) & (g191) & (g192)) + ((!shiftx4x) & (shiftx5x) & (!g186) & (g187) & (g191) & (!g192)) + ((!shiftx4x) & (shiftx5x) & (!g186) & (g187) & (g191) & (g192)) + ((!shiftx4x) & (shiftx5x) & (g186) & (!g187) & (g191) & (!g192)) + ((!shiftx4x) & (shiftx5x) & (g186) & (!g187) & (g191) & (g192)) + ((!shiftx4x) & (shiftx5x) & (g186) & (g187) & (g191) & (!g192)) + ((!shiftx4x) & (shiftx5x) & (g186) & (g187) & (g191) & (g192)) + ((shiftx4x) & (!shiftx5x) & (!g186) & (g187) & (!g191) & (!g192)) + ((shiftx4x) & (!shiftx5x) & (!g186) & (g187) & (!g191) & (g192)) + ((shiftx4x) & (!shiftx5x) & (!g186) & (g187) & (g191) & (!g192)) + ((shiftx4x) & (!shiftx5x) & (!g186) & (g187) & (g191) & (g192)) + ((shiftx4x) & (!shiftx5x) & (g186) & (g187) & (!g191) & (!g192)) + ((shiftx4x) & (!shiftx5x) & (g186) & (g187) & (!g191) & (g192)) + ((shiftx4x) & (!shiftx5x) & (g186) & (g187) & (g191) & (!g192)) + ((shiftx4x) & (!shiftx5x) & (g186) & (g187) & (g191) & (g192)) + ((shiftx4x) & (shiftx5x) & (!g186) & (!g187) & (!g191) & (g192)) + ((shiftx4x) & (shiftx5x) & (!g186) & (!g187) & (g191) & (g192)) + ((shiftx4x) & (shiftx5x) & (!g186) & (g187) & (!g191) & (g192)) + ((shiftx4x) & (shiftx5x) & (!g186) & (g187) & (g191) & (g192)) + ((shiftx4x) & (shiftx5x) & (g186) & (!g187) & (!g191) & (g192)) + ((shiftx4x) & (shiftx5x) & (g186) & (!g187) & (g191) & (g192)) + ((shiftx4x) & (shiftx5x) & (g186) & (g187) & (!g191) & (g192)) + ((shiftx4x) & (shiftx5x) & (g186) & (g187) & (g191) & (g192)));
	assign resultx37x = (((!sk[113]) & (shiftx6x) & (!g368) & (!g369)) + ((!sk[113]) & (shiftx6x) & (!g368) & (g369)) + ((!sk[113]) & (shiftx6x) & (g368) & (!g369)) + ((!sk[113]) & (shiftx6x) & (g368) & (g369)) + ((sk[113]) & (!shiftx6x) & (!g368) & (g369)) + ((sk[113]) & (!shiftx6x) & (g368) & (g369)) + ((sk[113]) & (shiftx6x) & (g368) & (!g369)) + ((sk[113]) & (shiftx6x) & (g368) & (g369)));
	assign g371 = (((!shiftx4x) & (!shiftx5x) & (!g195) & (!g196) & (!g200) & (g201)) + ((!shiftx4x) & (!shiftx5x) & (!g195) & (!g196) & (g200) & (g201)) + ((!shiftx4x) & (!shiftx5x) & (!g195) & (g196) & (!g200) & (g201)) + ((!shiftx4x) & (!shiftx5x) & (!g195) & (g196) & (g200) & (g201)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (!g196) & (!g200) & (g201)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (!g196) & (g200) & (g201)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (g196) & (!g200) & (g201)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (g196) & (g200) & (g201)) + ((!shiftx4x) & (shiftx5x) & (!g195) & (g196) & (!g200) & (!g201)) + ((!shiftx4x) & (shiftx5x) & (!g195) & (g196) & (!g200) & (g201)) + ((!shiftx4x) & (shiftx5x) & (!g195) & (g196) & (g200) & (!g201)) + ((!shiftx4x) & (shiftx5x) & (!g195) & (g196) & (g200) & (g201)) + ((!shiftx4x) & (shiftx5x) & (g195) & (g196) & (!g200) & (!g201)) + ((!shiftx4x) & (shiftx5x) & (g195) & (g196) & (!g200) & (g201)) + ((!shiftx4x) & (shiftx5x) & (g195) & (g196) & (g200) & (!g201)) + ((!shiftx4x) & (shiftx5x) & (g195) & (g196) & (g200) & (g201)) + ((shiftx4x) & (!shiftx5x) & (!g195) & (!g196) & (g200) & (!g201)) + ((shiftx4x) & (!shiftx5x) & (!g195) & (!g196) & (g200) & (g201)) + ((shiftx4x) & (!shiftx5x) & (!g195) & (g196) & (g200) & (!g201)) + ((shiftx4x) & (!shiftx5x) & (!g195) & (g196) & (g200) & (g201)) + ((shiftx4x) & (!shiftx5x) & (g195) & (!g196) & (g200) & (!g201)) + ((shiftx4x) & (!shiftx5x) & (g195) & (!g196) & (g200) & (g201)) + ((shiftx4x) & (!shiftx5x) & (g195) & (g196) & (g200) & (!g201)) + ((shiftx4x) & (!shiftx5x) & (g195) & (g196) & (g200) & (g201)) + ((shiftx4x) & (shiftx5x) & (g195) & (!g196) & (!g200) & (!g201)) + ((shiftx4x) & (shiftx5x) & (g195) & (!g196) & (!g200) & (g201)) + ((shiftx4x) & (shiftx5x) & (g195) & (!g196) & (g200) & (!g201)) + ((shiftx4x) & (shiftx5x) & (g195) & (!g196) & (g200) & (g201)) + ((shiftx4x) & (shiftx5x) & (g195) & (g196) & (!g200) & (!g201)) + ((shiftx4x) & (shiftx5x) & (g195) & (g196) & (!g200) & (g201)) + ((shiftx4x) & (shiftx5x) & (g195) & (g196) & (g200) & (!g201)) + ((shiftx4x) & (shiftx5x) & (g195) & (g196) & (g200) & (g201)));
	assign g372 = (((!shiftx4x) & (!shiftx5x) & (g197) & (!g198) & (!g202) & (!g203)) + ((!shiftx4x) & (!shiftx5x) & (g197) & (!g198) & (!g202) & (g203)) + ((!shiftx4x) & (!shiftx5x) & (g197) & (!g198) & (g202) & (!g203)) + ((!shiftx4x) & (!shiftx5x) & (g197) & (!g198) & (g202) & (g203)) + ((!shiftx4x) & (!shiftx5x) & (g197) & (g198) & (!g202) & (!g203)) + ((!shiftx4x) & (!shiftx5x) & (g197) & (g198) & (!g202) & (g203)) + ((!shiftx4x) & (!shiftx5x) & (g197) & (g198) & (g202) & (!g203)) + ((!shiftx4x) & (!shiftx5x) & (g197) & (g198) & (g202) & (g203)) + ((!shiftx4x) & (shiftx5x) & (!g197) & (!g198) & (g202) & (!g203)) + ((!shiftx4x) & (shiftx5x) & (!g197) & (!g198) & (g202) & (g203)) + ((!shiftx4x) & (shiftx5x) & (!g197) & (g198) & (g202) & (!g203)) + ((!shiftx4x) & (shiftx5x) & (!g197) & (g198) & (g202) & (g203)) + ((!shiftx4x) & (shiftx5x) & (g197) & (!g198) & (g202) & (!g203)) + ((!shiftx4x) & (shiftx5x) & (g197) & (!g198) & (g202) & (g203)) + ((!shiftx4x) & (shiftx5x) & (g197) & (g198) & (g202) & (!g203)) + ((!shiftx4x) & (shiftx5x) & (g197) & (g198) & (g202) & (g203)) + ((shiftx4x) & (!shiftx5x) & (!g197) & (g198) & (!g202) & (!g203)) + ((shiftx4x) & (!shiftx5x) & (!g197) & (g198) & (!g202) & (g203)) + ((shiftx4x) & (!shiftx5x) & (!g197) & (g198) & (g202) & (!g203)) + ((shiftx4x) & (!shiftx5x) & (!g197) & (g198) & (g202) & (g203)) + ((shiftx4x) & (!shiftx5x) & (g197) & (g198) & (!g202) & (!g203)) + ((shiftx4x) & (!shiftx5x) & (g197) & (g198) & (!g202) & (g203)) + ((shiftx4x) & (!shiftx5x) & (g197) & (g198) & (g202) & (!g203)) + ((shiftx4x) & (!shiftx5x) & (g197) & (g198) & (g202) & (g203)) + ((shiftx4x) & (shiftx5x) & (!g197) & (!g198) & (!g202) & (g203)) + ((shiftx4x) & (shiftx5x) & (!g197) & (!g198) & (g202) & (g203)) + ((shiftx4x) & (shiftx5x) & (!g197) & (g198) & (!g202) & (g203)) + ((shiftx4x) & (shiftx5x) & (!g197) & (g198) & (g202) & (g203)) + ((shiftx4x) & (shiftx5x) & (g197) & (!g198) & (!g202) & (g203)) + ((shiftx4x) & (shiftx5x) & (g197) & (!g198) & (g202) & (g203)) + ((shiftx4x) & (shiftx5x) & (g197) & (g198) & (!g202) & (g203)) + ((shiftx4x) & (shiftx5x) & (g197) & (g198) & (g202) & (g203)));
	assign resultx38x = (((!shiftx6x) & (!g371) & (sk[116]) & (g372)) + ((!shiftx6x) & (g371) & (sk[116]) & (g372)) + ((shiftx6x) & (!g371) & (!sk[116]) & (!g372)) + ((shiftx6x) & (!g371) & (!sk[116]) & (g372)) + ((shiftx6x) & (g371) & (!sk[116]) & (!g372)) + ((shiftx6x) & (g371) & (!sk[116]) & (g372)) + ((shiftx6x) & (g371) & (sk[116]) & (!g372)) + ((shiftx6x) & (g371) & (sk[116]) & (g372)));
	assign g374 = (((!shiftx4x) & (!shiftx5x) & (!g206) & (!g207) & (!g211) & (g212)) + ((!shiftx4x) & (!shiftx5x) & (!g206) & (!g207) & (g211) & (g212)) + ((!shiftx4x) & (!shiftx5x) & (!g206) & (g207) & (!g211) & (g212)) + ((!shiftx4x) & (!shiftx5x) & (!g206) & (g207) & (g211) & (g212)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (!g207) & (!g211) & (g212)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (!g207) & (g211) & (g212)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (g207) & (!g211) & (g212)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (g207) & (g211) & (g212)) + ((!shiftx4x) & (shiftx5x) & (!g206) & (g207) & (!g211) & (!g212)) + ((!shiftx4x) & (shiftx5x) & (!g206) & (g207) & (!g211) & (g212)) + ((!shiftx4x) & (shiftx5x) & (!g206) & (g207) & (g211) & (!g212)) + ((!shiftx4x) & (shiftx5x) & (!g206) & (g207) & (g211) & (g212)) + ((!shiftx4x) & (shiftx5x) & (g206) & (g207) & (!g211) & (!g212)) + ((!shiftx4x) & (shiftx5x) & (g206) & (g207) & (!g211) & (g212)) + ((!shiftx4x) & (shiftx5x) & (g206) & (g207) & (g211) & (!g212)) + ((!shiftx4x) & (shiftx5x) & (g206) & (g207) & (g211) & (g212)) + ((shiftx4x) & (!shiftx5x) & (!g206) & (!g207) & (g211) & (!g212)) + ((shiftx4x) & (!shiftx5x) & (!g206) & (!g207) & (g211) & (g212)) + ((shiftx4x) & (!shiftx5x) & (!g206) & (g207) & (g211) & (!g212)) + ((shiftx4x) & (!shiftx5x) & (!g206) & (g207) & (g211) & (g212)) + ((shiftx4x) & (!shiftx5x) & (g206) & (!g207) & (g211) & (!g212)) + ((shiftx4x) & (!shiftx5x) & (g206) & (!g207) & (g211) & (g212)) + ((shiftx4x) & (!shiftx5x) & (g206) & (g207) & (g211) & (!g212)) + ((shiftx4x) & (!shiftx5x) & (g206) & (g207) & (g211) & (g212)) + ((shiftx4x) & (shiftx5x) & (g206) & (!g207) & (!g211) & (!g212)) + ((shiftx4x) & (shiftx5x) & (g206) & (!g207) & (!g211) & (g212)) + ((shiftx4x) & (shiftx5x) & (g206) & (!g207) & (g211) & (!g212)) + ((shiftx4x) & (shiftx5x) & (g206) & (!g207) & (g211) & (g212)) + ((shiftx4x) & (shiftx5x) & (g206) & (g207) & (!g211) & (!g212)) + ((shiftx4x) & (shiftx5x) & (g206) & (g207) & (!g211) & (g212)) + ((shiftx4x) & (shiftx5x) & (g206) & (g207) & (g211) & (!g212)) + ((shiftx4x) & (shiftx5x) & (g206) & (g207) & (g211) & (g212)));
	assign g375 = (((!shiftx4x) & (!shiftx5x) & (g208) & (!g209) & (!g213) & (!g214)) + ((!shiftx4x) & (!shiftx5x) & (g208) & (!g209) & (!g213) & (g214)) + ((!shiftx4x) & (!shiftx5x) & (g208) & (!g209) & (g213) & (!g214)) + ((!shiftx4x) & (!shiftx5x) & (g208) & (!g209) & (g213) & (g214)) + ((!shiftx4x) & (!shiftx5x) & (g208) & (g209) & (!g213) & (!g214)) + ((!shiftx4x) & (!shiftx5x) & (g208) & (g209) & (!g213) & (g214)) + ((!shiftx4x) & (!shiftx5x) & (g208) & (g209) & (g213) & (!g214)) + ((!shiftx4x) & (!shiftx5x) & (g208) & (g209) & (g213) & (g214)) + ((!shiftx4x) & (shiftx5x) & (!g208) & (!g209) & (g213) & (!g214)) + ((!shiftx4x) & (shiftx5x) & (!g208) & (!g209) & (g213) & (g214)) + ((!shiftx4x) & (shiftx5x) & (!g208) & (g209) & (g213) & (!g214)) + ((!shiftx4x) & (shiftx5x) & (!g208) & (g209) & (g213) & (g214)) + ((!shiftx4x) & (shiftx5x) & (g208) & (!g209) & (g213) & (!g214)) + ((!shiftx4x) & (shiftx5x) & (g208) & (!g209) & (g213) & (g214)) + ((!shiftx4x) & (shiftx5x) & (g208) & (g209) & (g213) & (!g214)) + ((!shiftx4x) & (shiftx5x) & (g208) & (g209) & (g213) & (g214)) + ((shiftx4x) & (!shiftx5x) & (!g208) & (g209) & (!g213) & (!g214)) + ((shiftx4x) & (!shiftx5x) & (!g208) & (g209) & (!g213) & (g214)) + ((shiftx4x) & (!shiftx5x) & (!g208) & (g209) & (g213) & (!g214)) + ((shiftx4x) & (!shiftx5x) & (!g208) & (g209) & (g213) & (g214)) + ((shiftx4x) & (!shiftx5x) & (g208) & (g209) & (!g213) & (!g214)) + ((shiftx4x) & (!shiftx5x) & (g208) & (g209) & (!g213) & (g214)) + ((shiftx4x) & (!shiftx5x) & (g208) & (g209) & (g213) & (!g214)) + ((shiftx4x) & (!shiftx5x) & (g208) & (g209) & (g213) & (g214)) + ((shiftx4x) & (shiftx5x) & (!g208) & (!g209) & (!g213) & (g214)) + ((shiftx4x) & (shiftx5x) & (!g208) & (!g209) & (g213) & (g214)) + ((shiftx4x) & (shiftx5x) & (!g208) & (g209) & (!g213) & (g214)) + ((shiftx4x) & (shiftx5x) & (!g208) & (g209) & (g213) & (g214)) + ((shiftx4x) & (shiftx5x) & (g208) & (!g209) & (!g213) & (g214)) + ((shiftx4x) & (shiftx5x) & (g208) & (!g209) & (g213) & (g214)) + ((shiftx4x) & (shiftx5x) & (g208) & (g209) & (!g213) & (g214)) + ((shiftx4x) & (shiftx5x) & (g208) & (g209) & (g213) & (g214)));
	assign resultx39x = (((!sk[119]) & (shiftx6x) & (!g374) & (!g375)) + ((!sk[119]) & (shiftx6x) & (!g374) & (g375)) + ((!sk[119]) & (shiftx6x) & (g374) & (!g375)) + ((!sk[119]) & (shiftx6x) & (g374) & (g375)) + ((sk[119]) & (!shiftx6x) & (!g374) & (g375)) + ((sk[119]) & (!shiftx6x) & (g374) & (g375)) + ((sk[119]) & (shiftx6x) & (g374) & (!g375)) + ((sk[119]) & (shiftx6x) & (g374) & (g375)));
	assign g377 = (((!shiftx4x) & (!shiftx5x) & (!g217) & (!g218) & (!g222) & (g223)) + ((!shiftx4x) & (!shiftx5x) & (!g217) & (!g218) & (g222) & (g223)) + ((!shiftx4x) & (!shiftx5x) & (!g217) & (g218) & (!g222) & (g223)) + ((!shiftx4x) & (!shiftx5x) & (!g217) & (g218) & (g222) & (g223)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (!g218) & (!g222) & (g223)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (!g218) & (g222) & (g223)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (g218) & (!g222) & (g223)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (g218) & (g222) & (g223)) + ((!shiftx4x) & (shiftx5x) & (!g217) & (g218) & (!g222) & (!g223)) + ((!shiftx4x) & (shiftx5x) & (!g217) & (g218) & (!g222) & (g223)) + ((!shiftx4x) & (shiftx5x) & (!g217) & (g218) & (g222) & (!g223)) + ((!shiftx4x) & (shiftx5x) & (!g217) & (g218) & (g222) & (g223)) + ((!shiftx4x) & (shiftx5x) & (g217) & (g218) & (!g222) & (!g223)) + ((!shiftx4x) & (shiftx5x) & (g217) & (g218) & (!g222) & (g223)) + ((!shiftx4x) & (shiftx5x) & (g217) & (g218) & (g222) & (!g223)) + ((!shiftx4x) & (shiftx5x) & (g217) & (g218) & (g222) & (g223)) + ((shiftx4x) & (!shiftx5x) & (!g217) & (!g218) & (g222) & (!g223)) + ((shiftx4x) & (!shiftx5x) & (!g217) & (!g218) & (g222) & (g223)) + ((shiftx4x) & (!shiftx5x) & (!g217) & (g218) & (g222) & (!g223)) + ((shiftx4x) & (!shiftx5x) & (!g217) & (g218) & (g222) & (g223)) + ((shiftx4x) & (!shiftx5x) & (g217) & (!g218) & (g222) & (!g223)) + ((shiftx4x) & (!shiftx5x) & (g217) & (!g218) & (g222) & (g223)) + ((shiftx4x) & (!shiftx5x) & (g217) & (g218) & (g222) & (!g223)) + ((shiftx4x) & (!shiftx5x) & (g217) & (g218) & (g222) & (g223)) + ((shiftx4x) & (shiftx5x) & (g217) & (!g218) & (!g222) & (!g223)) + ((shiftx4x) & (shiftx5x) & (g217) & (!g218) & (!g222) & (g223)) + ((shiftx4x) & (shiftx5x) & (g217) & (!g218) & (g222) & (!g223)) + ((shiftx4x) & (shiftx5x) & (g217) & (!g218) & (g222) & (g223)) + ((shiftx4x) & (shiftx5x) & (g217) & (g218) & (!g222) & (!g223)) + ((shiftx4x) & (shiftx5x) & (g217) & (g218) & (!g222) & (g223)) + ((shiftx4x) & (shiftx5x) & (g217) & (g218) & (g222) & (!g223)) + ((shiftx4x) & (shiftx5x) & (g217) & (g218) & (g222) & (g223)));
	assign g378 = (((!shiftx4x) & (!shiftx5x) & (g219) & (!g220) & (!g224) & (!g225)) + ((!shiftx4x) & (!shiftx5x) & (g219) & (!g220) & (!g224) & (g225)) + ((!shiftx4x) & (!shiftx5x) & (g219) & (!g220) & (g224) & (!g225)) + ((!shiftx4x) & (!shiftx5x) & (g219) & (!g220) & (g224) & (g225)) + ((!shiftx4x) & (!shiftx5x) & (g219) & (g220) & (!g224) & (!g225)) + ((!shiftx4x) & (!shiftx5x) & (g219) & (g220) & (!g224) & (g225)) + ((!shiftx4x) & (!shiftx5x) & (g219) & (g220) & (g224) & (!g225)) + ((!shiftx4x) & (!shiftx5x) & (g219) & (g220) & (g224) & (g225)) + ((!shiftx4x) & (shiftx5x) & (!g219) & (!g220) & (g224) & (!g225)) + ((!shiftx4x) & (shiftx5x) & (!g219) & (!g220) & (g224) & (g225)) + ((!shiftx4x) & (shiftx5x) & (!g219) & (g220) & (g224) & (!g225)) + ((!shiftx4x) & (shiftx5x) & (!g219) & (g220) & (g224) & (g225)) + ((!shiftx4x) & (shiftx5x) & (g219) & (!g220) & (g224) & (!g225)) + ((!shiftx4x) & (shiftx5x) & (g219) & (!g220) & (g224) & (g225)) + ((!shiftx4x) & (shiftx5x) & (g219) & (g220) & (g224) & (!g225)) + ((!shiftx4x) & (shiftx5x) & (g219) & (g220) & (g224) & (g225)) + ((shiftx4x) & (!shiftx5x) & (!g219) & (g220) & (!g224) & (!g225)) + ((shiftx4x) & (!shiftx5x) & (!g219) & (g220) & (!g224) & (g225)) + ((shiftx4x) & (!shiftx5x) & (!g219) & (g220) & (g224) & (!g225)) + ((shiftx4x) & (!shiftx5x) & (!g219) & (g220) & (g224) & (g225)) + ((shiftx4x) & (!shiftx5x) & (g219) & (g220) & (!g224) & (!g225)) + ((shiftx4x) & (!shiftx5x) & (g219) & (g220) & (!g224) & (g225)) + ((shiftx4x) & (!shiftx5x) & (g219) & (g220) & (g224) & (!g225)) + ((shiftx4x) & (!shiftx5x) & (g219) & (g220) & (g224) & (g225)) + ((shiftx4x) & (shiftx5x) & (!g219) & (!g220) & (!g224) & (g225)) + ((shiftx4x) & (shiftx5x) & (!g219) & (!g220) & (g224) & (g225)) + ((shiftx4x) & (shiftx5x) & (!g219) & (g220) & (!g224) & (g225)) + ((shiftx4x) & (shiftx5x) & (!g219) & (g220) & (g224) & (g225)) + ((shiftx4x) & (shiftx5x) & (g219) & (!g220) & (!g224) & (g225)) + ((shiftx4x) & (shiftx5x) & (g219) & (!g220) & (g224) & (g225)) + ((shiftx4x) & (shiftx5x) & (g219) & (g220) & (!g224) & (g225)) + ((shiftx4x) & (shiftx5x) & (g219) & (g220) & (g224) & (g225)));
	assign resultx40x = (((!sk[122]) & (shiftx6x) & (!g377) & (!g378)) + ((!sk[122]) & (shiftx6x) & (!g377) & (g378)) + ((!sk[122]) & (shiftx6x) & (g377) & (!g378)) + ((!sk[122]) & (shiftx6x) & (g377) & (g378)) + ((sk[122]) & (!shiftx6x) & (!g377) & (g378)) + ((sk[122]) & (!shiftx6x) & (g377) & (g378)) + ((sk[122]) & (shiftx6x) & (g377) & (!g378)) + ((sk[122]) & (shiftx6x) & (g377) & (g378)));
	assign g380 = (((!shiftx4x) & (!shiftx5x) & (!g228) & (!g229) & (!g233) & (g234)) + ((!shiftx4x) & (!shiftx5x) & (!g228) & (!g229) & (g233) & (g234)) + ((!shiftx4x) & (!shiftx5x) & (!g228) & (g229) & (!g233) & (g234)) + ((!shiftx4x) & (!shiftx5x) & (!g228) & (g229) & (g233) & (g234)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (!g229) & (!g233) & (g234)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (!g229) & (g233) & (g234)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (g229) & (!g233) & (g234)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (g229) & (g233) & (g234)) + ((!shiftx4x) & (shiftx5x) & (!g228) & (g229) & (!g233) & (!g234)) + ((!shiftx4x) & (shiftx5x) & (!g228) & (g229) & (!g233) & (g234)) + ((!shiftx4x) & (shiftx5x) & (!g228) & (g229) & (g233) & (!g234)) + ((!shiftx4x) & (shiftx5x) & (!g228) & (g229) & (g233) & (g234)) + ((!shiftx4x) & (shiftx5x) & (g228) & (g229) & (!g233) & (!g234)) + ((!shiftx4x) & (shiftx5x) & (g228) & (g229) & (!g233) & (g234)) + ((!shiftx4x) & (shiftx5x) & (g228) & (g229) & (g233) & (!g234)) + ((!shiftx4x) & (shiftx5x) & (g228) & (g229) & (g233) & (g234)) + ((shiftx4x) & (!shiftx5x) & (!g228) & (!g229) & (g233) & (!g234)) + ((shiftx4x) & (!shiftx5x) & (!g228) & (!g229) & (g233) & (g234)) + ((shiftx4x) & (!shiftx5x) & (!g228) & (g229) & (g233) & (!g234)) + ((shiftx4x) & (!shiftx5x) & (!g228) & (g229) & (g233) & (g234)) + ((shiftx4x) & (!shiftx5x) & (g228) & (!g229) & (g233) & (!g234)) + ((shiftx4x) & (!shiftx5x) & (g228) & (!g229) & (g233) & (g234)) + ((shiftx4x) & (!shiftx5x) & (g228) & (g229) & (g233) & (!g234)) + ((shiftx4x) & (!shiftx5x) & (g228) & (g229) & (g233) & (g234)) + ((shiftx4x) & (shiftx5x) & (g228) & (!g229) & (!g233) & (!g234)) + ((shiftx4x) & (shiftx5x) & (g228) & (!g229) & (!g233) & (g234)) + ((shiftx4x) & (shiftx5x) & (g228) & (!g229) & (g233) & (!g234)) + ((shiftx4x) & (shiftx5x) & (g228) & (!g229) & (g233) & (g234)) + ((shiftx4x) & (shiftx5x) & (g228) & (g229) & (!g233) & (!g234)) + ((shiftx4x) & (shiftx5x) & (g228) & (g229) & (!g233) & (g234)) + ((shiftx4x) & (shiftx5x) & (g228) & (g229) & (g233) & (!g234)) + ((shiftx4x) & (shiftx5x) & (g228) & (g229) & (g233) & (g234)));
	assign g381 = (((!shiftx4x) & (!shiftx5x) & (g230) & (!g231) & (!g235) & (!g236)) + ((!shiftx4x) & (!shiftx5x) & (g230) & (!g231) & (!g235) & (g236)) + ((!shiftx4x) & (!shiftx5x) & (g230) & (!g231) & (g235) & (!g236)) + ((!shiftx4x) & (!shiftx5x) & (g230) & (!g231) & (g235) & (g236)) + ((!shiftx4x) & (!shiftx5x) & (g230) & (g231) & (!g235) & (!g236)) + ((!shiftx4x) & (!shiftx5x) & (g230) & (g231) & (!g235) & (g236)) + ((!shiftx4x) & (!shiftx5x) & (g230) & (g231) & (g235) & (!g236)) + ((!shiftx4x) & (!shiftx5x) & (g230) & (g231) & (g235) & (g236)) + ((!shiftx4x) & (shiftx5x) & (!g230) & (!g231) & (g235) & (!g236)) + ((!shiftx4x) & (shiftx5x) & (!g230) & (!g231) & (g235) & (g236)) + ((!shiftx4x) & (shiftx5x) & (!g230) & (g231) & (g235) & (!g236)) + ((!shiftx4x) & (shiftx5x) & (!g230) & (g231) & (g235) & (g236)) + ((!shiftx4x) & (shiftx5x) & (g230) & (!g231) & (g235) & (!g236)) + ((!shiftx4x) & (shiftx5x) & (g230) & (!g231) & (g235) & (g236)) + ((!shiftx4x) & (shiftx5x) & (g230) & (g231) & (g235) & (!g236)) + ((!shiftx4x) & (shiftx5x) & (g230) & (g231) & (g235) & (g236)) + ((shiftx4x) & (!shiftx5x) & (!g230) & (g231) & (!g235) & (!g236)) + ((shiftx4x) & (!shiftx5x) & (!g230) & (g231) & (!g235) & (g236)) + ((shiftx4x) & (!shiftx5x) & (!g230) & (g231) & (g235) & (!g236)) + ((shiftx4x) & (!shiftx5x) & (!g230) & (g231) & (g235) & (g236)) + ((shiftx4x) & (!shiftx5x) & (g230) & (g231) & (!g235) & (!g236)) + ((shiftx4x) & (!shiftx5x) & (g230) & (g231) & (!g235) & (g236)) + ((shiftx4x) & (!shiftx5x) & (g230) & (g231) & (g235) & (!g236)) + ((shiftx4x) & (!shiftx5x) & (g230) & (g231) & (g235) & (g236)) + ((shiftx4x) & (shiftx5x) & (!g230) & (!g231) & (!g235) & (g236)) + ((shiftx4x) & (shiftx5x) & (!g230) & (!g231) & (g235) & (g236)) + ((shiftx4x) & (shiftx5x) & (!g230) & (g231) & (!g235) & (g236)) + ((shiftx4x) & (shiftx5x) & (!g230) & (g231) & (g235) & (g236)) + ((shiftx4x) & (shiftx5x) & (g230) & (!g231) & (!g235) & (g236)) + ((shiftx4x) & (shiftx5x) & (g230) & (!g231) & (g235) & (g236)) + ((shiftx4x) & (shiftx5x) & (g230) & (g231) & (!g235) & (g236)) + ((shiftx4x) & (shiftx5x) & (g230) & (g231) & (g235) & (g236)));
	assign resultx41x = (((!sk[125]) & (shiftx6x) & (!g380) & (!g381)) + ((!sk[125]) & (shiftx6x) & (!g380) & (g381)) + ((!sk[125]) & (shiftx6x) & (g380) & (!g381)) + ((!sk[125]) & (shiftx6x) & (g380) & (g381)) + ((sk[125]) & (!shiftx6x) & (!g380) & (g381)) + ((sk[125]) & (!shiftx6x) & (g380) & (g381)) + ((sk[125]) & (shiftx6x) & (g380) & (!g381)) + ((sk[125]) & (shiftx6x) & (g380) & (g381)));
	assign g383 = (((!shiftx4x) & (!shiftx5x) & (!g239) & (!g240) & (!g244) & (g245)) + ((!shiftx4x) & (!shiftx5x) & (!g239) & (!g240) & (g244) & (g245)) + ((!shiftx4x) & (!shiftx5x) & (!g239) & (g240) & (!g244) & (g245)) + ((!shiftx4x) & (!shiftx5x) & (!g239) & (g240) & (g244) & (g245)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (!g240) & (!g244) & (g245)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (!g240) & (g244) & (g245)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (g240) & (!g244) & (g245)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (g240) & (g244) & (g245)) + ((!shiftx4x) & (shiftx5x) & (!g239) & (g240) & (!g244) & (!g245)) + ((!shiftx4x) & (shiftx5x) & (!g239) & (g240) & (!g244) & (g245)) + ((!shiftx4x) & (shiftx5x) & (!g239) & (g240) & (g244) & (!g245)) + ((!shiftx4x) & (shiftx5x) & (!g239) & (g240) & (g244) & (g245)) + ((!shiftx4x) & (shiftx5x) & (g239) & (g240) & (!g244) & (!g245)) + ((!shiftx4x) & (shiftx5x) & (g239) & (g240) & (!g244) & (g245)) + ((!shiftx4x) & (shiftx5x) & (g239) & (g240) & (g244) & (!g245)) + ((!shiftx4x) & (shiftx5x) & (g239) & (g240) & (g244) & (g245)) + ((shiftx4x) & (!shiftx5x) & (!g239) & (!g240) & (g244) & (!g245)) + ((shiftx4x) & (!shiftx5x) & (!g239) & (!g240) & (g244) & (g245)) + ((shiftx4x) & (!shiftx5x) & (!g239) & (g240) & (g244) & (!g245)) + ((shiftx4x) & (!shiftx5x) & (!g239) & (g240) & (g244) & (g245)) + ((shiftx4x) & (!shiftx5x) & (g239) & (!g240) & (g244) & (!g245)) + ((shiftx4x) & (!shiftx5x) & (g239) & (!g240) & (g244) & (g245)) + ((shiftx4x) & (!shiftx5x) & (g239) & (g240) & (g244) & (!g245)) + ((shiftx4x) & (!shiftx5x) & (g239) & (g240) & (g244) & (g245)) + ((shiftx4x) & (shiftx5x) & (g239) & (!g240) & (!g244) & (!g245)) + ((shiftx4x) & (shiftx5x) & (g239) & (!g240) & (!g244) & (g245)) + ((shiftx4x) & (shiftx5x) & (g239) & (!g240) & (g244) & (!g245)) + ((shiftx4x) & (shiftx5x) & (g239) & (!g240) & (g244) & (g245)) + ((shiftx4x) & (shiftx5x) & (g239) & (g240) & (!g244) & (!g245)) + ((shiftx4x) & (shiftx5x) & (g239) & (g240) & (!g244) & (g245)) + ((shiftx4x) & (shiftx5x) & (g239) & (g240) & (g244) & (!g245)) + ((shiftx4x) & (shiftx5x) & (g239) & (g240) & (g244) & (g245)));
	assign g384 = (((!shiftx4x) & (!shiftx5x) & (g241) & (!g242) & (!g246) & (!g247)) + ((!shiftx4x) & (!shiftx5x) & (g241) & (!g242) & (!g246) & (g247)) + ((!shiftx4x) & (!shiftx5x) & (g241) & (!g242) & (g246) & (!g247)) + ((!shiftx4x) & (!shiftx5x) & (g241) & (!g242) & (g246) & (g247)) + ((!shiftx4x) & (!shiftx5x) & (g241) & (g242) & (!g246) & (!g247)) + ((!shiftx4x) & (!shiftx5x) & (g241) & (g242) & (!g246) & (g247)) + ((!shiftx4x) & (!shiftx5x) & (g241) & (g242) & (g246) & (!g247)) + ((!shiftx4x) & (!shiftx5x) & (g241) & (g242) & (g246) & (g247)) + ((!shiftx4x) & (shiftx5x) & (!g241) & (!g242) & (g246) & (!g247)) + ((!shiftx4x) & (shiftx5x) & (!g241) & (!g242) & (g246) & (g247)) + ((!shiftx4x) & (shiftx5x) & (!g241) & (g242) & (g246) & (!g247)) + ((!shiftx4x) & (shiftx5x) & (!g241) & (g242) & (g246) & (g247)) + ((!shiftx4x) & (shiftx5x) & (g241) & (!g242) & (g246) & (!g247)) + ((!shiftx4x) & (shiftx5x) & (g241) & (!g242) & (g246) & (g247)) + ((!shiftx4x) & (shiftx5x) & (g241) & (g242) & (g246) & (!g247)) + ((!shiftx4x) & (shiftx5x) & (g241) & (g242) & (g246) & (g247)) + ((shiftx4x) & (!shiftx5x) & (!g241) & (g242) & (!g246) & (!g247)) + ((shiftx4x) & (!shiftx5x) & (!g241) & (g242) & (!g246) & (g247)) + ((shiftx4x) & (!shiftx5x) & (!g241) & (g242) & (g246) & (!g247)) + ((shiftx4x) & (!shiftx5x) & (!g241) & (g242) & (g246) & (g247)) + ((shiftx4x) & (!shiftx5x) & (g241) & (g242) & (!g246) & (!g247)) + ((shiftx4x) & (!shiftx5x) & (g241) & (g242) & (!g246) & (g247)) + ((shiftx4x) & (!shiftx5x) & (g241) & (g242) & (g246) & (!g247)) + ((shiftx4x) & (!shiftx5x) & (g241) & (g242) & (g246) & (g247)) + ((shiftx4x) & (shiftx5x) & (!g241) & (!g242) & (!g246) & (g247)) + ((shiftx4x) & (shiftx5x) & (!g241) & (!g242) & (g246) & (g247)) + ((shiftx4x) & (shiftx5x) & (!g241) & (g242) & (!g246) & (g247)) + ((shiftx4x) & (shiftx5x) & (!g241) & (g242) & (g246) & (g247)) + ((shiftx4x) & (shiftx5x) & (g241) & (!g242) & (!g246) & (g247)) + ((shiftx4x) & (shiftx5x) & (g241) & (!g242) & (g246) & (g247)) + ((shiftx4x) & (shiftx5x) & (g241) & (g242) & (!g246) & (g247)) + ((shiftx4x) & (shiftx5x) & (g241) & (g242) & (g246) & (g247)));
	assign resultx42x = (((!sk[0]) & (shiftx6x) & (!g383) & (!g384)) + ((!sk[0]) & (shiftx6x) & (!g383) & (g384)) + ((!sk[0]) & (shiftx6x) & (g383) & (!g384)) + ((!sk[0]) & (shiftx6x) & (g383) & (g384)) + ((sk[0]) & (!shiftx6x) & (!g383) & (g384)) + ((sk[0]) & (!shiftx6x) & (g383) & (g384)) + ((sk[0]) & (shiftx6x) & (g383) & (!g384)) + ((sk[0]) & (shiftx6x) & (g383) & (g384)));
	assign g386 = (((!shiftx4x) & (!shiftx5x) & (!g250) & (!g251) & (!g255) & (g256)) + ((!shiftx4x) & (!shiftx5x) & (!g250) & (!g251) & (g255) & (g256)) + ((!shiftx4x) & (!shiftx5x) & (!g250) & (g251) & (!g255) & (g256)) + ((!shiftx4x) & (!shiftx5x) & (!g250) & (g251) & (g255) & (g256)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (!g251) & (!g255) & (g256)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (!g251) & (g255) & (g256)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (g251) & (!g255) & (g256)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (g251) & (g255) & (g256)) + ((!shiftx4x) & (shiftx5x) & (!g250) & (g251) & (!g255) & (!g256)) + ((!shiftx4x) & (shiftx5x) & (!g250) & (g251) & (!g255) & (g256)) + ((!shiftx4x) & (shiftx5x) & (!g250) & (g251) & (g255) & (!g256)) + ((!shiftx4x) & (shiftx5x) & (!g250) & (g251) & (g255) & (g256)) + ((!shiftx4x) & (shiftx5x) & (g250) & (g251) & (!g255) & (!g256)) + ((!shiftx4x) & (shiftx5x) & (g250) & (g251) & (!g255) & (g256)) + ((!shiftx4x) & (shiftx5x) & (g250) & (g251) & (g255) & (!g256)) + ((!shiftx4x) & (shiftx5x) & (g250) & (g251) & (g255) & (g256)) + ((shiftx4x) & (!shiftx5x) & (!g250) & (!g251) & (g255) & (!g256)) + ((shiftx4x) & (!shiftx5x) & (!g250) & (!g251) & (g255) & (g256)) + ((shiftx4x) & (!shiftx5x) & (!g250) & (g251) & (g255) & (!g256)) + ((shiftx4x) & (!shiftx5x) & (!g250) & (g251) & (g255) & (g256)) + ((shiftx4x) & (!shiftx5x) & (g250) & (!g251) & (g255) & (!g256)) + ((shiftx4x) & (!shiftx5x) & (g250) & (!g251) & (g255) & (g256)) + ((shiftx4x) & (!shiftx5x) & (g250) & (g251) & (g255) & (!g256)) + ((shiftx4x) & (!shiftx5x) & (g250) & (g251) & (g255) & (g256)) + ((shiftx4x) & (shiftx5x) & (g250) & (!g251) & (!g255) & (!g256)) + ((shiftx4x) & (shiftx5x) & (g250) & (!g251) & (!g255) & (g256)) + ((shiftx4x) & (shiftx5x) & (g250) & (!g251) & (g255) & (!g256)) + ((shiftx4x) & (shiftx5x) & (g250) & (!g251) & (g255) & (g256)) + ((shiftx4x) & (shiftx5x) & (g250) & (g251) & (!g255) & (!g256)) + ((shiftx4x) & (shiftx5x) & (g250) & (g251) & (!g255) & (g256)) + ((shiftx4x) & (shiftx5x) & (g250) & (g251) & (g255) & (!g256)) + ((shiftx4x) & (shiftx5x) & (g250) & (g251) & (g255) & (g256)));
	assign g387 = (((!shiftx4x) & (!shiftx5x) & (g252) & (!g253) & (!g257) & (!g258)) + ((!shiftx4x) & (!shiftx5x) & (g252) & (!g253) & (!g257) & (g258)) + ((!shiftx4x) & (!shiftx5x) & (g252) & (!g253) & (g257) & (!g258)) + ((!shiftx4x) & (!shiftx5x) & (g252) & (!g253) & (g257) & (g258)) + ((!shiftx4x) & (!shiftx5x) & (g252) & (g253) & (!g257) & (!g258)) + ((!shiftx4x) & (!shiftx5x) & (g252) & (g253) & (!g257) & (g258)) + ((!shiftx4x) & (!shiftx5x) & (g252) & (g253) & (g257) & (!g258)) + ((!shiftx4x) & (!shiftx5x) & (g252) & (g253) & (g257) & (g258)) + ((!shiftx4x) & (shiftx5x) & (!g252) & (!g253) & (g257) & (!g258)) + ((!shiftx4x) & (shiftx5x) & (!g252) & (!g253) & (g257) & (g258)) + ((!shiftx4x) & (shiftx5x) & (!g252) & (g253) & (g257) & (!g258)) + ((!shiftx4x) & (shiftx5x) & (!g252) & (g253) & (g257) & (g258)) + ((!shiftx4x) & (shiftx5x) & (g252) & (!g253) & (g257) & (!g258)) + ((!shiftx4x) & (shiftx5x) & (g252) & (!g253) & (g257) & (g258)) + ((!shiftx4x) & (shiftx5x) & (g252) & (g253) & (g257) & (!g258)) + ((!shiftx4x) & (shiftx5x) & (g252) & (g253) & (g257) & (g258)) + ((shiftx4x) & (!shiftx5x) & (!g252) & (g253) & (!g257) & (!g258)) + ((shiftx4x) & (!shiftx5x) & (!g252) & (g253) & (!g257) & (g258)) + ((shiftx4x) & (!shiftx5x) & (!g252) & (g253) & (g257) & (!g258)) + ((shiftx4x) & (!shiftx5x) & (!g252) & (g253) & (g257) & (g258)) + ((shiftx4x) & (!shiftx5x) & (g252) & (g253) & (!g257) & (!g258)) + ((shiftx4x) & (!shiftx5x) & (g252) & (g253) & (!g257) & (g258)) + ((shiftx4x) & (!shiftx5x) & (g252) & (g253) & (g257) & (!g258)) + ((shiftx4x) & (!shiftx5x) & (g252) & (g253) & (g257) & (g258)) + ((shiftx4x) & (shiftx5x) & (!g252) & (!g253) & (!g257) & (g258)) + ((shiftx4x) & (shiftx5x) & (!g252) & (!g253) & (g257) & (g258)) + ((shiftx4x) & (shiftx5x) & (!g252) & (g253) & (!g257) & (g258)) + ((shiftx4x) & (shiftx5x) & (!g252) & (g253) & (g257) & (g258)) + ((shiftx4x) & (shiftx5x) & (g252) & (!g253) & (!g257) & (g258)) + ((shiftx4x) & (shiftx5x) & (g252) & (!g253) & (g257) & (g258)) + ((shiftx4x) & (shiftx5x) & (g252) & (g253) & (!g257) & (g258)) + ((shiftx4x) & (shiftx5x) & (g252) & (g253) & (g257) & (g258)));
	assign resultx43x = (((!shiftx6x) & (sk[3]) & (!g386) & (g387)) + ((!shiftx6x) & (sk[3]) & (g386) & (g387)) + ((shiftx6x) & (!sk[3]) & (!g386) & (!g387)) + ((shiftx6x) & (!sk[3]) & (!g386) & (g387)) + ((shiftx6x) & (!sk[3]) & (g386) & (!g387)) + ((shiftx6x) & (!sk[3]) & (g386) & (g387)) + ((shiftx6x) & (sk[3]) & (g386) & (!g387)) + ((shiftx6x) & (sk[3]) & (g386) & (g387)));
	assign g389 = (((!shiftx4x) & (!shiftx5x) & (!g261) & (!g262) & (!g266) & (g267)) + ((!shiftx4x) & (!shiftx5x) & (!g261) & (!g262) & (g266) & (g267)) + ((!shiftx4x) & (!shiftx5x) & (!g261) & (g262) & (!g266) & (g267)) + ((!shiftx4x) & (!shiftx5x) & (!g261) & (g262) & (g266) & (g267)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (!g262) & (!g266) & (g267)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (!g262) & (g266) & (g267)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (g262) & (!g266) & (g267)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (g262) & (g266) & (g267)) + ((!shiftx4x) & (shiftx5x) & (!g261) & (g262) & (!g266) & (!g267)) + ((!shiftx4x) & (shiftx5x) & (!g261) & (g262) & (!g266) & (g267)) + ((!shiftx4x) & (shiftx5x) & (!g261) & (g262) & (g266) & (!g267)) + ((!shiftx4x) & (shiftx5x) & (!g261) & (g262) & (g266) & (g267)) + ((!shiftx4x) & (shiftx5x) & (g261) & (g262) & (!g266) & (!g267)) + ((!shiftx4x) & (shiftx5x) & (g261) & (g262) & (!g266) & (g267)) + ((!shiftx4x) & (shiftx5x) & (g261) & (g262) & (g266) & (!g267)) + ((!shiftx4x) & (shiftx5x) & (g261) & (g262) & (g266) & (g267)) + ((shiftx4x) & (!shiftx5x) & (!g261) & (!g262) & (g266) & (!g267)) + ((shiftx4x) & (!shiftx5x) & (!g261) & (!g262) & (g266) & (g267)) + ((shiftx4x) & (!shiftx5x) & (!g261) & (g262) & (g266) & (!g267)) + ((shiftx4x) & (!shiftx5x) & (!g261) & (g262) & (g266) & (g267)) + ((shiftx4x) & (!shiftx5x) & (g261) & (!g262) & (g266) & (!g267)) + ((shiftx4x) & (!shiftx5x) & (g261) & (!g262) & (g266) & (g267)) + ((shiftx4x) & (!shiftx5x) & (g261) & (g262) & (g266) & (!g267)) + ((shiftx4x) & (!shiftx5x) & (g261) & (g262) & (g266) & (g267)) + ((shiftx4x) & (shiftx5x) & (g261) & (!g262) & (!g266) & (!g267)) + ((shiftx4x) & (shiftx5x) & (g261) & (!g262) & (!g266) & (g267)) + ((shiftx4x) & (shiftx5x) & (g261) & (!g262) & (g266) & (!g267)) + ((shiftx4x) & (shiftx5x) & (g261) & (!g262) & (g266) & (g267)) + ((shiftx4x) & (shiftx5x) & (g261) & (g262) & (!g266) & (!g267)) + ((shiftx4x) & (shiftx5x) & (g261) & (g262) & (!g266) & (g267)) + ((shiftx4x) & (shiftx5x) & (g261) & (g262) & (g266) & (!g267)) + ((shiftx4x) & (shiftx5x) & (g261) & (g262) & (g266) & (g267)));
	assign g390 = (((!shiftx4x) & (!shiftx5x) & (g263) & (!g264) & (!g268) & (!g269)) + ((!shiftx4x) & (!shiftx5x) & (g263) & (!g264) & (!g268) & (g269)) + ((!shiftx4x) & (!shiftx5x) & (g263) & (!g264) & (g268) & (!g269)) + ((!shiftx4x) & (!shiftx5x) & (g263) & (!g264) & (g268) & (g269)) + ((!shiftx4x) & (!shiftx5x) & (g263) & (g264) & (!g268) & (!g269)) + ((!shiftx4x) & (!shiftx5x) & (g263) & (g264) & (!g268) & (g269)) + ((!shiftx4x) & (!shiftx5x) & (g263) & (g264) & (g268) & (!g269)) + ((!shiftx4x) & (!shiftx5x) & (g263) & (g264) & (g268) & (g269)) + ((!shiftx4x) & (shiftx5x) & (!g263) & (!g264) & (g268) & (!g269)) + ((!shiftx4x) & (shiftx5x) & (!g263) & (!g264) & (g268) & (g269)) + ((!shiftx4x) & (shiftx5x) & (!g263) & (g264) & (g268) & (!g269)) + ((!shiftx4x) & (shiftx5x) & (!g263) & (g264) & (g268) & (g269)) + ((!shiftx4x) & (shiftx5x) & (g263) & (!g264) & (g268) & (!g269)) + ((!shiftx4x) & (shiftx5x) & (g263) & (!g264) & (g268) & (g269)) + ((!shiftx4x) & (shiftx5x) & (g263) & (g264) & (g268) & (!g269)) + ((!shiftx4x) & (shiftx5x) & (g263) & (g264) & (g268) & (g269)) + ((shiftx4x) & (!shiftx5x) & (!g263) & (g264) & (!g268) & (!g269)) + ((shiftx4x) & (!shiftx5x) & (!g263) & (g264) & (!g268) & (g269)) + ((shiftx4x) & (!shiftx5x) & (!g263) & (g264) & (g268) & (!g269)) + ((shiftx4x) & (!shiftx5x) & (!g263) & (g264) & (g268) & (g269)) + ((shiftx4x) & (!shiftx5x) & (g263) & (g264) & (!g268) & (!g269)) + ((shiftx4x) & (!shiftx5x) & (g263) & (g264) & (!g268) & (g269)) + ((shiftx4x) & (!shiftx5x) & (g263) & (g264) & (g268) & (!g269)) + ((shiftx4x) & (!shiftx5x) & (g263) & (g264) & (g268) & (g269)) + ((shiftx4x) & (shiftx5x) & (!g263) & (!g264) & (!g268) & (g269)) + ((shiftx4x) & (shiftx5x) & (!g263) & (!g264) & (g268) & (g269)) + ((shiftx4x) & (shiftx5x) & (!g263) & (g264) & (!g268) & (g269)) + ((shiftx4x) & (shiftx5x) & (!g263) & (g264) & (g268) & (g269)) + ((shiftx4x) & (shiftx5x) & (g263) & (!g264) & (!g268) & (g269)) + ((shiftx4x) & (shiftx5x) & (g263) & (!g264) & (g268) & (g269)) + ((shiftx4x) & (shiftx5x) & (g263) & (g264) & (!g268) & (g269)) + ((shiftx4x) & (shiftx5x) & (g263) & (g264) & (g268) & (g269)));
	assign resultx44x = (((!shiftx6x) & (!g389) & (sk[6]) & (g390)) + ((!shiftx6x) & (g389) & (sk[6]) & (g390)) + ((shiftx6x) & (!g389) & (!sk[6]) & (!g390)) + ((shiftx6x) & (!g389) & (!sk[6]) & (g390)) + ((shiftx6x) & (g389) & (!sk[6]) & (!g390)) + ((shiftx6x) & (g389) & (!sk[6]) & (g390)) + ((shiftx6x) & (g389) & (sk[6]) & (!g390)) + ((shiftx6x) & (g389) & (sk[6]) & (g390)));
	assign g392 = (((!shiftx4x) & (!shiftx5x) & (!g272) & (!g273) & (!g277) & (g278)) + ((!shiftx4x) & (!shiftx5x) & (!g272) & (!g273) & (g277) & (g278)) + ((!shiftx4x) & (!shiftx5x) & (!g272) & (g273) & (!g277) & (g278)) + ((!shiftx4x) & (!shiftx5x) & (!g272) & (g273) & (g277) & (g278)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (!g273) & (!g277) & (g278)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (!g273) & (g277) & (g278)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (g273) & (!g277) & (g278)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (g273) & (g277) & (g278)) + ((!shiftx4x) & (shiftx5x) & (!g272) & (g273) & (!g277) & (!g278)) + ((!shiftx4x) & (shiftx5x) & (!g272) & (g273) & (!g277) & (g278)) + ((!shiftx4x) & (shiftx5x) & (!g272) & (g273) & (g277) & (!g278)) + ((!shiftx4x) & (shiftx5x) & (!g272) & (g273) & (g277) & (g278)) + ((!shiftx4x) & (shiftx5x) & (g272) & (g273) & (!g277) & (!g278)) + ((!shiftx4x) & (shiftx5x) & (g272) & (g273) & (!g277) & (g278)) + ((!shiftx4x) & (shiftx5x) & (g272) & (g273) & (g277) & (!g278)) + ((!shiftx4x) & (shiftx5x) & (g272) & (g273) & (g277) & (g278)) + ((shiftx4x) & (!shiftx5x) & (!g272) & (!g273) & (g277) & (!g278)) + ((shiftx4x) & (!shiftx5x) & (!g272) & (!g273) & (g277) & (g278)) + ((shiftx4x) & (!shiftx5x) & (!g272) & (g273) & (g277) & (!g278)) + ((shiftx4x) & (!shiftx5x) & (!g272) & (g273) & (g277) & (g278)) + ((shiftx4x) & (!shiftx5x) & (g272) & (!g273) & (g277) & (!g278)) + ((shiftx4x) & (!shiftx5x) & (g272) & (!g273) & (g277) & (g278)) + ((shiftx4x) & (!shiftx5x) & (g272) & (g273) & (g277) & (!g278)) + ((shiftx4x) & (!shiftx5x) & (g272) & (g273) & (g277) & (g278)) + ((shiftx4x) & (shiftx5x) & (g272) & (!g273) & (!g277) & (!g278)) + ((shiftx4x) & (shiftx5x) & (g272) & (!g273) & (!g277) & (g278)) + ((shiftx4x) & (shiftx5x) & (g272) & (!g273) & (g277) & (!g278)) + ((shiftx4x) & (shiftx5x) & (g272) & (!g273) & (g277) & (g278)) + ((shiftx4x) & (shiftx5x) & (g272) & (g273) & (!g277) & (!g278)) + ((shiftx4x) & (shiftx5x) & (g272) & (g273) & (!g277) & (g278)) + ((shiftx4x) & (shiftx5x) & (g272) & (g273) & (g277) & (!g278)) + ((shiftx4x) & (shiftx5x) & (g272) & (g273) & (g277) & (g278)));
	assign g393 = (((!shiftx4x) & (!shiftx5x) & (g274) & (!g275) & (!g279) & (!g280)) + ((!shiftx4x) & (!shiftx5x) & (g274) & (!g275) & (!g279) & (g280)) + ((!shiftx4x) & (!shiftx5x) & (g274) & (!g275) & (g279) & (!g280)) + ((!shiftx4x) & (!shiftx5x) & (g274) & (!g275) & (g279) & (g280)) + ((!shiftx4x) & (!shiftx5x) & (g274) & (g275) & (!g279) & (!g280)) + ((!shiftx4x) & (!shiftx5x) & (g274) & (g275) & (!g279) & (g280)) + ((!shiftx4x) & (!shiftx5x) & (g274) & (g275) & (g279) & (!g280)) + ((!shiftx4x) & (!shiftx5x) & (g274) & (g275) & (g279) & (g280)) + ((!shiftx4x) & (shiftx5x) & (!g274) & (!g275) & (g279) & (!g280)) + ((!shiftx4x) & (shiftx5x) & (!g274) & (!g275) & (g279) & (g280)) + ((!shiftx4x) & (shiftx5x) & (!g274) & (g275) & (g279) & (!g280)) + ((!shiftx4x) & (shiftx5x) & (!g274) & (g275) & (g279) & (g280)) + ((!shiftx4x) & (shiftx5x) & (g274) & (!g275) & (g279) & (!g280)) + ((!shiftx4x) & (shiftx5x) & (g274) & (!g275) & (g279) & (g280)) + ((!shiftx4x) & (shiftx5x) & (g274) & (g275) & (g279) & (!g280)) + ((!shiftx4x) & (shiftx5x) & (g274) & (g275) & (g279) & (g280)) + ((shiftx4x) & (!shiftx5x) & (!g274) & (g275) & (!g279) & (!g280)) + ((shiftx4x) & (!shiftx5x) & (!g274) & (g275) & (!g279) & (g280)) + ((shiftx4x) & (!shiftx5x) & (!g274) & (g275) & (g279) & (!g280)) + ((shiftx4x) & (!shiftx5x) & (!g274) & (g275) & (g279) & (g280)) + ((shiftx4x) & (!shiftx5x) & (g274) & (g275) & (!g279) & (!g280)) + ((shiftx4x) & (!shiftx5x) & (g274) & (g275) & (!g279) & (g280)) + ((shiftx4x) & (!shiftx5x) & (g274) & (g275) & (g279) & (!g280)) + ((shiftx4x) & (!shiftx5x) & (g274) & (g275) & (g279) & (g280)) + ((shiftx4x) & (shiftx5x) & (!g274) & (!g275) & (!g279) & (g280)) + ((shiftx4x) & (shiftx5x) & (!g274) & (!g275) & (g279) & (g280)) + ((shiftx4x) & (shiftx5x) & (!g274) & (g275) & (!g279) & (g280)) + ((shiftx4x) & (shiftx5x) & (!g274) & (g275) & (g279) & (g280)) + ((shiftx4x) & (shiftx5x) & (g274) & (!g275) & (!g279) & (g280)) + ((shiftx4x) & (shiftx5x) & (g274) & (!g275) & (g279) & (g280)) + ((shiftx4x) & (shiftx5x) & (g274) & (g275) & (!g279) & (g280)) + ((shiftx4x) & (shiftx5x) & (g274) & (g275) & (g279) & (g280)));
	assign resultx45x = (((!sk[9]) & (shiftx6x) & (!g392) & (!g393)) + ((!sk[9]) & (shiftx6x) & (!g392) & (g393)) + ((!sk[9]) & (shiftx6x) & (g392) & (!g393)) + ((!sk[9]) & (shiftx6x) & (g392) & (g393)) + ((sk[9]) & (!shiftx6x) & (!g392) & (g393)) + ((sk[9]) & (!shiftx6x) & (g392) & (g393)) + ((sk[9]) & (shiftx6x) & (g392) & (!g393)) + ((sk[9]) & (shiftx6x) & (g392) & (g393)));
	assign g395 = (((!shiftx4x) & (!shiftx5x) & (!g283) & (!g284) & (!g288) & (g289)) + ((!shiftx4x) & (!shiftx5x) & (!g283) & (!g284) & (g288) & (g289)) + ((!shiftx4x) & (!shiftx5x) & (!g283) & (g284) & (!g288) & (g289)) + ((!shiftx4x) & (!shiftx5x) & (!g283) & (g284) & (g288) & (g289)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (!g284) & (!g288) & (g289)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (!g284) & (g288) & (g289)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (g284) & (!g288) & (g289)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (g284) & (g288) & (g289)) + ((!shiftx4x) & (shiftx5x) & (!g283) & (g284) & (!g288) & (!g289)) + ((!shiftx4x) & (shiftx5x) & (!g283) & (g284) & (!g288) & (g289)) + ((!shiftx4x) & (shiftx5x) & (!g283) & (g284) & (g288) & (!g289)) + ((!shiftx4x) & (shiftx5x) & (!g283) & (g284) & (g288) & (g289)) + ((!shiftx4x) & (shiftx5x) & (g283) & (g284) & (!g288) & (!g289)) + ((!shiftx4x) & (shiftx5x) & (g283) & (g284) & (!g288) & (g289)) + ((!shiftx4x) & (shiftx5x) & (g283) & (g284) & (g288) & (!g289)) + ((!shiftx4x) & (shiftx5x) & (g283) & (g284) & (g288) & (g289)) + ((shiftx4x) & (!shiftx5x) & (!g283) & (!g284) & (g288) & (!g289)) + ((shiftx4x) & (!shiftx5x) & (!g283) & (!g284) & (g288) & (g289)) + ((shiftx4x) & (!shiftx5x) & (!g283) & (g284) & (g288) & (!g289)) + ((shiftx4x) & (!shiftx5x) & (!g283) & (g284) & (g288) & (g289)) + ((shiftx4x) & (!shiftx5x) & (g283) & (!g284) & (g288) & (!g289)) + ((shiftx4x) & (!shiftx5x) & (g283) & (!g284) & (g288) & (g289)) + ((shiftx4x) & (!shiftx5x) & (g283) & (g284) & (g288) & (!g289)) + ((shiftx4x) & (!shiftx5x) & (g283) & (g284) & (g288) & (g289)) + ((shiftx4x) & (shiftx5x) & (g283) & (!g284) & (!g288) & (!g289)) + ((shiftx4x) & (shiftx5x) & (g283) & (!g284) & (!g288) & (g289)) + ((shiftx4x) & (shiftx5x) & (g283) & (!g284) & (g288) & (!g289)) + ((shiftx4x) & (shiftx5x) & (g283) & (!g284) & (g288) & (g289)) + ((shiftx4x) & (shiftx5x) & (g283) & (g284) & (!g288) & (!g289)) + ((shiftx4x) & (shiftx5x) & (g283) & (g284) & (!g288) & (g289)) + ((shiftx4x) & (shiftx5x) & (g283) & (g284) & (g288) & (!g289)) + ((shiftx4x) & (shiftx5x) & (g283) & (g284) & (g288) & (g289)));
	assign g396 = (((!shiftx4x) & (!shiftx5x) & (g285) & (!g286) & (!g290) & (!g291)) + ((!shiftx4x) & (!shiftx5x) & (g285) & (!g286) & (!g290) & (g291)) + ((!shiftx4x) & (!shiftx5x) & (g285) & (!g286) & (g290) & (!g291)) + ((!shiftx4x) & (!shiftx5x) & (g285) & (!g286) & (g290) & (g291)) + ((!shiftx4x) & (!shiftx5x) & (g285) & (g286) & (!g290) & (!g291)) + ((!shiftx4x) & (!shiftx5x) & (g285) & (g286) & (!g290) & (g291)) + ((!shiftx4x) & (!shiftx5x) & (g285) & (g286) & (g290) & (!g291)) + ((!shiftx4x) & (!shiftx5x) & (g285) & (g286) & (g290) & (g291)) + ((!shiftx4x) & (shiftx5x) & (!g285) & (!g286) & (g290) & (!g291)) + ((!shiftx4x) & (shiftx5x) & (!g285) & (!g286) & (g290) & (g291)) + ((!shiftx4x) & (shiftx5x) & (!g285) & (g286) & (g290) & (!g291)) + ((!shiftx4x) & (shiftx5x) & (!g285) & (g286) & (g290) & (g291)) + ((!shiftx4x) & (shiftx5x) & (g285) & (!g286) & (g290) & (!g291)) + ((!shiftx4x) & (shiftx5x) & (g285) & (!g286) & (g290) & (g291)) + ((!shiftx4x) & (shiftx5x) & (g285) & (g286) & (g290) & (!g291)) + ((!shiftx4x) & (shiftx5x) & (g285) & (g286) & (g290) & (g291)) + ((shiftx4x) & (!shiftx5x) & (!g285) & (g286) & (!g290) & (!g291)) + ((shiftx4x) & (!shiftx5x) & (!g285) & (g286) & (!g290) & (g291)) + ((shiftx4x) & (!shiftx5x) & (!g285) & (g286) & (g290) & (!g291)) + ((shiftx4x) & (!shiftx5x) & (!g285) & (g286) & (g290) & (g291)) + ((shiftx4x) & (!shiftx5x) & (g285) & (g286) & (!g290) & (!g291)) + ((shiftx4x) & (!shiftx5x) & (g285) & (g286) & (!g290) & (g291)) + ((shiftx4x) & (!shiftx5x) & (g285) & (g286) & (g290) & (!g291)) + ((shiftx4x) & (!shiftx5x) & (g285) & (g286) & (g290) & (g291)) + ((shiftx4x) & (shiftx5x) & (!g285) & (!g286) & (!g290) & (g291)) + ((shiftx4x) & (shiftx5x) & (!g285) & (!g286) & (g290) & (g291)) + ((shiftx4x) & (shiftx5x) & (!g285) & (g286) & (!g290) & (g291)) + ((shiftx4x) & (shiftx5x) & (!g285) & (g286) & (g290) & (g291)) + ((shiftx4x) & (shiftx5x) & (g285) & (!g286) & (!g290) & (g291)) + ((shiftx4x) & (shiftx5x) & (g285) & (!g286) & (g290) & (g291)) + ((shiftx4x) & (shiftx5x) & (g285) & (g286) & (!g290) & (g291)) + ((shiftx4x) & (shiftx5x) & (g285) & (g286) & (g290) & (g291)));
	assign resultx46x = (((!shiftx6x) & (sk[12]) & (!g395) & (g396)) + ((!shiftx6x) & (sk[12]) & (g395) & (g396)) + ((shiftx6x) & (!sk[12]) & (!g395) & (!g396)) + ((shiftx6x) & (!sk[12]) & (!g395) & (g396)) + ((shiftx6x) & (!sk[12]) & (g395) & (!g396)) + ((shiftx6x) & (!sk[12]) & (g395) & (g396)) + ((shiftx6x) & (sk[12]) & (g395) & (!g396)) + ((shiftx6x) & (sk[12]) & (g395) & (g396)));
	assign g398 = (((!shiftx4x) & (!shiftx5x) & (!g294) & (!g295) & (!g299) & (g300)) + ((!shiftx4x) & (!shiftx5x) & (!g294) & (!g295) & (g299) & (g300)) + ((!shiftx4x) & (!shiftx5x) & (!g294) & (g295) & (!g299) & (g300)) + ((!shiftx4x) & (!shiftx5x) & (!g294) & (g295) & (g299) & (g300)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (!g295) & (!g299) & (g300)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (!g295) & (g299) & (g300)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (g295) & (!g299) & (g300)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (g295) & (g299) & (g300)) + ((!shiftx4x) & (shiftx5x) & (!g294) & (g295) & (!g299) & (!g300)) + ((!shiftx4x) & (shiftx5x) & (!g294) & (g295) & (!g299) & (g300)) + ((!shiftx4x) & (shiftx5x) & (!g294) & (g295) & (g299) & (!g300)) + ((!shiftx4x) & (shiftx5x) & (!g294) & (g295) & (g299) & (g300)) + ((!shiftx4x) & (shiftx5x) & (g294) & (g295) & (!g299) & (!g300)) + ((!shiftx4x) & (shiftx5x) & (g294) & (g295) & (!g299) & (g300)) + ((!shiftx4x) & (shiftx5x) & (g294) & (g295) & (g299) & (!g300)) + ((!shiftx4x) & (shiftx5x) & (g294) & (g295) & (g299) & (g300)) + ((shiftx4x) & (!shiftx5x) & (!g294) & (!g295) & (g299) & (!g300)) + ((shiftx4x) & (!shiftx5x) & (!g294) & (!g295) & (g299) & (g300)) + ((shiftx4x) & (!shiftx5x) & (!g294) & (g295) & (g299) & (!g300)) + ((shiftx4x) & (!shiftx5x) & (!g294) & (g295) & (g299) & (g300)) + ((shiftx4x) & (!shiftx5x) & (g294) & (!g295) & (g299) & (!g300)) + ((shiftx4x) & (!shiftx5x) & (g294) & (!g295) & (g299) & (g300)) + ((shiftx4x) & (!shiftx5x) & (g294) & (g295) & (g299) & (!g300)) + ((shiftx4x) & (!shiftx5x) & (g294) & (g295) & (g299) & (g300)) + ((shiftx4x) & (shiftx5x) & (g294) & (!g295) & (!g299) & (!g300)) + ((shiftx4x) & (shiftx5x) & (g294) & (!g295) & (!g299) & (g300)) + ((shiftx4x) & (shiftx5x) & (g294) & (!g295) & (g299) & (!g300)) + ((shiftx4x) & (shiftx5x) & (g294) & (!g295) & (g299) & (g300)) + ((shiftx4x) & (shiftx5x) & (g294) & (g295) & (!g299) & (!g300)) + ((shiftx4x) & (shiftx5x) & (g294) & (g295) & (!g299) & (g300)) + ((shiftx4x) & (shiftx5x) & (g294) & (g295) & (g299) & (!g300)) + ((shiftx4x) & (shiftx5x) & (g294) & (g295) & (g299) & (g300)));
	assign g399 = (((!shiftx4x) & (!shiftx5x) & (g296) & (!g297) & (!g301) & (!g302)) + ((!shiftx4x) & (!shiftx5x) & (g296) & (!g297) & (!g301) & (g302)) + ((!shiftx4x) & (!shiftx5x) & (g296) & (!g297) & (g301) & (!g302)) + ((!shiftx4x) & (!shiftx5x) & (g296) & (!g297) & (g301) & (g302)) + ((!shiftx4x) & (!shiftx5x) & (g296) & (g297) & (!g301) & (!g302)) + ((!shiftx4x) & (!shiftx5x) & (g296) & (g297) & (!g301) & (g302)) + ((!shiftx4x) & (!shiftx5x) & (g296) & (g297) & (g301) & (!g302)) + ((!shiftx4x) & (!shiftx5x) & (g296) & (g297) & (g301) & (g302)) + ((!shiftx4x) & (shiftx5x) & (!g296) & (!g297) & (g301) & (!g302)) + ((!shiftx4x) & (shiftx5x) & (!g296) & (!g297) & (g301) & (g302)) + ((!shiftx4x) & (shiftx5x) & (!g296) & (g297) & (g301) & (!g302)) + ((!shiftx4x) & (shiftx5x) & (!g296) & (g297) & (g301) & (g302)) + ((!shiftx4x) & (shiftx5x) & (g296) & (!g297) & (g301) & (!g302)) + ((!shiftx4x) & (shiftx5x) & (g296) & (!g297) & (g301) & (g302)) + ((!shiftx4x) & (shiftx5x) & (g296) & (g297) & (g301) & (!g302)) + ((!shiftx4x) & (shiftx5x) & (g296) & (g297) & (g301) & (g302)) + ((shiftx4x) & (!shiftx5x) & (!g296) & (g297) & (!g301) & (!g302)) + ((shiftx4x) & (!shiftx5x) & (!g296) & (g297) & (!g301) & (g302)) + ((shiftx4x) & (!shiftx5x) & (!g296) & (g297) & (g301) & (!g302)) + ((shiftx4x) & (!shiftx5x) & (!g296) & (g297) & (g301) & (g302)) + ((shiftx4x) & (!shiftx5x) & (g296) & (g297) & (!g301) & (!g302)) + ((shiftx4x) & (!shiftx5x) & (g296) & (g297) & (!g301) & (g302)) + ((shiftx4x) & (!shiftx5x) & (g296) & (g297) & (g301) & (!g302)) + ((shiftx4x) & (!shiftx5x) & (g296) & (g297) & (g301) & (g302)) + ((shiftx4x) & (shiftx5x) & (!g296) & (!g297) & (!g301) & (g302)) + ((shiftx4x) & (shiftx5x) & (!g296) & (!g297) & (g301) & (g302)) + ((shiftx4x) & (shiftx5x) & (!g296) & (g297) & (!g301) & (g302)) + ((shiftx4x) & (shiftx5x) & (!g296) & (g297) & (g301) & (g302)) + ((shiftx4x) & (shiftx5x) & (g296) & (!g297) & (!g301) & (g302)) + ((shiftx4x) & (shiftx5x) & (g296) & (!g297) & (g301) & (g302)) + ((shiftx4x) & (shiftx5x) & (g296) & (g297) & (!g301) & (g302)) + ((shiftx4x) & (shiftx5x) & (g296) & (g297) & (g301) & (g302)));
	assign resultx47x = (((!shiftx6x) & (sk[15]) & (!g398) & (g399)) + ((!shiftx6x) & (sk[15]) & (g398) & (g399)) + ((shiftx6x) & (!sk[15]) & (!g398) & (!g399)) + ((shiftx6x) & (!sk[15]) & (!g398) & (g399)) + ((shiftx6x) & (!sk[15]) & (g398) & (!g399)) + ((shiftx6x) & (!sk[15]) & (g398) & (g399)) + ((shiftx6x) & (sk[15]) & (g398) & (!g399)) + ((shiftx6x) & (sk[15]) & (g398) & (g399)));
	assign g401 = (((!shiftx4x) & (!shiftx5x) & (!g15) & (!g26) & (!g31) & (g41)) + ((!shiftx4x) & (!shiftx5x) & (!g15) & (!g26) & (g31) & (g41)) + ((!shiftx4x) & (!shiftx5x) & (!g15) & (g26) & (!g31) & (g41)) + ((!shiftx4x) & (!shiftx5x) & (!g15) & (g26) & (g31) & (g41)) + ((!shiftx4x) & (!shiftx5x) & (g15) & (!g26) & (!g31) & (g41)) + ((!shiftx4x) & (!shiftx5x) & (g15) & (!g26) & (g31) & (g41)) + ((!shiftx4x) & (!shiftx5x) & (g15) & (g26) & (!g31) & (g41)) + ((!shiftx4x) & (!shiftx5x) & (g15) & (g26) & (g31) & (g41)) + ((!shiftx4x) & (shiftx5x) & (!g15) & (g26) & (!g31) & (!g41)) + ((!shiftx4x) & (shiftx5x) & (!g15) & (g26) & (!g31) & (g41)) + ((!shiftx4x) & (shiftx5x) & (!g15) & (g26) & (g31) & (!g41)) + ((!shiftx4x) & (shiftx5x) & (!g15) & (g26) & (g31) & (g41)) + ((!shiftx4x) & (shiftx5x) & (g15) & (g26) & (!g31) & (!g41)) + ((!shiftx4x) & (shiftx5x) & (g15) & (g26) & (!g31) & (g41)) + ((!shiftx4x) & (shiftx5x) & (g15) & (g26) & (g31) & (!g41)) + ((!shiftx4x) & (shiftx5x) & (g15) & (g26) & (g31) & (g41)) + ((shiftx4x) & (!shiftx5x) & (!g15) & (!g26) & (g31) & (!g41)) + ((shiftx4x) & (!shiftx5x) & (!g15) & (!g26) & (g31) & (g41)) + ((shiftx4x) & (!shiftx5x) & (!g15) & (g26) & (g31) & (!g41)) + ((shiftx4x) & (!shiftx5x) & (!g15) & (g26) & (g31) & (g41)) + ((shiftx4x) & (!shiftx5x) & (g15) & (!g26) & (g31) & (!g41)) + ((shiftx4x) & (!shiftx5x) & (g15) & (!g26) & (g31) & (g41)) + ((shiftx4x) & (!shiftx5x) & (g15) & (g26) & (g31) & (!g41)) + ((shiftx4x) & (!shiftx5x) & (g15) & (g26) & (g31) & (g41)) + ((shiftx4x) & (shiftx5x) & (g15) & (!g26) & (!g31) & (!g41)) + ((shiftx4x) & (shiftx5x) & (g15) & (!g26) & (!g31) & (g41)) + ((shiftx4x) & (shiftx5x) & (g15) & (!g26) & (g31) & (!g41)) + ((shiftx4x) & (shiftx5x) & (g15) & (!g26) & (g31) & (g41)) + ((shiftx4x) & (shiftx5x) & (g15) & (g26) & (!g31) & (!g41)) + ((shiftx4x) & (shiftx5x) & (g15) & (g26) & (!g31) & (g41)) + ((shiftx4x) & (shiftx5x) & (g15) & (g26) & (g31) & (!g41)) + ((shiftx4x) & (shiftx5x) & (g15) & (g26) & (g31) & (g41)));
	assign g402 = (((!shiftx4x) & (!shiftx5x) & (!g5) & (!g10) & (g20) & (!g36)) + ((!shiftx4x) & (!shiftx5x) & (!g5) & (!g10) & (g20) & (g36)) + ((!shiftx4x) & (!shiftx5x) & (!g5) & (g10) & (g20) & (!g36)) + ((!shiftx4x) & (!shiftx5x) & (!g5) & (g10) & (g20) & (g36)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (!g10) & (g20) & (!g36)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (!g10) & (g20) & (g36)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (g10) & (g20) & (!g36)) + ((!shiftx4x) & (!shiftx5x) & (g5) & (g10) & (g20) & (g36)) + ((!shiftx4x) & (shiftx5x) & (g5) & (!g10) & (!g20) & (!g36)) + ((!shiftx4x) & (shiftx5x) & (g5) & (!g10) & (!g20) & (g36)) + ((!shiftx4x) & (shiftx5x) & (g5) & (!g10) & (g20) & (!g36)) + ((!shiftx4x) & (shiftx5x) & (g5) & (!g10) & (g20) & (g36)) + ((!shiftx4x) & (shiftx5x) & (g5) & (g10) & (!g20) & (!g36)) + ((!shiftx4x) & (shiftx5x) & (g5) & (g10) & (!g20) & (g36)) + ((!shiftx4x) & (shiftx5x) & (g5) & (g10) & (g20) & (!g36)) + ((!shiftx4x) & (shiftx5x) & (g5) & (g10) & (g20) & (g36)) + ((shiftx4x) & (!shiftx5x) & (!g5) & (g10) & (!g20) & (!g36)) + ((shiftx4x) & (!shiftx5x) & (!g5) & (g10) & (!g20) & (g36)) + ((shiftx4x) & (!shiftx5x) & (!g5) & (g10) & (g20) & (!g36)) + ((shiftx4x) & (!shiftx5x) & (!g5) & (g10) & (g20) & (g36)) + ((shiftx4x) & (!shiftx5x) & (g5) & (g10) & (!g20) & (!g36)) + ((shiftx4x) & (!shiftx5x) & (g5) & (g10) & (!g20) & (g36)) + ((shiftx4x) & (!shiftx5x) & (g5) & (g10) & (g20) & (!g36)) + ((shiftx4x) & (!shiftx5x) & (g5) & (g10) & (g20) & (g36)) + ((shiftx4x) & (shiftx5x) & (!g5) & (!g10) & (!g20) & (g36)) + ((shiftx4x) & (shiftx5x) & (!g5) & (!g10) & (g20) & (g36)) + ((shiftx4x) & (shiftx5x) & (!g5) & (g10) & (!g20) & (g36)) + ((shiftx4x) & (shiftx5x) & (!g5) & (g10) & (g20) & (g36)) + ((shiftx4x) & (shiftx5x) & (g5) & (!g10) & (!g20) & (g36)) + ((shiftx4x) & (shiftx5x) & (g5) & (!g10) & (g20) & (g36)) + ((shiftx4x) & (shiftx5x) & (g5) & (g10) & (!g20) & (g36)) + ((shiftx4x) & (shiftx5x) & (g5) & (g10) & (g20) & (g36)));
	assign resultx48x = (((!shiftx6x) & (!g401) & (sk[18]) & (g402)) + ((!shiftx6x) & (g401) & (sk[18]) & (g402)) + ((shiftx6x) & (!g401) & (!sk[18]) & (!g402)) + ((shiftx6x) & (!g401) & (!sk[18]) & (g402)) + ((shiftx6x) & (g401) & (!sk[18]) & (!g402)) + ((shiftx6x) & (g401) & (!sk[18]) & (g402)) + ((shiftx6x) & (g401) & (sk[18]) & (!g402)) + ((shiftx6x) & (g401) & (sk[18]) & (g402)));
	assign g404 = (((!shiftx4x) & (!shiftx5x) & (!g48) & (!g69) & (!g74) & (g84)) + ((!shiftx4x) & (!shiftx5x) & (!g48) & (!g69) & (g74) & (g84)) + ((!shiftx4x) & (!shiftx5x) & (!g48) & (g69) & (!g74) & (g84)) + ((!shiftx4x) & (!shiftx5x) & (!g48) & (g69) & (g74) & (g84)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (!g69) & (!g74) & (g84)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (!g69) & (g74) & (g84)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (g69) & (!g74) & (g84)) + ((!shiftx4x) & (!shiftx5x) & (g48) & (g69) & (g74) & (g84)) + ((!shiftx4x) & (shiftx5x) & (!g48) & (g69) & (!g74) & (!g84)) + ((!shiftx4x) & (shiftx5x) & (!g48) & (g69) & (!g74) & (g84)) + ((!shiftx4x) & (shiftx5x) & (!g48) & (g69) & (g74) & (!g84)) + ((!shiftx4x) & (shiftx5x) & (!g48) & (g69) & (g74) & (g84)) + ((!shiftx4x) & (shiftx5x) & (g48) & (g69) & (!g74) & (!g84)) + ((!shiftx4x) & (shiftx5x) & (g48) & (g69) & (!g74) & (g84)) + ((!shiftx4x) & (shiftx5x) & (g48) & (g69) & (g74) & (!g84)) + ((!shiftx4x) & (shiftx5x) & (g48) & (g69) & (g74) & (g84)) + ((shiftx4x) & (!shiftx5x) & (!g48) & (!g69) & (g74) & (!g84)) + ((shiftx4x) & (!shiftx5x) & (!g48) & (!g69) & (g74) & (g84)) + ((shiftx4x) & (!shiftx5x) & (!g48) & (g69) & (g74) & (!g84)) + ((shiftx4x) & (!shiftx5x) & (!g48) & (g69) & (g74) & (g84)) + ((shiftx4x) & (!shiftx5x) & (g48) & (!g69) & (g74) & (!g84)) + ((shiftx4x) & (!shiftx5x) & (g48) & (!g69) & (g74) & (g84)) + ((shiftx4x) & (!shiftx5x) & (g48) & (g69) & (g74) & (!g84)) + ((shiftx4x) & (!shiftx5x) & (g48) & (g69) & (g74) & (g84)) + ((shiftx4x) & (shiftx5x) & (g48) & (!g69) & (!g74) & (!g84)) + ((shiftx4x) & (shiftx5x) & (g48) & (!g69) & (!g74) & (g84)) + ((shiftx4x) & (shiftx5x) & (g48) & (!g69) & (g74) & (!g84)) + ((shiftx4x) & (shiftx5x) & (g48) & (!g69) & (g74) & (g84)) + ((shiftx4x) & (shiftx5x) & (g48) & (g69) & (!g74) & (!g84)) + ((shiftx4x) & (shiftx5x) & (g48) & (g69) & (!g74) & (g84)) + ((shiftx4x) & (shiftx5x) & (g48) & (g69) & (g74) & (!g84)) + ((shiftx4x) & (shiftx5x) & (g48) & (g69) & (g74) & (g84)));
	assign g405 = (((!shiftx4x) & (!shiftx5x) & (!g53) & (g58) & (!g63) & (!g79)) + ((!shiftx4x) & (!shiftx5x) & (!g53) & (g58) & (!g63) & (g79)) + ((!shiftx4x) & (!shiftx5x) & (!g53) & (g58) & (g63) & (!g79)) + ((!shiftx4x) & (!shiftx5x) & (!g53) & (g58) & (g63) & (g79)) + ((!shiftx4x) & (!shiftx5x) & (g53) & (g58) & (!g63) & (!g79)) + ((!shiftx4x) & (!shiftx5x) & (g53) & (g58) & (!g63) & (g79)) + ((!shiftx4x) & (!shiftx5x) & (g53) & (g58) & (g63) & (!g79)) + ((!shiftx4x) & (!shiftx5x) & (g53) & (g58) & (g63) & (g79)) + ((!shiftx4x) & (shiftx5x) & (g53) & (!g58) & (!g63) & (!g79)) + ((!shiftx4x) & (shiftx5x) & (g53) & (!g58) & (!g63) & (g79)) + ((!shiftx4x) & (shiftx5x) & (g53) & (!g58) & (g63) & (!g79)) + ((!shiftx4x) & (shiftx5x) & (g53) & (!g58) & (g63) & (g79)) + ((!shiftx4x) & (shiftx5x) & (g53) & (g58) & (!g63) & (!g79)) + ((!shiftx4x) & (shiftx5x) & (g53) & (g58) & (!g63) & (g79)) + ((!shiftx4x) & (shiftx5x) & (g53) & (g58) & (g63) & (!g79)) + ((!shiftx4x) & (shiftx5x) & (g53) & (g58) & (g63) & (g79)) + ((shiftx4x) & (!shiftx5x) & (!g53) & (!g58) & (g63) & (!g79)) + ((shiftx4x) & (!shiftx5x) & (!g53) & (!g58) & (g63) & (g79)) + ((shiftx4x) & (!shiftx5x) & (!g53) & (g58) & (g63) & (!g79)) + ((shiftx4x) & (!shiftx5x) & (!g53) & (g58) & (g63) & (g79)) + ((shiftx4x) & (!shiftx5x) & (g53) & (!g58) & (g63) & (!g79)) + ((shiftx4x) & (!shiftx5x) & (g53) & (!g58) & (g63) & (g79)) + ((shiftx4x) & (!shiftx5x) & (g53) & (g58) & (g63) & (!g79)) + ((shiftx4x) & (!shiftx5x) & (g53) & (g58) & (g63) & (g79)) + ((shiftx4x) & (shiftx5x) & (!g53) & (!g58) & (!g63) & (g79)) + ((shiftx4x) & (shiftx5x) & (!g53) & (!g58) & (g63) & (g79)) + ((shiftx4x) & (shiftx5x) & (!g53) & (g58) & (!g63) & (g79)) + ((shiftx4x) & (shiftx5x) & (!g53) & (g58) & (g63) & (g79)) + ((shiftx4x) & (shiftx5x) & (g53) & (!g58) & (!g63) & (g79)) + ((shiftx4x) & (shiftx5x) & (g53) & (!g58) & (g63) & (g79)) + ((shiftx4x) & (shiftx5x) & (g53) & (g58) & (!g63) & (g79)) + ((shiftx4x) & (shiftx5x) & (g53) & (g58) & (g63) & (g79)));
	assign resultx49x = (((!sk[21]) & (shiftx6x) & (!g404) & (!g405)) + ((!sk[21]) & (shiftx6x) & (!g404) & (g405)) + ((!sk[21]) & (shiftx6x) & (g404) & (!g405)) + ((!sk[21]) & (shiftx6x) & (g404) & (g405)) + ((sk[21]) & (!shiftx6x) & (!g404) & (g405)) + ((sk[21]) & (!shiftx6x) & (g404) & (g405)) + ((sk[21]) & (shiftx6x) & (g404) & (!g405)) + ((sk[21]) & (shiftx6x) & (g404) & (g405)));
	assign g407 = (((!shiftx4x) & (!shiftx5x) & (!g91) & (!g112) & (!g117) & (g127)) + ((!shiftx4x) & (!shiftx5x) & (!g91) & (!g112) & (g117) & (g127)) + ((!shiftx4x) & (!shiftx5x) & (!g91) & (g112) & (!g117) & (g127)) + ((!shiftx4x) & (!shiftx5x) & (!g91) & (g112) & (g117) & (g127)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (!g112) & (!g117) & (g127)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (!g112) & (g117) & (g127)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (g112) & (!g117) & (g127)) + ((!shiftx4x) & (!shiftx5x) & (g91) & (g112) & (g117) & (g127)) + ((!shiftx4x) & (shiftx5x) & (!g91) & (g112) & (!g117) & (!g127)) + ((!shiftx4x) & (shiftx5x) & (!g91) & (g112) & (!g117) & (g127)) + ((!shiftx4x) & (shiftx5x) & (!g91) & (g112) & (g117) & (!g127)) + ((!shiftx4x) & (shiftx5x) & (!g91) & (g112) & (g117) & (g127)) + ((!shiftx4x) & (shiftx5x) & (g91) & (g112) & (!g117) & (!g127)) + ((!shiftx4x) & (shiftx5x) & (g91) & (g112) & (!g117) & (g127)) + ((!shiftx4x) & (shiftx5x) & (g91) & (g112) & (g117) & (!g127)) + ((!shiftx4x) & (shiftx5x) & (g91) & (g112) & (g117) & (g127)) + ((shiftx4x) & (!shiftx5x) & (!g91) & (!g112) & (g117) & (!g127)) + ((shiftx4x) & (!shiftx5x) & (!g91) & (!g112) & (g117) & (g127)) + ((shiftx4x) & (!shiftx5x) & (!g91) & (g112) & (g117) & (!g127)) + ((shiftx4x) & (!shiftx5x) & (!g91) & (g112) & (g117) & (g127)) + ((shiftx4x) & (!shiftx5x) & (g91) & (!g112) & (g117) & (!g127)) + ((shiftx4x) & (!shiftx5x) & (g91) & (!g112) & (g117) & (g127)) + ((shiftx4x) & (!shiftx5x) & (g91) & (g112) & (g117) & (!g127)) + ((shiftx4x) & (!shiftx5x) & (g91) & (g112) & (g117) & (g127)) + ((shiftx4x) & (shiftx5x) & (g91) & (!g112) & (!g117) & (!g127)) + ((shiftx4x) & (shiftx5x) & (g91) & (!g112) & (!g117) & (g127)) + ((shiftx4x) & (shiftx5x) & (g91) & (!g112) & (g117) & (!g127)) + ((shiftx4x) & (shiftx5x) & (g91) & (!g112) & (g117) & (g127)) + ((shiftx4x) & (shiftx5x) & (g91) & (g112) & (!g117) & (!g127)) + ((shiftx4x) & (shiftx5x) & (g91) & (g112) & (!g117) & (g127)) + ((shiftx4x) & (shiftx5x) & (g91) & (g112) & (g117) & (!g127)) + ((shiftx4x) & (shiftx5x) & (g91) & (g112) & (g117) & (g127)));
	assign g408 = (((!shiftx4x) & (!shiftx5x) & (!g96) & (g101) & (!g106) & (!g122)) + ((!shiftx4x) & (!shiftx5x) & (!g96) & (g101) & (!g106) & (g122)) + ((!shiftx4x) & (!shiftx5x) & (!g96) & (g101) & (g106) & (!g122)) + ((!shiftx4x) & (!shiftx5x) & (!g96) & (g101) & (g106) & (g122)) + ((!shiftx4x) & (!shiftx5x) & (g96) & (g101) & (!g106) & (!g122)) + ((!shiftx4x) & (!shiftx5x) & (g96) & (g101) & (!g106) & (g122)) + ((!shiftx4x) & (!shiftx5x) & (g96) & (g101) & (g106) & (!g122)) + ((!shiftx4x) & (!shiftx5x) & (g96) & (g101) & (g106) & (g122)) + ((!shiftx4x) & (shiftx5x) & (g96) & (!g101) & (!g106) & (!g122)) + ((!shiftx4x) & (shiftx5x) & (g96) & (!g101) & (!g106) & (g122)) + ((!shiftx4x) & (shiftx5x) & (g96) & (!g101) & (g106) & (!g122)) + ((!shiftx4x) & (shiftx5x) & (g96) & (!g101) & (g106) & (g122)) + ((!shiftx4x) & (shiftx5x) & (g96) & (g101) & (!g106) & (!g122)) + ((!shiftx4x) & (shiftx5x) & (g96) & (g101) & (!g106) & (g122)) + ((!shiftx4x) & (shiftx5x) & (g96) & (g101) & (g106) & (!g122)) + ((!shiftx4x) & (shiftx5x) & (g96) & (g101) & (g106) & (g122)) + ((shiftx4x) & (!shiftx5x) & (!g96) & (!g101) & (g106) & (!g122)) + ((shiftx4x) & (!shiftx5x) & (!g96) & (!g101) & (g106) & (g122)) + ((shiftx4x) & (!shiftx5x) & (!g96) & (g101) & (g106) & (!g122)) + ((shiftx4x) & (!shiftx5x) & (!g96) & (g101) & (g106) & (g122)) + ((shiftx4x) & (!shiftx5x) & (g96) & (!g101) & (g106) & (!g122)) + ((shiftx4x) & (!shiftx5x) & (g96) & (!g101) & (g106) & (g122)) + ((shiftx4x) & (!shiftx5x) & (g96) & (g101) & (g106) & (!g122)) + ((shiftx4x) & (!shiftx5x) & (g96) & (g101) & (g106) & (g122)) + ((shiftx4x) & (shiftx5x) & (!g96) & (!g101) & (!g106) & (g122)) + ((shiftx4x) & (shiftx5x) & (!g96) & (!g101) & (g106) & (g122)) + ((shiftx4x) & (shiftx5x) & (!g96) & (g101) & (!g106) & (g122)) + ((shiftx4x) & (shiftx5x) & (!g96) & (g101) & (g106) & (g122)) + ((shiftx4x) & (shiftx5x) & (g96) & (!g101) & (!g106) & (g122)) + ((shiftx4x) & (shiftx5x) & (g96) & (!g101) & (g106) & (g122)) + ((shiftx4x) & (shiftx5x) & (g96) & (g101) & (!g106) & (g122)) + ((shiftx4x) & (shiftx5x) & (g96) & (g101) & (g106) & (g122)));
	assign resultx50x = (((!shiftx6x) & (sk[24]) & (!g407) & (g408)) + ((!shiftx6x) & (sk[24]) & (g407) & (g408)) + ((shiftx6x) & (!sk[24]) & (!g407) & (!g408)) + ((shiftx6x) & (!sk[24]) & (!g407) & (g408)) + ((shiftx6x) & (!sk[24]) & (g407) & (!g408)) + ((shiftx6x) & (!sk[24]) & (g407) & (g408)) + ((shiftx6x) & (sk[24]) & (g407) & (!g408)) + ((shiftx6x) & (sk[24]) & (g407) & (g408)));
	assign g410 = (((!shiftx4x) & (!shiftx5x) & (!g134) & (g155) & (!g160) & (!g170)) + ((!shiftx4x) & (!shiftx5x) & (!g134) & (g155) & (!g160) & (g170)) + ((!shiftx4x) & (!shiftx5x) & (!g134) & (g155) & (g160) & (!g170)) + ((!shiftx4x) & (!shiftx5x) & (!g134) & (g155) & (g160) & (g170)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (g155) & (!g160) & (!g170)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (g155) & (!g160) & (g170)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (g155) & (g160) & (!g170)) + ((!shiftx4x) & (!shiftx5x) & (g134) & (g155) & (g160) & (g170)) + ((!shiftx4x) & (shiftx5x) & (!g134) & (!g155) & (!g160) & (g170)) + ((!shiftx4x) & (shiftx5x) & (!g134) & (!g155) & (g160) & (g170)) + ((!shiftx4x) & (shiftx5x) & (!g134) & (g155) & (!g160) & (g170)) + ((!shiftx4x) & (shiftx5x) & (!g134) & (g155) & (g160) & (g170)) + ((!shiftx4x) & (shiftx5x) & (g134) & (!g155) & (!g160) & (g170)) + ((!shiftx4x) & (shiftx5x) & (g134) & (!g155) & (g160) & (g170)) + ((!shiftx4x) & (shiftx5x) & (g134) & (g155) & (!g160) & (g170)) + ((!shiftx4x) & (shiftx5x) & (g134) & (g155) & (g160) & (g170)) + ((shiftx4x) & (!shiftx5x) & (!g134) & (!g155) & (g160) & (!g170)) + ((shiftx4x) & (!shiftx5x) & (!g134) & (!g155) & (g160) & (g170)) + ((shiftx4x) & (!shiftx5x) & (!g134) & (g155) & (g160) & (!g170)) + ((shiftx4x) & (!shiftx5x) & (!g134) & (g155) & (g160) & (g170)) + ((shiftx4x) & (!shiftx5x) & (g134) & (!g155) & (g160) & (!g170)) + ((shiftx4x) & (!shiftx5x) & (g134) & (!g155) & (g160) & (g170)) + ((shiftx4x) & (!shiftx5x) & (g134) & (g155) & (g160) & (!g170)) + ((shiftx4x) & (!shiftx5x) & (g134) & (g155) & (g160) & (g170)) + ((shiftx4x) & (shiftx5x) & (g134) & (!g155) & (!g160) & (!g170)) + ((shiftx4x) & (shiftx5x) & (g134) & (!g155) & (!g160) & (g170)) + ((shiftx4x) & (shiftx5x) & (g134) & (!g155) & (g160) & (!g170)) + ((shiftx4x) & (shiftx5x) & (g134) & (!g155) & (g160) & (g170)) + ((shiftx4x) & (shiftx5x) & (g134) & (g155) & (!g160) & (!g170)) + ((shiftx4x) & (shiftx5x) & (g134) & (g155) & (!g160) & (g170)) + ((shiftx4x) & (shiftx5x) & (g134) & (g155) & (g160) & (!g170)) + ((shiftx4x) & (shiftx5x) & (g134) & (g155) & (g160) & (g170)));
	assign g411 = (((!shiftx4x) & (!shiftx5x) & (g139) & (!g144) & (!g149) & (!g165)) + ((!shiftx4x) & (!shiftx5x) & (g139) & (!g144) & (!g149) & (g165)) + ((!shiftx4x) & (!shiftx5x) & (g139) & (!g144) & (g149) & (!g165)) + ((!shiftx4x) & (!shiftx5x) & (g139) & (!g144) & (g149) & (g165)) + ((!shiftx4x) & (!shiftx5x) & (g139) & (g144) & (!g149) & (!g165)) + ((!shiftx4x) & (!shiftx5x) & (g139) & (g144) & (!g149) & (g165)) + ((!shiftx4x) & (!shiftx5x) & (g139) & (g144) & (g149) & (!g165)) + ((!shiftx4x) & (!shiftx5x) & (g139) & (g144) & (g149) & (g165)) + ((!shiftx4x) & (shiftx5x) & (!g139) & (g144) & (!g149) & (!g165)) + ((!shiftx4x) & (shiftx5x) & (!g139) & (g144) & (!g149) & (g165)) + ((!shiftx4x) & (shiftx5x) & (!g139) & (g144) & (g149) & (!g165)) + ((!shiftx4x) & (shiftx5x) & (!g139) & (g144) & (g149) & (g165)) + ((!shiftx4x) & (shiftx5x) & (g139) & (g144) & (!g149) & (!g165)) + ((!shiftx4x) & (shiftx5x) & (g139) & (g144) & (!g149) & (g165)) + ((!shiftx4x) & (shiftx5x) & (g139) & (g144) & (g149) & (!g165)) + ((!shiftx4x) & (shiftx5x) & (g139) & (g144) & (g149) & (g165)) + ((shiftx4x) & (!shiftx5x) & (!g139) & (!g144) & (g149) & (!g165)) + ((shiftx4x) & (!shiftx5x) & (!g139) & (!g144) & (g149) & (g165)) + ((shiftx4x) & (!shiftx5x) & (!g139) & (g144) & (g149) & (!g165)) + ((shiftx4x) & (!shiftx5x) & (!g139) & (g144) & (g149) & (g165)) + ((shiftx4x) & (!shiftx5x) & (g139) & (!g144) & (g149) & (!g165)) + ((shiftx4x) & (!shiftx5x) & (g139) & (!g144) & (g149) & (g165)) + ((shiftx4x) & (!shiftx5x) & (g139) & (g144) & (g149) & (!g165)) + ((shiftx4x) & (!shiftx5x) & (g139) & (g144) & (g149) & (g165)) + ((shiftx4x) & (shiftx5x) & (!g139) & (!g144) & (!g149) & (g165)) + ((shiftx4x) & (shiftx5x) & (!g139) & (!g144) & (g149) & (g165)) + ((shiftx4x) & (shiftx5x) & (!g139) & (g144) & (!g149) & (g165)) + ((shiftx4x) & (shiftx5x) & (!g139) & (g144) & (g149) & (g165)) + ((shiftx4x) & (shiftx5x) & (g139) & (!g144) & (!g149) & (g165)) + ((shiftx4x) & (shiftx5x) & (g139) & (!g144) & (g149) & (g165)) + ((shiftx4x) & (shiftx5x) & (g139) & (g144) & (!g149) & (g165)) + ((shiftx4x) & (shiftx5x) & (g139) & (g144) & (g149) & (g165)));
	assign resultx51x = (((!shiftx6x) & (!g410) & (sk[27]) & (g411)) + ((!shiftx6x) & (g410) & (sk[27]) & (g411)) + ((shiftx6x) & (!g410) & (!sk[27]) & (!g411)) + ((shiftx6x) & (!g410) & (!sk[27]) & (g411)) + ((shiftx6x) & (g410) & (!sk[27]) & (!g411)) + ((shiftx6x) & (g410) & (!sk[27]) & (g411)) + ((shiftx6x) & (g410) & (sk[27]) & (!g411)) + ((shiftx6x) & (g410) & (sk[27]) & (g411)));
	assign g413 = (((!shiftx4x) & (!shiftx5x) & (!g174) & (!g178) & (!g179) & (g181)) + ((!shiftx4x) & (!shiftx5x) & (!g174) & (!g178) & (g179) & (g181)) + ((!shiftx4x) & (!shiftx5x) & (!g174) & (g178) & (!g179) & (g181)) + ((!shiftx4x) & (!shiftx5x) & (!g174) & (g178) & (g179) & (g181)) + ((!shiftx4x) & (!shiftx5x) & (g174) & (!g178) & (!g179) & (g181)) + ((!shiftx4x) & (!shiftx5x) & (g174) & (!g178) & (g179) & (g181)) + ((!shiftx4x) & (!shiftx5x) & (g174) & (g178) & (!g179) & (g181)) + ((!shiftx4x) & (!shiftx5x) & (g174) & (g178) & (g179) & (g181)) + ((!shiftx4x) & (shiftx5x) & (!g174) & (g178) & (!g179) & (!g181)) + ((!shiftx4x) & (shiftx5x) & (!g174) & (g178) & (!g179) & (g181)) + ((!shiftx4x) & (shiftx5x) & (!g174) & (g178) & (g179) & (!g181)) + ((!shiftx4x) & (shiftx5x) & (!g174) & (g178) & (g179) & (g181)) + ((!shiftx4x) & (shiftx5x) & (g174) & (g178) & (!g179) & (!g181)) + ((!shiftx4x) & (shiftx5x) & (g174) & (g178) & (!g179) & (g181)) + ((!shiftx4x) & (shiftx5x) & (g174) & (g178) & (g179) & (!g181)) + ((!shiftx4x) & (shiftx5x) & (g174) & (g178) & (g179) & (g181)) + ((shiftx4x) & (!shiftx5x) & (!g174) & (!g178) & (g179) & (!g181)) + ((shiftx4x) & (!shiftx5x) & (!g174) & (!g178) & (g179) & (g181)) + ((shiftx4x) & (!shiftx5x) & (!g174) & (g178) & (g179) & (!g181)) + ((shiftx4x) & (!shiftx5x) & (!g174) & (g178) & (g179) & (g181)) + ((shiftx4x) & (!shiftx5x) & (g174) & (!g178) & (g179) & (!g181)) + ((shiftx4x) & (!shiftx5x) & (g174) & (!g178) & (g179) & (g181)) + ((shiftx4x) & (!shiftx5x) & (g174) & (g178) & (g179) & (!g181)) + ((shiftx4x) & (!shiftx5x) & (g174) & (g178) & (g179) & (g181)) + ((shiftx4x) & (shiftx5x) & (g174) & (!g178) & (!g179) & (!g181)) + ((shiftx4x) & (shiftx5x) & (g174) & (!g178) & (!g179) & (g181)) + ((shiftx4x) & (shiftx5x) & (g174) & (!g178) & (g179) & (!g181)) + ((shiftx4x) & (shiftx5x) & (g174) & (!g178) & (g179) & (g181)) + ((shiftx4x) & (shiftx5x) & (g174) & (g178) & (!g179) & (!g181)) + ((shiftx4x) & (shiftx5x) & (g174) & (g178) & (!g179) & (g181)) + ((shiftx4x) & (shiftx5x) & (g174) & (g178) & (g179) & (!g181)) + ((shiftx4x) & (shiftx5x) & (g174) & (g178) & (g179) & (g181)));
	assign g414 = (((!shiftx4x) & (!shiftx5x) & (g173) & (!g175) & (!g176) & (!g180)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (!g175) & (!g176) & (g180)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (!g175) & (g176) & (!g180)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (!g175) & (g176) & (g180)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (g175) & (!g176) & (!g180)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (g175) & (!g176) & (g180)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (g175) & (g176) & (!g180)) + ((!shiftx4x) & (!shiftx5x) & (g173) & (g175) & (g176) & (g180)) + ((!shiftx4x) & (shiftx5x) & (!g173) & (!g175) & (g176) & (!g180)) + ((!shiftx4x) & (shiftx5x) & (!g173) & (!g175) & (g176) & (g180)) + ((!shiftx4x) & (shiftx5x) & (!g173) & (g175) & (g176) & (!g180)) + ((!shiftx4x) & (shiftx5x) & (!g173) & (g175) & (g176) & (g180)) + ((!shiftx4x) & (shiftx5x) & (g173) & (!g175) & (g176) & (!g180)) + ((!shiftx4x) & (shiftx5x) & (g173) & (!g175) & (g176) & (g180)) + ((!shiftx4x) & (shiftx5x) & (g173) & (g175) & (g176) & (!g180)) + ((!shiftx4x) & (shiftx5x) & (g173) & (g175) & (g176) & (g180)) + ((shiftx4x) & (!shiftx5x) & (!g173) & (g175) & (!g176) & (!g180)) + ((shiftx4x) & (!shiftx5x) & (!g173) & (g175) & (!g176) & (g180)) + ((shiftx4x) & (!shiftx5x) & (!g173) & (g175) & (g176) & (!g180)) + ((shiftx4x) & (!shiftx5x) & (!g173) & (g175) & (g176) & (g180)) + ((shiftx4x) & (!shiftx5x) & (g173) & (g175) & (!g176) & (!g180)) + ((shiftx4x) & (!shiftx5x) & (g173) & (g175) & (!g176) & (g180)) + ((shiftx4x) & (!shiftx5x) & (g173) & (g175) & (g176) & (!g180)) + ((shiftx4x) & (!shiftx5x) & (g173) & (g175) & (g176) & (g180)) + ((shiftx4x) & (shiftx5x) & (!g173) & (!g175) & (!g176) & (g180)) + ((shiftx4x) & (shiftx5x) & (!g173) & (!g175) & (g176) & (g180)) + ((shiftx4x) & (shiftx5x) & (!g173) & (g175) & (!g176) & (g180)) + ((shiftx4x) & (shiftx5x) & (!g173) & (g175) & (g176) & (g180)) + ((shiftx4x) & (shiftx5x) & (g173) & (!g175) & (!g176) & (g180)) + ((shiftx4x) & (shiftx5x) & (g173) & (!g175) & (g176) & (g180)) + ((shiftx4x) & (shiftx5x) & (g173) & (g175) & (!g176) & (g180)) + ((shiftx4x) & (shiftx5x) & (g173) & (g175) & (g176) & (g180)));
	assign resultx52x = (((!shiftx6x) & (!g413) & (sk[30]) & (g414)) + ((!shiftx6x) & (g413) & (sk[30]) & (g414)) + ((shiftx6x) & (!g413) & (!sk[30]) & (!g414)) + ((shiftx6x) & (!g413) & (!sk[30]) & (g414)) + ((shiftx6x) & (g413) & (!sk[30]) & (!g414)) + ((shiftx6x) & (g413) & (!sk[30]) & (g414)) + ((shiftx6x) & (g413) & (sk[30]) & (!g414)) + ((shiftx6x) & (g413) & (sk[30]) & (g414)));
	assign g416 = (((!shiftx4x) & (!shiftx5x) & (!g185) & (!g189) & (!g190) & (g192)) + ((!shiftx4x) & (!shiftx5x) & (!g185) & (!g189) & (g190) & (g192)) + ((!shiftx4x) & (!shiftx5x) & (!g185) & (g189) & (!g190) & (g192)) + ((!shiftx4x) & (!shiftx5x) & (!g185) & (g189) & (g190) & (g192)) + ((!shiftx4x) & (!shiftx5x) & (g185) & (!g189) & (!g190) & (g192)) + ((!shiftx4x) & (!shiftx5x) & (g185) & (!g189) & (g190) & (g192)) + ((!shiftx4x) & (!shiftx5x) & (g185) & (g189) & (!g190) & (g192)) + ((!shiftx4x) & (!shiftx5x) & (g185) & (g189) & (g190) & (g192)) + ((!shiftx4x) & (shiftx5x) & (!g185) & (g189) & (!g190) & (!g192)) + ((!shiftx4x) & (shiftx5x) & (!g185) & (g189) & (!g190) & (g192)) + ((!shiftx4x) & (shiftx5x) & (!g185) & (g189) & (g190) & (!g192)) + ((!shiftx4x) & (shiftx5x) & (!g185) & (g189) & (g190) & (g192)) + ((!shiftx4x) & (shiftx5x) & (g185) & (g189) & (!g190) & (!g192)) + ((!shiftx4x) & (shiftx5x) & (g185) & (g189) & (!g190) & (g192)) + ((!shiftx4x) & (shiftx5x) & (g185) & (g189) & (g190) & (!g192)) + ((!shiftx4x) & (shiftx5x) & (g185) & (g189) & (g190) & (g192)) + ((shiftx4x) & (!shiftx5x) & (!g185) & (!g189) & (g190) & (!g192)) + ((shiftx4x) & (!shiftx5x) & (!g185) & (!g189) & (g190) & (g192)) + ((shiftx4x) & (!shiftx5x) & (!g185) & (g189) & (g190) & (!g192)) + ((shiftx4x) & (!shiftx5x) & (!g185) & (g189) & (g190) & (g192)) + ((shiftx4x) & (!shiftx5x) & (g185) & (!g189) & (g190) & (!g192)) + ((shiftx4x) & (!shiftx5x) & (g185) & (!g189) & (g190) & (g192)) + ((shiftx4x) & (!shiftx5x) & (g185) & (g189) & (g190) & (!g192)) + ((shiftx4x) & (!shiftx5x) & (g185) & (g189) & (g190) & (g192)) + ((shiftx4x) & (shiftx5x) & (g185) & (!g189) & (!g190) & (!g192)) + ((shiftx4x) & (shiftx5x) & (g185) & (!g189) & (!g190) & (g192)) + ((shiftx4x) & (shiftx5x) & (g185) & (!g189) & (g190) & (!g192)) + ((shiftx4x) & (shiftx5x) & (g185) & (!g189) & (g190) & (g192)) + ((shiftx4x) & (shiftx5x) & (g185) & (g189) & (!g190) & (!g192)) + ((shiftx4x) & (shiftx5x) & (g185) & (g189) & (!g190) & (g192)) + ((shiftx4x) & (shiftx5x) & (g185) & (g189) & (g190) & (!g192)) + ((shiftx4x) & (shiftx5x) & (g185) & (g189) & (g190) & (g192)));
	assign g417 = (((!shiftx4x) & (!shiftx5x) & (g184) & (!g186) & (!g187) & (!g191)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (!g186) & (!g187) & (g191)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (!g186) & (g187) & (!g191)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (!g186) & (g187) & (g191)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (g186) & (!g187) & (!g191)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (g186) & (!g187) & (g191)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (g186) & (g187) & (!g191)) + ((!shiftx4x) & (!shiftx5x) & (g184) & (g186) & (g187) & (g191)) + ((!shiftx4x) & (shiftx5x) & (!g184) & (!g186) & (g187) & (!g191)) + ((!shiftx4x) & (shiftx5x) & (!g184) & (!g186) & (g187) & (g191)) + ((!shiftx4x) & (shiftx5x) & (!g184) & (g186) & (g187) & (!g191)) + ((!shiftx4x) & (shiftx5x) & (!g184) & (g186) & (g187) & (g191)) + ((!shiftx4x) & (shiftx5x) & (g184) & (!g186) & (g187) & (!g191)) + ((!shiftx4x) & (shiftx5x) & (g184) & (!g186) & (g187) & (g191)) + ((!shiftx4x) & (shiftx5x) & (g184) & (g186) & (g187) & (!g191)) + ((!shiftx4x) & (shiftx5x) & (g184) & (g186) & (g187) & (g191)) + ((shiftx4x) & (!shiftx5x) & (!g184) & (g186) & (!g187) & (!g191)) + ((shiftx4x) & (!shiftx5x) & (!g184) & (g186) & (!g187) & (g191)) + ((shiftx4x) & (!shiftx5x) & (!g184) & (g186) & (g187) & (!g191)) + ((shiftx4x) & (!shiftx5x) & (!g184) & (g186) & (g187) & (g191)) + ((shiftx4x) & (!shiftx5x) & (g184) & (g186) & (!g187) & (!g191)) + ((shiftx4x) & (!shiftx5x) & (g184) & (g186) & (!g187) & (g191)) + ((shiftx4x) & (!shiftx5x) & (g184) & (g186) & (g187) & (!g191)) + ((shiftx4x) & (!shiftx5x) & (g184) & (g186) & (g187) & (g191)) + ((shiftx4x) & (shiftx5x) & (!g184) & (!g186) & (!g187) & (g191)) + ((shiftx4x) & (shiftx5x) & (!g184) & (!g186) & (g187) & (g191)) + ((shiftx4x) & (shiftx5x) & (!g184) & (g186) & (!g187) & (g191)) + ((shiftx4x) & (shiftx5x) & (!g184) & (g186) & (g187) & (g191)) + ((shiftx4x) & (shiftx5x) & (g184) & (!g186) & (!g187) & (g191)) + ((shiftx4x) & (shiftx5x) & (g184) & (!g186) & (g187) & (g191)) + ((shiftx4x) & (shiftx5x) & (g184) & (g186) & (!g187) & (g191)) + ((shiftx4x) & (shiftx5x) & (g184) & (g186) & (g187) & (g191)));
	assign resultx53x = (((!sk[33]) & (shiftx6x) & (!g416) & (!g417)) + ((!sk[33]) & (shiftx6x) & (!g416) & (g417)) + ((!sk[33]) & (shiftx6x) & (g416) & (!g417)) + ((!sk[33]) & (shiftx6x) & (g416) & (g417)) + ((sk[33]) & (!shiftx6x) & (!g416) & (g417)) + ((sk[33]) & (!shiftx6x) & (g416) & (g417)) + ((sk[33]) & (shiftx6x) & (g416) & (!g417)) + ((sk[33]) & (shiftx6x) & (g416) & (g417)));
	assign g419 = (((!shiftx4x) & (!shiftx5x) & (!g196) & (!g200) & (!g201) & (g203)) + ((!shiftx4x) & (!shiftx5x) & (!g196) & (!g200) & (g201) & (g203)) + ((!shiftx4x) & (!shiftx5x) & (!g196) & (g200) & (!g201) & (g203)) + ((!shiftx4x) & (!shiftx5x) & (!g196) & (g200) & (g201) & (g203)) + ((!shiftx4x) & (!shiftx5x) & (g196) & (!g200) & (!g201) & (g203)) + ((!shiftx4x) & (!shiftx5x) & (g196) & (!g200) & (g201) & (g203)) + ((!shiftx4x) & (!shiftx5x) & (g196) & (g200) & (!g201) & (g203)) + ((!shiftx4x) & (!shiftx5x) & (g196) & (g200) & (g201) & (g203)) + ((!shiftx4x) & (shiftx5x) & (!g196) & (g200) & (!g201) & (!g203)) + ((!shiftx4x) & (shiftx5x) & (!g196) & (g200) & (!g201) & (g203)) + ((!shiftx4x) & (shiftx5x) & (!g196) & (g200) & (g201) & (!g203)) + ((!shiftx4x) & (shiftx5x) & (!g196) & (g200) & (g201) & (g203)) + ((!shiftx4x) & (shiftx5x) & (g196) & (g200) & (!g201) & (!g203)) + ((!shiftx4x) & (shiftx5x) & (g196) & (g200) & (!g201) & (g203)) + ((!shiftx4x) & (shiftx5x) & (g196) & (g200) & (g201) & (!g203)) + ((!shiftx4x) & (shiftx5x) & (g196) & (g200) & (g201) & (g203)) + ((shiftx4x) & (!shiftx5x) & (!g196) & (!g200) & (g201) & (!g203)) + ((shiftx4x) & (!shiftx5x) & (!g196) & (!g200) & (g201) & (g203)) + ((shiftx4x) & (!shiftx5x) & (!g196) & (g200) & (g201) & (!g203)) + ((shiftx4x) & (!shiftx5x) & (!g196) & (g200) & (g201) & (g203)) + ((shiftx4x) & (!shiftx5x) & (g196) & (!g200) & (g201) & (!g203)) + ((shiftx4x) & (!shiftx5x) & (g196) & (!g200) & (g201) & (g203)) + ((shiftx4x) & (!shiftx5x) & (g196) & (g200) & (g201) & (!g203)) + ((shiftx4x) & (!shiftx5x) & (g196) & (g200) & (g201) & (g203)) + ((shiftx4x) & (shiftx5x) & (g196) & (!g200) & (!g201) & (!g203)) + ((shiftx4x) & (shiftx5x) & (g196) & (!g200) & (!g201) & (g203)) + ((shiftx4x) & (shiftx5x) & (g196) & (!g200) & (g201) & (!g203)) + ((shiftx4x) & (shiftx5x) & (g196) & (!g200) & (g201) & (g203)) + ((shiftx4x) & (shiftx5x) & (g196) & (g200) & (!g201) & (!g203)) + ((shiftx4x) & (shiftx5x) & (g196) & (g200) & (!g201) & (g203)) + ((shiftx4x) & (shiftx5x) & (g196) & (g200) & (g201) & (!g203)) + ((shiftx4x) & (shiftx5x) & (g196) & (g200) & (g201) & (g203)));
	assign g420 = (((!shiftx4x) & (!shiftx5x) & (g195) & (!g197) & (!g198) & (!g202)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (!g197) & (!g198) & (g202)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (!g197) & (g198) & (!g202)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (!g197) & (g198) & (g202)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (g197) & (!g198) & (!g202)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (g197) & (!g198) & (g202)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (g197) & (g198) & (!g202)) + ((!shiftx4x) & (!shiftx5x) & (g195) & (g197) & (g198) & (g202)) + ((!shiftx4x) & (shiftx5x) & (!g195) & (!g197) & (g198) & (!g202)) + ((!shiftx4x) & (shiftx5x) & (!g195) & (!g197) & (g198) & (g202)) + ((!shiftx4x) & (shiftx5x) & (!g195) & (g197) & (g198) & (!g202)) + ((!shiftx4x) & (shiftx5x) & (!g195) & (g197) & (g198) & (g202)) + ((!shiftx4x) & (shiftx5x) & (g195) & (!g197) & (g198) & (!g202)) + ((!shiftx4x) & (shiftx5x) & (g195) & (!g197) & (g198) & (g202)) + ((!shiftx4x) & (shiftx5x) & (g195) & (g197) & (g198) & (!g202)) + ((!shiftx4x) & (shiftx5x) & (g195) & (g197) & (g198) & (g202)) + ((shiftx4x) & (!shiftx5x) & (!g195) & (g197) & (!g198) & (!g202)) + ((shiftx4x) & (!shiftx5x) & (!g195) & (g197) & (!g198) & (g202)) + ((shiftx4x) & (!shiftx5x) & (!g195) & (g197) & (g198) & (!g202)) + ((shiftx4x) & (!shiftx5x) & (!g195) & (g197) & (g198) & (g202)) + ((shiftx4x) & (!shiftx5x) & (g195) & (g197) & (!g198) & (!g202)) + ((shiftx4x) & (!shiftx5x) & (g195) & (g197) & (!g198) & (g202)) + ((shiftx4x) & (!shiftx5x) & (g195) & (g197) & (g198) & (!g202)) + ((shiftx4x) & (!shiftx5x) & (g195) & (g197) & (g198) & (g202)) + ((shiftx4x) & (shiftx5x) & (!g195) & (!g197) & (!g198) & (g202)) + ((shiftx4x) & (shiftx5x) & (!g195) & (!g197) & (g198) & (g202)) + ((shiftx4x) & (shiftx5x) & (!g195) & (g197) & (!g198) & (g202)) + ((shiftx4x) & (shiftx5x) & (!g195) & (g197) & (g198) & (g202)) + ((shiftx4x) & (shiftx5x) & (g195) & (!g197) & (!g198) & (g202)) + ((shiftx4x) & (shiftx5x) & (g195) & (!g197) & (g198) & (g202)) + ((shiftx4x) & (shiftx5x) & (g195) & (g197) & (!g198) & (g202)) + ((shiftx4x) & (shiftx5x) & (g195) & (g197) & (g198) & (g202)));
	assign resultx54x = (((!shiftx6x) & (!g419) & (sk[36]) & (g420)) + ((!shiftx6x) & (g419) & (sk[36]) & (g420)) + ((shiftx6x) & (!g419) & (!sk[36]) & (!g420)) + ((shiftx6x) & (!g419) & (!sk[36]) & (g420)) + ((shiftx6x) & (g419) & (!sk[36]) & (!g420)) + ((shiftx6x) & (g419) & (!sk[36]) & (g420)) + ((shiftx6x) & (g419) & (sk[36]) & (!g420)) + ((shiftx6x) & (g419) & (sk[36]) & (g420)));
	assign g422 = (((!shiftx4x) & (!shiftx5x) & (!g207) & (!g211) & (!g212) & (g214)) + ((!shiftx4x) & (!shiftx5x) & (!g207) & (!g211) & (g212) & (g214)) + ((!shiftx4x) & (!shiftx5x) & (!g207) & (g211) & (!g212) & (g214)) + ((!shiftx4x) & (!shiftx5x) & (!g207) & (g211) & (g212) & (g214)) + ((!shiftx4x) & (!shiftx5x) & (g207) & (!g211) & (!g212) & (g214)) + ((!shiftx4x) & (!shiftx5x) & (g207) & (!g211) & (g212) & (g214)) + ((!shiftx4x) & (!shiftx5x) & (g207) & (g211) & (!g212) & (g214)) + ((!shiftx4x) & (!shiftx5x) & (g207) & (g211) & (g212) & (g214)) + ((!shiftx4x) & (shiftx5x) & (!g207) & (g211) & (!g212) & (!g214)) + ((!shiftx4x) & (shiftx5x) & (!g207) & (g211) & (!g212) & (g214)) + ((!shiftx4x) & (shiftx5x) & (!g207) & (g211) & (g212) & (!g214)) + ((!shiftx4x) & (shiftx5x) & (!g207) & (g211) & (g212) & (g214)) + ((!shiftx4x) & (shiftx5x) & (g207) & (g211) & (!g212) & (!g214)) + ((!shiftx4x) & (shiftx5x) & (g207) & (g211) & (!g212) & (g214)) + ((!shiftx4x) & (shiftx5x) & (g207) & (g211) & (g212) & (!g214)) + ((!shiftx4x) & (shiftx5x) & (g207) & (g211) & (g212) & (g214)) + ((shiftx4x) & (!shiftx5x) & (!g207) & (!g211) & (g212) & (!g214)) + ((shiftx4x) & (!shiftx5x) & (!g207) & (!g211) & (g212) & (g214)) + ((shiftx4x) & (!shiftx5x) & (!g207) & (g211) & (g212) & (!g214)) + ((shiftx4x) & (!shiftx5x) & (!g207) & (g211) & (g212) & (g214)) + ((shiftx4x) & (!shiftx5x) & (g207) & (!g211) & (g212) & (!g214)) + ((shiftx4x) & (!shiftx5x) & (g207) & (!g211) & (g212) & (g214)) + ((shiftx4x) & (!shiftx5x) & (g207) & (g211) & (g212) & (!g214)) + ((shiftx4x) & (!shiftx5x) & (g207) & (g211) & (g212) & (g214)) + ((shiftx4x) & (shiftx5x) & (g207) & (!g211) & (!g212) & (!g214)) + ((shiftx4x) & (shiftx5x) & (g207) & (!g211) & (!g212) & (g214)) + ((shiftx4x) & (shiftx5x) & (g207) & (!g211) & (g212) & (!g214)) + ((shiftx4x) & (shiftx5x) & (g207) & (!g211) & (g212) & (g214)) + ((shiftx4x) & (shiftx5x) & (g207) & (g211) & (!g212) & (!g214)) + ((shiftx4x) & (shiftx5x) & (g207) & (g211) & (!g212) & (g214)) + ((shiftx4x) & (shiftx5x) & (g207) & (g211) & (g212) & (!g214)) + ((shiftx4x) & (shiftx5x) & (g207) & (g211) & (g212) & (g214)));
	assign g423 = (((!shiftx4x) & (!shiftx5x) & (g206) & (!g208) & (!g209) & (!g213)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (!g208) & (!g209) & (g213)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (!g208) & (g209) & (!g213)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (!g208) & (g209) & (g213)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (g208) & (!g209) & (!g213)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (g208) & (!g209) & (g213)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (g208) & (g209) & (!g213)) + ((!shiftx4x) & (!shiftx5x) & (g206) & (g208) & (g209) & (g213)) + ((!shiftx4x) & (shiftx5x) & (!g206) & (!g208) & (g209) & (!g213)) + ((!shiftx4x) & (shiftx5x) & (!g206) & (!g208) & (g209) & (g213)) + ((!shiftx4x) & (shiftx5x) & (!g206) & (g208) & (g209) & (!g213)) + ((!shiftx4x) & (shiftx5x) & (!g206) & (g208) & (g209) & (g213)) + ((!shiftx4x) & (shiftx5x) & (g206) & (!g208) & (g209) & (!g213)) + ((!shiftx4x) & (shiftx5x) & (g206) & (!g208) & (g209) & (g213)) + ((!shiftx4x) & (shiftx5x) & (g206) & (g208) & (g209) & (!g213)) + ((!shiftx4x) & (shiftx5x) & (g206) & (g208) & (g209) & (g213)) + ((shiftx4x) & (!shiftx5x) & (!g206) & (g208) & (!g209) & (!g213)) + ((shiftx4x) & (!shiftx5x) & (!g206) & (g208) & (!g209) & (g213)) + ((shiftx4x) & (!shiftx5x) & (!g206) & (g208) & (g209) & (!g213)) + ((shiftx4x) & (!shiftx5x) & (!g206) & (g208) & (g209) & (g213)) + ((shiftx4x) & (!shiftx5x) & (g206) & (g208) & (!g209) & (!g213)) + ((shiftx4x) & (!shiftx5x) & (g206) & (g208) & (!g209) & (g213)) + ((shiftx4x) & (!shiftx5x) & (g206) & (g208) & (g209) & (!g213)) + ((shiftx4x) & (!shiftx5x) & (g206) & (g208) & (g209) & (g213)) + ((shiftx4x) & (shiftx5x) & (!g206) & (!g208) & (!g209) & (g213)) + ((shiftx4x) & (shiftx5x) & (!g206) & (!g208) & (g209) & (g213)) + ((shiftx4x) & (shiftx5x) & (!g206) & (g208) & (!g209) & (g213)) + ((shiftx4x) & (shiftx5x) & (!g206) & (g208) & (g209) & (g213)) + ((shiftx4x) & (shiftx5x) & (g206) & (!g208) & (!g209) & (g213)) + ((shiftx4x) & (shiftx5x) & (g206) & (!g208) & (g209) & (g213)) + ((shiftx4x) & (shiftx5x) & (g206) & (g208) & (!g209) & (g213)) + ((shiftx4x) & (shiftx5x) & (g206) & (g208) & (g209) & (g213)));
	assign resultx55x = (((!sk[39]) & (shiftx6x) & (!g422) & (!g423)) + ((!sk[39]) & (shiftx6x) & (!g422) & (g423)) + ((!sk[39]) & (shiftx6x) & (g422) & (!g423)) + ((!sk[39]) & (shiftx6x) & (g422) & (g423)) + ((sk[39]) & (!shiftx6x) & (!g422) & (g423)) + ((sk[39]) & (!shiftx6x) & (g422) & (g423)) + ((sk[39]) & (shiftx6x) & (g422) & (!g423)) + ((sk[39]) & (shiftx6x) & (g422) & (g423)));
	assign g425 = (((!shiftx4x) & (!shiftx5x) & (!g218) & (!g222) & (!g223) & (g225)) + ((!shiftx4x) & (!shiftx5x) & (!g218) & (!g222) & (g223) & (g225)) + ((!shiftx4x) & (!shiftx5x) & (!g218) & (g222) & (!g223) & (g225)) + ((!shiftx4x) & (!shiftx5x) & (!g218) & (g222) & (g223) & (g225)) + ((!shiftx4x) & (!shiftx5x) & (g218) & (!g222) & (!g223) & (g225)) + ((!shiftx4x) & (!shiftx5x) & (g218) & (!g222) & (g223) & (g225)) + ((!shiftx4x) & (!shiftx5x) & (g218) & (g222) & (!g223) & (g225)) + ((!shiftx4x) & (!shiftx5x) & (g218) & (g222) & (g223) & (g225)) + ((!shiftx4x) & (shiftx5x) & (!g218) & (g222) & (!g223) & (!g225)) + ((!shiftx4x) & (shiftx5x) & (!g218) & (g222) & (!g223) & (g225)) + ((!shiftx4x) & (shiftx5x) & (!g218) & (g222) & (g223) & (!g225)) + ((!shiftx4x) & (shiftx5x) & (!g218) & (g222) & (g223) & (g225)) + ((!shiftx4x) & (shiftx5x) & (g218) & (g222) & (!g223) & (!g225)) + ((!shiftx4x) & (shiftx5x) & (g218) & (g222) & (!g223) & (g225)) + ((!shiftx4x) & (shiftx5x) & (g218) & (g222) & (g223) & (!g225)) + ((!shiftx4x) & (shiftx5x) & (g218) & (g222) & (g223) & (g225)) + ((shiftx4x) & (!shiftx5x) & (!g218) & (!g222) & (g223) & (!g225)) + ((shiftx4x) & (!shiftx5x) & (!g218) & (!g222) & (g223) & (g225)) + ((shiftx4x) & (!shiftx5x) & (!g218) & (g222) & (g223) & (!g225)) + ((shiftx4x) & (!shiftx5x) & (!g218) & (g222) & (g223) & (g225)) + ((shiftx4x) & (!shiftx5x) & (g218) & (!g222) & (g223) & (!g225)) + ((shiftx4x) & (!shiftx5x) & (g218) & (!g222) & (g223) & (g225)) + ((shiftx4x) & (!shiftx5x) & (g218) & (g222) & (g223) & (!g225)) + ((shiftx4x) & (!shiftx5x) & (g218) & (g222) & (g223) & (g225)) + ((shiftx4x) & (shiftx5x) & (g218) & (!g222) & (!g223) & (!g225)) + ((shiftx4x) & (shiftx5x) & (g218) & (!g222) & (!g223) & (g225)) + ((shiftx4x) & (shiftx5x) & (g218) & (!g222) & (g223) & (!g225)) + ((shiftx4x) & (shiftx5x) & (g218) & (!g222) & (g223) & (g225)) + ((shiftx4x) & (shiftx5x) & (g218) & (g222) & (!g223) & (!g225)) + ((shiftx4x) & (shiftx5x) & (g218) & (g222) & (!g223) & (g225)) + ((shiftx4x) & (shiftx5x) & (g218) & (g222) & (g223) & (!g225)) + ((shiftx4x) & (shiftx5x) & (g218) & (g222) & (g223) & (g225)));
	assign g426 = (((!shiftx4x) & (!shiftx5x) & (g217) & (!g219) & (!g220) & (!g224)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (!g219) & (!g220) & (g224)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (!g219) & (g220) & (!g224)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (!g219) & (g220) & (g224)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (g219) & (!g220) & (!g224)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (g219) & (!g220) & (g224)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (g219) & (g220) & (!g224)) + ((!shiftx4x) & (!shiftx5x) & (g217) & (g219) & (g220) & (g224)) + ((!shiftx4x) & (shiftx5x) & (!g217) & (!g219) & (g220) & (!g224)) + ((!shiftx4x) & (shiftx5x) & (!g217) & (!g219) & (g220) & (g224)) + ((!shiftx4x) & (shiftx5x) & (!g217) & (g219) & (g220) & (!g224)) + ((!shiftx4x) & (shiftx5x) & (!g217) & (g219) & (g220) & (g224)) + ((!shiftx4x) & (shiftx5x) & (g217) & (!g219) & (g220) & (!g224)) + ((!shiftx4x) & (shiftx5x) & (g217) & (!g219) & (g220) & (g224)) + ((!shiftx4x) & (shiftx5x) & (g217) & (g219) & (g220) & (!g224)) + ((!shiftx4x) & (shiftx5x) & (g217) & (g219) & (g220) & (g224)) + ((shiftx4x) & (!shiftx5x) & (!g217) & (g219) & (!g220) & (!g224)) + ((shiftx4x) & (!shiftx5x) & (!g217) & (g219) & (!g220) & (g224)) + ((shiftx4x) & (!shiftx5x) & (!g217) & (g219) & (g220) & (!g224)) + ((shiftx4x) & (!shiftx5x) & (!g217) & (g219) & (g220) & (g224)) + ((shiftx4x) & (!shiftx5x) & (g217) & (g219) & (!g220) & (!g224)) + ((shiftx4x) & (!shiftx5x) & (g217) & (g219) & (!g220) & (g224)) + ((shiftx4x) & (!shiftx5x) & (g217) & (g219) & (g220) & (!g224)) + ((shiftx4x) & (!shiftx5x) & (g217) & (g219) & (g220) & (g224)) + ((shiftx4x) & (shiftx5x) & (!g217) & (!g219) & (!g220) & (g224)) + ((shiftx4x) & (shiftx5x) & (!g217) & (!g219) & (g220) & (g224)) + ((shiftx4x) & (shiftx5x) & (!g217) & (g219) & (!g220) & (g224)) + ((shiftx4x) & (shiftx5x) & (!g217) & (g219) & (g220) & (g224)) + ((shiftx4x) & (shiftx5x) & (g217) & (!g219) & (!g220) & (g224)) + ((shiftx4x) & (shiftx5x) & (g217) & (!g219) & (g220) & (g224)) + ((shiftx4x) & (shiftx5x) & (g217) & (g219) & (!g220) & (g224)) + ((shiftx4x) & (shiftx5x) & (g217) & (g219) & (g220) & (g224)));
	assign resultx56x = (((!sk[42]) & (shiftx6x) & (!g425) & (!g426)) + ((!sk[42]) & (shiftx6x) & (!g425) & (g426)) + ((!sk[42]) & (shiftx6x) & (g425) & (!g426)) + ((!sk[42]) & (shiftx6x) & (g425) & (g426)) + ((sk[42]) & (!shiftx6x) & (!g425) & (g426)) + ((sk[42]) & (!shiftx6x) & (g425) & (g426)) + ((sk[42]) & (shiftx6x) & (g425) & (!g426)) + ((sk[42]) & (shiftx6x) & (g425) & (g426)));
	assign g428 = (((!shiftx4x) & (!shiftx5x) & (!g229) & (!g233) & (!g234) & (g236)) + ((!shiftx4x) & (!shiftx5x) & (!g229) & (!g233) & (g234) & (g236)) + ((!shiftx4x) & (!shiftx5x) & (!g229) & (g233) & (!g234) & (g236)) + ((!shiftx4x) & (!shiftx5x) & (!g229) & (g233) & (g234) & (g236)) + ((!shiftx4x) & (!shiftx5x) & (g229) & (!g233) & (!g234) & (g236)) + ((!shiftx4x) & (!shiftx5x) & (g229) & (!g233) & (g234) & (g236)) + ((!shiftx4x) & (!shiftx5x) & (g229) & (g233) & (!g234) & (g236)) + ((!shiftx4x) & (!shiftx5x) & (g229) & (g233) & (g234) & (g236)) + ((!shiftx4x) & (shiftx5x) & (!g229) & (g233) & (!g234) & (!g236)) + ((!shiftx4x) & (shiftx5x) & (!g229) & (g233) & (!g234) & (g236)) + ((!shiftx4x) & (shiftx5x) & (!g229) & (g233) & (g234) & (!g236)) + ((!shiftx4x) & (shiftx5x) & (!g229) & (g233) & (g234) & (g236)) + ((!shiftx4x) & (shiftx5x) & (g229) & (g233) & (!g234) & (!g236)) + ((!shiftx4x) & (shiftx5x) & (g229) & (g233) & (!g234) & (g236)) + ((!shiftx4x) & (shiftx5x) & (g229) & (g233) & (g234) & (!g236)) + ((!shiftx4x) & (shiftx5x) & (g229) & (g233) & (g234) & (g236)) + ((shiftx4x) & (!shiftx5x) & (!g229) & (!g233) & (g234) & (!g236)) + ((shiftx4x) & (!shiftx5x) & (!g229) & (!g233) & (g234) & (g236)) + ((shiftx4x) & (!shiftx5x) & (!g229) & (g233) & (g234) & (!g236)) + ((shiftx4x) & (!shiftx5x) & (!g229) & (g233) & (g234) & (g236)) + ((shiftx4x) & (!shiftx5x) & (g229) & (!g233) & (g234) & (!g236)) + ((shiftx4x) & (!shiftx5x) & (g229) & (!g233) & (g234) & (g236)) + ((shiftx4x) & (!shiftx5x) & (g229) & (g233) & (g234) & (!g236)) + ((shiftx4x) & (!shiftx5x) & (g229) & (g233) & (g234) & (g236)) + ((shiftx4x) & (shiftx5x) & (g229) & (!g233) & (!g234) & (!g236)) + ((shiftx4x) & (shiftx5x) & (g229) & (!g233) & (!g234) & (g236)) + ((shiftx4x) & (shiftx5x) & (g229) & (!g233) & (g234) & (!g236)) + ((shiftx4x) & (shiftx5x) & (g229) & (!g233) & (g234) & (g236)) + ((shiftx4x) & (shiftx5x) & (g229) & (g233) & (!g234) & (!g236)) + ((shiftx4x) & (shiftx5x) & (g229) & (g233) & (!g234) & (g236)) + ((shiftx4x) & (shiftx5x) & (g229) & (g233) & (g234) & (!g236)) + ((shiftx4x) & (shiftx5x) & (g229) & (g233) & (g234) & (g236)));
	assign g429 = (((!shiftx4x) & (!shiftx5x) & (g228) & (!g230) & (!g231) & (!g235)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (!g230) & (!g231) & (g235)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (!g230) & (g231) & (!g235)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (!g230) & (g231) & (g235)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (g230) & (!g231) & (!g235)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (g230) & (!g231) & (g235)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (g230) & (g231) & (!g235)) + ((!shiftx4x) & (!shiftx5x) & (g228) & (g230) & (g231) & (g235)) + ((!shiftx4x) & (shiftx5x) & (!g228) & (!g230) & (g231) & (!g235)) + ((!shiftx4x) & (shiftx5x) & (!g228) & (!g230) & (g231) & (g235)) + ((!shiftx4x) & (shiftx5x) & (!g228) & (g230) & (g231) & (!g235)) + ((!shiftx4x) & (shiftx5x) & (!g228) & (g230) & (g231) & (g235)) + ((!shiftx4x) & (shiftx5x) & (g228) & (!g230) & (g231) & (!g235)) + ((!shiftx4x) & (shiftx5x) & (g228) & (!g230) & (g231) & (g235)) + ((!shiftx4x) & (shiftx5x) & (g228) & (g230) & (g231) & (!g235)) + ((!shiftx4x) & (shiftx5x) & (g228) & (g230) & (g231) & (g235)) + ((shiftx4x) & (!shiftx5x) & (!g228) & (g230) & (!g231) & (!g235)) + ((shiftx4x) & (!shiftx5x) & (!g228) & (g230) & (!g231) & (g235)) + ((shiftx4x) & (!shiftx5x) & (!g228) & (g230) & (g231) & (!g235)) + ((shiftx4x) & (!shiftx5x) & (!g228) & (g230) & (g231) & (g235)) + ((shiftx4x) & (!shiftx5x) & (g228) & (g230) & (!g231) & (!g235)) + ((shiftx4x) & (!shiftx5x) & (g228) & (g230) & (!g231) & (g235)) + ((shiftx4x) & (!shiftx5x) & (g228) & (g230) & (g231) & (!g235)) + ((shiftx4x) & (!shiftx5x) & (g228) & (g230) & (g231) & (g235)) + ((shiftx4x) & (shiftx5x) & (!g228) & (!g230) & (!g231) & (g235)) + ((shiftx4x) & (shiftx5x) & (!g228) & (!g230) & (g231) & (g235)) + ((shiftx4x) & (shiftx5x) & (!g228) & (g230) & (!g231) & (g235)) + ((shiftx4x) & (shiftx5x) & (!g228) & (g230) & (g231) & (g235)) + ((shiftx4x) & (shiftx5x) & (g228) & (!g230) & (!g231) & (g235)) + ((shiftx4x) & (shiftx5x) & (g228) & (!g230) & (g231) & (g235)) + ((shiftx4x) & (shiftx5x) & (g228) & (g230) & (!g231) & (g235)) + ((shiftx4x) & (shiftx5x) & (g228) & (g230) & (g231) & (g235)));
	assign resultx57x = (((!shiftx6x) & (!g428) & (sk[45]) & (g429)) + ((!shiftx6x) & (g428) & (sk[45]) & (g429)) + ((shiftx6x) & (!g428) & (!sk[45]) & (!g429)) + ((shiftx6x) & (!g428) & (!sk[45]) & (g429)) + ((shiftx6x) & (g428) & (!sk[45]) & (!g429)) + ((shiftx6x) & (g428) & (!sk[45]) & (g429)) + ((shiftx6x) & (g428) & (sk[45]) & (!g429)) + ((shiftx6x) & (g428) & (sk[45]) & (g429)));
	assign g431 = (((!shiftx4x) & (!shiftx5x) & (!g240) & (!g244) & (!g245) & (g247)) + ((!shiftx4x) & (!shiftx5x) & (!g240) & (!g244) & (g245) & (g247)) + ((!shiftx4x) & (!shiftx5x) & (!g240) & (g244) & (!g245) & (g247)) + ((!shiftx4x) & (!shiftx5x) & (!g240) & (g244) & (g245) & (g247)) + ((!shiftx4x) & (!shiftx5x) & (g240) & (!g244) & (!g245) & (g247)) + ((!shiftx4x) & (!shiftx5x) & (g240) & (!g244) & (g245) & (g247)) + ((!shiftx4x) & (!shiftx5x) & (g240) & (g244) & (!g245) & (g247)) + ((!shiftx4x) & (!shiftx5x) & (g240) & (g244) & (g245) & (g247)) + ((!shiftx4x) & (shiftx5x) & (!g240) & (g244) & (!g245) & (!g247)) + ((!shiftx4x) & (shiftx5x) & (!g240) & (g244) & (!g245) & (g247)) + ((!shiftx4x) & (shiftx5x) & (!g240) & (g244) & (g245) & (!g247)) + ((!shiftx4x) & (shiftx5x) & (!g240) & (g244) & (g245) & (g247)) + ((!shiftx4x) & (shiftx5x) & (g240) & (g244) & (!g245) & (!g247)) + ((!shiftx4x) & (shiftx5x) & (g240) & (g244) & (!g245) & (g247)) + ((!shiftx4x) & (shiftx5x) & (g240) & (g244) & (g245) & (!g247)) + ((!shiftx4x) & (shiftx5x) & (g240) & (g244) & (g245) & (g247)) + ((shiftx4x) & (!shiftx5x) & (!g240) & (!g244) & (g245) & (!g247)) + ((shiftx4x) & (!shiftx5x) & (!g240) & (!g244) & (g245) & (g247)) + ((shiftx4x) & (!shiftx5x) & (!g240) & (g244) & (g245) & (!g247)) + ((shiftx4x) & (!shiftx5x) & (!g240) & (g244) & (g245) & (g247)) + ((shiftx4x) & (!shiftx5x) & (g240) & (!g244) & (g245) & (!g247)) + ((shiftx4x) & (!shiftx5x) & (g240) & (!g244) & (g245) & (g247)) + ((shiftx4x) & (!shiftx5x) & (g240) & (g244) & (g245) & (!g247)) + ((shiftx4x) & (!shiftx5x) & (g240) & (g244) & (g245) & (g247)) + ((shiftx4x) & (shiftx5x) & (g240) & (!g244) & (!g245) & (!g247)) + ((shiftx4x) & (shiftx5x) & (g240) & (!g244) & (!g245) & (g247)) + ((shiftx4x) & (shiftx5x) & (g240) & (!g244) & (g245) & (!g247)) + ((shiftx4x) & (shiftx5x) & (g240) & (!g244) & (g245) & (g247)) + ((shiftx4x) & (shiftx5x) & (g240) & (g244) & (!g245) & (!g247)) + ((shiftx4x) & (shiftx5x) & (g240) & (g244) & (!g245) & (g247)) + ((shiftx4x) & (shiftx5x) & (g240) & (g244) & (g245) & (!g247)) + ((shiftx4x) & (shiftx5x) & (g240) & (g244) & (g245) & (g247)));
	assign g432 = (((!shiftx4x) & (!shiftx5x) & (g239) & (!g241) & (!g242) & (!g246)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (!g241) & (!g242) & (g246)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (!g241) & (g242) & (!g246)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (!g241) & (g242) & (g246)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (g241) & (!g242) & (!g246)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (g241) & (!g242) & (g246)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (g241) & (g242) & (!g246)) + ((!shiftx4x) & (!shiftx5x) & (g239) & (g241) & (g242) & (g246)) + ((!shiftx4x) & (shiftx5x) & (!g239) & (!g241) & (g242) & (!g246)) + ((!shiftx4x) & (shiftx5x) & (!g239) & (!g241) & (g242) & (g246)) + ((!shiftx4x) & (shiftx5x) & (!g239) & (g241) & (g242) & (!g246)) + ((!shiftx4x) & (shiftx5x) & (!g239) & (g241) & (g242) & (g246)) + ((!shiftx4x) & (shiftx5x) & (g239) & (!g241) & (g242) & (!g246)) + ((!shiftx4x) & (shiftx5x) & (g239) & (!g241) & (g242) & (g246)) + ((!shiftx4x) & (shiftx5x) & (g239) & (g241) & (g242) & (!g246)) + ((!shiftx4x) & (shiftx5x) & (g239) & (g241) & (g242) & (g246)) + ((shiftx4x) & (!shiftx5x) & (!g239) & (g241) & (!g242) & (!g246)) + ((shiftx4x) & (!shiftx5x) & (!g239) & (g241) & (!g242) & (g246)) + ((shiftx4x) & (!shiftx5x) & (!g239) & (g241) & (g242) & (!g246)) + ((shiftx4x) & (!shiftx5x) & (!g239) & (g241) & (g242) & (g246)) + ((shiftx4x) & (!shiftx5x) & (g239) & (g241) & (!g242) & (!g246)) + ((shiftx4x) & (!shiftx5x) & (g239) & (g241) & (!g242) & (g246)) + ((shiftx4x) & (!shiftx5x) & (g239) & (g241) & (g242) & (!g246)) + ((shiftx4x) & (!shiftx5x) & (g239) & (g241) & (g242) & (g246)) + ((shiftx4x) & (shiftx5x) & (!g239) & (!g241) & (!g242) & (g246)) + ((shiftx4x) & (shiftx5x) & (!g239) & (!g241) & (g242) & (g246)) + ((shiftx4x) & (shiftx5x) & (!g239) & (g241) & (!g242) & (g246)) + ((shiftx4x) & (shiftx5x) & (!g239) & (g241) & (g242) & (g246)) + ((shiftx4x) & (shiftx5x) & (g239) & (!g241) & (!g242) & (g246)) + ((shiftx4x) & (shiftx5x) & (g239) & (!g241) & (g242) & (g246)) + ((shiftx4x) & (shiftx5x) & (g239) & (g241) & (!g242) & (g246)) + ((shiftx4x) & (shiftx5x) & (g239) & (g241) & (g242) & (g246)));
	assign resultx58x = (((!shiftx6x) & (sk[48]) & (!g431) & (g432)) + ((!shiftx6x) & (sk[48]) & (g431) & (g432)) + ((shiftx6x) & (!sk[48]) & (!g431) & (!g432)) + ((shiftx6x) & (!sk[48]) & (!g431) & (g432)) + ((shiftx6x) & (!sk[48]) & (g431) & (!g432)) + ((shiftx6x) & (!sk[48]) & (g431) & (g432)) + ((shiftx6x) & (sk[48]) & (g431) & (!g432)) + ((shiftx6x) & (sk[48]) & (g431) & (g432)));
	assign g434 = (((!shiftx4x) & (!shiftx5x) & (!g251) & (!g255) & (!g256) & (g258)) + ((!shiftx4x) & (!shiftx5x) & (!g251) & (!g255) & (g256) & (g258)) + ((!shiftx4x) & (!shiftx5x) & (!g251) & (g255) & (!g256) & (g258)) + ((!shiftx4x) & (!shiftx5x) & (!g251) & (g255) & (g256) & (g258)) + ((!shiftx4x) & (!shiftx5x) & (g251) & (!g255) & (!g256) & (g258)) + ((!shiftx4x) & (!shiftx5x) & (g251) & (!g255) & (g256) & (g258)) + ((!shiftx4x) & (!shiftx5x) & (g251) & (g255) & (!g256) & (g258)) + ((!shiftx4x) & (!shiftx5x) & (g251) & (g255) & (g256) & (g258)) + ((!shiftx4x) & (shiftx5x) & (!g251) & (g255) & (!g256) & (!g258)) + ((!shiftx4x) & (shiftx5x) & (!g251) & (g255) & (!g256) & (g258)) + ((!shiftx4x) & (shiftx5x) & (!g251) & (g255) & (g256) & (!g258)) + ((!shiftx4x) & (shiftx5x) & (!g251) & (g255) & (g256) & (g258)) + ((!shiftx4x) & (shiftx5x) & (g251) & (g255) & (!g256) & (!g258)) + ((!shiftx4x) & (shiftx5x) & (g251) & (g255) & (!g256) & (g258)) + ((!shiftx4x) & (shiftx5x) & (g251) & (g255) & (g256) & (!g258)) + ((!shiftx4x) & (shiftx5x) & (g251) & (g255) & (g256) & (g258)) + ((shiftx4x) & (!shiftx5x) & (!g251) & (!g255) & (g256) & (!g258)) + ((shiftx4x) & (!shiftx5x) & (!g251) & (!g255) & (g256) & (g258)) + ((shiftx4x) & (!shiftx5x) & (!g251) & (g255) & (g256) & (!g258)) + ((shiftx4x) & (!shiftx5x) & (!g251) & (g255) & (g256) & (g258)) + ((shiftx4x) & (!shiftx5x) & (g251) & (!g255) & (g256) & (!g258)) + ((shiftx4x) & (!shiftx5x) & (g251) & (!g255) & (g256) & (g258)) + ((shiftx4x) & (!shiftx5x) & (g251) & (g255) & (g256) & (!g258)) + ((shiftx4x) & (!shiftx5x) & (g251) & (g255) & (g256) & (g258)) + ((shiftx4x) & (shiftx5x) & (g251) & (!g255) & (!g256) & (!g258)) + ((shiftx4x) & (shiftx5x) & (g251) & (!g255) & (!g256) & (g258)) + ((shiftx4x) & (shiftx5x) & (g251) & (!g255) & (g256) & (!g258)) + ((shiftx4x) & (shiftx5x) & (g251) & (!g255) & (g256) & (g258)) + ((shiftx4x) & (shiftx5x) & (g251) & (g255) & (!g256) & (!g258)) + ((shiftx4x) & (shiftx5x) & (g251) & (g255) & (!g256) & (g258)) + ((shiftx4x) & (shiftx5x) & (g251) & (g255) & (g256) & (!g258)) + ((shiftx4x) & (shiftx5x) & (g251) & (g255) & (g256) & (g258)));
	assign g435 = (((!shiftx4x) & (!shiftx5x) & (g250) & (!g252) & (!g253) & (!g257)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (!g252) & (!g253) & (g257)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (!g252) & (g253) & (!g257)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (!g252) & (g253) & (g257)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (g252) & (!g253) & (!g257)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (g252) & (!g253) & (g257)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (g252) & (g253) & (!g257)) + ((!shiftx4x) & (!shiftx5x) & (g250) & (g252) & (g253) & (g257)) + ((!shiftx4x) & (shiftx5x) & (!g250) & (!g252) & (g253) & (!g257)) + ((!shiftx4x) & (shiftx5x) & (!g250) & (!g252) & (g253) & (g257)) + ((!shiftx4x) & (shiftx5x) & (!g250) & (g252) & (g253) & (!g257)) + ((!shiftx4x) & (shiftx5x) & (!g250) & (g252) & (g253) & (g257)) + ((!shiftx4x) & (shiftx5x) & (g250) & (!g252) & (g253) & (!g257)) + ((!shiftx4x) & (shiftx5x) & (g250) & (!g252) & (g253) & (g257)) + ((!shiftx4x) & (shiftx5x) & (g250) & (g252) & (g253) & (!g257)) + ((!shiftx4x) & (shiftx5x) & (g250) & (g252) & (g253) & (g257)) + ((shiftx4x) & (!shiftx5x) & (!g250) & (g252) & (!g253) & (!g257)) + ((shiftx4x) & (!shiftx5x) & (!g250) & (g252) & (!g253) & (g257)) + ((shiftx4x) & (!shiftx5x) & (!g250) & (g252) & (g253) & (!g257)) + ((shiftx4x) & (!shiftx5x) & (!g250) & (g252) & (g253) & (g257)) + ((shiftx4x) & (!shiftx5x) & (g250) & (g252) & (!g253) & (!g257)) + ((shiftx4x) & (!shiftx5x) & (g250) & (g252) & (!g253) & (g257)) + ((shiftx4x) & (!shiftx5x) & (g250) & (g252) & (g253) & (!g257)) + ((shiftx4x) & (!shiftx5x) & (g250) & (g252) & (g253) & (g257)) + ((shiftx4x) & (shiftx5x) & (!g250) & (!g252) & (!g253) & (g257)) + ((shiftx4x) & (shiftx5x) & (!g250) & (!g252) & (g253) & (g257)) + ((shiftx4x) & (shiftx5x) & (!g250) & (g252) & (!g253) & (g257)) + ((shiftx4x) & (shiftx5x) & (!g250) & (g252) & (g253) & (g257)) + ((shiftx4x) & (shiftx5x) & (g250) & (!g252) & (!g253) & (g257)) + ((shiftx4x) & (shiftx5x) & (g250) & (!g252) & (g253) & (g257)) + ((shiftx4x) & (shiftx5x) & (g250) & (g252) & (!g253) & (g257)) + ((shiftx4x) & (shiftx5x) & (g250) & (g252) & (g253) & (g257)));
	assign resultx59x = (((!sk[51]) & (shiftx6x) & (!g434) & (!g435)) + ((!sk[51]) & (shiftx6x) & (!g434) & (g435)) + ((!sk[51]) & (shiftx6x) & (g434) & (!g435)) + ((!sk[51]) & (shiftx6x) & (g434) & (g435)) + ((sk[51]) & (!shiftx6x) & (!g434) & (g435)) + ((sk[51]) & (!shiftx6x) & (g434) & (g435)) + ((sk[51]) & (shiftx6x) & (g434) & (!g435)) + ((sk[51]) & (shiftx6x) & (g434) & (g435)));
	assign g437 = (((!shiftx4x) & (!shiftx5x) & (!g262) & (!g266) & (!g267) & (g269)) + ((!shiftx4x) & (!shiftx5x) & (!g262) & (!g266) & (g267) & (g269)) + ((!shiftx4x) & (!shiftx5x) & (!g262) & (g266) & (!g267) & (g269)) + ((!shiftx4x) & (!shiftx5x) & (!g262) & (g266) & (g267) & (g269)) + ((!shiftx4x) & (!shiftx5x) & (g262) & (!g266) & (!g267) & (g269)) + ((!shiftx4x) & (!shiftx5x) & (g262) & (!g266) & (g267) & (g269)) + ((!shiftx4x) & (!shiftx5x) & (g262) & (g266) & (!g267) & (g269)) + ((!shiftx4x) & (!shiftx5x) & (g262) & (g266) & (g267) & (g269)) + ((!shiftx4x) & (shiftx5x) & (!g262) & (g266) & (!g267) & (!g269)) + ((!shiftx4x) & (shiftx5x) & (!g262) & (g266) & (!g267) & (g269)) + ((!shiftx4x) & (shiftx5x) & (!g262) & (g266) & (g267) & (!g269)) + ((!shiftx4x) & (shiftx5x) & (!g262) & (g266) & (g267) & (g269)) + ((!shiftx4x) & (shiftx5x) & (g262) & (g266) & (!g267) & (!g269)) + ((!shiftx4x) & (shiftx5x) & (g262) & (g266) & (!g267) & (g269)) + ((!shiftx4x) & (shiftx5x) & (g262) & (g266) & (g267) & (!g269)) + ((!shiftx4x) & (shiftx5x) & (g262) & (g266) & (g267) & (g269)) + ((shiftx4x) & (!shiftx5x) & (!g262) & (!g266) & (g267) & (!g269)) + ((shiftx4x) & (!shiftx5x) & (!g262) & (!g266) & (g267) & (g269)) + ((shiftx4x) & (!shiftx5x) & (!g262) & (g266) & (g267) & (!g269)) + ((shiftx4x) & (!shiftx5x) & (!g262) & (g266) & (g267) & (g269)) + ((shiftx4x) & (!shiftx5x) & (g262) & (!g266) & (g267) & (!g269)) + ((shiftx4x) & (!shiftx5x) & (g262) & (!g266) & (g267) & (g269)) + ((shiftx4x) & (!shiftx5x) & (g262) & (g266) & (g267) & (!g269)) + ((shiftx4x) & (!shiftx5x) & (g262) & (g266) & (g267) & (g269)) + ((shiftx4x) & (shiftx5x) & (g262) & (!g266) & (!g267) & (!g269)) + ((shiftx4x) & (shiftx5x) & (g262) & (!g266) & (!g267) & (g269)) + ((shiftx4x) & (shiftx5x) & (g262) & (!g266) & (g267) & (!g269)) + ((shiftx4x) & (shiftx5x) & (g262) & (!g266) & (g267) & (g269)) + ((shiftx4x) & (shiftx5x) & (g262) & (g266) & (!g267) & (!g269)) + ((shiftx4x) & (shiftx5x) & (g262) & (g266) & (!g267) & (g269)) + ((shiftx4x) & (shiftx5x) & (g262) & (g266) & (g267) & (!g269)) + ((shiftx4x) & (shiftx5x) & (g262) & (g266) & (g267) & (g269)));
	assign g438 = (((!shiftx4x) & (!shiftx5x) & (g261) & (!g263) & (!g264) & (!g268)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (!g263) & (!g264) & (g268)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (!g263) & (g264) & (!g268)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (!g263) & (g264) & (g268)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (g263) & (!g264) & (!g268)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (g263) & (!g264) & (g268)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (g263) & (g264) & (!g268)) + ((!shiftx4x) & (!shiftx5x) & (g261) & (g263) & (g264) & (g268)) + ((!shiftx4x) & (shiftx5x) & (!g261) & (!g263) & (g264) & (!g268)) + ((!shiftx4x) & (shiftx5x) & (!g261) & (!g263) & (g264) & (g268)) + ((!shiftx4x) & (shiftx5x) & (!g261) & (g263) & (g264) & (!g268)) + ((!shiftx4x) & (shiftx5x) & (!g261) & (g263) & (g264) & (g268)) + ((!shiftx4x) & (shiftx5x) & (g261) & (!g263) & (g264) & (!g268)) + ((!shiftx4x) & (shiftx5x) & (g261) & (!g263) & (g264) & (g268)) + ((!shiftx4x) & (shiftx5x) & (g261) & (g263) & (g264) & (!g268)) + ((!shiftx4x) & (shiftx5x) & (g261) & (g263) & (g264) & (g268)) + ((shiftx4x) & (!shiftx5x) & (!g261) & (g263) & (!g264) & (!g268)) + ((shiftx4x) & (!shiftx5x) & (!g261) & (g263) & (!g264) & (g268)) + ((shiftx4x) & (!shiftx5x) & (!g261) & (g263) & (g264) & (!g268)) + ((shiftx4x) & (!shiftx5x) & (!g261) & (g263) & (g264) & (g268)) + ((shiftx4x) & (!shiftx5x) & (g261) & (g263) & (!g264) & (!g268)) + ((shiftx4x) & (!shiftx5x) & (g261) & (g263) & (!g264) & (g268)) + ((shiftx4x) & (!shiftx5x) & (g261) & (g263) & (g264) & (!g268)) + ((shiftx4x) & (!shiftx5x) & (g261) & (g263) & (g264) & (g268)) + ((shiftx4x) & (shiftx5x) & (!g261) & (!g263) & (!g264) & (g268)) + ((shiftx4x) & (shiftx5x) & (!g261) & (!g263) & (g264) & (g268)) + ((shiftx4x) & (shiftx5x) & (!g261) & (g263) & (!g264) & (g268)) + ((shiftx4x) & (shiftx5x) & (!g261) & (g263) & (g264) & (g268)) + ((shiftx4x) & (shiftx5x) & (g261) & (!g263) & (!g264) & (g268)) + ((shiftx4x) & (shiftx5x) & (g261) & (!g263) & (g264) & (g268)) + ((shiftx4x) & (shiftx5x) & (g261) & (g263) & (!g264) & (g268)) + ((shiftx4x) & (shiftx5x) & (g261) & (g263) & (g264) & (g268)));
	assign resultx60x = (((!shiftx6x) & (!g437) & (sk[54]) & (g438)) + ((!shiftx6x) & (g437) & (sk[54]) & (g438)) + ((shiftx6x) & (!g437) & (!sk[54]) & (!g438)) + ((shiftx6x) & (!g437) & (!sk[54]) & (g438)) + ((shiftx6x) & (g437) & (!sk[54]) & (!g438)) + ((shiftx6x) & (g437) & (!sk[54]) & (g438)) + ((shiftx6x) & (g437) & (sk[54]) & (!g438)) + ((shiftx6x) & (g437) & (sk[54]) & (g438)));
	assign g440 = (((!shiftx4x) & (!shiftx5x) & (!g273) & (!g277) & (!g278) & (g280)) + ((!shiftx4x) & (!shiftx5x) & (!g273) & (!g277) & (g278) & (g280)) + ((!shiftx4x) & (!shiftx5x) & (!g273) & (g277) & (!g278) & (g280)) + ((!shiftx4x) & (!shiftx5x) & (!g273) & (g277) & (g278) & (g280)) + ((!shiftx4x) & (!shiftx5x) & (g273) & (!g277) & (!g278) & (g280)) + ((!shiftx4x) & (!shiftx5x) & (g273) & (!g277) & (g278) & (g280)) + ((!shiftx4x) & (!shiftx5x) & (g273) & (g277) & (!g278) & (g280)) + ((!shiftx4x) & (!shiftx5x) & (g273) & (g277) & (g278) & (g280)) + ((!shiftx4x) & (shiftx5x) & (!g273) & (g277) & (!g278) & (!g280)) + ((!shiftx4x) & (shiftx5x) & (!g273) & (g277) & (!g278) & (g280)) + ((!shiftx4x) & (shiftx5x) & (!g273) & (g277) & (g278) & (!g280)) + ((!shiftx4x) & (shiftx5x) & (!g273) & (g277) & (g278) & (g280)) + ((!shiftx4x) & (shiftx5x) & (g273) & (g277) & (!g278) & (!g280)) + ((!shiftx4x) & (shiftx5x) & (g273) & (g277) & (!g278) & (g280)) + ((!shiftx4x) & (shiftx5x) & (g273) & (g277) & (g278) & (!g280)) + ((!shiftx4x) & (shiftx5x) & (g273) & (g277) & (g278) & (g280)) + ((shiftx4x) & (!shiftx5x) & (!g273) & (!g277) & (g278) & (!g280)) + ((shiftx4x) & (!shiftx5x) & (!g273) & (!g277) & (g278) & (g280)) + ((shiftx4x) & (!shiftx5x) & (!g273) & (g277) & (g278) & (!g280)) + ((shiftx4x) & (!shiftx5x) & (!g273) & (g277) & (g278) & (g280)) + ((shiftx4x) & (!shiftx5x) & (g273) & (!g277) & (g278) & (!g280)) + ((shiftx4x) & (!shiftx5x) & (g273) & (!g277) & (g278) & (g280)) + ((shiftx4x) & (!shiftx5x) & (g273) & (g277) & (g278) & (!g280)) + ((shiftx4x) & (!shiftx5x) & (g273) & (g277) & (g278) & (g280)) + ((shiftx4x) & (shiftx5x) & (g273) & (!g277) & (!g278) & (!g280)) + ((shiftx4x) & (shiftx5x) & (g273) & (!g277) & (!g278) & (g280)) + ((shiftx4x) & (shiftx5x) & (g273) & (!g277) & (g278) & (!g280)) + ((shiftx4x) & (shiftx5x) & (g273) & (!g277) & (g278) & (g280)) + ((shiftx4x) & (shiftx5x) & (g273) & (g277) & (!g278) & (!g280)) + ((shiftx4x) & (shiftx5x) & (g273) & (g277) & (!g278) & (g280)) + ((shiftx4x) & (shiftx5x) & (g273) & (g277) & (g278) & (!g280)) + ((shiftx4x) & (shiftx5x) & (g273) & (g277) & (g278) & (g280)));
	assign g441 = (((!shiftx4x) & (!shiftx5x) & (g272) & (!g274) & (!g275) & (!g279)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (!g274) & (!g275) & (g279)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (!g274) & (g275) & (!g279)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (!g274) & (g275) & (g279)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (g274) & (!g275) & (!g279)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (g274) & (!g275) & (g279)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (g274) & (g275) & (!g279)) + ((!shiftx4x) & (!shiftx5x) & (g272) & (g274) & (g275) & (g279)) + ((!shiftx4x) & (shiftx5x) & (!g272) & (!g274) & (g275) & (!g279)) + ((!shiftx4x) & (shiftx5x) & (!g272) & (!g274) & (g275) & (g279)) + ((!shiftx4x) & (shiftx5x) & (!g272) & (g274) & (g275) & (!g279)) + ((!shiftx4x) & (shiftx5x) & (!g272) & (g274) & (g275) & (g279)) + ((!shiftx4x) & (shiftx5x) & (g272) & (!g274) & (g275) & (!g279)) + ((!shiftx4x) & (shiftx5x) & (g272) & (!g274) & (g275) & (g279)) + ((!shiftx4x) & (shiftx5x) & (g272) & (g274) & (g275) & (!g279)) + ((!shiftx4x) & (shiftx5x) & (g272) & (g274) & (g275) & (g279)) + ((shiftx4x) & (!shiftx5x) & (!g272) & (g274) & (!g275) & (!g279)) + ((shiftx4x) & (!shiftx5x) & (!g272) & (g274) & (!g275) & (g279)) + ((shiftx4x) & (!shiftx5x) & (!g272) & (g274) & (g275) & (!g279)) + ((shiftx4x) & (!shiftx5x) & (!g272) & (g274) & (g275) & (g279)) + ((shiftx4x) & (!shiftx5x) & (g272) & (g274) & (!g275) & (!g279)) + ((shiftx4x) & (!shiftx5x) & (g272) & (g274) & (!g275) & (g279)) + ((shiftx4x) & (!shiftx5x) & (g272) & (g274) & (g275) & (!g279)) + ((shiftx4x) & (!shiftx5x) & (g272) & (g274) & (g275) & (g279)) + ((shiftx4x) & (shiftx5x) & (!g272) & (!g274) & (!g275) & (g279)) + ((shiftx4x) & (shiftx5x) & (!g272) & (!g274) & (g275) & (g279)) + ((shiftx4x) & (shiftx5x) & (!g272) & (g274) & (!g275) & (g279)) + ((shiftx4x) & (shiftx5x) & (!g272) & (g274) & (g275) & (g279)) + ((shiftx4x) & (shiftx5x) & (g272) & (!g274) & (!g275) & (g279)) + ((shiftx4x) & (shiftx5x) & (g272) & (!g274) & (g275) & (g279)) + ((shiftx4x) & (shiftx5x) & (g272) & (g274) & (!g275) & (g279)) + ((shiftx4x) & (shiftx5x) & (g272) & (g274) & (g275) & (g279)));
	assign resultx61x = (((!shiftx6x) & (sk[57]) & (!g440) & (g441)) + ((!shiftx6x) & (sk[57]) & (g440) & (g441)) + ((shiftx6x) & (!sk[57]) & (!g440) & (!g441)) + ((shiftx6x) & (!sk[57]) & (!g440) & (g441)) + ((shiftx6x) & (!sk[57]) & (g440) & (!g441)) + ((shiftx6x) & (!sk[57]) & (g440) & (g441)) + ((shiftx6x) & (sk[57]) & (g440) & (!g441)) + ((shiftx6x) & (sk[57]) & (g440) & (g441)));
	assign g443 = (((!shiftx4x) & (!shiftx5x) & (!g284) & (!g288) & (!g289) & (g291)) + ((!shiftx4x) & (!shiftx5x) & (!g284) & (!g288) & (g289) & (g291)) + ((!shiftx4x) & (!shiftx5x) & (!g284) & (g288) & (!g289) & (g291)) + ((!shiftx4x) & (!shiftx5x) & (!g284) & (g288) & (g289) & (g291)) + ((!shiftx4x) & (!shiftx5x) & (g284) & (!g288) & (!g289) & (g291)) + ((!shiftx4x) & (!shiftx5x) & (g284) & (!g288) & (g289) & (g291)) + ((!shiftx4x) & (!shiftx5x) & (g284) & (g288) & (!g289) & (g291)) + ((!shiftx4x) & (!shiftx5x) & (g284) & (g288) & (g289) & (g291)) + ((!shiftx4x) & (shiftx5x) & (!g284) & (g288) & (!g289) & (!g291)) + ((!shiftx4x) & (shiftx5x) & (!g284) & (g288) & (!g289) & (g291)) + ((!shiftx4x) & (shiftx5x) & (!g284) & (g288) & (g289) & (!g291)) + ((!shiftx4x) & (shiftx5x) & (!g284) & (g288) & (g289) & (g291)) + ((!shiftx4x) & (shiftx5x) & (g284) & (g288) & (!g289) & (!g291)) + ((!shiftx4x) & (shiftx5x) & (g284) & (g288) & (!g289) & (g291)) + ((!shiftx4x) & (shiftx5x) & (g284) & (g288) & (g289) & (!g291)) + ((!shiftx4x) & (shiftx5x) & (g284) & (g288) & (g289) & (g291)) + ((shiftx4x) & (!shiftx5x) & (!g284) & (!g288) & (g289) & (!g291)) + ((shiftx4x) & (!shiftx5x) & (!g284) & (!g288) & (g289) & (g291)) + ((shiftx4x) & (!shiftx5x) & (!g284) & (g288) & (g289) & (!g291)) + ((shiftx4x) & (!shiftx5x) & (!g284) & (g288) & (g289) & (g291)) + ((shiftx4x) & (!shiftx5x) & (g284) & (!g288) & (g289) & (!g291)) + ((shiftx4x) & (!shiftx5x) & (g284) & (!g288) & (g289) & (g291)) + ((shiftx4x) & (!shiftx5x) & (g284) & (g288) & (g289) & (!g291)) + ((shiftx4x) & (!shiftx5x) & (g284) & (g288) & (g289) & (g291)) + ((shiftx4x) & (shiftx5x) & (g284) & (!g288) & (!g289) & (!g291)) + ((shiftx4x) & (shiftx5x) & (g284) & (!g288) & (!g289) & (g291)) + ((shiftx4x) & (shiftx5x) & (g284) & (!g288) & (g289) & (!g291)) + ((shiftx4x) & (shiftx5x) & (g284) & (!g288) & (g289) & (g291)) + ((shiftx4x) & (shiftx5x) & (g284) & (g288) & (!g289) & (!g291)) + ((shiftx4x) & (shiftx5x) & (g284) & (g288) & (!g289) & (g291)) + ((shiftx4x) & (shiftx5x) & (g284) & (g288) & (g289) & (!g291)) + ((shiftx4x) & (shiftx5x) & (g284) & (g288) & (g289) & (g291)));
	assign g444 = (((!shiftx4x) & (!shiftx5x) & (g283) & (!g285) & (!g286) & (!g290)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (!g285) & (!g286) & (g290)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (!g285) & (g286) & (!g290)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (!g285) & (g286) & (g290)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (g285) & (!g286) & (!g290)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (g285) & (!g286) & (g290)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (g285) & (g286) & (!g290)) + ((!shiftx4x) & (!shiftx5x) & (g283) & (g285) & (g286) & (g290)) + ((!shiftx4x) & (shiftx5x) & (!g283) & (!g285) & (g286) & (!g290)) + ((!shiftx4x) & (shiftx5x) & (!g283) & (!g285) & (g286) & (g290)) + ((!shiftx4x) & (shiftx5x) & (!g283) & (g285) & (g286) & (!g290)) + ((!shiftx4x) & (shiftx5x) & (!g283) & (g285) & (g286) & (g290)) + ((!shiftx4x) & (shiftx5x) & (g283) & (!g285) & (g286) & (!g290)) + ((!shiftx4x) & (shiftx5x) & (g283) & (!g285) & (g286) & (g290)) + ((!shiftx4x) & (shiftx5x) & (g283) & (g285) & (g286) & (!g290)) + ((!shiftx4x) & (shiftx5x) & (g283) & (g285) & (g286) & (g290)) + ((shiftx4x) & (!shiftx5x) & (!g283) & (g285) & (!g286) & (!g290)) + ((shiftx4x) & (!shiftx5x) & (!g283) & (g285) & (!g286) & (g290)) + ((shiftx4x) & (!shiftx5x) & (!g283) & (g285) & (g286) & (!g290)) + ((shiftx4x) & (!shiftx5x) & (!g283) & (g285) & (g286) & (g290)) + ((shiftx4x) & (!shiftx5x) & (g283) & (g285) & (!g286) & (!g290)) + ((shiftx4x) & (!shiftx5x) & (g283) & (g285) & (!g286) & (g290)) + ((shiftx4x) & (!shiftx5x) & (g283) & (g285) & (g286) & (!g290)) + ((shiftx4x) & (!shiftx5x) & (g283) & (g285) & (g286) & (g290)) + ((shiftx4x) & (shiftx5x) & (!g283) & (!g285) & (!g286) & (g290)) + ((shiftx4x) & (shiftx5x) & (!g283) & (!g285) & (g286) & (g290)) + ((shiftx4x) & (shiftx5x) & (!g283) & (g285) & (!g286) & (g290)) + ((shiftx4x) & (shiftx5x) & (!g283) & (g285) & (g286) & (g290)) + ((shiftx4x) & (shiftx5x) & (g283) & (!g285) & (!g286) & (g290)) + ((shiftx4x) & (shiftx5x) & (g283) & (!g285) & (g286) & (g290)) + ((shiftx4x) & (shiftx5x) & (g283) & (g285) & (!g286) & (g290)) + ((shiftx4x) & (shiftx5x) & (g283) & (g285) & (g286) & (g290)));
	assign resultx62x = (((!sk[60]) & (shiftx6x) & (!g443) & (!g444)) + ((!sk[60]) & (shiftx6x) & (!g443) & (g444)) + ((!sk[60]) & (shiftx6x) & (g443) & (!g444)) + ((!sk[60]) & (shiftx6x) & (g443) & (g444)) + ((sk[60]) & (!shiftx6x) & (!g443) & (g444)) + ((sk[60]) & (!shiftx6x) & (g443) & (g444)) + ((sk[60]) & (shiftx6x) & (g443) & (!g444)) + ((sk[60]) & (shiftx6x) & (g443) & (g444)));
	assign g446 = (((!shiftx4x) & (!shiftx5x) & (!g295) & (!g299) & (!g300) & (g302)) + ((!shiftx4x) & (!shiftx5x) & (!g295) & (!g299) & (g300) & (g302)) + ((!shiftx4x) & (!shiftx5x) & (!g295) & (g299) & (!g300) & (g302)) + ((!shiftx4x) & (!shiftx5x) & (!g295) & (g299) & (g300) & (g302)) + ((!shiftx4x) & (!shiftx5x) & (g295) & (!g299) & (!g300) & (g302)) + ((!shiftx4x) & (!shiftx5x) & (g295) & (!g299) & (g300) & (g302)) + ((!shiftx4x) & (!shiftx5x) & (g295) & (g299) & (!g300) & (g302)) + ((!shiftx4x) & (!shiftx5x) & (g295) & (g299) & (g300) & (g302)) + ((!shiftx4x) & (shiftx5x) & (!g295) & (g299) & (!g300) & (!g302)) + ((!shiftx4x) & (shiftx5x) & (!g295) & (g299) & (!g300) & (g302)) + ((!shiftx4x) & (shiftx5x) & (!g295) & (g299) & (g300) & (!g302)) + ((!shiftx4x) & (shiftx5x) & (!g295) & (g299) & (g300) & (g302)) + ((!shiftx4x) & (shiftx5x) & (g295) & (g299) & (!g300) & (!g302)) + ((!shiftx4x) & (shiftx5x) & (g295) & (g299) & (!g300) & (g302)) + ((!shiftx4x) & (shiftx5x) & (g295) & (g299) & (g300) & (!g302)) + ((!shiftx4x) & (shiftx5x) & (g295) & (g299) & (g300) & (g302)) + ((shiftx4x) & (!shiftx5x) & (!g295) & (!g299) & (g300) & (!g302)) + ((shiftx4x) & (!shiftx5x) & (!g295) & (!g299) & (g300) & (g302)) + ((shiftx4x) & (!shiftx5x) & (!g295) & (g299) & (g300) & (!g302)) + ((shiftx4x) & (!shiftx5x) & (!g295) & (g299) & (g300) & (g302)) + ((shiftx4x) & (!shiftx5x) & (g295) & (!g299) & (g300) & (!g302)) + ((shiftx4x) & (!shiftx5x) & (g295) & (!g299) & (g300) & (g302)) + ((shiftx4x) & (!shiftx5x) & (g295) & (g299) & (g300) & (!g302)) + ((shiftx4x) & (!shiftx5x) & (g295) & (g299) & (g300) & (g302)) + ((shiftx4x) & (shiftx5x) & (g295) & (!g299) & (!g300) & (!g302)) + ((shiftx4x) & (shiftx5x) & (g295) & (!g299) & (!g300) & (g302)) + ((shiftx4x) & (shiftx5x) & (g295) & (!g299) & (g300) & (!g302)) + ((shiftx4x) & (shiftx5x) & (g295) & (!g299) & (g300) & (g302)) + ((shiftx4x) & (shiftx5x) & (g295) & (g299) & (!g300) & (!g302)) + ((shiftx4x) & (shiftx5x) & (g295) & (g299) & (!g300) & (g302)) + ((shiftx4x) & (shiftx5x) & (g295) & (g299) & (g300) & (!g302)) + ((shiftx4x) & (shiftx5x) & (g295) & (g299) & (g300) & (g302)));
	assign g447 = (((!shiftx4x) & (!shiftx5x) & (g294) & (!g296) & (!g297) & (!g301)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (!g296) & (!g297) & (g301)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (!g296) & (g297) & (!g301)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (!g296) & (g297) & (g301)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (g296) & (!g297) & (!g301)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (g296) & (!g297) & (g301)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (g296) & (g297) & (!g301)) + ((!shiftx4x) & (!shiftx5x) & (g294) & (g296) & (g297) & (g301)) + ((!shiftx4x) & (shiftx5x) & (!g294) & (!g296) & (g297) & (!g301)) + ((!shiftx4x) & (shiftx5x) & (!g294) & (!g296) & (g297) & (g301)) + ((!shiftx4x) & (shiftx5x) & (!g294) & (g296) & (g297) & (!g301)) + ((!shiftx4x) & (shiftx5x) & (!g294) & (g296) & (g297) & (g301)) + ((!shiftx4x) & (shiftx5x) & (g294) & (!g296) & (g297) & (!g301)) + ((!shiftx4x) & (shiftx5x) & (g294) & (!g296) & (g297) & (g301)) + ((!shiftx4x) & (shiftx5x) & (g294) & (g296) & (g297) & (!g301)) + ((!shiftx4x) & (shiftx5x) & (g294) & (g296) & (g297) & (g301)) + ((shiftx4x) & (!shiftx5x) & (!g294) & (g296) & (!g297) & (!g301)) + ((shiftx4x) & (!shiftx5x) & (!g294) & (g296) & (!g297) & (g301)) + ((shiftx4x) & (!shiftx5x) & (!g294) & (g296) & (g297) & (!g301)) + ((shiftx4x) & (!shiftx5x) & (!g294) & (g296) & (g297) & (g301)) + ((shiftx4x) & (!shiftx5x) & (g294) & (g296) & (!g297) & (!g301)) + ((shiftx4x) & (!shiftx5x) & (g294) & (g296) & (!g297) & (g301)) + ((shiftx4x) & (!shiftx5x) & (g294) & (g296) & (g297) & (!g301)) + ((shiftx4x) & (!shiftx5x) & (g294) & (g296) & (g297) & (g301)) + ((shiftx4x) & (shiftx5x) & (!g294) & (!g296) & (!g297) & (g301)) + ((shiftx4x) & (shiftx5x) & (!g294) & (!g296) & (g297) & (g301)) + ((shiftx4x) & (shiftx5x) & (!g294) & (g296) & (!g297) & (g301)) + ((shiftx4x) & (shiftx5x) & (!g294) & (g296) & (g297) & (g301)) + ((shiftx4x) & (shiftx5x) & (g294) & (!g296) & (!g297) & (g301)) + ((shiftx4x) & (shiftx5x) & (g294) & (!g296) & (g297) & (g301)) + ((shiftx4x) & (shiftx5x) & (g294) & (g296) & (!g297) & (g301)) + ((shiftx4x) & (shiftx5x) & (g294) & (g296) & (g297) & (g301)));
	assign resultx63x = (((!shiftx6x) & (sk[63]) & (!g446) & (g447)) + ((!shiftx6x) & (sk[63]) & (g446) & (g447)) + ((shiftx6x) & (!sk[63]) & (!g446) & (!g447)) + ((shiftx6x) & (!sk[63]) & (!g446) & (g447)) + ((shiftx6x) & (!sk[63]) & (g446) & (!g447)) + ((shiftx6x) & (!sk[63]) & (g446) & (g447)) + ((shiftx6x) & (sk[63]) & (g446) & (!g447)) + ((shiftx6x) & (sk[63]) & (g446) & (g447)));
	assign resultx64x = (((!sk[64]) & (shiftx6x) & (!g21) & (!g42)) + ((!sk[64]) & (shiftx6x) & (!g21) & (g42)) + ((!sk[64]) & (shiftx6x) & (g21) & (!g42)) + ((!sk[64]) & (shiftx6x) & (g21) & (g42)) + ((sk[64]) & (!shiftx6x) & (g21) & (!g42)) + ((sk[64]) & (!shiftx6x) & (g21) & (g42)) + ((sk[64]) & (shiftx6x) & (!g21) & (g42)) + ((sk[64]) & (shiftx6x) & (g21) & (g42)));
	assign resultx65x = (((!sk[65]) & (shiftx6x) & (!g64) & (!g85)) + ((!sk[65]) & (shiftx6x) & (!g64) & (g85)) + ((!sk[65]) & (shiftx6x) & (g64) & (!g85)) + ((!sk[65]) & (shiftx6x) & (g64) & (g85)) + ((sk[65]) & (!shiftx6x) & (g64) & (!g85)) + ((sk[65]) & (!shiftx6x) & (g64) & (g85)) + ((sk[65]) & (shiftx6x) & (!g64) & (g85)) + ((sk[65]) & (shiftx6x) & (g64) & (g85)));
	assign resultx66x = (((!sk[66]) & (shiftx6x) & (!g107) & (!g128)) + ((!sk[66]) & (shiftx6x) & (!g107) & (g128)) + ((!sk[66]) & (shiftx6x) & (g107) & (!g128)) + ((!sk[66]) & (shiftx6x) & (g107) & (g128)) + ((sk[66]) & (!shiftx6x) & (g107) & (!g128)) + ((sk[66]) & (!shiftx6x) & (g107) & (g128)) + ((sk[66]) & (shiftx6x) & (!g107) & (g128)) + ((sk[66]) & (shiftx6x) & (g107) & (g128)));
	assign resultx67x = (((!shiftx6x) & (sk[67]) & (g150) & (!g171)) + ((!shiftx6x) & (sk[67]) & (g150) & (g171)) + ((shiftx6x) & (!sk[67]) & (!g150) & (!g171)) + ((shiftx6x) & (!sk[67]) & (!g150) & (g171)) + ((shiftx6x) & (!sk[67]) & (g150) & (!g171)) + ((shiftx6x) & (!sk[67]) & (g150) & (g171)) + ((shiftx6x) & (sk[67]) & (!g150) & (g171)) + ((shiftx6x) & (sk[67]) & (g150) & (g171)));
	assign resultx68x = (((!sk[68]) & (shiftx6x) & (!g177) & (!g182)) + ((!sk[68]) & (shiftx6x) & (!g177) & (g182)) + ((!sk[68]) & (shiftx6x) & (g177) & (!g182)) + ((!sk[68]) & (shiftx6x) & (g177) & (g182)) + ((sk[68]) & (!shiftx6x) & (g177) & (!g182)) + ((sk[68]) & (!shiftx6x) & (g177) & (g182)) + ((sk[68]) & (shiftx6x) & (!g177) & (g182)) + ((sk[68]) & (shiftx6x) & (g177) & (g182)));
	assign resultx69x = (((!sk[69]) & (shiftx6x) & (!g188) & (!g193)) + ((!sk[69]) & (shiftx6x) & (!g188) & (g193)) + ((!sk[69]) & (shiftx6x) & (g188) & (!g193)) + ((!sk[69]) & (shiftx6x) & (g188) & (g193)) + ((sk[69]) & (!shiftx6x) & (g188) & (!g193)) + ((sk[69]) & (!shiftx6x) & (g188) & (g193)) + ((sk[69]) & (shiftx6x) & (!g188) & (g193)) + ((sk[69]) & (shiftx6x) & (g188) & (g193)));
	assign resultx70x = (((!sk[70]) & (shiftx6x) & (!g199) & (!g204)) + ((!sk[70]) & (shiftx6x) & (!g199) & (g204)) + ((!sk[70]) & (shiftx6x) & (g199) & (!g204)) + ((!sk[70]) & (shiftx6x) & (g199) & (g204)) + ((sk[70]) & (!shiftx6x) & (g199) & (!g204)) + ((sk[70]) & (!shiftx6x) & (g199) & (g204)) + ((sk[70]) & (shiftx6x) & (!g199) & (g204)) + ((sk[70]) & (shiftx6x) & (g199) & (g204)));
	assign resultx71x = (((!shiftx6x) & (g210) & (sk[71]) & (!g215)) + ((!shiftx6x) & (g210) & (sk[71]) & (g215)) + ((shiftx6x) & (!g210) & (!sk[71]) & (!g215)) + ((shiftx6x) & (!g210) & (!sk[71]) & (g215)) + ((shiftx6x) & (!g210) & (sk[71]) & (g215)) + ((shiftx6x) & (g210) & (!sk[71]) & (!g215)) + ((shiftx6x) & (g210) & (!sk[71]) & (g215)) + ((shiftx6x) & (g210) & (sk[71]) & (g215)));
	assign resultx72x = (((!shiftx6x) & (sk[72]) & (g221) & (!g226)) + ((!shiftx6x) & (sk[72]) & (g221) & (g226)) + ((shiftx6x) & (!sk[72]) & (!g221) & (!g226)) + ((shiftx6x) & (!sk[72]) & (!g221) & (g226)) + ((shiftx6x) & (!sk[72]) & (g221) & (!g226)) + ((shiftx6x) & (!sk[72]) & (g221) & (g226)) + ((shiftx6x) & (sk[72]) & (!g221) & (g226)) + ((shiftx6x) & (sk[72]) & (g221) & (g226)));
	assign resultx73x = (((!shiftx6x) & (sk[73]) & (g232) & (!g237)) + ((!shiftx6x) & (sk[73]) & (g232) & (g237)) + ((shiftx6x) & (!sk[73]) & (!g232) & (!g237)) + ((shiftx6x) & (!sk[73]) & (!g232) & (g237)) + ((shiftx6x) & (!sk[73]) & (g232) & (!g237)) + ((shiftx6x) & (!sk[73]) & (g232) & (g237)) + ((shiftx6x) & (sk[73]) & (!g232) & (g237)) + ((shiftx6x) & (sk[73]) & (g232) & (g237)));
	assign resultx74x = (((!sk[74]) & (shiftx6x) & (!g243) & (!g248)) + ((!sk[74]) & (shiftx6x) & (!g243) & (g248)) + ((!sk[74]) & (shiftx6x) & (g243) & (!g248)) + ((!sk[74]) & (shiftx6x) & (g243) & (g248)) + ((sk[74]) & (!shiftx6x) & (g243) & (!g248)) + ((sk[74]) & (!shiftx6x) & (g243) & (g248)) + ((sk[74]) & (shiftx6x) & (!g243) & (g248)) + ((sk[74]) & (shiftx6x) & (g243) & (g248)));
	assign resultx75x = (((!shiftx6x) & (g254) & (sk[75]) & (!g259)) + ((!shiftx6x) & (g254) & (sk[75]) & (g259)) + ((shiftx6x) & (!g254) & (!sk[75]) & (!g259)) + ((shiftx6x) & (!g254) & (!sk[75]) & (g259)) + ((shiftx6x) & (!g254) & (sk[75]) & (g259)) + ((shiftx6x) & (g254) & (!sk[75]) & (!g259)) + ((shiftx6x) & (g254) & (!sk[75]) & (g259)) + ((shiftx6x) & (g254) & (sk[75]) & (g259)));
	assign resultx76x = (((!shiftx6x) & (g265) & (sk[76]) & (!g270)) + ((!shiftx6x) & (g265) & (sk[76]) & (g270)) + ((shiftx6x) & (!g265) & (!sk[76]) & (!g270)) + ((shiftx6x) & (!g265) & (!sk[76]) & (g270)) + ((shiftx6x) & (!g265) & (sk[76]) & (g270)) + ((shiftx6x) & (g265) & (!sk[76]) & (!g270)) + ((shiftx6x) & (g265) & (!sk[76]) & (g270)) + ((shiftx6x) & (g265) & (sk[76]) & (g270)));
	assign resultx77x = (((!shiftx6x) & (sk[77]) & (g276) & (!g281)) + ((!shiftx6x) & (sk[77]) & (g276) & (g281)) + ((shiftx6x) & (!sk[77]) & (!g276) & (!g281)) + ((shiftx6x) & (!sk[77]) & (!g276) & (g281)) + ((shiftx6x) & (!sk[77]) & (g276) & (!g281)) + ((shiftx6x) & (!sk[77]) & (g276) & (g281)) + ((shiftx6x) & (sk[77]) & (!g276) & (g281)) + ((shiftx6x) & (sk[77]) & (g276) & (g281)));
	assign resultx78x = (((!sk[78]) & (shiftx6x) & (!g287) & (!g292)) + ((!sk[78]) & (shiftx6x) & (!g287) & (g292)) + ((!sk[78]) & (shiftx6x) & (g287) & (!g292)) + ((!sk[78]) & (shiftx6x) & (g287) & (g292)) + ((sk[78]) & (!shiftx6x) & (g287) & (!g292)) + ((sk[78]) & (!shiftx6x) & (g287) & (g292)) + ((sk[78]) & (shiftx6x) & (!g287) & (g292)) + ((sk[78]) & (shiftx6x) & (g287) & (g292)));
	assign resultx79x = (((!sk[79]) & (shiftx6x) & (!g298) & (!g303)) + ((!sk[79]) & (shiftx6x) & (!g298) & (g303)) + ((!sk[79]) & (shiftx6x) & (g298) & (!g303)) + ((!sk[79]) & (shiftx6x) & (g298) & (g303)) + ((sk[79]) & (!shiftx6x) & (g298) & (!g303)) + ((sk[79]) & (!shiftx6x) & (g298) & (g303)) + ((sk[79]) & (shiftx6x) & (!g298) & (g303)) + ((sk[79]) & (shiftx6x) & (g298) & (g303)));
	assign resultx80x = (((!shiftx6x) & (sk[80]) & (g305) & (!g306)) + ((!shiftx6x) & (sk[80]) & (g305) & (g306)) + ((shiftx6x) & (!sk[80]) & (!g305) & (!g306)) + ((shiftx6x) & (!sk[80]) & (!g305) & (g306)) + ((shiftx6x) & (!sk[80]) & (g305) & (!g306)) + ((shiftx6x) & (!sk[80]) & (g305) & (g306)) + ((shiftx6x) & (sk[80]) & (!g305) & (g306)) + ((shiftx6x) & (sk[80]) & (g305) & (g306)));
	assign resultx81x = (((!shiftx6x) & (g308) & (sk[81]) & (!g309)) + ((!shiftx6x) & (g308) & (sk[81]) & (g309)) + ((shiftx6x) & (!g308) & (!sk[81]) & (!g309)) + ((shiftx6x) & (!g308) & (!sk[81]) & (g309)) + ((shiftx6x) & (!g308) & (sk[81]) & (g309)) + ((shiftx6x) & (g308) & (!sk[81]) & (!g309)) + ((shiftx6x) & (g308) & (!sk[81]) & (g309)) + ((shiftx6x) & (g308) & (sk[81]) & (g309)));
	assign resultx82x = (((!sk[82]) & (shiftx6x) & (!g311) & (!g312)) + ((!sk[82]) & (shiftx6x) & (!g311) & (g312)) + ((!sk[82]) & (shiftx6x) & (g311) & (!g312)) + ((!sk[82]) & (shiftx6x) & (g311) & (g312)) + ((sk[82]) & (!shiftx6x) & (g311) & (!g312)) + ((sk[82]) & (!shiftx6x) & (g311) & (g312)) + ((sk[82]) & (shiftx6x) & (!g311) & (g312)) + ((sk[82]) & (shiftx6x) & (g311) & (g312)));
	assign resultx83x = (((!shiftx6x) & (g314) & (sk[83]) & (!g315)) + ((!shiftx6x) & (g314) & (sk[83]) & (g315)) + ((shiftx6x) & (!g314) & (!sk[83]) & (!g315)) + ((shiftx6x) & (!g314) & (!sk[83]) & (g315)) + ((shiftx6x) & (!g314) & (sk[83]) & (g315)) + ((shiftx6x) & (g314) & (!sk[83]) & (!g315)) + ((shiftx6x) & (g314) & (!sk[83]) & (g315)) + ((shiftx6x) & (g314) & (sk[83]) & (g315)));
	assign resultx84x = (((!shiftx6x) & (g317) & (sk[84]) & (!g318)) + ((!shiftx6x) & (g317) & (sk[84]) & (g318)) + ((shiftx6x) & (!g317) & (!sk[84]) & (!g318)) + ((shiftx6x) & (!g317) & (!sk[84]) & (g318)) + ((shiftx6x) & (!g317) & (sk[84]) & (g318)) + ((shiftx6x) & (g317) & (!sk[84]) & (!g318)) + ((shiftx6x) & (g317) & (!sk[84]) & (g318)) + ((shiftx6x) & (g317) & (sk[84]) & (g318)));
	assign resultx85x = (((!shiftx6x) & (sk[85]) & (g320) & (!g321)) + ((!shiftx6x) & (sk[85]) & (g320) & (g321)) + ((shiftx6x) & (!sk[85]) & (!g320) & (!g321)) + ((shiftx6x) & (!sk[85]) & (!g320) & (g321)) + ((shiftx6x) & (!sk[85]) & (g320) & (!g321)) + ((shiftx6x) & (!sk[85]) & (g320) & (g321)) + ((shiftx6x) & (sk[85]) & (!g320) & (g321)) + ((shiftx6x) & (sk[85]) & (g320) & (g321)));
	assign resultx86x = (((!shiftx6x) & (g323) & (sk[86]) & (!g324)) + ((!shiftx6x) & (g323) & (sk[86]) & (g324)) + ((shiftx6x) & (!g323) & (!sk[86]) & (!g324)) + ((shiftx6x) & (!g323) & (!sk[86]) & (g324)) + ((shiftx6x) & (!g323) & (sk[86]) & (g324)) + ((shiftx6x) & (g323) & (!sk[86]) & (!g324)) + ((shiftx6x) & (g323) & (!sk[86]) & (g324)) + ((shiftx6x) & (g323) & (sk[86]) & (g324)));
	assign resultx87x = (((!shiftx6x) & (sk[87]) & (g326) & (!g327)) + ((!shiftx6x) & (sk[87]) & (g326) & (g327)) + ((shiftx6x) & (!sk[87]) & (!g326) & (!g327)) + ((shiftx6x) & (!sk[87]) & (!g326) & (g327)) + ((shiftx6x) & (!sk[87]) & (g326) & (!g327)) + ((shiftx6x) & (!sk[87]) & (g326) & (g327)) + ((shiftx6x) & (sk[87]) & (!g326) & (g327)) + ((shiftx6x) & (sk[87]) & (g326) & (g327)));
	assign resultx88x = (((!shiftx6x) & (sk[88]) & (g329) & (!g330)) + ((!shiftx6x) & (sk[88]) & (g329) & (g330)) + ((shiftx6x) & (!sk[88]) & (!g329) & (!g330)) + ((shiftx6x) & (!sk[88]) & (!g329) & (g330)) + ((shiftx6x) & (!sk[88]) & (g329) & (!g330)) + ((shiftx6x) & (!sk[88]) & (g329) & (g330)) + ((shiftx6x) & (sk[88]) & (!g329) & (g330)) + ((shiftx6x) & (sk[88]) & (g329) & (g330)));
	assign resultx89x = (((!shiftx6x) & (sk[89]) & (g332) & (!g333)) + ((!shiftx6x) & (sk[89]) & (g332) & (g333)) + ((shiftx6x) & (!sk[89]) & (!g332) & (!g333)) + ((shiftx6x) & (!sk[89]) & (!g332) & (g333)) + ((shiftx6x) & (!sk[89]) & (g332) & (!g333)) + ((shiftx6x) & (!sk[89]) & (g332) & (g333)) + ((shiftx6x) & (sk[89]) & (!g332) & (g333)) + ((shiftx6x) & (sk[89]) & (g332) & (g333)));
	assign resultx90x = (((!shiftx6x) & (g335) & (sk[90]) & (!g336)) + ((!shiftx6x) & (g335) & (sk[90]) & (g336)) + ((shiftx6x) & (!g335) & (!sk[90]) & (!g336)) + ((shiftx6x) & (!g335) & (!sk[90]) & (g336)) + ((shiftx6x) & (!g335) & (sk[90]) & (g336)) + ((shiftx6x) & (g335) & (!sk[90]) & (!g336)) + ((shiftx6x) & (g335) & (!sk[90]) & (g336)) + ((shiftx6x) & (g335) & (sk[90]) & (g336)));
	assign resultx91x = (((!sk[91]) & (shiftx6x) & (!g338) & (!g339)) + ((!sk[91]) & (shiftx6x) & (!g338) & (g339)) + ((!sk[91]) & (shiftx6x) & (g338) & (!g339)) + ((!sk[91]) & (shiftx6x) & (g338) & (g339)) + ((sk[91]) & (!shiftx6x) & (g338) & (!g339)) + ((sk[91]) & (!shiftx6x) & (g338) & (g339)) + ((sk[91]) & (shiftx6x) & (!g338) & (g339)) + ((sk[91]) & (shiftx6x) & (g338) & (g339)));
	assign resultx92x = (((!shiftx6x) & (sk[92]) & (g341) & (!g342)) + ((!shiftx6x) & (sk[92]) & (g341) & (g342)) + ((shiftx6x) & (!sk[92]) & (!g341) & (!g342)) + ((shiftx6x) & (!sk[92]) & (!g341) & (g342)) + ((shiftx6x) & (!sk[92]) & (g341) & (!g342)) + ((shiftx6x) & (!sk[92]) & (g341) & (g342)) + ((shiftx6x) & (sk[92]) & (!g341) & (g342)) + ((shiftx6x) & (sk[92]) & (g341) & (g342)));
	assign resultx93x = (((!shiftx6x) & (sk[93]) & (g344) & (!g345)) + ((!shiftx6x) & (sk[93]) & (g344) & (g345)) + ((shiftx6x) & (!sk[93]) & (!g344) & (!g345)) + ((shiftx6x) & (!sk[93]) & (!g344) & (g345)) + ((shiftx6x) & (!sk[93]) & (g344) & (!g345)) + ((shiftx6x) & (!sk[93]) & (g344) & (g345)) + ((shiftx6x) & (sk[93]) & (!g344) & (g345)) + ((shiftx6x) & (sk[93]) & (g344) & (g345)));
	assign resultx94x = (((!shiftx6x) & (sk[94]) & (g347) & (!g348)) + ((!shiftx6x) & (sk[94]) & (g347) & (g348)) + ((shiftx6x) & (!sk[94]) & (!g347) & (!g348)) + ((shiftx6x) & (!sk[94]) & (!g347) & (g348)) + ((shiftx6x) & (!sk[94]) & (g347) & (!g348)) + ((shiftx6x) & (!sk[94]) & (g347) & (g348)) + ((shiftx6x) & (sk[94]) & (!g347) & (g348)) + ((shiftx6x) & (sk[94]) & (g347) & (g348)));
	assign resultx95x = (((!shiftx6x) & (g350) & (sk[95]) & (!g351)) + ((!shiftx6x) & (g350) & (sk[95]) & (g351)) + ((shiftx6x) & (!g350) & (!sk[95]) & (!g351)) + ((shiftx6x) & (!g350) & (!sk[95]) & (g351)) + ((shiftx6x) & (!g350) & (sk[95]) & (g351)) + ((shiftx6x) & (g350) & (!sk[95]) & (!g351)) + ((shiftx6x) & (g350) & (!sk[95]) & (g351)) + ((shiftx6x) & (g350) & (sk[95]) & (g351)));
	assign resultx96x = (((!shiftx6x) & (g353) & (sk[96]) & (!g354)) + ((!shiftx6x) & (g353) & (sk[96]) & (g354)) + ((shiftx6x) & (!g353) & (!sk[96]) & (!g354)) + ((shiftx6x) & (!g353) & (!sk[96]) & (g354)) + ((shiftx6x) & (!g353) & (sk[96]) & (g354)) + ((shiftx6x) & (g353) & (!sk[96]) & (!g354)) + ((shiftx6x) & (g353) & (!sk[96]) & (g354)) + ((shiftx6x) & (g353) & (sk[96]) & (g354)));
	assign resultx97x = (((!shiftx6x) & (g356) & (sk[97]) & (!g357)) + ((!shiftx6x) & (g356) & (sk[97]) & (g357)) + ((shiftx6x) & (!g356) & (!sk[97]) & (!g357)) + ((shiftx6x) & (!g356) & (!sk[97]) & (g357)) + ((shiftx6x) & (!g356) & (sk[97]) & (g357)) + ((shiftx6x) & (g356) & (!sk[97]) & (!g357)) + ((shiftx6x) & (g356) & (!sk[97]) & (g357)) + ((shiftx6x) & (g356) & (sk[97]) & (g357)));
	assign resultx98x = (((!sk[98]) & (shiftx6x) & (!g359) & (!g360)) + ((!sk[98]) & (shiftx6x) & (!g359) & (g360)) + ((!sk[98]) & (shiftx6x) & (g359) & (!g360)) + ((!sk[98]) & (shiftx6x) & (g359) & (g360)) + ((sk[98]) & (!shiftx6x) & (g359) & (!g360)) + ((sk[98]) & (!shiftx6x) & (g359) & (g360)) + ((sk[98]) & (shiftx6x) & (!g359) & (g360)) + ((sk[98]) & (shiftx6x) & (g359) & (g360)));
	assign resultx99x = (((!shiftx6x) & (sk[99]) & (g362) & (!g363)) + ((!shiftx6x) & (sk[99]) & (g362) & (g363)) + ((shiftx6x) & (!sk[99]) & (!g362) & (!g363)) + ((shiftx6x) & (!sk[99]) & (!g362) & (g363)) + ((shiftx6x) & (!sk[99]) & (g362) & (!g363)) + ((shiftx6x) & (!sk[99]) & (g362) & (g363)) + ((shiftx6x) & (sk[99]) & (!g362) & (g363)) + ((shiftx6x) & (sk[99]) & (g362) & (g363)));
	assign resultx100x = (((!sk[100]) & (shiftx6x) & (!g365) & (!g366)) + ((!sk[100]) & (shiftx6x) & (!g365) & (g366)) + ((!sk[100]) & (shiftx6x) & (g365) & (!g366)) + ((!sk[100]) & (shiftx6x) & (g365) & (g366)) + ((sk[100]) & (!shiftx6x) & (g365) & (!g366)) + ((sk[100]) & (!shiftx6x) & (g365) & (g366)) + ((sk[100]) & (shiftx6x) & (!g365) & (g366)) + ((sk[100]) & (shiftx6x) & (g365) & (g366)));
	assign resultx101x = (((!sk[101]) & (shiftx6x) & (!g368) & (!g369)) + ((!sk[101]) & (shiftx6x) & (!g368) & (g369)) + ((!sk[101]) & (shiftx6x) & (g368) & (!g369)) + ((!sk[101]) & (shiftx6x) & (g368) & (g369)) + ((sk[101]) & (!shiftx6x) & (g368) & (!g369)) + ((sk[101]) & (!shiftx6x) & (g368) & (g369)) + ((sk[101]) & (shiftx6x) & (!g368) & (g369)) + ((sk[101]) & (shiftx6x) & (g368) & (g369)));
	assign resultx102x = (((!sk[102]) & (shiftx6x) & (!g371) & (!g372)) + ((!sk[102]) & (shiftx6x) & (!g371) & (g372)) + ((!sk[102]) & (shiftx6x) & (g371) & (!g372)) + ((!sk[102]) & (shiftx6x) & (g371) & (g372)) + ((sk[102]) & (!shiftx6x) & (g371) & (!g372)) + ((sk[102]) & (!shiftx6x) & (g371) & (g372)) + ((sk[102]) & (shiftx6x) & (!g371) & (g372)) + ((sk[102]) & (shiftx6x) & (g371) & (g372)));
	assign resultx103x = (((!shiftx6x) & (sk[103]) & (g374) & (!g375)) + ((!shiftx6x) & (sk[103]) & (g374) & (g375)) + ((shiftx6x) & (!sk[103]) & (!g374) & (!g375)) + ((shiftx6x) & (!sk[103]) & (!g374) & (g375)) + ((shiftx6x) & (!sk[103]) & (g374) & (!g375)) + ((shiftx6x) & (!sk[103]) & (g374) & (g375)) + ((shiftx6x) & (sk[103]) & (!g374) & (g375)) + ((shiftx6x) & (sk[103]) & (g374) & (g375)));
	assign resultx104x = (((!sk[104]) & (shiftx6x) & (!g377) & (!g378)) + ((!sk[104]) & (shiftx6x) & (!g377) & (g378)) + ((!sk[104]) & (shiftx6x) & (g377) & (!g378)) + ((!sk[104]) & (shiftx6x) & (g377) & (g378)) + ((sk[104]) & (!shiftx6x) & (g377) & (!g378)) + ((sk[104]) & (!shiftx6x) & (g377) & (g378)) + ((sk[104]) & (shiftx6x) & (!g377) & (g378)) + ((sk[104]) & (shiftx6x) & (g377) & (g378)));
	assign resultx105x = (((!shiftx6x) & (sk[105]) & (g380) & (!g381)) + ((!shiftx6x) & (sk[105]) & (g380) & (g381)) + ((shiftx6x) & (!sk[105]) & (!g380) & (!g381)) + ((shiftx6x) & (!sk[105]) & (!g380) & (g381)) + ((shiftx6x) & (!sk[105]) & (g380) & (!g381)) + ((shiftx6x) & (!sk[105]) & (g380) & (g381)) + ((shiftx6x) & (sk[105]) & (!g380) & (g381)) + ((shiftx6x) & (sk[105]) & (g380) & (g381)));
	assign resultx106x = (((!sk[106]) & (shiftx6x) & (!g383) & (!g384)) + ((!sk[106]) & (shiftx6x) & (!g383) & (g384)) + ((!sk[106]) & (shiftx6x) & (g383) & (!g384)) + ((!sk[106]) & (shiftx6x) & (g383) & (g384)) + ((sk[106]) & (!shiftx6x) & (g383) & (!g384)) + ((sk[106]) & (!shiftx6x) & (g383) & (g384)) + ((sk[106]) & (shiftx6x) & (!g383) & (g384)) + ((sk[106]) & (shiftx6x) & (g383) & (g384)));
	assign resultx107x = (((!sk[107]) & (shiftx6x) & (!g386) & (!g387)) + ((!sk[107]) & (shiftx6x) & (!g386) & (g387)) + ((!sk[107]) & (shiftx6x) & (g386) & (!g387)) + ((!sk[107]) & (shiftx6x) & (g386) & (g387)) + ((sk[107]) & (!shiftx6x) & (g386) & (!g387)) + ((sk[107]) & (!shiftx6x) & (g386) & (g387)) + ((sk[107]) & (shiftx6x) & (!g386) & (g387)) + ((sk[107]) & (shiftx6x) & (g386) & (g387)));
	assign resultx108x = (((!shiftx6x) & (g389) & (sk[108]) & (!g390)) + ((!shiftx6x) & (g389) & (sk[108]) & (g390)) + ((shiftx6x) & (!g389) & (!sk[108]) & (!g390)) + ((shiftx6x) & (!g389) & (!sk[108]) & (g390)) + ((shiftx6x) & (!g389) & (sk[108]) & (g390)) + ((shiftx6x) & (g389) & (!sk[108]) & (!g390)) + ((shiftx6x) & (g389) & (!sk[108]) & (g390)) + ((shiftx6x) & (g389) & (sk[108]) & (g390)));
	assign resultx109x = (((!shiftx6x) & (g392) & (sk[109]) & (!g393)) + ((!shiftx6x) & (g392) & (sk[109]) & (g393)) + ((shiftx6x) & (!g392) & (!sk[109]) & (!g393)) + ((shiftx6x) & (!g392) & (!sk[109]) & (g393)) + ((shiftx6x) & (!g392) & (sk[109]) & (g393)) + ((shiftx6x) & (g392) & (!sk[109]) & (!g393)) + ((shiftx6x) & (g392) & (!sk[109]) & (g393)) + ((shiftx6x) & (g392) & (sk[109]) & (g393)));
	assign resultx110x = (((!shiftx6x) & (sk[110]) & (g395) & (!g396)) + ((!shiftx6x) & (sk[110]) & (g395) & (g396)) + ((shiftx6x) & (!sk[110]) & (!g395) & (!g396)) + ((shiftx6x) & (!sk[110]) & (!g395) & (g396)) + ((shiftx6x) & (!sk[110]) & (g395) & (!g396)) + ((shiftx6x) & (!sk[110]) & (g395) & (g396)) + ((shiftx6x) & (sk[110]) & (!g395) & (g396)) + ((shiftx6x) & (sk[110]) & (g395) & (g396)));
	assign resultx111x = (((!shiftx6x) & (sk[111]) & (g398) & (!g399)) + ((!shiftx6x) & (sk[111]) & (g398) & (g399)) + ((shiftx6x) & (!sk[111]) & (!g398) & (!g399)) + ((shiftx6x) & (!sk[111]) & (!g398) & (g399)) + ((shiftx6x) & (!sk[111]) & (g398) & (!g399)) + ((shiftx6x) & (!sk[111]) & (g398) & (g399)) + ((shiftx6x) & (sk[111]) & (!g398) & (g399)) + ((shiftx6x) & (sk[111]) & (g398) & (g399)));
	assign resultx112x = (((!shiftx6x) & (g401) & (sk[112]) & (!g402)) + ((!shiftx6x) & (g401) & (sk[112]) & (g402)) + ((shiftx6x) & (!g401) & (!sk[112]) & (!g402)) + ((shiftx6x) & (!g401) & (!sk[112]) & (g402)) + ((shiftx6x) & (!g401) & (sk[112]) & (g402)) + ((shiftx6x) & (g401) & (!sk[112]) & (!g402)) + ((shiftx6x) & (g401) & (!sk[112]) & (g402)) + ((shiftx6x) & (g401) & (sk[112]) & (g402)));
	assign resultx113x = (((!shiftx6x) & (sk[113]) & (g404) & (!g405)) + ((!shiftx6x) & (sk[113]) & (g404) & (g405)) + ((shiftx6x) & (!sk[113]) & (!g404) & (!g405)) + ((shiftx6x) & (!sk[113]) & (!g404) & (g405)) + ((shiftx6x) & (!sk[113]) & (g404) & (!g405)) + ((shiftx6x) & (!sk[113]) & (g404) & (g405)) + ((shiftx6x) & (sk[113]) & (!g404) & (g405)) + ((shiftx6x) & (sk[113]) & (g404) & (g405)));
	assign resultx114x = (((!shiftx6x) & (sk[114]) & (g407) & (!g408)) + ((!shiftx6x) & (sk[114]) & (g407) & (g408)) + ((shiftx6x) & (!sk[114]) & (!g407) & (!g408)) + ((shiftx6x) & (!sk[114]) & (!g407) & (g408)) + ((shiftx6x) & (!sk[114]) & (g407) & (!g408)) + ((shiftx6x) & (!sk[114]) & (g407) & (g408)) + ((shiftx6x) & (sk[114]) & (!g407) & (g408)) + ((shiftx6x) & (sk[114]) & (g407) & (g408)));
	assign resultx115x = (((!shiftx6x) & (g410) & (sk[115]) & (!g411)) + ((!shiftx6x) & (g410) & (sk[115]) & (g411)) + ((shiftx6x) & (!g410) & (!sk[115]) & (!g411)) + ((shiftx6x) & (!g410) & (!sk[115]) & (g411)) + ((shiftx6x) & (!g410) & (sk[115]) & (g411)) + ((shiftx6x) & (g410) & (!sk[115]) & (!g411)) + ((shiftx6x) & (g410) & (!sk[115]) & (g411)) + ((shiftx6x) & (g410) & (sk[115]) & (g411)));
	assign resultx116x = (((!sk[116]) & (shiftx6x) & (!g413) & (!g414)) + ((!sk[116]) & (shiftx6x) & (!g413) & (g414)) + ((!sk[116]) & (shiftx6x) & (g413) & (!g414)) + ((!sk[116]) & (shiftx6x) & (g413) & (g414)) + ((sk[116]) & (!shiftx6x) & (g413) & (!g414)) + ((sk[116]) & (!shiftx6x) & (g413) & (g414)) + ((sk[116]) & (shiftx6x) & (!g413) & (g414)) + ((sk[116]) & (shiftx6x) & (g413) & (g414)));
	assign resultx117x = (((!shiftx6x) & (sk[117]) & (g416) & (!g417)) + ((!shiftx6x) & (sk[117]) & (g416) & (g417)) + ((shiftx6x) & (!sk[117]) & (!g416) & (!g417)) + ((shiftx6x) & (!sk[117]) & (!g416) & (g417)) + ((shiftx6x) & (!sk[117]) & (g416) & (!g417)) + ((shiftx6x) & (!sk[117]) & (g416) & (g417)) + ((shiftx6x) & (sk[117]) & (!g416) & (g417)) + ((shiftx6x) & (sk[117]) & (g416) & (g417)));
	assign resultx118x = (((!shiftx6x) & (g419) & (sk[118]) & (!g420)) + ((!shiftx6x) & (g419) & (sk[118]) & (g420)) + ((shiftx6x) & (!g419) & (!sk[118]) & (!g420)) + ((shiftx6x) & (!g419) & (!sk[118]) & (g420)) + ((shiftx6x) & (!g419) & (sk[118]) & (g420)) + ((shiftx6x) & (g419) & (!sk[118]) & (!g420)) + ((shiftx6x) & (g419) & (!sk[118]) & (g420)) + ((shiftx6x) & (g419) & (sk[118]) & (g420)));
	assign resultx119x = (((!shiftx6x) & (g422) & (sk[119]) & (!g423)) + ((!shiftx6x) & (g422) & (sk[119]) & (g423)) + ((shiftx6x) & (!g422) & (!sk[119]) & (!g423)) + ((shiftx6x) & (!g422) & (!sk[119]) & (g423)) + ((shiftx6x) & (!g422) & (sk[119]) & (g423)) + ((shiftx6x) & (g422) & (!sk[119]) & (!g423)) + ((shiftx6x) & (g422) & (!sk[119]) & (g423)) + ((shiftx6x) & (g422) & (sk[119]) & (g423)));
	assign resultx120x = (((!shiftx6x) & (sk[120]) & (g425) & (!g426)) + ((!shiftx6x) & (sk[120]) & (g425) & (g426)) + ((shiftx6x) & (!sk[120]) & (!g425) & (!g426)) + ((shiftx6x) & (!sk[120]) & (!g425) & (g426)) + ((shiftx6x) & (!sk[120]) & (g425) & (!g426)) + ((shiftx6x) & (!sk[120]) & (g425) & (g426)) + ((shiftx6x) & (sk[120]) & (!g425) & (g426)) + ((shiftx6x) & (sk[120]) & (g425) & (g426)));
	assign resultx121x = (((!shiftx6x) & (g428) & (sk[121]) & (!g429)) + ((!shiftx6x) & (g428) & (sk[121]) & (g429)) + ((shiftx6x) & (!g428) & (!sk[121]) & (!g429)) + ((shiftx6x) & (!g428) & (!sk[121]) & (g429)) + ((shiftx6x) & (!g428) & (sk[121]) & (g429)) + ((shiftx6x) & (g428) & (!sk[121]) & (!g429)) + ((shiftx6x) & (g428) & (!sk[121]) & (g429)) + ((shiftx6x) & (g428) & (sk[121]) & (g429)));
	assign resultx122x = (((!shiftx6x) & (g431) & (sk[122]) & (!g432)) + ((!shiftx6x) & (g431) & (sk[122]) & (g432)) + ((shiftx6x) & (!g431) & (!sk[122]) & (!g432)) + ((shiftx6x) & (!g431) & (!sk[122]) & (g432)) + ((shiftx6x) & (!g431) & (sk[122]) & (g432)) + ((shiftx6x) & (g431) & (!sk[122]) & (!g432)) + ((shiftx6x) & (g431) & (!sk[122]) & (g432)) + ((shiftx6x) & (g431) & (sk[122]) & (g432)));
	assign resultx123x = (((!shiftx6x) & (g434) & (sk[123]) & (!g435)) + ((!shiftx6x) & (g434) & (sk[123]) & (g435)) + ((shiftx6x) & (!g434) & (!sk[123]) & (!g435)) + ((shiftx6x) & (!g434) & (!sk[123]) & (g435)) + ((shiftx6x) & (!g434) & (sk[123]) & (g435)) + ((shiftx6x) & (g434) & (!sk[123]) & (!g435)) + ((shiftx6x) & (g434) & (!sk[123]) & (g435)) + ((shiftx6x) & (g434) & (sk[123]) & (g435)));
	assign resultx124x = (((!shiftx6x) & (sk[124]) & (g437) & (!g438)) + ((!shiftx6x) & (sk[124]) & (g437) & (g438)) + ((shiftx6x) & (!sk[124]) & (!g437) & (!g438)) + ((shiftx6x) & (!sk[124]) & (!g437) & (g438)) + ((shiftx6x) & (!sk[124]) & (g437) & (!g438)) + ((shiftx6x) & (!sk[124]) & (g437) & (g438)) + ((shiftx6x) & (sk[124]) & (!g437) & (g438)) + ((shiftx6x) & (sk[124]) & (g437) & (g438)));
	assign resultx125x = (((!sk[125]) & (shiftx6x) & (!g440) & (!g441)) + ((!sk[125]) & (shiftx6x) & (!g440) & (g441)) + ((!sk[125]) & (shiftx6x) & (g440) & (!g441)) + ((!sk[125]) & (shiftx6x) & (g440) & (g441)) + ((sk[125]) & (!shiftx6x) & (g440) & (!g441)) + ((sk[125]) & (!shiftx6x) & (g440) & (g441)) + ((sk[125]) & (shiftx6x) & (!g440) & (g441)) + ((sk[125]) & (shiftx6x) & (g440) & (g441)));
	assign resultx126x = (((!sk[126]) & (shiftx6x) & (!g443) & (!g444)) + ((!sk[126]) & (shiftx6x) & (!g443) & (g444)) + ((!sk[126]) & (shiftx6x) & (g443) & (!g444)) + ((!sk[126]) & (shiftx6x) & (g443) & (g444)) + ((sk[126]) & (!shiftx6x) & (g443) & (!g444)) + ((sk[126]) & (!shiftx6x) & (g443) & (g444)) + ((sk[126]) & (shiftx6x) & (!g443) & (g444)) + ((sk[126]) & (shiftx6x) & (g443) & (g444)));
	assign resultx127x = (((!sk[127]) & (shiftx6x) & (!g446) & (!g447)) + ((!sk[127]) & (shiftx6x) & (!g446) & (g447)) + ((!sk[127]) & (shiftx6x) & (g446) & (!g447)) + ((!sk[127]) & (shiftx6x) & (g446) & (g447)) + ((sk[127]) & (!shiftx6x) & (g446) & (!g447)) + ((sk[127]) & (!shiftx6x) & (g446) & (g447)) + ((sk[127]) & (shiftx6x) & (!g446) & (g447)) + ((sk[127]) & (shiftx6x) & (g446) & (g447)));

endmodule