module apex2x6xv (i_30_, i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_27_, i_14_, i_3_, i_28_, i_13_, i_4_, i_25_, i_12_, i_1_, i_26_, i_11_, i_2_, i_23_, i_18_, i_24_, i_17_, i_0_, i_21_, i_16_, i_22_, i_15_, i_32_, i_31_, i_34_, i_33_, i_19_, i_36_, i_35_, i_38_, i_29_, i_37_, o_1_, o_2_, o_0_);

	input i_30_;
	input i_20_;
	input i_9_;
	input i_10_;
	input i_7_;
	input i_8_;
	input i_5_;
	input i_6_;
	input i_27_;
	input i_14_;
	input i_3_;
	input i_28_;
	input i_13_;
	input i_4_;
	input i_25_;
	input i_12_;
	input i_1_;
	input i_26_;
	input i_11_;
	input i_2_;
	input i_23_;
	input i_18_;
	input i_24_;
	input i_17_;
	input i_0_;
	input i_21_;
	input i_16_;
	input i_22_;
	input i_15_;
	input i_32_;
	input i_31_;
	input i_34_;
	input i_33_;
	input i_19_;
	input i_36_;
	input i_35_;
	input i_38_;
	input i_29_;
	input i_37_;
	output o_1_;
	output o_2_;
	output o_0_;

	wire [1347 : 0] sk /* synthesis noprune */;

	lut_sub lut_3 ({sk[0], x7257x, x7252x, x7044x, x7045x, x7248x, x7249x}, o_1_);
	defparam lut_3.LUT_SIZE = 7;
	defparam lut_3.mask = 128'h0f0fffffffffffff7fffffffffffffff;

	lut_sub lut_10 ({sk[1], x7747x, n_n1827, x7486x, x7487x, n_n1811, x7743x}, o_2_);
	defparam lut_10.LUT_SIZE = 7;
	defparam lut_10.mask = 128'h57ffffff57ffffff7fffffffffffffff;

	lut_sub lut_17 ({sk[2], x8080x, x8054x, x8052x, x8053x, x8096x, x8097x}, o_0_);
	defparam lut_17.LUT_SIZE = 7;
	defparam lut_17.mask = 128'h57ffffff57ffffff7fffffffffffffff;

	lut_sub lut_24 ({sk[3], x1757x, x6898x, x1747x, x6919x, x1465x}, x7257x);
	defparam lut_24.LUT_SIZE = 6;
	defparam lut_24.mask = 64'h3f3fffff7fffffff;

	lut_sub lut_30 ({sk[4], n_n1697, n_n1690, n_n1687, x7238x, x7239x}, x7252x);
	defparam lut_30.LUT_SIZE = 6;
	defparam lut_30.mask = 64'h3f3fffff7fffffff;

	lut_sub lut_36 ({sk[5], n_n1718, n_n1719, n_n1720, x7043x}, x7044x);
	defparam lut_36.LUT_SIZE = 5;
	defparam lut_36.mask = 32'h77777fff;

	lut_sub lut_41 ({sk[6], n_n1716, n_n1715, x7022x, n_n1723}, x7045x);
	defparam lut_41.LUT_SIZE = 5;
	defparam lut_41.mask = 32'h77777fff;

	lut_sub lut_46 ({sk[7], x7111x, n_n1713, n_n1712, x1587x, x7110x}, x7248x);
	defparam lut_46.LUT_SIZE = 6;
	defparam lut_46.mask = 64'h3f3fffff7fffffff;

	lut_sub lut_52 ({sk[8], x6933x, x6934x, x6942x, x6943x, x1597x, x7104x}, x7249x);
	defparam lut_52.LUT_SIZE = 7;
	defparam lut_52.mask = 128'h57ffffff57ffffff7fffffffffffffff;

	lut_sub lut_59 ({sk[9], x7349x, n_n1829, n_n1820, x7441x, n_n1824, x7348x}, x7747x);
	defparam lut_59.LUT_SIZE = 7;
	defparam lut_59.mask = 128'h57ffffff57ffffff7fffffffffffffff;

	lut_sub lut_66 ({sk[10], n_n1862, x7370x, x7371x, x7381x, x7382x}, n_n1827);
	defparam lut_66.LUT_SIZE = 6;
	defparam lut_66.mask = 64'h3f3fffff7fffffff;

	lut_sub lut_72 ({sk[11], i_31_, n_n1850, x651x, x7452x, x1240x, x7483x}, x7486x);
	defparam lut_72.LUT_SIZE = 7;
	defparam lut_72.mask = 128'h57ffffff57ffffff7fffffff7f7fffff;

	lut_sub lut_78 ({sk[12], n_n1847, n_n1846, n_n1848, x7463x, n_n1844, x7477x}, x7487x);
	defparam lut_78.LUT_SIZE = 7;
	defparam lut_78.mask = 128'h57ffffff57ffffff7fffffffffffffff;

	lut_sub lut_85 ({sk[13], n_n1834, x7598x, x7711x, x7712x, x9194x}, n_n1811);
	defparam lut_85.LUT_SIZE = 6;
	defparam lut_85.mask = 64'h3f3fffffbfffffff;

	lut_sub lut_91 ({sk[14], x7719x, x7720x, n_n1865, x7740x, x7741x}, x7743x);
	defparam lut_91.LUT_SIZE = 6;
	defparam lut_91.mask = 64'h3f3fffff7fffffff;

	lut_sub lut_97 ({sk[15], n_n1549, x7882x, x7883x, n_n1556, x7922x, x8078x}, x8080x);
	defparam lut_97.LUT_SIZE = 7;
	defparam lut_97.mask = 128'h57ffffff57ffffff7fffffffffffffff;

	lut_sub lut_104 ({sk[16], n_n1574, n_n1575, n_n1577, x8037x, x8038x}, x8054x);
	defparam lut_104.LUT_SIZE = 6;
	defparam lut_104.mask = 64'h3f3fffff7fffffff;

	lut_sub lut_110 ({sk[17], i_21_, x8025x, x8026x, x8048x, x730x}, x8052x);
	defparam lut_110.LUT_SIZE = 6;
	defparam lut_110.mask = 64'h3f3fffff3fff7fff;

	lut_sub lut_115 ({sk[18], n_n1578, n_n1576, x8016x, x8017x}, x8053x);
	defparam lut_115.LUT_SIZE = 5;
	defparam lut_115.mask = 32'h77777fff;

	lut_sub lut_120 ({sk[19], i_17_, x7781x, x43x, x569x, x8093x, x8094x}, x8096x);
	defparam lut_120.LUT_SIZE = 7;
	defparam lut_120.mask = 128'h57ffffff57ffffff777fffff7777ffff;

	lut_sub lut_125 ({sk[20], i_36_, x7760x, x7771x, x548x, x566x}, x8097x);
	defparam lut_125.LUT_SIZE = 6;
	defparam lut_125.mask = 64'h3f3fffff0fff7fff;

	lut_sub lut_130 ({sk[21], x10x, n_n1318, x604x, x1761x, x1762x, x6889x}, x1757x);
	defparam lut_130.LUT_SIZE = 7;
	defparam lut_130.mask = 128'h57ffffff57ffffff0000005500003f7f;

	lut_sub lut_134 ({sk[22], x19x, x1765x, x1766x, x492x, x1755x, x6884x}, x6898x);
	defparam lut_134.LUT_SIZE = 7;
	defparam lut_134.mask = 128'h57ffffff57ffffff337777773f7f7f7f;

	lut_sub lut_139 ({sk[23], n_n26, x1753x, x1754x, x6912x, x1749x, x1750x}, x1747x);
	defparam lut_139.LUT_SIZE = 7;
	defparam lut_139.mask = 128'h57ffffff57ffffff00000000777f7f7f;

	lut_sub lut_144 ({sk[24], x1743x, x1744x, x1745x, x1746x}, x6919x);
	defparam lut_144.LUT_SIZE = 5;
	defparam lut_144.mask = 32'h77777fff;

	lut_sub lut_149 ({sk[25], i_9_, i_13_, x59x, x1470x, x1471x, x1472x}, x1465x);
	defparam lut_149.LUT_SIZE = 7;
	defparam lut_149.mask = 128'h57ffffff57ffffff007f000f000f000f;

	lut_sub lut_153 ({sk[26], x1457x, x7267x, n_n1856, x1392x, x7339x, x7290x}, x7349x);
	defparam lut_153.LUT_SIZE = 7;
	defparam lut_153.mask = 128'h57ffffff57ffffff7fffffffffffffff;

	lut_sub lut_160 ({sk[27], i_38_, x1347x, x7396x, n_n1870, x627x, x7406x}, n_n1829);
	defparam lut_160.LUT_SIZE = 7;
	defparam lut_160.mask = 128'h57ffffff57ffffff5fffffff7fffffff;

	lut_sub lut_166 ({sk[28], x1318x, x7422x, n_n1843, x7434x}, n_n1820);
	defparam lut_166.LUT_SIZE = 5;
	defparam lut_166.mask = 32'h77777fff;

	lut_sub lut_171 ({sk[29], n_n1839, x1296x, x7439x}, x7441x);
	defparam lut_171.LUT_SIZE = 4;
	defparam lut_171.mask = 16'h557f;

	lut_sub lut_175 ({sk[30], i_31_, x42x, x7313x, x7315x, x623x, x1408x}, n_n1824);
	defparam lut_175.LUT_SIZE = 7;
	defparam lut_175.mask = 128'h57ffffff57ffffff5fff7fff5fff5fff;

	lut_sub lut_180 ({sk[31], i_32_, x7327x, x7346x, x7347x, x611x}, x7348x);
	defparam lut_180.LUT_SIZE = 6;
	defparam lut_180.mask = 64'h3f3fffff7fff3fff;

	lut_sub lut_185 ({sk[32], i_14_, i_16_}, x10x);
	defparam lut_185.LUT_SIZE = 3;
	defparam lut_185.mask = 8'h38;

	lut_sub lut_187 ({sk[33], i_35_, i_37_}, n_n1318);
	defparam lut_187.LUT_SIZE = 3;
	defparam lut_187.mask = 8'h34;

	lut_sub lut_189 ({sk[34], i_5_, i_3_, i_4_, i_0_, x361x, x353x}, x604x);
	defparam lut_189.LUT_SIZE = 7;
	defparam lut_189.mask = 128'h57ffffff57ffffff3000700000005000;

	lut_sub lut_192 ({sk[35], i_20_, i_18_, i_17_, x46x, n_n26, x6891x}, x1761x);
	defparam lut_192.LUT_SIZE = 7;
	defparam lut_192.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_194 ({sk[36], i_20_, i_11_, i_17_, i_19_, x46x, x487x}, x1762x);
	defparam lut_194.LUT_SIZE = 7;
	defparam lut_194.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_196 ({sk[37], i_28_, i_17_, i_32_, i_29_, x10x, x6886x}, x6889x);
	defparam lut_196.LUT_SIZE = 7;
	defparam lut_196.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_198 ({sk[38], n_n1278, n_n787, n_n180, x14x, n_n179, x326x}, x19x);
	defparam lut_198.LUT_SIZE = 7;
	defparam lut_198.mask = 128'h57ffffff57ffffff0505050505050537;

	lut_sub lut_201 ({sk[39], i_9_, i_13_, i_11_, i_19_, x263x, x376x}, x1765x);
	defparam lut_201.LUT_SIZE = 7;
	defparam lut_201.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_203 ({sk[40], i_8_, i_13_, i_18_, n_n1278, x263x, x404x}, x1766x);
	defparam lut_203.LUT_SIZE = 7;
	defparam lut_203.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_205 ({sk[41], i_32_, i_34_, i_33_, i_35_, i_37_, n_n1375}, x492x);
	defparam lut_205.LUT_SIZE = 7;
	defparam lut_205.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_207 ({sk[42], i_20_, x263x, n_n245, x46x, x6876x, x6879x}, x1755x);
	defparam lut_207.LUT_SIZE = 7;
	defparam lut_207.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_209 ({sk[43], i_34_, i_33_, i_35_, i_29_, i_37_, n_n793}, x6884x);
	defparam lut_209.LUT_SIZE = 7;
	defparam lut_209.mask = 128'h57ffffff57ffffff0010000000000000;

	lut_sub lut_211 ({sk[44], i_3_, i_4_, i_0_}, n_n26);
	defparam lut_211.LUT_SIZE = 4;
	defparam lut_211.mask = 16'h5508;

	lut_sub lut_213 ({sk[45], i_20_, i_14_, i_29_, n_n1441, x54x, x413x}, x1753x);
	defparam lut_213.LUT_SIZE = 7;
	defparam lut_213.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_215 ({sk[46], i_20_, i_18_, i_17_, i_32_, x10x, x46x}, x1754x);
	defparam lut_215.LUT_SIZE = 7;
	defparam lut_215.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_217 ({sk[47], i_9_, i_7_, i_5_, i_6_, i_37_}, x6912x);
	defparam lut_217.LUT_SIZE = 6;
	defparam lut_217.mask = 64'h3f3fffff40000000;

	lut_sub lut_219 ({sk[48], i_20_, n_n180, x46x, x6890x, x1751x, x1752x}, x1749x);
	defparam lut_219.LUT_SIZE = 7;
	defparam lut_219.mask = 128'h57ffffff57ffffff0000000700000000;

	lut_sub lut_222 ({sk[49], i_28_, i_32_, i_29_, x6886x, x461x, x353x}, x1750x);
	defparam lut_222.LUT_SIZE = 7;
	defparam lut_222.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_224 ({sk[50], n_n1303, n_n245, x431x, x44x, x6899x, x6900x}, x1743x);
	defparam lut_224.LUT_SIZE = 7;
	defparam lut_224.mask = 128'h57ffffff57ffffff0000000000000001;

	lut_sub lut_226 ({sk[51], i_20_, n_n504, x46x, n_n178, x6893x, x487x}, x1744x);
	defparam lut_226.LUT_SIZE = 7;
	defparam lut_226.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_228 ({sk[52], n_n1443, n_n504, n_n245, n_n460, x6886x, x361x}, x1745x);
	defparam lut_228.LUT_SIZE = 7;
	defparam lut_228.mask = 128'h57ffffff57ffffff0000000000000001;

	lut_sub lut_230 ({sk[53], i_20_, n_n245, x46x, x6893x, x6908x, x6906x}, x1746x);
	defparam lut_230.LUT_SIZE = 7;
	defparam lut_230.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_232 ({sk[54], i_5_, i_4_, i_0_, x636x, x7133x}, n_n1697);
	defparam lut_232.LUT_SIZE = 6;
	defparam lut_232.mask = 64'h3f3fffff75555555;

	lut_sub lut_235 ({sk[55], i_37_, x7062x, x1619x, x7077x, x768x, x7093x}, n_n1690);
	defparam lut_235.LUT_SIZE = 7;
	defparam lut_235.mask = 128'h57ffffff57ffffff5fffffff7fffffff;

	lut_sub lut_241 ({sk[56], x1501x, x7207x, x7221x, x7222x, x7233x, x7234x}, n_n1687);
	defparam lut_241.LUT_SIZE = 7;
	defparam lut_241.mask = 128'h57ffffff57ffffff7fffffffffffffff;

	lut_sub lut_248 ({sk[57], i_33_, i_37_, x685x, x7157x, x7192x, x7193x}, x7238x);
	defparam lut_248.LUT_SIZE = 7;
	defparam lut_248.mask = 128'h57ffffff57ffffff7f7f7fff7f7f7f7f;

	lut_sub lut_253 ({sk[58], x7142x, x7143x, x1536x, x7172x, x1525x, x7184x}, x7239x);
	defparam lut_253.LUT_SIZE = 7;
	defparam lut_253.mask = 128'h57ffffff57ffffff7fffffffffffffff;

	lut_sub lut_260 ({sk[59], i_33_, i_37_}, x59x);
	defparam lut_260.LUT_SIZE = 3;
	defparam lut_260.mask = 8'h34;

	lut_sub lut_262 ({sk[60], i_5_, i_4_, i_0_}, n_n245);
	defparam lut_262.LUT_SIZE = 4;
	defparam lut_262.mask = 16'h5580;

	lut_sub lut_264 ({sk[61], i_27_, i_28_, i_26_, i_23_, i_24_, i_29_}, x46x);
	defparam lut_264.LUT_SIZE = 7;
	defparam lut_264.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_266 ({sk[62], i_13_, i_11_, i_16_}, n_n178);
	defparam lut_266.LUT_SIZE = 4;
	defparam lut_266.mask = 16'h5580;

	lut_sub lut_268 ({sk[63], i_17_, i_19_}, x6893x);
	defparam lut_268.LUT_SIZE = 3;
	defparam lut_268.mask = 8'h38;

	lut_sub lut_270 ({sk[64], i_9_, i_7_, i_6_, i_32_}, x6906x);
	defparam lut_270.LUT_SIZE = 5;
	defparam lut_270.mask = 32'h77778000;

	lut_sub lut_272 ({sk[65], i_20_, n_n245, x46x, n_n178, x6893x, x6906x}, x1470x);
	defparam lut_272.LUT_SIZE = 7;
	defparam lut_272.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_274 ({sk[66], i_28_, i_22_, i_38_, n_n1454, x1462x, x581x}, x1457x);
	defparam lut_274.LUT_SIZE = 7;
	defparam lut_274.mask = 128'h57ffffff57ffffff0037003300330033;

	lut_sub lut_277 ({sk[67], i_9_, x204x, n_n416, x70x, x376x, x1456x}, x7267x);
	defparam lut_277.LUT_SIZE = 7;
	defparam lut_277.mask = 128'h57ffffff57ffffff555f575f555f555f;

	lut_sub lut_281 ({sk[68], i_24_, x801x, x1447x, x1448x, x7275x, x1450x}, n_n1856);
	defparam lut_281.LUT_SIZE = 7;
	defparam lut_281.mask = 128'h57ffffff57ffffff5fff7fff5fff5fff;

	lut_sub lut_286 ({sk[69], i_24_, i_32_, x42x, n_n416, x800x, x7332x}, x1392x);
	defparam lut_286.LUT_SIZE = 7;
	defparam lut_286.mask = 128'h57ffffff57ffffff0015000500000000;

	lut_sub lut_289 ({sk[70], x1393x, x1394x, x1395x, x1396x, x7335x}, x7339x);
	defparam lut_289.LUT_SIZE = 6;
	defparam lut_289.mask = 64'h3f3fffff7fffffff;

	lut_sub lut_295 ({sk[71], i_9_, x204x, x376x, x1437x, x7286x, x1439x}, x7290x);
	defparam lut_295.LUT_SIZE = 7;
	defparam lut_295.mask = 128'h57ffffff57ffffff5f5f5f7f5f5f5f5f;

	lut_sub lut_299 ({sk[72], x1372x, x1373x, x1374x, x1375x, x1376x, x1377x}, n_n1862);
	defparam lut_299.LUT_SIZE = 7;
	defparam lut_299.mask = 128'h57ffffff57ffffff7fffffffffffffff;

	lut_sub lut_306 ({sk[73], i_32_, i_31_, x53x, x218x, x1370x, x1371x}, x7370x);
	defparam lut_306.LUT_SIZE = 7;
	defparam lut_306.mask = 128'h57ffffff57ffffff777f777777777777;

	lut_sub lut_310 ({sk[74], x243x, x311x, x26x, x1366x, x1369x, x7366x}, x7371x);
	defparam lut_310.LUT_SIZE = 7;
	defparam lut_310.mask = 128'h57ffffff57ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_315 ({sk[75], x223x, n_n1133, x218x, x315x, x387x, x1353x}, x7381x);
	defparam lut_315.LUT_SIZE = 7;
	defparam lut_315.mask = 128'h57ffffff57ffffff5555555f7777777f;

	lut_sub lut_319 ({sk[76], i_22_, x73x, x7287x, x625x, x1355x, x1358x}, x7382x);
	defparam lut_319.LUT_SIZE = 7;
	defparam lut_319.mask = 128'h57ffffff57ffffff7777777f77777777;

	lut_sub lut_323 ({sk[77], i_33_, i_35_, i_38_, x1352x, x1350x, x7392x}, x1347x);
	defparam lut_323.LUT_SIZE = 7;
	defparam lut_323.mask = 128'h57ffffff57ffffff007f000000000000;

	lut_sub lut_327 ({sk[78], i_24_, n_n1353, x11x, x7386x, x1348x, x7394x}, x7396x);
	defparam lut_327.LUT_SIZE = 7;
	defparam lut_327.mask = 128'h57ffffff57ffffff7777777f77777777;

	lut_sub lut_331 ({sk[79], i_13_, x15x, x388x, x1335x, x1334x, x1337x}, n_n1870);
	defparam lut_331.LUT_SIZE = 7;
	defparam lut_331.mask = 128'h57ffffff57ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_336 ({sk[80], i_9_, i_10_, i_13_, x52x, x376x, x1330x}, x627x);
	defparam lut_336.LUT_SIZE = 7;
	defparam lut_336.mask = 128'h57ffffff57ffffff5757555755555555;

	lut_sub lut_340 ({sk[81], i_13_, i_24_, i_38_, x85x, x78x, x1325x}, x7406x);
	defparam lut_340.LUT_SIZE = 7;
	defparam lut_340.mask = 128'h57ffffff57ffffff5555555555575555;

	lut_sub lut_343 ({sk[82], i_28_, i_33_, n_n1361, n_n1523, x1320x, x7421x}, x1318x);
	defparam lut_343.LUT_SIZE = 7;
	defparam lut_343.mask = 128'h57ffffff57ffffff0007000000000000;

	lut_sub lut_346 ({sk[83], i_35_, i_38_, x476x, n_n338, x28x, x752x}, x7422x);
	defparam lut_346.LUT_SIZE = 7;
	defparam lut_346.mask = 128'h57ffffff57ffffff0303035703030303;

	lut_sub lut_349 ({sk[84], i_32_, x53x, x253x, x755x, x754x, x1316x}, n_n1843);
	defparam lut_349.LUT_SIZE = 7;
	defparam lut_349.mask = 128'h57ffffff57ffffff55775f7f55775577;

	lut_sub lut_353 ({sk[85], n_n300, x654x, x1308x, x1309x, x1311x}, x7434x);
	defparam lut_353.LUT_SIZE = 6;
	defparam lut_353.mask = 64'h3f3fffff7f7f7fff;

	lut_sub lut_358 ({sk[86], n_n300, x53x, x675x, x674x, x1305x}, n_n1839);
	defparam lut_358.LUT_SIZE = 6;
	defparam lut_358.mask = 64'h3f3fffff55775f7f;

	lut_sub lut_362 ({sk[87], i_19_, x12x, x21x, x28x, x78x, x7438x}, x1296x);
	defparam lut_362.LUT_SIZE = 7;
	defparam lut_362.mask = 128'h57ffffff57ffffff0000003300001333;

	lut_sub lut_366 ({sk[88], i_32_, x208x, x53x, x7427x, x656x}, x7439x);
	defparam lut_366.LUT_SIZE = 6;
	defparam lut_366.mask = 64'h3f3fffff05070003;

	lut_sub lut_369 ({sk[89], x24x, x381x, x1293x, x7442x, x7443x, x1292x}, n_n1850);
	defparam lut_369.LUT_SIZE = 7;
	defparam lut_369.mask = 128'h57ffffff57ffffff577757775777ffff;

	lut_sub lut_374 ({sk[90], i_28_, i_25_, i_29_, n_n805, x30x, x1288x}, x651x);
	defparam lut_374.LUT_SIZE = 7;
	defparam lut_374.mask = 128'h57ffffff57ffffff5755555555555555;

	lut_sub lut_377 ({sk[91], x204x, n_n416, x15x, x387x, x1284x, x1285x}, x7452x);
	defparam lut_377.LUT_SIZE = 7;
	defparam lut_377.mask = 128'h57ffffff57ffffff77777f7f777f7f7f;

	lut_sub lut_382 ({sk[92], i_25_, x204x, x42x, n_n416, x15x, n_n1419}, x1240x);
	defparam lut_382.LUT_SIZE = 7;
	defparam lut_382.mask = 128'h57ffffff57ffffff0005001500000000;

	lut_sub lut_385 ({sk[93], n_n1288, x14x, x1238x, x7480x, x1241x, x1242x}, x7483x);
	defparam lut_385.LUT_SIZE = 7;
	defparam lut_385.mask = 128'h57ffffff57ffffff77ff77ff77ff7fff;

	lut_sub lut_390 ({sk[94], x11x, x7423x, x253x, x24x, x1281x, x1283x}, n_n1847);
	defparam lut_390.LUT_SIZE = 7;
	defparam lut_390.mask = 128'h57ffffff57ffffff777f777f777f77ff;

	lut_sub lut_395 ({sk[95], n_n1486, x28x, x371x, x1265x, x1266x, x1267x}, n_n1846);
	defparam lut_395.LUT_SIZE = 7;
	defparam lut_395.mask = 128'h57ffffff57ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_400 ({sk[96], x20x, x381x, x1277x, x671x, x7456x, x1275x}, n_n1848);
	defparam lut_400.LUT_SIZE = 7;
	defparam lut_400.mask = 128'h57ffffff57ffffff55775f7f77777f7f;

	lut_sub lut_405 ({sk[97], n_n1497, x7444x, x676x, x1268x, x1270x, x1271x}, x7463x);
	defparam lut_405.LUT_SIZE = 7;
	defparam lut_405.mask = 128'h57ffffff57ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_410 ({sk[98], x12x, x21x, x7431x, x1256x, x1257x, x1259x}, n_n1844);
	defparam lut_410.LUT_SIZE = 7;
	defparam lut_410.mask = 128'h57ffffff57ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_415 ({sk[99], i_35_, i_38_, x476x, x677x, x1247x, x1249x}, x7477x);
	defparam lut_415.LUT_SIZE = 7;
	defparam lut_415.mask = 128'h57ffffff57ffffff7777777f77777777;

	lut_sub lut_419 ({sk[100], i_9_, i_12_, n_n1884, x760x, x7669x, x7680x}, n_n1834);
	defparam lut_419.LUT_SIZE = 7;
	defparam lut_419.mask = 128'h57ffffff57ffffff77ff77ff77ff7fff;

	lut_sub lut_424 ({sk[101], i_25_, x42x, n_n1871, x700x, x7529x, n_n1873}, x7598x);
	defparam lut_424.LUT_SIZE = 7;
	defparam lut_424.mask = 128'h57ffffff57ffffff77ff7fff77ff77ff;

	lut_sub lut_429 ({sk[102], n_n1881, n_n1882, n_n1880}, x7711x);
	defparam lut_429.LUT_SIZE = 4;
	defparam lut_429.mask = 16'h557f;

	lut_sub lut_433 ({sk[103], n_n1889, x7622x, n_n1837, n_n1887, x7709x, x7642x}, x7712x);
	defparam lut_433.LUT_SIZE = 7;
	defparam lut_433.mask = 128'h57ffffff57ffffff7fffffffffffffff;

	lut_sub lut_440 ({sk[104], n_n1875, n_n1876, n_n1877, n_n1878, x7570x, x7595x}, x9194x);
	defparam lut_440.LUT_SIZE = 7;
	defparam lut_440.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_442 ({sk[105], i_11_, i_19_}, x204x);
	defparam lut_442.LUT_SIZE = 3;
	defparam lut_442.mask = 8'h38;

	lut_sub lut_444 ({sk[106], i_7_, i_8_, i_5_, i_6_, i_18_, x404x}, n_n416);
	defparam lut_444.LUT_SIZE = 7;
	defparam lut_444.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_446 ({sk[107], i_9_, i_5_, i_6_, i_4_, i_2_, x13x}, x15x);
	defparam lut_446.LUT_SIZE = 7;
	defparam lut_446.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_448 ({sk[108], i_28_, i_24_, i_31_, i_33_, i_29_, n_n805}, x66x);
	defparam lut_448.LUT_SIZE = 7;
	defparam lut_448.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_450 ({sk[109], i_10_, i_13_, i_32_, n_n1307, x41x, n_n839}, x750x);
	defparam lut_450.LUT_SIZE = 7;
	defparam lut_450.mask = 128'h57ffffff57ffffff3733373305003733;

	lut_sub lut_454 ({sk[110], i_28_, i_26_, i_24_, i_33_, i_38_, i_29_}, x7715x);
	defparam lut_454.LUT_SIZE = 7;
	defparam lut_454.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_456 ({sk[111], x204x, n_n416, x15x, x66x, x750x, x7715x}, x7719x);
	defparam lut_456.LUT_SIZE = 7;
	defparam lut_456.mask = 128'h57ffffff57ffffff0303575703575757;

	lut_sub lut_460 ({sk[112], i_34_, i_35_, i_38_}, n_n805);
	defparam lut_460.LUT_SIZE = 4;
	defparam lut_460.mask = 16'h5504;

	lut_sub lut_462 ({sk[113], i_28_, i_26_, i_33_, i_38_, i_29_}, x380x);
	defparam lut_462.LUT_SIZE = 6;
	defparam lut_462.mask = 64'h3f3fffff20000000;

	lut_sub lut_464 ({sk[114], i_9_, i_18_, x204x, n_n1278, n_n787, x14x}, x800x);
	defparam lut_464.LUT_SIZE = 7;
	defparam lut_464.mask = 128'h57ffffff57ffffff0357005500550055;

	lut_sub lut_467 ({sk[115], i_8_, i_24_, x230x, x11x, n_n1302, x7717x}, x749x);
	defparam lut_467.LUT_SIZE = 7;
	defparam lut_467.mask = 128'h57ffffff57ffffff0007000000050000;

	lut_sub lut_470 ({sk[116], i_24_, i_32_, n_n805, x380x, x800x, x749x}, x7720x);
	defparam lut_470.LUT_SIZE = 7;
	defparam lut_470.mask = 128'h57ffffff57ffffff0357005500550055;

	lut_sub lut_473 ({sk[117], i_10_, i_28_, i_24_, n_n805, n_n1305, x229x}, x982x);
	defparam lut_473.LUT_SIZE = 7;
	defparam lut_473.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_475 ({sk[118], i_9_, i_22_, n_n1497, x343x, x764x, x7724x}, x983x);
	defparam lut_475.LUT_SIZE = 7;
	defparam lut_475.mask = 128'h57ffffff57ffffff0005000000150011;

	lut_sub lut_478 ({sk[119], i_28_, i_25_, i_24_, n_n805, n_n1133, x207x}, x984x);
	defparam lut_478.LUT_SIZE = 7;
	defparam lut_478.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_480 ({sk[120], i_9_, i_10_, i_28_, i_32_, x11x, x389x}, x985x);
	defparam lut_480.LUT_SIZE = 7;
	defparam lut_480.mask = 128'h57ffffff57ffffff0000000010000000;

	lut_sub lut_482 ({sk[121], i_10_, i_35_, i_38_, x42x, x14x, n_n1311}, x986x);
	defparam lut_482.LUT_SIZE = 7;
	defparam lut_482.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_484 ({sk[122], i_9_, i_10_, i_8_, i_24_, x11x, x271x}, x987x);
	defparam lut_484.LUT_SIZE = 7;
	defparam lut_484.mask = 128'h57ffffff57ffffff0000000010000000;

	lut_sub lut_486 ({sk[123], x982x, x983x, x984x, x985x, x986x, x987x}, n_n1865);
	defparam lut_486.LUT_SIZE = 7;
	defparam lut_486.mask = 128'h57ffffff57ffffff7fffffffffffffff;

	lut_sub lut_493 ({sk[124], i_10_, n_n1486, x50x, x229x, n_n1359, x7736x}, x791x);
	defparam lut_493.LUT_SIZE = 7;
	defparam lut_493.mask = 128'h57ffffff57ffffff0505053700000033;

	lut_sub lut_496 ({sk[125], i_10_, i_13_, i_31_, x41x, x71x, x12x}, x976x);
	defparam lut_496.LUT_SIZE = 7;
	defparam lut_496.mask = 128'h57ffffff57ffffff0100010000000100;

	lut_sub lut_499 ({sk[126], i_33_, i_35_, i_38_, x791x, x976x}, x7740x);
	defparam lut_499.LUT_SIZE = 6;
	defparam lut_499.mask = 64'h3f3fffff57555555;

	lut_sub lut_502 ({sk[127], i_9_, i_10_, i_5_, i_6_, i_4_, i_2_}, x207x);
	defparam lut_502.LUT_SIZE = 7;
	defparam lut_502.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_504 ({sk[128], i_10_, i_24_, i_32_, n_n1361, x229x, x71x}, x971x);
	defparam lut_504.LUT_SIZE = 7;
	defparam lut_504.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_506 ({sk[129], i_28_, i_31_, i_29_, n_n1307, n_n839, x270x}, x974x);
	defparam lut_506.LUT_SIZE = 7;
	defparam lut_506.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_508 ({sk[130], n_n805, x11x, x50x, n_n1359, x344x, x7732x}, x7737x);
	defparam lut_508.LUT_SIZE = 7;
	defparam lut_508.mask = 128'h57ffffff57ffffff0005000500050307;

	lut_sub lut_511 ({sk[131], i_32_, x207x, x66x, x971x, x974x, x7737x}, x7741x);
	defparam lut_511.LUT_SIZE = 7;
	defparam lut_511.mask = 128'h57ffffff57ffffff7f7f7fff7f7f7f7f;

	lut_sub lut_516 ({sk[132], i_27_, i_28_, i_26_, i_24_, i_29_}, x45x);
	defparam lut_516.LUT_SIZE = 6;
	defparam lut_516.mask = 64'h3f3fffff40000000;

	lut_sub lut_518 ({sk[133], i_13_, i_23_, i_17_, i_21_, i_16_}, x7752x);
	defparam lut_518.LUT_SIZE = 6;
	defparam lut_518.mask = 64'h3f3fffff80000000;

	lut_sub lut_520 ({sk[134], i_9_, i_8_, i_6_, x204x, n_n461, x338x}, x547x);
	defparam lut_520.LUT_SIZE = 7;
	defparam lut_520.mask = 128'h57ffffff57ffffff5703000000000000;

	lut_sub lut_523 ({sk[135], i_21_, x232x, x54x, x549x, x44x, x7750x}, x960x);
	defparam lut_523.LUT_SIZE = 7;
	defparam lut_523.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_525 ({sk[136], i_36_, i_35_, x45x, x7752x, x547x, x960x}, x7760x);
	defparam lut_525.LUT_SIZE = 7;
	defparam lut_525.mask = 128'h57ffffff57ffffff5555555555575555;

	lut_sub lut_528 ({sk[137], i_9_, i_8_, i_5_, i_6_, i_4_, i_2_}, x41x);
	defparam lut_528.LUT_SIZE = 7;
	defparam lut_528.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_530 ({sk[138], i_34_, i_36_, i_35_, i_29_, n_n1216}, x396x);
	defparam lut_530.LUT_SIZE = 6;
	defparam lut_530.mask = 64'h3f3fffff00000040;

	lut_sub lut_532 ({sk[139], i_23_, i_18_, i_17_, n_n787, n_n1118, n_n180}, x498x);
	defparam lut_532.LUT_SIZE = 7;
	defparam lut_532.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_534 ({sk[140], i_13_, i_11_, i_23_, i_17_, i_16_, i_19_}, x326x);
	defparam lut_534.LUT_SIZE = 7;
	defparam lut_534.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_536 ({sk[141], i_9_, i_13_, n_n461, x10x, x45x, x7762x}, x952x);
	defparam lut_536.LUT_SIZE = 7;
	defparam lut_536.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_538 ({sk[142], i_21_, x232x, x54x, x420x, x7769x, x44x}, x955x);
	defparam lut_538.LUT_SIZE = 7;
	defparam lut_538.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_540 ({sk[143], x41x, x396x, x498x, x326x, x952x, x955x}, x7771x);
	defparam lut_540.LUT_SIZE = 7;
	defparam lut_540.mask = 128'h57ffffff57ffffff777777ff77777fff;

	lut_sub lut_545 ({sk[144], i_9_, i_5_, i_6_, i_4_}, x232x);
	defparam lut_545.LUT_SIZE = 5;
	defparam lut_545.mask = 32'h77778000;

	lut_sub lut_547 ({sk[145], i_28_, i_29_}, x42x);
	defparam lut_547.LUT_SIZE = 3;
	defparam lut_547.mask = 8'h38;

	lut_sub lut_549 ({sk[146], i_27_, i_26_, i_24_, i_36_, i_35_}, x368x);
	defparam lut_549.LUT_SIZE = 6;
	defparam lut_549.mask = 64'h3f3fffff20000000;

	lut_sub lut_551 ({sk[147], n_n787, n_n1118, n_n180, n_n179, x41x, x326x}, x570x);
	defparam lut_551.LUT_SIZE = 7;
	defparam lut_551.mask = 128'h57ffffff57ffffff111111111111111f;

	lut_sub lut_554 ({sk[148], n_n301, x46x, n_n576, x45x, x7762x, x7776x}, x568x);
	defparam lut_554.LUT_SIZE = 7;
	defparam lut_554.mask = 128'h57ffffff57ffffff0000005503030357;

	lut_sub lut_557 ({sk[149], i_21_, x232x, x54x, x571x, x44x, x7772x}, x942x);
	defparam lut_557.LUT_SIZE = 7;
	defparam lut_557.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_559 ({sk[150], x232x, x42x, x368x, x570x, x568x, x942x}, x7781x);
	defparam lut_559.LUT_SIZE = 7;
	defparam lut_559.mask = 128'h57ffffff57ffffff5555555f7777777f;

	lut_sub lut_563 ({sk[151], x7825x, x7826x, x7839x, x7840x, x7852x}, n_n1549);
	defparam lut_563.LUT_SIZE = 6;
	defparam lut_563.mask = 64'h3f3fffff7fffffff;

	lut_sub lut_569 ({sk[152], i_27_, i_28_, i_31_, x47x, x542x, x7881x}, x7882x);
	defparam lut_569.LUT_SIZE = 7;
	defparam lut_569.mask = 128'h57ffffff57ffffff5557555555555555;

	lut_sub lut_572 ({sk[153], i_36_, x877x, x7866x, x7876x, x563x, x863x}, x7883x);
	defparam lut_572.LUT_SIZE = 7;
	defparam lut_572.mask = 128'h57ffffff57ffffff5fffffff7fffffff;

	lut_sub lut_578 ({sk[154], n_n1443, n_n1429, n_n1585, x1662x, x308x, x7938x}, n_n1556);
	defparam lut_578.LUT_SIZE = 7;
	defparam lut_578.mask = 128'h57ffffff57ffffff5fff7fff7fff7fff;

	lut_sub lut_584 ({sk[155], x843x, x7895x, x834x, x7909x, x7919x, x7920x}, x7922x);
	defparam lut_584.LUT_SIZE = 7;
	defparam lut_584.mask = 128'h57ffffff57ffffff7fffffffffffffff;

	lut_sub lut_591 ({sk[156], n_n1580, n_n1579, n_n1581, n_n1583, n_n1582, n_n1584}, x8078x);
	defparam lut_591.LUT_SIZE = 7;
	defparam lut_591.mask = 128'h57ffffff57ffffff7fffffffffffffff;

	lut_sub lut_598 ({sk[157], i_7_, i_5_, i_6_}, n_n1278);
	defparam lut_598.LUT_SIZE = 4;
	defparam lut_598.mask = 16'h5580;

	lut_sub lut_600 ({sk[158], i_3_, i_4_, i_2_}, n_n787);
	defparam lut_600.LUT_SIZE = 4;
	defparam lut_600.mask = 16'h5508;

	lut_sub lut_602 ({sk[159], i_9_, i_13_, i_16_}, n_n180);
	defparam lut_602.LUT_SIZE = 4;
	defparam lut_602.mask = 16'h5580;

	lut_sub lut_604 ({sk[160], i_9_, i_7_, i_5_, i_6_, i_4_, i_2_}, x14x);
	defparam lut_604.LUT_SIZE = 7;
	defparam lut_604.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_606 ({sk[161], i_23_, i_18_, i_17_}, n_n179);
	defparam lut_606.LUT_SIZE = 4;
	defparam lut_606.mask = 16'h5580;

	lut_sub lut_608 ({sk[162], i_17_, i_16_}, x263x);
	defparam lut_608.LUT_SIZE = 3;
	defparam lut_608.mask = 8'h38;

	lut_sub lut_610 ({sk[163], i_7_, i_8_, i_5_, i_6_, i_4_, i_2_}, x376x);
	defparam lut_610.LUT_SIZE = 7;
	defparam lut_610.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_612 ({sk[164], i_9_, i_3_, i_4_, i_2_}, x404x);
	defparam lut_612.LUT_SIZE = 5;
	defparam lut_612.mask = 32'h77770800;

	lut_sub lut_614 ({sk[165], i_5_, i_6_, i_4_}, n_n461);
	defparam lut_614.LUT_SIZE = 4;
	defparam lut_614.mask = 16'h5580;

	lut_sub lut_616 ({sk[166], i_27_, i_28_, i_23_}, n_n793);
	defparam lut_616.LUT_SIZE = 4;
	defparam lut_616.mask = 16'h5580;

	lut_sub lut_618 ({sk[167], i_27_, i_26_, i_24_, i_36_}, x79x);
	defparam lut_618.LUT_SIZE = 5;
	defparam lut_618.mask = 32'h77774000;

	lut_sub lut_620 ({sk[168], i_27_, i_28_, i_29_}, n_n1375);
	defparam lut_620.LUT_SIZE = 4;
	defparam lut_620.mask = 16'h5580;

	lut_sub lut_622 ({sk[169], i_32_, i_34_, i_36_, i_35_}, x227x);
	defparam lut_622.LUT_SIZE = 5;
	defparam lut_622.mask = 32'h77771000;

	lut_sub lut_624 ({sk[170], i_5_, i_3_, i_4_, i_18_}, x338x);
	defparam lut_624.LUT_SIZE = 5;
	defparam lut_624.mask = 32'h77770800;

	lut_sub lut_626 ({sk[171], i_7_, i_8_, i_13_, i_11_, i_16_, i_19_}, x8087x);
	defparam lut_626.LUT_SIZE = 7;
	defparam lut_626.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_628 ({sk[172], i_9_, i_7_, i_8_, i_6_, i_13_, i_16_}, x8088x);
	defparam lut_628.LUT_SIZE = 7;
	defparam lut_628.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_630 ({sk[173], i_17_, i_36_}, x8089x);
	defparam lut_630.LUT_SIZE = 3;
	defparam lut_630.mask = 8'h34;

	lut_sub lut_632 ({sk[174], x232x, x46x, x338x, x8087x, x8088x, x8089x}, x101x);
	defparam lut_632.LUT_SIZE = 7;
	defparam lut_632.mask = 128'h57ffffff57ffffff0000001100000515;

	lut_sub lut_635 ({sk[175], i_13_, i_17_, i_16_}, n_n1443);
	defparam lut_635.LUT_SIZE = 4;
	defparam lut_635.mask = 16'h5580;

	lut_sub lut_637 ({sk[176], i_9_, i_7_, i_6_}, n_n1100);
	defparam lut_637.LUT_SIZE = 4;
	defparam lut_637.mask = 16'h5580;

	lut_sub lut_639 ({sk[177], i_28_, i_32_, i_29_}, n_n460);
	defparam lut_639.LUT_SIZE = 4;
	defparam lut_639.mask = 16'h5540;

	lut_sub lut_641 ({sk[178], i_23_, x79x, n_n1443, n_n1100, n_n460, x338x}, x102x);
	defparam lut_641.LUT_SIZE = 7;
	defparam lut_641.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_643 ({sk[179], i_28_, i_26_}, x58x);
	defparam lut_643.LUT_SIZE = 3;
	defparam lut_643.mask = 8'h38;

	lut_sub lut_645 ({sk[180], i_27_, i_28_, i_26_}, n_n1441);
	defparam lut_645.LUT_SIZE = 4;
	defparam lut_645.mask = 16'h5580;

	lut_sub lut_647 ({sk[181], i_13_, i_16_}, x43x);
	defparam lut_647.LUT_SIZE = 3;
	defparam lut_647.mask = 8'h38;

	lut_sub lut_649 ({sk[182], i_32_, i_31_}, x302x);
	defparam lut_649.LUT_SIZE = 3;
	defparam lut_649.mask = 8'h38;

	lut_sub lut_651 ({sk[183], i_23_, i_24_}, x54x);
	defparam lut_651.LUT_SIZE = 3;
	defparam lut_651.mask = 8'h38;

	lut_sub lut_653 ({sk[184], i_25_, i_23_, i_24_}, n_n1396);
	defparam lut_653.LUT_SIZE = 4;
	defparam lut_653.mask = 16'h5508;

	lut_sub lut_655 ({sk[185], i_14_, i_12_, i_16_}, n_n1404);
	defparam lut_655.LUT_SIZE = 4;
	defparam lut_655.mask = 16'h5580;

	lut_sub lut_657 ({sk[186], i_23_, i_24_, i_16_}, n_n1390);
	defparam lut_657.LUT_SIZE = 4;
	defparam lut_657.mask = 16'h5580;

	lut_sub lut_659 ({sk[187], i_14_, i_12_}, x415x);
	defparam lut_659.LUT_SIZE = 3;
	defparam lut_659.mask = 8'h38;

	lut_sub lut_661 ({sk[188], i_26_, i_24_}, x73x);
	defparam lut_661.LUT_SIZE = 3;
	defparam lut_661.mask = 8'h38;

	lut_sub lut_663 ({sk[189], i_27_, i_26_, i_24_}, n_n1369);
	defparam lut_663.LUT_SIZE = 4;
	defparam lut_663.mask = 16'h5580;

	lut_sub lut_665 ({sk[190], i_13_, i_12_, i_16_}, n_n1429);
	defparam lut_665.LUT_SIZE = 4;
	defparam lut_665.mask = 16'h5580;

	lut_sub lut_667 ({sk[191], i_25_, i_26_, i_24_}, n_n1454);
	defparam lut_667.LUT_SIZE = 4;
	defparam lut_667.mask = 16'h5580;

	lut_sub lut_669 ({sk[192], i_30_, i_28_, i_29_}, n_n1489);
	defparam lut_669.LUT_SIZE = 4;
	defparam lut_669.mask = 16'h5580;

	lut_sub lut_671 ({sk[193], i_9_, i_10_}, x230x);
	defparam lut_671.LUT_SIZE = 3;
	defparam lut_671.mask = 8'h32;

	lut_sub lut_673 ({sk[194], i_9_, i_10_, i_8_}, n_n1353);
	defparam lut_673.LUT_SIZE = 4;
	defparam lut_673.mask = 16'h5508;

	lut_sub lut_675 ({sk[195], i_35_, i_38_}, n_n1361);
	defparam lut_675.LUT_SIZE = 3;
	defparam lut_675.mask = 8'h34;

	lut_sub lut_677 ({sk[196], i_30_, i_32_}, x3x);
	defparam lut_677.LUT_SIZE = 3;
	defparam lut_677.mask = 8'h37;

	lut_sub lut_680 ({sk[197], i_30_, i_32_, i_31_}, n_n1438);
	defparam lut_680.LUT_SIZE = 4;
	defparam lut_680.mask = 16'h5580;

	lut_sub lut_682 ({sk[198], i_34_, i_35_}, n_n1397);
	defparam lut_682.LUT_SIZE = 3;
	defparam lut_682.mask = 8'h34;

	lut_sub lut_684 ({sk[199], i_23_, i_17_}, x242x);
	defparam lut_684.LUT_SIZE = 3;
	defparam lut_684.mask = 8'h38;

	lut_sub lut_686 ({sk[200], i_20_, i_23_, i_17_}, n_n1274);
	defparam lut_686.LUT_SIZE = 4;
	defparam lut_686.mask = 16'h5580;

	lut_sub lut_688 ({sk[201], i_31_, i_34_}, n_n1334);
	defparam lut_688.LUT_SIZE = 3;
	defparam lut_688.mask = 8'h31;

	lut_sub lut_690 ({sk[202], i_28_, i_29_}, n_n1368);
	defparam lut_690.LUT_SIZE = 3;
	defparam lut_690.mask = 8'h34;

	lut_sub lut_692 ({sk[203], i_27_, i_28_, i_24_}, n_n1216);
	defparam lut_692.LUT_SIZE = 4;
	defparam lut_692.mask = 16'h5580;

	lut_sub lut_694 ({sk[204], i_4_, i_2_}, x292x);
	defparam lut_694.LUT_SIZE = 3;
	defparam lut_694.mask = 8'h38;

	lut_sub lut_696 ({sk[205], i_5_, i_4_, i_2_}, n_n1307);
	defparam lut_696.LUT_SIZE = 4;
	defparam lut_696.mask = 16'h5580;

	lut_sub lut_698 ({sk[206], i_34_, i_33_}, n_n1374);
	defparam lut_698.LUT_SIZE = 3;
	defparam lut_698.mask = 8'h31;

	lut_sub lut_700 ({sk[207], i_31_, i_34_, i_35_}, n_n1504);
	defparam lut_700.LUT_SIZE = 4;
	defparam lut_700.mask = 16'h5504;

	lut_sub lut_702 ({sk[208], i_9_, i_10_, i_6_}, n_n853);
	defparam lut_702.LUT_SIZE = 4;
	defparam lut_702.mask = 16'h5580;

	lut_sub lut_704 ({sk[209], i_20_, i_23_, i_21_}, n_n1092);
	defparam lut_704.LUT_SIZE = 4;
	defparam lut_704.mask = 16'h5508;

	lut_sub lut_706 ({sk[210], i_27_, i_28_, i_29_}, n_n1406);
	defparam lut_706.LUT_SIZE = 4;
	defparam lut_706.mask = 16'h5540;

	lut_sub lut_708 ({sk[211], i_33_, i_35_, i_38_}, n_n1197);
	defparam lut_708.LUT_SIZE = 4;
	defparam lut_708.mask = 16'h5540;

	lut_sub lut_710 ({sk[212], i_30_, i_32_, i_33_, i_35_, i_38_}, n_n762);
	defparam lut_710.LUT_SIZE = 6;
	defparam lut_710.mask = 64'h3f3fffff40000000;

	lut_sub lut_712 ({sk[213], i_9_, i_8_, i_3_}, n_n1038);
	defparam lut_712.LUT_SIZE = 4;
	defparam lut_712.mask = 16'h5508;

	lut_sub lut_714 ({sk[214], i_13_, i_23_, i_16_}, n_n1314);
	defparam lut_714.LUT_SIZE = 4;
	defparam lut_714.mask = 16'h5580;

	lut_sub lut_716 ({sk[215], i_7_, i_8_}, x13x);
	defparam lut_716.LUT_SIZE = 3;
	defparam lut_716.mask = 8'h38;

	lut_sub lut_718 ({sk[216], i_7_, i_8_, i_12_}, n_n1141);
	defparam lut_718.LUT_SIZE = 4;
	defparam lut_718.mask = 16'h5580;

	lut_sub lut_720 ({sk[217], i_5_, i_6_, i_4_, i_12_, i_2_}, x11x);
	defparam lut_720.LUT_SIZE = 6;
	defparam lut_720.mask = 64'h3f3fffff80000000;

	lut_sub lut_722 ({sk[218], i_28_, i_26_, i_29_}, n_n1486);
	defparam lut_722.LUT_SIZE = 4;
	defparam lut_722.mask = 16'h5580;

	lut_sub lut_724 ({sk[219], i_14_, i_17_, i_16_}, n_n1408);
	defparam lut_724.LUT_SIZE = 4;
	defparam lut_724.mask = 16'h5580;

	lut_sub lut_726 ({sk[220], i_33_, i_35_, i_37_}, n_n504);
	defparam lut_726.LUT_SIZE = 4;
	defparam lut_726.mask = 16'h5540;

	lut_sub lut_728 ({sk[221], i_32_, i_29_}, x243x);
	defparam lut_728.LUT_SIZE = 3;
	defparam lut_728.mask = 8'h38;

	lut_sub lut_730 ({sk[222], i_32_, i_33_, i_29_}, n_n1305);
	defparam lut_730.LUT_SIZE = 4;
	defparam lut_730.mask = 16'h5580;

	lut_sub lut_732 ({sk[223], i_8_, i_5_, i_6_}, n_n1118);
	defparam lut_732.LUT_SIZE = 4;
	defparam lut_732.mask = 16'h5580;

	lut_sub lut_734 ({sk[224], i_7_, i_5_, i_6_, i_4_, i_1_, i_2_}, x49x);
	defparam lut_734.LUT_SIZE = 7;
	defparam lut_734.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_736 ({sk[225], i_9_, i_13_}, x279x);
	defparam lut_736.LUT_SIZE = 3;
	defparam lut_736.mask = 8'h32;

	lut_sub lut_738 ({sk[226], i_9_, i_13_, i_18_}, n_n1048);
	defparam lut_738.LUT_SIZE = 4;
	defparam lut_738.mask = 16'h5504;

	lut_sub lut_740 ({sk[227], i_8_, i_5_, i_6_, i_4_, i_12_, i_2_}, x76x);
	defparam lut_740.LUT_SIZE = 7;
	defparam lut_740.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_742 ({sk[228], i_14_, i_23_, i_16_}, n_n1263);
	defparam lut_742.LUT_SIZE = 4;
	defparam lut_742.mask = 16'h5580;

	lut_sub lut_744 ({sk[229], i_7_, i_6_, i_12_}, n_n1306);
	defparam lut_744.LUT_SIZE = 4;
	defparam lut_744.mask = 16'h5580;

	lut_sub lut_746 ({sk[230], i_7_, i_5_, i_6_, i_4_, i_12_, i_2_}, x321x);
	defparam lut_746.LUT_SIZE = 7;
	defparam lut_746.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_748 ({sk[231], i_7_, i_6_, i_12_, i_23_, x10x, n_n1307}, n_n620);
	defparam lut_748.LUT_SIZE = 7;
	defparam lut_748.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_750 ({sk[232], i_28_, i_32_, i_29_}, n_n1288);
	defparam lut_750.LUT_SIZE = 4;
	defparam lut_750.mask = 16'h5580;

	lut_sub lut_752 ({sk[233], i_3_, i_13_, i_4_, i_12_, i_2_}, x213x);
	defparam lut_752.LUT_SIZE = 6;
	defparam lut_752.mask = 64'h3f3fffff80000000;

	lut_sub lut_754 ({sk[234], i_9_, i_5_, i_6_, i_11_}, x7425x);
	defparam lut_754.LUT_SIZE = 5;
	defparam lut_754.mask = 32'h77770040;

	lut_sub lut_756 ({sk[235], i_9_, i_13_, i_11_, i_18_}, x7426x);
	defparam lut_756.LUT_SIZE = 5;
	defparam lut_756.mask = 32'h77770010;

	lut_sub lut_758 ({sk[236], i_9_, i_13_, i_11_}, n_n1055);
	defparam lut_758.LUT_SIZE = 4;
	defparam lut_758.mask = 16'h5504;

	lut_sub lut_760 ({sk[237], i_5_, i_6_, i_3_, i_4_, i_1_, i_2_}, x208x);
	defparam lut_760.LUT_SIZE = 7;
	defparam lut_760.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_762 ({sk[238], i_32_, i_35_, i_38_}, n_n1179);
	defparam lut_762.LUT_SIZE = 4;
	defparam lut_762.mask = 16'h5540;

	lut_sub lut_764 ({sk[239], i_24_, i_22_}, x205x);
	defparam lut_764.LUT_SIZE = 3;
	defparam lut_764.mask = 8'h38;

	lut_sub lut_766 ({sk[240], i_28_, i_25_, i_26_, i_24_, i_22_}, x257x);
	defparam lut_766.LUT_SIZE = 6;
	defparam lut_766.mask = 64'h3f3fffff80000000;

	lut_sub lut_768 ({sk[241], i_25_, i_24_, i_22_, i_32_, x58x, n_n1361}, n_n300);
	defparam lut_768.LUT_SIZE = 7;
	defparam lut_768.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_770 ({sk[242], i_28_, i_34_, i_29_}, n_n1225);
	defparam lut_770.LUT_SIZE = 4;
	defparam lut_770.mask = 16'h5520;

	lut_sub lut_772 ({sk[243], i_10_, i_13_, i_16_}, n_n301);
	defparam lut_772.LUT_SIZE = 4;
	defparam lut_772.mask = 16'h5580;

	lut_sub lut_774 ({sk[244], i_5_, i_6_, i_4_, i_1_, i_2_}, x51x);
	defparam lut_774.LUT_SIZE = 6;
	defparam lut_774.mask = 64'h3f3fffff80000000;

	lut_sub lut_776 ({sk[245], i_23_, i_17_, i_16_}, n_n1322);
	defparam lut_776.LUT_SIZE = 4;
	defparam lut_776.mask = 16'h5580;

	lut_sub lut_778 ({sk[246], i_14_, i_23_, i_17_, i_16_}, x260x);
	defparam lut_778.LUT_SIZE = 5;
	defparam lut_778.mask = 32'h77778000;

	lut_sub lut_780 ({sk[247], i_27_, i_23_, i_17_}, n_n1258);
	defparam lut_780.LUT_SIZE = 4;
	defparam lut_780.mask = 16'h5580;

	lut_sub lut_782 ({sk[248], i_34_, i_33_, i_35_}, n_n1437);
	defparam lut_782.LUT_SIZE = 4;
	defparam lut_782.mask = 16'h5508;

	lut_sub lut_784 ({sk[249], i_32_, i_34_, i_33_}, n_n1340);
	defparam lut_784.LUT_SIZE = 4;
	defparam lut_784.mask = 16'h5520;

	lut_sub lut_786 ({sk[250], i_4_, i_1_, i_0_}, n_n152);
	defparam lut_786.LUT_SIZE = 4;
	defparam lut_786.mask = 16'h5580;

	lut_sub lut_788 ({sk[251], i_33_, i_38_}, n_n1300);
	defparam lut_788.LUT_SIZE = 3;
	defparam lut_788.mask = 8'h34;

	lut_sub lut_790 ({sk[252], i_8_, i_5_, i_6_, i_4_, i_1_, i_2_}, x50x);
	defparam lut_790.LUT_SIZE = 7;
	defparam lut_790.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_792 ({sk[253], i_28_, i_25_, i_26_, i_24_, i_22_}, x52x);
	defparam lut_792.LUT_SIZE = 6;
	defparam lut_792.mask = 64'h3f3fffff80000000;

	lut_sub lut_794 ({sk[254], i_9_, i_7_, i_6_, i_32_, n_n1307}, x85x);
	defparam lut_794.LUT_SIZE = 6;
	defparam lut_794.mask = 64'h3f3fffff40000000;

	lut_sub lut_796 ({sk[255], i_9_, i_10_, i_7_, i_8_, i_6_, n_n1307}, x223x);
	defparam lut_796.LUT_SIZE = 7;
	defparam lut_796.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_798 ({sk[256], i_28_, i_24_, i_34_, i_33_, i_35_, i_38_}, x237x);
	defparam lut_798.LUT_SIZE = 7;
	defparam lut_798.mask = 128'h57ffffff57ffffff0040000000000000;

	lut_sub lut_800 ({sk[257], i_31_, i_35_, i_38_}, x264x);
	defparam lut_800.LUT_SIZE = 4;
	defparam lut_800.mask = 16'h5540;

	lut_sub lut_802 ({sk[258], i_28_, i_26_, i_24_, i_22_}, x61x);
	defparam lut_802.LUT_SIZE = 5;
	defparam lut_802.mask = 32'h77778000;

	lut_sub lut_804 ({sk[259], i_28_, i_26_, i_24_, i_22_, i_33_, i_38_}, x388x);
	defparam lut_804.LUT_SIZE = 7;
	defparam lut_804.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_806 ({sk[260], i_32_, i_31_, i_35_, i_38_}, x446x);
	defparam lut_806.LUT_SIZE = 5;
	defparam lut_806.mask = 32'h77774000;

	lut_sub lut_808 ({sk[261], i_10_, i_24_, i_22_}, n_n1191);
	defparam lut_808.LUT_SIZE = 4;
	defparam lut_808.mask = 16'h5580;

	lut_sub lut_810 ({sk[262], i_10_, i_28_, i_26_, i_24_, i_22_}, x518x);
	defparam lut_810.LUT_SIZE = 6;
	defparam lut_810.mask = 64'h3f3fffff80000000;

	lut_sub lut_812 ({sk[263], i_9_, i_3_, i_13_, i_11_}, x262x);
	defparam lut_812.LUT_SIZE = 5;
	defparam lut_812.mask = 32'h77770040;

	lut_sub lut_814 ({sk[264], i_9_, i_3_, i_13_, i_11_, i_18_, i_19_}, x529x);
	defparam lut_814.LUT_SIZE = 7;
	defparam lut_814.mask = 128'h57ffffff57ffffff000000005f001300;

	lut_sub lut_819 ({sk[265], i_30_, i_32_, i_29_, x237x, x529x}, x1215x);
	defparam lut_819.LUT_SIZE = 6;
	defparam lut_819.mask = 64'h3f3fffff10000000;

	lut_sub lut_821 ({sk[266], i_32_, i_33_, i_38_, x58x, x14x, n_n1191}, x1216x);
	defparam lut_821.LUT_SIZE = 7;
	defparam lut_821.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_823 ({sk[267], i_32_, i_31_, i_35_, i_38_, x51x, x52x}, x1217x);
	defparam lut_823.LUT_SIZE = 7;
	defparam lut_823.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_825 ({sk[268], i_9_, i_13_, i_24_, n_n1307, n_n1303, x7509x}, x1218x);
	defparam lut_825.LUT_SIZE = 7;
	defparam lut_825.mask = 128'h57ffffff57ffffff0000010000000000;

	lut_sub lut_827 ({sk[269], i_31_, i_35_, i_38_, x257x, x50x}, x1219x);
	defparam lut_827.LUT_SIZE = 6;
	defparam lut_827.mask = 64'h3f3fffff01000000;

	lut_sub lut_829 ({sk[270], i_9_, i_10_, i_33_, i_38_, x61x, x376x}, x1220x);
	defparam lut_829.LUT_SIZE = 7;
	defparam lut_829.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_831 ({sk[271], x1215x, x1216x, x1217x, x1218x, x1219x, x1220x}, n_n1871);
	defparam lut_831.LUT_SIZE = 7;
	defparam lut_831.mask = 128'h57ffffff57ffffff7fffffffffffffff;

	lut_sub lut_838 ({sk[272], i_7_, i_13_, i_12_}, n_n1147);
	defparam lut_838.LUT_SIZE = 4;
	defparam lut_838.mask = 16'h5580;

	lut_sub lut_840 ({sk[273], i_7_, i_14_, i_12_}, n_n1089);
	defparam lut_840.LUT_SIZE = 4;
	defparam lut_840.mask = 16'h5580;

	lut_sub lut_842 ({sk[274], i_24_, i_34_}, x298x);
	defparam lut_842.LUT_SIZE = 3;
	defparam lut_842.mask = 8'h34;

	lut_sub lut_844 ({sk[275], i_27_, i_28_, i_26_, i_36_}, x7791x);
	defparam lut_844.LUT_SIZE = 5;
	defparam lut_844.mask = 32'h77774000;

	lut_sub lut_846 ({sk[276], i_30_, i_23_, i_24_, i_16_, i_32_, i_29_}, x7792x);
	defparam lut_846.LUT_SIZE = 7;
	defparam lut_846.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_848 ({sk[277], i_30_, i_34_, i_36_, i_29_}, x7784x);
	defparam lut_848.LUT_SIZE = 5;
	defparam lut_848.mask = 32'h77770200;

	lut_sub lut_850 ({sk[278], i_27_, i_28_, i_23_, i_24_, i_17_, i_29_}, x48x);
	defparam lut_850.LUT_SIZE = 7;
	defparam lut_850.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_852 ({sk[279], i_30_, i_7_, i_32_, i_34_, i_36_}, x7790x);
	defparam lut_852.LUT_SIZE = 6;
	defparam lut_852.mask = 64'h3f3fffff10000000;

	lut_sub lut_854 ({sk[280], i_30_, i_32_, i_34_, i_36_}, x7787x);
	defparam lut_854.LUT_SIZE = 5;
	defparam lut_854.mask = 32'h77771000;

	lut_sub lut_856 ({sk[281], i_27_, i_28_, i_23_, i_24_, i_16_, i_29_}, x7788x);
	defparam lut_856.LUT_SIZE = 7;
	defparam lut_856.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_858 ({sk[282], i_27_, i_28_, i_26_, i_23_, i_24_, i_17_}, x74x);
	defparam lut_858.LUT_SIZE = 7;
	defparam lut_858.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_860 ({sk[283], i_30_, i_7_, i_32_, i_36_, i_29_}, x7786x);
	defparam lut_860.LUT_SIZE = 6;
	defparam lut_860.mask = 64'h3f3fffff20000000;

	lut_sub lut_862 ({sk[284], i_7_, i_8_, i_14_, i_12_, i_23_, i_16_}, x324x);
	defparam lut_862.LUT_SIZE = 7;
	defparam lut_862.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_864 ({sk[285], i_30_, i_28_, i_29_, x13x, x260x, x324x}, x531x);
	defparam lut_864.LUT_SIZE = 7;
	defparam lut_864.mask = 128'h57ffffff57ffffff5700000000000000;

	lut_sub lut_867 ({sk[286], i_7_, i_8_, i_13_, i_12_, i_23_, i_16_}, x323x);
	defparam lut_867.LUT_SIZE = 7;
	defparam lut_867.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_869 ({sk[287], i_7_, i_8_, i_13_, i_23_, i_17_, i_16_}, x291x);
	defparam lut_869.LUT_SIZE = 7;
	defparam lut_869.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_871 ({sk[288], n_n1216, x7784x, x323x, x291x, x7782x, x7783x}, x7793x);
	defparam lut_871.LUT_SIZE = 7;
	defparam lut_871.mask = 128'h57ffffff57ffffff1111111111111fff;

	lut_sub lut_875 ({sk[289], x10x, n_n1147, x7787x, x7788x, x74x, x7786x}, x7794x);
	defparam lut_875.LUT_SIZE = 7;
	defparam lut_875.mask = 128'h57ffffff57ffffff0000000f1111111f;

	lut_sub lut_878 ({sk[290], x43x, n_n1089, x7791x, x7792x, x48x, x7790x}, x7795x);
	defparam lut_878.LUT_SIZE = 7;
	defparam lut_878.mask = 128'h57ffffff57ffffff0000000f1111111f;

	lut_sub lut_881 ({sk[291], i_36_, n_n1369, x531x, x7793x, x7794x, x7795x}, n_n1580);
	defparam lut_881.LUT_SIZE = 7;
	defparam lut_881.mask = 128'h57ffffff57ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_886 ({sk[292], i_28_, i_34_, i_29_}, n_n1326);
	defparam lut_886.LUT_SIZE = 4;
	defparam lut_886.mask = 16'h5540;

	lut_sub lut_888 ({sk[293], i_27_, i_28_, i_24_, i_34_, i_29_}, x7804x);
	defparam lut_888.LUT_SIZE = 6;
	defparam lut_888.mask = 64'h3f3fffff10000000;

	lut_sub lut_890 ({sk[294], i_23_, i_24_, i_21_, i_34_}, x245x);
	defparam lut_890.LUT_SIZE = 5;
	defparam lut_890.mask = 32'h77771000;

	lut_sub lut_892 ({sk[295], i_30_, i_28_}, x277x);
	defparam lut_892.LUT_SIZE = 3;
	defparam lut_892.mask = 8'h38;

	lut_sub lut_894 ({sk[296], i_28_, i_31_, i_34_}, n_n1511);
	defparam lut_894.LUT_SIZE = 4;
	defparam lut_894.mask = 16'h5510;

	lut_sub lut_896 ({sk[297], i_27_, i_23_, i_24_, i_21_}, x7802x);
	defparam lut_896.LUT_SIZE = 5;
	defparam lut_896.mask = 32'h77774000;

	lut_sub lut_898 ({sk[298], i_32_, i_31_, i_33_}, n_n1393);
	defparam lut_898.LUT_SIZE = 4;
	defparam lut_898.mask = 16'h5540;

	lut_sub lut_900 ({sk[299], i_14_, i_32_, i_31_, i_33_}, x340x);
	defparam lut_900.LUT_SIZE = 5;
	defparam lut_900.mask = 32'h77770040;

	lut_sub lut_902 ({sk[300], i_20_, i_26_, i_2_, i_21_, x54x, n_n1406}, x432x);
	defparam lut_902.LUT_SIZE = 7;
	defparam lut_902.mask = 128'h57ffffff57ffffff0010000000000000;

	lut_sub lut_904 ({sk[301], i_13_, i_12_, i_17_, i_16_}, x533x);
	defparam lut_904.LUT_SIZE = 5;
	defparam lut_904.mask = 32'h7777a800;

	lut_sub lut_907 ({sk[302], i_9_, i_7_, i_13_, i_12_, i_17_, i_16_}, x532x);
	defparam lut_907.LUT_SIZE = 7;
	defparam lut_907.mask = 128'h57ffffff57ffffff0000a80000000000;

	lut_sub lut_910 ({sk[303], n_n1438, n_n1216, x7784x, n_n1326, x7798x, x7800x}, x7805x);
	defparam lut_910.LUT_SIZE = 7;
	defparam lut_910.mask = 128'h57ffffff57ffffff0000005503030357;

	lut_sub lut_913 ({sk[304], x245x, x277x, n_n1511, x7802x, x340x, x532x}, x7806x);
	defparam lut_913.LUT_SIZE = 7;
	defparam lut_913.mask = 128'h57ffffff57ffffff0005000500053337;

	lut_sub lut_916 ({sk[305], x10x, n_n1092, x48x, x7790x, x7804x, x533x}, x7807x);
	defparam lut_916.LUT_SIZE = 7;
	defparam lut_916.mask = 128'h57ffffff57ffffff00001111000f111f;

	lut_sub lut_919 ({sk[306], i_12_, x10x, x432x, x7805x, x7806x, x7807x}, n_n1579);
	defparam lut_919.LUT_SIZE = 7;
	defparam lut_919.mask = 128'h57ffffff57ffffff7f7f7fff7f7f7f7f;

	lut_sub lut_924 ({sk[307], i_27_, i_28_, i_24_, i_29_}, x80x);
	defparam lut_924.LUT_SIZE = 5;
	defparam lut_924.mask = 32'h77778000;

	lut_sub lut_926 ({sk[308], i_9_, i_7_, i_14_, i_12_, i_23_, i_16_}, x922x);
	defparam lut_926.LUT_SIZE = 7;
	defparam lut_926.mask = 128'h57ffffff57ffffff0000800000000000;

	lut_sub lut_928 ({sk[309], i_9_, i_7_, i_14_, i_23_, i_17_, i_16_}, x923x);
	defparam lut_928.LUT_SIZE = 7;
	defparam lut_928.mask = 128'h57ffffff57ffffff0000800000000000;

	lut_sub lut_930 ({sk[310], i_31_, i_34_, i_29_, n_n1216, x922x, x923x}, x914x);
	defparam lut_930.LUT_SIZE = 7;
	defparam lut_930.mask = 128'h57ffffff57ffffff0000000000000700;

	lut_sub lut_933 ({sk[311], i_27_, i_36_, x73x, n_n1489, x323x, x291x}, x915x);
	defparam lut_933.LUT_SIZE = 7;
	defparam lut_933.mask = 128'h57ffffff57ffffff0000000700000000;

	lut_sub lut_936 ({sk[312], i_21_, x54x, n_n1404, x47x, x485x, x6999x}, x916x);
	defparam lut_936.LUT_SIZE = 7;
	defparam lut_936.mask = 128'h57ffffff57ffffff0005000500050037;

	lut_sub lut_939 ({sk[313], x43x, n_n1147, x7791x, x7792x, x74x, x7786x}, x7813x);
	defparam lut_939.LUT_SIZE = 7;
	defparam lut_939.mask = 128'h57ffffff57ffffff0000000f1111111f;

	lut_sub lut_942 ({sk[314], n_n1429, x432x, x914x, x915x, x916x, x7813x}, n_n1581);
	defparam lut_942.LUT_SIZE = 7;
	defparam lut_942.mask = 128'h57ffffff57ffffff7fff7fff7fffffff;

	lut_sub lut_948 ({sk[315], i_12_, i_24_, i_17_}, n_n1519);
	defparam lut_948.LUT_SIZE = 4;
	defparam lut_948.mask = 16'h5504;

	lut_sub lut_950 ({sk[316], i_34_, i_35_, i_38_}, n_n1419);
	defparam lut_950.LUT_SIZE = 4;
	defparam lut_950.mask = 16'h5510;

	lut_sub lut_952 ({sk[317], i_28_, i_33_, i_29_}, n_n1302);
	defparam lut_952.LUT_SIZE = 4;
	defparam lut_952.mask = 16'h5580;

	lut_sub lut_954 ({sk[318], i_9_, i_7_, i_13_}, n_n1323);
	defparam lut_954.LUT_SIZE = 4;
	defparam lut_954.mask = 16'h5520;

	lut_sub lut_956 ({sk[319], i_32_, i_31_, i_29_}, n_n1133);
	defparam lut_956.LUT_SIZE = 4;
	defparam lut_956.mask = 16'h5580;

	lut_sub lut_958 ({sk[320], i_28_, i_31_, i_29_}, n_n1128);
	defparam lut_958.LUT_SIZE = 4;
	defparam lut_958.mask = 16'h5580;

	lut_sub lut_960 ({sk[321], i_7_, i_8_, i_6_}, n_n1303);
	defparam lut_960.LUT_SIZE = 4;
	defparam lut_960.mask = 16'h5580;

	lut_sub lut_962 ({sk[322], i_26_, i_24_, i_22_}, n_n1523);
	defparam lut_962.LUT_SIZE = 4;
	defparam lut_962.mask = 16'h5580;

	lut_sub lut_964 ({sk[323], i_7_, i_6_, i_12_, i_23_, x43x, n_n1307}, n_n269);
	defparam lut_964.LUT_SIZE = 7;
	defparam lut_964.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_966 ({sk[324], i_8_, i_13_, i_16_}, x259x);
	defparam lut_966.LUT_SIZE = 4;
	defparam lut_966.mask = 16'h5580;

	lut_sub lut_968 ({sk[325], i_7_, i_5_, i_6_, i_1_, x292x, x259x}, n_n242);
	defparam lut_968.LUT_SIZE = 7;
	defparam lut_968.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_970 ({sk[326], i_32_, i_34_, i_35_}, n_n1202);
	defparam lut_970.LUT_SIZE = 4;
	defparam lut_970.mask = 16'h5540;

	lut_sub lut_972 ({sk[327], i_8_, i_14_, i_16_}, x258x);
	defparam lut_972.LUT_SIZE = 4;
	defparam lut_972.mask = 16'h5580;

	lut_sub lut_974 ({sk[328], i_7_, i_5_, i_6_, i_1_, x292x, x258x}, n_n355);
	defparam lut_974.LUT_SIZE = 7;
	defparam lut_974.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_976 ({sk[329], i_30_, i_28_, i_31_}, n_n1345);
	defparam lut_976.LUT_SIZE = 4;
	defparam lut_976.mask = 16'h5580;

	lut_sub lut_978 ({sk[330], i_9_, i_5_, i_6_, i_4_, i_1_, i_2_}, x229x);
	defparam lut_978.LUT_SIZE = 7;
	defparam lut_978.mask = 128'h57ffffff57ffffff0000000080000000;

	lut_sub lut_980 ({sk[331], i_13_, i_18_}, x347x);
	defparam lut_980.LUT_SIZE = 3;
	defparam lut_980.mask = 8'h34;

	lut_sub lut_982 ({sk[332], i_26_, i_24_, i_22_, i_33_, i_35_, i_38_}, x389x);
	defparam lut_982.LUT_SIZE = 7;
	defparam lut_982.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_984 ({sk[333], i_28_, i_26_, i_24_, i_22_, i_33_, n_n1361}, x53x);
	defparam lut_984.LUT_SIZE = 7;
	defparam lut_984.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_986 ({sk[334], i_9_, i_13_, i_18_, i_19_}, x7423x);
	defparam lut_986.LUT_SIZE = 5;
	defparam lut_986.mask = 32'h77770010;

	lut_sub lut_988 ({sk[335], i_32_, i_33_, i_35_}, n_n1458);
	defparam lut_988.LUT_SIZE = 4;
	defparam lut_988.mask = 16'h5580;

	lut_sub lut_990 ({sk[336], i_30_, i_28_, i_32_}, n_n1431);
	defparam lut_990.LUT_SIZE = 4;
	defparam lut_990.mask = 16'h5580;

	lut_sub lut_992 ({sk[337], i_20_, i_21_, i_22_}, x7491x);
	defparam lut_992.LUT_SIZE = 4;
	defparam lut_992.mask = 16'h5508;

	lut_sub lut_994 ({sk[338], i_20_, i_26_, i_21_, i_22_, x54x, n_n1406}, x62x);
	defparam lut_994.LUT_SIZE = 7;
	defparam lut_994.mask = 128'h57ffffff57ffffff0000000010000000;

	lut_sub lut_996 ({sk[339], i_28_, i_26_, i_24_, i_22_, i_33_, i_38_}, x70x);
	defparam lut_996.LUT_SIZE = 7;
	defparam lut_996.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_998 ({sk[340], i_8_, i_24_, i_38_}, x7492x);
	defparam lut_998.LUT_SIZE = 4;
	defparam lut_998.mask = 16'h5540;

	lut_sub lut_1000 ({sk[341], i_25_, i_24_, i_38_}, x239x);
	defparam lut_1000.LUT_SIZE = 4;
	defparam lut_1000.mask = 16'h5540;

	lut_sub lut_1002 ({sk[342], i_28_, i_34_, i_33_, i_29_}, x288x);
	defparam lut_1002.LUT_SIZE = 5;
	defparam lut_1002.mask = 32'h77770800;

	lut_sub lut_1004 ({sk[343], i_28_, i_25_, i_24_, i_32_, i_34_, i_29_}, x476x);
	defparam lut_1004.LUT_SIZE = 7;
	defparam lut_1004.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_1006 ({sk[344], i_24_, i_38_, x42x, x49x, n_n1340, x476x}, x1232x);
	defparam lut_1006.LUT_SIZE = 7;
	defparam lut_1006.mask = 128'h57ffffff57ffffff0000050700000505;

	lut_sub lut_1009 ({sk[345], i_12_, i_32_, n_n1307, n_n1306, n_n1303, x70x}, x1233x);
	defparam lut_1009.LUT_SIZE = 7;
	defparam lut_1009.mask = 128'h57ffffff57ffffff0015001100050000;

	lut_sub lut_1012 ({sk[346], i_20_, i_21_, i_22_, n_n1443, n_n1429, x46x}, x1234x);
	defparam lut_1012.LUT_SIZE = 7;
	defparam lut_1012.mask = 128'h57ffffff57ffffff0000000015000000;

	lut_sub lut_1015 ({sk[347], i_28_, i_34_, i_33_, i_29_, x49x, x7492x}, x1235x);
	defparam lut_1015.LUT_SIZE = 7;
	defparam lut_1015.mask = 128'h57ffffff57ffffff0000100000000000;

	lut_sub lut_1017 ({sk[348], i_12_, n_n1225, x389x, x376x, x239x, x7489x}, x7493x);
	defparam lut_1017.LUT_SIZE = 7;
	defparam lut_1017.mask = 128'h57ffffff57ffffff0055035700550055;

	lut_sub lut_1020 ({sk[349], x1232x, x1233x, x1234x, x1235x, x7493x}, n_n1881);
	defparam lut_1020.LUT_SIZE = 6;
	defparam lut_1020.mask = 64'h3f3fffff7fffffff;

	lut_sub lut_1026 ({sk[350], i_32_, i_36_, i_35_}, n_n576);
	defparam lut_1026.LUT_SIZE = 4;
	defparam lut_1026.mask = 16'h5520;

	lut_sub lut_1028 ({sk[351], i_28_, i_31_, i_29_}, n_n1499);
	defparam lut_1028.LUT_SIZE = 4;
	defparam lut_1028.mask = 16'h5520;

	lut_sub lut_1030 ({sk[352], n_n1443, n_n301, x48x, x41x, x207x, x221x}, x576x);
	defparam lut_1030.LUT_SIZE = 7;
	defparam lut_1030.mask = 128'h57ffffff57ffffff0000000f1111111f;

	lut_sub lut_1033 ({sk[353], i_23_, i_17_, i_21_, x43x, x45x, x7817x}, x902x);
	defparam lut_1033.LUT_SIZE = 7;
	defparam lut_1033.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_1035 ({sk[354], i_28_, i_21_, x79x, x242x, x49x, x258x}, x907x);
	defparam lut_1035.LUT_SIZE = 7;
	defparam lut_1035.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1037 ({sk[355], i_34_, i_36_, i_35_, x576x, x902x, x907x}, x7825x);
	defparam lut_1037.LUT_SIZE = 7;
	defparam lut_1037.mask = 128'h57ffffff57ffffff7777777777777f77;

	lut_sub lut_1041 ({sk[356], n_n1443, n_n1408, x50x, n_n576, x265x, x218x}, x577x);
	defparam lut_1041.LUT_SIZE = 7;
	defparam lut_1041.mask = 128'h57ffffff57ffffff0000050500330537;

	lut_sub lut_1044 ({sk[357], i_23_, i_21_, i_16_, x45x, x7818x, x7820x}, x903x);
	defparam lut_1044.LUT_SIZE = 7;
	defparam lut_1044.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_1046 ({sk[358], i_36_, i_35_, i_29_, x74x, x41x, n_n916}, x904x);
	defparam lut_1046.LUT_SIZE = 7;
	defparam lut_1046.mask = 128'h57ffffff57ffffff0000000001000000;

	lut_sub lut_1048 ({sk[359], i_26_, n_n1375, x54x, x577x, x903x, x904x}, x7826x);
	defparam lut_1048.LUT_SIZE = 7;
	defparam lut_1048.mask = 128'h57ffffff57ffffff7777777f77777777;

	lut_sub lut_1052 ({sk[360], i_27_, i_28_, i_23_, i_24_, i_31_, i_34_}, x84x);
	defparam lut_1052.LUT_SIZE = 7;
	defparam lut_1052.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_1054 ({sk[361], i_10_, i_7_, i_11_, i_21_, i_19_}, x440x);
	defparam lut_1054.LUT_SIZE = 6;
	defparam lut_1054.mask = 64'h3f3fffff00000020;

	lut_sub lut_1056 ({sk[362], i_28_, i_31_, n_n1397, n_n1080, x325x, x328x}, x893x);
	defparam lut_1056.LUT_SIZE = 7;
	defparam lut_1056.mask = 128'h57ffffff57ffffff0000000700000000;

	lut_sub lut_1059 ({sk[363], i_17_, i_32_, i_36_, x43x, x49x, x228x}, x894x);
	defparam lut_1059.LUT_SIZE = 7;
	defparam lut_1059.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1061 ({sk[364], i_36_, i_29_, n_n793, n_n1404, n_n1397, x376x}, x896x);
	defparam lut_1061.LUT_SIZE = 7;
	defparam lut_1061.mask = 128'h57ffffff57ffffff0000000000010000;

	lut_sub lut_1063 ({sk[365], n_n1429, x84x, x440x, x893x, x894x, x896x}, x7839x);
	defparam lut_1063.LUT_SIZE = 7;
	defparam lut_1063.mask = 128'h57ffffff57ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_1068 ({sk[366], n_n1408, x49x, x48x, x258x, x244x, x221x}, x897x);
	defparam lut_1068.LUT_SIZE = 7;
	defparam lut_1068.mask = 128'h57ffffff57ffffff0000000300001113;

	lut_sub lut_1071 ({sk[367], i_28_, i_21_, x79x, x242x, x49x, x259x}, x899x);
	defparam lut_1071.LUT_SIZE = 7;
	defparam lut_1071.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1073 ({sk[368], i_36_, n_n1375, n_n620, n_n1202, x897x, x899x}, x7840x);
	defparam lut_1073.LUT_SIZE = 7;
	defparam lut_1073.mask = 128'h57ffffff57ffffff777777777777777f;

	lut_sub lut_1077 ({sk[369], i_10_, i_7_, i_3_, i_18_}, x437x);
	defparam lut_1077.LUT_SIZE = 5;
	defparam lut_1077.mask = 32'h77770002;

	lut_sub lut_1079 ({sk[370], i_10_, i_7_, i_3_, i_11_, i_18_, i_19_}, x16x);
	defparam lut_1079.LUT_SIZE = 7;
	defparam lut_1079.mask = 128'h57ffffff57ffffff000000000000a0ec;

	lut_sub lut_1082 ({sk[371], i_23_, i_34_, i_35_}, x47x);
	defparam lut_1082.LUT_SIZE = 4;
	defparam lut_1082.mask = 16'h5540;

	lut_sub lut_1084 ({sk[372], i_27_, i_28_, i_26_, i_23_, i_24_, i_21_}, x228x);
	defparam lut_1084.LUT_SIZE = 7;
	defparam lut_1084.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_1086 ({sk[373], i_27_, i_28_, i_26_, i_29_}, x44x);
	defparam lut_1086.LUT_SIZE = 5;
	defparam lut_1086.mask = 32'h77774000;

	lut_sub lut_1088 ({sk[374], i_21_, i_31_, n_n461, x54x, n_n576, x44x}, x307x);
	defparam lut_1088.LUT_SIZE = 7;
	defparam lut_1088.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1090 ({sk[375], i_13_, i_23_, i_17_, i_16_}, x6920x);
	defparam lut_1090.LUT_SIZE = 5;
	defparam lut_1090.mask = 32'h77778000;

	lut_sub lut_1092 ({sk[376], i_27_, i_28_, i_26_, i_24_, i_31_, i_29_}, x468x);
	defparam lut_1092.LUT_SIZE = 7;
	defparam lut_1092.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_1094 ({sk[377], i_27_, i_28_, i_26_, i_23_, i_24_, i_29_}, x67x);
	defparam lut_1094.LUT_SIZE = 7;
	defparam lut_1094.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_1096 ({sk[378], n_n1443, x51x, x6920x, x468x, x67x, x207x}, x540x);
	defparam lut_1096.LUT_SIZE = 7;
	defparam lut_1096.mask = 128'h57ffffff57ffffff0000000f1111111f;

	lut_sub lut_1099 ({sk[379], i_27_, n_n1443, n_n1429, n_n1499, x16x, x47x}, x882x);
	defparam lut_1099.LUT_SIZE = 7;
	defparam lut_1099.mask = 128'h57ffffff57ffffff0001010100000000;

	lut_sub lut_1102 ({sk[380], i_17_, i_32_, i_36_, x10x, x49x, x228x}, x883x);
	defparam lut_1102.LUT_SIZE = 7;
	defparam lut_1102.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1104 ({sk[381], i_36_, i_35_, i_29_, n_n301, x74x, x41x}, x884x);
	defparam lut_1104.LUT_SIZE = 7;
	defparam lut_1104.mask = 128'h57ffffff57ffffff0000000001000000;

	lut_sub lut_1106 ({sk[382], i_21_, x54x, n_n1429, n_n576, x44x, x7847x}, x886x);
	defparam lut_1106.LUT_SIZE = 7;
	defparam lut_1106.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_1108 ({sk[383], n_n576, x540x, x882x, x883x, x884x, x886x}, x7852x);
	defparam lut_1108.LUT_SIZE = 7;
	defparam lut_1108.mask = 128'h57ffffff57ffffff7fff7fff7fffffff;

	lut_sub lut_1114 ({sk[384], i_9_, i_10_, i_6_, i_13_, n_n1307, x13x}, n_n82);
	defparam lut_1114.LUT_SIZE = 7;
	defparam lut_1114.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_1116 ({sk[385], i_14_, i_13_, i_16_}, n_n916);
	defparam lut_1116.LUT_SIZE = 4;
	defparam lut_1116.mask = 16'h5520;

	lut_sub lut_1118 ({sk[386], i_9_, i_14_, i_13_, n_n1322, x80x, x376x}, x878x);
	defparam lut_1118.LUT_SIZE = 7;
	defparam lut_1118.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1120 ({sk[387], i_34_, i_36_, x85x, x48x, n_n916, x878x}, x877x);
	defparam lut_1120.LUT_SIZE = 7;
	defparam lut_1120.mask = 128'h57ffffff57ffffff0000000000005557;

	lut_sub lut_1123 ({sk[388], i_27_, i_36_, x242x, x49x, x258x, x214x}, x873x);
	defparam lut_1123.LUT_SIZE = 7;
	defparam lut_1123.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_1125 ({sk[389], i_17_, x43x, x10x, x50x, x228x, x265x}, x874x);
	defparam lut_1125.LUT_SIZE = 7;
	defparam lut_1125.mask = 128'h57ffffff57ffffff0001010100000000;

	lut_sub lut_1128 ({sk[390], x51x, x46x, x7862x, x7858x, x7861x, x7857x}, x875x);
	defparam lut_1128.LUT_SIZE = 7;
	defparam lut_1128.mask = 128'h57ffffff57ffffff0000003300050037;

	lut_sub lut_1131 ({sk[391], i_27_, i_28_, i_23_, i_36_, i_29_, n_n1202}, x7863x);
	defparam lut_1131.LUT_SIZE = 7;
	defparam lut_1131.mask = 128'h57ffffff57ffffff0400000000000000;

	lut_sub lut_1133 ({sk[392], n_n1408, x49x, x873x, x874x, x875x, x7863x}, x7866x);
	defparam lut_1133.LUT_SIZE = 7;
	defparam lut_1133.mask = 128'h57ffffff57ffffff3fff3fff3fff7fff;

	lut_sub lut_1138 ({sk[393], i_27_, x73x, x51x, x260x, n_n1128, n_n576}, x862x);
	defparam lut_1138.LUT_SIZE = 7;
	defparam lut_1138.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_1140 ({sk[394], i_27_, n_n1443, x54x, x50x, n_n1128, x86x}, x865x);
	defparam lut_1140.LUT_SIZE = 7;
	defparam lut_1140.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_1142 ({sk[395], i_13_, n_n1216, x51x, n_n1322, n_n1133, x86x}, x866x);
	defparam lut_1142.LUT_SIZE = 7;
	defparam lut_1142.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_1144 ({sk[396], i_12_, x10x, x307x, x862x, x865x, x866x}, x7876x);
	defparam lut_1144.LUT_SIZE = 7;
	defparam lut_1144.mask = 128'h57ffffff57ffffff7f7f7fff7f7f7f7f;

	lut_sub lut_1149 ({sk[397], i_34_, i_36_, i_35_}, x86x);
	defparam lut_1149.LUT_SIZE = 4;
	defparam lut_1149.mask = 16'h5502;

	lut_sub lut_1151 ({sk[398], i_34_, i_36_}, x244x);
	defparam lut_1151.LUT_SIZE = 3;
	defparam lut_1151.mask = 8'h31;

	lut_sub lut_1153 ({sk[399], i_27_, i_28_, i_23_, i_31_, i_34_, i_35_}, x275x);
	defparam lut_1153.LUT_SIZE = 7;
	defparam lut_1153.mask = 128'h57ffffff57ffffff0400000000000000;

	lut_sub lut_1155 ({sk[400], i_9_, i_5_, i_6_, i_13_, i_4_, i_2_}, x218x);
	defparam lut_1155.LUT_SIZE = 7;
	defparam lut_1155.mask = 128'h57ffffff57ffffff0800000000000000;

	lut_sub lut_1157 ({sk[401], i_27_, i_28_, i_23_, i_24_, i_32_, i_29_}, x221x);
	defparam lut_1157.LUT_SIZE = 7;
	defparam lut_1157.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_1159 ({sk[402], n_n1408, x48x, x41x, n_n916, x218x, x221x}, x543x);
	defparam lut_1159.LUT_SIZE = 7;
	defparam lut_1159.mask = 128'h57ffffff57ffffff0000000f1111111f;

	lut_sub lut_1162 ({sk[403], i_10_, i_7_, i_11_}, n_n712);
	defparam lut_1162.LUT_SIZE = 4;
	defparam lut_1162.mask = 16'h5502;

	lut_sub lut_1164 ({sk[404], i_21_, i_19_, n_n1443, n_n1429, x437x, n_n712}, x542x);
	defparam lut_1164.LUT_SIZE = 7;
	defparam lut_1164.mask = 128'h57ffffff57ffffff0000000007770333;

	lut_sub lut_1169 ({sk[405], n_n82, x86x, x543x, x7878x, x852x, x853x}, x7881x);
	defparam lut_1169.LUT_SIZE = 7;
	defparam lut_1169.mask = 128'h57ffffff57ffffff777777ff7f7f7fff;

	lut_sub lut_1174 ({sk[406], i_34_, n_n301, x85x, x48x, x871x, x872x}, x563x);
	defparam lut_1174.LUT_SIZE = 7;
	defparam lut_1174.mask = 128'h57ffffff57ffffff777777777777777f;

	lut_sub lut_1178 ({sk[407], i_17_, x10x, x50x, x265x, x868x, x67x}, x863x);
	defparam lut_1178.LUT_SIZE = 7;
	defparam lut_1178.mask = 128'h57ffffff57ffffff0303030703030303;

	lut_sub lut_1181 ({sk[408], i_14_, i_21_, i_16_, n_n461, n_n1141, x46x}, x846x);
	defparam lut_1181.LUT_SIZE = 7;
	defparam lut_1181.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_1183 ({sk[409], i_27_, i_34_, n_n1443, x54x, x49x, n_n1288}, x844x);
	defparam lut_1183.LUT_SIZE = 7;
	defparam lut_1183.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_1185 ({sk[410], i_36_, i_29_, x74x, n_n355, x846x, x844x}, x843x);
	defparam lut_1185.LUT_SIZE = 7;
	defparam lut_1185.mask = 128'h57ffffff57ffffff00000000777f7777;

	lut_sub lut_1189 ({sk[411], i_27_, i_14_, n_n1390, x42x, x11x, x7884x}, x839x);
	defparam lut_1189.LUT_SIZE = 7;
	defparam lut_1189.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1191 ({sk[412], i_21_, n_n1443, n_n1429, x437x, x16x, x84x}, x840x);
	defparam lut_1191.LUT_SIZE = 7;
	defparam lut_1191.mask = 128'h57ffffff57ffffff0000000000051115;

	lut_sub lut_1194 ({sk[413], i_31_, i_29_, n_n1216, x76x, n_n1263, x86x}, x841x);
	defparam lut_1194.LUT_SIZE = 7;
	defparam lut_1194.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1196 ({sk[414], x48x, n_n242, x244x, x839x, x840x, x841x}, x7895x);
	defparam lut_1196.LUT_SIZE = 7;
	defparam lut_1196.mask = 128'h57ffffff57ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_1201 ({sk[415], i_13_, i_21_, i_16_, n_n461, n_n1141, x46x}, x838x);
	defparam lut_1201.LUT_SIZE = 7;
	defparam lut_1201.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_1203 ({sk[416], i_26_, i_32_, n_n1375, n_n1443, x54x, x49x}, x836x);
	defparam lut_1203.LUT_SIZE = 7;
	defparam lut_1203.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1205 ({sk[417], i_36_, i_29_, x74x, n_n242, x838x, x836x}, x834x);
	defparam lut_1205.LUT_SIZE = 7;
	defparam lut_1205.mask = 128'h57ffffff57ffffff00000000777f7777;

	lut_sub lut_1209 ({sk[418], i_31_, i_29_, n_n793, n_n1397, x325x, x328x}, x830x);
	defparam lut_1209.LUT_SIZE = 7;
	defparam lut_1209.mask = 128'h57ffffff57ffffff0000000000070000;

	lut_sub lut_1212 ({sk[419], i_36_, i_35_, n_n1369, n_n1314, x76x, n_n1128}, x831x);
	defparam lut_1212.LUT_SIZE = 7;
	defparam lut_1212.mask = 128'h57ffffff57ffffff0000000000010000;

	lut_sub lut_1214 ({sk[420], i_27_, i_28_, i_29_, n_n1429, n_n1334, x393x}, x832x);
	defparam lut_1214.LUT_SIZE = 7;
	defparam lut_1214.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_1216 ({sk[421], i_10_, i_21_, n_n1443, x54x, x7900x, x44x}, x833x);
	defparam lut_1216.LUT_SIZE = 7;
	defparam lut_1216.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1218 ({sk[422], i_36_, n_n461, n_n1369, n_n1147, n_n460, n_n1254}, x835x);
	defparam lut_1218.LUT_SIZE = 7;
	defparam lut_1218.mask = 128'h57ffffff57ffffff0000000000000001;

	lut_sub lut_1220 ({sk[423], x830x, x831x, x832x, x833x, x835x}, x7909x);
	defparam lut_1220.LUT_SIZE = 6;
	defparam lut_1220.mask = 64'h3f3fffff7fffffff;

	lut_sub lut_1226 ({sk[424], i_17_, i_32_, i_36_, x10x, x49x, x67x}, x820x);
	defparam lut_1226.LUT_SIZE = 7;
	defparam lut_1226.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1228 ({sk[425], i_31_, i_29_, n_n1216, n_n1314, x76x, x86x}, x821x);
	defparam lut_1228.LUT_SIZE = 7;
	defparam lut_1228.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1230 ({sk[426], i_36_, i_29_, n_n793, n_n1429, n_n1397, x376x}, x822x);
	defparam lut_1230.LUT_SIZE = 7;
	defparam lut_1230.mask = 128'h57ffffff57ffffff0000000000010000;

	lut_sub lut_1232 ({sk[427], n_n1375, x227x, n_n269, x820x, x821x, x822x}, x7919x);
	defparam lut_1232.LUT_SIZE = 7;
	defparam lut_1232.mask = 128'h57ffffff57ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_1237 ({sk[428], i_27_, i_31_, x73x, x42x, x76x, n_n1263}, x829x);
	defparam lut_1237.LUT_SIZE = 7;
	defparam lut_1237.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1239 ({sk[429], i_14_, i_13_, n_n1390, x11x, x7913x, x7914x}, x7915x);
	defparam lut_1239.LUT_SIZE = 7;
	defparam lut_1239.mask = 128'h57ffffff57ffffff0007000300050000;

	lut_sub lut_1242 ({sk[430], i_13_, i_21_, x54x, n_n1408, x7900x, x44x}, x825x);
	defparam lut_1242.LUT_SIZE = 7;
	defparam lut_1242.mask = 128'h57ffffff57ffffff0000000000010000;

	lut_sub lut_1244 ({sk[431], i_7_, n_n461, x79x, x415x, n_n460, n_n1254}, x826x);
	defparam lut_1244.LUT_SIZE = 7;
	defparam lut_1244.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_1246 ({sk[432], i_36_, i_35_, x829x, x7915x, x825x, x826x}, x7920x);
	defparam lut_1246.LUT_SIZE = 7;
	defparam lut_1246.mask = 128'h57ffffff57ffffff777777777fff7777;

	lut_sub lut_1251 ({sk[433], i_28_, i_26_, i_24_}, n_n1497);
	defparam lut_1251.LUT_SIZE = 4;
	defparam lut_1251.mask = 16'h5580;

	lut_sub lut_1253 ({sk[434], i_9_, i_6_, i_13_}, n_n839);
	defparam lut_1253.LUT_SIZE = 4;
	defparam lut_1253.mask = 16'h5540;

	lut_sub lut_1255 ({sk[435], i_32_, i_34_, i_33_}, n_n1311);
	defparam lut_1255.LUT_SIZE = 4;
	defparam lut_1255.mask = 16'h5580;

	lut_sub lut_1257 ({sk[436], i_9_, i_8_, i_5_, i_6_}, x7420x);
	defparam lut_1257.LUT_SIZE = 5;
	defparam lut_1257.mask = 32'h77770080;

	lut_sub lut_1259 ({sk[437], i_9_, i_5_, i_6_, i_19_}, x7424x);
	defparam lut_1259.LUT_SIZE = 5;
	defparam lut_1259.mask = 32'h77770040;

	lut_sub lut_1261 ({sk[438], i_9_, i_8_, i_13_}, n_n1028);
	defparam lut_1261.LUT_SIZE = 4;
	defparam lut_1261.mask = 16'h5508;

	lut_sub lut_1263 ({sk[439], i_30_, i_29_}, x57x);
	defparam lut_1263.LUT_SIZE = 3;
	defparam lut_1263.mask = 8'h38;

	lut_sub lut_1265 ({sk[440], i_30_, i_7_, i_8_}, x77x);
	defparam lut_1265.LUT_SIZE = 4;
	defparam lut_1265.mask = 16'h5580;

	lut_sub lut_1267 ({sk[441], i_28_, i_34_, i_35_, i_29_}, x372x);
	defparam lut_1267.LUT_SIZE = 5;
	defparam lut_1267.mask = 32'h77771000;

	lut_sub lut_1269 ({sk[442], i_28_, i_25_, i_26_, i_29_}, x71x);
	defparam lut_1269.LUT_SIZE = 5;
	defparam lut_1269.mask = 32'h77778000;

	lut_sub lut_1271 ({sk[443], i_28_, i_25_, i_26_, i_24_, i_38_, i_29_}, x395x);
	defparam lut_1271.LUT_SIZE = 7;
	defparam lut_1271.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_1273 ({sk[444], i_7_, i_32_}, x211x);
	defparam lut_1273.LUT_SIZE = 3;
	defparam lut_1273.mask = 8'h38;

	lut_sub lut_1275 ({sk[445], i_30_, i_7_, i_28_, i_32_, i_29_}, x474x);
	defparam lut_1275.LUT_SIZE = 6;
	defparam lut_1275.mask = 64'h3f3fffff80000000;

	lut_sub lut_1277 ({sk[446], i_14_, i_34_, i_33_, i_35_}, x1137x);
	defparam lut_1277.LUT_SIZE = 5;
	defparam lut_1277.mask = 32'h77770010;

	lut_sub lut_1279 ({sk[447], i_27_, i_23_, i_16_, i_31_, i_34_, i_35_}, x1138x);
	defparam lut_1279.LUT_SIZE = 7;
	defparam lut_1279.mask = 128'h57ffffff57ffffff0004040404040404;

	lut_sub lut_1283 ({sk[448], i_30_, i_7_, i_32_}, x7602x);
	defparam lut_1283.LUT_SIZE = 4;
	defparam lut_1283.mask = 16'h5580;

	lut_sub lut_1285 ({sk[449], i_28_, i_22_, x395x, x1137x, x1138x, x7602x}, x7608x);
	defparam lut_1285.LUT_SIZE = 7;
	defparam lut_1285.mask = 128'h57ffffff57ffffff00553f7f00550055;

	lut_sub lut_1289 ({sk[450], i_14_, i_13_, i_16_}, n_n1387);
	defparam lut_1289.LUT_SIZE = 4;
	defparam lut_1289.mask = 16'h5508;

	lut_sub lut_1291 ({sk[451], i_9_, i_10_, i_24_}, n_n1359);
	defparam lut_1291.LUT_SIZE = 4;
	defparam lut_1291.mask = 16'h5508;

	lut_sub lut_1293 ({sk[452], i_27_, i_23_, i_21_}, n_n1080);
	defparam lut_1293.LUT_SIZE = 4;
	defparam lut_1293.mask = 16'h5540;

	lut_sub lut_1295 ({sk[453], i_23_, i_21_, i_16_}, n_n1254);
	defparam lut_1295.LUT_SIZE = 4;
	defparam lut_1295.mask = 16'h5580;

	lut_sub lut_1297 ({sk[454], i_30_, i_32_, i_31_, i_34_, i_33_, i_35_}, x479x);
	defparam lut_1297.LUT_SIZE = 7;
	defparam lut_1297.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_1299 ({sk[455], i_25_, i_26_, i_23_, i_24_, i_34_}, x806x);
	defparam lut_1299.LUT_SIZE = 6;
	defparam lut_1299.mask = 64'h3f3fffff0000c840;

	lut_sub lut_1302 ({sk[456], i_30_, i_28_, i_32_, i_31_, i_33_, i_29_}, x6950x);
	defparam lut_1302.LUT_SIZE = 7;
	defparam lut_1302.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_1304 ({sk[457], i_14_, i_25_, x42x, x479x, x806x, x6950x}, x7928x);
	defparam lut_1304.LUT_SIZE = 7;
	defparam lut_1304.mask = 128'h57ffffff57ffffff1111111f111f111f;

	lut_sub lut_1308 ({sk[458], i_34_, x302x, x54x, n_n1489, n_n1438, x214x}, x564x);
	defparam lut_1308.LUT_SIZE = 7;
	defparam lut_1308.mask = 128'h57ffffff57ffffff111111111111111f;

	lut_sub lut_1311 ({sk[459], n_n1375, n_n1374, x340x, x1038x, x1039x, x7925x}, x7927x);
	defparam lut_1311.LUT_SIZE = 7;
	defparam lut_1311.mask = 128'h57ffffff57ffffff0055005500553f7f;

	lut_sub lut_1315 ({sk[460], i_7_, i_36_, x7928x, x564x, x7927x}, n_n1585);
	defparam lut_1315.LUT_SIZE = 6;
	defparam lut_1315.mask = 64'h3f3fffff5f7f5f5f;

	lut_sub lut_1319 ({sk[461], i_32_, i_34_, i_35_}, n_n1422);
	defparam lut_1319.LUT_SIZE = 4;
	defparam lut_1319.mask = 16'h5520;

	lut_sub lut_1321 ({sk[462], i_14_, i_12_, i_17_, i_16_}, x8x);
	defparam lut_1321.LUT_SIZE = 5;
	defparam lut_1321.mask = 32'h7777a800;

	lut_sub lut_1324 ({sk[463], i_14_, i_13_, i_23_, i_24_, i_17_, i_16_}, x1038x);
	defparam lut_1324.LUT_SIZE = 7;
	defparam lut_1324.mask = 128'h57ffffff57ffffff0000000080000000;

	lut_sub lut_1326 ({sk[464], i_14_, i_13_, i_12_, i_23_, i_24_, i_16_}, x1039x);
	defparam lut_1326.LUT_SIZE = 7;
	defparam lut_1326.mask = 128'h57ffffff57ffffff0000000080000000;

	lut_sub lut_1328 ({sk[465], x54x, x215x, x398x, x44x, x805x, x7026x}, x803x);
	defparam lut_1328.LUT_SIZE = 7;
	defparam lut_1328.mask = 128'h57ffffff57ffffff0000555503ff57ff;

	lut_sub lut_1332 ({sk[466], i_22_, x803x}, x1662x);
	defparam lut_1332.LUT_SIZE = 3;
	defparam lut_1332.mask = 8'h31;

	lut_sub lut_1334 ({sk[467], i_30_, i_28_, i_23_, i_24_, i_34_, i_29_}, x7683x);
	defparam lut_1334.LUT_SIZE = 7;
	defparam lut_1334.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_1336 ({sk[468], i_30_, i_22_, i_32_, i_31_}, x7029x);
	defparam lut_1336.LUT_SIZE = 5;
	defparam lut_1336.mask = 32'h77770800;

	lut_sub lut_1338 ({sk[469], i_23_, i_24_, i_22_, i_34_}, x7025x);
	defparam lut_1338.LUT_SIZE = 5;
	defparam lut_1338.mask = 32'h77771000;

	lut_sub lut_1340 ({sk[470], i_27_, i_28_, i_22_, i_34_, i_29_, x54x}, x308x);
	defparam lut_1340.LUT_SIZE = 7;
	defparam lut_1340.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1342 ({sk[471], i_27_, i_28_, i_26_, i_33_}, x6958x);
	defparam lut_1342.LUT_SIZE = 5;
	defparam lut_1342.mask = 32'h77774000;

	lut_sub lut_1344 ({sk[472], i_27_, i_28_, i_25_, i_26_, i_33_, x54x}, x309x);
	defparam lut_1344.LUT_SIZE = 7;
	defparam lut_1344.mask = 128'h57ffffff57ffffff0010000000000000;

	lut_sub lut_1346 ({sk[473], i_30_, i_31_, i_29_}, n_n1459);
	defparam lut_1346.LUT_SIZE = 4;
	defparam lut_1346.mask = 16'h5580;

	lut_sub lut_1348 ({sk[474], i_30_, i_28_, i_23_, i_24_, i_31_, i_29_}, x419x);
	defparam lut_1348.LUT_SIZE = 7;
	defparam lut_1348.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_1350 ({sk[475], i_30_, i_28_, i_26_, i_24_, i_31_, i_29_}, x513x);
	defparam lut_1350.LUT_SIZE = 7;
	defparam lut_1350.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_1352 ({sk[476], n_n1404, n_n1408, x309x, x7933x, x7934x, x7935x}, x7938x);
	defparam lut_1352.LUT_SIZE = 7;
	defparam lut_1352.mask = 128'h57ffffff57ffffff7f7f7fff7fff7fff;

	lut_sub lut_1358 ({sk[477], i_24_, i_35_, i_38_}, x12x);
	defparam lut_1358.LUT_SIZE = 4;
	defparam lut_1358.mask = 16'h5540;

	lut_sub lut_1360 ({sk[478], i_28_, i_34_, i_33_, i_19_, i_29_, x12x}, n_n338);
	defparam lut_1360.LUT_SIZE = 7;
	defparam lut_1360.mask = 128'h57ffffff57ffffff0000040000000000;

	lut_sub lut_1362 ({sk[479], i_11_, i_17_, i_16_, i_19_}, x431x);
	defparam lut_1362.LUT_SIZE = 5;
	defparam lut_1362.mask = 32'h77778000;

	lut_sub lut_1364 ({sk[480], i_3_, i_11_, i_18_, i_17_, i_16_, i_19_}, x549x);
	defparam lut_1364.LUT_SIZE = 7;
	defparam lut_1364.mask = 128'h57ffffff57ffffff80800000c080c000;

	lut_sub lut_1367 ({sk[481], i_27_, i_28_, i_23_, i_24_, i_34_, i_29_}, x273x);
	defparam lut_1367.LUT_SIZE = 7;
	defparam lut_1367.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_1369 ({sk[482], i_9_, i_14_, i_13_, n_n1397, x376x, x220x}, x966x);
	defparam lut_1369.LUT_SIZE = 7;
	defparam lut_1369.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1371 ({sk[483], n_n1288, x14x, n_n916, x318x, x256x, x326x}, x7758x);
	defparam lut_1371.LUT_SIZE = 7;
	defparam lut_1371.mask = 128'h57ffffff57ffffff000011110000111f;

	lut_sub lut_1374 ({sk[484], x1765x, x1766x, x273x, x966x, x7758x}, x548x);
	defparam lut_1374.LUT_SIZE = 6;
	defparam lut_1374.mask = 64'h3f3fffff777f7f7f;

	lut_sub lut_1379 ({sk[485], n_n1375, n_n1322, x211x, x496x, x7944x, x7945x}, x573x);
	defparam lut_1379.LUT_SIZE = 7;
	defparam lut_1379.mask = 128'h57ffffff57ffffff0005000500053337;

	lut_sub lut_1382 ({sk[486], i_13_, i_23_, i_21_, i_16_, x368x, x7946x}, x459x);
	defparam lut_1382.LUT_SIZE = 7;
	defparam lut_1382.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_1384 ({sk[487], i_7_, i_36_, x10x, n_n1489, n_n1258, n_n1202}, x469x);
	defparam lut_1384.LUT_SIZE = 7;
	defparam lut_1384.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_1386 ({sk[488], n_n793, n_n1375, n_n846, x7942x, x342x, x572x}, x7952x);
	defparam lut_1386.LUT_SIZE = 7;
	defparam lut_1386.mask = 128'h57ffffff57ffffff0000003305050537;

	lut_sub lut_1389 ({sk[489], n_n1443, n_n1429, n_n1406, x228x, x7951x, x7948x}, x7953x);
	defparam lut_1389.LUT_SIZE = 7;
	defparam lut_1389.mask = 128'h57ffffff57ffffff0000050500330537;

	lut_sub lut_1392 ({sk[490], i_14_, x573x, x459x, x469x, x7952x, x7953x}, n_n1574);
	defparam lut_1392.LUT_SIZE = 7;
	defparam lut_1392.mask = 128'h57ffffff57ffffff7fffffff7fff7fff;

	lut_sub lut_1398 ({sk[491], i_30_, i_36_, n_n1397, x323x, n_n846, x348x}, x574x);
	defparam lut_1398.LUT_SIZE = 7;
	defparam lut_1398.mask = 128'h57ffffff57ffffff1111111f11111111;

	lut_sub lut_1401 ({sk[492], i_13_, x211x, x496x, x220x, x7944x, x7961x}, x412x);
	defparam lut_1401.LUT_SIZE = 7;
	defparam lut_1401.mask = 128'h57ffffff57ffffff0303035700000000;

	lut_sub lut_1404 ({sk[493], i_7_, i_36_, x43x, n_n1489, n_n1258, n_n1202}, x424x);
	defparam lut_1404.LUT_SIZE = 7;
	defparam lut_1404.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_1406 ({sk[494], n_n1441, x228x, x77x, x342x, x385x, x7957x}, x7963x);
	defparam lut_1406.LUT_SIZE = 7;
	defparam lut_1406.mask = 128'h57ffffff57ffffff0000005503030357;

	lut_sub lut_1409 ({sk[495], x227x, n_n1147, x48x, x258x, n_n846, x7962x}, x7964x);
	defparam lut_1409.LUT_SIZE = 7;
	defparam lut_1409.mask = 128'h57ffffff57ffffff0003000300035557;

	lut_sub lut_1412 ({sk[496], n_n1375, x574x, x412x, x424x, x7963x, x7964x}, n_n1575);
	defparam lut_1412.LUT_SIZE = 7;
	defparam lut_1412.mask = 128'h57ffffff57ffffff7fff7fff7fffffff;

	lut_sub lut_1418 ({sk[497], i_30_, i_31_, n_n1202, x7969x, x7972x, x7973x}, x7978x);
	defparam lut_1418.LUT_SIZE = 7;
	defparam lut_1418.mask = 128'h57ffffff57ffffff111f111111111111;

	lut_sub lut_1421 ({sk[498], n_n1216, x7784x, x324x, x325x, x328x, x7974x}, x7979x);
	defparam lut_1421.LUT_SIZE = 7;
	defparam lut_1421.mask = 128'h57ffffff57ffffff15151515151515ff;

	lut_sub lut_1425 ({sk[499], x79x, n_n1147, n_n1089, x7787x, x7788x, x7975x}, x7980x);
	defparam lut_1425.LUT_SIZE = 7;
	defparam lut_1425.mask = 128'h57ffffff57ffffff0003000300035557;

	lut_sub lut_1428 ({sk[500], i_14_, x43x, n_n1393, x441x, x496x, x7977x}, x7981x);
	defparam lut_1428.LUT_SIZE = 7;
	defparam lut_1428.mask = 128'h57ffffff57ffffff00001111000f111f;

	lut_sub lut_1431 ({sk[501], x7978x, x7979x, x7980x, x7981x}, n_n1578);
	defparam lut_1431.LUT_SIZE = 5;
	defparam lut_1431.mask = 32'h77777fff;

	lut_sub lut_1436 ({sk[502], i_27_, x58x, x74x, x258x, x385x, x348x}, x195x);
	defparam lut_1436.LUT_SIZE = 7;
	defparam lut_1436.mask = 128'h57ffffff57ffffff0003111300030003;

	lut_sub lut_1439 ({sk[503], i_25_, i_21_, x220x, x505x, x668x, x7987x}, x7989x);
	defparam lut_1439.LUT_SIZE = 7;
	defparam lut_1439.mask = 128'h57ffffff57ffffff0055005500550357;

	lut_sub lut_1442 ({sk[504], x79x, n_n1089, x48x, x259x, n_n846, x7975x}, x7990x);
	defparam lut_1442.LUT_SIZE = 7;
	defparam lut_1442.mask = 128'h57ffffff57ffffff0003000300035557;

	lut_sub lut_1445 ({sk[505], i_23_, n_n1375, x10x, x496x, x7977x, x7988x}, x7991x);
	defparam lut_1445.LUT_SIZE = 7;
	defparam lut_1445.mask = 128'h57ffffff57ffffff0003005700030003;

	lut_sub lut_1448 ({sk[506], x195x, x7989x, x7990x, x7991x}, n_n1576);
	defparam lut_1448.LUT_SIZE = 5;
	defparam lut_1448.mask = 32'h77777fff;

	lut_sub lut_1453 ({sk[507], i_23_, i_16_, n_n1374, x7997x, x7998x, x8000x}, x188x);
	defparam lut_1453.LUT_SIZE = 7;
	defparam lut_1453.mask = 128'h57ffffff57ffffff0357000003030000;

	lut_sub lut_1456 ({sk[508], i_14_, i_28_, i_31_, i_33_, x3x, n_n1397}, x189x);
	defparam lut_1456.LUT_SIZE = 7;
	defparam lut_1456.mask = 128'h57ffffff57ffffff0000000004000000;

	lut_sub lut_1458 ({sk[509], i_9_, i_7_, i_12_, n_n1375, n_n1504, n_n1314}, x187x);
	defparam lut_1458.LUT_SIZE = 7;
	defparam lut_1458.mask = 128'h57ffffff57ffffff0000010000000000;

	lut_sub lut_1460 ({sk[510], n_n1375, n_n1322, x74x, x259x, x385x, x7996x}, x8001x);
	defparam lut_1460.LUT_SIZE = 7;
	defparam lut_1460.mask = 128'h57ffffff57ffffff0003000300035557;

	lut_sub lut_1463 ({sk[511], n_n1092, x7804x, n_n1511, x7802x, x687x, x7995x}, x8002x);
	defparam lut_1463.LUT_SIZE = 7;
	defparam lut_1463.mask = 128'h57ffffff57ffffff0005000500053337;

	lut_sub lut_1466 ({sk[512], i_21_, x188x, x189x, x187x, x8001x, x8002x}, n_n1577);
	defparam lut_1466.LUT_SIZE = 7;
	defparam lut_1466.mask = 128'h57ffffff57ffffff7f7f7f7f7fffffff;

	lut_sub lut_1472 ({sk[513], i_20_, i_23_, i_21_, i_34_, i_35_}, x7951x);
	defparam lut_1472.LUT_SIZE = 6;
	defparam lut_1472.mask = 64'h3f3fffff00004000;

	lut_sub lut_1474 ({sk[514], i_27_, i_28_, i_31_, x245x, x325x}, x172x);
	defparam lut_1474.LUT_SIZE = 6;
	defparam lut_1474.mask = 64'h3f3fffff01000000;

	lut_sub lut_1476 ({sk[515], i_27_, i_36_, x73x, n_n1263, x321x, n_n1288}, x173x);
	defparam lut_1476.LUT_SIZE = 7;
	defparam lut_1476.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_1478 ({sk[516], i_14_, i_23_, i_21_, i_16_, x368x, x7946x}, x175x);
	defparam lut_1478.LUT_SIZE = 7;
	defparam lut_1478.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_1480 ({sk[517], n_n1404, n_n1406, x7951x, x172x, x173x, x175x}, x8016x);
	defparam lut_1480.LUT_SIZE = 7;
	defparam lut_1480.mask = 128'h57ffffff57ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_1485 ({sk[518], i_8_, i_31_, i_36_, i_35_, x496x, x8008x}, x352x);
	defparam lut_1485.LUT_SIZE = 7;
	defparam lut_1485.mask = 128'h57ffffff57ffffff0010000000000000;

	lut_sub lut_1487 ({sk[519], i_27_, i_26_, x54x, n_n1404, x42x, x376x}, x181x);
	defparam lut_1487.LUT_SIZE = 7;
	defparam lut_1487.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1489 ({sk[520], n_n1429, n_n1314, x321x, x376x, x273x, x256x}, x8007x);
	defparam lut_1489.LUT_SIZE = 7;
	defparam lut_1489.mask = 128'h57ffffff57ffffff0000005503030357;

	lut_sub lut_1492 ({sk[521], i_2_, i_21_, x43x, n_n1369, x242x, x8011x}, x177x);
	defparam lut_1492.LUT_SIZE = 7;
	defparam lut_1492.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1494 ({sk[522], i_13_, i_36_, x352x, x181x, x8007x, x177x}, x8017x);
	defparam lut_1494.LUT_SIZE = 7;
	defparam lut_1494.mask = 128'h57ffffff57ffffff55ff7fff55557f7f;

	lut_sub lut_1499 ({sk[523], i_13_, i_12_, i_17_, i_16_, x393x, x382x}, x711x);
	defparam lut_1499.LUT_SIZE = 7;
	defparam lut_1499.mask = 128'h57ffffff57ffffff7050700000000000;

	lut_sub lut_1503 ({sk[524], i_13_, i_16_, x54x, x11x, n_n1133, x8018x}, x162x);
	defparam lut_1503.LUT_SIZE = 7;
	defparam lut_1503.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1505 ({sk[525], i_27_, i_28_, i_31_, x245x, x328x}, x163x);
	defparam lut_1505.LUT_SIZE = 6;
	defparam lut_1505.mask = 64'h3f3fffff01000000;

	lut_sub lut_1507 ({sk[526], i_27_, x42x, n_n1334, x711x, x162x, x163x}, x8025x);
	defparam lut_1507.LUT_SIZE = 7;
	defparam lut_1507.mask = 128'h57ffffff57ffffff7777777f77777777;

	lut_sub lut_1511 ({sk[527], i_27_, i_2_, i_21_, x73x, x242x, x8011x}, x295x);
	defparam lut_1511.LUT_SIZE = 7;
	defparam lut_1511.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_1513 ({sk[528], n_n1404, n_n1263, x321x, x376x, x273x, x256x}, x712x);
	defparam lut_1513.LUT_SIZE = 7;
	defparam lut_1513.mask = 128'h57ffffff57ffffff0000005503030357;

	lut_sub lut_1516 ({sk[529], i_14_, i_16_, i_36_, x295x, x352x, x712x}, x8026x);
	defparam lut_1516.LUT_SIZE = 7;
	defparam lut_1516.mask = 128'h57ffffff57ffffff3f7f337700550055;

	lut_sub lut_1520 ({sk[530], i_27_, i_34_, x54x, n_n1499, x325x, x328x}, x155x);
	defparam lut_1520.LUT_SIZE = 7;
	defparam lut_1520.mask = 128'h57ffffff57ffffff0000000700000000;

	lut_sub lut_1523 ({sk[531], i_30_, i_27_, i_36_, x42x, n_n1397, x324x}, x158x);
	defparam lut_1523.LUT_SIZE = 7;
	defparam lut_1523.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1525 ({sk[532], i_27_, n_n1429, n_n1368, x7951x, x155x, x158x}, x8037x);
	defparam lut_1525.LUT_SIZE = 7;
	defparam lut_1525.mask = 128'h57ffffff57ffffff7777777f77777777;

	lut_sub lut_1529 ({sk[533], i_27_, i_28_, i_26_, i_31_}, x305x);
	defparam lut_1529.LUT_SIZE = 5;
	defparam lut_1529.mask = 32'h77774000;

	lut_sub lut_1531 ({sk[534], i_10_, i_7_, i_11_, i_19_, x54x, x8021x}, x723x);
	defparam lut_1531.LUT_SIZE = 7;
	defparam lut_1531.mask = 128'h57ffffff57ffffff0000000000003111;

	lut_sub lut_1534 ({sk[535], i_2_, i_17_, i_36_, x10x, x228x, x77x}, x156x);
	defparam lut_1534.LUT_SIZE = 7;
	defparam lut_1534.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1536 ({sk[536], i_27_, i_36_, x73x, n_n1314, x321x, n_n1288}, x159x);
	defparam lut_1536.LUT_SIZE = 7;
	defparam lut_1536.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_1538 ({sk[537], i_7_, i_36_, x415x, n_n1489, n_n1202, n_n1251}, x160x);
	defparam lut_1538.LUT_SIZE = 7;
	defparam lut_1538.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_1540 ({sk[538], n_n1443, x305x, x723x, x156x, x159x, x160x}, x8038x);
	defparam lut_1540.LUT_SIZE = 7;
	defparam lut_1540.mask = 128'h57ffffff57ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_1545 ({sk[539], i_21_, i_36_, i_35_, n_n1441, x54x, n_n1438}, x478x);
	defparam lut_1545.LUT_SIZE = 7;
	defparam lut_1545.mask = 128'h57ffffff57ffffff0000010000000000;

	lut_sub lut_1547 ({sk[540], i_27_, i_31_, x58x, n_n1429, x393x, x382x}, x141x);
	defparam lut_1547.LUT_SIZE = 7;
	defparam lut_1547.mask = 128'h57ffffff57ffffff0000000700000000;

	lut_sub lut_1550 ({sk[541], i_9_, i_7_, i_12_, n_n793, x10x, x7942x}, x142x);
	defparam lut_1550.LUT_SIZE = 7;
	defparam lut_1550.mask = 128'h57ffffff57ffffff0000010000000000;

	lut_sub lut_1552 ({sk[542], i_26_, i_36_, n_n1375, x54x, n_n1429, x376x}, x146x);
	defparam lut_1552.LUT_SIZE = 7;
	defparam lut_1552.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_1554 ({sk[543], i_20_, i_23_, i_21_, n_n1397, n_n1406, n_n1408}, x150x);
	defparam lut_1554.LUT_SIZE = 7;
	defparam lut_1554.mask = 128'h57ffffff57ffffff0000000001000000;

	lut_sub lut_1556 ({sk[544], n_n1404, x478x, x141x, x142x, x146x, x150x}, x8048x);
	defparam lut_1556.LUT_SIZE = 7;
	defparam lut_1556.mask = 128'h57ffffff57ffffff7fff7fff7fffffff;

	lut_sub lut_1562 ({sk[545], i_27_, i_16_}, x103x);
	defparam lut_1562.LUT_SIZE = 3;
	defparam lut_1562.mask = 8'h37;

	lut_sub lut_1565 ({sk[546], i_27_, i_23_, i_16_}, n_n1251);
	defparam lut_1565.LUT_SIZE = 4;
	defparam lut_1565.mask = 16'h5580;

	lut_sub lut_1567 ({sk[547], i_27_, i_23_, i_22_, i_35_}, x6947x);
	defparam lut_1567.LUT_SIZE = 5;
	defparam lut_1567.mask = 32'h77771000;

	lut_sub lut_1569 ({sk[548], i_27_, i_23_, i_17_, i_34_, i_35_}, x318x);
	defparam lut_1569.LUT_SIZE = 6;
	defparam lut_1569.mask = 64'h3f3fffff40000000;

	lut_sub lut_1571 ({sk[549], i_27_, i_14_, i_13_, i_12_, i_23_, i_16_}, x7499x);
	defparam lut_1571.LUT_SIZE = 7;
	defparam lut_1571.mask = 128'h57ffffff57ffffff0000800000000000;

	lut_sub lut_1573 ({sk[550], i_27_, i_28_, i_26_, i_24_, i_31_}, x236x);
	defparam lut_1573.LUT_SIZE = 6;
	defparam lut_1573.mask = 64'h3f3fffff40000000;

	lut_sub lut_1575 ({sk[551], i_27_, i_28_, i_26_, i_24_, i_0_, i_29_}, x355x);
	defparam lut_1575.LUT_SIZE = 7;
	defparam lut_1575.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_1577 ({sk[552], i_30_, i_28_, i_26_, i_24_, i_21_, i_34_}, x441x);
	defparam lut_1577.LUT_SIZE = 7;
	defparam lut_1577.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_1579 ({sk[553], i_30_, i_28_, i_26_, i_24_, i_34_}, x215x);
	defparam lut_1579.LUT_SIZE = 6;
	defparam lut_1579.mask = 64'h3f3fffff80000000;

	lut_sub lut_1581 ({sk[554], i_30_, i_28_, i_21_, i_34_, x54x, x215x}, x551x);
	defparam lut_1581.LUT_SIZE = 7;
	defparam lut_1581.mask = 128'h57ffffff57ffffff0057005500550055;

	lut_sub lut_1584 ({sk[555], i_13_, i_12_, i_23_, i_21_, i_16_}, x137x);
	defparam lut_1584.LUT_SIZE = 6;
	defparam lut_1584.mask = 64'h3f3fffff80000000;

	lut_sub lut_1586 ({sk[556], i_14_, i_23_, i_17_, i_21_, i_16_}, x138x);
	defparam lut_1586.LUT_SIZE = 6;
	defparam lut_1586.mask = 64'h3f3fffff80000000;

	lut_sub lut_1588 ({sk[557], i_33_, x42x, n_n1397, n_n1258, n_n1387, x7499x}, x8059x);
	defparam lut_1588.LUT_SIZE = 7;
	defparam lut_1588.mask = 128'h57ffffff57ffffff0000000000000057;

	lut_sub lut_1591 ({sk[558], i_34_, n_n1404, n_n1368, x6947x, x236x, x8058x}, x8060x);
	defparam lut_1591.LUT_SIZE = 7;
	defparam lut_1591.mask = 128'h57ffffff57ffffff1111111f11111111;

	lut_sub lut_1594 ({sk[559], n_n1443, x46x, x7491x, x355x, x137x, x138x}, x8061x);
	defparam lut_1594.LUT_SIZE = 7;
	defparam lut_1594.mask = 128'h57ffffff57ffffff07070707070707ff;

	lut_sub lut_1598 ({sk[560], i_25_, n_n1393, x551x, x8059x, x8060x, x8061x}, n_n1583);
	defparam lut_1598.LUT_SIZE = 7;
	defparam lut_1598.mask = 128'h57ffffff57ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_1603 ({sk[561], i_21_, x54x, n_n1408, x47x, x485x, x6999x}, x119x);
	defparam lut_1603.LUT_SIZE = 7;
	defparam lut_1603.mask = 128'h57ffffff57ffffff0005000500050037;

	lut_sub lut_1606 ({sk[562], i_29_, n_n1334, n_n1216, n_n1322, n_n1323, x8066x}, x120x);
	defparam lut_1606.LUT_SIZE = 7;
	defparam lut_1606.mask = 128'h57ffffff57ffffff0000005700000000;

	lut_sub lut_1609 ({sk[563], i_28_, i_25_, i_21_, x355x, x479x, x8064x}, x8067x);
	defparam lut_1609.LUT_SIZE = 7;
	defparam lut_1609.mask = 128'h57ffffff57ffffff0505053705050505;

	lut_sub lut_1612 ({sk[564], n_n1429, x62x, x8x, x119x, x120x, x8067x}, n_n1582);
	defparam lut_1612.LUT_SIZE = 7;
	defparam lut_1612.mask = 128'h57ffffff57ffffff7f7f7fff7f7fffff;

	lut_sub lut_1618 ({sk[565], i_25_, i_23_, i_24_, i_34_, i_33_}, x6944x);
	defparam lut_1618.LUT_SIZE = 6;
	defparam lut_1618.mask = 64'h3f3fffff00001000;

	lut_sub lut_1620 ({sk[566], n_n1375, n_n1443, n_n1408, n_n1326, x6947x, x6944x}, x104x);
	defparam lut_1620.LUT_SIZE = 7;
	defparam lut_1620.mask = 128'h57ffffff57ffffff0000030300550357;

	lut_sub lut_1623 ({sk[567], i_9_, i_7_, i_13_, i_12_, i_23_, i_16_}, x115x);
	defparam lut_1623.LUT_SIZE = 7;
	defparam lut_1623.mask = 128'h57ffffff57ffffff0000800000000000;

	lut_sub lut_1625 ({sk[568], i_28_, i_31_, n_n1369, n_n1322, x115x, x557x}, x109x);
	defparam lut_1625.LUT_SIZE = 7;
	defparam lut_1625.mask = 128'h57ffffff57ffffff0000003700000000;

	lut_sub lut_1628 ({sk[569], n_n1429, n_n1408, n_n1326, x6947x, x355x, x8070x}, x8071x);
	defparam lut_1628.LUT_SIZE = 7;
	defparam lut_1628.mask = 128'h57ffffff57ffffff1111111f111f111f;

	lut_sub lut_1632 ({sk[570], n_n1375, n_n1404, x104x, x6944x, x109x, x8071x}, n_n1584);
	defparam lut_1632.LUT_SIZE = 7;
	defparam lut_1632.mask = 128'h57ffffff57ffffff77ff77ff77ff7fff;

	lut_sub lut_1637 ({sk[571], i_28_, i_34_, i_35_, i_29_}, x214x);
	defparam lut_1637.LUT_SIZE = 5;
	defparam lut_1637.mask = 32'h77772000;

	lut_sub lut_1639 ({sk[572], i_31_, i_36_, i_35_}, x265x);
	defparam lut_1639.LUT_SIZE = 4;
	defparam lut_1639.mask = 16'h5520;

	lut_sub lut_1641 ({sk[573], i_17_, i_29_, n_n793, x43x, x49x, n_n1202}, x871x);
	defparam lut_1641.LUT_SIZE = 7;
	defparam lut_1641.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1643 ({sk[574], i_27_, i_23_, i_17_, x49x, x259x, x214x}, x872x);
	defparam lut_1643.LUT_SIZE = 7;
	defparam lut_1643.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_1645 ({sk[575], i_8_, i_5_, i_6_, i_4_, i_12_}, x7818x);
	defparam lut_1645.LUT_SIZE = 6;
	defparam lut_1645.mask = 64'h3f3fffff80000000;

	lut_sub lut_1647 ({sk[576], i_14_, i_23_, i_21_, i_16_, x45x, x7818x}, x868x);
	defparam lut_1647.LUT_SIZE = 7;
	defparam lut_1647.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_1649 ({sk[577], i_7_, i_8_, i_23_, i_17_, i_21_, i_36_}, x7762x);
	defparam lut_1649.LUT_SIZE = 7;
	defparam lut_1649.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_1651 ({sk[578], i_14_, i_13_, i_17_, i_16_}, x420x);
	defparam lut_1651.LUT_SIZE = 5;
	defparam lut_1651.mask = 32'h77770800;

	lut_sub lut_1653 ({sk[579], i_7_, i_32_, i_36_}, x7769x);
	defparam lut_1653.LUT_SIZE = 4;
	defparam lut_1653.mask = 16'h5540;

	lut_sub lut_1655 ({sk[580], i_28_, i_32_, i_29_, x14x, x318x}, x87x);
	defparam lut_1655.LUT_SIZE = 6;
	defparam lut_1655.mask = 64'h3f3fffff10000000;

	lut_sub lut_1657 ({sk[581], i_27_, i_28_, i_34_, i_35_, i_29_, n_n1322}, x373x);
	defparam lut_1657.LUT_SIZE = 7;
	defparam lut_1657.mask = 128'h57ffffff57ffffff0400000000000000;

	lut_sub lut_1659 ({sk[582], n_n1422, x7145x, x7146x, x7148x, x7149x, x7764x}, x956x);
	defparam lut_1659.LUT_SIZE = 7;
	defparam lut_1659.mask = 128'h57ffffff57ffffff0000000001010155;

	lut_sub lut_1662 ({sk[583], i_9_, x43x, n_n1278, n_n787, n_n179, x256x}, x957x);
	defparam lut_1662.LUT_SIZE = 7;
	defparam lut_1662.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_1664 ({sk[584], n_n301, n_n82, x87x, x373x, x956x, x957x}, x566x);
	defparam lut_1664.LUT_SIZE = 7;
	defparam lut_1664.mask = 128'h57ffffff57ffffff77777f7f77ff7fff;

	lut_sub lut_1669 ({sk[585], i_10_, i_14_, i_13_, i_17_, i_16_}, x571x);
	defparam lut_1669.LUT_SIZE = 6;
	defparam lut_1669.mask = 64'h3f3fffff88800800;

	lut_sub lut_1672 ({sk[586], i_10_, i_21_, x232x, x54x, x7769x, x44x}, x949x);
	defparam lut_1672.LUT_SIZE = 7;
	defparam lut_1672.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1674 ({sk[587], i_9_, i_5_, i_6_, x54x, x7146x, x7149x}, x7x);
	defparam lut_1674.LUT_SIZE = 7;
	defparam lut_1674.mask = 128'h57ffffff57ffffff0700030005000000;

	lut_sub lut_1677 ({sk[588], i_27_, i_29_, x58x, n_n576, x949x, x7x}, x569x);
	defparam lut_1677.LUT_SIZE = 7;
	defparam lut_1677.mask = 128'h57ffffff57ffffff3337333333333333;

	lut_sub lut_1680 ({sk[589], i_14_, i_13_, i_17_, i_21_, i_16_}, x7776x);
	defparam lut_1680.LUT_SIZE = 6;
	defparam lut_1680.mask = 64'h3f3fffff00800000;

	lut_sub lut_1682 ({sk[590], i_34_, i_33_, i_35_, i_38_}, n_n1059);
	defparam lut_1682.LUT_SIZE = 5;
	defparam lut_1682.mask = 32'h77771000;

	lut_sub lut_1684 ({sk[591], i_30_, i_31_, i_34_, i_36_, i_35_}, n_n846);
	defparam lut_1684.LUT_SIZE = 6;
	defparam lut_1684.mask = 64'h3f3fffff02000000;

	lut_sub lut_1686 ({sk[592], i_18_, i_17_}, x6890x);
	defparam lut_1686.LUT_SIZE = 3;
	defparam lut_1686.mask = 8'h38;

	lut_sub lut_1688 ({sk[593], i_21_, i_31_, i_34_, i_35_}, x7942x);
	defparam lut_1688.LUT_SIZE = 5;
	defparam lut_1688.mask = 32'h77770004;

	lut_sub lut_1690 ({sk[594], i_8_, i_14_, i_12_, i_23_, i_24_, i_16_}, x342x);
	defparam lut_1690.LUT_SIZE = 7;
	defparam lut_1690.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_1692 ({sk[595], i_30_, i_32_, i_31_, i_36_, i_35_}, x7948x);
	defparam lut_1692.LUT_SIZE = 6;
	defparam lut_1692.mask = 64'h3f3fffff20000000;

	lut_sub lut_1694 ({sk[596], i_30_, i_8_, i_28_, i_12_, i_31_}, x7946x);
	defparam lut_1694.LUT_SIZE = 6;
	defparam lut_1694.mask = 64'h3f3fffff80000000;

	lut_sub lut_1696 ({sk[597], i_30_, i_27_, i_28_, i_26_, i_23_, i_24_}, x496x);
	defparam lut_1696.LUT_SIZE = 7;
	defparam lut_1696.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_1698 ({sk[598], i_30_, i_7_, i_8_, i_34_, i_36_, i_35_}, x7944x);
	defparam lut_1698.LUT_SIZE = 7;
	defparam lut_1698.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_1700 ({sk[599], i_2_, i_17_, i_21_, i_16_, i_36_}, x7945x);
	defparam lut_1700.LUT_SIZE = 6;
	defparam lut_1700.mask = 64'h3f3fffff40000000;

	lut_sub lut_1702 ({sk[600], i_9_, i_7_, i_13_, i_12_, i_17_, i_16_}, x572x);
	defparam lut_1702.LUT_SIZE = 7;
	defparam lut_1702.mask = 128'h57ffffff57ffffff0000a80000000000;

	lut_sub lut_1705 ({sk[601], i_30_, i_31_, i_36_, i_35_, i_29_}, x385x);
	defparam lut_1705.LUT_SIZE = 6;
	defparam lut_1705.mask = 64'h3f3fffff08000000;

	lut_sub lut_1707 ({sk[602], i_30_, i_27_, i_28_, i_23_, i_16_, i_29_}, x7962x);
	defparam lut_1707.LUT_SIZE = 7;
	defparam lut_1707.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_1709 ({sk[603], i_8_, i_13_, i_12_, i_23_, i_24_, i_16_}, x348x);
	defparam lut_1709.LUT_SIZE = 7;
	defparam lut_1709.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_1711 ({sk[604], i_9_, i_8_, i_18_, n_n1278, n_n787, x257x}, x1462x);
	defparam lut_1711.LUT_SIZE = 7;
	defparam lut_1711.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_1713 ({sk[605], i_18_, i_32_, x204x, n_n1278, x14x, x404x}, x581x);
	defparam lut_1713.LUT_SIZE = 7;
	defparam lut_1713.mask = 128'h57ffffff57ffffff0537000000330000;

	lut_sub lut_1716 ({sk[606], i_12_, n_n762, x61x, x262x, x582x, x7261x}, x1456x);
	defparam lut_1716.LUT_SIZE = 7;
	defparam lut_1716.mask = 128'h57ffffff57ffffff000011110000111f;

	lut_sub lut_1719 ({sk[607], i_9_, i_8_, i_13_, i_11_}, x7427x);
	defparam lut_1719.LUT_SIZE = 5;
	defparam lut_1719.mask = 32'h77770040;

	lut_sub lut_1721 ({sk[608], i_9_, i_13_, i_11_, i_18_}, x7428x);
	defparam lut_1721.LUT_SIZE = 5;
	defparam lut_1721.mask = 32'h77770010;

	lut_sub lut_1723 ({sk[609], i_1_, x292x, n_n1118, x208x, x7427x, x7428x}, x20x);
	defparam lut_1723.LUT_SIZE = 7;
	defparam lut_1723.mask = 128'h57ffffff57ffffff0303035703030303;

	lut_sub lut_1726 ({sk[610], i_3_, i_13_, i_18_, i_22_, i_19_}, x5x);
	defparam lut_1726.LUT_SIZE = 6;
	defparam lut_1726.mask = 64'h3f3fffff44000400;

	lut_sub lut_1729 ({sk[611], i_3_, i_13_, i_11_, i_18_, i_22_, i_19_}, x23x);
	defparam lut_1729.LUT_SIZE = 7;
	defparam lut_1729.mask = 128'h57ffffff57ffffff444c0000040c0000;

	lut_sub lut_1733 ({sk[612], i_28_, i_24_, i_35_, i_38_, i_29_, n_n1340}, x253x);
	defparam lut_1733.LUT_SIZE = 7;
	defparam lut_1733.mask = 128'h57ffffff57ffffff0400000000000000;

	lut_sub lut_1735 ({sk[613], i_28_, i_26_, i_24_, i_33_, i_35_, i_38_}, x509x);
	defparam lut_1735.LUT_SIZE = 7;
	defparam lut_1735.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_1737 ({sk[614], i_11_, x11x, n_n1048, x213x, x7425x, x7424x}, x24x);
	defparam lut_1737.LUT_SIZE = 7;
	defparam lut_1737.mask = 128'h57ffffff57ffffff07070707070707ff;

	lut_sub lut_1741 ({sk[615], i_10_, i_12_, i_31_, x3x, x23x, x509x}, x1281x);
	defparam lut_1741.LUT_SIZE = 7;
	defparam lut_1741.mask = 128'h57ffffff57ffffff0000000000001000;

	lut_sub lut_1743 ({sk[616], x208x, x50x, x71x, x12x, x7427x, x7428x}, x1283x);
	defparam lut_1743.LUT_SIZE = 7;
	defparam lut_1743.mask = 128'h57ffffff57ffffff0000000500030007;

	lut_sub lut_1746 ({sk[617], i_30_, i_28_, i_22_, i_32_}, x7612x);
	defparam lut_1746.LUT_SIZE = 5;
	defparam lut_1746.mask = 32'h77771030;

	lut_sub lut_1749 ({sk[618], i_28_, i_25_, i_24_, i_38_, i_29_}, x7613x);
	defparam lut_1749.LUT_SIZE = 6;
	defparam lut_1749.mask = 64'h3f3fffff20000000;

	lut_sub lut_1751 ({sk[619], i_12_, i_24_, i_17_, x77x, x7612x, x7613x}, x7614x);
	defparam lut_1751.LUT_SIZE = 7;
	defparam lut_1751.mask = 128'h57ffffff57ffffff0505050505370505;

	lut_sub lut_1754 ({sk[620], i_14_, i_13_, i_12_, i_17_}, x585x);
	defparam lut_1754.LUT_SIZE = 5;
	defparam lut_1754.mask = 32'h7777111f;

	lut_sub lut_1757 ({sk[621], i_30_, i_14_, i_28_, i_13_, i_22_, i_32_}, x1127x);
	defparam lut_1757.LUT_SIZE = 7;
	defparam lut_1757.mask = 128'h57ffffff57ffffff0000010000000300;

	lut_sub lut_1760 ({sk[622], i_30_, i_7_, i_8_, i_28_, i_29_}, x369x);
	defparam lut_1760.LUT_SIZE = 6;
	defparam lut_1760.mask = 64'h3f3fffff80000000;

	lut_sub lut_1762 ({sk[623], i_28_, i_31_, i_34_, i_35_, i_29_}, x7610x);
	defparam lut_1762.LUT_SIZE = 6;
	defparam lut_1762.mask = 64'h3f3fffff00200000;

	lut_sub lut_1764 ({sk[624], n_n1300, x298x, x585x, x1127x, x369x, x7610x}, x7615x);
	defparam lut_1764.LUT_SIZE = 7;
	defparam lut_1764.mask = 128'h57ffffff57ffffff00550f5f00553f7f;

	lut_sub lut_1768 ({sk[625], i_34_, n_n1489, x239x, x211x, x7614x, x7615x}, n_n1889);
	defparam lut_1768.LUT_SIZE = 7;
	defparam lut_1768.mask = 128'h57ffffff57ffffff555555557777777f;

	lut_sub lut_1772 ({sk[626], i_14_, i_13_, i_12_, i_24_, i_17_}, x588x);
	defparam lut_1772.LUT_SIZE = 6;
	defparam lut_1772.mask = 64'h3f3fffff040404cc;

	lut_sub lut_1775 ({sk[627], i_30_, i_27_, i_23_, i_16_, i_32_}, x587x);
	defparam lut_1775.LUT_SIZE = 6;
	defparam lut_1775.mask = 64'h3f3fffff15553fff;

	lut_sub lut_1782 ({sk[628], i_28_, i_25_, i_26_, x57x, x7600x, x1134x}, x7606x);
	defparam lut_1782.LUT_SIZE = 7;
	defparam lut_1782.mask = 128'h57ffffff57ffffff5755555555555555;

	lut_sub lut_1785 ({sk[629], i_26_, i_24_, x42x, n_n1300, x77x, x474x}, x7607x);
	defparam lut_1785.LUT_SIZE = 7;
	defparam lut_1785.mask = 128'h57ffffff57ffffff0507000000000000;

	lut_sub lut_1788 ({sk[630], x588x, x587x, x7616x, x7617x, x7618x, x7619x}, x7621x);
	defparam lut_1788.LUT_SIZE = 7;
	defparam lut_1788.mask = 128'h57ffffff57ffffff000f333f555f777f;

	lut_sub lut_1792 ({sk[631], x7608x, x7606x, x7607x, x7621x}, x7622x);
	defparam lut_1792.LUT_SIZE = 5;
	defparam lut_1792.mask = 32'h77777fff;

	lut_sub lut_1797 ({sk[632], i_9_, i_18_, x204x, n_n787, n_n1118, x41x}, x801x);
	defparam lut_1797.LUT_SIZE = 7;
	defparam lut_1797.mask = 128'h57ffffff57ffffff0357005500550055;

	lut_sub lut_1800 ({sk[633], i_18_, i_24_, x204x, n_n1118, x404x, x41x}, x30x);
	defparam lut_1800.LUT_SIZE = 7;
	defparam lut_1800.mask = 128'h57ffffff57ffffff0357000000550000;

	lut_sub lut_1803 ({sk[634], i_30_, i_28_, i_25_, i_26_, i_24_, i_22_}, x313x);
	defparam lut_1803.LUT_SIZE = 7;
	defparam lut_1803.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_1805 ({sk[635], i_30_, i_25_, i_24_, i_22_, x58x, n_n1361}, x56x);
	defparam lut_1805.LUT_SIZE = 7;
	defparam lut_1805.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_1807 ({sk[636], i_10_, i_3_, i_13_, i_12_, i_11_}, x210x);
	defparam lut_1807.LUT_SIZE = 6;
	defparam lut_1807.mask = 64'h3f3fffff00001000;

	lut_sub lut_1809 ({sk[637], i_31_, i_33_, i_35_, i_38_}, x226x);
	defparam lut_1809.LUT_SIZE = 5;
	defparam lut_1809.mask = 32'h77774000;

	lut_sub lut_1811 ({sk[638], i_26_, i_24_, i_32_, i_33_, i_35_, i_38_}, x294x);
	defparam lut_1811.LUT_SIZE = 7;
	defparam lut_1811.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_1813 ({sk[639], n_n1307, n_n787, n_n1128, x294x, x361x, x353x}, x1447x);
	defparam lut_1813.LUT_SIZE = 7;
	defparam lut_1813.mask = 128'h57ffffff57ffffff0000000500030007;

	lut_sub lut_1816 ({sk[640], i_7_, i_33_, i_38_, n_n1523, n_n1431, x210x}, x1448x);
	defparam lut_1816.LUT_SIZE = 7;
	defparam lut_1816.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1818 ({sk[641], i_26_, i_31_, i_33_, i_35_, i_38_, x42x}, x7275x);
	defparam lut_1818.LUT_SIZE = 7;
	defparam lut_1818.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_1820 ({sk[642], n_n1361, n_n1038, x313x, x414x, x590x, x1452x}, x1450x);
	defparam lut_1820.LUT_SIZE = 7;
	defparam lut_1820.mask = 128'h57ffffff57ffffff00000000005f007f;

	lut_sub lut_1824 ({sk[643], i_25_, i_26_, i_24_, i_35_, i_38_}, x81x);
	defparam lut_1824.LUT_SIZE = 6;
	defparam lut_1824.mask = 64'h3f3fffff40000000;

	lut_sub lut_1826 ({sk[644], i_30_, i_28_, i_33_, i_35_, i_38_}, x7287x);
	defparam lut_1826.LUT_SIZE = 6;
	defparam lut_1826.mask = 64'h3f3fffff40000000;

	lut_sub lut_1828 ({sk[645], i_9_, i_3_, i_13_, i_12_, i_11_, i_22_}, x1442x);
	defparam lut_1828.LUT_SIZE = 7;
	defparam lut_1828.mask = 128'h57ffffff57ffffff0000000002000000;

	lut_sub lut_1830 ({sk[646], i_3_, i_13_, i_12_, i_11_, i_18_, i_19_}, x807x);
	defparam lut_1830.LUT_SIZE = 7;
	defparam lut_1830.mask = 128'h57ffffff57ffffff0057000000130000;

	lut_sub lut_1834 ({sk[647], i_10_, i_38_, x211x, x313x, x210x, x807x}, x1431x);
	defparam lut_1834.LUT_SIZE = 7;
	defparam lut_1834.mask = 128'h57ffffff57ffffff0000000300000007;

	lut_sub lut_1837 ({sk[648], i_9_, i_18_, x204x, n_n1278, n_n787, x14x}, x36x);
	defparam lut_1837.LUT_SIZE = 7;
	defparam lut_1837.mask = 128'h57ffffff57ffffff0357005500550055;

	lut_sub lut_1840 ({sk[649], i_28_, i_25_, i_26_, i_22_, x7292x, x7306x}, x1418x);
	defparam lut_1840.LUT_SIZE = 7;
	defparam lut_1840.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_1842 ({sk[650], n_n1307, n_n787, x237x, n_n1133, x361x, x353x}, x1420x);
	defparam lut_1842.LUT_SIZE = 7;
	defparam lut_1842.mask = 128'h57ffffff57ffffff0000000500030007;

	lut_sub lut_1845 ({sk[651], i_28_, n_n1305, n_n1419, x36x, x1418x, x1420x}, x7313x);
	defparam lut_1845.LUT_SIZE = 7;
	defparam lut_1845.mask = 128'h57ffffff57ffffff7777777f77777777;

	lut_sub lut_1849 ({sk[652], i_24_, i_32_, i_31_, i_35_, i_38_}, x7314x);
	defparam lut_1849.LUT_SIZE = 6;
	defparam lut_1849.mask = 64'h3f3fffff40000000;

	lut_sub lut_1851 ({sk[653], i_10_, i_7_, n_n1523, n_n1431, x807x}, x1413x);
	defparam lut_1851.LUT_SIZE = 6;
	defparam lut_1851.mask = 64'h3f3fffff00000100;

	lut_sub lut_1853 ({sk[654], n_n1307, n_n787, x71x, x7314x, x361x, x353x}, x1409x);
	defparam lut_1853.LUT_SIZE = 7;
	defparam lut_1853.mask = 128'h57ffffff57ffffff0000000500030007;

	lut_sub lut_1856 ({sk[655], i_28_, i_25_, i_26_, i_22_, x7292x, x7294x}, x1428x);
	defparam lut_1856.LUT_SIZE = 7;
	defparam lut_1856.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_1858 ({sk[656], i_25_, i_31_, i_35_, i_38_, i_29_, x58x}, x7296x);
	defparam lut_1858.LUT_SIZE = 7;
	defparam lut_1858.mask = 128'h57ffffff57ffffff0400000000000000;

	lut_sub lut_1860 ({sk[657], i_10_, x13x, x205x, x210x, x7300x, x7298x}, x1430x);
	defparam lut_1860.LUT_SIZE = 7;
	defparam lut_1860.mask = 128'h57ffffff57ffffff0000000300000013;

	lut_sub lut_1863 ({sk[658], x30x, x1431x, x1409x, x1428x, x7296x, x1430x}, x7315x);
	defparam lut_1863.LUT_SIZE = 7;
	defparam lut_1863.mask = 128'h57ffffff57ffffff5fffffff7fffffff;

	lut_sub lut_1869 ({sk[659], i_34_, i_33_, i_35_, i_38_, x30x, x1422x}, x623x);
	defparam lut_1869.LUT_SIZE = 7;
	defparam lut_1869.mask = 128'h57ffffff57ffffff5555555557555555;

	lut_sub lut_1872 ({sk[660], i_30_, i_33_, i_38_, x58x, x1413x, x595x}, x1408x);
	defparam lut_1872.LUT_SIZE = 7;
	defparam lut_1872.mask = 128'h57ffffff57ffffff0037000000330000;

	lut_sub lut_1875 ({sk[661], i_28_, i_25_, i_24_, i_34_, i_38_, i_29_}, x7318x);
	defparam lut_1875.LUT_SIZE = 7;
	defparam lut_1875.mask = 128'h57ffffff57ffffff0200000000000000;

	lut_sub lut_1877 ({sk[662], i_28_, i_24_, i_34_, i_33_, i_38_, i_29_}, x7323x);
	defparam lut_1877.LUT_SIZE = 7;
	defparam lut_1877.mask = 128'h57ffffff57ffffff0020000000000000;

	lut_sub lut_1879 ({sk[663], x50x, x52x, n_n1191, x229x, x7321x, x7319x}, x7325x);
	defparam lut_1879.LUT_SIZE = 7;
	defparam lut_1879.mask = 128'h57ffffff57ffffff0003000300035557;

	lut_sub lut_1882 ({sk[664], x204x, n_n416, x15x, x7318x, x7323x, x7325x}, x7327x);
	defparam lut_1882.LUT_SIZE = 7;
	defparam lut_1882.mask = 128'h57ffffff57ffffff55555f5f557f5f7f;

	lut_sub lut_1887 ({sk[665], i_34_, i_33_, i_38_}, x7332x);
	defparam lut_1887.LUT_SIZE = 4;
	defparam lut_1887.mask = 16'h5504;

	lut_sub lut_1889 ({sk[666], i_9_, i_10_, i_33_, n_n1361, x50x, x61x}, x1393x);
	defparam lut_1889.LUT_SIZE = 7;
	defparam lut_1889.mask = 128'h57ffffff57ffffff0000000001000000;

	lut_sub lut_1891 ({sk[667], i_32_, i_31_, n_n1361, n_n1307, x257x, n_n839}, x1394x);
	defparam lut_1891.LUT_SIZE = 7;
	defparam lut_1891.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_1893 ({sk[668], i_9_, i_13_, i_25_, x42x, n_n1419, x376x}, x1395x);
	defparam lut_1893.LUT_SIZE = 7;
	defparam lut_1893.mask = 128'h57ffffff57ffffff0000010000000000;

	lut_sub lut_1895 ({sk[669], i_13_, i_24_, i_31_, n_n1361, x41x, x78x}, x1396x);
	defparam lut_1895.LUT_SIZE = 7;
	defparam lut_1895.mask = 128'h57ffffff57ffffff0000000001000000;

	lut_sub lut_1897 ({sk[670], x58x, n_n1191, x229x, x41x, x7328x, x7330x}, x7335x);
	defparam lut_1897.LUT_SIZE = 7;
	defparam lut_1897.mask = 128'h57ffffff57ffffff0000050500000537;

	lut_sub lut_1900 ({sk[671], i_9_, i_10_, i_8_, n_n1361, x11x, x52x}, x1380x);
	defparam lut_1900.LUT_SIZE = 7;
	defparam lut_1900.mask = 128'h57ffffff57ffffff0000000001000000;

	lut_sub lut_1902 ({sk[672], i_9_, i_10_, i_24_, x50x, x271x}, x1384x);
	defparam lut_1902.LUT_SIZE = 6;
	defparam lut_1902.mask = 64'h3f3fffff00001000;

	lut_sub lut_1904 ({sk[673], i_31_, n_n1307, n_n853, n_n300, x1380x, x1384x}, x7346x);
	defparam lut_1904.LUT_SIZE = 7;
	defparam lut_1904.mask = 128'h57ffffff57ffffff7777777f77777777;

	lut_sub lut_1908 ({sk[674], i_13_, x1388x, x1389x, x1385x, x1387x}, x726x);
	defparam lut_1908.LUT_SIZE = 6;
	defparam lut_1908.mask = 64'h3f3fffff7fff7777;

	lut_sub lut_1913 ({sk[675], i_9_, i_10_, i_13_, i_32_, x14x, x376x}, x725x);
	defparam lut_1913.LUT_SIZE = 7;
	defparam lut_1913.mask = 128'h57ffffff57ffffff5575003000300030;

	lut_sub lut_1916 ({sk[676], i_25_, x42x, n_n1419, x56x, x726x, x725x}, x7347x);
	defparam lut_1916.LUT_SIZE = 7;
	defparam lut_1916.mask = 128'h57ffffff57ffffff0303035703030303;

	lut_sub lut_1919 ({sk[677], i_20_, i_7_, i_13_, i_17_, i_16_}, x399x);
	defparam lut_1919.LUT_SIZE = 6;
	defparam lut_1919.mask = 64'h3f3fffff00000080;

	lut_sub lut_1921 ({sk[678], i_30_, i_28_, i_26_, i_23_, i_24_, i_34_}, x599x);
	defparam lut_1921.LUT_SIZE = 7;
	defparam lut_1921.mask = 128'h57ffffff57ffffffc840000000000000;

	lut_sub lut_1924 ({sk[679], i_28_, i_21_, i_34_, i_35_, i_29_}, x1712x);
	defparam lut_1924.LUT_SIZE = 6;
	defparam lut_1924.mask = 64'h3f3fffff00100000;

	lut_sub lut_1926 ({sk[680], n_n1396, n_n1429, n_n1406, n_n1408, x245x, x6958x}, x6963x);
	defparam lut_1926.LUT_SIZE = 7;
	defparam lut_1926.mask = 128'h57ffffff57ffffff0003003300035577;

	lut_sub lut_1930 ({sk[681], i_20_, i_2_, i_23_, i_17_, x10x, x45x}, x1706x);
	defparam lut_1930.LUT_SIZE = 7;
	defparam lut_1930.mask = 128'h57ffffff57ffffff0000100000000000;

	lut_sub lut_1932 ({sk[682], i_28_, i_33_, i_29_, n_n1438, x1712x, x6957x}, x1707x);
	defparam lut_1932.LUT_SIZE = 7;
	defparam lut_1932.mask = 128'h57ffffff57ffffff0703030303030303;

	lut_sub lut_1935 ({sk[683], i_20_, i_25_, n_n1393, x84x, x399x, x599x}, x6961x);
	defparam lut_1935.LUT_SIZE = 7;
	defparam lut_1935.mask = 128'h57ffffff57ffffff0303030303030357;

	lut_sub lut_1938 ({sk[684], x6963x, x1706x, x1707x, x6961x}, n_n1718);
	defparam lut_1938.LUT_SIZE = 5;
	defparam lut_1938.mask = 32'h77777fff;

	lut_sub lut_1943 ({sk[685], i_27_, i_28_, i_24_, i_34_, i_37_}, x316x);
	defparam lut_1943.LUT_SIZE = 6;
	defparam lut_1943.mask = 64'h3f3fffff10000000;

	lut_sub lut_1945 ({sk[686], i_27_, i_23_, i_24_, i_34_, i_37_}, x6929x);
	defparam lut_1945.LUT_SIZE = 6;
	defparam lut_1945.mask = 64'h3f3fffff10000000;

	lut_sub lut_1947 ({sk[687], i_28_, i_33_, i_29_, x6929x}, x317x);
	defparam lut_1947.LUT_SIZE = 5;
	defparam lut_1947.mask = 32'h77774000;

	lut_sub lut_1949 ({sk[688], i_8_, i_17_, x10x, x49x, x48x, x221x}, x601x);
	defparam lut_1949.LUT_SIZE = 7;
	defparam lut_1949.mask = 128'h57ffffff57ffffff0007000300050000;

	lut_sub lut_1952 ({sk[689], i_27_, i_28_, i_24_, i_32_, i_34_, i_29_}, x256x);
	defparam lut_1952.LUT_SIZE = 7;
	defparam lut_1952.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_1954 ({sk[690], n_n1408, x51x, x260x, x50x, x273x, x256x}, x600x);
	defparam lut_1954.LUT_SIZE = 7;
	defparam lut_1954.mask = 128'h57ffffff57ffffff0000005503030357;

	lut_sub lut_1957 ({sk[691], i_23_, i_37_, n_n1375, x10x, x321x, n_n1202}, x1734x);
	defparam lut_1957.LUT_SIZE = 7;
	defparam lut_1957.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_1959 ({sk[692], i_32_, i_33_, i_29_, n_n1314, x321x, x316x}, x1735x);
	defparam lut_1959.LUT_SIZE = 7;
	defparam lut_1959.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_1961 ({sk[693], i_35_, i_37_, x600x, x1734x, x1735x}, x6933x);
	defparam lut_1961.LUT_SIZE = 6;
	defparam lut_1961.mask = 64'h3f3fffff777f7777;

	lut_sub lut_1965 ({sk[694], i_28_, i_32_, i_29_, x51x, x6920x, x6921x}, x1732x);
	defparam lut_1965.LUT_SIZE = 7;
	defparam lut_1965.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_1967 ({sk[695], i_29_, i_37_, n_n793, n_n1404, n_n1397, x376x}, x1733x);
	defparam lut_1967.LUT_SIZE = 7;
	defparam lut_1967.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_1969 ({sk[696], i_28_, i_33_, i_29_, n_n1429, x376x, x6929x}, x1738x);
	defparam lut_1969.LUT_SIZE = 7;
	defparam lut_1969.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_1971 ({sk[697], i_34_, i_37_, x601x, x1732x, x1733x, x1738x}, x6934x);
	defparam lut_1971.LUT_SIZE = 7;
	defparam lut_1971.mask = 128'h57ffffff57ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_1976 ({sk[698], i_9_, i_7_, i_8_, i_6_}, x6876x);
	defparam lut_1976.LUT_SIZE = 5;
	defparam lut_1976.mask = 32'h77778000;

	lut_sub lut_1978 ({sk[699], i_34_, i_33_, i_35_, i_37_}, x246x);
	defparam lut_1978.LUT_SIZE = 5;
	defparam lut_1978.mask = 32'h77771000;

	lut_sub lut_1980 ({sk[700], i_20_, i_27_, i_26_, i_23_, i_24_}, x6886x);
	defparam lut_1980.LUT_SIZE = 6;
	defparam lut_1980.mask = 64'h3f3fffff80000000;

	lut_sub lut_1982 ({sk[701], i_14_, i_16_, i_37_}, x268x);
	defparam lut_1982.LUT_SIZE = 4;
	defparam lut_1982.mask = 16'h5540;

	lut_sub lut_1984 ({sk[702], i_9_, i_6_, i_11_, i_19_}, x361x);
	defparam lut_1984.LUT_SIZE = 5;
	defparam lut_1984.mask = 32'h77778000;

	lut_sub lut_1986 ({sk[703], i_13_, i_17_, i_16_, i_33_, i_35_, i_37_}, x461x);
	defparam lut_1986.LUT_SIZE = 7;
	defparam lut_1986.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_1988 ({sk[704], i_9_, i_8_, i_5_, i_6_, i_4_, i_0_}, x487x);
	defparam lut_1988.LUT_SIZE = 7;
	defparam lut_1988.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_1990 ({sk[705], i_20_, i_23_, i_24_}, x6899x);
	defparam lut_1990.LUT_SIZE = 4;
	defparam lut_1990.mask = 16'h5580;

	lut_sub lut_1992 ({sk[706], i_7_, i_8_, i_6_, n_n245, x44x, x6899x}, x508x);
	defparam lut_1992.LUT_SIZE = 7;
	defparam lut_1992.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_1994 ({sk[707], i_7_, i_8_, i_12_, i_21_, i_36_}, x7977x);
	defparam lut_1994.LUT_SIZE = 6;
	defparam lut_1994.mask = 64'h3f3fffff40000000;

	lut_sub lut_1996 ({sk[708], i_30_, i_28_, i_23_, i_21_, i_16_, i_32_}, x7975x);
	defparam lut_1996.LUT_SIZE = 7;
	defparam lut_1996.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_1998 ({sk[709], i_10_, i_7_, i_14_, i_13_, i_17_, i_16_}, x325x);
	defparam lut_1998.LUT_SIZE = 7;
	defparam lut_1998.mask = 128'h57ffffff57ffffff0000000000000800;

	lut_sub lut_2000 ({sk[710], i_10_, i_7_, i_14_, i_13_, i_12_, i_16_}, x328x);
	defparam lut_2000.LUT_SIZE = 7;
	defparam lut_2000.mask = 128'h57ffffff57ffffff0000000000000800;

	lut_sub lut_2002 ({sk[711], i_32_, i_31_, i_33_, i_35_, i_38_}, n_n1149);
	defparam lut_2002.LUT_SIZE = 6;
	defparam lut_2002.mask = 64'h3f3fffff40000000;

	lut_sub lut_2004 ({sk[712], i_28_, i_24_, i_34_, i_29_}, x447x);
	defparam lut_2004.LUT_SIZE = 5;
	defparam lut_2004.mask = 32'h77772000;

	lut_sub lut_2006 ({sk[713], i_18_, x204x, n_n1278, x14x, x388x, x404x}, x1405x);
	defparam lut_2006.LUT_SIZE = 7;
	defparam lut_2006.mask = 128'h57ffffff57ffffff0011031300000303;

	lut_sub lut_2009 ({sk[714], i_18_, i_24_, x204x, n_n1278, x14x, x404x}, x26x);
	defparam lut_2009.LUT_SIZE = 7;
	defparam lut_2009.mask = 128'h57ffffff57ffffff0537000000330000;

	lut_sub lut_2012 ({sk[715], i_25_, i_34_, i_38_, x42x, x1405x, x26x}, x611x);
	defparam lut_2012.LUT_SIZE = 7;
	defparam lut_2012.mask = 128'h57ffffff57ffffff3333333733333333;

	lut_sub lut_2015 ({sk[716], i_9_, i_8_, i_5_, i_6_, i_3_, i_11_}, x7416x);
	defparam lut_2015.LUT_SIZE = 7;
	defparam lut_2015.mask = 128'h57ffffff57ffffff0000000040000000;

	lut_sub lut_2017 ({sk[717], i_9_, i_8_, i_13_, i_11_, i_18_}, x7418x);
	defparam lut_2017.LUT_SIZE = 6;
	defparam lut_2017.mask = 64'h3f3fffff00001000;

	lut_sub lut_2019 ({sk[718], i_13_, i_12_, x292x, x11x, x7416x, x7418x}, x21x);
	defparam lut_2019.LUT_SIZE = 7;
	defparam lut_2019.mask = 128'h57ffffff57ffffff0537050505050505;

	lut_sub lut_2022 ({sk[719], i_9_, i_8_, i_13_, i_18_, x208x, x50x}, x28x);
	defparam lut_2022.LUT_SIZE = 7;
	defparam lut_2022.mask = 128'h57ffffff57ffffff0000000037000500;

	lut_sub lut_2025 ({sk[720], i_30_, i_8_, i_28_, i_31_}, x7466x);
	defparam lut_2025.LUT_SIZE = 5;
	defparam lut_2025.mask = 32'h77778000;

	lut_sub lut_2027 ({sk[721], i_25_, i_24_, i_19_, i_35_, i_38_}, x371x);
	defparam lut_2027.LUT_SIZE = 6;
	defparam lut_2027.mask = 64'h3f3fffff04000000;

	lut_sub lut_2029 ({sk[722], i_10_, i_8_, n_n1345, x389x, x210x, x807x}, x1265x);
	defparam lut_2029.LUT_SIZE = 7;
	defparam lut_2029.mask = 128'h57ffffff57ffffff0003000000070000;

	lut_sub lut_2032 ({sk[723], x11x, x288x, x12x, x7415x, x7416x, x7418x}, x1266x);
	defparam lut_2032.LUT_SIZE = 7;
	defparam lut_2032.mask = 128'h57ffffff57ffffff0000000300000057;

	lut_sub lut_2035 ({sk[724], i_9_, i_19_, n_n1118, x213x, x288x, x12x}, x1267x);
	defparam lut_2035.LUT_SIZE = 7;
	defparam lut_2035.mask = 128'h57ffffff57ffffff0000000000000001;

	lut_sub lut_2037 ({sk[725], i_30_, i_28_, i_32_, i_31_, i_34_, i_29_}, x616x);
	defparam lut_2037.LUT_SIZE = 7;
	defparam lut_2037.mask = 128'h57ffffff57ffffff0222000022220000;

	lut_sub lut_2041 ({sk[726], i_14_, i_13_, i_12_, i_24_, i_17_}, x614x);
	defparam lut_2041.LUT_SIZE = 6;
	defparam lut_2041.mask = 64'h3f3fffff040404cc;

	lut_sub lut_2044 ({sk[727], i_14_, i_13_, i_12_, i_17_, i_29_}, x7623x);
	defparam lut_2044.LUT_SIZE = 6;
	defparam lut_2044.mask = 64'h3f3fffff01010155;

	lut_sub lut_2047 ({sk[728], i_28_, i_21_, i_22_, i_34_, i_35_, i_29_}, x1106x);
	defparam lut_2047.LUT_SIZE = 7;
	defparam lut_2047.mask = 128'h57ffffff57ffffff0000100000000000;

	lut_sub lut_2049 ({sk[729], i_22_, n_n1497, x616x, x614x, x7623x, x1106x}, n_n1892);
	defparam lut_2049.LUT_SIZE = 7;
	defparam lut_2049.mask = 128'h57ffffff57ffffff555f777f555f555f;

	lut_sub lut_2053 ({sk[730], i_30_, i_27_, i_16_, i_32_}, x35x);
	defparam lut_2053.LUT_SIZE = 5;
	defparam lut_2053.mask = 32'h7777151f;

	lut_sub lut_2057 ({sk[731], i_30_, i_14_, i_16_, i_34_, i_33_}, x620x);
	defparam lut_2057.LUT_SIZE = 6;
	defparam lut_2057.mask = 64'h3f3fffff00110313;

	lut_sub lut_2060 ({sk[732], i_27_, i_28_, i_16_, i_22_, n_n1334, x620x}, x619x);
	defparam lut_2060.LUT_SIZE = 7;
	defparam lut_2060.mask = 128'h57ffffff57ffffff0507000007070000;

	lut_sub lut_2064 ({sk[733], i_30_, i_27_, i_23_, i_16_, i_32_}, x618x);
	defparam lut_2064.LUT_SIZE = 6;
	defparam lut_2064.mask = 64'h3f3fffff15553fff;

	lut_sub lut_2071 ({sk[734], i_28_, i_22_, x298x, n_n1519, x35x, x7627x}, x7631x);
	defparam lut_2071.LUT_SIZE = 7;
	defparam lut_2071.mask = 128'h57ffffff57ffffff0505053705050505;

	lut_sub lut_2074 ({sk[735], i_28_, i_31_, i_29_, n_n1397, n_n1251, x618x}, x7632x);
	defparam lut_2074.LUT_SIZE = 7;
	defparam lut_2074.mask = 128'h57ffffff57ffffff05000d0000000000;

	lut_sub lut_2077 ({sk[736], i_24_, n_n1892, x619x, x7631x, x7632x}, n_n1837);
	defparam lut_2077.LUT_SIZE = 6;
	defparam lut_2077.mask = 64'h3f3fffff7fff77ff;

	lut_sub lut_2082 ({sk[737], i_28_, i_25_, i_26_, i_38_}, x311x);
	defparam lut_2082.LUT_SIZE = 5;
	defparam lut_2082.mask = 32'h77774000;

	lut_sub lut_2084 ({sk[738], i_28_, i_25_, i_26_, i_22_}, x78x);
	defparam lut_2084.LUT_SIZE = 5;
	defparam lut_2084.mask = 32'h77778000;

	lut_sub lut_2086 ({sk[739], i_30_, i_7_, i_8_, i_24_, i_38_}, x7292x);
	defparam lut_2086.LUT_SIZE = 6;
	defparam lut_2086.mask = 64'h3f3fffff40000000;

	lut_sub lut_2088 ({sk[740], i_28_, i_32_, i_33_, i_29_}, x344x);
	defparam lut_2088.LUT_SIZE = 5;
	defparam lut_2088.mask = 32'h77778000;

	lut_sub lut_2090 ({sk[741], i_9_, i_5_, i_6_, i_18_}, x353x);
	defparam lut_2090.LUT_SIZE = 5;
	defparam lut_2090.mask = 32'h77778000;

	lut_sub lut_2092 ({sk[742], n_n1307, n_n787, x239x, n_n1422, x361x, x353x}, x1422x);
	defparam lut_2092.LUT_SIZE = 7;
	defparam lut_2092.mask = 128'h57ffffff57ffffff0000000500030007;

	lut_sub lut_2095 ({sk[743], i_9_, i_2_, n_n1431, x23x, x81x, x1378x}, x1372x);
	defparam lut_2095.LUT_SIZE = 7;
	defparam lut_2095.mask = 128'h57ffffff57ffffff0011000000130000;

	lut_sub lut_2098 ({sk[744], i_10_, i_25_, i_32_, x42x, x14x, n_n1419}, x1373x);
	defparam lut_2098.LUT_SIZE = 7;
	defparam lut_2098.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2100 ({sk[745], i_10_, i_28_, i_32_, i_29_, x229x, x238x}, x1374x);
	defparam lut_2100.LUT_SIZE = 7;
	defparam lut_2100.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_2102 ({sk[746], i_9_, i_10_, i_24_, x11x, n_n1179, x78x}, x1375x);
	defparam lut_2102.LUT_SIZE = 7;
	defparam lut_2102.mask = 128'h57ffffff57ffffff0000000001000000;

	lut_sub lut_2104 ({sk[747], i_9_, i_38_, x204x, n_n1454, x42x, x376x}, x1376x);
	defparam lut_2104.LUT_SIZE = 7;
	defparam lut_2104.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_2106 ({sk[748], i_28_, i_13_, i_31_, x389x, x41x}, x1377x);
	defparam lut_2106.LUT_SIZE = 6;
	defparam lut_2106.mask = 64'h3f3fffff00100000;

	lut_sub lut_2108 ({sk[749], i_9_, i_8_, i_18_, n_n1278, n_n787, x456x}, x1370x);
	defparam lut_2108.LUT_SIZE = 7;
	defparam lut_2108.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2110 ({sk[750], i_9_, i_13_, i_38_, n_n1397, n_n1302, x376x}, x1371x);
	defparam lut_2110.LUT_SIZE = 7;
	defparam lut_2110.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_2112 ({sk[751], i_9_, i_10_, i_24_, n_n805, x50x, n_n1302}, x1366x);
	defparam lut_2112.LUT_SIZE = 7;
	defparam lut_2112.mask = 128'h57ffffff57ffffff0000000001000000;

	lut_sub lut_2114 ({sk[752], i_24_, i_22_, x58x, n_n1353, n_n1197, x11x}, x1369x);
	defparam lut_2114.LUT_SIZE = 7;
	defparam lut_2114.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_2116 ({sk[753], i_13_, x518x, n_n1128, x41x, x226x, x238x}, x7366x);
	defparam lut_2116.LUT_SIZE = 7;
	defparam lut_2116.mask = 128'h57ffffff57ffffff0000030300050307;

	lut_sub lut_2119 ({sk[754], i_25_, i_24_, i_34_, i_35_, i_38_}, x238x);
	defparam lut_2119.LUT_SIZE = 6;
	defparam lut_2119.mask = 64'h3f3fffff04000000;

	lut_sub lut_2121 ({sk[755], i_28_, i_25_, i_24_, i_34_, i_35_, i_38_}, x315x);
	defparam lut_2121.LUT_SIZE = 7;
	defparam lut_2121.mask = 128'h57ffffff57ffffff0400000000000000;

	lut_sub lut_2123 ({sk[756], i_28_, i_34_, i_33_, i_35_, i_38_, i_29_}, x387x);
	defparam lut_2123.LUT_SIZE = 7;
	defparam lut_2123.mask = 128'h57ffffff57ffffff0200000000000000;

	lut_sub lut_2125 ({sk[757], i_9_, i_8_, i_11_, i_2_, i_18_}, x1388x);
	defparam lut_2125.LUT_SIZE = 6;
	defparam lut_2125.mask = 64'h3f3fffff00000400;

	lut_sub lut_2127 ({sk[758], i_9_, i_8_, i_3_, i_2_, i_19_}, x1389x);
	defparam lut_2127.LUT_SIZE = 6;
	defparam lut_2127.mask = 64'h3f3fffff00004000;

	lut_sub lut_2129 ({sk[759], i_9_, i_8_, i_3_, i_13_, i_11_, i_2_}, x1361x);
	defparam lut_2129.LUT_SIZE = 7;
	defparam lut_2129.mask = 128'h57ffffff57ffffff0000000020000000;

	lut_sub lut_2131 ({sk[760], i_9_, i_8_, i_13_, i_2_, i_18_, i_19_}, x1363x);
	defparam lut_2131.LUT_SIZE = 7;
	defparam lut_2131.mask = 128'h57ffffff57ffffff0000000010000000;

	lut_sub lut_2133 ({sk[761], i_13_, x1388x, x1389x, x1361x, x1363x}, x625x);
	defparam lut_2133.LUT_SIZE = 6;
	defparam lut_2133.mask = 64'h3f3fffff7fff7777;

	lut_sub lut_2138 ({sk[762], i_28_, i_26_, i_24_, i_29_, n_n1353, x11x}, x1352x);
	defparam lut_2138.LUT_SIZE = 7;
	defparam lut_2138.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_2140 ({sk[763], i_9_, i_10_, i_26_, i_24_, x11x, n_n1288}, x1350x);
	defparam lut_2140.LUT_SIZE = 7;
	defparam lut_2140.mask = 128'h57ffffff57ffffff0000000010000000;

	lut_sub lut_2142 ({sk[764], n_n1133, n_n1128, x41x, n_n1497, x207x, x7388x}, x7392x);
	defparam lut_2142.LUT_SIZE = 7;
	defparam lut_2142.mask = 128'h57ffffff57ffffff0000005503030357;

	lut_sub lut_2145 ({sk[765], i_28_, i_25_, i_26_, i_35_, i_38_, i_29_}, x7386x);
	defparam lut_2145.LUT_SIZE = 7;
	defparam lut_2145.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_2147 ({sk[766], i_9_, i_10_, i_24_, x11x, n_n1179, x71x}, x1348x);
	defparam lut_2147.LUT_SIZE = 7;
	defparam lut_2147.mask = 128'h57ffffff57ffffff0000000001000000;

	lut_sub lut_2149 ({sk[767], n_n1133, n_n1128, x509x, x207x, x218x, x270x}, x7394x);
	defparam lut_2149.LUT_SIZE = 7;
	defparam lut_2149.mask = 128'h57ffffff57ffffff0000050500330537;

	lut_sub lut_2152 ({sk[768], i_9_, i_8_, i_3_, i_13_, i_11_, i_18_}, x425x);
	defparam lut_2152.LUT_SIZE = 7;
	defparam lut_2152.mask = 128'h57ffffff57ffffff0000000030100000;

	lut_sub lut_2155 ({sk[769], i_9_, i_8_, i_3_, i_13_, i_18_, i_19_}, x454x);
	defparam lut_2155.LUT_SIZE = 7;
	defparam lut_2155.mask = 128'h57ffffff57ffffff0000000050100000;

	lut_sub lut_2158 ({sk[770], i_9_, i_3_, i_13_, i_11_, i_18_}, x785x);
	defparam lut_2158.LUT_SIZE = 6;
	defparam lut_2158.mask = 64'h3f3fffff00003010;

	lut_sub lut_2161 ({sk[771], i_25_, i_24_, i_32_, i_34_, i_35_, i_38_}, x7398x);
	defparam lut_2161.LUT_SIZE = 7;
	defparam lut_2161.mask = 128'h57ffffff57ffffff0400000000000000;

	lut_sub lut_2163 ({sk[772], i_24_, i_34_, i_33_, i_35_, i_38_}, x7399x);
	defparam lut_2163.LUT_SIZE = 6;
	defparam lut_2163.mask = 64'h3f3fffff00400000;

	lut_sub lut_2165 ({sk[773], n_n1489, x425x, x454x, x785x, x7398x, x7399x}, x1335x);
	defparam lut_2165.LUT_SIZE = 7;
	defparam lut_2165.mask = 128'h57ffffff57ffffff0000000003575757;

	lut_sub lut_2169 ({sk[774], i_25_, i_32_, i_38_, x58x, x14x, n_n1191}, x1334x);
	defparam lut_2169.LUT_SIZE = 7;
	defparam lut_2169.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_2171 ({sk[775], i_13_, i_32_, x14x, x70x}, x1337x);
	defparam lut_2171.LUT_SIZE = 5;
	defparam lut_2171.mask = 32'h77770010;

	lut_sub lut_2173 ({sk[776], i_28_, i_25_, i_34_, i_35_, i_38_, i_29_}, x271x);
	defparam lut_2173.LUT_SIZE = 7;
	defparam lut_2173.mask = 128'h57ffffff57ffffff0020000000000000;

	lut_sub lut_2175 ({sk[777], i_9_, i_3_, i_13_, i_18_}, x18x);
	defparam lut_2175.LUT_SIZE = 5;
	defparam lut_2175.mask = 32'h777700c4;

	lut_sub lut_2178 ({sk[778], i_25_, i_24_, i_19_, n_n1489, n_n1422, x18x}, x1330x);
	defparam lut_2178.LUT_SIZE = 7;
	defparam lut_2178.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_2180 ({sk[779], i_14_, i_35_, i_37_}, x416x);
	defparam lut_2180.LUT_SIZE = 4;
	defparam lut_2180.mask = 16'h5540;

	lut_sub lut_2182 ({sk[780], i_14_, i_12_, i_17_, i_16_}, x629x);
	defparam lut_2182.LUT_SIZE = 5;
	defparam lut_2182.mask = 32'h7777a800;

	lut_sub lut_2185 ({sk[781], x54x, n_n1489, n_n1438, x6971x, x6967x, x6970x}, x1716x);
	defparam lut_2185.LUT_SIZE = 7;
	defparam lut_2185.mask = 128'h57ffffff57ffffff0005000500050307;

	lut_sub lut_2188 ({sk[782], i_17_, x43x, n_n1396, n_n1406, x245x, x6958x}, x1720x);
	defparam lut_2188.LUT_SIZE = 7;
	defparam lut_2188.mask = 128'h57ffffff57ffffff0000035700000000;

	lut_sub lut_2191 ({sk[783], n_n1375, x302x, n_n1489, n_n1334, x6966x, x6972x}, x6974x);
	defparam lut_2191.LUT_SIZE = 7;
	defparam lut_2191.mask = 128'h57ffffff57ffffff0000003305050537;

	lut_sub lut_2194 ({sk[784], n_n1274, n_n1326, x45x, x6947x, x629x, x6973x}, x6975x);
	defparam lut_2194.LUT_SIZE = 7;
	defparam lut_2194.mask = 128'h57ffffff57ffffff0000030300550357;

	lut_sub lut_2197 ({sk[785], x1716x, x1720x, x6974x, x6975x}, n_n1719);
	defparam lut_2197.LUT_SIZE = 5;
	defparam lut_2197.mask = 32'h77777fff;

	lut_sub lut_2202 ({sk[786], i_14_, i_17_, i_16_, i_32_, i_35_, i_37_}, x303x);
	defparam lut_2202.LUT_SIZE = 7;
	defparam lut_2202.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_2204 ({sk[787], i_9_, i_10_, i_6_, i_13_}, x635x);
	defparam lut_2204.LUT_SIZE = 5;
	defparam lut_2204.mask = 32'h7777c400;

	lut_sub lut_2207 ({sk[788], n_n1443, n_n1307, n_n504, x50x, x303x, x635x}, x633x);
	defparam lut_2207.LUT_SIZE = 7;
	defparam lut_2207.mask = 128'h57ffffff57ffffff00001111000f111f;

	lut_sub lut_2210 ({sk[789], i_27_, i_28_, i_23_, i_24_, i_33_, i_29_}, x6937x);
	defparam lut_2210.LUT_SIZE = 7;
	defparam lut_2210.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_2212 ({sk[790], i_27_, i_28_, i_24_, i_32_, i_33_, i_29_}, x6938x);
	defparam lut_2212.LUT_SIZE = 7;
	defparam lut_2212.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_2214 ({sk[791], n_n1443, x51x, x50x, x6920x, x6937x, x6938x}, x632x);
	defparam lut_2214.LUT_SIZE = 7;
	defparam lut_2214.mask = 128'h57ffffff57ffffff0000050500330537;

	lut_sub lut_2217 ({sk[792], i_17_, i_29_, n_n1441, x54x, x41x, x6935x}, x1723x);
	defparam lut_2217.LUT_SIZE = 7;
	defparam lut_2217.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_2219 ({sk[793], i_12_, i_29_, n_n793, x43x, x376x, x246x}, x1724x);
	defparam lut_2219.LUT_SIZE = 7;
	defparam lut_2219.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_2221 ({sk[794], i_23_, x43x, x321x, x492x, x1723x, x1724x}, x6942x);
	defparam lut_2221.LUT_SIZE = 7;
	defparam lut_2221.mask = 128'h57ffffff57ffffff7777777f77777777;

	lut_sub lut_2225 ({sk[795], i_34_, i_35_, i_37_, x67x, x633x, x632x}, x6943x);
	defparam lut_2225.LUT_SIZE = 7;
	defparam lut_2225.mask = 128'h57ffffff57ffffff0303030303570303;

	lut_sub lut_2228 ({sk[796], i_8_, i_18_, i_17_, i_16_}, x413x);
	defparam lut_2228.LUT_SIZE = 5;
	defparam lut_2228.mask = 32'h77778000;

	lut_sub lut_2230 ({sk[797], i_9_, n_n1278, n_n787, x376x, x431x, x413x}, x31x);
	defparam lut_2230.LUT_SIZE = 7;
	defparam lut_2230.mask = 128'h57ffffff57ffffff0303035700000000;

	lut_sub lut_2233 ({sk[798], i_11_, i_23_, i_17_, i_19_, x14x, x268x}, x351x);
	defparam lut_2233.LUT_SIZE = 7;
	defparam lut_2233.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_2235 ({sk[799], i_11_, i_23_, i_17_, i_19_}, x7121x);
	defparam lut_2235.LUT_SIZE = 5;
	defparam lut_2235.mask = 32'h77778000;

	lut_sub lut_2237 ({sk[800], i_14_, i_23_, i_18_, i_17_, i_16_, i_37_}, x7124x);
	defparam lut_2237.LUT_SIZE = 7;
	defparam lut_2237.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_2239 ({sk[801], n_n1278, x14x, x404x, x268x, x7121x, x7124x}, x637x);
	defparam lut_2239.LUT_SIZE = 7;
	defparam lut_2239.mask = 128'h57ffffff57ffffff0000030300550357;

	lut_sub lut_2242 ({sk[802], i_14_, i_13_, i_37_}, x7128x);
	defparam lut_2242.LUT_SIZE = 4;
	defparam lut_2242.mask = 16'h5510;

	lut_sub lut_2244 ({sk[803], i_20_, i_17_, i_16_, x46x, x6876x, x7128x}, x1568x);
	defparam lut_2244.LUT_SIZE = 7;
	defparam lut_2244.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2246 ({sk[804], i_28_, i_32_, i_29_, i_37_, n_n916, x7129x}, x1570x);
	defparam lut_2246.LUT_SIZE = 7;
	defparam lut_2246.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_2248 ({sk[805], x59x, n_n301, n_n460, x45x, x7129x, x7131x}, x1571x);
	defparam lut_2248.LUT_SIZE = 7;
	defparam lut_2248.mask = 128'h57ffffff57ffffff0000050500000537;

	lut_sub lut_2251 ({sk[806], i_20_, i_23_, i_17_, x1568x, x1570x, x1571x}, x636x);
	defparam lut_2251.LUT_SIZE = 7;
	defparam lut_2251.mask = 128'h57ffffff57ffffff7f0f0f0f0f0f0f0f;

	lut_sub lut_2255 ({sk[807], i_20_, x54x, n_n245, x461x, x44x, x7119x}, x1564x);
	defparam lut_2255.LUT_SIZE = 7;
	defparam lut_2255.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_2257 ({sk[808], i_14_, i_34_, i_35_, i_29_, i_37_, n_n793}, x7126x);
	defparam lut_2257.LUT_SIZE = 7;
	defparam lut_2257.mask = 128'h57ffffff57ffffff0010000000000000;

	lut_sub lut_2259 ({sk[809], n_n1375, n_n1202, x31x, x637x, x1564x, x7126x}, x7133x);
	defparam lut_2259.LUT_SIZE = 7;
	defparam lut_2259.mask = 128'h57ffffff57ffffff3377337733773f7f;

	lut_sub lut_2263 ({sk[810], i_25_, i_34_, i_33_, n_n1375, x54x, n_n1404}, x1703x);
	defparam lut_2263.LUT_SIZE = 7;
	defparam lut_2263.mask = 128'h57ffffff57ffffff0000000000000001;

	lut_sub lut_2265 ({sk[811], i_31_, i_34_, n_n1375, x513x, x6978x, x6980x}, x6985x);
	defparam lut_2265.LUT_SIZE = 7;
	defparam lut_2265.mask = 128'h57ffffff57ffffff0303030303030357;

	lut_sub lut_2268 ({sk[812], i_35_, i_37_, n_n1340, x48x, x419x, x6981x}, x6986x);
	defparam lut_2268.LUT_SIZE = 7;
	defparam lut_2268.mask = 128'h57ffffff57ffffff0505053705050505;

	lut_sub lut_2271 ({sk[813], i_21_, x54x, n_n1429, n_n1326, x6947x, x398x}, x6987x);
	defparam lut_2271.LUT_SIZE = 7;
	defparam lut_2271.mask = 128'h57ffffff57ffffff0003000300035557;

	lut_sub lut_2274 ({sk[814], i_29_, x302x, n_n1489, x441x, x416x, x6983x}, x6988x);
	defparam lut_2274.LUT_SIZE = 7;
	defparam lut_2274.mask = 128'h57ffffff57ffffff0011001100110f1f;

	lut_sub lut_2277 ({sk[815], x1703x, x6985x, x6986x, x6987x, x6988x}, n_n1720);
	defparam lut_2277.LUT_SIZE = 6;
	defparam lut_2277.mask = 64'h3f3fffff7fffffff;

	lut_sub lut_2283 ({sk[816], i_8_, n_n1441, x10x, x74x, x342x, x6994x}, x1687x);
	defparam lut_2283.LUT_SIZE = 7;
	defparam lut_2283.mask = 128'h57ffffff57ffffff0005111500001111;

	lut_sub lut_2286 ({sk[817], i_7_, x10x, n_n1499, x318x, x661x, x6995x}, x1688x);
	defparam lut_2286.LUT_SIZE = 7;
	defparam lut_2286.mask = 128'h57ffffff57ffffff001100110011001f;

	lut_sub lut_2289 ({sk[818], i_20_, x54x, n_n1404, x47x, x485x, x6999x}, x1689x);
	defparam lut_2289.LUT_SIZE = 7;
	defparam lut_2289.mask = 128'h57ffffff57ffffff0005000500050037;

	lut_sub lut_2292 ({sk[819], i_17_, i_34_, i_33_, n_n1375, x43x, n_n1396}, x1691x);
	defparam lut_2292.LUT_SIZE = 7;
	defparam lut_2292.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_2294 ({sk[820], n_n1429, x432x, x1687x, x1688x, x1689x, x1691x}, n_n1716);
	defparam lut_2294.LUT_SIZE = 7;
	defparam lut_2294.mask = 128'h57ffffff57ffffff7fff7fff7fffffff;

	lut_sub lut_2300 ({sk[821], i_8_, n_n1375, x10x, x48x, x342x, x7004x}, x1679x);
	defparam lut_2300.LUT_SIZE = 7;
	defparam lut_2300.mask = 128'h57ffffff57ffffff0005111500001111;

	lut_sub lut_2303 ({sk[822], i_35_, n_n1375, n_n1429, n_n1326, n_n1080, x6944x}, x1682x);
	defparam lut_2303.LUT_SIZE = 7;
	defparam lut_2303.mask = 128'h57ffffff57ffffff0000005500030057;

	lut_sub lut_2306 ({sk[823], i_27_, i_23_, i_21_, i_35_, n_n1443, n_n1326}, x1684x);
	defparam lut_2306.LUT_SIZE = 7;
	defparam lut_2306.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_2308 ({sk[824], x57x, x67x, x316x, x7006x, x7005x, x7007x}, x7010x);
	defparam lut_2308.LUT_SIZE = 7;
	defparam lut_2308.mask = 128'h57ffffff57ffffff0000050500330537;

	lut_sub lut_2311 ({sk[825], n_n1404, x432x, x1679x, x1682x, x1684x, x7010x}, n_n1715);
	defparam lut_2311.LUT_SIZE = 7;
	defparam lut_2311.mask = 128'h57ffffff57ffffff7fff7fff7fffffff;

	lut_sub lut_2317 ({sk[826], i_20_, i_7_, i_13_, i_12_, i_16_}, x401x);
	defparam lut_2317.LUT_SIZE = 6;
	defparam lut_2317.mask = 64'h3f3fffff00000080;

	lut_sub lut_2319 ({sk[827], i_27_, i_28_, i_25_, i_34_, i_33_}, x485x);
	defparam lut_2319.LUT_SIZE = 6;
	defparam lut_2319.mask = 64'h3f3fffff01000000;

	lut_sub lut_2321 ({sk[828], i_27_, i_28_, i_25_, i_33_, i_29_}, x6999x);
	defparam lut_2321.LUT_SIZE = 6;
	defparam lut_2321.mask = 64'h3f3fffff02000000;

	lut_sub lut_2323 ({sk[829], i_20_, i_23_, i_24_, n_n1397, x485x, x6999x}, x640x);
	defparam lut_2323.LUT_SIZE = 7;
	defparam lut_2323.mask = 128'h57ffffff57ffffff0505000037050000;

	lut_sub lut_2326 ({sk[830], i_20_, i_28_, i_25_, x479x, x84x, x94x}, x1670x);
	defparam lut_2326.LUT_SIZE = 7;
	defparam lut_2326.mask = 128'h57ffffff57ffffff00000000111f1111;

	lut_sub lut_2329 ({sk[831], i_7_, x43x, n_n1499, x318x, x7014x, x7015x}, x7018x);
	defparam lut_2329.LUT_SIZE = 7;
	defparam lut_2329.mask = 128'h57ffffff57ffffff111111111111111f;

	lut_sub lut_2332 ({sk[832], i_12_, x10x, n_n1406, x245x, x84x, x401x}, x7019x);
	defparam lut_2332.LUT_SIZE = 7;
	defparam lut_2332.mask = 128'h57ffffff57ffffff1111111f11111111;

	lut_sub lut_2335 ({sk[833], i_17_, x10x, x640x, x1670x, x7018x, x7019x}, x7022x);
	defparam lut_2335.LUT_SIZE = 7;
	defparam lut_2335.mask = 128'h57ffffff57ffffff7f7f7fff7f7f7f7f;

	lut_sub lut_2340 ({sk[834], i_7_, i_17_, i_31_, n_n1441, x43x, x54x}, x1659x);
	defparam lut_2340.LUT_SIZE = 7;
	defparam lut_2340.mask = 128'h57ffffff57ffffff0000000000010000;

	lut_sub lut_2342 ({sk[835], i_22_, n_n1443, n_n1429, x308x, x1659x, x803x}, n_n1723);
	defparam lut_2342.LUT_SIZE = 7;
	defparam lut_2342.mask = 128'h57ffffff57ffffff333f3f3f777f7f7f;

	lut_sub lut_2347 ({sk[836], i_23_, i_21_, i_22_}, x7033x);
	defparam lut_2347.LUT_SIZE = 4;
	defparam lut_2347.mask = 16'h5520;

	lut_sub lut_2349 ({sk[837], i_14_, i_12_, i_17_, i_16_}, x716x);
	defparam lut_2349.LUT_SIZE = 5;
	defparam lut_2349.mask = 32'h7777a800;

	lut_sub lut_2352 ({sk[838], n_n1443, n_n1396, x6958x, x45x, x7033x, x716x}, x7036x);
	defparam lut_2352.LUT_SIZE = 7;
	defparam lut_2352.mask = 128'h57ffffff57ffffff0000005503030357;

	lut_sub lut_2355 ({sk[839], i_27_, i_23_, i_21_, i_22_, x73x, n_n1368}, x55x);
	defparam lut_2355.LUT_SIZE = 7;
	defparam lut_2355.mask = 128'h57ffffff57ffffff0010000000000000;

	lut_sub lut_2357 ({sk[840], x104x, x7036x, x7034x, x7035x, x7039x, x7040x}, x7043x);
	defparam lut_2357.LUT_SIZE = 7;
	defparam lut_2357.mask = 128'h57ffffff57ffffff7fffffffffffffff;

	lut_sub lut_2364 ({sk[841], i_30_, i_28_, i_22_, i_32_, x298x, n_n1497}, x646x);
	defparam lut_2364.LUT_SIZE = 7;
	defparam lut_2364.mask = 128'h57ffffff57ffffff0537050555775555;

	lut_sub lut_2368 ({sk[842], i_30_, i_27_, i_16_, i_31_, i_34_}, x645x);
	defparam lut_2368.LUT_SIZE = 6;
	defparam lut_2368.mask = 64'h3f3fffff01110515;

	lut_sub lut_2372 ({sk[843], i_28_, i_24_, i_34_, i_29_, x35x, x645x}, x7635x);
	defparam lut_2372.LUT_SIZE = 7;
	defparam lut_2372.mask = 128'h57ffffff57ffffff5070000000000000;

	lut_sub lut_2375 ({sk[844], i_30_, i_27_, i_14_, i_16_, i_32_, i_33_}, x7637x);
	defparam lut_2375.LUT_SIZE = 7;
	defparam lut_2375.mask = 128'h57ffffff57ffffff035733770f5fffff;

	lut_sub lut_2381 ({sk[845], i_23_, i_31_, n_n1497, x103x, x447x, x7637x}, n_n1897);
	defparam lut_2381.LUT_SIZE = 7;
	defparam lut_2381.mask = 128'h57ffffff57ffffff0055005f337733ff;

	lut_sub lut_2386 ({sk[846], i_32_, i_33_, i_35_, i_38_, i_29_}, x7444x);
	defparam lut_2386.LUT_SIZE = 6;
	defparam lut_2386.mask = 64'h3f3fffff20000000;

	lut_sub lut_2388 ({sk[847], i_25_, i_32_, i_35_, i_38_, x73x, x42x}, x381x);
	defparam lut_2388.LUT_SIZE = 7;
	defparam lut_2388.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2390 ({sk[848], i_9_, i_19_, n_n1118, n_n1048, x76x, x213x}, x1293x);
	defparam lut_2390.LUT_SIZE = 7;
	defparam lut_2390.mask = 128'h57ffffff57ffffff0000030300000357;

	lut_sub lut_2393 ({sk[849], i_13_, i_12_, x292x, x11x, x7416x, x7418x}, x7442x);
	defparam lut_2393.LUT_SIZE = 7;
	defparam lut_2393.mask = 128'h57ffffff57ffffff0537050505050505;

	lut_sub lut_2396 ({sk[850], i_26_, i_24_, i_33_, i_35_, i_38_, x42x}, x7443x);
	defparam lut_2396.LUT_SIZE = 7;
	defparam lut_2396.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_2398 ({sk[851], x11x, x213x, x7423x, n_n1497, x7424x, x7444x}, x1292x);
	defparam lut_2398.LUT_SIZE = 7;
	defparam lut_2398.mask = 128'h57ffffff57ffffff0000010100050105;

	lut_sub lut_2401 ({sk[852], i_28_, i_26_, i_24_, i_22_, i_38_}, x7449x);
	defparam lut_2401.LUT_SIZE = 6;
	defparam lut_2401.mask = 64'h3f3fffff40000000;

	lut_sub lut_2403 ({sk[853], n_n1307, n_n787, n_n1458, x361x, x353x, x7449x}, x1288x);
	defparam lut_2403.LUT_SIZE = 7;
	defparam lut_2403.mask = 128'h57ffffff57ffffff0000001100050015;

	lut_sub lut_2406 ({sk[854], x204x, x61x, x404x, x41x, x226x, x7274x}, x1284x);
	defparam lut_2406.LUT_SIZE = 7;
	defparam lut_2406.mask = 128'h57ffffff57ffffff0000001100000313;

	lut_sub lut_2409 ({sk[855], i_25_, i_18_, n_n1278, n_n1288, n_n1419, x404x}, x1285x);
	defparam lut_2409.LUT_SIZE = 7;
	defparam lut_2409.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_2411 ({sk[856], i_9_, i_19_, n_n1118, n_n1048, x76x, x213x}, x1320x);
	defparam lut_2411.LUT_SIZE = 7;
	defparam lut_2411.mask = 128'h57ffffff57ffffff0000030300000357;

	lut_sub lut_2414 ({sk[857], i_13_, i_12_, x292x, x11x, x7416x, x7418x}, x7421x);
	defparam lut_2414.LUT_SIZE = 7;
	defparam lut_2414.mask = 128'h57ffffff57ffffff0537050505050505;

	lut_sub lut_2417 ({sk[858], i_11_, i_19_, x279x, x208x, x229x, x347x}, x752x);
	defparam lut_2417.LUT_SIZE = 7;
	defparam lut_2417.mask = 128'h57ffffff57ffffff0000000f111f111f;

	lut_sub lut_2421 ({sk[859], x11x, x213x, x7425x, x7426x, x7423x, x7424x}, x755x);
	defparam lut_2421.LUT_SIZE = 7;
	defparam lut_2421.mask = 128'h57ffffff57ffffff000055ff3f3f7fff;

	lut_sub lut_2426 ({sk[860], i_11_, i_19_, x279x, x208x, x229x, x347x}, x754x);
	defparam lut_2426.LUT_SIZE = 7;
	defparam lut_2426.mask = 128'h57ffffff57ffffff0000111f1111111f;

	lut_sub lut_2430 ({sk[861], x208x, x50x, x288x, x12x, x7427x, x7428x}, x1316x);
	defparam lut_2430.LUT_SIZE = 7;
	defparam lut_2430.mask = 128'h57ffffff57ffffff0000000500030007;

	lut_sub lut_2433 ({sk[862], i_28_, i_25_, i_34_, i_29_}, x7431x);
	defparam lut_2433.LUT_SIZE = 5;
	defparam lut_2433.mask = 32'h77772000;

	lut_sub lut_2435 ({sk[863], x11x, x213x, x7425x, x7426x, x7423x, x7424x}, x654x);
	defparam lut_2435.LUT_SIZE = 7;
	defparam lut_2435.mask = 128'h57ffffff57ffffff000055ff3f3f7fff;

	lut_sub lut_2440 ({sk[864], n_n1048, x208x, n_n1225, x50x, n_n1028, x371x}, x1308x);
	defparam lut_2440.LUT_SIZE = 7;
	defparam lut_2440.mask = 128'h57ffffff57ffffff0000001100050015;

	lut_sub lut_2443 ({sk[865], x208x, x50x, x12x, x7431x, x7427x, x7428x}, x1309x);
	defparam lut_2443.LUT_SIZE = 7;
	defparam lut_2443.mask = 128'h57ffffff57ffffff0000000500030007;

	lut_sub lut_2446 ({sk[866], i_13_, i_18_, i_19_, n_n1361, x229x, x476x}, x1311x);
	defparam lut_2446.LUT_SIZE = 7;
	defparam lut_2446.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_2448 ({sk[867], i_11_, i_19_, x279x, x208x, x229x, x347x}, x675x);
	defparam lut_2448.LUT_SIZE = 7;
	defparam lut_2448.mask = 128'h57ffffff57ffffff0000111f111f111f;

	lut_sub lut_2453 ({sk[868], i_19_, n_n1048, x208x, x50x, n_n1028, x7428x}, x674x);
	defparam lut_2453.LUT_SIZE = 7;
	defparam lut_2453.mask = 128'h57ffffff57ffffff0505050505370f3f;

	lut_sub lut_2457 ({sk[869], x208x, x50x, x12x, x78x, x7427x, x7428x}, x1305x);
	defparam lut_2457.LUT_SIZE = 7;
	defparam lut_2457.mask = 128'h57ffffff57ffffff0000000500030007;

	lut_sub lut_2460 ({sk[870], i_11_, i_19_, x279x, x208x, x229x, x347x}, x656x);
	defparam lut_2460.LUT_SIZE = 7;
	defparam lut_2460.mask = 128'h57ffffff57ffffff0000111f111f111f;

	lut_sub lut_2465 ({sk[871], i_9_, i_7_, i_6_, i_27_, i_26_, i_24_}, x7129x);
	defparam lut_2465.LUT_SIZE = 7;
	defparam lut_2465.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_2467 ({sk[872], i_20_, i_23_, i_17_, x10x, n_n460, x7129x}, x1562x);
	defparam lut_2467.LUT_SIZE = 7;
	defparam lut_2467.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2469 ({sk[873], i_20_, i_14_, i_17_, i_16_, x46x, x6876x}, x1563x);
	defparam lut_2469.LUT_SIZE = 7;
	defparam lut_2469.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_2471 ({sk[874], i_10_, i_14_, i_13_, i_16_}, x663x);
	defparam lut_2471.LUT_SIZE = 5;
	defparam lut_2471.mask = 32'h7777a020;

	lut_sub lut_2474 ({sk[875], i_9_, i_13_, i_11_, i_19_, x263x, x376x}, x1560x);
	defparam lut_2474.LUT_SIZE = 7;
	defparam lut_2474.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_2476 ({sk[876], i_8_, i_13_, i_18_, n_n1278, x263x, x404x}, x1561x);
	defparam lut_2476.LUT_SIZE = 7;
	defparam lut_2476.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2478 ({sk[877], i_35_, i_37_, n_n1274, x45x, x487x, x663x}, x1555x);
	defparam lut_2478.LUT_SIZE = 7;
	defparam lut_2478.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_2480 ({sk[878], i_20_, x54x, n_n245, n_n839, x303x, x44x}, x1558x);
	defparam lut_2480.LUT_SIZE = 7;
	defparam lut_2480.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_2482 ({sk[879], i_33_, x19x, x243x, x316x, x1555x, x1558x}, x7142x);
	defparam lut_2482.LUT_SIZE = 7;
	defparam lut_2482.mask = 128'h57ffffff57ffffff7777777f77777777;

	lut_sub lut_2486 ({sk[880], i_10_, i_5_, i_4_, i_0_, i_37_}, x7138x);
	defparam lut_2486.LUT_SIZE = 6;
	defparam lut_2486.mask = 64'h3f3fffff40000000;

	lut_sub lut_2488 ({sk[881], x317x, x1562x, x1563x, x1560x, x1561x, x7138x}, x7143x);
	defparam lut_2488.LUT_SIZE = 7;
	defparam lut_2488.mask = 128'h57ffffff57ffffff005555553f7f7f7f;

	lut_sub lut_2493 ({sk[882], i_20_, i_27_, i_28_, i_25_, i_33_, x47x}, x331x);
	defparam lut_2493.LUT_SIZE = 7;
	defparam lut_2493.mask = 128'h57ffffff57ffffff0000000001000000;

	lut_sub lut_2495 ({sk[883], i_30_, i_7_, i_8_, i_13_, x246x, x220x}, x1628x);
	defparam lut_2495.LUT_SIZE = 7;
	defparam lut_2495.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_2497 ({sk[884], i_34_, i_35_, i_37_, x76x, n_n1263, x80x}, x1629x);
	defparam lut_2497.LUT_SIZE = 7;
	defparam lut_2497.mask = 128'h57ffffff57ffffff0000000000010000;

	lut_sub lut_2499 ({sk[885], i_14_, i_37_, n_n1375, n_n1390, x11x, n_n1422}, x1630x);
	defparam lut_2499.LUT_SIZE = 7;
	defparam lut_2499.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_2501 ({sk[886], i_12_, x43x, x331x, x1628x, x1629x, x1630x}, x7062x);
	defparam lut_2501.LUT_SIZE = 7;
	defparam lut_2501.mask = 128'h57ffffff57ffffff7f7f7fff7f7f7f7f;

	lut_sub lut_2506 ({sk[887], i_20_, i_8_, n_n1404, n_n1431, x496x, x7068x}, x1624x);
	defparam lut_2506.LUT_SIZE = 7;
	defparam lut_2506.mask = 128'h57ffffff57ffffff0037000500000000;

	lut_sub lut_2509 ({sk[888], i_8_, n_n1274, n_n1431, x496x, x7066x, x7070x}, x7071x);
	defparam lut_2509.LUT_SIZE = 7;
	defparam lut_2509.mask = 128'h57ffffff57ffffff0505053700000033;

	lut_sub lut_2512 ({sk[889], i_0_, i_35_, i_37_, x1624x, x7071x}, x1619x);
	defparam lut_2512.LUT_SIZE = 6;
	defparam lut_2512.mask = 64'h3f3fffff07000000;

	lut_sub lut_2515 ({sk[890], i_12_, i_17_, i_37_, x10x, n_n1202, x445x}, x1618x);
	defparam lut_2515.LUT_SIZE = 7;
	defparam lut_2515.mask = 128'h57ffffff57ffffff0001000100010000;

	lut_sub lut_2518 ({sk[891], i_28_, i_23_, i_29_, x10x, x76x, x269x}, x1620x);
	defparam lut_2518.LUT_SIZE = 7;
	defparam lut_2518.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2520 ({sk[892], i_14_, i_32_, i_29_, n_n1390, x11x, x366x}, x1621x);
	defparam lut_2520.LUT_SIZE = 7;
	defparam lut_2520.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2522 ({sk[893], i_17_, x43x, x331x, x1618x, x1620x, x1621x}, x7077x);
	defparam lut_2522.LUT_SIZE = 7;
	defparam lut_2522.mask = 128'h57ffffff57ffffff7f7f7fff7f7f7f7f;

	lut_sub lut_2527 ({sk[894], i_13_, i_12_, i_17_, i_16_}, x29x);
	defparam lut_2527.LUT_SIZE = 5;
	defparam lut_2527.mask = 32'h7777a800;

	lut_sub lut_2530 ({sk[895], i_27_, i_26_, i_24_, i_35_, i_37_}, x269x);
	defparam lut_2530.LUT_SIZE = 6;
	defparam lut_2530.mask = 64'h3f3fffff40000000;

	lut_sub lut_2532 ({sk[896], i_27_, i_28_, i_26_, i_35_, i_37_}, x366x);
	defparam lut_2532.LUT_SIZE = 6;
	defparam lut_2532.mask = 64'h3f3fffff40000000;

	lut_sub lut_2534 ({sk[897], i_30_, i_27_, i_28_, i_23_, i_31_, i_29_}, x445x);
	defparam lut_2534.LUT_SIZE = 7;
	defparam lut_2534.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_2536 ({sk[898], i_0_, n_n1404, n_n620, x256x, x7057x, x770x}, x768x);
	defparam lut_2536.LUT_SIZE = 7;
	defparam lut_2536.mask = 128'h57ffffff57ffffff333f777f000f000f;

	lut_sub lut_2540 ({sk[899], x1608x, x1609x, x1610x, x1611x, x7089x}, x7093x);
	defparam lut_2540.LUT_SIZE = 6;
	defparam lut_2540.mask = 64'h3f3fffff7fffffff;

	lut_sub lut_2546 ({sk[900], i_27_, i_28_, i_23_, i_17_, i_16_, i_29_}, x220x);
	defparam lut_2546.LUT_SIZE = 7;
	defparam lut_2546.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_2548 ({sk[901], i_9_, i_7_, i_12_, i_31_, i_34_, i_35_}, x7988x);
	defparam lut_2548.LUT_SIZE = 7;
	defparam lut_2548.mask = 128'h57ffffff57ffffff0000040000000000;

	lut_sub lut_2550 ({sk[902], i_27_, i_28_, i_23_, i_34_, i_33_, i_35_}, x505x);
	defparam lut_2550.LUT_SIZE = 7;
	defparam lut_2550.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_2552 ({sk[903], i_14_, i_12_, i_17_, i_16_}, x668x);
	defparam lut_2552.LUT_SIZE = 5;
	defparam lut_2552.mask = 32'h7777a800;

	lut_sub lut_2555 ({sk[904], i_9_, i_2_}, x7900x);
	defparam lut_2555.LUT_SIZE = 3;
	defparam lut_2555.mask = 8'h34;

	lut_sub lut_2557 ({sk[905], i_10_, i_7_, i_11_, i_23_, i_24_, i_19_}, x393x);
	defparam lut_2557.LUT_SIZE = 7;
	defparam lut_2557.mask = 128'h57ffffff57ffffff0000000000008000;

	lut_sub lut_2559 ({sk[906], i_8_, i_18_, i_19_, x279x, x208x, x50x}, x1277x);
	defparam lut_2559.LUT_SIZE = 7;
	defparam lut_2559.mask = 128'h57ffffff57ffffff0003000700000005;

	lut_sub lut_2562 ({sk[907], i_11_, i_19_, x279x, x208x, x229x, x347x}, x671x);
	defparam lut_2562.LUT_SIZE = 7;
	defparam lut_2562.mask = 128'h57ffffff57ffffff0000111f111f111f;

	lut_sub lut_2567 ({sk[908], i_26_, i_24_, i_33_, i_35_, i_38_, x42x}, x7456x);
	defparam lut_2567.LUT_SIZE = 7;
	defparam lut_2567.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_2569 ({sk[909], i_24_, i_22_, x58x, n_n1438, n_n1197, x210x}, x1275x);
	defparam lut_2569.LUT_SIZE = 7;
	defparam lut_2569.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_2571 ({sk[910], i_11_, i_19_, x279x, x208x, x229x, x347x}, x676x);
	defparam lut_2571.LUT_SIZE = 7;
	defparam lut_2571.mask = 128'h57ffffff57ffffff0000111f111f111f;

	lut_sub lut_2576 ({sk[911], n_n1486, n_n1048, x76x, x213x, x7420x, x371x}, x1268x);
	defparam lut_2576.LUT_SIZE = 7;
	defparam lut_2576.mask = 128'h57ffffff57ffffff0000000001010155;

	lut_sub lut_2579 ({sk[912], i_28_, i_32_, i_29_, x11x, x7423x, x81x}, x1270x);
	defparam lut_2579.LUT_SIZE = 7;
	defparam lut_2579.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2581 ({sk[913], x11x, x71x, x12x, x7415x, x7416x, x7418x}, x1271x);
	defparam lut_2581.LUT_SIZE = 7;
	defparam lut_2581.mask = 128'h57ffffff57ffffff0000000300000057;

	lut_sub lut_2584 ({sk[914], i_8_, i_31_}, x284x);
	defparam lut_2584.LUT_SIZE = 3;
	defparam lut_2584.mask = 8'h38;

	lut_sub lut_2586 ({sk[915], i_10_, i_13_, i_12_, i_18_, i_19_}, x1261x);
	defparam lut_2586.LUT_SIZE = 6;
	defparam lut_2586.mask = 64'h3f3fffff00000100;

	lut_sub lut_2588 ({sk[916], i_3_, i_13_, i_12_, i_11_, i_18_, i_19_}, x766x);
	defparam lut_2588.LUT_SIZE = 7;
	defparam lut_2588.mask = 128'h57ffffff57ffffff005f000000030000;

	lut_sub lut_2592 ({sk[917], i_10_, n_n1361, x313x, x284x, x1261x, x766x}, x1256x);
	defparam lut_2592.LUT_SIZE = 7;
	defparam lut_2592.mask = 128'h57ffffff57ffffff0000000300000007;

	lut_sub lut_2595 ({sk[918], n_n1048, x76x, x213x, n_n1225, x7420x, x371x}, x1257x);
	defparam lut_2595.LUT_SIZE = 7;
	defparam lut_2595.mask = 128'h57ffffff57ffffff0001000100010505;

	lut_sub lut_2598 ({sk[919], i_24_, x42x, n_n1361, n_n1055, x208x, n_n1340}, x1259x);
	defparam lut_2598.LUT_SIZE = 7;
	defparam lut_2598.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_2600 ({sk[920], i_25_, i_26_, i_24_, i_32_, i_35_, i_38_}, x270x);
	defparam lut_2600.LUT_SIZE = 7;
	defparam lut_2600.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_2602 ({sk[921], x11x, x213x, x7425x, x7426x, x7423x, x7424x}, x677x);
	defparam lut_2602.LUT_SIZE = 7;
	defparam lut_2602.mask = 128'h57ffffff57ffffff000055ff3f3f7fff;

	lut_sub lut_2607 ({sk[922], i_10_, i_12_, n_n1345, x5x, x270x, x679x}, x1247x);
	defparam lut_2607.LUT_SIZE = 7;
	defparam lut_2607.mask = 128'h57ffffff57ffffff0000000000110013;

	lut_sub lut_2610 ({sk[923], i_24_, i_19_, n_n1361, n_n1048, x76x, x288x}, x1249x);
	defparam lut_2610.LUT_SIZE = 7;
	defparam lut_2610.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_2612 ({sk[924], i_27_, i_28_, i_24_, i_35_, i_37_}, x7101x);
	defparam lut_2612.LUT_SIZE = 6;
	defparam lut_2612.mask = 64'h3f3fffff40000000;

	lut_sub lut_2614 ({sk[925], i_34_, i_33_, i_29_, x7101x}, x482x);
	defparam lut_2614.LUT_SIZE = 5;
	defparam lut_2614.mask = 32'h77770040;

	lut_sub lut_2616 ({sk[926], i_32_, i_34_, i_33_, i_35_, i_37_}, x499x);
	defparam lut_2616.LUT_SIZE = 6;
	defparam lut_2616.mask = 64'h3f3fffff00400000;

	lut_sub lut_2618 ({sk[927], n_n1443, x211x, x496x, x7055x, x7056x, x683x}, x682x);
	defparam lut_2618.LUT_SIZE = 7;
	defparam lut_2618.mask = 128'h57ffffff57ffffff0000005503030357;

	lut_sub lut_2621 ({sk[928], i_8_, i_33_, i_35_, i_37_, x496x, x402x}, x1599x);
	defparam lut_2621.LUT_SIZE = 7;
	defparam lut_2621.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2623 ({sk[929], i_20_, i_33_, i_37_, x54x, n_n1429, x7056x}, x1601x);
	defparam lut_2623.LUT_SIZE = 7;
	defparam lut_2623.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_2625 ({sk[930], i_0_, i_33_, i_37_, x682x, x1599x, x1601x}, x1597x);
	defparam lut_2625.LUT_SIZE = 7;
	defparam lut_2625.mask = 128'h57ffffff57ffffff777f777700000000;

	lut_sub lut_2629 ({sk[931], i_13_, i_16_, n_n1375, x54x, x11x, x499x}, x1594x);
	defparam lut_2629.LUT_SIZE = 7;
	defparam lut_2629.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_2631 ({sk[932], i_28_, i_32_, i_29_, x51x, x260x, x269x}, x1595x);
	defparam lut_2631.LUT_SIZE = 7;
	defparam lut_2631.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2633 ({sk[933], i_17_, i_35_, i_37_, x10x, x50x, x67x}, x1596x);
	defparam lut_2633.LUT_SIZE = 7;
	defparam lut_2633.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_2635 ({sk[934], i_34_, i_33_, i_29_, n_n1314, x76x, x7101x}, x1598x);
	defparam lut_2635.LUT_SIZE = 7;
	defparam lut_2635.mask = 128'h57ffffff57ffffff0000000001000000;

	lut_sub lut_2637 ({sk[935], x1594x, x1595x, x1596x, x1598x}, x7104x);
	defparam lut_2637.LUT_SIZE = 5;
	defparam lut_2637.mask = 32'h77777fff;

	lut_sub lut_2642 ({sk[936], i_5_, i_4_, i_11_, i_2_, i_19_}, x7146x);
	defparam lut_2642.LUT_SIZE = 6;
	defparam lut_2642.mask = 64'h3f3fffff80000000;

	lut_sub lut_2644 ({sk[937], i_9_, i_3_, i_4_, i_2_, i_18_}, x7149x);
	defparam lut_2644.LUT_SIZE = 6;
	defparam lut_2644.mask = 64'h3f3fffff00800000;

	lut_sub lut_2646 ({sk[938], i_9_, i_10_, i_13_, n_n1397, x376x, x220x}, x1551x);
	defparam lut_2646.LUT_SIZE = 7;
	defparam lut_2646.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2648 ({sk[939], n_n1274, x259x, x45x, x44x, x6899x, x7153x}, x686x);
	defparam lut_2648.LUT_SIZE = 7;
	defparam lut_2648.mask = 128'h57ffffff57ffffff01010101010101ff;

	lut_sub lut_2651 ({sk[940], n_n1278, n_n301, n_n152, x1551x, x87x, x686x}, x685x);
	defparam lut_2651.LUT_SIZE = 7;
	defparam lut_2651.mask = 128'h57ffffff57ffffff0f0f3f3f0f5f3f7f;

	lut_sub lut_2655 ({sk[941], x499x, x7145x, x7146x, x7148x, x7149x, x7150x}, x1546x);
	defparam lut_2655.LUT_SIZE = 7;
	defparam lut_2655.mask = 128'h57ffffff57ffffff0000000001010155;

	lut_sub lut_2658 ({sk[942], i_20_, x54x, n_n853, n_n245, x303x, x44x}, x1547x);
	defparam lut_2658.LUT_SIZE = 7;
	defparam lut_2658.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_2660 ({sk[943], x41x, x498x, x482x, x326x, x1546x, x1547x}, x7157x);
	defparam lut_2660.LUT_SIZE = 7;
	defparam lut_2660.mask = 128'h57ffffff57ffffff777777ff777f77ff;

	lut_sub lut_2665 ({sk[944], i_27_, i_23_, i_24_, i_17_}, x7997x);
	defparam lut_2665.LUT_SIZE = 5;
	defparam lut_2665.mask = 32'h77778000;

	lut_sub lut_2667 ({sk[945], i_9_, i_7_, i_14_, i_28_, i_31_, i_34_}, x7998x);
	defparam lut_2667.LUT_SIZE = 7;
	defparam lut_2667.mask = 128'h57ffffff57ffffff0000100000000000;

	lut_sub lut_2669 ({sk[946], i_27_, i_14_, i_28_, i_13_, i_12_, i_24_}, x8000x);
	defparam lut_2669.LUT_SIZE = 7;
	defparam lut_2669.mask = 128'h57ffffff57ffffff0000800000000000;

	lut_sub lut_2671 ({sk[947], i_14_, i_12_, i_17_, i_16_}, x687x);
	defparam lut_2671.LUT_SIZE = 5;
	defparam lut_2671.mask = 32'h7777a800;

	lut_sub lut_2674 ({sk[948], i_27_, i_28_, i_26_, i_32_, i_31_, i_29_}, x7913x);
	defparam lut_2674.LUT_SIZE = 7;
	defparam lut_2674.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_2676 ({sk[949], i_27_, i_28_, i_32_, i_31_, i_34_, i_29_}, x7914x);
	defparam lut_2676.LUT_SIZE = 7;
	defparam lut_2676.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_2678 ({sk[950], i_9_, i_12_}, x68x);
	defparam lut_2678.LUT_SIZE = 3;
	defparam lut_2678.mask = 8'h31;

	lut_sub lut_2680 ({sk[951], i_28_, i_25_, i_26_, i_33_, i_29_}, x691x);
	defparam lut_2680.LUT_SIZE = 6;
	defparam lut_2680.mask = 64'h3f3fffffa0800000;

	lut_sub lut_2683 ({sk[952], i_24_, i_38_, x42x, x321x, n_n1340, x476x}, x1225x);
	defparam lut_2683.LUT_SIZE = 7;
	defparam lut_2683.mask = 128'h57ffffff57ffffff0000050700000505;

	lut_sub lut_2686 ({sk[953], i_12_, i_24_, i_38_, n_n1307, n_n1303, x288x}, x1226x);
	defparam lut_2686.LUT_SIZE = 7;
	defparam lut_2686.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_2688 ({sk[954], i_9_, i_12_, i_24_, i_38_, x77x, x78x}, x1227x);
	defparam lut_2688.LUT_SIZE = 7;
	defparam lut_2688.mask = 128'h57ffffff57ffffff0000000000000100;

	lut_sub lut_2690 ({sk[955], i_33_, x42x, n_n1397, n_n1387, x318x, x7499x}, x7501x);
	defparam lut_2690.LUT_SIZE = 7;
	defparam lut_2690.mask = 128'h57ffffff57ffffff0000000000000357;

	lut_sub lut_2693 ({sk[956], i_38_, n_n1454, x49x, n_n1288, x7492x, x691x}, x7502x);
	defparam lut_2693.LUT_SIZE = 7;
	defparam lut_2693.mask = 128'h57ffffff57ffffff001100110011001f;

	lut_sub lut_2696 ({sk[957], x1225x, x1226x, x1227x, x7501x, x7502x}, n_n1882);
	defparam lut_2696.LUT_SIZE = 6;
	defparam lut_2696.mask = 64'h3f3fffff7fffffff;

	lut_sub lut_2702 ({sk[958], i_32_, i_31_, i_34_, i_37_}, x7108x);
	defparam lut_2702.LUT_SIZE = 5;
	defparam lut_2702.mask = 32'h77770100;

	lut_sub lut_2704 ({sk[959], i_30_, i_27_, i_28_, i_23_, i_24_, i_29_}, x7109x);
	defparam lut_2704.LUT_SIZE = 7;
	defparam lut_2704.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_2706 ({sk[960], i_14_, i_12_, i_17_, i_16_}, x694x);
	defparam lut_2706.LUT_SIZE = 5;
	defparam lut_2706.mask = 32'h7777a800;

	lut_sub lut_2709 ({sk[961], i_20_, i_7_, i_13_, i_12_, i_17_, i_16_}, x693x);
	defparam lut_2709.LUT_SIZE = 7;
	defparam lut_2709.mask = 128'h57ffffff57ffffff000000000000a800;

	lut_sub lut_2712 ({sk[962], x57x, x8x, x316x, x324x, x7108x, x7109x}, x7111x);
	defparam lut_2712.LUT_SIZE = 7;
	defparam lut_2712.mask = 128'h57ffffff57ffffff00001111000f111f;

	lut_sub lut_2715 ({sk[963], i_5_, i_4_, i_0_, i_32_}, x7161x);
	defparam lut_2715.LUT_SIZE = 5;
	defparam lut_2715.mask = 32'h77778000;

	lut_sub lut_2717 ({sk[964], i_20_, i_7_, i_6_, i_12_, x46x, x7161x}, x358x);
	defparam lut_2717.LUT_SIZE = 7;
	defparam lut_2717.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_2719 ({sk[965], i_13_, i_12_, i_16_, i_33_, i_37_}, x470x);
	defparam lut_2719.LUT_SIZE = 6;
	defparam lut_2719.mask = 64'h3f3fffff40000000;

	lut_sub lut_2721 ({sk[966], i_8_, i_6_, i_13_, i_12_, i_16_}, x7158x);
	defparam lut_2721.LUT_SIZE = 6;
	defparam lut_2721.mask = 64'h3f3fffff80000000;

	lut_sub lut_2723 ({sk[967], i_6_, i_13_, i_12_, i_16_}, x7159x);
	defparam lut_2723.LUT_SIZE = 5;
	defparam lut_2723.mask = 32'h77778000;

	lut_sub lut_2725 ({sk[968], i_20_, x46x, n_n460, x6886x, x7158x, x7159x}, x696x);
	defparam lut_2725.LUT_SIZE = 7;
	defparam lut_2725.mask = 128'h57ffffff57ffffff0005333700050005;

	lut_sub lut_2728 ({sk[969], n_n1443, n_n301, x48x, x41x, x207x, x221x}, x698x);
	defparam lut_2728.LUT_SIZE = 7;
	defparam lut_2728.mask = 128'h57ffffff57ffffff0000000f1111111f;

	lut_sub lut_2731 ({sk[970], i_17_, n_n793, x43x, n_n1397, n_n1305, x49x}, x1540x);
	defparam lut_2731.LUT_SIZE = 7;
	defparam lut_2731.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_2733 ({sk[971], i_17_, n_n1375, x54x, n_n301, n_n1340, x14x}, x1541x);
	defparam lut_2733.LUT_SIZE = 7;
	defparam lut_2733.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_2735 ({sk[972], i_28_, i_33_, i_29_, x49x, x259x, x318x}, x1542x);
	defparam lut_2735.LUT_SIZE = 7;
	defparam lut_2735.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2737 ({sk[973], i_37_, n_n1437, x698x, x1540x, x1541x, x1542x}, x1536x);
	defparam lut_2737.LUT_SIZE = 7;
	defparam lut_2737.mask = 128'h57ffffff57ffffff000000007f7f7fff;

	lut_sub lut_2742 ({sk[974], i_20_, x59x, x43x, n_n1306, x46x, x7161x}, x1535x);
	defparam lut_2742.LUT_SIZE = 7;
	defparam lut_2742.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_2744 ({sk[975], n_n504, n_n245, x508x, x470x, x696x, x1535x}, x7172x);
	defparam lut_2744.LUT_SIZE = 7;
	defparam lut_2744.mask = 128'h57ffffff57ffffff555f555f555f777f;

	lut_sub lut_2748 ({sk[976], i_30_, i_28_, i_32_, i_31_, i_36_, i_35_}, x8011x);
	defparam lut_2748.LUT_SIZE = 7;
	defparam lut_2748.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_2750 ({sk[977], i_2_, i_17_, i_21_, i_16_}, x8008x);
	defparam lut_2750.LUT_SIZE = 5;
	defparam lut_2750.mask = 32'h77778000;

	lut_sub lut_2752 ({sk[978], i_28_, i_24_, i_34_, i_38_, n_n1305, x14x}, x286x);
	defparam lut_2752.LUT_SIZE = 7;
	defparam lut_2752.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_2754 ({sk[979], i_24_, i_34_, i_38_, x49x, x223x, n_n1202}, x700x);
	defparam lut_2754.LUT_SIZE = 7;
	defparam lut_2754.mask = 128'h57ffffff57ffffff0005003700050005;

	lut_sub lut_2757 ({sk[980], i_9_, i_13_, i_24_, n_n1307, n_n1303, x7520x}, x1208x);
	defparam lut_2757.LUT_SIZE = 7;
	defparam lut_2757.mask = 128'h57ffffff57ffffff0000010000000000;

	lut_sub lut_2759 ({sk[981], i_28_, i_26_, i_24_, i_22_, x51x, n_n1149}, x1209x);
	defparam lut_2759.LUT_SIZE = 7;
	defparam lut_2759.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_2761 ({sk[982], i_28_, i_1_, i_31_, x292x, n_n1118, x389x}, x1210x);
	defparam lut_2761.LUT_SIZE = 7;
	defparam lut_2761.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2763 ({sk[983], i_38_, x49x, n_n1288, x14x, x7516x, x7519x}, x7525x);
	defparam lut_2763.LUT_SIZE = 7;
	defparam lut_2763.mask = 128'h57ffffff57ffffff0003000300035557;

	lut_sub lut_2766 ({sk[984], i_13_, x286x, x1208x, x1209x, x1210x, x7525x}, x7529x);
	defparam lut_2766.LUT_SIZE = 7;
	defparam lut_2766.mask = 128'h57ffffff57ffffff7fff7fff7fffffff;

	lut_sub lut_2772 ({sk[985], i_30_, i_32_, i_31_}, x7006x);
	defparam lut_2772.LUT_SIZE = 4;
	defparam lut_2772.mask = 16'h5540;

	lut_sub lut_2774 ({sk[986], i_30_, i_28_, i_32_, i_31_, i_34_, i_29_}, x398x);
	defparam lut_2774.LUT_SIZE = 7;
	defparam lut_2774.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_2776 ({sk[987], i_23_, i_24_, i_32_, i_31_, i_34_}, x6983x);
	defparam lut_2776.LUT_SIZE = 6;
	defparam lut_2776.mask = 64'h3f3fffff40000000;

	lut_sub lut_2778 ({sk[988], i_9_, i_14_, i_13_, n_n1322, x80x, x376x}, x1532x);
	defparam lut_2778.LUT_SIZE = 7;
	defparam lut_2778.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_2780 ({sk[989], i_17_, x43x, n_n1307, n_n853, n_n1458, x67x}, x1526x);
	defparam lut_2780.LUT_SIZE = 7;
	defparam lut_2780.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_2782 ({sk[990], i_9_, i_10_, i_14_, n_n1322, x80x, x376x}, x1531x);
	defparam lut_2782.LUT_SIZE = 7;
	defparam lut_2782.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2784 ({sk[991], i_10_, i_13_, i_32_, x10x, x14x, x48x}, x7181x);
	defparam lut_2784.LUT_SIZE = 7;
	defparam lut_2784.mask = 128'h57ffffff57ffffff0100010000000100;

	lut_sub lut_2787 ({sk[992], i_34_, i_37_, x1532x, x1531x, x7181x}, x1525x);
	defparam lut_2787.LUT_SIZE = 6;
	defparam lut_2787.mask = 64'h3f3fffff0000007f;

	lut_sub lut_2791 ({sk[993], n_n1408, x49x, x258x, x7175x, x7173x, x7174x}, x1522x);
	defparam lut_2791.LUT_SIZE = 7;
	defparam lut_2791.mask = 128'h57ffffff57ffffff0000000500000307;

	lut_sub lut_2794 ({sk[994], i_10_, i_29_, x43x, n_n504, x74x, x41x}, x1523x);
	defparam lut_2794.LUT_SIZE = 7;
	defparam lut_2794.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_2796 ({sk[995], i_37_, n_n1404, x508x, x1526x, x1522x, x1523x}, x7184x);
	defparam lut_2796.LUT_SIZE = 7;
	defparam lut_2796.mask = 128'h57ffffff57ffffff777777777f7f7fff;

	lut_sub lut_2801 ({sk[996], i_17_, x10x, n_n1307, n_n853, n_n839, x221x}, x1518x);
	defparam lut_2801.LUT_SIZE = 7;
	defparam lut_2801.mask = 128'h57ffffff57ffffff0000001500000000;

	lut_sub lut_2804 ({sk[997], i_10_, i_14_, i_13_, i_16_, x48x, x41x}, x7191x);
	defparam lut_2804.LUT_SIZE = 7;
	defparam lut_2804.mask = 128'h57ffffff57ffffff1010000000100000;

	lut_sub lut_2807 ({sk[998], i_8_, i_6_, i_14_, i_12_, i_16_}, x7185x);
	defparam lut_2807.LUT_SIZE = 6;
	defparam lut_2807.mask = 64'h3f3fffff80000000;

	lut_sub lut_2809 ({sk[999], i_6_, i_14_, i_12_, i_16_}, x7186x);
	defparam lut_2809.LUT_SIZE = 5;
	defparam lut_2809.mask = 32'h77778000;

	lut_sub lut_2811 ({sk[1000], i_20_, x46x, n_n460, x6886x, x7185x, x7186x}, x707x);
	defparam lut_2811.LUT_SIZE = 7;
	defparam lut_2811.mask = 128'h57ffffff57ffffff0005333700050005;

	lut_sub lut_2814 ({sk[1001], i_35_, i_37_, x10x, n_n245, x358x, x707x}, x7192x);
	defparam lut_2814.LUT_SIZE = 7;
	defparam lut_2814.mask = 128'h57ffffff57ffffff0000053700000033;

	lut_sub lut_2817 ({sk[1002], n_n1443, x49x, x48x, x259x, x221x, x7188x}, x1510x);
	defparam lut_2817.LUT_SIZE = 7;
	defparam lut_2817.mask = 128'h57ffffff57ffffff0000000500001115;

	lut_sub lut_2820 ({sk[1003], i_34_, i_35_, i_37_, x1518x, x7191x, x1510x}, x7193x);
	defparam lut_2820.LUT_SIZE = 7;
	defparam lut_2820.mask = 128'h57ffffff57ffffff55555555557f5555;

	lut_sub lut_2824 ({sk[1004], i_10_, i_7_, i_3_, i_23_, i_18_, i_24_}, x382x);
	defparam lut_2824.LUT_SIZE = 7;
	defparam lut_2824.mask = 128'h57ffffff57ffffff0000000000000080;

	lut_sub lut_2826 ({sk[1005], i_28_, i_25_, i_26_, i_24_, i_38_, i_29_}, x456x);
	defparam lut_2826.LUT_SIZE = 7;
	defparam lut_2826.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_2828 ({sk[1006], i_9_, i_3_, i_13_, i_11_, i_22_}, x1378x);
	defparam lut_2828.LUT_SIZE = 6;
	defparam lut_2828.mask = 64'h3f3fffff00002000;

	lut_sub lut_2830 ({sk[1007], i_7_, i_14_, i_13_, i_12_}, x717x);
	defparam lut_2830.LUT_SIZE = 5;
	defparam lut_2830.mask = 32'h777700a8;

	lut_sub lut_2833 ({sk[1008], i_9_, i_6_, i_23_, i_24_}, x7145x);
	defparam lut_2833.LUT_SIZE = 5;
	defparam lut_2833.mask = 32'h77778000;

	lut_sub lut_2835 ({sk[1009], i_5_, i_6_, i_23_, i_24_}, x7148x);
	defparam lut_2835.LUT_SIZE = 5;
	defparam lut_2835.mask = 32'h77778000;

	lut_sub lut_2837 ({sk[1010], n_n1408, n_n1422, x7145x, x7146x, x7148x, x7149x}, x1502x);
	defparam lut_2837.LUT_SIZE = 7;
	defparam lut_2837.mask = 128'h57ffffff57ffffff000000000000111f;

	lut_sub lut_2840 ({sk[1011], i_9_, i_14_, i_13_, n_n1397, n_n1322, x376x}, x1503x);
	defparam lut_2840.LUT_SIZE = 7;
	defparam lut_2840.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_2842 ({sk[1012], i_8_, i_14_, i_16_, n_n1274, x45x, x7202x}, x1504x);
	defparam lut_2842.LUT_SIZE = 7;
	defparam lut_2842.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2844 ({sk[1013], i_9_, i_10_, i_14_, n_n1397, x376x, x220x}, x1505x);
	defparam lut_2844.LUT_SIZE = 7;
	defparam lut_2844.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2846 ({sk[1014], i_13_, i_37_, x10x, x87x, x1504x, x1505x}, x1501x);
	defparam lut_2846.LUT_SIZE = 7;
	defparam lut_2846.mask = 128'h57ffffff57ffffff000077770000777f;

	lut_sub lut_2850 ({sk[1015], i_37_, x10x, n_n1278, x404x, n_n179, x256x}, x1498x);
	defparam lut_2850.LUT_SIZE = 7;
	defparam lut_2850.mask = 128'h57ffffff57ffffff0000000000000001;

	lut_sub lut_2852 ({sk[1016], x80x, x404x, x41x, x7196x, x7197x, x7198x}, x1499x);
	defparam lut_2852.LUT_SIZE = 7;
	defparam lut_2852.mask = 128'h57ffffff57ffffff0000000000110515;

	lut_sub lut_2855 ({sk[1017], i_37_, n_n1375, x1502x, x1503x, x1498x, x1499x}, x7207x);
	defparam lut_2855.LUT_SIZE = 7;
	defparam lut_2855.mask = 128'h57ffffff57ffffff7777777777777fff;

	lut_sub lut_2860 ({sk[1018], i_5_, i_6_, i_4_, i_1_, i_0_}, x7213x);
	defparam lut_2860.LUT_SIZE = 6;
	defparam lut_2860.mask = 64'h3f3fffff80000000;

	lut_sub lut_2862 ({sk[1019], i_7_, i_5_, i_6_, i_32_, i_37_}, x1496x);
	defparam lut_2862.LUT_SIZE = 6;
	defparam lut_2862.mask = 64'h3f3fffff40000000;

	lut_sub lut_2864 ({sk[1020], i_8_, i_5_, i_6_, i_35_, i_37_}, x1497x);
	defparam lut_2864.LUT_SIZE = 6;
	defparam lut_2864.mask = 64'h3f3fffff40000000;

	lut_sub lut_2866 ({sk[1021], i_20_, x54x, n_n152, x44x, x1496x, x1497x}, x1494x);
	defparam lut_2866.LUT_SIZE = 7;
	defparam lut_2866.mask = 128'h57ffffff57ffffff0000000700000000;

	lut_sub lut_2869 ({sk[1022], x243x, x366x, x7145x, x7146x, x7148x, x7149x}, x1495x);
	defparam lut_2869.LUT_SIZE = 7;
	defparam lut_2869.mask = 128'h57ffffff57ffffff000000000000111f;

	lut_sub lut_2872 ({sk[1023], i_9_, i_10_, i_13_, x376x, x7208x, x7209x}, x1489x);
	defparam lut_2872.LUT_SIZE = 7;
	defparam lut_2872.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2874 ({sk[1024], i_10_, i_14_, i_16_, i_37_, x87x, x1489x}, x7221x);
	defparam lut_2874.LUT_SIZE = 7;
	defparam lut_2874.mask = 128'h57ffffff57ffffff5755555555555555;

	lut_sub lut_2877 ({sk[1025], x404x, x41x, x269x, x7196x, x7197x, x7211x}, x1490x);
	defparam lut_2877.LUT_SIZE = 7;
	defparam lut_2877.mask = 128'h57ffffff57ffffff0000001100050015;

	lut_sub lut_2880 ({sk[1026], i_20_, i_17_, i_16_, x46x, x7213x, x7215x}, x1491x);
	defparam lut_2880.LUT_SIZE = 7;
	defparam lut_2880.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2882 ({sk[1027], i_17_, x10x, x1494x, x1495x, x1490x, x1491x}, x7222x);
	defparam lut_2882.LUT_SIZE = 7;
	defparam lut_2882.mask = 128'h57ffffff57ffffff77777fff77777777;

	lut_sub lut_2887 ({sk[1028], n_n787, n_n1118, n_n180, n_n179, x41x, x326x}, x722x);
	defparam lut_2887.LUT_SIZE = 7;
	defparam lut_2887.mask = 128'h57ffffff57ffffff111111111111111f;

	lut_sub lut_2890 ({sk[1029], i_14_, i_37_, x31x, x273x, x722x, x7229x}, x7233x);
	defparam lut_2890.LUT_SIZE = 7;
	defparam lut_2890.mask = 128'h57ffffff57ffffff1111111f11111111;

	lut_sub lut_2893 ({sk[1030], x351x, x256x, x1481x, x1482x, x1483x}, x7234x);
	defparam lut_2893.LUT_SIZE = 6;
	defparam lut_2893.mask = 64'h3f3fffff7f7f7fff;

	lut_sub lut_2898 ({sk[1031], i_3_, i_18_}, x8021x);
	defparam lut_2898.LUT_SIZE = 3;
	defparam lut_2898.mask = 8'h32;

	lut_sub lut_2900 ({sk[1032], i_9_, i_8_, i_3_, i_13_, i_11_, i_2_}, x1385x);
	defparam lut_2900.LUT_SIZE = 7;
	defparam lut_2900.mask = 128'h57ffffff57ffffff0000000020000000;

	lut_sub lut_2902 ({sk[1033], i_9_, i_8_, i_13_, i_2_, i_18_, i_19_}, x1387x);
	defparam lut_2902.LUT_SIZE = 7;
	defparam lut_2902.mask = 128'h57ffffff57ffffff0000000010000000;

	lut_sub lut_2904 ({sk[1034], i_7_, i_14_, i_12_, i_17_, i_16_}, x94x);
	defparam lut_2904.LUT_SIZE = 6;
	defparam lut_2904.mask = 64'h3f3fffff0000a800;

	lut_sub lut_2907 ({sk[1035], i_20_, x59x, x54x, x67x, x7006x, x485x}, x728x);
	defparam lut_2907.LUT_SIZE = 7;
	defparam lut_2907.mask = 128'h57ffffff57ffffff0000030300550357;

	lut_sub lut_2910 ({sk[1036], i_14_, i_12_, i_17_, i_16_}, x727x);
	defparam lut_2910.LUT_SIZE = 5;
	defparam lut_2910.mask = 32'h7777a800;

	lut_sub lut_2913 ({sk[1037], i_8_, n_n1375, x43x, x48x, x348x, x7114x}, x1578x);
	defparam lut_2913.LUT_SIZE = 7;
	defparam lut_2913.mask = 128'h57ffffff57ffffff0005111500001111;

	lut_sub lut_2916 ({sk[1038], i_20_, i_12_, i_23_, i_24_, x43x, x485x}, x1582x);
	defparam lut_2916.LUT_SIZE = 7;
	defparam lut_2916.mask = 128'h57ffffff57ffffff0000000010000000;

	lut_sub lut_2918 ({sk[1039], i_20_, i_25_, x275x, x505x, x94x, x727x}, x7116x);
	defparam lut_2918.LUT_SIZE = 7;
	defparam lut_2918.mask = 128'h57ffffff57ffffff0000000000330537;

	lut_sub lut_2921 ({sk[1040], i_17_, x43x, x728x, x1578x, x1582x, x7116x}, n_n1713);
	defparam lut_2921.LUT_SIZE = 7;
	defparam lut_2921.mask = 128'h57ffffff57ffffff7f7f7fff7f7f7f7f;

	lut_sub lut_2926 ({sk[1041], i_14_, i_13_, i_12_, i_16_}, x8042x);
	defparam lut_2926.LUT_SIZE = 5;
	defparam lut_2926.mask = 32'h77770080;

	lut_sub lut_2928 ({sk[1042], i_16_, i_31_, i_34_, i_35_}, x8043x);
	defparam lut_2928.LUT_SIZE = 5;
	defparam lut_2928.mask = 32'h77770400;

	lut_sub lut_2930 ({sk[1043], i_9_, i_7_, i_27_, i_14_, i_28_, i_23_}, x8044x);
	defparam lut_2930.LUT_SIZE = 7;
	defparam lut_2930.mask = 128'h57ffffff57ffffff0000800000000000;

	lut_sub lut_2932 ({sk[1044], i_17_, n_n1387, x505x, x8042x, x8043x, x8044x}, x730x);
	defparam lut_2932.LUT_SIZE = 7;
	defparam lut_2932.mask = 128'h57ffffff57ffffff111f11ff000f000f;

	lut_sub lut_2936 ({sk[1045], i_30_, i_14_, i_28_, i_13_, i_22_, i_32_}, x1028x);
	defparam lut_2936.LUT_SIZE = 7;
	defparam lut_2936.mask = 128'h57ffffff57ffffff0000010000000300;

	lut_sub lut_2939 ({sk[1046], i_25_, i_34_, i_33_, i_35_, i_38_}, x733x);
	defparam lut_2939.LUT_SIZE = 6;
	defparam lut_2939.mask = 64'h3f3fffff11001000;

	lut_sub lut_2942 ({sk[1047], i_7_, i_8_, i_31_, n_n1489, x238x, x733x}, x7688x);
	defparam lut_2942.LUT_SIZE = 7;
	defparam lut_2942.mask = 128'h57ffffff57ffffff0705000003000000;

	lut_sub lut_2945 ({sk[1048], i_28_, i_32_, i_31_, i_34_, i_33_, i_29_}, x7546x);
	defparam lut_2945.LUT_SIZE = 7;
	defparam lut_2945.mask = 128'h57ffffff57ffffff0800000000000000;

	lut_sub lut_2947 ({sk[1049], i_9_, i_8_, i_13_, i_18_, i_19_}, x1196x);
	defparam lut_2947.LUT_SIZE = 6;
	defparam lut_2947.mask = 64'h3f3fffff00001000;

	lut_sub lut_2949 ({sk[1050], i_13_, i_26_, x42x, x1196x, x737x, x7542x}, x1190x);
	defparam lut_2949.LUT_SIZE = 7;
	defparam lut_2949.mask = 128'h57ffffff57ffffff0015000000050000;

	lut_sub lut_2952 ({sk[1051], i_9_, i_13_, i_24_, i_29_, x376x, x311x}, x1191x);
	defparam lut_2952.LUT_SIZE = 7;
	defparam lut_2952.mask = 128'h57ffffff57ffffff0000100000000000;

	lut_sub lut_2954 ({sk[1052], i_28_, i_31_, i_33_, n_n1361, x76x, n_n1523}, x1194x);
	defparam lut_2954.LUT_SIZE = 7;
	defparam lut_2954.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2956 ({sk[1053], x11x, x51x, x61x, x12x, n_n1149, x7546x}, x7548x);
	defparam lut_2956.LUT_SIZE = 7;
	defparam lut_2956.mask = 128'h57ffffff57ffffff0000050500330537;

	lut_sub lut_2959 ({sk[1054], x50x, x66x, x1190x, x1191x, x1194x, x7548x}, n_n1875);
	defparam lut_2959.LUT_SIZE = 7;
	defparam lut_2959.mask = 128'h57ffffff57ffffff7fff7fff7fffffff;

	lut_sub lut_2965 ({sk[1055], i_30_, i_13_, i_29_, x454x, x375x, x17x}, x1202x);
	defparam lut_2965.LUT_SIZE = 7;
	defparam lut_2965.mask = 128'h57ffffff57ffffff1300030000000000;

	lut_sub lut_2968 ({sk[1056], i_9_, i_10_, i_24_, n_n1307, n_n1303, x7535x}, x1203x);
	defparam lut_2968.LUT_SIZE = 7;
	defparam lut_2968.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2970 ({sk[1057], i_31_, i_35_, i_38_, x76x, x257x}, x1204x);
	defparam lut_2970.LUT_SIZE = 6;
	defparam lut_2970.mask = 64'h3f3fffff01000000;

	lut_sub lut_2972 ({sk[1058], x49x, x50x, n_n1059, x315x, x7530x, x7532x}, x7537x);
	defparam lut_2972.LUT_SIZE = 7;
	defparam lut_2972.mask = 128'h57ffffff57ffffff0000030300550357;

	lut_sub lut_2975 ({sk[1059], i_10_, x286x, x1202x, x1203x, x1204x, x7537x}, n_n1873);
	defparam lut_2975.LUT_SIZE = 7;
	defparam lut_2975.mask = 128'h57ffffff57ffffff7fffffff7fff7fff;

	lut_sub lut_2981 ({sk[1060], i_28_, i_25_, i_24_, i_31_, n_n805, x76x}, x1188x);
	defparam lut_2981.LUT_SIZE = 7;
	defparam lut_2981.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_2983 ({sk[1061], i_9_, i_10_, i_24_, n_n1307, n_n1303, x311x}, x1189x);
	defparam lut_2983.LUT_SIZE = 7;
	defparam lut_2983.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_2985 ({sk[1062], i_26_, i_24_, i_38_, n_n1489, n_n1458, x744x}, x1182x);
	defparam lut_2985.LUT_SIZE = 7;
	defparam lut_2985.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_2987 ({sk[1063], i_12_, i_32_, x42x, x321x, x376x, n_n1059}, x1183x);
	defparam lut_2987.LUT_SIZE = 7;
	defparam lut_2987.mask = 128'h57ffffff57ffffff0015001100050000;

	lut_sub lut_2990 ({sk[1064], i_13_, i_24_, i_32_, i_38_, x14x, x71x}, x1185x);
	defparam lut_2990.LUT_SIZE = 7;
	defparam lut_2990.mask = 128'h57ffffff57ffffff0000000001000000;

	lut_sub lut_2992 ({sk[1065], i_29_, x1188x, x1189x, x1182x, x1183x, x1185x}, n_n1876);
	defparam lut_2992.LUT_SIZE = 7;
	defparam lut_2992.mask = 128'h57ffffff57ffffff7fffffff7f7f7f7f;

	lut_sub lut_2998 ({sk[1066], i_10_, i_24_, i_32_, i_38_, x14x, x71x}, x1154x);
	defparam lut_2998.LUT_SIZE = 7;
	defparam lut_2998.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_3000 ({sk[1067], i_31_, i_35_, i_38_, n_n1454, x42x, x50x}, x1155x);
	defparam lut_3000.LUT_SIZE = 7;
	defparam lut_3000.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_3002 ({sk[1068], i_9_, i_10_, i_13_, i_24_, x376x, x380x}, x1156x);
	defparam lut_3002.LUT_SIZE = 7;
	defparam lut_3002.mask = 128'h57ffffff57ffffff1010001000000000;

	lut_sub lut_3005 ({sk[1069], i_31_, x42x, x11x, n_n1340, x12x, x7564x}, x1157x);
	defparam lut_3005.LUT_SIZE = 7;
	defparam lut_3005.mask = 128'h57ffffff57ffffff0011001300110011;

	lut_sub lut_3008 ({sk[1070], i_24_, i_31_, i_33_, x42x, n_n805, x76x}, x1158x);
	defparam lut_3008.LUT_SIZE = 7;
	defparam lut_3008.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_3010 ({sk[1071], n_n1288, x14x, x12x, x78x, x7583x, x7584x}, x7587x);
	defparam lut_3010.LUT_SIZE = 7;
	defparam lut_3010.mask = 128'h57ffffff57ffffff0003000300035557;

	lut_sub lut_3013 ({sk[1072], x1154x, x1155x, x1156x, x1157x, x1158x, x7587x}, n_n1877);
	defparam lut_3013.LUT_SIZE = 7;
	defparam lut_3013.mask = 128'h57ffffff57ffffff7fffffffffffffff;

	lut_sub lut_3020 ({sk[1073], i_20_, i_24_, i_21_, i_22_, i_34_}, x1078x);
	defparam lut_3020.LUT_SIZE = 6;
	defparam lut_3020.mask = 64'h3f3fffff04004400;

	lut_sub lut_3023 ({sk[1074], i_27_, i_26_, i_23_, i_24_, i_16_, i_22_}, x1079x);
	defparam lut_3023.LUT_SIZE = 7;
	defparam lut_3023.mask = 128'h57ffffff57ffffff20a00000a0a00000;

	lut_sub lut_3027 ({sk[1075], i_30_, i_14_, i_13_, i_24_, i_32_, i_31_}, x1076x);
	defparam lut_3027.LUT_SIZE = 7;
	defparam lut_3027.mask = 128'h57ffffff57ffffff00000070000000f0;

	lut_sub lut_3031 ({sk[1076], i_12_, i_24_, i_17_, i_31_}, x1077x);
	defparam lut_3031.LUT_SIZE = 5;
	defparam lut_3031.mask = 32'h77770010;

	lut_sub lut_3033 ({sk[1077], i_38_, n_n1307, x49x, n_n1306, x257x, x70x}, x788x);
	defparam lut_3033.LUT_SIZE = 7;
	defparam lut_3033.mask = 128'h57ffffff57ffffff0055005500770377;

	lut_sub lut_3037 ({sk[1078], i_12_, i_24_, i_38_, n_n1307, n_n1303, x78x}, x1065x);
	defparam lut_3037.LUT_SIZE = 7;
	defparam lut_3037.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_3039 ({sk[1079], i_25_, x49x, n_n1225, x7492x, x313x, x7645x}, x7649x);
	defparam lut_3039.LUT_SIZE = 7;
	defparam lut_3039.mask = 128'h57ffffff57ffffff1111111f11111111;

	lut_sub lut_3042 ({sk[1080], i_8_, x49x, x70x, x1066x, x1067x, x7646x}, x7650x);
	defparam lut_3042.LUT_SIZE = 7;
	defparam lut_3042.mask = 128'h57ffffff57ffffff151515ff15151515;

	lut_sub lut_3046 ({sk[1081], i_32_, x788x, x1065x, x7649x, x7650x}, n_n1880);
	defparam lut_3046.LUT_SIZE = 6;
	defparam lut_3046.mask = 64'h3f3fffff7fff7f7f;

	lut_sub lut_3051 ({sk[1082], i_24_, x230x, x747x, x1052x, x1053x, x7660x}, n_n1884);
	defparam lut_3051.LUT_SIZE = 7;
	defparam lut_3051.mask = 128'h57ffffff57ffffff7f7f7fff7f7f7f7f;

	lut_sub lut_3056 ({sk[1083], i_7_, i_32_, i_33_, i_38_, x313x, x761x}, x760x);
	defparam lut_3056.LUT_SIZE = 7;
	defparam lut_3056.mask = 128'h57ffffff57ffffff0703050005000500;

	lut_sub lut_3059 ({sk[1084], i_12_, x376x, x395x, x1040x, x1044x, x7666x}, x7669x);
	defparam lut_3059.LUT_SIZE = 7;
	defparam lut_3059.mask = 128'h57ffffff57ffffff7f7f7fff7f7f7f7f;

	lut_sub lut_3064 ({sk[1085], n_n1443, n_n1429, x55x, x7675x, x7676x, x7677x}, x7680x);
	defparam lut_3064.LUT_SIZE = 7;
	defparam lut_3064.mask = 128'h57ffffff57ffffff7f7f7fff7fff7fff;

	lut_sub lut_3070 ({sk[1086], i_24_, x42x, n_n1438, n_n1437, n_n1459, x7692x}, x7696x);
	defparam lut_3070.LUT_SIZE = 7;
	defparam lut_3070.mask = 128'h57ffffff57ffffff1111111f11111111;

	lut_sub lut_3073 ({sk[1087], i_7_, i_8_, i_22_, n_n1454, n_n1431, x313x}, x795x);
	defparam lut_3073.LUT_SIZE = 7;
	defparam lut_3073.mask = 128'h57ffffff57ffffff5755030000000000;

	lut_sub lut_3076 ({sk[1088], i_8_, i_2_, x237x, x70x, x77x, n_n1459}, x7697x);
	defparam lut_3076.LUT_SIZE = 7;
	defparam lut_3076.mask = 128'h57ffffff57ffffff0357005503030000;

	lut_sub lut_3079 ({sk[1089], i_31_, i_33_, i_38_, n_n1397, x474x, x793x}, x7698x);
	defparam lut_3079.LUT_SIZE = 7;
	defparam lut_3079.mask = 128'h57ffffff57ffffff0003000005070505;

	lut_sub lut_3082 ({sk[1090], i_2_, i_38_, x7696x, x795x, x7697x, x7698x}, n_n1887);
	defparam lut_3082.LUT_SIZE = 7;
	defparam lut_3082.mask = 128'h57ffffff57ffffff77777fff777777ff;

	lut_sub lut_3087 ({sk[1091], i_8_, i_31_, x73x, n_n1489, n_n1197, x270x}, x1002x);
	defparam lut_3087.LUT_SIZE = 7;
	defparam lut_3087.mask = 128'h57ffffff57ffffff0507000005050000;

	lut_sub lut_3090 ({sk[1092], i_28_, i_22_, i_34_, i_35_, x1028x, x7686x}, x1025x);
	defparam lut_3090.LUT_SIZE = 7;
	defparam lut_3090.mask = 128'h57ffffff57ffffff0300070003000300;

	lut_sub lut_3093 ({sk[1093], i_14_, i_25_, n_n1393, n_n1419, x7683x, x7684x}, x7687x);
	defparam lut_3093.LUT_SIZE = 7;
	defparam lut_3093.mask = 128'h57ffffff57ffffff0505000005370033;

	lut_sub lut_3096 ({sk[1094], i_38_, n_n1458, n_n1497, n_n1459, x214x, x797x}, x7705x);
	defparam lut_3096.LUT_SIZE = 7;
	defparam lut_3096.mask = 128'h57ffffff57ffffff111111111111111f;

	lut_sub lut_3099 ({sk[1095], i_24_, n_n1361, x388x, x71x, x7701x, x7703x}, x7706x);
	defparam lut_3099.LUT_SIZE = 7;
	defparam lut_3099.mask = 128'h57ffffff57ffffff0033053700330033;

	lut_sub lut_3102 ({sk[1096], x7688x, x1002x, x1025x, x7687x, x7705x, x7706x}, x7709x);
	defparam lut_3102.LUT_SIZE = 7;
	defparam lut_3102.mask = 128'h57ffffff57ffffff7fffffffffffffff;

	lut_sub lut_3109 ({sk[1097], i_9_, i_3_, i_13_, i_11_, i_18_, i_19_}, x744x);
	defparam lut_3109.LUT_SIZE = 7;
	defparam lut_3109.mask = 128'h57ffffff57ffffff000000005f001300;

	lut_sub lut_3114 ({sk[1098], i_28_, i_25_, i_26_, i_35_, i_38_}, x370x);
	defparam lut_3114.LUT_SIZE = 6;
	defparam lut_3114.mask = 64'h3f3fffff40000000;

	lut_sub lut_3116 ({sk[1099], i_30_, i_28_, i_35_, i_38_, i_29_}, x7658x);
	defparam lut_3116.LUT_SIZE = 6;
	defparam lut_3116.mask = 64'h3f3fffff20000000;

	lut_sub lut_3118 ({sk[1100], i_29_, x3x, n_n1340, x271x, x370x, x7658x}, x747x);
	defparam lut_3118.LUT_SIZE = 7;
	defparam lut_3118.mask = 128'h57ffffff57ffffff3f7f00550f5f0055;

	lut_sub lut_3122 ({sk[1101], i_23_, i_21_, i_22_, n_n1404, n_n1408, x45x}, x1052x);
	defparam lut_3122.LUT_SIZE = 7;
	defparam lut_3122.mask = 128'h57ffffff57ffffff0000150000000000;

	lut_sub lut_3125 ({sk[1102], i_30_, x42x, n_n1353, n_n805, x81x, x7547x}, x1053x);
	defparam lut_3125.LUT_SIZE = 7;
	defparam lut_3125.mask = 128'h57ffffff57ffffff0005003700000000;

	lut_sub lut_3128 ({sk[1103], i_2_, n_n1438, x12x, x81x, x78x, x7656x}, x7660x);
	defparam lut_3128.LUT_SIZE = 7;
	defparam lut_3128.mask = 128'h57ffffff57ffffff0505053705050505;

	lut_sub lut_3131 ({sk[1104], i_28_, i_25_, i_26_, i_24_, i_35_, i_38_}, x375x);
	defparam lut_3131.LUT_SIZE = 7;
	defparam lut_3131.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_3133 ({sk[1105], i_28_, i_25_, i_32_, i_29_}, x7717x);
	defparam lut_3133.LUT_SIZE = 5;
	defparam lut_3133.mask = 32'h77778000;

	lut_sub lut_3135 ({sk[1106], i_28_, i_25_, i_32_, i_31_, i_34_, i_29_}, x7564x);
	defparam lut_3135.LUT_SIZE = 7;
	defparam lut_3135.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_3137 ({sk[1107], i_23_, x43x, n_n1141, x291x, x57x, x316x}, x1479x);
	defparam lut_3137.LUT_SIZE = 7;
	defparam lut_3137.mask = 128'h57ffffff57ffffff0101011101010101;

	lut_sub lut_3140 ({sk[1108], i_27_, n_n1443, x54x, n_n1429, n_n1489, x7108x}, x1480x);
	defparam lut_3140.LUT_SIZE = 7;
	defparam lut_3140.mask = 128'h57ffffff57ffffff0001001100000000;

	lut_sub lut_3143 ({sk[1109], i_30_, i_7_, i_8_, x260x, x324x, x7242x}, x1473x);
	defparam lut_3143.LUT_SIZE = 7;
	defparam lut_3143.mask = 128'h57ffffff57ffffff1511111100000000;

	lut_sub lut_3146 ({sk[1110], x47x, x67x, x29x, x470x, x7006x, x6999x}, x7244x);
	defparam lut_3146.LUT_SIZE = 7;
	defparam lut_3146.mask = 128'h57ffffff57ffffff0000030300550357;

	lut_sub lut_3149 ({sk[1111], i_33_, x1479x, x1480x, x1473x, x7244x}, n_n1712);
	defparam lut_3149.LUT_SIZE = 6;
	defparam lut_3149.mask = 64'h3f3fffff7fff7777;

	lut_sub lut_3154 ({sk[1112], i_7_, i_8_, i_22_, x73x, n_n1431, x466x}, x761x);
	defparam lut_3154.LUT_SIZE = 7;
	defparam lut_3154.mask = 128'h57ffffff57ffffff5755030000000000;

	lut_sub lut_3157 ({sk[1113], i_24_, i_38_, x58x, n_n1305, x49x, x321x}, x1040x);
	defparam lut_3157.LUT_SIZE = 7;
	defparam lut_3157.mask = 128'h57ffffff57ffffff0000000700000000;

	lut_sub lut_3160 ({sk[1114], i_12_, i_26_, i_24_, i_38_, n_n1302, x376x}, x1044x);
	defparam lut_3160.LUT_SIZE = 7;
	defparam lut_3160.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_3162 ({sk[1115], i_38_, n_n1353, x321x, x57x, x315x, x7665x}, x7666x);
	defparam lut_3162.LUT_SIZE = 7;
	defparam lut_3162.mask = 128'h57ffffff57ffffff0000030300550357;

	lut_sub lut_3165 ({sk[1116], n_n1408, x211x, x496x, x7055x, x7056x, x7054x}, x7057x);
	defparam lut_3165.LUT_SIZE = 7;
	defparam lut_3165.mask = 128'h57ffffff57ffffff0000005503030357;

	lut_sub lut_3168 ({sk[1117], i_20_, i_23_, i_24_, x211x, x496x, x7056x}, x770x);
	defparam lut_3168.LUT_SIZE = 7;
	defparam lut_3168.mask = 128'h57ffffff57ffffff5703030300000000;

	lut_sub lut_3171 ({sk[1118], i_27_, i_26_, i_23_, i_24_}, x7068x);
	defparam lut_3171.LUT_SIZE = 5;
	defparam lut_3171.mask = 32'h77778000;

	lut_sub lut_3173 ({sk[1119], i_27_, i_14_, i_26_, i_24_, i_16_}, x7066x);
	defparam lut_3173.LUT_SIZE = 6;
	defparam lut_3173.mask = 64'h3f3fffff80000000;

	lut_sub lut_3175 ({sk[1120], i_20_, i_14_, i_17_, i_16_}, x7070x);
	defparam lut_3175.LUT_SIZE = 5;
	defparam lut_3175.mask = 32'h77778000;

	lut_sub lut_3177 ({sk[1121], i_30_, i_28_, i_26_, i_24_, i_22_}, x466x);
	defparam lut_3177.LUT_SIZE = 6;
	defparam lut_3177.mask = 64'h3f3fffff80000000;

	lut_sub lut_3179 ({sk[1122], i_10_, i_32_, n_n1361, x389x, n_n1431, x313x}, x1167x);
	defparam lut_3179.LUT_SIZE = 7;
	defparam lut_3179.mask = 128'h57ffffff57ffffff0357030300000000;

	lut_sub lut_3182 ({sk[1123], i_30_, i_28_, i_22_, i_31_}, x7577x);
	defparam lut_3182.LUT_SIZE = 5;
	defparam lut_3182.mask = 32'h77778000;

	lut_sub lut_3184 ({sk[1124], i_8_, i_31_, n_n1361, x313x, x270x, x7577x}, x7578x);
	defparam lut_3184.LUT_SIZE = 7;
	defparam lut_3184.mask = 128'h57ffffff57ffffff111f111111111111;

	lut_sub lut_3187 ({sk[1125], i_31_, i_33_, i_29_, n_n1361, x50x, n_n1497}, x1161x);
	defparam lut_3187.LUT_SIZE = 7;
	defparam lut_3187.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_3189 ({sk[1126], i_24_, n_n1486, x51x, n_n1133, n_n1149, x375x}, x1162x);
	defparam lut_3189.LUT_SIZE = 7;
	defparam lut_3189.mask = 128'h57ffffff57ffffff0005003700050005;

	lut_sub lut_3192 ({sk[1127], n_n1197, n_n1288, x14x, x466x, x7572x, x7574x}, x7579x);
	defparam lut_3192.LUT_SIZE = 7;
	defparam lut_3192.mask = 128'h57ffffff57ffffff0000005503030357;

	lut_sub lut_3195 ({sk[1128], x68x, x1167x, x7578x, x1161x, x1162x, x7579x}, n_n1878);
	defparam lut_3195.LUT_SIZE = 7;
	defparam lut_3195.mask = 128'h57ffffff57ffffff7f7f7f7f7fffffff;

	lut_sub lut_3201 ({sk[1129], i_22_, n_n1438, n_n1197, n_n1523, n_n1497, x7466x}, x782x);
	defparam lut_3201.LUT_SIZE = 7;
	defparam lut_3201.mask = 128'h57ffffff57ffffff0005003700050005;

	lut_sub lut_3204 ({sk[1130], i_30_, i_28_, i_25_, i_26_, i_35_, i_38_}, x1066x);
	defparam lut_3204.LUT_SIZE = 7;
	defparam lut_3204.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_3206 ({sk[1131], i_30_, i_28_, i_26_, i_33_, i_35_, i_38_}, x1067x);
	defparam lut_3206.LUT_SIZE = 7;
	defparam lut_3206.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_3208 ({sk[1132], i_28_, i_26_, i_24_, i_32_, i_29_}, x7736x);
	defparam lut_3208.LUT_SIZE = 6;
	defparam lut_3208.mask = 64'h3f3fffff80000000;

	lut_sub lut_3210 ({sk[1133], i_28_, i_25_, i_24_, i_32_, i_34_, i_35_}, x7692x);
	defparam lut_3210.LUT_SIZE = 7;
	defparam lut_3210.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_3212 ({sk[1134], i_14_, i_28_, i_13_, i_12_, i_17_, i_22_}, x793x);
	defparam lut_3212.LUT_SIZE = 7;
	defparam lut_3212.mask = 128'h57ffffff57ffffff0101000001550000;

	lut_sub lut_3215 ({sk[1135], i_30_, i_14_, i_13_, i_12_, i_17_, i_32_}, x797x);
	defparam lut_3215.LUT_SIZE = 7;
	defparam lut_3215.mask = 128'h57ffffff57ffffff01010155030303ff;

	lut_sub lut_3220 ({sk[1136], i_9_, i_8_, i_3_, i_11_, i_18_}, x17x);
	defparam lut_3220.LUT_SIZE = 6;
	defparam lut_3220.mask = 64'h3f3fffff00003100;

	lut_sub lut_3223 ({sk[1137], i_13_, i_4_, i_12_, i_2_}, x7415x);
	defparam lut_3223.LUT_SIZE = 5;
	defparam lut_3223.mask = 32'h77778000;

	lut_sub lut_3225 ({sk[1138], i_28_, i_24_, i_33_, i_29_}, x7547x);
	defparam lut_3225.LUT_SIZE = 5;
	defparam lut_3225.mask = 32'h77778000;

	lut_sub lut_3227 ({sk[1139], i_9_, i_13_, i_11_, i_18_}, x436x);
	defparam lut_3227.LUT_SIZE = 5;
	defparam lut_3227.mask = 32'h77770010;

	lut_sub lut_3229 ({sk[1140], i_14_, i_13_, i_12_, i_17_, i_16_}, x805x);
	defparam lut_3229.LUT_SIZE = 6;
	defparam lut_3229.mask = 64'h3f3fffffa8a8a800;

	lut_sub lut_3234 ({sk[1141], i_32_, i_31_, i_29_}, x7026x);
	defparam lut_3234.LUT_SIZE = 4;
	defparam lut_3234.mask = 16'h5540;

	lut_sub lut_3236 ({sk[1142], i_8_, i_5_, i_6_, i_18_}, x7274x);
	defparam lut_3236.LUT_SIZE = 5;
	defparam lut_3236.mask = 32'h77778000;

	lut_sub lut_3238 ({sk[1143], i_20_, i_23_, i_24_}, x7055x);
	defparam lut_3238.LUT_SIZE = 4;
	defparam lut_3238.mask = 16'h5580;

	lut_sub lut_3240 ({sk[1144], i_30_, i_7_, i_8_, i_27_, i_28_, i_26_}, x7056x);
	defparam lut_3240.LUT_SIZE = 7;
	defparam lut_3240.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_3242 ({sk[1145], i_9_, i_3_, i_13_, i_11_}, x343x);
	defparam lut_3242.LUT_SIZE = 5;
	defparam lut_3242.mask = 32'h77770040;

	lut_sub lut_3244 ({sk[1146], i_20_, i_13_, i_12_, i_16_}, x402x);
	defparam lut_3244.LUT_SIZE = 5;
	defparam lut_3244.mask = 32'h77778000;

	lut_sub lut_3246 ({sk[1147], i_9_, i_8_, i_13_, i_12_, i_18_, i_19_}, x414x);
	defparam lut_3246.LUT_SIZE = 7;
	defparam lut_3246.mask = 128'h57ffffff57ffffff0000000001000000;

	lut_sub lut_3248 ({sk[1148], i_7_, i_5_, i_6_, i_3_, i_4_, i_0_}, x7253x);
	defparam lut_3248.LUT_SIZE = 7;
	defparam lut_3248.mask = 128'h57ffffff57ffffff0800000000000000;

	lut_sub lut_3250 ({sk[1149], i_20_, i_29_, n_n1441, x54x, x413x, x7253x}, x1471x);
	defparam lut_3250.LUT_SIZE = 7;
	defparam lut_3250.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_3252 ({sk[1150], i_20_, x54x, n_n1303, n_n245, x431x, x44x}, x1472x);
	defparam lut_3252.LUT_SIZE = 7;
	defparam lut_3252.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_3254 ({sk[1151], i_9_, i_7_, i_14_, i_13_}, x557x);
	defparam lut_3254.LUT_SIZE = 5;
	defparam lut_3254.mask = 32'h77770e00;

	lut_sub lut_3257 ({sk[1152], i_3_, i_13_, i_11_, i_18_, i_22_, i_19_}, x582x);
	defparam lut_3257.LUT_SIZE = 7;
	defparam lut_3257.mask = 128'h57ffffff57ffffff444c0000040c0000;

	lut_sub lut_3261 ({sk[1153], i_13_, i_12_, i_11_, i_19_}, x590x);
	defparam lut_3261.LUT_SIZE = 5;
	defparam lut_3261.mask = 32'h77770700;

	lut_sub lut_3264 ({sk[1154], i_13_, i_12_, i_11_, i_19_}, x593x);
	defparam lut_3264.LUT_SIZE = 5;
	defparam lut_3264.mask = 32'h77770700;

	lut_sub lut_3267 ({sk[1155], i_13_, i_12_, i_11_, i_18_, i_19_}, x596x);
	defparam lut_3267.LUT_SIZE = 6;
	defparam lut_3267.mask = 64'h3f3fffff00130000;

	lut_sub lut_3270 ({sk[1156], i_3_, i_13_, i_12_, i_19_}, x7298x);
	defparam lut_3270.LUT_SIZE = 5;
	defparam lut_3270.mask = 32'h77771000;

	lut_sub lut_3272 ({sk[1157], i_10_, x13x, x205x, x210x, x596x, x7298x}, x595x);
	defparam lut_3272.LUT_SIZE = 7;
	defparam lut_3272.mask = 128'h57ffffff57ffffff0000000f0000007f;

	lut_sub lut_3276 ({sk[1158], i_9_, i_8_, i_5_, i_6_}, x6891x);
	defparam lut_3276.LUT_SIZE = 5;
	defparam lut_3276.mask = 32'h77778000;

	lut_sub lut_3278 ({sk[1159], i_7_, i_5_, i_6_, i_32_, i_33_, i_37_}, x1751x);
	defparam lut_3278.LUT_SIZE = 7;
	defparam lut_3278.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_3280 ({sk[1160], i_8_, i_5_, i_6_, i_33_, i_35_, i_37_}, x1752x);
	defparam lut_3280.LUT_SIZE = 7;
	defparam lut_3280.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_3282 ({sk[1161], i_9_, i_8_, i_6_, i_33_, i_35_, i_37_}, x7131x);
	defparam lut_3282.LUT_SIZE = 7;
	defparam lut_3282.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_3284 ({sk[1162], i_9_, i_13_, i_18_, n_n1118, x76x, x213x}, x7438x);
	defparam lut_3284.LUT_SIZE = 7;
	defparam lut_3284.mask = 128'h57ffffff57ffffff0000000005370505;

	lut_sub lut_3287 ({sk[1163], i_7_, i_14_, i_13_, i_12_}, x661x);
	defparam lut_3287.LUT_SIZE = 5;
	defparam lut_3287.mask = 32'h777700a8;

	lut_sub lut_3290 ({sk[1164], i_20_, i_13_, i_12_, i_23_, i_17_, i_16_}, x666x);
	defparam lut_3290.LUT_SIZE = 7;
	defparam lut_3290.mask = 128'h57ffffff57ffffffa080000000000000;

	lut_sub lut_3293 ({sk[1165], i_3_, i_13_, i_12_, i_11_, i_18_, i_22_}, x679x);
	defparam lut_3293.LUT_SIZE = 7;
	defparam lut_3293.mask = 128'h57ffffff57ffffff000a000000020000;

	lut_sub lut_3296 ({sk[1166], i_20_, i_13_, i_12_, i_17_, i_16_}, x683x);
	defparam lut_3296.LUT_SIZE = 6;
	defparam lut_3296.mask = 64'h3f3fffffa8000000;

	lut_sub lut_3299 ({sk[1167], i_13_, i_17_, i_16_, i_32_}, x7153x);
	defparam lut_3299.LUT_SIZE = 5;
	defparam lut_3299.mask = 32'h77778000;

	lut_sub lut_3301 ({sk[1168], i_9_, i_8_, i_3_, i_11_, i_18_, i_19_}, x737x);
	defparam lut_3301.LUT_SIZE = 7;
	defparam lut_3301.mask = 128'h57ffffff57ffffff000000005f030000;

	lut_sub lut_3305 ({sk[1169], i_3_, i_13_, i_11_, i_18_, i_22_, i_19_}, x764x);
	defparam lut_3305.LUT_SIZE = 7;
	defparam lut_3305.mask = 128'h57ffffff57ffffff444c0000040c0000;

	lut_sub lut_3309 ({sk[1170], i_20_, i_14_, i_17_, i_16_}, x7054x);
	defparam lut_3309.LUT_SIZE = 5;
	defparam lut_3309.mask = 32'h77778000;

	lut_sub lut_3311 ({sk[1171], i_7_, i_11_, i_23_, i_21_, i_19_}, x8083x);
	defparam lut_3311.LUT_SIZE = 6;
	defparam lut_3311.mask = 64'h3f3fffff80000000;

	lut_sub lut_3313 ({sk[1172], i_36_, x232x, n_n1443, n_n1369, n_n460, x8083x}, x6x);
	defparam lut_3313.LUT_SIZE = 7;
	defparam lut_3313.mask = 128'h57ffffff57ffffff0000000000000001;

	lut_sub lut_3315 ({sk[1173], i_27_, i_28_, i_23_, i_36_, i_29_, n_n1397}, x8085x);
	defparam lut_3315.LUT_SIZE = 7;
	defparam lut_3315.mask = 128'h57ffffff57ffffff0400000000000000;

	lut_sub lut_3317 ({sk[1174], i_13_, i_23_, i_17_, i_21_, i_16_}, x8070x);
	defparam lut_3317.LUT_SIZE = 6;
	defparam lut_3317.mask = 64'h3f3fffff80000000;

	lut_sub lut_3319 ({sk[1175], i_14_, i_12_, i_23_, i_21_, i_16_}, x8064x);
	defparam lut_3319.LUT_SIZE = 6;
	defparam lut_3319.mask = 64'h3f3fffff80000000;

	lut_sub lut_3321 ({sk[1176], i_9_, i_7_, i_13_, i_12_, i_23_, i_16_}, x8066x);
	defparam lut_3321.LUT_SIZE = 7;
	defparam lut_3321.mask = 128'h57ffffff57ffffff0000800000000000;

	lut_sub lut_3323 ({sk[1177], i_9_, i_7_, i_14_, i_12_, i_23_, i_16_}, x8058x);
	defparam lut_3323.LUT_SIZE = 7;
	defparam lut_3323.mask = 128'h57ffffff57ffffff0000800000000000;

	lut_sub lut_3325 ({sk[1178], i_27_, i_28_, i_26_, i_36_, i_35_}, x8018x);
	defparam lut_3325.LUT_SIZE = 6;
	defparam lut_3325.mask = 64'h3f3fffff20000000;

	lut_sub lut_3327 ({sk[1179], i_9_, i_7_, i_14_, i_12_, i_16_}, x7995x);
	defparam lut_3327.LUT_SIZE = 6;
	defparam lut_3327.mask = 64'h3f3fffff00800000;

	lut_sub lut_3329 ({sk[1180], i_9_, i_7_, i_13_, i_31_, i_34_, i_35_}, x7996x);
	defparam lut_3329.LUT_SIZE = 7;
	defparam lut_3329.mask = 128'h57ffffff57ffffff0000040000000000;

	lut_sub lut_3331 ({sk[1181], i_9_, i_7_, i_14_, i_31_, i_34_, i_35_}, x7987x);
	defparam lut_3331.LUT_SIZE = 7;
	defparam lut_3331.mask = 128'h57ffffff57ffffff0000040000000000;

	lut_sub lut_3333 ({sk[1182], i_20_, i_28_, i_21_, i_29_}, x7969x);
	defparam lut_3333.LUT_SIZE = 5;
	defparam lut_3333.mask = 32'h77770040;

	lut_sub lut_3335 ({sk[1183], i_27_, i_28_, i_24_, i_34_, i_33_}, x7972x);
	defparam lut_3335.LUT_SIZE = 6;
	defparam lut_3335.mask = 64'h3f3fffff10000000;

	lut_sub lut_3337 ({sk[1184], i_14_, i_13_, i_23_, i_17_, i_21_, i_16_}, x7973x);
	defparam lut_3337.LUT_SIZE = 7;
	defparam lut_3337.mask = 128'h57ffffff57ffffff0000000020000000;

	lut_sub lut_3339 ({sk[1185], i_27_, i_28_, i_26_, i_23_, i_24_, i_31_}, x7974x);
	defparam lut_3339.LUT_SIZE = 7;
	defparam lut_3339.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_3341 ({sk[1186], i_13_, i_2_, i_17_, i_16_, i_36_}, x7957x);
	defparam lut_3341.LUT_SIZE = 6;
	defparam lut_3341.mask = 64'h3f3fffff40000000;

	lut_sub lut_3343 ({sk[1187], i_2_, i_17_, i_21_, i_16_, i_36_}, x7961x);
	defparam lut_3343.LUT_SIZE = 6;
	defparam lut_3343.mask = 64'h3f3fffff40000000;

	lut_sub lut_3345 ({sk[1188], i_27_, i_28_, i_26_, i_33_}, x7932x);
	defparam lut_3345.LUT_SIZE = 5;
	defparam lut_3345.mask = 32'h77774000;

	lut_sub lut_3347 ({sk[1189], i_30_, i_28_, i_26_, i_24_, i_34_, i_29_}, x7925x);
	defparam lut_3347.LUT_SIZE = 7;
	defparam lut_3347.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_3349 ({sk[1190], i_32_, i_31_, i_34_, i_36_, i_35_}, x7884x);
	defparam lut_3349.LUT_SIZE = 6;
	defparam lut_3349.mask = 64'h3f3fffff02000000;

	lut_sub lut_3351 ({sk[1191], i_16_, i_34_, i_36_, i_29_, x242x, n_n1216}, x7878x);
	defparam lut_3351.LUT_SIZE = 7;
	defparam lut_3351.mask = 128'h57ffffff57ffffff0000001000000000;

	lut_sub lut_3353 ({sk[1192], i_27_, x54x, n_n1408, x50x, n_n1128, x86x}, x852x);
	defparam lut_3353.LUT_SIZE = 7;
	defparam lut_3353.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_3355 ({sk[1193], i_31_, n_n1216, x243x, x51x, x260x, x86x}, x853x);
	defparam lut_3355.LUT_SIZE = 7;
	defparam lut_3355.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_3357 ({sk[1194], i_17_, i_21_, i_16_, i_32_, i_36_, i_35_}, x7862x);
	defparam lut_3357.LUT_SIZE = 7;
	defparam lut_3357.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_3359 ({sk[1195], i_14_, i_13_, i_26_, i_23_, i_24_}, x7858x);
	defparam lut_3359.LUT_SIZE = 6;
	defparam lut_3359.mask = 64'h3f3fffff80808000;

	lut_sub lut_3362 ({sk[1196], i_9_, i_10_, i_5_, i_6_, i_13_, i_4_}, x7861x);
	defparam lut_3362.LUT_SIZE = 7;
	defparam lut_3362.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_3364 ({sk[1197], i_27_, i_28_, i_31_}, x7857x);
	defparam lut_3364.LUT_SIZE = 4;
	defparam lut_3364.mask = 16'h5580;

	lut_sub lut_3366 ({sk[1198], i_5_, i_6_, i_4_, i_31_}, x7847x);
	defparam lut_3366.LUT_SIZE = 5;
	defparam lut_3366.mask = 32'h77778000;

	lut_sub lut_3368 ({sk[1199], i_9_, i_3_, i_11_, i_2_, i_18_, i_19_}, x7817x);
	defparam lut_3368.LUT_SIZE = 7;
	defparam lut_3368.mask = 128'h57ffffff57ffffff0a000e0c00000000;

	lut_sub lut_3371 ({sk[1200], i_13_, i_31_, i_36_, i_35_}, x7820x);
	defparam lut_3371.LUT_SIZE = 5;
	defparam lut_3371.mask = 32'h77772000;

	lut_sub lut_3373 ({sk[1201], i_20_, i_26_, i_24_, i_21_}, x7798x);
	defparam lut_3373.LUT_SIZE = 5;
	defparam lut_3373.mask = 32'h77770080;

	lut_sub lut_3375 ({sk[1202], i_7_, i_8_, i_14_, i_23_, i_17_, i_16_}, x7800x);
	defparam lut_3375.LUT_SIZE = 7;
	defparam lut_3375.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_3377 ({sk[1203], i_28_, i_24_, i_34_, i_29_}, x7782x);
	defparam lut_3377.LUT_SIZE = 5;
	defparam lut_3377.mask = 32'h77771000;

	lut_sub lut_3379 ({sk[1204], i_30_, i_20_, i_23_, i_21_, i_32_, i_31_}, x7783x);
	defparam lut_3379.LUT_SIZE = 7;
	defparam lut_3379.mask = 128'h57ffffff57ffffff0000800000000000;

	lut_sub lut_3381 ({sk[1205], i_8_, i_36_, i_35_}, x7772x);
	defparam lut_3381.LUT_SIZE = 4;
	defparam lut_3381.mask = 16'h5520;

	lut_sub lut_3383 ({sk[1206], i_27_, i_28_, i_13_, i_17_, i_16_, i_29_}, x7764x);
	defparam lut_3383.LUT_SIZE = 7;
	defparam lut_3383.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_3385 ({sk[1207], i_13_, i_32_, i_36_, i_35_}, x7750x);
	defparam lut_3385.LUT_SIZE = 5;
	defparam lut_3385.mask = 32'h77772000;

	lut_sub lut_3387 ({sk[1208], i_28_, i_25_, i_26_, i_35_, i_38_, i_29_}, x7732x);
	defparam lut_3387.LUT_SIZE = 7;
	defparam lut_3387.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_3389 ({sk[1209], i_30_, i_2_, i_32_, i_33_, i_35_, i_38_}, x7724x);
	defparam lut_3389.LUT_SIZE = 7;
	defparam lut_3389.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_3391 ({sk[1210], i_30_, i_7_, i_2_, i_32_}, x7701x);
	defparam lut_3391.LUT_SIZE = 5;
	defparam lut_3391.mask = 32'h77778000;

	lut_sub lut_3393 ({sk[1211], i_30_, i_8_, i_31_}, x7703x);
	defparam lut_3393.LUT_SIZE = 4;
	defparam lut_3393.mask = 16'h5580;

	lut_sub lut_3395 ({sk[1212], i_30_, i_7_, i_28_, i_32_, i_29_}, x7684x);
	defparam lut_3395.LUT_SIZE = 6;
	defparam lut_3395.mask = 64'h3f3fffff80000000;

	lut_sub lut_3397 ({sk[1213], i_30_, i_12_, i_17_, i_32_}, x7686x);
	defparam lut_3397.LUT_SIZE = 5;
	defparam lut_3397.mask = 32'h77770103;

	lut_sub lut_3400 ({sk[1214], i_9_, i_10_, i_28_, i_26_, i_24_, i_29_}, x7674x);
	defparam lut_3400.LUT_SIZE = 7;
	defparam lut_3400.mask = 128'h57ffffff57ffffff0000000080000000;

	lut_sub lut_3402 ({sk[1215], i_28_, i_25_, i_26_, i_24_, i_32_, i_29_}, x7665x);
	defparam lut_3402.LUT_SIZE = 7;
	defparam lut_3402.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_3404 ({sk[1216], i_30_, i_8_, i_28_, i_2_, i_22_, i_31_}, x7656x);
	defparam lut_3404.LUT_SIZE = 7;
	defparam lut_3404.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_3406 ({sk[1217], i_9_, i_10_, i_2_, i_32_, i_35_, i_38_}, x7645x);
	defparam lut_3406.LUT_SIZE = 7;
	defparam lut_3406.mask = 128'h57ffffff57ffffff0000000040000000;

	lut_sub lut_3408 ({sk[1218], i_9_, i_10_, i_8_, i_2_, i_24_, i_22_}, x7646x);
	defparam lut_3408.LUT_SIZE = 7;
	defparam lut_3408.mask = 128'h57ffffff57ffffff0000000080000000;

	lut_sub lut_3410 ({sk[1219], i_30_, i_28_, i_26_, i_32_}, x7627x);
	defparam lut_3410.LUT_SIZE = 5;
	defparam lut_3410.mask = 32'h777740c0;

	lut_sub lut_3413 ({sk[1220], i_24_, i_34_, i_33_, i_38_}, x7616x);
	defparam lut_3413.LUT_SIZE = 5;
	defparam lut_3413.mask = 32'h77770400;

	lut_sub lut_3415 ({sk[1221], i_30_, i_7_, i_28_, i_32_, i_29_}, x7617x);
	defparam lut_3415.LUT_SIZE = 6;
	defparam lut_3415.mask = 64'h3f3fffff80000000;

	lut_sub lut_3417 ({sk[1222], i_28_, i_22_, i_34_, i_35_}, x7618x);
	defparam lut_3417.LUT_SIZE = 5;
	defparam lut_3417.mask = 32'h77770400;

	lut_sub lut_3419 ({sk[1223], i_28_, i_22_, i_31_, i_34_}, x7619x);
	defparam lut_3419.LUT_SIZE = 5;
	defparam lut_3419.mask = 32'h77770100;

	lut_sub lut_3421 ({sk[1224], i_7_, i_8_, i_24_, i_38_}, x7600x);
	defparam lut_3421.LUT_SIZE = 5;
	defparam lut_3421.mask = 32'h77774000;

	lut_sub lut_3423 ({sk[1225], i_20_, i_28_, i_22_, i_34_, i_35_, i_29_}, x1134x);
	defparam lut_3423.LUT_SIZE = 7;
	defparam lut_3423.mask = 128'h57ffffff57ffffff0000000010000000;

	lut_sub lut_3425 ({sk[1226], i_29_, x76x, n_n1128, n_n1497, x226x, x81x}, x1139x);
	defparam lut_3425.LUT_SIZE = 7;
	defparam lut_3425.mask = 128'h57ffffff57ffffff0000035700000055;

	lut_sub lut_3428 ({sk[1227], i_24_, x11x, n_n1486, n_n1133, n_n1149, x375x}, x1141x);
	defparam lut_3428.LUT_SIZE = 7;
	defparam lut_3428.mask = 128'h57ffffff57ffffff0000053700000505;

	lut_sub lut_3431 ({sk[1228], i_30_, i_9_, i_10_, i_8_, i_12_}, x7583x);
	defparam lut_3431.LUT_SIZE = 6;
	defparam lut_3431.mask = 64'h3f3fffff00400000;

	lut_sub lut_3433 ({sk[1229], i_13_, i_26_, i_24_, i_33_, i_38_}, x7584x);
	defparam lut_3433.LUT_SIZE = 6;
	defparam lut_3433.mask = 64'h3f3fffff00004000;

	lut_sub lut_3435 ({sk[1230], i_9_, i_10_, i_8_, i_12_}, x7572x);
	defparam lut_3435.LUT_SIZE = 5;
	defparam lut_3435.mask = 32'h77770040;

	lut_sub lut_3437 ({sk[1231], i_10_, i_26_, i_24_, i_33_, i_38_}, x7574x);
	defparam lut_3437.LUT_SIZE = 6;
	defparam lut_3437.mask = 64'h3f3fffff40000000;

	lut_sub lut_3439 ({sk[1232], i_28_, i_25_, i_34_, i_35_, i_38_, i_29_}, x7556x);
	defparam lut_3439.LUT_SIZE = 7;
	defparam lut_3439.mask = 128'h57ffffff57ffffff0200000000000000;

	lut_sub lut_3441 ({sk[1233], i_30_, i_32_, i_35_, i_38_}, x7559x);
	defparam lut_3441.LUT_SIZE = 5;
	defparam lut_3441.mask = 32'h77774000;

	lut_sub lut_3443 ({sk[1234], i_28_, i_25_, i_26_, i_24_, i_19_, i_29_}, x7558x);
	defparam lut_3443.LUT_SIZE = 7;
	defparam lut_3443.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_3445 ({sk[1235], i_24_, x71x, x18x, x436x, x7559x, x7558x}, x1172x);
	defparam lut_3445.LUT_SIZE = 7;
	defparam lut_3445.mask = 128'h57ffffff57ffffff0011031300110011;

	lut_sub lut_3448 ({sk[1236], i_30_, i_9_, i_3_, i_13_, i_11_, i_24_}, x7560x);
	defparam lut_3448.LUT_SIZE = 7;
	defparam lut_3448.mask = 128'h57ffffff57ffffff0000200000000000;

	lut_sub lut_3450 ({sk[1237], i_28_, i_25_, i_32_, i_34_, i_35_, i_29_}, x7562x);
	defparam lut_3450.LUT_SIZE = 7;
	defparam lut_3450.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_3452 ({sk[1238], i_30_, i_24_, i_33_, i_35_, i_38_}, x7542x);
	defparam lut_3452.LUT_SIZE = 6;
	defparam lut_3452.mask = 64'h3f3fffff40000000;

	lut_sub lut_3454 ({sk[1239], i_28_, i_34_, i_33_, i_38_, i_29_}, x7535x);
	defparam lut_3454.LUT_SIZE = 6;
	defparam lut_3454.mask = 64'h3f3fffff00200000;

	lut_sub lut_3456 ({sk[1240], i_10_, i_13_, i_25_, i_24_, i_34_, i_38_}, x7516x);
	defparam lut_3456.LUT_SIZE = 7;
	defparam lut_3456.mask = 128'h57ffffff57ffffff1000100000001000;

	lut_sub lut_3459 ({sk[1241], i_8_, i_28_, i_25_, i_34_, i_35_, i_29_}, x7519x);
	defparam lut_3459.LUT_SIZE = 7;
	defparam lut_3459.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_3461 ({sk[1242], i_28_, i_34_, i_33_, i_38_, i_29_}, x7520x);
	defparam lut_3461.LUT_SIZE = 6;
	defparam lut_3461.mask = 64'h3f3fffff00200000;

	lut_sub lut_3463 ({sk[1243], i_28_, i_25_, i_34_, i_38_, i_29_}, x7509x);
	defparam lut_3463.LUT_SIZE = 6;
	defparam lut_3463.mask = 64'h3f3fffff02000000;

	lut_sub lut_3465 ({sk[1244], i_30_, i_9_, i_10_, i_28_, i_2_, i_32_}, x7489x);
	defparam lut_3465.LUT_SIZE = 7;
	defparam lut_3465.mask = 128'h57ffffff57ffffff0000800000000000;

	lut_sub lut_3467 ({sk[1245], x204x, x52x, x264x, x404x, x41x, x7274x}, x1238x);
	defparam lut_3467.LUT_SIZE = 7;
	defparam lut_3467.mask = 128'h57ffffff57ffffff0000000500000037;

	lut_sub lut_3470 ({sk[1246], i_25_, i_11_, i_34_, i_19_, i_35_, i_38_}, x7480x);
	defparam lut_3470.LUT_SIZE = 7;
	defparam lut_3470.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_3472 ({sk[1247], n_n1307, n_n787, x7314x, x361x, x78x, x353x}, x1241x);
	defparam lut_3472.LUT_SIZE = 7;
	defparam lut_3472.mask = 128'h57ffffff57ffffff0000001100030013;

	lut_sub lut_3475 ({sk[1248], x11x, x213x, x7425x, x7426x, n_n1497, x7444x}, x1242x);
	defparam lut_3475.LUT_SIZE = 7;
	defparam lut_3475.mask = 128'h57ffffff57ffffff0000001101010111;

	lut_sub lut_3478 ({sk[1249], i_30_, i_13_, i_24_, x271x, x454x, x17x}, x1325x);
	defparam lut_3478.LUT_SIZE = 7;
	defparam lut_3478.mask = 128'h57ffffff57ffffff0700030000000000;

	lut_sub lut_3481 ({sk[1250], i_10_, i_28_, i_31_, i_29_, x41x, x238x}, x1353x);
	defparam lut_3481.LUT_SIZE = 7;
	defparam lut_3481.mask = 128'h57ffffff57ffffff1000000000000000;

	lut_sub lut_3483 ({sk[1251], i_28_, i_32_, i_31_, n_n1307, n_n853, x389x}, x1355x);
	defparam lut_3483.LUT_SIZE = 7;
	defparam lut_3483.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_3485 ({sk[1252], i_13_, i_35_, i_38_, x42x, x14x, n_n1311}, x1358x);
	defparam lut_3485.LUT_SIZE = 7;
	defparam lut_3485.mask = 128'h57ffffff57ffffff0000000000000001;

	lut_sub lut_3487 ({sk[1253], i_32_, i_33_, i_35_, i_38_}, x7328x);
	defparam lut_3487.LUT_SIZE = 5;
	defparam lut_3487.mask = 32'h77774000;

	lut_sub lut_3489 ({sk[1254], i_28_, i_25_, i_26_, i_31_, i_35_, i_38_}, x7330x);
	defparam lut_3489.LUT_SIZE = 7;
	defparam lut_3489.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_3491 ({sk[1255], i_28_, i_25_, i_26_, i_32_, i_35_, i_38_}, x7321x);
	defparam lut_3491.LUT_SIZE = 7;
	defparam lut_3491.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_3493 ({sk[1256], i_10_, i_13_, i_12_, i_18_, i_19_}, x7306x);
	defparam lut_3493.LUT_SIZE = 6;
	defparam lut_3493.mask = 64'h3f3fffff00000100;

	lut_sub lut_3495 ({sk[1257], i_10_, i_13_, i_12_, i_11_, i_18_}, x7294x);
	defparam lut_3495.LUT_SIZE = 6;
	defparam lut_3495.mask = 64'h3f3fffff00000100;

	lut_sub lut_3497 ({sk[1258], i_30_, i_28_, i_25_, i_26_, i_38_}, x7300x);
	defparam lut_3497.LUT_SIZE = 6;
	defparam lut_3497.mask = 64'h3f3fffff40000000;

	lut_sub lut_3499 ({sk[1259], i_9_, i_12_, n_n1431, x23x, x81x, x1442x}, x1437x);
	defparam lut_3499.LUT_SIZE = 7;
	defparam lut_3499.mask = 128'h57ffffff57ffffff0011001100110013;

	lut_sub lut_3502 ({sk[1260], i_28_, i_25_, i_26_, i_24_, i_22_, i_38_}, x7286x);
	defparam lut_3502.LUT_SIZE = 7;
	defparam lut_3502.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_3504 ({sk[1261], i_9_, i_8_, i_13_, i_12_, i_11_, i_18_}, x1445x);
	defparam lut_3504.LUT_SIZE = 7;
	defparam lut_3504.mask = 128'h57ffffff57ffffff0000000001000000;

	lut_sub lut_3506 ({sk[1262], n_n1038, n_n1523, x7287x, x414x, x593x, x1445x}, x1439x);
	defparam lut_3506.LUT_SIZE = 7;
	defparam lut_3506.mask = 128'h57ffffff57ffffff0000005f0000007f;

	lut_sub lut_3510 ({sk[1263], i_9_, i_8_, i_13_, i_12_, i_11_, i_18_}, x1452x);
	defparam lut_3510.LUT_SIZE = 7;
	defparam lut_3510.mask = 128'h57ffffff57ffffff0000000001000000;

	lut_sub lut_3512 ({sk[1264], i_9_, i_28_, i_12_, i_26_, i_24_}, x7261x);
	defparam lut_3512.LUT_SIZE = 6;
	defparam lut_3512.mask = 64'h3f3fffff00000800;

	lut_sub lut_3514 ({sk[1265], i_27_, i_28_, i_34_, i_35_, i_29_, i_37_}, x7242x);
	defparam lut_3514.LUT_SIZE = 7;
	defparam lut_3514.mask = 128'h57ffffff57ffffff0400000000000000;

	lut_sub lut_3516 ({sk[1266], i_20_, x54x, n_n1118, n_n152, x461x, x44x}, x1481x);
	defparam lut_3516.LUT_SIZE = 7;
	defparam lut_3516.mask = 128'h57ffffff57ffffff0000000100000000;

	lut_sub lut_3518 ({sk[1267], i_13_, i_32_, i_33_, i_35_, i_37_}, x7226x);
	defparam lut_3518.LUT_SIZE = 6;
	defparam lut_3518.mask = 64'h3f3fffff40000000;

	lut_sub lut_3520 ({sk[1268], i_20_, i_17_, i_16_, x46x, x7213x, x7226x}, x1482x);
	defparam lut_3520.LUT_SIZE = 7;
	defparam lut_3520.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_3522 ({sk[1269], i_13_, i_17_, i_16_, i_32_, i_33_, i_29_}, x7227x);
	defparam lut_3522.LUT_SIZE = 7;
	defparam lut_3522.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_3524 ({sk[1270], x366x, x7145x, x7146x, x7148x, x7149x, x7227x}, x1483x);
	defparam lut_3524.LUT_SIZE = 7;
	defparam lut_3524.mask = 128'h57ffffff57ffffff0000000001010155;

	lut_sub lut_3527 ({sk[1271], i_28_, i_33_, i_29_, x269x}, x7229x);
	defparam lut_3527.LUT_SIZE = 5;
	defparam lut_3527.mask = 32'h77774000;

	lut_sub lut_3529 ({sk[1272], i_27_, i_28_, i_24_, i_37_}, x7208x);
	defparam lut_3529.LUT_SIZE = 5;
	defparam lut_3529.mask = 32'h77774000;

	lut_sub lut_3531 ({sk[1273], i_23_, i_17_, i_16_, i_34_, i_33_, i_29_}, x7209x);
	defparam lut_3531.LUT_SIZE = 7;
	defparam lut_3531.mask = 128'h57ffffff57ffffff0800000000000000;

	lut_sub lut_3533 ({sk[1274], i_8_, i_5_, i_6_, i_23_, i_18_, i_17_}, x7196x);
	defparam lut_3533.LUT_SIZE = 7;
	defparam lut_3533.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_3535 ({sk[1275], i_11_, i_23_, i_17_, i_19_}, x7197x);
	defparam lut_3535.LUT_SIZE = 5;
	defparam lut_3535.mask = 32'h77778000;

	lut_sub lut_3537 ({sk[1276], i_14_, i_28_, i_16_, i_29_}, x7211x);
	defparam lut_3537.LUT_SIZE = 5;
	defparam lut_3537.mask = 32'h77778000;

	lut_sub lut_3539 ({sk[1277], i_14_, i_32_, i_35_, i_37_}, x7215x);
	defparam lut_3539.LUT_SIZE = 5;
	defparam lut_3539.mask = 32'h77774000;

	lut_sub lut_3541 ({sk[1278], i_14_, i_16_, i_34_, i_35_, i_37_}, x7198x);
	defparam lut_3541.LUT_SIZE = 6;
	defparam lut_3541.mask = 64'h3f3fffff04000000;

	lut_sub lut_3543 ({sk[1279], i_7_, i_5_, i_6_, i_4_, i_1_, i_0_}, x7202x);
	defparam lut_3543.LUT_SIZE = 7;
	defparam lut_3543.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_3545 ({sk[1280], i_34_, i_33_, i_37_}, x7188x);
	defparam lut_3545.LUT_SIZE = 4;
	defparam lut_3545.mask = 16'h5504;

	lut_sub lut_3547 ({sk[1281], i_34_, i_35_, i_37_}, x7175x);
	defparam lut_3547.LUT_SIZE = 4;
	defparam lut_3547.mask = 16'h5510;

	lut_sub lut_3549 ({sk[1282], i_27_, i_28_, i_23_, i_32_, i_29_}, x7173x);
	defparam lut_3549.LUT_SIZE = 6;
	defparam lut_3549.mask = 64'h3f3fffff80000000;

	lut_sub lut_3551 ({sk[1283], i_27_, i_28_, i_23_, i_17_, i_29_}, x7174x);
	defparam lut_3551.LUT_SIZE = 6;
	defparam lut_3551.mask = 64'h3f3fffff80000000;

	lut_sub lut_3553 ({sk[1284], i_27_, i_28_, i_13_, i_17_, i_16_, i_29_}, x7150x);
	defparam lut_3553.LUT_SIZE = 7;
	defparam lut_3553.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_3555 ({sk[1285], i_9_, i_10_, i_6_, i_32_}, x7119x);
	defparam lut_3555.LUT_SIZE = 5;
	defparam lut_3555.mask = 32'h77778000;

	lut_sub lut_3557 ({sk[1286], i_30_, i_34_, i_33_, i_35_, i_37_}, x7114x);
	defparam lut_3557.LUT_SIZE = 6;
	defparam lut_3557.mask = 64'h3f3fffff00400000;

	lut_sub lut_3559 ({sk[1287], i_30_, i_33_, i_35_, i_29_, i_37_}, x7106x);
	defparam lut_3559.LUT_SIZE = 6;
	defparam lut_3559.mask = 64'h3f3fffff40000000;

	lut_sub lut_3561 ({sk[1288], i_8_, n_n1441, x43x, x74x, x348x, x7106x}, x1587x);
	defparam lut_3561.LUT_SIZE = 7;
	defparam lut_3561.mask = 128'h57ffffff57ffffff0005111500001111;

	lut_sub lut_3564 ({sk[1289], i_32_, i_34_, i_33_, i_35_, i_37_}, x7078x);
	defparam lut_3564.LUT_SIZE = 6;
	defparam lut_3564.mask = 64'h3f3fffff10000000;

	lut_sub lut_3566 ({sk[1290], i_30_, i_27_, i_28_, i_29_}, x7080x);
	defparam lut_3566.LUT_SIZE = 5;
	defparam lut_3566.mask = 32'h77778000;

	lut_sub lut_3568 ({sk[1291], i_0_, i_33_, i_35_, i_37_}, x7084x);
	defparam lut_3568.LUT_SIZE = 5;
	defparam lut_3568.mask = 32'h77774000;

	lut_sub lut_3570 ({sk[1292], i_30_, i_27_, i_28_, i_26_, i_24_, i_32_}, x7082x);
	defparam lut_3570.LUT_SIZE = 7;
	defparam lut_3570.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_3572 ({sk[1293], i_20_, i_13_, i_17_, i_16_}, x7083x);
	defparam lut_3572.LUT_SIZE = 5;
	defparam lut_3572.mask = 32'h77778000;

	lut_sub lut_3574 ({sk[1294], i_8_, x496x, x666x, x7084x, x7082x, x7083x}, x1608x);
	defparam lut_3574.LUT_SIZE = 7;
	defparam lut_3574.mask = 128'h57ffffff57ffffff0003050700030003;

	lut_sub lut_3577 ({sk[1295], i_28_, i_33_, i_29_, n_n1314, x76x, x269x}, x1609x);
	defparam lut_3577.LUT_SIZE = 7;
	defparam lut_3577.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_3579 ({sk[1296], i_13_, i_16_, x54x, x11x, n_n1305, x366x}, x1610x);
	defparam lut_3579.LUT_SIZE = 7;
	defparam lut_3579.mask = 128'h57ffffff57ffffff0001000000000000;

	lut_sub lut_3581 ({sk[1297], i_14_, i_12_, i_16_, i_37_, x376x, x273x}, x1611x);
	defparam lut_3581.LUT_SIZE = 7;
	defparam lut_3581.mask = 128'h57ffffff57ffffff0100000000000000;

	lut_sub lut_3583 ({sk[1298], i_7_, i_13_, i_16_, i_31_, i_34_}, x7038x);
	defparam lut_3583.LUT_SIZE = 6;
	defparam lut_3583.mask = 64'h3f3fffff00001000;

	lut_sub lut_3585 ({sk[1299], i_7_, i_14_, i_28_, i_37_}, x7014x);
	defparam lut_3585.LUT_SIZE = 5;
	defparam lut_3585.mask = 32'h77774000;

	lut_sub lut_3587 ({sk[1300], i_30_, i_32_, i_31_, i_34_, i_35_, i_29_}, x7015x);
	defparam lut_3587.LUT_SIZE = 7;
	defparam lut_3587.mask = 128'h57ffffff57ffffff2000000000000000;

	lut_sub lut_3589 ({sk[1301], i_30_, i_34_, i_35_, i_37_}, x7004x);
	defparam lut_3589.LUT_SIZE = 5;
	defparam lut_3589.mask = 32'h77770400;

	lut_sub lut_3591 ({sk[1302], i_7_, i_8_, i_14_, i_23_, i_17_, i_16_}, x7005x);
	defparam lut_3591.LUT_SIZE = 7;
	defparam lut_3591.mask = 128'h57ffffff57ffffff8000000000000000;

	lut_sub lut_3593 ({sk[1303], i_14_, i_12_, i_17_, i_16_, i_37_}, x7007x);
	defparam lut_3593.LUT_SIZE = 6;
	defparam lut_3593.mask = 64'h3f3fffff44400000;

	lut_sub lut_3596 ({sk[1304], i_30_, i_35_, i_29_, i_37_}, x6994x);
	defparam lut_3596.LUT_SIZE = 5;
	defparam lut_3596.mask = 32'h77774000;

	lut_sub lut_3598 ({sk[1305], i_27_, i_23_, i_16_, i_34_, i_35_}, x6995x);
	defparam lut_3598.LUT_SIZE = 6;
	defparam lut_3598.mask = 64'h3f3fffff40000000;

	lut_sub lut_3600 ({sk[1306], i_32_, i_34_, i_33_, i_35_, i_37_}, x6978x);
	defparam lut_3600.LUT_SIZE = 6;
	defparam lut_3600.mask = 64'h3f3fffff40000000;

	lut_sub lut_3602 ({sk[1307], i_7_, i_13_, i_12_, i_23_, i_24_, i_16_}, x6980x);
	defparam lut_3602.LUT_SIZE = 7;
	defparam lut_3602.mask = 128'h57ffffff57ffffff0000000080000000;

	lut_sub lut_3604 ({sk[1308], i_7_, i_14_, i_16_, i_31_, i_34_}, x6981x);
	defparam lut_3604.LUT_SIZE = 6;
	defparam lut_3604.mask = 64'h3f3fffff00001000;

	lut_sub lut_3606 ({sk[1309], i_7_, i_34_, i_35_, i_37_}, x6957x);
	defparam lut_3606.LUT_SIZE = 5;
	defparam lut_3606.mask = 32'h77771000;

	lut_sub lut_3608 ({sk[1310], i_14_, i_26_, i_24_, i_34_, i_35_, i_37_}, x6966x);
	defparam lut_3608.LUT_SIZE = 7;
	defparam lut_3608.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_3610 ({sk[1311], i_7_, i_34_, i_37_}, x6971x);
	defparam lut_3610.LUT_SIZE = 4;
	defparam lut_3610.mask = 16'h5510;

	lut_sub lut_3612 ({sk[1312], i_32_, i_31_, i_33_}, x6967x);
	defparam lut_3612.LUT_SIZE = 4;
	defparam lut_3612.mask = 16'h5580;

	lut_sub lut_3614 ({sk[1313], i_14_, i_28_, i_23_, i_24_, i_29_}, x6970x);
	defparam lut_3614.LUT_SIZE = 6;
	defparam lut_3614.mask = 64'h3f3fffff80000000;

	lut_sub lut_3616 ({sk[1314], i_7_, i_14_, i_12_, i_23_, i_24_, i_16_}, x6972x);
	defparam lut_3616.LUT_SIZE = 7;
	defparam lut_3616.mask = 128'h57ffffff57ffffff0000000080000000;

	lut_sub lut_3618 ({sk[1315], i_13_, i_2_, i_16_}, x6973x);
	defparam lut_3618.LUT_SIZE = 4;
	defparam lut_3618.mask = 16'h5520;

	lut_sub lut_3620 ({sk[1316], i_10_, i_14_, i_13_, i_16_, i_35_, i_37_}, x6935x);
	defparam lut_3620.LUT_SIZE = 7;
	defparam lut_3620.mask = 128'h57ffffff57ffffff4040000000400000;

	lut_sub lut_3623 ({sk[1317], i_27_, i_26_, i_24_, i_33_, i_35_, i_37_}, x6921x);
	defparam lut_3623.LUT_SIZE = 7;
	defparam lut_3623.mask = 128'h57ffffff57ffffff4000000000000000;

	lut_sub lut_3625 ({sk[1318], i_9_, i_14_, i_37_}, x6900x);
	defparam lut_3625.LUT_SIZE = 4;
	defparam lut_3625.mask = 16'h5540;

	lut_sub lut_3627 ({sk[1319], i_14_, i_11_, i_16_, i_37_}, x6908x);
	defparam lut_3627.LUT_SIZE = 5;
	defparam lut_3627.mask = 32'h77774000;

	lut_sub lut_3629 ({sk[1320], i_10_, i_13_, i_33_, i_37_}, x6879x);
	defparam lut_3629.LUT_SIZE = 5;
	defparam lut_3629.mask = 32'h77774000;

	lut_sub lut_3631 ({sk[1321], i_7_, i_31_, x10x, x74x, x372x, x7029x}, x7034x);
	defparam lut_3631.LUT_SIZE = 7;
	defparam lut_3631.mask = 128'h57ffffff57ffffff111111111111111f;

	lut_sub lut_3634 ({sk[1322], n_n1390, n_n1406, x8x, x7025x, x305x, x717x}, x7035x);
	defparam lut_3634.LUT_SIZE = 7;
	defparam lut_3634.mask = 128'h57ffffff57ffffff0000000f1111111f;

	lut_sub lut_3637 ({sk[1323], i_28_, i_25_, i_29_, x48x, x479x, x7038x}, x7039x);
	defparam lut_3637.LUT_SIZE = 7;
	defparam lut_3637.mask = 128'h57ffffff57ffffff0505370505050505;

	lut_sub lut_3640 ({sk[1324], n_n1429, x8x, x45x, x806x, x6950x, x7033x}, x7040x);
	defparam lut_3640.LUT_SIZE = 7;
	defparam lut_3640.mask = 128'h57ffffff57ffffff0303035703570357;

	lut_sub lut_3644 ({sk[1325], x323x, x246x, x29x, x445x, x7078x, x7080x}, x7089x);
	defparam lut_3644.LUT_SIZE = 7;
	defparam lut_3644.mask = 128'h57ffffff57ffffff0003000300035557;

	lut_sub lut_3647 ({sk[1326], i_35_, n_n1326, x275x, n_n1080, x694x, x693x}, x7110x);
	defparam lut_3647.LUT_SIZE = 7;
	defparam lut_3647.mask = 128'h57ffffff57ffffff0055005500550357;

	lut_sub lut_3650 ({sk[1327], i_9_, i_10_, i_35_, i_38_}, x7319x);
	defparam lut_3650.LUT_SIZE = 5;
	defparam lut_3650.mask = 32'h77770040;

	lut_sub lut_3652 ({sk[1328], i_10_, i_13_, i_26_, i_24_}, x7388x);
	defparam lut_3652.LUT_SIZE = 5;
	defparam lut_3652.mask = 32'h77778808;

	lut_sub lut_3655 ({sk[1329], i_31_, i_29_}, x7530x);
	defparam lut_3655.LUT_SIZE = 3;
	defparam lut_3655.mask = 8'h38;

	lut_sub lut_3657 ({sk[1330], i_8_, i_28_, i_29_}, x7532x);
	defparam lut_3657.LUT_SIZE = 4;
	defparam lut_3657.mask = 16'h5580;

	lut_sub lut_3659 ({sk[1331], i_12_, n_n1179, x376x, x71x, x7556x, x7560x}, x7565x);
	defparam lut_3659.LUT_SIZE = 7;
	defparam lut_3659.mask = 128'h57ffffff57ffffff0033053700000505;

	lut_sub lut_3662 ({sk[1332], i_38_, x11x, x321x, x52x, x446x, x7562x}, x7566x);
	defparam lut_3662.LUT_SIZE = 7;
	defparam lut_3662.mask = 128'h57ffffff57ffffff0000030300550357;

	lut_sub lut_3665 ({sk[1333], x49x, n_n1288, x51x, x12x, n_n1059, x7564x}, x7567x);
	defparam lut_3665.LUT_SIZE = 7;
	defparam lut_3665.mask = 128'h57ffffff57ffffff0005000500053337;

	lut_sub lut_3668 ({sk[1334], x1172x, x7565x, x7566x, x7567x}, x7570x);
	defparam lut_3668.LUT_SIZE = 5;
	defparam lut_3668.mask = 32'h77777fff;

	lut_sub lut_3673 ({sk[1335], x49x, x46x, x7491x, x7492x, x8x, x78x}, x7592x);
	defparam lut_3673.LUT_SIZE = 7;
	defparam lut_3673.mask = 128'h57ffffff57ffffff0000003305050537;

	lut_sub lut_3676 ({sk[1336], i_9_, i_12_, x782x, x1139x, x1141x, x7592x}, x7595x);
	defparam lut_3676.LUT_SIZE = 7;
	defparam lut_3676.mask = 128'h57ffffff57ffffff7f7f7f7f7f7f7fff;

	lut_sub lut_3681 ({sk[1337], x58x, n_n1368, x1078x, x1079x, x1076x, x1077x}, x7640x);
	defparam lut_3681.LUT_SIZE = 7;
	defparam lut_3681.mask = 128'h57ffffff57ffffff00000fff77777fff;

	lut_sub lut_3686 ({sk[1338], i_23_, x646x, x7635x, n_n1897, x7640x}, x7642x);
	defparam lut_3686.LUT_SIZE = 6;
	defparam lut_3686.mask = 64'h3f3fffff7f7f7fff;

	lut_sub lut_3691 ({sk[1339], i_30_, i_8_, i_2_}, x7670x);
	defparam lut_3691.LUT_SIZE = 4;
	defparam lut_3691.mask = 16'h5580;

	lut_sub lut_3693 ({sk[1340], i_14_, x42x, n_n1353, x57x, x479x, x509x}, x7675x);
	defparam lut_3693.LUT_SIZE = 7;
	defparam lut_3693.mask = 128'h57ffffff57ffffff0005000500053337;

	lut_sub lut_3696 ({sk[1341], n_n1375, n_n1374, n_n762, x1038x, x1039x, x7674x}, x7676x);
	defparam lut_3696.LUT_SIZE = 7;
	defparam lut_3696.mask = 128'h00ff00ffffffffff0055005500553f7f;

	lut_sub lut_3700 ({sk[1342], i_2_, i_32_, x61x, x226x, x466x, x7670x}, x7677x);
	defparam lut_3700.LUT_SIZE = 7;
	defparam lut_3700.mask = 128'h00ff00ffffffffff0307000500050005;

	lut_sub lut_3703 ({sk[1343], i_34_, x54x, n_n1489, x340x, x372x, x7029x}, x7933x);
	defparam lut_3703.LUT_SIZE = 7;
	defparam lut_3703.mask = 128'h00ff00ffffffffff111111111111111f;

	lut_sub lut_3706 ({sk[1344], i_32_, i_34_, i_36_, i_35_, x419x, x513x}, x7934x);
	defparam lut_3706.LUT_SIZE = 7;
	defparam lut_3706.mask = 128'h00ff00ffffffffff0050003000000000;

	lut_sub lut_3709 ({sk[1345], n_n1406, x8x, x1038x, x1039x, x7025x, x7932x}, x7935x);
	defparam lut_3709.LUT_SIZE = 7;
	defparam lut_3709.mask = 128'h00ff00ffffffffff0555055505553777;

	lut_sub lut_3713 ({sk[1346], i_27_, i_36_, x19x, x42x, n_n1202, x6x}, x8093x);
	defparam lut_3713.LUT_SIZE = 7;
	defparam lut_3713.mask = 128'h00ff00ffffffffff5555555755555555;

	lut_sub lut_3716 ({sk[1347], i_21_, x1765x, x1766x, x101x, x102x, x8085x}, x8094x);
	defparam lut_3716.LUT_SIZE = 7;
	defparam lut_3716.mask = 128'h77ff77ff77ff77ff3f7f7f7f00555555;


endmodule