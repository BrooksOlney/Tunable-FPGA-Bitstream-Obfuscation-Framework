module ks_misex3_qmap_map (sk, b, e, f, g, n, m, k, j, l, h, i, d, c, a, r2, s2, t2, u2, n2, o2, p2, q2, h2, i2, j2, k2, m2, l2);

	input b;
	input e;
	input f;
	input g;
	input n;
	input m;
	input k;
	input j;
	input l;
	input h;
	input i;
	input d;
	input c;
	input a;
	output r2;
	output s2;
	output t2;
	output u2;
	output n2;
	output o2;
	output p2;
	output q2;
	output h2;
	output i2;
	output j2;
	output k2;
	output m2;
	output l2;

	input [127 : 0] sk /* synthesis noprune */;


	wire g53, g103, g129, g173, g217, g235, g252, g274, g295, g328, g339, g345, g351, g1, g2, g3, g4, g5, g6, g7, g8;
	wire g9, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g20, g21, g22, g23, g24, g25, g26, g27, g28, g29;
	wire g30, g31, g32, g33, g34, g35, g36, g37, g38, g39, g40, g41, g42, g43, g44, g45, g46, g47, g48, g49, g50;
	wire g51, g455, g52, g54, g55, g56, g57, g58, g59, g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g70, g71;
	wire g72, g73, g74, g75, g76, g77, g78, g79, g80, g81, g82, g83, g84, g85, g86, g87, g88, g89, g90, g91, g92;
	wire g93, g94, g95, g96, g97, g98, g99, g100, g101, g539, g102, g104, g105, g106, g107, g108, g109, g110, g111, g112, g113;
	wire g114, g115, g116, g117, g118, g119, g120, g121, g122, g123, g124, g125, g126, g127, g128, g130, g131, g132, g532, g133, g134;
	wire g135, g136, g137, g138, g139, g140, g141, g142, g525, g143, g144, g145, g146, g147, g148, g149, g150, g151, g152, g153, g154;
	wire g155, g156, g157, g158, g159, g160, g161, g162, g163, g164, g165, g166, g167, g168, g169, g511, g170, g171, g172, g518, g174;
	wire g175, g176, g504, g177, g178, g179, g180, g181, g182, g183, g184, g185, g186, g187, g188, g189, g190, g191, g192, g193, g194;
	wire g195, g196, g197, g198, g199, g200, g201, g202, g203, g204, g205, g206, g207, g208, g497, g209, g210, g211, g212, g213, g214;
	wire g215, g216, g218, g219, g220, g221, g222, g223, g224, g225, g226, g227, g228, g229, g230, g231, g232, g233, g234, g236, g237;
	wire g238, g239, g240, g241, g242, g243, g244, g245, g246, g247, g248, g249, g250, g251, g253, g254, g255, g256, g257, g258, g259;
	wire g260, g261, g262, g263, g264, g265, g266, g267, g268, g269, g270, g271, g479, g272, g273, g486, g275, g276, g277, g278, g279;
	wire g280, g281, g282, g283, g284, g285, g286, g287, g472, g288, g289, g290, g291, g292, g293, g294, g296, g297, g298, g299, g300;
	wire g301, g302, g303, g304, g305, g306, g307, g308, g309, g310, g311, g312, g313, g314, g315, g316, g317, g318, g319, g320, g321;
	wire g322, g323, g324, g325, g326, g327, g329, g330, g331, g332, g333, g334, g335, g336, g337, g338, g340, g341, g342, g343, g344;
	wire g346, g347, g348, g349, g350, g352, g353, g354, g355, g356, g357, g358, g359, g360, g361, g362, g363, g364, g365, g366, g367;
	wire g368, g369, g370, g371, g372, g373, g374, g375, g376, g377, g378, g379, g380, g381, g462, g382, g383, g384, g385, g386, g387;
	wire g388, g389, g390, g391, g392, g393, g394, g395, g396, g397, g398, g399, g400, g401, g402, g403, g404, g405, g406, g407, g408;
	wire g409, g410, g411, g412, g413, g414, g415, g416, g417, g418, g419, g420, g421, g422, g423, g424, g425, g426, g427, g428, g429;
	wire g430, g431, g432, g433, g434, g435, g436, g437, g438, g439, g440, g441, g442, g443, g444, g445, g446, g456, g447, g448, g449;
	wire g450, g451, g453, g454, g457, g458, g459, g460, g461, g463, g464, g465, g468, g466, g467, g469, g470, g471, g473, g474, g475;
	wire g476, g477, g478, g480, g481, g482, g483, g484, g485, g487, g488, g489, g492, g490, g491, g494, g495, g493, g496, g498, g499;
	wire g500, g501, g502, g503, g505, g506, g507, g508, g509, g510, g512, g513, g514, g515, g516, g517, g519, g520, g521, g522, g523;
	wire g524, g526, g527, g528, g529, g530, g531, g533, g534, g535, g536, g537, g538, g540, g541, g542, g545, g543, g544, g547, g548;
	wire g546, g549;

	assign r2 = (((sk[0]) & (!g53)));
	assign s2 = (((sk[1]) & (!g103)));
	assign t2 = (((sk[2]) & (!g129)));
	assign u2 = (((sk[3]) & (!g173)));
	assign n2 = (((sk[4]) & (!g217)));
	assign o2 = (((sk[5]) & (!g235)));
	assign p2 = (((sk[6]) & (!g252)));
	assign q2 = (((sk[7]) & (!g274)));
	assign h2 = (((sk[8]) & (!g295)));
	assign i2 = (((sk[9]) & (!g328)));
	assign j2 = (((sk[10]) & (!g339)));
	assign k2 = (((sk[11]) & (!g345)));
	assign m2 = (((sk[12]) & (!g351)));
	assign g1 = (((!n) & (!sk[13]) & (m)) + ((n) & (sk[13]) & (!m)));
	assign g2 = (((!sk[14]) & (!n) & (!m) & (j) & (!l)) + ((!sk[14]) & (!n) & (!m) & (!j) & (l)) + ((!sk[14]) & (n) & (!m) & (!j) & (l)));
	assign g3 = (((!sk[15]) & (!k) & (g1) & (!g2)) + ((sk[15]) & (!k) & (!g1) & (!g2)) + ((!sk[15]) & (!k) & (g1) & (!g2)));
	assign g4 = (((k) & (!sk[16]) & (g1)) + ((!k) & (!sk[16]) & (g1)));
	assign g5 = (((h) & (!g) & (!j) & (!i) & (!sk[17]) & (!g4)) + ((!h) & (!g) & (j) & (!i) & (!sk[17]) & (!g4)) + ((!h) & (!g) & (!j) & (!i) & (!sk[17]) & (g4)) + ((!h) & (!g) & (!j) & (i) & (sk[17]) & (!g4)) + ((h) & (!g) & (!j) & (!i) & (!sk[17]) & (g4)) + ((!h) & (!g) & (!j) & (i) & (!sk[17]) & (g4)));
	assign g6 = (((!h) & (!j) & (!sk[18]) & (k) & (!l)) + ((!h) & (!j) & (!sk[18]) & (!k) & (l)) + ((h) & (!j) & (!sk[18]) & (k) & (!l)) + ((h) & (j) & (sk[18]) & (!k) & (!l)));
	assign g7 = (((!sk[19]) & (g) & (!g1) & (!g3) & (!g5) & (!g6)) + ((!sk[19]) & (!g) & (!g1) & (g3) & (!g5) & (!g6)) + ((!sk[19]) & (!g) & (!g1) & (!g3) & (!g5) & (g6)) + ((sk[19]) & (!g) & (!g1) & (!g3) & (g5) & (!g6)) + ((!sk[19]) & (!g) & (g1) & (!g3) & (!g5) & (g6)));
	assign g8 = (((!e) & (f) & (!sk[20]) & (!g7)) + ((!e) & (f) & (!sk[20]) & (g7)));
	assign g9 = (((!sk[21]) & (!n) & (m)) + ((sk[21]) & (!n) & (!m)));
	assign g10 = (((!h) & (!sk[22]) & (i)) + ((!h) & (!sk[22]) & (i)));
	assign g11 = (((!sk[23]) & (h) & (!j) & (!k) & (!i) & (!l)) + ((!sk[23]) & (!h) & (!j) & (k) & (!i) & (!l)) + ((!sk[23]) & (!h) & (!j) & (!k) & (!i) & (l)) + ((!sk[23]) & (h) & (j) & (!k) & (!i) & (!l)) + ((!sk[23]) & (!h) & (!j) & (k) & (i) & (!l)) + ((!sk[23]) & (h) & (!j) & (k) & (!i) & (!l)) + ((!sk[23]) & (h) & (!j) & (k) & (!i) & (!l)) + ((!sk[23]) & (!h) & (!j) & (k) & (i) & (!l)));
	assign g12 = (((j) & (!sk[24]) & (!l) & (!g9) & (!g10) & (!g11)) + ((!j) & (!sk[24]) & (!l) & (g9) & (!g10) & (!g11)) + ((!j) & (!sk[24]) & (!l) & (!g9) & (!g10) & (g11)) + ((!j) & (!sk[24]) & (!l) & (g9) & (!g10) & (g11)) + ((!j) & (!sk[24]) & (l) & (g9) & (g10) & (!g11)));
	assign g13 = (((!sk[25]) & (d) & (!e) & (!f) & (!g12) & (!c)) + ((!sk[25]) & (!d) & (!e) & (f) & (!g12) & (!c)) + ((!sk[25]) & (!d) & (!e) & (!f) & (!g12) & (c)) + ((!sk[25]) & (!d) & (!e) & (f) & (g12) & (c)) + ((!sk[25]) & (!d) & (!e) & (f) & (g12) & (c)));
	assign g14 = (((h) & (!sk[26]) & (!j) & (k) & (!l)) + ((!h) & (!sk[26]) & (!j) & (k) & (!l)) + ((!h) & (!sk[26]) & (!j) & (!k) & (l)) + ((h) & (!sk[26]) & (!j) & (!k) & (l)));
	assign g15 = (((!sk[27]) & (!n) & (m)) + ((!sk[27]) & (!n) & (m)));
	assign g16 = (((!sk[28]) & (!b) & (d) & (!a)) + ((!sk[28]) & (b) & (d) & (a)));
	assign g17 = (((!sk[29]) & (h) & (!j) & (!k) & (!i) & (!l)) + ((!sk[29]) & (!h) & (!j) & (k) & (!i) & (!l)) + ((!sk[29]) & (!h) & (!j) & (!k) & (!i) & (l)) + ((!sk[29]) & (h) & (!j) & (k) & (i) & (l)) + ((!sk[29]) & (!h) & (!j) & (!k) & (!i) & (l)) + ((sk[29]) & (!h) & (!j) & (!k) & (!i) & (!l)) + ((!sk[29]) & (h) & (!j) & (!k) & (i) & (!l)) + ((!sk[29]) & (h) & (!j) & (!k) & (!i) & (!l)) + ((!sk[29]) & (!h) & (j) & (k) & (!i) & (!l)));
	assign g18 = (((!j) & (!k) & (!sk[30]) & (i) & (!g17)) + ((!j) & (!k) & (!sk[30]) & (!i) & (g17)) + ((j) & (k) & (!sk[30]) & (!i) & (g17)) + ((!j) & (!k) & (!sk[30]) & (i) & (g17)) + ((!j) & (!k) & (!sk[30]) & (!i) & (g17)));
	assign g19 = (((!e) & (!g) & (g14) & (g15) & (g16) & (!g18)) + ((!e) & (g) & (!g14) & (g15) & (g16) & (!g18)));
	assign g20 = (((!d) & (!sk[32]) & (e) & (!c)) + ((d) & (!sk[32]) & (e) & (c)));
	assign g21 = (((n) & (!m) & (!j) & (!k) & (!sk[33]) & (!l)) + ((!n) & (!m) & (j) & (!k) & (!sk[33]) & (!l)) + ((!n) & (!m) & (!j) & (!k) & (!sk[33]) & (l)) + ((!n) & (!m) & (!j) & (k) & (sk[33]) & (!l)) + ((!n) & (!m) & (!j) & (!k) & (!sk[33]) & (l)));
	assign g22 = (((!f) & (g10) & (!sk[34]) & (!g21)) + ((!f) & (g10) & (!sk[34]) & (g21)));
	assign g23 = (((!sk[35]) & (!f) & (h)) + ((!sk[35]) & (!f) & (h)));
	assign g24 = (((!j) & (k) & (!i) & (!l) & (g9) & (g23)) + ((j) & (!k) & (!i) & (!l) & (g9) & (g23)) + ((!j) & (k) & (!i) & (!l) & (g9) & (g23)) + ((!j) & (k) & (!i) & (!l) & (g9) & (g23)));
	assign g25 = (((!b) & (!sk[37]) & (!h) & (i) & (!g1)) + ((!b) & (!sk[37]) & (!h) & (!i) & (g1)) + ((b) & (!sk[37]) & (h) & (!i) & (g1)) + ((b) & (!sk[37]) & (!h) & (i) & (g1)));
	assign g26 = (((h) & (!j) & (!k) & (!i) & (!sk[38]) & (!l)) + ((!h) & (!j) & (k) & (!i) & (!sk[38]) & (!l)) + ((!h) & (!j) & (!k) & (!i) & (!sk[38]) & (l)) + ((h) & (!j) & (!k) & (!i) & (!sk[38]) & (!l)) + ((h) & (j) & (k) & (i) & (!sk[38]) & (l)) + ((!h) & (j) & (!k) & (!i) & (sk[38]) & (!l)) + ((!h) & (!j) & (!k) & (!i) & (sk[38]) & (!l)));
	assign g27 = (((e) & (!f) & (!c) & (!g25) & (!sk[39]) & (!g26)) + ((!e) & (!f) & (c) & (!g25) & (!sk[39]) & (!g26)) + ((!e) & (!f) & (!c) & (!g25) & (!sk[39]) & (g26)) + ((e) & (!f) & (c) & (g25) & (!sk[39]) & (!g26)));
	assign g28 = (((!sk[40]) & (g19) & (!g20) & (!g22) & (!g24) & (!g27)) + ((!sk[40]) & (!g19) & (!g20) & (g22) & (!g24) & (!g27)) + ((!sk[40]) & (!g19) & (!g20) & (!g22) & (!g24) & (g27)) + ((sk[40]) & (!g19) & (!g20) & (!g22) & (!g24) & (!g27)) + ((sk[40]) & (!g19) & (!g20) & (!g22) & (!g24) & (!g27)));
	assign g29 = (((!j) & (k) & (!sk[41]) & (!i)) + ((!j) & (k) & (!sk[41]) & (i)) + ((j) & (!k) & (sk[41]) & (!i)));
	assign g30 = (((b) & (!d) & (!e) & (!sk[42]) & (!c) & (!a)) + ((!b) & (!d) & (e) & (!sk[42]) & (!c) & (!a)) + ((!b) & (!d) & (!e) & (!sk[42]) & (!c) & (a)) + ((b) & (!d) & (e) & (!sk[42]) & (!c) & (!a)) + ((b) & (!d) & (e) & (!sk[42]) & (!c) & (!a)));
	assign g31 = (((n) & (!m) & (!j) & (k) & (!i) & (!l)) + ((n) & (!m) & (j) & (!k) & (!i) & (!l)) + ((n) & (!m) & (!j) & (k) & (!i) & (!l)) + ((n) & (!m) & (!j) & (k) & (!i) & (!l)));
	assign g32 = (((n) & (!m) & (!j) & (k) & (i) & (!l)) + ((n) & (!m) & (!j) & (!k) & (i) & (l)));
	assign g33 = (((!h) & (!sk[45]) & (g31) & (!g32)) + ((h) & (sk[45]) & (!g31) & (!g32)) + ((!h) & (sk[45]) & (!g31) & (!g32)));
	assign g34 = (((!e) & (!sk[46]) & (g)) + ((!e) & (!sk[46]) & (g)));
	assign g35 = (((b) & (!sk[47]) & (c)) + ((!b) & (!sk[47]) & (c)));
	assign g36 = (((!sk[48]) & (!d) & (g35)) + ((!sk[48]) & (!d) & (g35)));
	assign g37 = (((!b) & (!sk[49]) & (d) & (!c)) + ((b) & (!sk[49]) & (d) & (!c)));
	assign g38 = (((f) & (!g33) & (!sk[50]) & (!g34) & (!g36) & (!g37)) + ((!f) & (!g33) & (!sk[50]) & (g34) & (!g36) & (!g37)) + ((!f) & (!g33) & (!sk[50]) & (!g34) & (!g36) & (g37)) + ((!f) & (!g33) & (!sk[50]) & (g34) & (g36) & (!g37)) + ((f) & (!g33) & (!sk[50]) & (!g34) & (!g36) & (g37)));
	assign g39 = (((!sk[51]) & (!b) & (d) & (!e)) + ((sk[51]) & (!b) & (!d) & (!e)) + ((sk[51]) & (!b) & (!d) & (!e)));
	assign g40 = (((!f) & (!sk[52]) & (h) & (!g)) + ((f) & (!sk[52]) & (h) & (g)));
	assign g41 = (((!f) & (h) & (!sk[53]) & (!g)) + ((f) & (!h) & (sk[53]) & (g)));
	assign g42 = (((!g40) & (!g31) & (!sk[54]) & (g41) & (!g32)) + ((!g40) & (!g31) & (!sk[54]) & (!g41) & (g32)) + ((!g40) & (!g31) & (!sk[54]) & (g41) & (g32)) + ((g40) & (g31) & (sk[54]) & (!g41) & (!g32)));
	assign g43 = (((!b) & (d) & (!sk[55]) & (!e)) + ((b) & (d) & (!sk[55]) & (!e)));
	assign g44 = (((f) & (!sk[56]) & (h)) + ((!f) & (!sk[56]) & (h)));
	assign g45 = (((g44) & (!j) & (k) & (!i) & (!l) & (g1)) + ((g44) & (j) & (!k) & (!i) & (!l) & (g1)) + ((g44) & (!j) & (k) & (!i) & (!l) & (g1)) + ((g44) & (!j) & (k) & (!i) & (!l) & (g1)));
	assign g46 = (((!f) & (!g10) & (!g4) & (!g2) & (g43) & (g45)) + ((f) & (g10) & (g4) & (!g2) & (g43) & (!g45)) + ((f) & (g10) & (!g4) & (g2) & (g43) & (!g45)));
	assign g47 = (((!sk[59]) & (!g14) & (g15)) + ((!sk[59]) & (g14) & (g15)));
	assign g48 = (((!sk[60]) & (!g15) & (g29) & (!g17)) + ((!sk[60]) & (g15) & (g29) & (!g17)) + ((sk[60]) & (g15) & (!g29) & (!g17)));
	assign g49 = (((!d) & (a) & (!sk[61]) & (!g35)) + ((!d) & (a) & (!sk[61]) & (g35)));
	assign g50 = (((e) & (!g) & (!g47) & (!g48) & (!sk[62]) & (!g49)) + ((!e) & (!g) & (g47) & (!g48) & (!sk[62]) & (!g49)) + ((!e) & (!g) & (!g47) & (!g48) & (!sk[62]) & (g49)) + ((e) & (!g) & (g47) & (!g48) & (!sk[62]) & (g49)) + ((e) & (g) & (!g47) & (g48) & (!sk[62]) & (g49)));
	assign g51 = (((!sk[63]) & (!g39) & (!g42) & (g46) & (!g50)) + ((!sk[63]) & (!g39) & (!g42) & (!g46) & (g50)) + ((sk[63]) & (g39) & (!g42) & (!g46) & (!g50)) + ((sk[63]) & (!g39) & (!g42) & (!g46) & (!g50)));
	assign g52 = (((!g455) & (!g30) & (g38) & (!sk[64]) & (!g51)) + ((!g455) & (!g30) & (!g38) & (!sk[64]) & (g51)) + ((g455) & (!g30) & (!g38) & (!sk[64]) & (g51)) + ((!g455) & (!g30) & (!g38) & (!sk[64]) & (g51)));
	assign g53 = (((!sk[65]) & (b) & (!g8) & (!g13) & (!g28) & (!g52)) + ((!sk[65]) & (!b) & (!g8) & (g13) & (!g28) & (!g52)) + ((!sk[65]) & (!b) & (!g8) & (!g13) & (!g28) & (g52)) + ((!sk[65]) & (!b) & (!g8) & (!g13) & (g28) & (g52)) + ((!sk[65]) & (!b) & (!g8) & (!g13) & (g28) & (g52)));
	assign g54 = (((!n) & (!sk[66]) & (m) & (!k)) + ((!n) & (!sk[66]) & (m) & (k)));
	assign g55 = (((!h) & (!sk[67]) & (g) & (!g54)) + ((h) & (sk[67]) & (!g) & (g54)));
	assign g56 = (((!e) & (!sk[68]) & (g55)) + ((!e) & (!sk[68]) & (g55)));
	assign g57 = (((f) & (!sk[69]) & (g)) + ((!f) & (!sk[69]) & (g)));
	assign g58 = (((!j) & (!sk[70]) & (i)) + ((j) & (sk[70]) & (!i)));
	assign g59 = (((!m) & (!k) & (!sk[71]) & (l) & (!g58)) + ((!m) & (!k) & (!sk[71]) & (!l) & (g58)) + ((m) & (k) & (sk[71]) & (!l) & (!g58)));
	assign g60 = (((m) & (!j) & (!sk[72]) & (!k) & (!i) & (!l)) + ((!m) & (!j) & (!sk[72]) & (k) & (!i) & (!l)) + ((!m) & (!j) & (!sk[72]) & (!k) & (!i) & (l)) + ((m) & (j) & (!sk[72]) & (!k) & (!i) & (!l)) + ((m) & (j) & (!sk[72]) & (!k) & (!i) & (l)));
	assign g61 = (((!m) & (!sk[73]) & (k) & (!l)) + ((m) & (sk[73]) & (!k) & (l)));
	assign g62 = (((m) & (!sk[74]) & (l)) + ((!m) & (!sk[74]) & (l)));
	assign g63 = (((h) & (!j) & (!k) & (!i) & (!sk[75]) & (!g62)) + ((!h) & (!j) & (k) & (!i) & (!sk[75]) & (!g62)) + ((!h) & (!j) & (!k) & (!i) & (!sk[75]) & (g62)) + ((!h) & (j) & (!k) & (!i) & (!sk[75]) & (g62)) + ((!h) & (!j) & (!k) & (i) & (!sk[75]) & (g62)) + ((!h) & (j) & (!k) & (i) & (!sk[75]) & (g62)));
	assign g64 = (((!m) & (!sk[76]) & (j) & (!l)) + ((m) & (sk[76]) & (!j) & (l)));
	assign g65 = (((!sk[77]) & (!m) & (!j) & (i) & (!l)) + ((!sk[77]) & (!m) & (!j) & (!i) & (l)) + ((!sk[77]) & (m) & (!j) & (!i) & (l)) + ((sk[77]) & (m) & (j) & (!i) & (!l)));
	assign g66 = (((g44) & (!g) & (!g54) & (!sk[78]) & (!g64) & (!g65)) + ((!g44) & (!g) & (g54) & (!sk[78]) & (!g64) & (!g65)) + ((!g44) & (!g) & (!g54) & (!sk[78]) & (!g64) & (g65)) + ((g44) & (!g) & (g54) & (!sk[78]) & (!g64) & (!g65)) + ((g44) & (!g) & (!g54) & (!sk[78]) & (g64) & (!g65)) + ((g44) & (g) & (!g54) & (!sk[78]) & (!g64) & (g65)));
	assign g67 = (((!h) & (!g57) & (g61) & (!sk[79]) & (!g63) & (!g66)) + ((!h) & (!g57) & (!g61) & (!sk[79]) & (!g63) & (g66)) + ((h) & (!g57) & (!g61) & (!sk[79]) & (!g63) & (!g66)) + ((!h) & (!g57) & (!g61) & (sk[79]) & (!g63) & (!g66)) + ((!h) & (!g57) & (!g61) & (sk[79]) & (!g63) & (!g66)));
	assign g68 = (((n) & (!g57) & (!sk[80]) & (!g59) & (!g60) & (!g67)) + ((!n) & (!g57) & (!sk[80]) & (!g59) & (!g60) & (g67)) + ((!n) & (g57) & (!sk[80]) & (g59) & (!g60) & (!g67)) + ((!n) & (!g57) & (sk[80]) & (!g59) & (!g60) & (!g67)) + ((!n) & (!g57) & (!sk[80]) & (g59) & (!g60) & (!g67)) + ((!n) & (g57) & (!sk[80]) & (!g59) & (g60) & (g67)));
	assign g69 = (((!sk[81]) & (!j) & (g61)) + ((!sk[81]) & (j) & (g61)));
	assign g70 = (((h) & (!g34) & (!sk[82]) & (!g65) & (!g60) & (!g69)) + ((!h) & (!g34) & (!sk[82]) & (g65) & (!g60) & (!g69)) + ((!h) & (g34) & (!sk[82]) & (!g65) & (!g60) & (g69)) + ((!h) & (!g34) & (!sk[82]) & (!g65) & (!g60) & (g69)) + ((h) & (g34) & (!sk[82]) & (g65) & (!g60) & (!g69)) + ((!h) & (g34) & (sk[82]) & (!g65) & (g60) & (!g69)));
	assign g71 = (((!n) & (!m) & (k) & (!sk[83]) & (!l)) + ((!n) & (!m) & (!k) & (!sk[83]) & (l)) + ((!n) & (m) & (k) & (!sk[83]) & (!l)));
	assign g72 = (((!e) & (h) & (!g) & (!j) & (!i) & (g62)) + ((!e) & (!h) & (g) & (!j) & (i) & (g62)));
	assign g73 = (((!n) & (!g58) & (!g34) & (g70) & (!g71) & (!g72)) + ((!n) & (!g58) & (!g34) & (!g70) & (!g71) & (g72)) + ((!n) & (!g58) & (g34) & (!g70) & (g71) & (!g72)));
	assign g74 = (((!f) & (!g12) & (!a) & (!g56) & (!g68) & (!g73)) + ((!f) & (!g12) & (!a) & (!g56) & (!g68) & (!g73)) + ((!f) & (!g12) & (!a) & (!g56) & (!g68) & (!g73)) + ((!f) & (!g12) & (!a) & (!g56) & (!g68) & (!g73)));
	assign g75 = (((!e) & (h) & (!sk[87]) & (!g)) + ((e) & (h) & (!sk[87]) & (!g)));
	assign g76 = (((e) & (!sk[88]) & (g)) + ((!e) & (!sk[88]) & (g)));
	assign g77 = (((!m) & (j) & (!sk[89]) & (!k)) + ((m) & (!j) & (sk[89]) & (k)));
	assign g78 = (((!sk[90]) & (h) & (!i) & (!g76) & (!g62) & (!g77)) + ((!sk[90]) & (!h) & (!i) & (g76) & (!g62) & (!g77)) + ((!sk[90]) & (!h) & (!i) & (!g76) & (!g62) & (g77)) + ((!sk[90]) & (!h) & (i) & (g76) & (!g62) & (g77)) + ((!sk[90]) & (!h) & (i) & (g76) & (g62) & (!g77)));
	assign g79 = (((!h) & (g76) & (g59) & (!g65) & (!g60) & (!g69)) + ((!h) & (g76) & (!g59) & (!g65) & (g60) & (!g69)) + ((!h) & (g76) & (!g59) & (!g65) & (!g60) & (g69)) + ((h) & (g76) & (!g59) & (g65) & (!g60) & (!g69)));
	assign g80 = (((!n) & (!g54) & (!g75) & (!g64) & (g78) & (!g79)) + ((!n) & (!g54) & (!g75) & (!g64) & (!g78) & (g79)) + ((!n) & (g54) & (g75) & (!g64) & (!g78) & (!g79)) + ((!n) & (!g54) & (g75) & (g64) & (!g78) & (!g79)));
	assign g81 = (((!b) & (!c) & (sk[93]) & (!a)) + ((!b) & (c) & (!sk[93]) & (!a)) + ((b) & (!c) & (sk[93]) & (!a)) + ((!b) & (!c) & (sk[93]) & (!a)));
	assign g82 = (((!d) & (!sk[94]) & (e) & (!f)) + ((d) & (!sk[94]) & (e) & (f)));
	assign g83 = (((!g81) & (!sk[95]) & (g82) & (!g455)) + ((!g81) & (!sk[95]) & (g82) & (!g455)));
	assign g84 = (((!b) & (d) & (!sk[96]) & (!a)) + ((b) & (d) & (!sk[96]) & (!a)));
	assign g85 = (((e) & (!f) & (!sk[97]) & (!g) & (!g47) & (!g48)) + ((!e) & (!f) & (!sk[97]) & (g) & (!g47) & (!g48)) + ((!e) & (!f) & (!sk[97]) & (!g) & (!g47) & (g48)) + ((!e) & (f) & (!sk[97]) & (g) & (!g47) & (g48)) + ((!e) & (f) & (sk[97]) & (!g) & (g47) & (!g48)));
	assign g86 = (((!sk[98]) & (!j) & (i)) + ((!sk[98]) & (!j) & (i)));
	assign g87 = (((!n) & (!m) & (!sk[99]) & (k) & (!g86)) + ((!n) & (!m) & (!sk[99]) & (!k) & (g86)) + ((!n) & (m) & (!sk[99]) & (k) & (g86)));
	assign g88 = (((!sk[100]) & (!d) & (c) & (!a)) + ((sk[100]) & (!d) & (!c) & (!a)) + ((sk[100]) & (!d) & (!c) & (!a)));
	assign g89 = (((!g57) & (!sk[101]) & (!g34) & (g87) & (!g88)) + ((!g57) & (!sk[101]) & (!g34) & (!g87) & (g88)) + ((g57) & (!sk[101]) & (!g34) & (g87) & (!g88)) + ((!g57) & (!sk[101]) & (g34) & (g87) & (!g88)));
	assign g90 = (((!b) & (d) & (!sk[102]) & (!c)) + ((b) & (d) & (!sk[102]) & (c)));
	assign g91 = (((!e) & (!g44) & (g31) & (!sk[103]) & (!g90)) + ((!e) & (!g44) & (!g31) & (!sk[103]) & (g90)) + ((!e) & (g44) & (g31) & (!sk[103]) & (g90)));
	assign g92 = (((!sk[104]) & (e) & (!f) & (!h) & (!g32) & (!g90)) + ((!sk[104]) & (!e) & (!f) & (h) & (!g32) & (!g90)) + ((!sk[104]) & (!e) & (!f) & (!h) & (!g32) & (g90)) + ((!sk[104]) & (!e) & (f) & (!h) & (g32) & (g90)));
	assign g93 = (((!b) & (!sk[105]) & (f) & (!c)) + ((!b) & (!sk[105]) & (f) & (c)));
	assign g94 = (((j) & (!sk[106]) & (!l) & (!g1) & (!g10) & (!g11)) + ((!j) & (!sk[106]) & (!l) & (g1) & (!g10) & (!g11)) + ((!j) & (!sk[106]) & (!l) & (!g1) & (!g10) & (g11)) + ((!j) & (!sk[106]) & (!l) & (g1) & (!g10) & (g11)) + ((!j) & (!sk[106]) & (l) & (g1) & (g10) & (!g11)));
	assign g95 = (((f) & (!g34) & (!g36) & (!g93) & (!sk[107]) & (!g94)) + ((!f) & (!g34) & (g36) & (!g93) & (!sk[107]) & (!g94)) + ((!f) & (!g34) & (!g36) & (g93) & (!sk[107]) & (g94)) + ((!f) & (!g34) & (!g36) & (!g93) & (!sk[107]) & (g94)) + ((f) & (g34) & (g36) & (!g93) & (!sk[107]) & (g94)));
	assign g96 = (((g81) & (!g85) & (!g89) & (!g91) & (!g92) & (!g95)) + ((!g81) & (!g85) & (!g89) & (!g91) & (!g92) & (!g95)));
	assign g97 = (((d) & (!sk[109]) & (c)) + ((!d) & (!sk[109]) & (c)));
	assign g98 = (((!sk[110]) & (!g9) & (g6)) + ((!sk[110]) & (g9) & (g6)));
	assign g99 = (((!sk[111]) & (!j) & (i)) + ((!sk[111]) & (j) & (i)));
	assign g100 = (((!sk[112]) & (!g44) & (!k) & (g9) & (!g99)) + ((!sk[112]) & (!g44) & (!k) & (!g9) & (g99)) + ((!sk[112]) & (g44) & (k) & (g9) & (!g99)));
	assign g101 = (((f) & (!g10) & (!g21) & (!g98) & (!sk[113]) & (!g100)) + ((!f) & (!g10) & (!g21) & (!g98) & (!sk[113]) & (g100)) + ((!f) & (!g10) & (!g21) & (!g98) & (sk[113]) & (!g100)) + ((!f) & (!g10) & (g21) & (!g98) & (!sk[113]) & (!g100)) + ((!f) & (!g10) & (!g21) & (!g98) & (sk[113]) & (!g100)) + ((!f) & (!g10) & (!g21) & (!g98) & (sk[113]) & (!g100)));
	assign g102 = (((!g80) & (!g83) & (g28) & (!g84) & (g96) & (g539)) + ((!g80) & (!g83) & (g28) & (!g84) & (g96) & (g539)));
	assign g103 = (((d) & (!c) & (!sk[115]) & (!g8) & (!g74) & (!g102)) + ((!d) & (!c) & (!sk[115]) & (g8) & (!g74) & (!g102)) + ((!d) & (!c) & (!sk[115]) & (!g8) & (!g74) & (g102)) + ((!d) & (c) & (!sk[115]) & (!g8) & (!g74) & (g102)) + ((!d) & (!c) & (!sk[115]) & (!g8) & (g74) & (g102)));
	assign g104 = (((!f) & (!g10) & (!sk[116]) & (!g3) & (g45)) + ((!f) & (!g10) & (!sk[116]) & (g3) & (!g45)) + ((!f) & (!g10) & (sk[116]) & (!g3) & (!g45)) + ((!f) & (!g10) & (sk[116]) & (!g3) & (!g45)));
	assign g105 = (((f) & (!h) & (!sk[117]) & (!g) & (!g31) & (!g32)) + ((!f) & (!h) & (!sk[117]) & (g) & (!g31) & (!g32)) + ((!f) & (!h) & (!sk[117]) & (!g) & (!g31) & (g32)) + ((!f) & (h) & (!sk[117]) & (g) & (g31) & (!g32)) + ((!f) & (!h) & (!sk[117]) & (g) & (!g31) & (g32)));
	assign g106 = (((e) & (!f) & (!g37) & (!sk[118]) & (!g94) & (!g105)) + ((!e) & (!f) & (g37) & (!sk[118]) & (!g94) & (!g105)) + ((!e) & (!f) & (g37) & (!sk[118]) & (!g94) & (g105)) + ((!e) & (!f) & (!g37) & (!sk[118]) & (!g94) & (g105)) + ((e) & (f) & (g37) & (!sk[118]) & (g94) & (!g105)));
	assign g107 = (((!sk[119]) & (!b) & (e) & (!c)) + ((!sk[119]) & (!b) & (e) & (c)));
	assign g108 = (((!sk[120]) & (!e) & (!f) & (g12) & (!c)) + ((!sk[120]) & (!e) & (!f) & (!g12) & (c)) + ((!sk[120]) & (e) & (!f) & (g12) & (c)));
	assign g109 = (((!sk[121]) & (!g57) & (g87)) + ((!sk[121]) & (g57) & (g87)));
	assign g110 = (((b) & (!d) & (!e) & (!a) & (!sk[122]) & (!g109)) + ((!b) & (!d) & (e) & (!a) & (!sk[122]) & (!g109)) + ((!b) & (!d) & (!e) & (!a) & (!sk[122]) & (g109)) + ((!b) & (d) & (!e) & (a) & (!sk[122]) & (g109)) + ((b) & (!d) & (!e) & (!a) & (!sk[122]) & (g109)));
	assign g111 = (((!b) & (!sk[123]) & (!d) & (f) & (!a)) + ((!b) & (!sk[123]) & (!d) & (!f) & (a)) + ((!b) & (!sk[123]) & (d) & (f) & (a)));
	assign g112 = (((!sk[124]) & (f) & (!g) & (!g47) & (!g48) & (!g111)) + ((!sk[124]) & (!f) & (!g) & (g47) & (!g48) & (!g111)) + ((!sk[124]) & (!f) & (!g) & (!g47) & (!g48) & (g111)) + ((!sk[124]) & (!f) & (!g) & (g47) & (!g48) & (g111)) + ((!sk[124]) & (!f) & (!g) & (g47) & (g48) & (g111)) + ((!sk[124]) & (f) & (g) & (!g47) & (g48) & (g111)));
	assign g113 = (((!sk[125]) & (!b) & (c) & (!a)) + ((sk[125]) & (b) & (!c) & (a)));
	assign g114 = (((!sk[126]) & (!d) & (c) & (!a)) + ((!sk[126]) & (!d) & (c) & (a)));
	assign g115 = (((g) & (!sk[127]) & (!g14) & (!g15) & (!g29) & (!g17)) + ((!g) & (!sk[127]) & (!g14) & (g15) & (!g29) & (!g17)) + ((!g) & (!sk[127]) & (!g14) & (!g15) & (!g29) & (g17)) + ((!g) & (!sk[127]) & (g14) & (g15) & (!g29) & (!g17)) + ((g) & (!sk[127]) & (!g14) & (g15) & (g29) & (!g17)) + ((g) & (!sk[127]) & (!g14) & (g15) & (!g29) & (!g17)));
	assign g116 = (((!d) & (!e) & (f) & (g113) & (!g114) & (g115)) + ((!d) & (e) & (f) & (!g113) & (g114) & (g115)));
	assign g117 = (((g108) & (!sk[1]) & (!g110) & (!g27) & (!g112) & (!g116)) + ((!g108) & (!sk[1]) & (!g110) & (g27) & (!g112) & (!g116)) + ((!g108) & (!sk[1]) & (!g110) & (!g27) & (!g112) & (g116)) + ((!g108) & (sk[1]) & (!g110) & (!g27) & (!g112) & (!g116)));
	assign g118 = (((g) & (!sk[2]) & (g10)) + ((!g) & (!sk[2]) & (g10)));
	assign g119 = (((!h) & (!sk[3]) & (g) & (!j)) + ((h) & (!sk[3]) & (g) & (j)));
	assign g120 = (((!k) & (!sk[4]) & (g1) & (!g119)) + ((!k) & (!sk[4]) & (g1) & (g119)));
	assign g121 = (((h) & (!g) & (!k) & (!g1) & (!sk[5]) & (!g99)) + ((!h) & (!g) & (k) & (!g1) & (!sk[5]) & (!g99)) + ((!h) & (!g) & (!k) & (!g1) & (!sk[5]) & (g99)) + ((h) & (g) & (k) & (g1) & (!sk[5]) & (!g99)));
	assign g122 = (((!sk[6]) & (h) & (!g) & (!k) & (!l) & (!g1)) + ((!sk[6]) & (!h) & (!g) & (k) & (!l) & (!g1)) + ((!sk[6]) & (!h) & (!g) & (!k) & (!l) & (g1)) + ((!sk[6]) & (h) & (g) & (k) & (!l) & (g1)));
	assign g123 = (((g3) & (!sk[7]) & (!g118) & (!g120) & (!g121) & (!g122)) + ((!g3) & (!sk[7]) & (!g118) & (g120) & (!g121) & (!g122)) + ((!g3) & (!sk[7]) & (!g118) & (!g120) & (!g121) & (g122)) + ((g3) & (!sk[7]) & (!g118) & (!g120) & (!g121) & (!g122)) + ((!g3) & (sk[7]) & (!g118) & (!g120) & (!g121) & (!g122)));
	assign g124 = (((!j) & (k) & (!i) & (!l) & (g1) & (g23)) + ((j) & (!k) & (!i) & (!l) & (g1) & (g23)) + ((!j) & (k) & (!i) & (!l) & (g1) & (g23)) + ((!j) & (k) & (!i) & (!l) & (g1) & (g23)));
	assign g125 = (((!f) & (!g10) & (!g3) & (!sk[9]) & (g124)) + ((!f) & (!g10) & (g3) & (!sk[9]) & (!g124)) + ((f) & (!g10) & (!g3) & (sk[9]) & (!g124)) + ((!f) & (!g10) & (!g3) & (sk[9]) & (!g124)));
	assign g126 = (((!d) & (!sk[10]) & (!e) & (c) & (!g101)) + ((!d) & (!sk[10]) & (!e) & (!c) & (g101)) + ((!d) & (!sk[10]) & (e) & (c) & (!g101)) + ((d) & (sk[10]) & (e) & (!c) & (!g101)));
	assign g127 = (((!g39) & (!sk[11]) & (!g123) & (g125) & (!g126)) + ((!g39) & (!sk[11]) & (!g123) & (!g125) & (g126)) + ((g39) & (sk[11]) & (!g123) & (!g125) & (!g126)) + ((!g39) & (!sk[11]) & (g123) & (g125) & (!g126)));
	assign g128 = (((!b) & (d) & (!e) & (a) & (g68) & (!g109)) + ((b) & (!d) & (!e) & (!a) & (g68) & (!g109)) + ((b) & (!d) & (e) & (!a) & (g68) & (!g109)) + ((b) & (!d) & (e) & (!a) & (!g68) & (g109)));
	assign g129 = (((g104) & (!g106) & (!g107) & (g117) & (g127) & (!g128)) + ((!g104) & (!g106) & (!g107) & (g117) & (g127) & (!g128)));
	assign g130 = (((g75) & (!sk[14]) & (g114)) + ((!g75) & (!sk[14]) & (g114)));
	assign g131 = (((!sk[15]) & (!b) & (!d) & (!e) & (!c) & (a)) + ((!sk[15]) & (b) & (!d) & (!e) & (!c) & (!a)) + ((!sk[15]) & (!b) & (!d) & (e) & (!c) & (!a)) + ((sk[15]) & (!b) & (!d) & (!e) & (!c) & (!a)) + ((!sk[15]) & (!b) & (!d) & (!e) & (!c) & (a)) + ((!sk[15]) & (!b) & (d) & (!e) & (!c) & (a)));
	assign g132 = (((b) & (!d) & (!e) & (!sk[16]) & (!c) & (!a)) + ((!b) & (!d) & (!e) & (!sk[16]) & (!c) & (a)) + ((!b) & (!d) & (!e) & (sk[16]) & (!c) & (!a)) + ((b) & (!d) & (!e) & (!sk[16]) & (c) & (a)) + ((!b) & (!d) & (e) & (!sk[16]) & (!c) & (!a)) + ((!b) & (d) & (!e) & (sk[16]) & (!c) & (!a)) + ((b) & (!d) & (e) & (!sk[16]) & (c) & (a)) + ((!b) & (!d) & (!e) & (!sk[16]) & (!c) & (a)));
	assign g133 = (((!sk[17]) & (!g130) & (g532)) + ((!sk[17]) & (!g130) & (g532)));
	assign g134 = (((sk[18]) & (!b) & (!e) & (!f) & (!a)) + ((sk[18]) & (!b) & (!e) & (!f) & (!a)) + ((!sk[18]) & (!b) & (!e) & (f) & (!a)) + ((!sk[18]) & (!b) & (!e) & (!f) & (a)) + ((!sk[18]) & (!b) & (!e) & (f) & (a)));
	assign g135 = (((!h) & (!sk[19]) & (g) & (!i)) + ((h) & (sk[19]) & (!g) & (i)));
	assign g136 = (((!h) & (!sk[20]) & (g) & (!i)) + ((h) & (!sk[20]) & (g) & (i)));
	assign g137 = (((m) & (!j) & (!l) & (!sk[21]) & (!g135) & (!g136)) + ((!m) & (!j) & (l) & (!sk[21]) & (!g135) & (!g136)) + ((!m) & (!j) & (!l) & (!sk[21]) & (!g135) & (g136)) + ((m) & (!j) & (l) & (!sk[21]) & (g135) & (!g136)) + ((m) & (j) & (!l) & (!sk[21]) & (!g135) & (g136)));
	assign g138 = (((g) & (!g99) & (!sk[22]) & (!g61) & (!g134) & (!g137)) + ((!g) & (!g99) & (!sk[22]) & (g61) & (!g134) & (!g137)) + ((!g) & (!g99) & (!sk[22]) & (!g61) & (!g134) & (g137)) + ((!g) & (!g99) & (!sk[22]) & (!g61) & (!g134) & (g137)) + ((g) & (g99) & (!sk[22]) & (g61) & (!g134) & (!g137)));
	assign g139 = (((m) & (!j) & (!k) & (!sk[23]) & (!i) & (!l)) + ((!m) & (!j) & (!k) & (!sk[23]) & (!i) & (l)) + ((!m) & (!j) & (k) & (!sk[23]) & (!i) & (!l)) + ((!m) & (!j) & (k) & (!sk[23]) & (!i) & (!l)) + ((!m) & (j) & (!k) & (sk[23]) & (!i) & (!l)) + ((!m) & (j) & (!k) & (sk[23]) & (!i) & (!l)));
	assign g140 = (((!d) & (e) & (!sk[24]) & (!c)) + ((!d) & (e) & (!sk[24]) & (c)));
	assign g141 = (((!m) & (!k) & (!sk[25]) & (i) & (!g41)) + ((!m) & (!k) & (!sk[25]) & (!i) & (g41)) + ((!m) & (k) & (!sk[25]) & (i) & (g41)));
	assign g142 = (((!g40) & (!sk[26]) & (!g139) & (g140) & (!g141)) + ((!g40) & (!sk[26]) & (!g139) & (!g140) & (g141)) + ((!g40) & (!sk[26]) & (!g139) & (g140) & (g141)) + ((g40) & (!sk[26]) & (g139) & (g140) & (!g141)));
	assign g143 = (((i) & (!g62) & (!g138) & (!g525) & (!sk[27]) & (!g142)) + ((!i) & (!g62) & (g138) & (!g525) & (!sk[27]) & (!g142)) + ((!i) & (!g62) & (!g138) & (!g525) & (!sk[27]) & (g142)) + ((!i) & (!g62) & (!g138) & (!g525) & (sk[27]) & (!g142)) + ((!i) & (!g62) & (!g138) & (!g525) & (sk[27]) & (!g142)) + ((!i) & (!g62) & (!g138) & (g525) & (sk[27]) & (!g142)));
	assign g144 = (((m) & (!k) & (!i) & (!sk[28]) & (!g133) & (!g143)) + ((!m) & (!k) & (i) & (!sk[28]) & (!g133) & (!g143)) + ((!m) & (!k) & (!i) & (!sk[28]) & (!g133) & (g143)) + ((!m) & (!k) & (!i) & (!sk[28]) & (!g133) & (g143)) + ((!m) & (!k) & (!i) & (!sk[28]) & (!g133) & (g143)) + ((!m) & (!k) & (!i) & (!sk[28]) & (g133) & (g143)));
	assign g145 = (((!j) & (!sk[29]) & (k)) + ((j) & (sk[29]) & (!k)));
	assign g146 = (((!f) & (!sk[30]) & (h) & (!g)) + ((!f) & (!sk[30]) & (h) & (g)));
	assign g147 = (((d) & (!sk[31]) & (!e) & (!g) & (!c) & (!a)) + ((!d) & (!sk[31]) & (!e) & (g) & (!c) & (!a)) + ((!d) & (!sk[31]) & (!e) & (!g) & (!c) & (a)) + ((!d) & (!sk[31]) & (e) & (g) & (c) & (a)));
	assign g148 = (((h) & (!g40) & (!g34) & (!g88) & (g147) & (!g132)) + ((!h) & (g40) & (!g34) & (!g88) & (!g147) & (!g132)) + ((h) & (!g40) & (g34) & (!g88) & (!g147) & (!g132)));
	assign g149 = (((!g146) & (g131) & (!sk[33]) & (!g148)) + ((!g146) & (g131) & (!sk[33]) & (!g148)) + ((!g146) & (!g131) & (sk[33]) & (!g148)));
	assign g150 = (((!g34) & (!sk[34]) & (g88)) + ((g34) & (sk[34]) & (!g88)));
	assign g151 = (((!f) & (!g) & (!i) & (!g150) & (!g131) & (!g132)) + ((!f) & (!g) & (!i) & (!g150) & (!g131) & (!g132)) + ((!f) & (!g) & (!i) & (!g150) & (g131) & (!g132)) + ((f) & (!g) & (!i) & (!g150) & (!g131) & (g132)));
	assign g152 = (((!sk[36]) & (!g) & (g134)) + ((sk[36]) & (g) & (!g134)));
	assign g153 = (((g86) & (!sk[37]) & (g152)) + ((!g86) & (!sk[37]) & (g152)));
	assign g154 = (((g54) & (!sk[38]) & (g153)) + ((!g54) & (!sk[38]) & (g153)));
	assign g155 = (((!e) & (c) & (!sk[39]) & (!a)) + ((e) & (c) & (!sk[39]) & (a)));
	assign g156 = (((!sk[40]) & (f) & (!g) & (!g81) & (!g87) & (!g155)) + ((!sk[40]) & (!f) & (!g) & (g81) & (!g87) & (!g155)) + ((!sk[40]) & (!f) & (!g) & (!g81) & (!g87) & (g155)) + ((!sk[40]) & (f) & (g) & (!g81) & (g87) & (!g155)) + ((!sk[40]) & (!f) & (g) & (!g81) & (g87) & (g155)));
	assign g157 = (((f) & (!g) & (!g113) & (!sk[41]) & (!g16) & (!g87)) + ((!f) & (!g) & (g113) & (!sk[41]) & (!g16) & (!g87)) + ((!f) & (!g) & (!g113) & (!sk[41]) & (!g16) & (g87)) + ((f) & (g) & (g113) & (!sk[41]) & (!g16) & (g87)) + ((!f) & (g) & (!g113) & (!sk[41]) & (g16) & (g87)));
	assign g158 = (((!d) & (e) & (!f) & (g) & (a) & (g87)));
	assign g159 = (((!g87) & (!sk[43]) & (g158) & (!g147)) + ((!g87) & (sk[43]) & (!g158) & (!g147)) + ((!g87) & (sk[43]) & (!g158) & (!g147)));
	assign g160 = (((!g89) & (!g110) & (!g154) & (!g156) & (!g157) & (g159)));
	assign g161 = (((g33) & (!sk[45]) & (!g34) & (!g36) & (!g71) & (!g151)) + ((!g33) & (!sk[45]) & (!g34) & (g36) & (!g71) & (!g151)) + ((!g33) & (!sk[45]) & (!g34) & (!g36) & (!g71) & (g151)) + ((!g33) & (!sk[45]) & (g34) & (g36) & (!g71) & (!g151)) + ((!g33) & (sk[45]) & (!g34) & (!g36) & (g71) & (!g151)));
	assign g162 = (((!sk[46]) & (!l) & (g86) & (!g15)) + ((!sk[46]) & (l) & (g86) & (g15)));
	assign g163 = (((h) & (!sk[47]) & (!g) & (!k) & (!g9) & (!g99)) + ((!h) & (!sk[47]) & (!g) & (k) & (!g9) & (!g99)) + ((!h) & (!sk[47]) & (!g) & (!k) & (!g9) & (g99)) + ((h) & (!sk[47]) & (g) & (k) & (g9) & (!g99)));
	assign g164 = (((g) & (!g10) & (!g21) & (!g98) & (!sk[48]) & (!g163)) + ((!g) & (!g10) & (!g21) & (!g98) & (!sk[48]) & (g163)) + ((!g) & (!g10) & (!g21) & (!g98) & (sk[48]) & (!g163)) + ((!g) & (!g10) & (g21) & (!g98) & (!sk[48]) & (!g163)) + ((!g) & (!g10) & (!g21) & (!g98) & (sk[48]) & (!g163)) + ((!g) & (!g10) & (!g21) & (!g98) & (sk[48]) & (!g163)));
	assign g165 = (((d) & (!e) & (!f) & (!c) & (!sk[49]) & (!g164)) + ((!d) & (!e) & (f) & (!c) & (!sk[49]) & (!g164)) + ((!d) & (!e) & (!f) & (!c) & (!sk[49]) & (g164)) + ((!d) & (!e) & (f) & (c) & (!sk[49]) & (!g164)) + ((d) & (!e) & (!f) & (!c) & (!sk[49]) & (!g164)) + ((d) & (!e) & (f) & (!c) & (!sk[49]) & (!g164)) + ((!d) & (e) & (!f) & (c) & (sk[49]) & (!g164)));
	assign g166 = (((!h) & (!n) & (i) & (!g62) & (g71) & (g147)) + ((!h) & (!n) & (i) & (g62) & (!g71) & (g147)));
	assign g167 = (((!sk[51]) & (l) & (!g41) & (!g86) & (!g9) & (!g140)) + ((!sk[51]) & (!l) & (!g41) & (g86) & (!g9) & (!g140)) + ((!sk[51]) & (!l) & (!g41) & (!g86) & (!g9) & (g140)) + ((!sk[51]) & (l) & (g41) & (g86) & (g9) & (g140)));
	assign g168 = (((!sk[52]) & (!g54) & (!g134) & (g135) & (!g167)) + ((!sk[52]) & (!g54) & (!g134) & (!g135) & (g167)) + ((sk[52]) & (!g54) & (!g134) & (!g135) & (!g167)) + ((!sk[52]) & (!g54) & (!g134) & (g135) & (!g167)) + ((!sk[52]) & (!g54) & (g134) & (g135) & (!g167)));
	assign g169 = (((!b) & (!c) & (g76) & (!sk[53]) & (!g33)) + ((!b) & (!c) & (!g76) & (!sk[53]) & (g33)) + ((b) & (!c) & (g76) & (!sk[53]) & (!g33)));
	assign g170 = (((!g42) & (!g43) & (!g166) & (g511) & (g168) & (!g169)) + ((!g42) & (!g43) & (!g166) & (g511) & (g168) & (!g169)));
	assign g171 = (((b) & (!e) & (!f) & (!sk[55]) & (!c) & (!g123)) + ((!b) & (!e) & (f) & (!sk[55]) & (!c) & (!g123)) + ((!b) & (!e) & (!f) & (!sk[55]) & (!c) & (g123)) + ((b) & (e) & (!f) & (!sk[55]) & (!c) & (!g123)) + ((!b) & (!e) & (f) & (!sk[55]) & (c) & (!g123)) + ((!b) & (!e) & (!f) & (sk[55]) & (c) & (!g123)));
	assign g172 = (((g133) & (!g161) & (!g162) & (!g165) & (g170) & (!g171)) + ((!g133) & (!g161) & (!g162) & (!g165) & (g170) & (!g171)));
	assign g173 = (((n) & (!m) & (!g144) & (!g518) & (g160) & (g172)) + ((!n) & (!m) & (g144) & (!g518) & (g160) & (g172)) + ((!n) & (!m) & (g144) & (g518) & (g160) & (g172)));
	assign g174 = (((h) & (!i) & (!sk[58]) & (!g15) & (!g147) & (!g525)) + ((!h) & (!i) & (!sk[58]) & (g15) & (!g147) & (!g525)) + ((!h) & (!i) & (!sk[58]) & (!g15) & (!g147) & (g525)) + ((!h) & (i) & (!sk[58]) & (g15) & (!g147) & (!g525)) + ((!h) & (i) & (!sk[58]) & (g15) & (g147) & (!g525)));
	assign g175 = (((k) & (!sk[59]) & (g174)) + ((!k) & (!sk[59]) & (g174)));
	assign g176 = (((!b) & (!d) & (!e) & (!f) & (sk[60]) & (!c)) + ((b) & (!d) & (!e) & (!f) & (!sk[60]) & (!c)) + ((!b) & (!d) & (e) & (!f) & (!sk[60]) & (!c)) + ((!b) & (!d) & (e) & (!f) & (!sk[60]) & (!c)) + ((!b) & (!d) & (!e) & (!f) & (!sk[60]) & (c)) + ((!b) & (!d) & (!e) & (!f) & (sk[60]) & (!c)) + ((!b) & (!d) & (!e) & (!f) & (sk[60]) & (!c)));
	assign g177 = (((!g4) & (!sk[61]) & (g504)) + ((g4) & (sk[61]) & (!g504)));
	assign g178 = (((!d) & (e) & (!sk[62]) & (!c)) + ((!d) & (!e) & (sk[62]) & (!c)) + ((!d) & (!e) & (sk[62]) & (c)));
	assign g179 = (((n) & (!m) & (!sk[63]) & (!g145) & (!g136) & (!g178)) + ((!n) & (!m) & (!sk[63]) & (g145) & (!g136) & (!g178)) + ((!n) & (!m) & (!sk[63]) & (!g145) & (!g136) & (g178)) + ((!n) & (!m) & (!sk[63]) & (g145) & (g136) & (!g178)));
	assign g180 = (((d) & (!e) & (!f) & (!sk[64]) & (!g) & (!c)) + ((!d) & (!e) & (f) & (!sk[64]) & (!g) & (!c)) + ((!d) & (!e) & (!f) & (!sk[64]) & (!g) & (c)) + ((!d) & (e) & (!f) & (!sk[64]) & (!g) & (c)) + ((d) & (!e) & (f) & (!sk[64]) & (!g) & (!c)) + ((!d) & (!e) & (f) & (!sk[64]) & (!g) & (c)) + ((!d) & (!e) & (f) & (!sk[64]) & (!g) & (c)) + ((!d) & (!e) & (f) & (!sk[64]) & (!g) & (c)));
	assign g181 = (((h) & (!k) & (!sk[65]) & (!g9) & (!g99) & (!g180)) + ((!h) & (!k) & (!sk[65]) & (g9) & (!g99) & (!g180)) + ((!h) & (!k) & (!sk[65]) & (!g9) & (!g99) & (g180)) + ((h) & (!k) & (!sk[65]) & (g9) & (g99) & (g180)));
	assign g182 = (((!h) & (!sk[66]) & (j) & (!i)) + ((h) & (!sk[66]) & (j) & (i)));
	assign g183 = (((!k) & (!g1) & (g93) & (!sk[67]) & (!g182)) + ((!k) & (!g1) & (!g93) & (!sk[67]) & (g182)) + ((!k) & (g1) & (g93) & (!sk[67]) & (g182)));
	assign g184 = (((!g15) & (!sk[68]) & (g16) & (!g146)) + ((g15) & (!sk[68]) & (g16) & (g146)));
	assign g185 = (((d) & (!e) & (g40) & (!c) & (a) & (!g146)) + ((!d) & (e) & (!g40) & (!c) & (a) & (g146)) + ((!d) & (e) & (!g40) & (c) & (a) & (g146)));
	assign g186 = (((h) & (!g40) & (!g34) & (!sk[70]) & (!g88) & (!g147)) + ((!h) & (!g40) & (g34) & (!sk[70]) & (!g88) & (!g147)) + ((h) & (!g40) & (!g34) & (!sk[70]) & (!g88) & (g147)) + ((!h) & (!g40) & (!g34) & (!sk[70]) & (!g88) & (g147)) + ((h) & (!g40) & (g34) & (!sk[70]) & (!g88) & (!g147)) + ((!h) & (g40) & (!g34) & (sk[70]) & (!g88) & (!g147)));
	assign g187 = (((h) & (!g) & (!g184) & (!sk[71]) & (!g185) & (!g186)) + ((!h) & (!g) & (g184) & (!sk[71]) & (!g185) & (!g186)) + ((!h) & (!g) & (!g184) & (!sk[71]) & (!g185) & (g186)) + ((!h) & (!g) & (!g184) & (sk[71]) & (!g185) & (!g186)) + ((!h) & (!g) & (!g184) & (sk[71]) & (!g185) & (!g186)) + ((!h) & (!g) & (!g184) & (sk[71]) & (!g185) & (!g186)));
	assign g188 = (((b) & (!sk[72]) & (!d) & (!g40) & (!c) & (!a)) + ((!b) & (!sk[72]) & (!d) & (g40) & (!c) & (!a)) + ((!b) & (!sk[72]) & (!d) & (!g40) & (!c) & (a)) + ((!b) & (!sk[72]) & (!d) & (g40) & (c) & (a)) + ((b) & (!sk[72]) & (!d) & (g40) & (!c) & (a)) + ((b) & (!sk[72]) & (!d) & (g40) & (!c) & (!a)));
	assign g189 = (((b) & (e) & (!k) & (!a) & (g15) & (g119)));
	assign g190 = (((g145) & (!g15) & (!sk[74]) & (!g187) & (!g188) & (!g189)) + ((!g145) & (!g15) & (!sk[74]) & (!g187) & (!g188) & (g189)) + ((!g145) & (!g15) & (sk[74]) & (!g187) & (!g188) & (!g189)) + ((!g145) & (!g15) & (!sk[74]) & (g187) & (!g188) & (!g189)) + ((!g145) & (!g15) & (sk[74]) & (!g187) & (!g188) & (!g189)) + ((!g145) & (!g15) & (!sk[74]) & (g187) & (!g188) & (!g189)));
	assign g191 = (((!b) & (!d) & (e) & (!f) & (!sk[75]) & (!c)) + ((b) & (!d) & (!e) & (!f) & (!sk[75]) & (!c)) + ((!b) & (!d) & (!e) & (!f) & (!sk[75]) & (c)) + ((!b) & (!d) & (!e) & (!f) & (sk[75]) & (!c)) + ((b) & (d) & (!e) & (!f) & (!sk[75]) & (c)) + ((!b) & (d) & (e) & (f) & (!sk[75]) & (c)) + ((!b) & (!d) & (!e) & (!f) & (sk[75]) & (!c)));
	assign g192 = (((!sk[76]) & (!h) & (g) & (!g191)) + ((!sk[76]) & (h) & (g) & (!g191)));
	assign g193 = (((!m) & (g145) & (!sk[77]) & (!i)) + ((!m) & (g145) & (!sk[77]) & (i)));
	assign g194 = (((!sk[78]) & (b) & (!d) & (!e) & (!f) & (!h)) + ((!sk[78]) & (!b) & (!d) & (e) & (!f) & (!h)) + ((!sk[78]) & (!b) & (!d) & (!e) & (!f) & (h)) + ((!sk[78]) & (b) & (d) & (!e) & (f) & (h)) + ((!sk[78]) & (b) & (!d) & (e) & (!f) & (h)));
	assign g195 = (((n) & (!g135) & (!g176) & (g192) & (g193) & (!g194)) + ((n) & (!g135) & (!g176) & (!g192) & (g193) & (g194)) + ((n) & (g135) & (!g176) & (!g192) & (g193) & (!g194)));
	assign g196 = (((g179) & (!sk[80]) & (!g181) & (!g183) & (!g190) & (!g195)) + ((!g179) & (!sk[80]) & (!g181) & (g183) & (!g190) & (!g195)) + ((!g179) & (!sk[80]) & (!g181) & (!g183) & (!g190) & (g195)) + ((!g179) & (sk[80]) & (!g181) & (!g183) & (g190) & (!g195)));
	assign g197 = (((!sk[81]) & (n) & (!m) & (!k) & (!g178) & (!g191)) + ((!sk[81]) & (!n) & (!m) & (k) & (!g178) & (!g191)) + ((!sk[81]) & (!n) & (!m) & (!k) & (!g178) & (g191)) + ((!sk[81]) & (!n) & (!m) & (k) & (!g178) & (!g191)) + ((!sk[81]) & (n) & (!m) & (k) & (!g178) & (!g191)));
	assign g198 = (((!h) & (!g) & (g99) & (!sk[82]) & (!g197)) + ((!h) & (!g) & (!g99) & (!sk[82]) & (g197)) + ((h) & (g) & (!g99) & (!sk[82]) & (g197)));
	assign g199 = (((!sk[83]) & (!n) & (!m) & (g93) & (!g180)) + ((!sk[83]) & (!n) & (!m) & (!g93) & (g180)) + ((!sk[83]) & (n) & (!m) & (g93) & (!g180)) + ((!sk[83]) & (!n) & (!m) & (!g93) & (g180)));
	assign g200 = (((!h) & (!k) & (!sk[84]) & (g99) & (!g199)) + ((!h) & (!k) & (!sk[84]) & (!g99) & (g199)) + ((h) & (k) & (!sk[84]) & (!g99) & (g199)));
	assign g201 = (((!f) & (!g) & (!i) & (g150) & (!g131) & (!g132)) + ((!f) & (g) & (!i) & (!g150) & (!g131) & (!g132)) + ((f) & (g) & (!i) & (!g150) & (!g131) & (!g132)));
	assign g202 = (((!sk[86]) & (!j) & (k) & (!l)) + ((sk[86]) & (!j) & (!k) & (!l)) + ((!sk[86]) & (!j) & (k) & (!l)) + ((!sk[86]) & (!j) & (k) & (!l)));
	assign g203 = (((!sk[87]) & (!g15) & (g202)) + ((sk[87]) & (g15) & (!g202)));
	assign g204 = (((j) & (!k) & (!sk[88]) & (!l) & (!g15) & (!g152)) + ((!j) & (!k) & (!sk[88]) & (l) & (!g15) & (!g152)) + ((!j) & (!k) & (!sk[88]) & (!l) & (!g15) & (g152)) + ((!j) & (k) & (!sk[88]) & (!l) & (g15) & (g152)));
	assign g205 = (((!sk[89]) & (!n) & (!m) & (k) & (!g134)) + ((!sk[89]) & (!n) & (!m) & (!k) & (g134)) + ((!sk[89]) & (!n) & (m) & (k) & (!g134)));
	assign g206 = (((!g) & (!l) & (!sk[90]) & (g10) & (!g58)) + ((!g) & (!l) & (!sk[90]) & (!g10) & (g58)) + ((g) & (l) & (!sk[90]) & (g10) & (!g58)) + ((g) & (l) & (!sk[90]) & (!g10) & (g58)));
	assign g207 = (((!sk[91]) & (j) & (!g71) & (!g147) & (!g205) & (!g206)) + ((!sk[91]) & (!j) & (!g71) & (g147) & (!g205) & (!g206)) + ((!sk[91]) & (!j) & (!g71) & (!g147) & (!g205) & (g206)) + ((!sk[91]) & (!j) & (!g71) & (!g147) & (g205) & (g206)) + ((!sk[91]) & (!j) & (g71) & (g147) & (!g205) & (!g206)));
	assign g208 = (((!i) & (!g147) & (!g201) & (!g203) & (!g204) & (!g207)) + ((i) & (!g147) & (!g201) & (!g203) & (!g204) & (!g207)) + ((!i) & (!g147) & (!g201) & (!g203) & (!g204) & (!g207)));
	assign g209 = (((g4) & (!g198) & (!sk[93]) & (!g497) & (!g200) & (!g208)) + ((!g4) & (!g198) & (!sk[93]) & (g497) & (!g200) & (!g208)) + ((!g4) & (!g198) & (!sk[93]) & (!g497) & (!g200) & (g208)) + ((!g4) & (!g198) & (!sk[93]) & (!g497) & (!g200) & (g208)) + ((!g4) & (!g198) & (!sk[93]) & (g497) & (!g200) & (g208)));
	assign g210 = (((!sk[94]) & (f) & (!g) & (!g150) & (!g131) & (!g132)) + ((!sk[94]) & (!f) & (!g) & (g150) & (!g131) & (!g132)) + ((!sk[94]) & (!f) & (!g) & (!g150) & (!g131) & (g132)) + ((sk[94]) & (!f) & (!g) & (!g150) & (!g131) & (!g132)) + ((!sk[94]) & (f) & (!g) & (!g150) & (!g131) & (g132)) + ((sk[94]) & (!f) & (!g) & (!g150) & (g131) & (!g132)));
	assign g211 = (((!sk[95]) & (!h) & (g) & (!i)) + ((sk[95]) & (!h) & (!g) & (!i)) + ((!sk[95]) & (!h) & (g) & (!i)) + ((!sk[95]) & (!h) & (g) & (i)));
	assign g212 = (((!sk[96]) & (!j) & (i) & (!l)) + ((sk[96]) & (!j) & (!i) & (l)));
	assign g213 = (((!sk[97]) & (d) & (!e) & (!c) & (!a) & (!g146)) + ((!sk[97]) & (!d) & (!e) & (c) & (!a) & (!g146)) + ((!sk[97]) & (!d) & (!e) & (!c) & (!a) & (g146)) + ((!sk[97]) & (!d) & (e) & (!c) & (a) & (g146)) + ((!sk[97]) & (!d) & (e) & (c) & (a) & (g146)));
	assign g214 = (((!g15) & (!g148) & (g184) & (g212) & (!sk[98]) & (!g213)) + ((g15) & (!g148) & (!g184) & (!g212) & (!sk[98]) & (!g213)) + ((!g15) & (!g148) & (g184) & (!g212) & (!sk[98]) & (!g213)) + ((!g15) & (!g148) & (!g184) & (!g212) & (!sk[98]) & (g213)) + ((g15) & (g148) & (!g184) & (g212) & (!sk[98]) & (!g213)) + ((g15) & (!g148) & (!g184) & (g212) & (!sk[98]) & (g213)));
	assign g215 = (((!n) & (!sk[99]) & (!g211) & (g64) & (!g134) & (!g214)) + ((!n) & (!sk[99]) & (!g211) & (!g64) & (!g134) & (g214)) + ((n) & (!sk[99]) & (!g211) & (!g64) & (!g134) & (!g214)) + ((!n) & (sk[99]) & (!g211) & (!g64) & (!g134) & (!g214)) + ((!n) & (!sk[99]) & (g211) & (g64) & (!g134) & (!g214)) + ((!n) & (!sk[99]) & (!g211) & (g64) & (g134) & (!g214)));
	assign g216 = (((!j) & (!g71) & (!g118) & (!g134) & (!g210) & (g215)) + ((j) & (!g71) & (!g118) & (!g134) & (!g210) & (g215)) + ((j) & (!g71) & (!g118) & (g134) & (!g210) & (g215)) + ((!j) & (!g71) & (!g118) & (!g134) & (g210) & (g215)) + ((!j) & (!g71) & (!g118) & (g134) & (g210) & (g215)));
	assign g217 = (((!g175) & (!g177) & (g160) & (g196) & (g209) & (g216)));
	assign g218 = (((!sk[102]) & (!m) & (j) & (!k)) + ((sk[102]) & (!m) & (!j) & (k)));
	assign g219 = (((!n) & (g218) & (!sk[103]) & (!i)) + ((n) & (g218) & (!sk[103]) & (i)));
	assign g220 = (((k) & (!g10) & (!g199) & (!g194) & (!sk[104]) & (!g219)) + ((!k) & (!g10) & (g199) & (!g194) & (!sk[104]) & (!g219)) + ((!k) & (!g10) & (!g199) & (g194) & (!sk[104]) & (g219)) + ((!k) & (!g10) & (!g199) & (!g194) & (!sk[104]) & (g219)) + ((k) & (g10) & (g199) & (!g194) & (!sk[104]) & (!g219)));
	assign g221 = (((!g44) & (!j) & (g71) & (!sk[105]) & (!g132)) + ((!g44) & (!j) & (!g71) & (!sk[105]) & (g132)) + ((g44) & (!j) & (g71) & (!sk[105]) & (!g132)));
	assign g222 = (((!n) & (!sk[106]) & (!g218) & (!g135) & (!g176) & (g221)) + ((n) & (!sk[106]) & (!g218) & (!g135) & (!g176) & (!g221)) + ((!n) & (sk[106]) & (!g218) & (!g135) & (!g176) & (!g221)) + ((!n) & (!sk[106]) & (!g218) & (g135) & (!g176) & (!g221)) + ((!n) & (sk[106]) & (!g218) & (!g135) & (!g176) & (!g221)) + ((!n) & (!sk[106]) & (!g218) & (g135) & (g176) & (!g221)));
	assign g223 = (((!sk[107]) & (!k) & (l) & (!g15)) + ((!sk[107]) & (k) & (l) & (g15)));
	assign g224 = (((!sk[108]) & (!j) & (i) & (!g223)) + ((sk[108]) & (!j) & (!i) & (g223)));
	assign g225 = (((g39) & (!sk[109]) & (!f) & (!g) & (!g10) & (!g176)) + ((!g39) & (!sk[109]) & (!f) & (g) & (!g10) & (!g176)) + ((!g39) & (!sk[109]) & (!f) & (!g) & (!g10) & (g176)) + ((!g39) & (sk[109]) & (!f) & (!g) & (g10) & (!g176)) + ((!g39) & (sk[109]) & (!f) & (!g) & (g10) & (!g176)));
	assign g226 = (((!f) & (!g10) & (!sk[110]) & (g43) & (!g225)) + ((!f) & (!g10) & (!sk[110]) & (!g43) & (g225)) + ((!f) & (!g10) & (sk[110]) & (!g43) & (!g225)) + ((!f) & (!g10) & (!sk[110]) & (g43) & (!g225)) + ((!f) & (!g10) & (!sk[110]) & (g43) & (!g225)));
	assign g227 = (((!n) & (!sk[111]) & (g178) & (!g191)) + ((!n) & (!sk[111]) & (g178) & (!g191)) + ((n) & (sk[111]) & (!g178) & (g191)));
	assign g228 = (((g218) & (!g4) & (!g136) & (!sk[112]) & (!g226) & (!g227)) + ((!g218) & (!g4) & (g136) & (!sk[112]) & (!g226) & (!g227)) + ((!g218) & (!g4) & (!g136) & (!sk[112]) & (!g226) & (g227)) + ((!g218) & (g4) & (!g136) & (sk[112]) & (!g226) & (!g227)) + ((g218) & (!g4) & (g136) & (!sk[112]) & (!g226) & (!g227)));
	assign g229 = (((n) & (!m) & (!k) & (!sk[113]) & (!g93) & (!g180)) + ((!n) & (!m) & (k) & (!sk[113]) & (!g93) & (!g180)) + ((!n) & (!m) & (!k) & (!sk[113]) & (!g93) & (g180)) + ((n) & (!m) & (k) & (!sk[113]) & (g93) & (!g180)) + ((!n) & (!m) & (k) & (!sk[113]) & (!g93) & (g180)));
	assign g230 = (((f) & (!a) & (!g140) & (!g131) & (!sk[114]) & (!g178)) + ((f) & (!a) & (!g140) & (!g131) & (!sk[114]) & (!g178)) + ((!f) & (!a) & (g140) & (!g131) & (!sk[114]) & (!g178)) + ((!f) & (!a) & (!g140) & (!g131) & (!sk[114]) & (g178)) + ((!f) & (!a) & (!g140) & (g131) & (sk[114]) & (!g178)) + ((f) & (!a) & (!g140) & (!g131) & (!sk[114]) & (g178)) + ((!f) & (!a) & (!g140) & (g131) & (!sk[114]) & (g178)));
	assign g231 = (((h) & (!j) & (i) & (!g71) & (g229) & (!g230)) + ((h) & (!j) & (!i) & (g71) & (!g229) & (!g230)));
	assign g232 = (((!g15) & (!g29) & (g149) & (!g224) & (!g228) & (!g231)) + ((!g15) & (!g29) & (!g149) & (!g224) & (!g228) & (!g231)) + ((!g15) & (!g29) & (!g149) & (!g224) & (!g228) & (!g231)));
	assign g233 = (((!h) & (!g) & (!sk[117]) & (j) & (!g205)) + ((!h) & (!g) & (!sk[117]) & (!j) & (g205)) + ((h) & (!g) & (!sk[117]) & (!j) & (g205)) + ((h) & (!g) & (!sk[117]) & (!j) & (g205)));
	assign g234 = (((g54) & (!sk[118]) & (!g118) & (!g133) & (!g197) & (!g233)) + ((!g54) & (!sk[118]) & (!g118) & (g133) & (!g197) & (!g233)) + ((!g54) & (!sk[118]) & (!g118) & (!g133) & (!g197) & (g233)) + ((!g54) & (!sk[118]) & (!g118) & (g133) & (!g197) & (!g233)) + ((!g54) & (!sk[118]) & (!g118) & (g133) & (!g197) & (!g233)) + ((!g54) & (sk[118]) & (!g118) & (!g133) & (!g197) & (!g233)) + ((!g54) & (sk[118]) & (!g118) & (!g133) & (!g197) & (!g233)));
	assign g235 = (((!sk[119]) & (g196) & (!g220) & (!g222) & (!g232) & (!g234)) + ((!sk[119]) & (!g196) & (!g220) & (g222) & (!g232) & (!g234)) + ((!sk[119]) & (!g196) & (!g220) & (!g222) & (!g232) & (g234)) + ((!sk[119]) & (g196) & (!g220) & (g222) & (g232) & (g234)));
	assign g236 = (((!j) & (!k) & (!sk[120]) & (l) & (!g174)) + ((!j) & (!k) & (!sk[120]) & (!l) & (g174)) + ((j) & (k) & (!sk[120]) & (!l) & (g174)) + ((!j) & (!k) & (!sk[120]) & (l) & (g174)));
	assign g237 = (((n) & (!sk[121]) & (m) & (!g133)) + ((!n) & (!sk[121]) & (m) & (!g133)) + ((!n) & (!sk[121]) & (m) & (g133)));
	assign g238 = (((!n) & (!g118) & (!sk[122]) & (g226) & (!g227)) + ((!n) & (!g118) & (!sk[122]) & (!g226) & (g227)) + ((n) & (!g118) & (sk[122]) & (!g226) & (!g227)) + ((!n) & (g118) & (sk[122]) & (!g226) & (!g227)));
	assign g239 = (((!m) & (!sk[123]) & (g211) & (!g227)) + ((!m) & (!sk[123]) & (g211) & (!g227)) + ((!m) & (sk[123]) & (!g211) & (g227)));
	assign g240 = (((!n) & (j) & (k) & (!g497) & (g238) & (!g239)) + ((!n) & (j) & (k) & (!g497) & (!g238) & (!g239)) + ((n) & (j) & (k) & (!g497) & (!g238) & (!g239)));
	assign g241 = (((j) & (!sk[125]) & (!k) & (!l) & (!g15) & (!g118)) + ((!j) & (!sk[125]) & (!k) & (l) & (!g15) & (!g118)) + ((!j) & (!sk[125]) & (!k) & (!l) & (!g15) & (g118)) + ((j) & (!sk[125]) & (k) & (!l) & (g15) & (g118)) + ((!j) & (!sk[125]) & (!k) & (l) & (g15) & (g118)));
	assign g242 = (((g) & (!k) & (!sk[126]) & (!l) & (!g15) & (!g58)) + ((!g) & (!k) & (!sk[126]) & (l) & (!g15) & (!g58)) + ((!g) & (!k) & (!sk[126]) & (!l) & (!g15) & (g58)) + ((g) & (!k) & (!sk[126]) & (!l) & (g15) & (g58)) + ((g) & (!k) & (!sk[126]) & (l) & (g15) & (g58)));
	assign g243 = (((j) & (!g55) & (!sk[127]) & (!g134) & (!g241) & (!g242)) + ((!j) & (!g55) & (!sk[127]) & (g134) & (!g241) & (!g242)) + ((!j) & (!g55) & (!sk[127]) & (!g134) & (!g241) & (g242)) + ((j) & (g55) & (!sk[127]) & (!g134) & (!g241) & (!g242)) + ((!j) & (!g55) & (sk[127]) & (!g134) & (g241) & (!g242)));
	assign g244 = (((n) & (!m) & (!j) & (!k) & (!sk[0]) & (!l)) + ((!n) & (!m) & (j) & (!k) & (!sk[0]) & (!l)) + ((!n) & (!m) & (!j) & (!k) & (!sk[0]) & (l)) + ((!n) & (m) & (j) & (!k) & (!sk[0]) & (!l)) + ((!n) & (m) & (j) & (!k) & (!sk[0]) & (l)));
	assign g245 = (((!n) & (!sk[1]) & (g60) & (!g147)) + ((!n) & (!sk[1]) & (g60) & (g147)));
	assign g246 = (((!h) & (!g145) & (g199) & (!sk[2]) & (!g245)) + ((!h) & (!g145) & (!g199) & (!sk[2]) & (g245)) + ((!h) & (!g145) & (!g199) & (sk[2]) & (!g245)) + ((!h) & (!g145) & (!g199) & (sk[2]) & (!g245)) + ((!h) & (!g145) & (!g199) & (sk[2]) & (!g245)));
	assign g247 = (((h) & (!g) & (!sk[3]) & (!j) & (!g176) & (!g194)) + ((!h) & (!g) & (!sk[3]) & (j) & (!g176) & (!g194)) + ((!h) & (!g) & (!sk[3]) & (!j) & (!g176) & (g194)) + ((!h) & (!g) & (!sk[3]) & (j) & (!g176) & (g194)) + ((h) & (!g) & (!sk[3]) & (j) & (!g176) & (!g194)));
	assign g248 = (((!h) & (!sk[4]) & (!j) & (i) & (!g229)) + ((!h) & (!sk[4]) & (!j) & (!i) & (g229)) + ((!h) & (!sk[4]) & (j) & (i) & (g229)) + ((h) & (!sk[4]) & (j) & (!i) & (g229)));
	assign g249 = (((!n) & (!m) & (!k) & (g119) & (!g178) & (!g191)) + ((n) & (!m) & (!k) & (g119) & (!g178) & (!g191)));
	assign g250 = (((k) & (!sk[6]) & (!g1) & (!g247) & (!g248) & (!g249)) + ((!k) & (!sk[6]) & (!g1) & (g247) & (!g248) & (!g249)) + ((!k) & (!sk[6]) & (!g1) & (!g247) & (!g248) & (g249)) + ((k) & (!sk[6]) & (!g1) & (!g247) & (!g248) & (!g249)) + ((!k) & (sk[6]) & (!g1) & (!g247) & (!g248) & (!g249)) + ((!k) & (!sk[6]) & (!g1) & (g247) & (!g248) & (!g249)));
	assign g251 = (((g201) & (!g243) & (!g244) & (!sk[7]) & (!g246) & (!g250)) + ((!g201) & (!g243) & (g244) & (!sk[7]) & (!g246) & (!g250)) + ((!g201) & (!g243) & (!g244) & (!sk[7]) & (!g246) & (g250)) + ((!g201) & (!g243) & (!g244) & (!sk[7]) & (g246) & (g250)) + ((!g201) & (!g243) & (!g244) & (!sk[7]) & (g246) & (g250)));
	assign g252 = (((g236) & (!g237) & (!g190) & (!sk[8]) & (!g240) & (!g251)) + ((!g236) & (!g237) & (g190) & (!sk[8]) & (!g240) & (!g251)) + ((!g236) & (!g237) & (!g190) & (!sk[8]) & (!g240) & (g251)) + ((!g236) & (g237) & (g190) & (!sk[8]) & (!g240) & (g251)) + ((!g236) & (!g237) & (g190) & (!sk[8]) & (!g240) & (g251)));
	assign g253 = (((!sk[9]) & (!h) & (g147) & (!g525)) + ((sk[9]) & (!h) & (!g147) & (g525)) + ((!sk[9]) & (h) & (g147) & (g525)));
	assign g254 = (((h) & (!g) & (!j) & (!sk[10]) & (!k) & (!g134)) + ((!h) & (!g) & (j) & (!sk[10]) & (!k) & (!g134)) + ((!h) & (!g) & (!j) & (!sk[10]) & (!k) & (g134)) + ((h) & (!g) & (!j) & (!sk[10]) & (!k) & (!g134)) + ((h) & (!g) & (!j) & (!sk[10]) & (k) & (!g134)) + ((!h) & (g) & (j) & (!sk[10]) & (!k) & (!g134)));
	assign g255 = (((j) & (!l) & (!sk[11]) & (!g15) & (!g253) & (!g254)) + ((!j) & (!l) & (!sk[11]) & (g15) & (!g253) & (!g254)) + ((!j) & (!l) & (!sk[11]) & (!g15) & (!g253) & (g254)) + ((!j) & (l) & (!sk[11]) & (g15) & (!g253) & (g254)) + ((j) & (l) & (!sk[11]) & (g15) & (!g253) & (!g254)));
	assign g256 = (((!sk[12]) & (!m) & (k) & (!l)) + ((!sk[12]) & (m) & (k) & (l)));
	assign g257 = (((j) & (!k) & (!g62) & (!g532) & (!sk[13]) & (!g210)) + ((!j) & (!k) & (g62) & (!g532) & (!sk[13]) & (!g210)) + ((!j) & (!k) & (!g62) & (!g532) & (!sk[13]) & (g210)) + ((!j) & (!k) & (g62) & (!g532) & (!sk[13]) & (!g210)) + ((j) & (!k) & (g62) & (!g532) & (!sk[13]) & (!g210)));
	assign g258 = (((!sk[14]) & (!m) & (k) & (!l)) + ((!sk[14]) & (!m) & (k) & (l)));
	assign g259 = (((h) & (!sk[15]) & (!g) & (!j) & (!g62) & (!g134)) + ((!h) & (!sk[15]) & (!g) & (j) & (!g62) & (!g134)) + ((!h) & (!sk[15]) & (!g) & (!j) & (!g62) & (g134)) + ((!h) & (!sk[15]) & (g) & (j) & (g62) & (!g134)));
	assign g260 = (((!h) & (!n) & (!g58) & (!g180) & (!g258) & (!g259)) + ((!h) & (!n) & (!g58) & (!g180) & (!g258) & (!g259)) + ((!h) & (!n) & (!g58) & (!g180) & (!g258) & (!g259)) + ((!h) & (!n) & (!g58) & (!g180) & (!g258) & (!g259)));
	assign g261 = (((g153) & (!g133) & (!g256) & (!g257) & (!sk[17]) & (!g260)) + ((!g153) & (!g133) & (g256) & (!g257) & (!sk[17]) & (!g260)) + ((!g153) & (!g133) & (!g256) & (!g257) & (!sk[17]) & (g260)) + ((!g153) & (!g133) & (!g256) & (!g257) & (!sk[17]) & (g260)) + ((!g153) & (g133) & (!g256) & (!g257) & (!sk[17]) & (g260)));
	assign g262 = (((!m) & (!sk[18]) & (k) & (!l)) + ((!m) & (sk[18]) & (!k) & (l)));
	assign g263 = (((!h) & (!g58) & (g93) & (!sk[19]) & (!g504)) + ((!h) & (!g58) & (!g93) & (!sk[19]) & (g504)) + ((!h) & (!g58) & (!g93) & (!sk[19]) & (g504)) + ((!h) & (!g58) & (!g93) & (!sk[19]) & (g504)));
	assign g264 = (((n) & (!sk[20]) & (m) & (!j) & (!l) & (!g225)) + ((n) & (!sk[20]) & (!m) & (j) & (!l) & (!g225)) + ((!n) & (!sk[20]) & (!m) & (j) & (!l) & (!g225)) + ((n) & (!sk[20]) & (!m) & (!j) & (!l) & (!g225)) + ((!n) & (!sk[20]) & (!m) & (!j) & (!l) & (g225)) + ((n) & (!sk[20]) & (!m) & (!j) & (!l) & (!g225)));
	assign g265 = (((g247) & (!g258) & (!sk[21]) & (!g262) & (!g263) & (!g264)) + ((!g247) & (!g258) & (!sk[21]) & (g262) & (!g263) & (!g264)) + ((!g247) & (!g258) & (!sk[21]) & (!g262) & (!g263) & (g264)) + ((!g247) & (!g258) & (!sk[21]) & (!g262) & (!g263) & (g264)) + ((!g247) & (!g258) & (!sk[21]) & (!g262) & (!g263) & (g264)) + ((!g247) & (!g258) & (!sk[21]) & (!g262) & (g263) & (g264)) + ((!g247) & (!g258) & (!sk[21]) & (!g262) & (g263) & (g264)));
	assign g266 = (((j) & (!i) & (!g147) & (!sk[22]) & (!g151) & (!g223)) + ((!j) & (!i) & (g147) & (!sk[22]) & (!g151) & (!g223)) + ((!j) & (!i) & (!g147) & (!sk[22]) & (!g151) & (g223)) + ((!j) & (!i) & (!g147) & (!sk[22]) & (!g151) & (g223)) + ((!j) & (i) & (g147) & (!sk[22]) & (!g151) & (g223)));
	assign g267 = (((n) & (!g64) & (!g69) & (!sk[23]) & (!g147) & (!g130)) + ((!n) & (!g64) & (g69) & (!sk[23]) & (!g147) & (!g130)) + ((!n) & (!g64) & (!g69) & (!sk[23]) & (!g147) & (g130)) + ((!n) & (!g64) & (g69) & (!sk[23]) & (g147) & (!g130)) + ((!n) & (g64) & (!g69) & (!sk[23]) & (!g147) & (g130)));
	assign g268 = (((!h) & (!sk[24]) & (!j) & (k) & (!i)) + ((!h) & (!sk[24]) & (!j) & (!k) & (i)) + ((h) & (!sk[24]) & (!j) & (k) & (!i)) + ((!h) & (!sk[24]) & (!j) & (!k) & (i)) + ((!h) & (!sk[24]) & (!j) & (k) & (i)) + ((h) & (sk[24]) & (j) & (!k) & (!i)));
	assign g269 = (((n) & (!m) & (l) & (g93) & (!g180) & (g268)) + ((!n) & (!m) & (l) & (!g93) & (g180) & (g268)));
	assign g270 = (((!f) & (!g10) & (g2) & (!sk[26]) & (!g43)) + ((!f) & (!g10) & (!g2) & (!sk[26]) & (g43)) + ((f) & (g10) & (g2) & (!sk[26]) & (g43)));
	assign g271 = (((!g119) & (!sk[27]) & (!g270) & (g227) & (!g262)) + ((!g119) & (!sk[27]) & (!g270) & (g227) & (!g262)) + ((!g119) & (!sk[27]) & (!g270) & (!g227) & (g262)) + ((!g119) & (sk[27]) & (!g270) & (!g227) & (!g262)) + ((!g119) & (!sk[27]) & (!g270) & (!g227) & (g262)));
	assign g272 = (((!sk[28]) & (g227) & (!g479) & (!g267) & (!g269) & (!g271)) + ((!sk[28]) & (!g227) & (!g479) & (g267) & (!g269) & (!g271)) + ((!sk[28]) & (!g227) & (!g479) & (!g267) & (!g269) & (g271)) + ((!sk[28]) & (g227) & (!g479) & (!g267) & (!g269) & (g271)) + ((!sk[28]) & (!g227) & (g479) & (!g267) & (!g269) & (g271)));
	assign g273 = (((g238) & (!g258) & (!g266) & (!g215) & (!sk[29]) & (!g272)) + ((!g238) & (!g258) & (g266) & (!g215) & (!sk[29]) & (!g272)) + ((!g238) & (!g258) & (!g266) & (!g215) & (!sk[29]) & (g272)) + ((!g238) & (!g258) & (!g266) & (g215) & (!sk[29]) & (g272)) + ((!g238) & (!g258) & (!g266) & (g215) & (!sk[29]) & (g272)));
	assign g274 = (((g255) & (!g261) & (!sk[30]) & (!g265) & (!g486) & (!g273)) + ((!g255) & (!g261) & (!sk[30]) & (g265) & (!g486) & (!g273)) + ((!g255) & (!g261) & (!sk[30]) & (!g265) & (!g486) & (g273)) + ((!g255) & (g261) & (!sk[30]) & (!g265) & (g486) & (g273)) + ((!g255) & (!g261) & (!sk[30]) & (g265) & (g486) & (g273)));
	assign g275 = (((!g) & (!sk[31]) & (g23) & (!g54)) + ((!g) & (!sk[31]) & (g23) & (g54)));
	assign g276 = (((f) & (!h) & (!sk[32]) & (!g) & (!g61) & (!g63)) + ((!f) & (!h) & (!sk[32]) & (g) & (!g61) & (!g63)) + ((!f) & (!h) & (!sk[32]) & (!g) & (!g61) & (g63)) + ((!f) & (!h) & (!sk[32]) & (g) & (!g61) & (g63)) + ((!f) & (!h) & (!sk[32]) & (g) & (g61) & (g63)));
	assign g277 = (((!f) & (!h) & (g) & (g59) & (!g64) & (!g60)) + ((!f) & (!h) & (g) & (!g59) & (!g64) & (g60)) + ((!f) & (h) & (!g) & (!g59) & (g64) & (!g60)));
	assign g278 = (((n) & (!g65) & (!sk[34]) & (!g146) & (!g276) & (!g277)) + ((!n) & (!g65) & (!sk[34]) & (g146) & (!g276) & (!g277)) + ((!n) & (!g65) & (!sk[34]) & (!g146) & (!g276) & (g277)) + ((!n) & (g65) & (!sk[34]) & (g146) & (!g276) & (!g277)) + ((!n) & (!g65) & (sk[34]) & (!g146) & (g276) & (!g277)));
	assign g279 = (((!sk[35]) & (!g275) & (g278)) + ((sk[35]) & (!g275) & (!g278)));
	assign g280 = (((!g54) & (g75) & (!sk[36]) & (!g114)) + ((g54) & (g75) & (!sk[36]) & (g114)));
	assign g281 = (((!sk[37]) & (!d) & (c)) + ((sk[37]) & (!d) & (!c)));
	assign g282 = (((!sk[38]) & (!e) & (!l) & (g9) & (!g281)) + ((!sk[38]) & (!e) & (!l) & (!g9) & (g281)) + ((!sk[38]) & (e) & (l) & (g9) & (g281)));
	assign g283 = (((!g40) & (!sk[39]) & (!k) & (g86) & (!g282)) + ((!g40) & (!sk[39]) & (!k) & (!g86) & (g282)) + ((g40) & (!sk[39]) & (!k) & (g86) & (g282)));
	assign g284 = (((h) & (!n) & (!sk[40]) & (!g65) & (!g87) & (!g147)) + ((!h) & (!n) & (!sk[40]) & (g65) & (!g87) & (!g147)) + ((!h) & (!n) & (!sk[40]) & (!g65) & (!g87) & (g147)) + ((!h) & (!n) & (!sk[40]) & (!g65) & (g87) & (g147)) + ((h) & (!n) & (!sk[40]) & (g65) & (!g87) & (g147)));
	assign g285 = (((j) & (!g71) & (!g147) & (!g166) & (!sk[41]) & (!g284)) + ((!j) & (!g71) & (g147) & (!g166) & (!sk[41]) & (!g284)) + ((!j) & (!g71) & (!g147) & (!g166) & (!sk[41]) & (g284)) + ((j) & (!g71) & (!g147) & (!g166) & (!sk[41]) & (!g284)) + ((!j) & (!g71) & (!g147) & (!g166) & (sk[41]) & (!g284)) + ((!j) & (!g71) & (!g147) & (!g166) & (sk[41]) & (!g284)));
	assign g286 = (((g245) & (!g267) & (!g280) & (!g283) & (!sk[42]) & (!g285)) + ((!g245) & (!g267) & (g280) & (!g283) & (!sk[42]) & (!g285)) + ((!g245) & (!g267) & (!g280) & (!g283) & (!sk[42]) & (g285)) + ((!g245) & (!g267) & (!g280) & (!g283) & (!sk[42]) & (g285)));
	assign g287 = (((!d) & (!f) & (!a) & (g35) & (g80) & (!g115)) + ((!d) & (f) & (!a) & (g35) & (!g80) & (g115)));
	assign g288 = (((!g81) & (!g68) & (g156) & (!sk[44]) & (!g472)) + ((!g81) & (!g68) & (!g156) & (!sk[44]) & (g472)) + ((g81) & (!g68) & (!g156) & (!sk[44]) & (g472)) + ((!g81) & (!g68) & (!g156) & (!sk[44]) & (g472)));
	assign g289 = (((!sk[45]) & (!h) & (!g) & (i) & (!g9)) + ((!sk[45]) & (!h) & (!g) & (!i) & (g9)) + ((!sk[45]) & (!h) & (!g) & (!i) & (g9)));
	assign g290 = (((!g135) & (!sk[46]) & (g202)) + ((g135) & (sk[46]) & (!g202)));
	assign g291 = (((k) & (!l) & (!sk[47]) & (!g9) & (!g289) & (!g290)) + ((!k) & (!l) & (!sk[47]) & (g9) & (!g289) & (!g290)) + ((!k) & (!l) & (!sk[47]) & (!g9) & (!g289) & (g290)) + ((!k) & (!l) & (!sk[47]) & (g9) & (!g289) & (g290)) + ((!k) & (!l) & (sk[47]) & (!g9) & (g289) & (!g290)));
	assign g292 = (((!sk[48]) & (!f) & (g281) & (!g291)) + ((!sk[48]) & (!f) & (g281) & (g291)));
	assign g293 = (((!k) & (!sk[49]) & (!g41) & (g58) & (!g282)) + ((!k) & (!sk[49]) & (!g41) & (!g58) & (g282)) + ((k) & (!sk[49]) & (g41) & (g58) & (g282)));
	assign g294 = (((a) & (!g97) & (!sk[50]) & (!g85) & (!g292) & (!g293)) + ((!a) & (!g97) & (!sk[50]) & (g85) & (!g292) & (!g293)) + ((!a) & (!g97) & (!sk[50]) & (!g85) & (!g292) & (g293)) + ((!a) & (!g97) & (sk[50]) & (!g85) & (!g292) & (!g293)) + ((!a) & (!g97) & (sk[50]) & (!g85) & (!g292) & (!g293)) + ((!a) & (!g97) & (sk[50]) & (!g85) & (!g292) & (!g293)));
	assign g295 = (((!g155) & (!g279) & (g286) & (!g287) & (g288) & (g294)) + ((!g155) & (g279) & (g286) & (!g287) & (g288) & (g294)));
	assign g296 = (((d) & (!e) & (!sk[52]) & (!a) & (!g275) & (!g278)) + ((!d) & (!e) & (!sk[52]) & (a) & (!g275) & (!g278)) + ((!d) & (!e) & (!sk[52]) & (!a) & (!g275) & (g278)) + ((!d) & (e) & (!sk[52]) & (a) & (g275) & (!g278)) + ((!d) & (e) & (!sk[52]) & (a) & (!g275) & (g278)));
	assign g297 = (((h) & (!g) & (!i) & (!g1) & (!sk[53]) & (!c)) + ((!h) & (!g) & (i) & (!g1) & (!sk[53]) & (!c)) + ((!h) & (!g) & (!i) & (!g1) & (!sk[53]) & (c)) + ((!h) & (!g) & (i) & (g1) & (!sk[53]) & (c)));
	assign g298 = (((!sk[54]) & (j) & (!k) & (!l) & (!g105) & (!g297)) + ((!sk[54]) & (!j) & (!k) & (l) & (!g105) & (!g297)) + ((!sk[54]) & (!j) & (!k) & (!l) & (!g105) & (g297)) + ((!sk[54]) & (j) & (!k) & (!l) & (!g105) & (!g297)) + ((sk[54]) & (!j) & (!k) & (!l) & (!g105) & (!g297)) + ((!sk[54]) & (!j) & (!k) & (!l) & (!g105) & (g297)));
	assign g299 = (((f) & (!g) & (!g47) & (!sk[55]) & (!g48) & (!g81)) + ((!f) & (!g) & (g47) & (!sk[55]) & (!g48) & (!g81)) + ((!f) & (!g) & (!g47) & (!sk[55]) & (!g48) & (g81)) + ((!f) & (!g) & (g47) & (!sk[55]) & (!g48) & (!g81)) + ((!f) & (g) & (!g47) & (sk[55]) & (g48) & (!g81)));
	assign g300 = (((!sk[56]) & (b) & (!d) & (!e) & (!g298) & (!g299)) + ((!sk[56]) & (!b) & (!d) & (e) & (!g298) & (!g299)) + ((!sk[56]) & (!b) & (!d) & (!e) & (!g298) & (g299)) + ((!sk[56]) & (!b) & (!d) & (e) & (!g298) & (g299)) + ((!sk[56]) & (b) & (d) & (e) & (!g298) & (!g299)));
	assign g301 = (((!b) & (!sk[57]) & (!d) & (f) & (!g7)) + ((!b) & (!sk[57]) & (!d) & (!f) & (g7)) + ((b) & (!sk[57]) & (d) & (f) & (g7)));
	assign g302 = (((!sk[58]) & (b) & (!g33) & (!g34) & (!g97) & (!g104)) + ((!sk[58]) & (!b) & (!g33) & (g34) & (!g97) & (!g104)) + ((!sk[58]) & (!b) & (!g33) & (!g34) & (!g97) & (g104)) + ((!sk[58]) & (!b) & (!g33) & (g34) & (g97) & (!g104)) + ((sk[58]) & (!b) & (!g33) & (!g34) & (g97) & (!g104)));
	assign g303 = (((!sk[59]) & (!e) & (!l) & (g9) & (!g97)) + ((!sk[59]) & (!e) & (!l) & (!g9) & (g97)) + ((!sk[59]) & (!e) & (l) & (g9) & (g97)));
	assign g304 = (((f) & (!h) & (!g) & (!k) & (!sk[60]) & (!g58)) + ((!f) & (!h) & (g) & (!k) & (!sk[60]) & (!g58)) + ((!f) & (!h) & (!g) & (!k) & (!sk[60]) & (g58)) + ((!f) & (!h) & (g) & (k) & (!sk[60]) & (g58)));
	assign g305 = (((!sk[61]) & (!h) & (!g58) & (g34) & (!g258)) + ((!sk[61]) & (!h) & (!g58) & (!g34) & (g258)) + ((!sk[61]) & (!h) & (g58) & (g34) & (g258)));
	assign g306 = (((!f) & (!g90) & (g303) & (g304) & (!sk[62]) & (!g305)) + ((f) & (!g90) & (!g303) & (!g304) & (!sk[62]) & (!g305)) + ((!f) & (!g90) & (g303) & (!g304) & (!sk[62]) & (!g305)) + ((!f) & (!g90) & (!g303) & (!g304) & (!sk[62]) & (g305)) + ((!f) & (g90) & (!g303) & (!g304) & (!sk[62]) & (g305)));
	assign g307 = (((d) & (!e) & (!l) & (!g9) & (!sk[63]) & (!c)) + ((!d) & (!e) & (l) & (!g9) & (!sk[63]) & (!c)) + ((!d) & (!e) & (!l) & (!g9) & (!sk[63]) & (c)) + ((d) & (e) & (l) & (g9) & (!sk[63]) & (!c)));
	assign g308 = (((!sk[64]) & (b) & (!f) & (!n) & (!g76) & (!g97)) + ((!sk[64]) & (!b) & (!f) & (n) & (!g76) & (!g97)) + ((!sk[64]) & (!b) & (!f) & (!n) & (!g76) & (g97)) + ((!sk[64]) & (!b) & (!f) & (n) & (g76) & (g97)));
	assign g309 = (((!h) & (!g58) & (!g258) & (g304) & (g307) & (!g308)) + ((!h) & (g58) & (g258) & (!g304) & (!g307) & (g308)));
	assign g310 = (((!sk[66]) & (!k) & (g86) & (!g146)) + ((!sk[66]) & (!k) & (g86) & (g146)));
	assign g311 = (((!sk[67]) & (!h) & (g86) & (!g262)) + ((!sk[67]) & (h) & (g86) & (g262)));
	assign g312 = (((!f) & (!g34) & (!g90) & (g303) & (g310) & (!g311)) + ((!f) & (g34) & (g90) & (!g303) & (!g310) & (g311)));
	assign g313 = (((!sk[69]) & (!i) & (g9) & (!g281)) + ((!sk[69]) & (!i) & (g9) & (g281)));
	assign g314 = (((!sk[70]) & (!e) & (!f) & (h) & (!g)) + ((!sk[70]) & (!e) & (!f) & (!h) & (g)) + ((sk[70]) & (!e) & (!f) & (!h) & (!g)));
	assign g315 = (((!k) & (!l) & (g313) & (!sk[71]) & (!g314)) + ((!k) & (!l) & (!g313) & (!sk[71]) & (g314)) + ((!k) & (!l) & (g313) & (!sk[71]) & (g314)));
	assign g316 = (((!sk[72]) & (g46) & (!g19) & (!g158) & (!g312) & (!g315)) + ((!sk[72]) & (!g46) & (!g19) & (g158) & (!g312) & (!g315)) + ((!sk[72]) & (!g46) & (!g19) & (!g158) & (!g312) & (g315)) + ((sk[72]) & (!g46) & (!g19) & (!g158) & (!g312) & (!g315)));
	assign g317 = (((!k) & (!l) & (!sk[73]) & (g9) & (!g99)) + ((!k) & (!l) & (!sk[73]) & (!g9) & (g99)) + ((k) & (l) & (!sk[73]) & (g9) & (g99)));
	assign g318 = (((!g) & (!sk[74]) & (!g23) & (g281) & (!g317)) + ((!g) & (!sk[74]) & (!g23) & (!g281) & (g317)) + ((!g) & (!sk[74]) & (g23) & (g281) & (g317)));
	assign g319 = (((!f) & (!sk[75]) & (g76) & (!g90)) + ((f) & (!sk[75]) & (g76) & (g90)));
	assign g320 = (((k) & (!sk[76]) & (!l) & (!g41) & (!g58) & (!g20)) + ((!k) & (!sk[76]) & (!l) & (g41) & (!g58) & (!g20)) + ((!k) & (!sk[76]) & (!l) & (!g41) & (!g58) & (g20)) + ((!k) & (!sk[76]) & (!l) & (g41) & (g58) & (g20)));
	assign g321 = (((!h) & (!k) & (l) & (!sk[77]) & (!g58)) + ((!h) & (!k) & (!l) & (!sk[77]) & (g58)) + ((!h) & (!k) & (!l) & (!sk[77]) & (g58)));
	assign g322 = (((n) & (!sk[78]) & (!m) & (!g319) & (!g320) & (!g321)) + ((!n) & (!sk[78]) & (!m) & (g319) & (!g320) & (!g321)) + ((!n) & (!sk[78]) & (!m) & (!g319) & (!g320) & (g321)) + ((!n) & (!sk[78]) & (!m) & (g319) & (!g320) & (g321)) + ((!n) & (sk[78]) & (!m) & (!g319) & (g320) & (!g321)));
	assign g323 = (((!g31) & (g90) & (!sk[79]) & (!g75)) + ((g31) & (g90) & (!sk[79]) & (g75)));
	assign g324 = (((!sk[80]) & (!b) & (!d) & (c) & (!a)) + ((!sk[80]) & (!b) & (!d) & (!c) & (a)) + ((!sk[80]) & (!b) & (!d) & (c) & (a)) + ((!sk[80]) & (!b) & (d) & (!c) & (a)));
	assign g325 = (((!d) & (!e) & (f) & (g113) & (g115) & (!g324)) + ((!d) & (e) & (f) & (!g113) & (g115) & (g324)));
	assign g326 = (((e) & (!sk[82]) & (!g318) & (!g322) & (!g323) & (!g325)) + ((!e) & (!sk[82]) & (!g318) & (g322) & (!g323) & (!g325)) + ((!e) & (!sk[82]) & (!g318) & (!g322) & (!g323) & (g325)) + ((e) & (!sk[82]) & (!g318) & (!g322) & (!g323) & (!g325)) + ((!e) & (sk[82]) & (!g318) & (!g322) & (!g323) & (!g325)));
	assign g327 = (((!g37) & (!g123) & (!g306) & (!g309) & (g316) & (g326)) + ((!g37) & (g123) & (!g306) & (!g309) & (g316) & (g326)));
	assign g328 = (((!g296) & (!g300) & (g286) & (!g301) & (!g302) & (g327)));
	assign g329 = (((g310) & (!sk[85]) & (!g311) & (g307) & (!g308)) + ((!g310) & (!sk[85]) & (!g311) & (g307) & (!g308)) + ((!g310) & (!sk[85]) & (!g311) & (!g307) & (g308)) + ((!g310) & (!sk[85]) & (g311) & (!g307) & (g308)));
	assign g330 = (((!j) & (!sk[86]) & (k)) + ((!j) & (sk[86]) & (!k)));
	assign g331 = (((d) & (!sk[87]) & (!e) & (!f) & (!a) & (!g35)) + ((!d) & (!sk[87]) & (!e) & (f) & (!a) & (!g35)) + ((!d) & (!sk[87]) & (!e) & (!f) & (!a) & (g35)) + ((d) & (!sk[87]) & (!e) & (f) & (!a) & (g35)));
	assign g332 = (((!l) & (!g15) & (!g330) & (!g136) & (!g293) & (!g331)) + ((!l) & (!g15) & (!g330) & (!g136) & (!g293) & (!g331)) + ((!l) & (!g15) & (!g330) & (!g136) & (!g293) & (!g331)) + ((!l) & (!g15) & (!g330) & (!g136) & (!g293) & (!g331)) + ((!l) & (!g15) & (!g330) & (!g136) & (!g293) & (!g331)));
	assign g333 = (((!j) & (!sk[89]) & (!g10) & (g262) & (!g308)) + ((!j) & (!sk[89]) & (!g10) & (!g262) & (g308)) + ((j) & (!sk[89]) & (g10) & (g262) & (g308)));
	assign g334 = (((f) & (!sk[90]) & (!h) & (!g) & (!k) & (!g99)) + ((!f) & (!sk[90]) & (!h) & (g) & (!k) & (!g99)) + ((!f) & (!sk[90]) & (!h) & (!g) & (!k) & (g99)) + ((!f) & (!sk[90]) & (!h) & (g) & (!k) & (g99)));
	assign g335 = (((g145) & (!l) & (!g15) & (!g135) & (!sk[91]) & (!g331)) + ((!g145) & (!l) & (g15) & (!g135) & (!sk[91]) & (!g331)) + ((!g145) & (!l) & (!g15) & (!g135) & (!sk[91]) & (g331)) + ((g145) & (l) & (g15) & (g135) & (!sk[91]) & (g331)));
	assign g336 = (((g306) & (!g307) & (!sk[92]) & (!g333) & (!g334) & (!g335)) + ((!g306) & (!g307) & (!sk[92]) & (g333) & (!g334) & (!g335)) + ((!g306) & (!g307) & (!sk[92]) & (!g333) & (!g334) & (g335)) + ((!g306) & (!g307) & (sk[92]) & (!g333) & (!g334) & (!g335)) + ((!g306) & (!g307) & (sk[92]) & (!g333) & (!g334) & (!g335)));
	assign g337 = (((!sk[93]) & (!f) & (!l) & (g330) & (!g281)) + ((!sk[93]) & (!f) & (!l) & (!g330) & (g281)) + ((!sk[93]) & (!f) & (!l) & (g330) & (g281)));
	assign g338 = (((!e) & (!sk[94]) & (!g289) & (g318) & (!g337)) + ((!e) & (!sk[94]) & (!g289) & (g318) & (!g337)) + ((!e) & (!sk[94]) & (!g289) & (!g318) & (g337)) + ((!e) & (!sk[94]) & (g289) & (!g318) & (g337)));
	assign g339 = (((g312) & (!g329) & (!g332) & (!g336) & (!sk[95]) & (!g338)) + ((!g312) & (!g329) & (g332) & (!g336) & (!sk[95]) & (!g338)) + ((!g312) & (!g329) & (!g332) & (!g336) & (!sk[95]) & (g338)) + ((!g312) & (!g329) & (g332) & (g336) & (!sk[95]) & (!g338)));
	assign g340 = (((!a) & (!sk[96]) & (g35) & (!g82)) + ((a) & (!sk[96]) & (g35) & (g82)));
	assign g341 = (((!g136) & (g203) & (!sk[97]) & (!g340)) + ((g136) & (g203) & (!sk[97]) & (g340)));
	assign g342 = (((!g182) & (g258) & (!sk[98]) & (!g319)) + ((g182) & (g258) & (!sk[98]) & (g319)));
	assign g343 = (((g40) & (!g20) & (!g317) & (!sk[99]) & (!g309) & (!g342)) + ((!g40) & (!g20) & (g317) & (!sk[99]) & (!g309) & (!g342)) + ((!g40) & (!g20) & (!g317) & (!sk[99]) & (!g309) & (g342)) + ((!g40) & (!g20) & (!g317) & (sk[99]) & (!g309) & (!g342)) + ((!g40) & (!g20) & (!g317) & (sk[99]) & (!g309) & (!g342)) + ((!g40) & (!g20) & (!g317) & (sk[99]) & (!g309) & (!g342)));
	assign g344 = (((g312) & (!sk[100]) & (!g329) & (!g332) & (!g341) & (!g343)) + ((!g312) & (!sk[100]) & (!g329) & (g332) & (!g341) & (!g343)) + ((!g312) & (!sk[100]) & (!g329) & (!g332) & (!g341) & (g343)) + ((!g312) & (!sk[100]) & (!g329) & (g332) & (!g341) & (g343)));
	assign g345 = (((!e) & (!g318) & (g315) & (!sk[101]) & (!g344)) + ((!e) & (!g318) & (!g315) & (!sk[101]) & (g344)) + ((!e) & (!g318) & (!g315) & (!sk[101]) & (g344)) + ((!e) & (!g318) & (!g315) & (!sk[101]) & (g344)));
	assign g346 = (((h) & (g) & (!sk[102]) & (!a) & (!g36) & (!g223)) + ((h) & (!g) & (!sk[102]) & (!a) & (!g36) & (!g223)) + ((!h) & (g) & (!sk[102]) & (a) & (!g36) & (!g223)) + ((!h) & (!g) & (!sk[102]) & (a) & (!g36) & (!g223)) + ((!h) & (!g) & (!sk[102]) & (!a) & (!g36) & (g223)) + ((!h) & (g) & (sk[102]) & (!a) & (!g36) & (!g223)) + ((!h) & (g) & (!sk[102]) & (!a) & (!g36) & (g223)));
	assign g347 = (((b) & (!h) & (!sk[103]) & (!n) & (!k) & (!g97)) + ((!b) & (!h) & (!sk[103]) & (n) & (!k) & (!g97)) + ((!b) & (!h) & (!sk[103]) & (!n) & (!k) & (g97)) + ((!b) & (h) & (!sk[103]) & (!n) & (!k) & (g97)) + ((!b) & (h) & (!sk[103]) & (!n) & (!k) & (g97)));
	assign g348 = (((!g) & (!m) & (l) & (!sk[104]) & (!g347)) + ((!g) & (!m) & (!l) & (!sk[104]) & (g347)) + ((!g) & (m) & (!l) & (sk[104]) & (!g347)) + ((!g) & (!m) & (!l) & (sk[104]) & (!g347)) + ((!g) & (!m) & (!l) & (sk[104]) & (!g347)));
	assign g349 = (((!e) & (!f) & (j) & (!sk[105]) & (!i)) + ((!e) & (!f) & (!j) & (!sk[105]) & (i)) + ((!e) & (!f) & (!j) & (sk[105]) & (!i)));
	assign g350 = (((g322) & (!g346) & (!g348) & (!sk[106]) & (!g283) & (!g349)) + ((!g322) & (!g346) & (g348) & (!sk[106]) & (!g283) & (!g349)) + ((!g322) & (!g346) & (!g348) & (!sk[106]) & (!g283) & (g349)) + ((!g322) & (!g346) & (g348) & (!sk[106]) & (!g283) & (!g349)) + ((!g322) & (!g346) & (!g348) & (sk[106]) & (!g283) & (!g349)) + ((!g322) & (g346) & (!g348) & (!sk[106]) & (!g283) & (g349)));
	assign g351 = (((!g292) & (!g336) & (g344) & (!sk[107]) & (!g350)) + ((!g292) & (!g336) & (!g344) & (!sk[107]) & (g350)) + ((!g292) & (g336) & (g344) & (!sk[107]) & (g350)));
	assign g352 = (((h) & (!k) & (!l) & (!g9) & (!sk[108]) & (!g99)) + ((!h) & (!k) & (l) & (!g9) & (!sk[108]) & (!g99)) + ((!h) & (!k) & (!l) & (!g9) & (!sk[108]) & (g99)) + ((!h) & (!k) & (!l) & (g9) & (!sk[108]) & (g99)) + ((h) & (k) & (l) & (g9) & (!sk[108]) & (g99)));
	assign g353 = (((!h) & (!j) & (!sk[109]) & (k) & (!i)) + ((!h) & (!j) & (!sk[109]) & (!k) & (i)) + ((h) & (!j) & (!sk[109]) & (!k) & (i)));
	assign g354 = (((g15) & (!sk[110]) & (g353)) + ((!g15) & (!sk[110]) & (g353)));
	assign g355 = (((!e) & (!g) & (g1) & (!sk[111]) & (!g281)) + ((!e) & (!g) & (!g1) & (!sk[111]) & (g281)) + ((e) & (g) & (!g1) & (sk[111]) & (!g281)) + ((!e) & (g) & (!g1) & (sk[111]) & (!g281)) + ((!e) & (g) & (!g1) & (sk[111]) & (!g281)));
	assign g356 = (((e) & (!sk[112]) & (!h) & (!m) & (!i) & (!c)) + ((!e) & (!sk[112]) & (!h) & (m) & (!i) & (!c)) + ((!e) & (!sk[112]) & (!h) & (!m) & (!i) & (c)) + ((!e) & (sk[112]) & (!h) & (!m) & (!i) & (!c)));
	assign g357 = (((!sk[113]) & (b) & (!e) & (!h) & (!i) & (!g1)) + ((!sk[113]) & (!b) & (!e) & (h) & (!i) & (!g1)) + ((!sk[113]) & (!b) & (!e) & (!h) & (!i) & (g1)) + ((!sk[113]) & (!b) & (!e) & (!h) & (!i) & (g1)));
	assign g358 = (((g35) & (!g182) & (!g223) & (!sk[114]) & (!g356) & (!g357)) + ((!g35) & (!g182) & (g223) & (!sk[114]) & (!g356) & (!g357)) + ((!g35) & (!g182) & (!g223) & (!sk[114]) & (!g356) & (g357)) + ((g35) & (!g182) & (!g223) & (!sk[114]) & (!g356) & (!g357)) + ((!g35) & (!g182) & (!g223) & (sk[114]) & (!g356) & (!g357)) + ((!g35) & (!g182) & (!g223) & (sk[114]) & (!g356) & (!g357)));
	assign g359 = (((!f) & (!sk[115]) & (!g313) & (g355) & (!g358)) + ((!f) & (!sk[115]) & (!g313) & (!g355) & (g358)) + ((f) & (!sk[115]) & (!g313) & (g355) & (g358)) + ((!f) & (!sk[115]) & (!g313) & (g355) & (g358)));
	assign g360 = (((d) & (!a) & (!g35) & (!g352) & (!g354) & (g359)) + ((!d) & (!a) & (!g35) & (!g352) & (!g354) & (g359)) + ((d) & (!a) & (g35) & (!g352) & (!g354) & (g359)));
	assign g361 = (((!e) & (!sk[117]) & (f) & (!c)) + ((!e) & (sk[117]) & (!f) & (c)));
	assign g362 = (((e) & (!f) & (g145) & (!a) & (g15) & (!g90)) + ((!e) & (!f) & (g145) & (!a) & (g15) & (!g90)) + ((!e) & (!f) & (g145) & (a) & (g15) & (!g90)) + ((!e) & (!f) & (g145) & (!a) & (g15) & (!g90)));
	assign g363 = (((!sk[119]) & (!g9) & (c)) + ((!sk[119]) & (g9) & (c)));
	assign g364 = (((h) & (!i) & (!sk[120]) & (!g281) & (!g317) & (!g363)) + ((!h) & (!i) & (!sk[120]) & (g281) & (!g317) & (!g363)) + ((!h) & (!i) & (!sk[120]) & (!g281) & (!g317) & (g363)) + ((h) & (!i) & (!sk[120]) & (!g281) & (g317) & (!g363)) + ((!h) & (!i) & (!sk[120]) & (!g281) & (!g317) & (g363)));
	assign g365 = (((h) & (!g) & (!g54) & (!g362) & (!sk[121]) & (!g364)) + ((!h) & (!g) & (g54) & (!g362) & (!sk[121]) & (!g364)) + ((!h) & (!g) & (!g54) & (!g362) & (!sk[121]) & (g364)) + ((h) & (!g) & (!g54) & (!g362) & (!sk[121]) & (!g364)) + ((!h) & (!g) & (!g54) & (!g362) & (sk[121]) & (!g364)));
	assign g366 = (((i) & (!g9) & (!sk[122]) & (!g330) & (!g361) & (!g365)) + ((!i) & (!g9) & (!sk[122]) & (g330) & (!g361) & (!g365)) + ((!i) & (!g9) & (!sk[122]) & (!g330) & (!g361) & (g365)) + ((!i) & (!g9) & (!sk[122]) & (!g330) & (!g361) & (g365)) + ((!i) & (!g9) & (!sk[122]) & (!g330) & (!g361) & (g365)) + ((!i) & (!g9) & (!sk[122]) & (g330) & (!g361) & (g365)));
	assign g367 = (((b) & (!d) & (e) & (!l) & (!c) & (!g330)) + ((b) & (!d) & (e) & (!l) & (c) & (!g330)) + ((!b) & (!d) & (e) & (l) & (!c) & (g330)) + ((!b) & (!d) & (!e) & (l) & (c) & (g330)));
	assign g368 = (((!sk[124]) & (!e) & (c) & (!g90)) + ((!sk[124]) & (!e) & (c) & (g90)));
	assign g369 = (((!b) & (h) & (j) & (!k) & (!i) & (g368)) + ((!b) & (!h) & (!j) & (!k) & (!i) & (g368)) + ((b) & (!h) & (j) & (!k) & (i) & (!g368)) + ((!b) & (!h) & (!j) & (k) & (!i) & (g368)) + ((!b) & (!h) & (j) & (!k) & (i) & (g368)));
	assign g370 = (((!g) & (!g1) & (g367) & (!sk[126]) & (!g369)) + ((!g) & (g1) & (!g367) & (!sk[126]) & (g369)) + ((!g) & (!g1) & (!g367) & (!sk[126]) & (g369)) + ((!g) & (g1) & (!g367) & (sk[126]) & (!g369)));
	assign g371 = (((!d) & (!a) & (!sk[127]) & (g15) & (!g212)) + ((!d) & (!a) & (!sk[127]) & (!g15) & (g212)) + ((d) & (!a) & (!sk[127]) & (g15) & (g212)) + ((!d) & (a) & (!sk[127]) & (g15) & (g212)));
	assign g372 = (((!i) & (!l) & (!sk[0]) & (g1) & (!g371)) + ((!i) & (!l) & (!sk[0]) & (!g1) & (g371)) + ((!i) & (!l) & (sk[0]) & (!g1) & (!g371)) + ((i) & (!l) & (!sk[0]) & (g1) & (!g371)) + ((!i) & (l) & (!sk[0]) & (g1) & (!g371)));
	assign g373 = (((!sk[1]) & (!b) & (!h) & (k) & (!i)) + ((!sk[1]) & (!b) & (!h) & (!k) & (i)) + ((sk[1]) & (!b) & (!h) & (!k) & (!i)) + ((sk[1]) & (b) & (!h) & (!k) & (!i)));
	assign g374 = (((e) & (!g1) & (!c) & (!sk[2]) & (!g352) & (!g373)) + ((!e) & (!g1) & (c) & (!sk[2]) & (!g352) & (!g373)) + ((!e) & (!g1) & (c) & (!sk[2]) & (g352) & (!g373)) + ((!e) & (!g1) & (!c) & (!sk[2]) & (!g352) & (g373)) + ((e) & (g1) & (!c) & (!sk[2]) & (!g352) & (g373)));
	assign g375 = (((!sk[3]) & (f) & (!h) & (!g370) & (!g372) & (!g374)) + ((!sk[3]) & (!f) & (!h) & (g370) & (!g372) & (!g374)) + ((!sk[3]) & (!f) & (!h) & (!g370) & (!g372) & (g374)) + ((sk[3]) & (!f) & (!h) & (!g370) & (!g372) & (!g374)));
	assign g376 = (((!b) & (!k) & (!sk[4]) & (l) & (!g1)) + ((!b) & (!k) & (!sk[4]) & (!l) & (g1)) + ((!b) & (k) & (!sk[4]) & (!l) & (g1)) + ((!b) & (!k) & (!sk[4]) & (!l) & (g1)) + ((!b) & (!k) & (!sk[4]) & (l) & (g1)));
	assign g377 = (((h) & (!sk[5]) & (!n) & (!i) & (!g64) & (!g376)) + ((!h) & (!sk[5]) & (!n) & (i) & (!g64) & (!g376)) + ((!h) & (!sk[5]) & (!n) & (!i) & (!g64) & (g376)) + ((!h) & (sk[5]) & (!n) & (!i) & (g64) & (!g376)));
	assign g378 = (((e) & (!g) & (!n) & (!m) & (g281) & (!g353)) + ((!e) & (!g) & (!n) & (!m) & (g281) & (!g353)) + ((!e) & (!g) & (!n) & (!m) & (!g281) & (g353)));
	assign g379 = (((d) & (!e) & (!sk[7]) & (!h) & (!k) & (!a)) + ((!d) & (!e) & (!sk[7]) & (h) & (!k) & (!a)) + ((!d) & (!e) & (!sk[7]) & (!h) & (!k) & (a)) + ((d) & (!e) & (!sk[7]) & (!h) & (!k) & (!a)) + ((d) & (!e) & (!sk[7]) & (!h) & (k) & (!a)));
	assign g380 = (((!sk[8]) & (d) & (!e) & (!i) & (!a) & (!g35)) + ((!sk[8]) & (!d) & (!e) & (i) & (!a) & (!g35)) + ((!sk[8]) & (!d) & (!e) & (!i) & (!a) & (g35)) + ((!sk[8]) & (d) & (!e) & (!i) & (!a) & (!g35)) + ((!sk[8]) & (!d) & (!e) & (!i) & (a) & (g35)));
	assign g381 = (((b) & (!g15) & (!g281) & (!sk[9]) & (!g379) & (!g380)) + ((!b) & (!g15) & (g281) & (!sk[9]) & (!g379) & (!g380)) + ((!b) & (g15) & (!g281) & (!sk[9]) & (!g379) & (g380)) + ((!b) & (!g15) & (!g281) & (!sk[9]) & (!g379) & (g380)) + ((!b) & (g15) & (g281) & (!sk[9]) & (!g379) & (!g380)) + ((!b) & (g15) & (!g281) & (sk[9]) & (g379) & (!g380)));
	assign g382 = (((!k) & (!l) & (!sk[10]) & (!g182) & (!g462) & (g381)) + ((k) & (!l) & (!sk[10]) & (!g182) & (!g462) & (!g381)) + ((!k) & (!l) & (sk[10]) & (!g182) & (!g462) & (!g381)) + ((!k) & (!l) & (!sk[10]) & (g182) & (!g462) & (!g381)) + ((!k) & (!l) & (sk[10]) & (!g182) & (!g462) & (!g381)) + ((!k) & (!l) & (!sk[10]) & (g182) & (!g462) & (!g381)));
	assign g383 = (((!sk[11]) & (!h) & (!k) & (g34) & (!g99)) + ((!sk[11]) & (!h) & (!k) & (!g34) & (g99)) + ((!sk[11]) & (!h) & (!k) & (g34) & (g99)));
	assign g384 = (((!sk[12]) & (!g57) & (g20)) + ((!sk[12]) & (g57) & (g20)));
	assign g385 = (((j) & (!k) & (!sk[13]) & (!i) & (!l) & (!g384)) + ((!j) & (!k) & (!sk[13]) & (i) & (!l) & (!g384)) + ((!j) & (!k) & (!sk[13]) & (!i) & (!l) & (g384)) + ((!j) & (!k) & (!sk[13]) & (!i) & (l) & (g384)) + ((!j) & (!k) & (!sk[13]) & (i) & (!l) & (g384)) + ((!j) & (!k) & (!sk[13]) & (!i) & (l) & (g384)) + ((!j) & (k) & (!sk[13]) & (!i) & (!l) & (g384)));
	assign g386 = (((g) & (!l) & (!g211) & (!sk[14]) & (!g281) & (!g361)) + ((!g) & (!l) & (g211) & (!sk[14]) & (!g281) & (!g361)) + ((!g) & (!l) & (!g211) & (!sk[14]) & (!g281) & (g361)) + ((!g) & (!l) & (!g211) & (!sk[14]) & (!g281) & (g361)) + ((g) & (!l) & (!g211) & (!sk[14]) & (g281) & (!g361)));
	assign g387 = (((h) & (!g) & (!j) & (!k) & (!sk[15]) & (!i)) + ((!h) & (!g) & (j) & (!k) & (!sk[15]) & (!i)) + ((h) & (g) & (j) & (!k) & (!sk[15]) & (!i)) + ((!h) & (!g) & (!j) & (!k) & (!sk[15]) & (i)) + ((!h) & (g) & (!j) & (k) & (!sk[15]) & (i)));
	assign g388 = (((!e) & (f) & (!g) & (!j) & (!l) & (!c)) + ((!e) & (!f) & (g) & (!j) & (!l) & (!c)) + ((!e) & (!f) & (g) & (!j) & (!l) & (!c)));
	assign g389 = (((h) & (!sk[17]) & (!g40) & (!i) & (!g20) & (!g388)) + ((!h) & (!sk[17]) & (!g40) & (i) & (!g20) & (!g388)) + ((!h) & (!sk[17]) & (!g40) & (!i) & (!g20) & (g388)) + ((!h) & (sk[17]) & (g40) & (!i) & (g20) & (!g388)));
	assign g390 = (((e) & (!f) & (!c) & (!sk[18]) & (!g387) & (!g389)) + ((!e) & (!f) & (c) & (!sk[18]) & (!g387) & (!g389)) + ((!e) & (!f) & (!c) & (!sk[18]) & (!g387) & (g389)) + ((e) & (!f) & (c) & (!sk[18]) & (!g387) & (!g389)) + ((!e) & (!f) & (!c) & (sk[18]) & (!g387) & (!g389)) + ((!e) & (f) & (!c) & (sk[18]) & (!g387) & (!g389)) + ((!e) & (!f) & (!c) & (sk[18]) & (!g387) & (!g389)));
	assign g391 = (((g9) & (g383) & (!sk[19]) & (!g385) & (!g386) & (!g390)) + ((g9) & (!g383) & (!sk[19]) & (g385) & (!g386) & (!g390)) + ((!g9) & (!g383) & (!sk[19]) & (g385) & (!g386) & (!g390)) + ((g9) & (!g383) & (!sk[19]) & (!g385) & (g386) & (!g390)) + ((!g9) & (!g383) & (!sk[19]) & (!g385) & (!g386) & (g390)) + ((g9) & (!g383) & (!sk[19]) & (!g385) & (!g386) & (!g390)));
	assign g392 = (((f) & (!g377) & (!g378) & (!sk[20]) & (!g382) & (!g391)) + ((!f) & (!g377) & (!g378) & (!sk[20]) & (!g382) & (g391)) + ((!f) & (!g377) & (!g378) & (sk[20]) & (!g382) & (!g391)) + ((!f) & (!g377) & (g378) & (!sk[20]) & (!g382) & (!g391)) + ((!f) & (!g377) & (!g378) & (sk[20]) & (g382) & (!g391)));
	assign g393 = (((!f) & (!m) & (!sk[21]) & (g145) & (!g10)) + ((!f) & (!m) & (!sk[21]) & (!g145) & (g10)) + ((f) & (!m) & (!sk[21]) & (g145) & (g10)));
	assign g394 = (((g) & (!sk[22]) & (!m) & (!j) & (!i) & (!l)) + ((!g) & (!sk[22]) & (!m) & (j) & (!i) & (!l)) + ((!g) & (!sk[22]) & (!m) & (!j) & (!i) & (l)) + ((g) & (!sk[22]) & (!m) & (!j) & (!i) & (!l)) + ((!g) & (sk[22]) & (!m) & (!j) & (i) & (!l)) + ((!g) & (sk[22]) & (!m) & (!j) & (i) & (!l)));
	assign g395 = (((!h) & (!sk[23]) & (!k) & (g393) & (!g394)) + ((!h) & (!sk[23]) & (!k) & (!g393) & (g394)) + ((!h) & (sk[23]) & (!k) & (!g393) & (!g394)) + ((!h) & (!sk[23]) & (!k) & (!g393) & (g394)) + ((!h) & (!sk[23]) & (k) & (!g393) & (g394)));
	assign g396 = (((d) & (!e) & (!l) & (!sk[24]) & (!g57) & (!g182)) + ((!d) & (!e) & (l) & (!sk[24]) & (!g57) & (!g182)) + ((!d) & (!e) & (!l) & (!sk[24]) & (!g57) & (g182)) + ((!d) & (!e) & (l) & (!sk[24]) & (g57) & (g182)) + ((!d) & (!e) & (l) & (!sk[24]) & (g57) & (g182)));
	assign g397 = (((m) & (!j) & (!sk[25]) & (!k) & (!g340) & (!g396)) + ((!m) & (!j) & (!sk[25]) & (k) & (!g340) & (!g396)) + ((!m) & (!j) & (!sk[25]) & (!k) & (!g340) & (g396)) + ((m) & (!j) & (!sk[25]) & (k) & (!g340) & (g396)) + ((m) & (!j) & (!sk[25]) & (k) & (g340) & (!g396)));
	assign g398 = (((!d) & (!f) & (!h) & (g) & (!k) & (!c)) + ((d) & (f) & (!h) & (!g) & (!k) & (!c)) + ((d) & (!f) & (!h) & (!g) & (!k) & (!c)) + ((!d) & (!f) & (!h) & (g) & (!k) & (!c)));
	assign g399 = (((e) & (!f) & (!sk[27]) & (!h) & (!g) & (!c)) + ((!e) & (!f) & (!sk[27]) & (h) & (!g) & (!c)) + ((!e) & (!f) & (!sk[27]) & (!h) & (!g) & (c)) + ((e) & (!f) & (!sk[27]) & (!h) & (!g) & (c)) + ((e) & (!f) & (!sk[27]) & (h) & (!g) & (!c)) + ((!e) & (!f) & (!sk[27]) & (h) & (!g) & (!c)));
	assign g400 = (((!sk[28]) & (!m) & (!i) & (g398) & (!g399)) + ((!sk[28]) & (!m) & (!i) & (!g398) & (g399)) + ((!sk[28]) & (!m) & (!i) & (g398) & (!g399)) + ((!sk[28]) & (!m) & (!i) & (!g398) & (g399)));
	assign g401 = (((!g44) & (!g) & (!sk[29]) & (m) & (!g330)) + ((!g44) & (!g) & (!sk[29]) & (!m) & (g330)) + ((g44) & (!g) & (!sk[29]) & (!m) & (g330)));
	assign g402 = (((!sk[30]) & (h) & (!j) & (!k) & (!i) & (!l)) + ((!sk[30]) & (!h) & (!j) & (k) & (!i) & (!l)) + ((!sk[30]) & (!h) & (!j) & (!k) & (!i) & (l)) + ((!sk[30]) & (h) & (j) & (!k) & (i) & (!l)) + ((sk[30]) & (!h) & (!j) & (!k) & (!i) & (!l)));
	assign g403 = (((f) & (!g) & (!sk[31]) & (!m) & (!c) & (!g402)) + ((!f) & (!g) & (!sk[31]) & (m) & (!c) & (!g402)) + ((!f) & (!g) & (!sk[31]) & (!m) & (!c) & (g402)) + ((!f) & (!g) & (sk[31]) & (!m) & (!c) & (!g402)));
	assign g404 = (((!sk[32]) & (!f) & (!m) & (g86) & (!g281)) + ((!sk[32]) & (!f) & (!m) & (!g86) & (g281)) + ((!sk[32]) & (!f) & (!m) & (g86) & (g281)));
	assign g405 = (((!sk[33]) & (g193) & (!g384) & (!g401) & (!g403) & (!g404)) + ((!sk[33]) & (!g193) & (!g384) & (g401) & (!g403) & (!g404)) + ((!sk[33]) & (!g193) & (!g384) & (!g401) & (!g403) & (g404)) + ((sk[33]) & (!g193) & (!g384) & (!g401) & (!g403) & (!g404)) + ((!sk[33]) & (g193) & (!g384) & (!g401) & (!g403) & (!g404)));
	assign g406 = (((!sk[34]) & (d) & (!e) & (!f) & (!a) & (!g35)) + ((!sk[34]) & (!d) & (!e) & (f) & (!a) & (!g35)) + ((!sk[34]) & (!d) & (!e) & (!f) & (!a) & (g35)) + ((!sk[34]) & (d) & (!e) & (!f) & (!a) & (!g35)) + ((sk[34]) & (!d) & (!e) & (!f) & (!a) & (!g35)) + ((!sk[34]) & (d) & (e) & (f) & (a) & (g35)));
	assign g407 = (((!sk[35]) & (!g) & (!m) & (g145) & (!g406)) + ((!sk[35]) & (!g) & (!m) & (!g145) & (g406)) + ((!sk[35]) & (!g) & (m) & (!g145) & (g406)));
	assign g408 = (((g395) & (!g397) & (!g400) & (!sk[36]) & (!g405) & (!g407)) + ((!g395) & (!g397) & (g400) & (!sk[36]) & (!g405) & (!g407)) + ((!g395) & (!g397) & (!g400) & (!sk[36]) & (!g405) & (g407)) + ((g395) & (!g397) & (!g400) & (!sk[36]) & (g405) & (!g407)));
	assign g409 = (((!d) & (!e) & (f) & (!sk[37]) & (!a)) + ((!d) & (!e) & (!f) & (!sk[37]) & (a)) + ((!d) & (!e) & (!f) & (sk[37]) & (!a)) + ((!d) & (!e) & (!f) & (!sk[37]) & (a)));
	assign g410 = (((!b) & (!sk[38]) & (e) & (!f)) + ((!b) & (!sk[38]) & (e) & (!f)));
	assign g411 = (((!sk[39]) & (!g1) & (g410)) + ((!sk[39]) & (g1) & (g410)));
	assign g412 = (((!b) & (!e) & (!j) & (!k) & (g1) & (!g97)) + ((b) & (e) & (!j) & (!k) & (g1) & (!g97)));
	assign g413 = (((j) & (!g15) & (!sk[41]) & (!g409) & (!g411) & (!g412)) + ((!j) & (!g15) & (!sk[41]) & (g409) & (!g411) & (!g412)) + ((!j) & (!g15) & (!sk[41]) & (!g409) & (!g411) & (g412)) + ((!j) & (!g15) & (sk[41]) & (!g409) & (!g411) & (!g412)) + ((!j) & (!g15) & (!sk[41]) & (g409) & (!g411) & (!g412)) + ((!j) & (!g15) & (sk[41]) & (!g409) & (!g411) & (!g412)) + ((!j) & (!g15) & (sk[41]) & (!g409) & (!g411) & (!g412)));
	assign g414 = (((!sk[42]) & (!d) & (e) & (!f)) + ((sk[42]) & (d) & (!e) & (!f)) + ((!sk[42]) & (d) & (e) & (f)));
	assign g415 = (((b) & (!e) & (!n) & (!sk[43]) & (!i) & (!c)) + ((!b) & (!e) & (n) & (!sk[43]) & (!i) & (!c)) + ((!b) & (!e) & (!n) & (!sk[43]) & (!i) & (c)) + ((!b) & (!e) & (n) & (!sk[43]) & (i) & (!c)) + ((!b) & (!e) & (!n) & (sk[43]) & (i) & (!c)));
	assign g416 = (((m) & (!sk[44]) & (!g330) & (!g414) & (!g363) & (!g415)) + ((!m) & (!sk[44]) & (!g330) & (g414) & (!g363) & (!g415)) + ((!m) & (!sk[44]) & (!g330) & (!g414) & (!g363) & (g415)) + ((!m) & (!sk[44]) & (g330) & (!g414) & (!g363) & (g415)) + ((!m) & (sk[44]) & (g330) & (!g414) & (g363) & (!g415)));
	assign g417 = (((n) & (!m) & (!j) & (!i) & (!g97) & (!g61)) + ((!n) & (!m) & (!j) & (!i) & (!g97) & (g61)));
	assign g418 = (((!h) & (!n) & (k) & (!sk[46]) & (!i) & (!l)) + ((h) & (!n) & (!k) & (!sk[46]) & (!i) & (!l)) + ((!h) & (!n) & (!k) & (!sk[46]) & (!i) & (l)) + ((!h) & (n) & (!k) & (sk[46]) & (!i) & (!l)) + ((!h) & (!n) & (!k) & (sk[46]) & (!i) & (!l)));
	assign g419 = (((d) & (!sk[47]) & (!j) & (!i) & (!g9) & (!c)) + ((!d) & (!sk[47]) & (!j) & (i) & (!g9) & (!c)) + ((!d) & (!sk[47]) & (!j) & (!i) & (!g9) & (c)) + ((!d) & (!sk[47]) & (!j) & (!i) & (g9) & (c)) + ((!d) & (!sk[47]) & (!j) & (i) & (g9) & (!c)));
	assign g420 = (((j) & (!g411) & (!g417) & (!sk[48]) & (!g418) & (!g419)) + ((!j) & (!g411) & (g417) & (!sk[48]) & (!g418) & (!g419)) + ((!j) & (!g411) & (!g417) & (!sk[48]) & (!g418) & (g419)) + ((j) & (!g411) & (!g417) & (!sk[48]) & (g418) & (!g419)) + ((!j) & (!g411) & (!g417) & (sk[48]) & (g418) & (!g419)));
	assign g421 = (((b) & (!e) & (!f) & (!g) & (!sk[49]) & (!g145)) + ((!b) & (!e) & (f) & (!g) & (!sk[49]) & (!g145)) + ((!b) & (!e) & (!f) & (!g) & (!sk[49]) & (g145)) + ((!b) & (!e) & (!f) & (g) & (!sk[49]) & (g145)) + ((!b) & (!e) & (!f) & (!g) & (sk[49]) & (!g145)));
	assign g422 = (((!g) & (!k) & (!l) & (g1) & (!g58) & (g421)) + ((!g) & (!k) & (!l) & (g1) & (!g58) & (!g421)) + ((!g) & (!k) & (!l) & (g1) & (!g58) & (!g421)));
	assign g423 = (((!h) & (!g313) & (!g413) & (!g416) & (g420) & (!g422)) + ((h) & (!g313) & (g413) & (!g416) & (!g420) & (!g422)));
	assign g424 = (((!b) & (!sk[52]) & (!d) & (c) & (!g410)) + ((!b) & (!sk[52]) & (!d) & (!c) & (g410)) + ((!b) & (!sk[52]) & (!d) & (!c) & (g410)) + ((!b) & (sk[52]) & (!d) & (!c) & (!g410)));
	assign g425 = (((!j) & (g1) & (g290) & (!g319) & (!sk[53]) & (!g424)) + ((j) & (!g1) & (!g290) & (!g319) & (!sk[53]) & (!g424)) + ((!j) & (!g1) & (g290) & (!g319) & (!sk[53]) & (!g424)) + ((!j) & (g1) & (!g290) & (!g319) & (!sk[53]) & (g424)) + ((!j) & (!g1) & (!g290) & (!g319) & (!sk[53]) & (g424)) + ((!j) & (g1) & (!g290) & (g319) & (sk[53]) & (!g424)));
	assign g426 = (((!g44) & (!j) & (!sk[54]) & (k) & (!g1)) + ((!g44) & (!j) & (!sk[54]) & (!k) & (g1)) + ((g44) & (!j) & (!sk[54]) & (!k) & (g1)));
	assign g427 = (((b) & (!e) & (!sk[55]) & (!f) & (!c) & (!a)) + ((!b) & (!e) & (!sk[55]) & (f) & (!c) & (!a)) + ((!b) & (!e) & (!sk[55]) & (!f) & (!c) & (a)) + ((!b) & (!e) & (sk[55]) & (!f) & (c) & (!a)) + ((!b) & (!e) & (sk[55]) & (!f) & (!c) & (!a)));
	assign g428 = (((!h) & (!k) & (!g15) & (!g340) & (!g426) & (!g427)) + ((!h) & (!k) & (!g15) & (!g340) & (!g426) & (!g427)) + ((h) & (k) & (!g15) & (!g340) & (!g426) & (!g427)));
	assign g429 = (((!sk[57]) & (!d) & (!e) & (g) & (!g145)) + ((!sk[57]) & (!d) & (!e) & (!g) & (g145)) + ((!sk[57]) & (d) & (!e) & (g) & (g145)));
	assign g430 = (((i) & (!sk[58]) & (!a) & (!g35) & (!g82) & (!g429)) + ((!i) & (!sk[58]) & (!a) & (g35) & (!g82) & (!g429)) + ((!i) & (!sk[58]) & (!a) & (!g35) & (!g82) & (g429)) + ((!i) & (!sk[58]) & (!a) & (!g35) & (!g82) & (g429)) + ((!i) & (!sk[58]) & (a) & (g35) & (g82) & (!g429)));
	assign g431 = (((!sk[59]) & (!f) & (!h) & (!g) & (g409)) + ((!sk[59]) & (!f) & (!h) & (g) & (!g409)) + ((sk[59]) & (f) & (!h) & (!g) & (!g409)) + ((sk[59]) & (!f) & (h) & (!g) & (!g409)));
	assign g432 = (((!j) & (!l) & (!sk[60]) & (g406) & (!g431)) + ((!j) & (!l) & (!sk[60]) & (g406) & (!g431)) + ((!j) & (!l) & (!sk[60]) & (!g406) & (g431)) + ((j) & (!l) & (sk[60]) & (!g406) & (!g431)));
	assign g433 = (((!sk[61]) & (!f) & (h) & (!g)) + ((sk[61]) & (f) & (!h) & (!g)));
	assign g434 = (((!b) & (!sk[62]) & (!l) & (a) & (!g330)) + ((!b) & (!sk[62]) & (!l) & (!a) & (g330)) + ((!b) & (!sk[62]) & (!l) & (!a) & (g330)) + ((!b) & (sk[62]) & (!l) & (!a) & (!g330)));
	assign g435 = (((e) & (!f) & (!h) & (g) & (!g212) & (g353)) + ((e) & (!f) & (!h) & (!g) & (g212) & (!g353)));
	assign g436 = (((!d) & (!c) & (!g433) & (!g410) & (!g434) & (!g435)) + ((!d) & (c) & (!g433) & (!g410) & (!g434) & (!g435)) + ((!d) & (!c) & (!g433) & (!g410) & (!g434) & (!g435)));
	assign g437 = (((!sk[65]) & (!g99) & (g146) & (!g223)) + ((!sk[65]) & (g99) & (g146) & (g223)));
	assign g438 = (((h) & (!g58) & (!sk[66]) & (!g34) & (!g71) & (!g317)) + ((!h) & (!g58) & (!sk[66]) & (g34) & (!g71) & (!g317)) + ((!h) & (!g58) & (!sk[66]) & (!g34) & (!g71) & (g317)) + ((h) & (!g58) & (!sk[66]) & (g34) & (!g71) & (g317)) + ((!h) & (g58) & (sk[66]) & (!g34) & (g71) & (!g317)));
	assign g439 = (((!g15) & (!g430) & (!g432) & (!g436) & (!g437) & (!g438)) + ((!g15) & (!g430) & (!g432) & (g436) & (!g437) & (!g438)));
	assign g440 = (((n) & (!g408) & (g423) & (!g425) & (g428) & (g439)) + ((!n) & (g408) & (g423) & (!g425) & (g428) & (g439)));
	assign g441 = (((!sk[69]) & (!g) & (!j) & (g281) & (!g361)) + ((!sk[69]) & (!g) & (!j) & (!g281) & (g361)) + ((!sk[69]) & (!g) & (j) & (!g281) & (g361)) + ((!sk[69]) & (g) & (j) & (g281) & (!g361)));
	assign g442 = (((!g41) & (!g9) & (!sk[70]) & (g20) & (!g441)) + ((!g41) & (g9) & (!sk[70]) & (!g20) & (g441)) + ((!g41) & (!g9) & (!sk[70]) & (!g20) & (g441)) + ((g41) & (g9) & (!sk[70]) & (g20) & (!g441)));
	assign g443 = (((!k) & (!l) & (!sk[71]) & (g1) & (!g319)) + ((!k) & (!l) & (!sk[71]) & (!g1) & (g319)) + ((!k) & (!l) & (!sk[71]) & (g1) & (g319)) + ((!k) & (!l) & (!sk[71]) & (g1) & (g319)));
	assign g444 = (((h) & (!g1) & (!c) & (!sk[72]) & (!g82) & (!g202)) + ((!h) & (!g1) & (c) & (!sk[72]) & (!g82) & (!g202)) + ((!h) & (!g1) & (!c) & (!sk[72]) & (!g82) & (g202)) + ((h) & (g1) & (!c) & (!sk[72]) & (!g82) & (!g202)) + ((h) & (g1) & (!c) & (!sk[72]) & (!g82) & (!g202)));
	assign g445 = (((f) & (!sk[73]) & (!g) & (!k) & (!g9) & (!c)) + ((!f) & (!sk[73]) & (!g) & (k) & (!g9) & (!c)) + ((!f) & (!sk[73]) & (!g) & (!k) & (!g9) & (c)) + ((!f) & (sk[73]) & (!g) & (!k) & (g9) & (!c)));
	assign g446 = (((!n) & (!sk[74]) & (g218) & (!g281)) + ((!n) & (!sk[74]) & (g218) & (g281)));
	assign g447 = (((g443) & (!g444) & (!g445) & (!sk[75]) & (!g446) & (!g456)) + ((!g443) & (!g444) & (g445) & (!sk[75]) & (!g446) & (!g456)) + ((!g443) & (!g444) & (!g445) & (!sk[75]) & (!g446) & (g456)) + ((!g443) & (!g444) & (!g445) & (!sk[75]) & (!g446) & (g456)));
	assign g448 = (((h) & (!sk[76]) & (!k) & (i) & (!l)) + ((!h) & (!sk[76]) & (!k) & (i) & (!l)) + ((!h) & (!sk[76]) & (!k) & (!i) & (l)) + ((!h) & (sk[76]) & (!k) & (!i) & (!l)));
	assign g449 = (((!sk[77]) & (!m) & (!k) & (g58) & (!g410)) + ((!sk[77]) & (!m) & (!k) & (!g58) & (g410)) + ((!sk[77]) & (!m) & (k) & (!g58) & (g410)));
	assign g450 = (((m) & (!sk[78]) & (!g319) & (!g395) & (!g448) & (!g449)) + ((!m) & (!sk[78]) & (!g319) & (g395) & (!g448) & (!g449)) + ((!m) & (!sk[78]) & (!g319) & (!g395) & (!g448) & (g449)) + ((m) & (!sk[78]) & (!g319) & (g395) & (!g448) & (!g449)) + ((!m) & (!sk[78]) & (!g319) & (g395) & (!g448) & (!g449)) + ((!m) & (!sk[78]) & (!g319) & (g395) & (g448) & (!g449)));
	assign g451 = (((n) & (!i) & (!g442) & (!sk[79]) & (!g447) & (!g450)) + ((!n) & (!i) & (g442) & (!sk[79]) & (!g447) & (!g450)) + ((!n) & (!i) & (!g442) & (!sk[79]) & (!g447) & (g450)) + ((!n) & (!i) & (!g442) & (!sk[79]) & (!g447) & (g450)) + ((!n) & (!i) & (!g442) & (sk[79]) & (!g447) & (!g450)) + ((!n) & (!i) & (!g442) & (!sk[79]) & (g447) & (g450)) + ((!n) & (!i) & (!g442) & (sk[79]) & (g447) & (!g450)));
	assign l2 = (((!g360) & (!g366) & (g375) & (!g392) & (!g440) & (!g451)) + ((!g360) & (!g366) & (!g375) & (!g392) & (!g440) & (!g451)) + ((!g360) & (!g366) & (!g375) & (!g392) & (!g440) & (!g451)) + ((!g360) & (!g366) & (!g375) & (!g392) & (!g440) & (!g451)) + ((!g360) & (!g366) & (!g375) & (!g392) & (!g440) & (!g451)));
	assign g453 = (((h) & (!k) & (!j) & (!g15) & (!sk[81]) & (!l)) + ((!h) & (!k) & (j) & (!g15) & (!sk[81]) & (!l)) + ((!h) & (!k) & (!j) & (!g15) & (!sk[81]) & (l)) + ((h) & (k) & (!j) & (g15) & (!sk[81]) & (!l)) + ((h) & (!k) & (!j) & (g15) & (!sk[81]) & (l)));
	assign g454 = (((!h) & (!i) & (!k) & (j) & (g15) & (!l)) + ((!h) & (i) & (!k) & (!j) & (g15) & (l)) + ((h) & (!i) & (!k) & (!j) & (g15) & (l)) + ((!h) & (!i) & (k) & (!j) & (g15) & (!l)) + ((h) & (!i) & (!k) & (j) & (g15) & (!l)) + ((!h) & (i) & (k) & (!j) & (g15) & (!l)) + ((!h) & (!i) & (!k) & (j) & (g15) & (l)) + ((!h) & (i) & (k) & (!j) & (g15) & (!l)) + ((h) & (!i) & (!k) & (j) & (g15) & (!l)));
	assign g455 = (((!sk[83]) & (!g453) & (g454) & (!g)) + ((sk[83]) & (!g453) & (!g454) & (g)) + ((sk[83]) & (!g453) & (!g454) & (!g)));
	assign g456 = (((!sk[84]) & (!n) & (g457)) + ((sk[84]) & (!n) & (!g457)));
	assign g457 = (((!sk[85]) & (!n) & (g458)) + ((!sk[85]) & (!n) & (g458)));
	assign g458 = (((!sk[86]) & (!g459) & (g460)) + ((sk[86]) & (!g459) & (!g460)));
	assign g459 = (((!sk[87]) & (!m) & (g461)) + ((!sk[87]) & (!m) & (g461)));
	assign g460 = (((!sk[88]) & (!m) & (g431)) + ((!sk[88]) & (m) & (g431)));
	assign g461 = (((!g34) & (!c) & (!sk[89]) & (l) & (!f)) + ((!g34) & (!c) & (!sk[89]) & (!l) & (f)) + ((g34) & (!c) & (sk[89]) & (!l) & (!f)) + ((!g34) & (c) & (sk[89]) & (!l) & (!f)));
	assign g462 = (((!sk[90]) & (!g463) & (g464)) + ((sk[90]) & (!g463) & (!g464)));
	assign g463 = (((!sk[91]) & (!a) & (g465)) + ((!sk[91]) & (!a) & (g465)));
	assign g464 = (((a) & (!sk[92]) & (g468)) + ((!a) & (!sk[92]) & (g468)));
	assign g465 = (((!sk[93]) & (!g466) & (g467)) + ((sk[93]) & (!g466) & (!g467)));
	assign g466 = (((!sk[94]) & (!m) & (g469)) + ((!sk[94]) & (!m) & (g469)));
	assign g467 = (((m) & (!sk[95]) & (g470)) + ((!m) & (!sk[95]) & (g470)));
	assign g468 = (((!m) & (!sk[96]) & (g471)) + ((!m) & (!sk[96]) & (g471)));
	assign g469 = (((!c) & (!sk[97]) & (!l) & (b) & (!n)) + ((!c) & (!sk[97]) & (!l) & (!b) & (n)) + ((!c) & (sk[97]) & (!l) & (!b) & (!n)) + ((!c) & (!sk[97]) & (l) & (b) & (!n)));
	assign g470 = (((!g) & (!sk[98]) & (n)) + ((g) & (sk[98]) & (!n)));
	assign g471 = (((!sk[99]) & (!c) & (!l) & (b) & (!n)) + ((!sk[99]) & (!c) & (!l) & (!b) & (n)) + ((sk[99]) & (!c) & (!l) & (!b) & (!n)) + ((!sk[99]) & (!c) & (l) & (b) & (!n)));
	assign g472 = (((!sk[100]) & (!f) & (g473)) + ((sk[100]) & (!f) & (!g473)));
	assign g473 = (((!f) & (!sk[101]) & (g474)) + ((!f) & (!sk[101]) & (g474)));
	assign g474 = (((!sk[102]) & (!g475) & (g476)) + ((sk[102]) & (!g475) & (!g476)));
	assign g475 = (((!g) & (!sk[103]) & (g477)) + ((!g) & (!sk[103]) & (g477)));
	assign g476 = (((!sk[104]) & (!g) & (g478)) + ((!sk[104]) & (g) & (g478)));
	assign g477 = (((sk[105]) & (!g35) & (!a) & (!g47) & (!d)) + ((sk[105]) & (!g35) & (!a) & (!g47) & (!d)) + ((!sk[105]) & (!g35) & (!a) & (g47) & (!d)) + ((!sk[105]) & (!g35) & (!a) & (!g47) & (d)) + ((sk[105]) & (!g35) & (!a) & (!g47) & (!d)));
	assign g478 = (((!g35) & (!a) & (!sk[106]) & (g48) & (!d)) + ((!g35) & (!a) & (!sk[106]) & (!g48) & (d)) + ((!g35) & (!a) & (!sk[106]) & (!g48) & (d)) + ((!g35) & (!a) & (!sk[106]) & (!g48) & (d)) + ((!g35) & (!a) & (sk[106]) & (!g48) & (!d)));
	assign g479 = (((!sk[107]) & (!m) & (g480)) + ((sk[107]) & (!m) & (!g480)));
	assign g480 = (((!m) & (!sk[108]) & (g481)) + ((!m) & (!sk[108]) & (g481)));
	assign g481 = (((!g482) & (!sk[109]) & (g483)) + ((!g482) & (sk[109]) & (!g483)));
	assign g482 = (((!sk[110]) & (!h) & (g484)) + ((!sk[110]) & (!h) & (g484)));
	assign g483 = (((h) & (!sk[111]) & (g485)) + ((!h) & (!sk[111]) & (g485)));
	assign g484 = (((!sk[112]) & (!g) & (!l) & (!i) & (j)) + ((!sk[112]) & (!g) & (!l) & (i) & (!j)) + ((sk[112]) & (!g) & (!l) & (!i) & (!j)) + ((!sk[112]) & (!g) & (!l) & (i) & (!j)) + ((!sk[112]) & (!g) & (!l) & (i) & (!j)));
	assign g485 = (((!g) & (!l) & (!sk[113]) & (!k) & (j)) + ((!g) & (!l) & (!sk[113]) & (k) & (!j)) + ((!g) & (!l) & (sk[113]) & (!k) & (!j)) + ((!g) & (!l) & (!sk[113]) & (k) & (!j)) + ((!g) & (!l) & (!sk[113]) & (k) & (!j)));
	assign g486 = (((!sk[114]) & (!g487) & (g488)) + ((sk[114]) & (!g487) & (!g488)));
	assign g487 = (((!sk[115]) & (!g211) & (g489)) + ((!sk[115]) & (!g211) & (g489)));
	assign g488 = (((g211) & (!sk[116]) & (g492)) + ((!g211) & (!sk[116]) & (g492)));
	assign g489 = (((!sk[117]) & (!g490) & (g491)) + ((sk[117]) & (!g490) & (!g491)));
	assign g490 = (((!sk[118]) & (!n) & (g494)) + ((!sk[118]) & (!n) & (g494)));
	assign g491 = (((!sk[119]) & (!n) & (g495)) + ((!sk[119]) & (n) & (g495)));
	assign g492 = (((!n) & (!sk[120]) & (g493)) + ((n) & (sk[120]) & (!g493)));
	assign g493 = (((!sk[121]) & (!n) & (g496)) + ((!sk[121]) & (n) & (g496)));
	assign g494 = (((!sk[122]) & (!m) & (g202) & (!g178)) + ((sk[122]) & (m) & (!g202) & (!g178)) + ((sk[122]) & (!m) & (!g202) & (g178)));
	assign g495 = (((m) & (!g202) & (!g497) & (sk[123]) & (!g191)) + ((!m) & (g202) & (!g497) & (sk[123]) & (!g191)) + ((!m) & (!g202) & (g497) & (!sk[123]) & (!g191)) + ((!m) & (!g202) & (g497) & (!sk[123]) & (g191)) + ((!m) & (!g202) & (!g497) & (!sk[123]) & (g191)));
	assign g496 = (((!sk[124]) & (!m) & (g202) & (!g497)) + ((sk[124]) & (m) & (!g202) & (!g497)) + ((sk[124]) & (!m) & (!g202) & (g497)));
	assign g497 = (((!h) & (!sk[125]) & (g498)) + ((h) & (sk[125]) & (!g498)));
	assign g498 = (((!sk[126]) & (!h) & (g499)) + ((!sk[126]) & (h) & (g499)));
	assign g499 = (((!g500) & (!sk[127]) & (g501)) + ((!g500) & (sk[127]) & (!g501)));
	assign g500 = (((!sk[0]) & (!f) & (g502)) + ((!sk[0]) & (!f) & (g502)));
	assign g501 = (((f) & (!sk[1]) & (g503)) + ((!f) & (!sk[1]) & (g503)));
	assign g502 = (((!g176) & (!g) & (!g39) & (!sk[2]) & (i)) + ((g176) & (!g) & (g39) & (!sk[2]) & (!i)) + ((!g176) & (g) & (g39) & (!sk[2]) & (!i)) + ((!g176) & (!g) & (g39) & (!sk[2]) & (!i)));
	assign g503 = (((!sk[3]) & (!g176) & (!g) & (!g43) & (i)) + ((!sk[3]) & (!g176) & (!g) & (g43) & (!i)) + ((sk[3]) & (g176) & (!g) & (!g43) & (!i)) + ((sk[3]) & (!g176) & (g) & (!g43) & (!i)));
	assign g504 = (((!h) & (!sk[4]) & (g505)) + ((h) & (sk[4]) & (!g505)));
	assign g505 = (((!sk[5]) & (!h) & (g506)) + ((!sk[5]) & (h) & (g506)));
	assign g506 = (((!g507) & (!sk[6]) & (g508)) + ((!g507) & (sk[6]) & (!g508)));
	assign g507 = (((!f) & (!sk[7]) & (g509)) + ((!f) & (!sk[7]) & (g509)));
	assign g508 = (((!sk[8]) & (!f) & (g510)) + ((!sk[8]) & (f) & (g510)));
	assign g509 = (((sk[9]) & (!g176) & (j) & (!g39) & (!g)) + ((!sk[9]) & (!g176) & (!j) & (g39) & (!g)) + ((!sk[9]) & (g176) & (!j) & (g39) & (!g)) + ((!sk[9]) & (!g176) & (!j) & (!g39) & (g)) + ((!sk[9]) & (!g176) & (!j) & (g39) & (g)));
	assign g510 = (((sk[10]) & (!g176) & (j) & (!g43) & (!g)) + ((!sk[10]) & (!g176) & (!j) & (g43) & (!g)) + ((!sk[10]) & (!g176) & (!j) & (!g43) & (g)) + ((sk[10]) & (g176) & (!j) & (!g43) & (!g)));
	assign g511 = (((!sk[11]) & (!g15) & (g512)) + ((sk[11]) & (g15) & (!g512)));
	assign g512 = (((!sk[12]) & (!g15) & (g513)) + ((!sk[12]) & (g15) & (g513)));
	assign g513 = (((!g514) & (!sk[13]) & (g515)) + ((!g514) & (sk[13]) & (!g515)));
	assign g514 = (((!sk[14]) & (!l) & (g516)) + ((!sk[14]) & (!l) & (g516)));
	assign g515 = (((!sk[15]) & (!l) & (g517)) + ((!sk[15]) & (l) & (g517)));
	assign g516 = (((!i) & (sk[16]) & (g134) & (!k) & (!g)) + ((!i) & (!sk[16]) & (!g134) & (k) & (!g)) + ((!i) & (!sk[16]) & (!g134) & (!k) & (g)) + ((!i) & (!sk[16]) & (!g134) & (!k) & (g)) + ((!i) & (sk[16]) & (!g134) & (!k) & (!g)));
	assign g517 = (((!i) & (!g134) & (!sk[17]) & (h) & (!g)) + ((!i) & (!g134) & (!sk[17]) & (!h) & (g)) + ((!i) & (!g134) & (sk[17]) & (!h) & (!g)) + ((!i) & (!g134) & (!sk[17]) & (!h) & (g)) + ((!i) & (g134) & (!sk[17]) & (!h) & (g)));
	assign g518 = (((!j) & (!sk[18]) & (g519)) + ((j) & (sk[18]) & (!g519)));
	assign g519 = (((j) & (!sk[19]) & (g520)) + ((!j) & (!sk[19]) & (g520)));
	assign g520 = (((!sk[20]) & (!g521) & (g522)) + ((sk[20]) & (!g521) & (!g522)));
	assign g521 = (((!l) & (!sk[21]) & (g523)) + ((!l) & (!sk[21]) & (g523)));
	assign g522 = (((!sk[22]) & (!l) & (g524)) + ((!sk[22]) & (l) & (g524)));
	assign g523 = (((!sk[23]) & (!i) & (g149)) + ((sk[23]) & (!i) & (!g149)));
	assign g524 = (((!g147) & (!sk[24]) & (!i) & (!g151) & (k)) + ((!g147) & (!sk[24]) & (!i) & (g151) & (!k)) + ((!g147) & (!sk[24]) & (!i) & (g151) & (!k)) + ((!g147) & (!sk[24]) & (!i) & (g151) & (!k)));
	assign g525 = (((!h) & (!sk[25]) & (g526)) + ((!h) & (sk[25]) & (!g526)));
	assign g526 = (((!sk[26]) & (!h) & (g527)) + ((!sk[26]) & (!h) & (g527)));
	assign g527 = (((!sk[27]) & (!g528) & (g529)) + ((sk[27]) & (!g528) & (!g529)));
	assign g528 = (((!f) & (!sk[28]) & (g530)) + ((!f) & (!sk[28]) & (g530)));
	assign g529 = (((f) & (!sk[29]) & (g531)) + ((!f) & (!sk[29]) & (g531)));
	assign g530 = (((!g) & (!e) & (sk[30]) & (!g131) & (!g88)) + ((!g) & (e) & (!sk[30]) & (g131) & (!g88)) + ((!g) & (!e) & (!sk[30]) & (g131) & (!g88)) + ((!g) & (!e) & (!sk[30]) & (!g131) & (g88)) + ((!g) & (!e) & (!sk[30]) & (g131) & (g88)));
	assign g531 = (((!g) & (!e) & (sk[31]) & (!g132) & (!g88)) + ((!g) & (e) & (!sk[31]) & (g132) & (!g88)) + ((!g) & (!e) & (!sk[31]) & (g132) & (!g88)) + ((!g) & (!e) & (!sk[31]) & (!g132) & (g88)) + ((!g) & (!e) & (!sk[31]) & (g132) & (g88)));
	assign g532 = (((!h) & (!sk[32]) & (g533)) + ((h) & (sk[32]) & (!g533)));
	assign g533 = (((!sk[33]) & (!h) & (g534)) + ((!sk[33]) & (h) & (g534)));
	assign g534 = (((!sk[34]) & (!g535) & (g536)) + ((sk[34]) & (!g535) & (!g536)));
	assign g535 = (((!f) & (!sk[35]) & (g537)) + ((!f) & (!sk[35]) & (g537)));
	assign g536 = (((!sk[36]) & (!f) & (g538)) + ((!sk[36]) & (f) & (g538)));
	assign g537 = (((!g88) & (!e) & (!g131) & (!sk[37]) & (g)) + ((g88) & (!e) & (g131) & (!sk[37]) & (!g)) + ((!g88) & (e) & (g131) & (!sk[37]) & (!g)) + ((!g88) & (!e) & (g131) & (!sk[37]) & (!g)));
	assign g538 = (((!g88) & (!e) & (!sk[38]) & (!g132) & (g)) + ((g88) & (!e) & (!sk[38]) & (g132) & (!g)) + ((!g88) & (e) & (!sk[38]) & (g132) & (!g)) + ((!g88) & (!e) & (!sk[38]) & (g132) & (!g)));
	assign g539 = (((!g540) & (!sk[39]) & (g541)) + ((!g540) & (sk[39]) & (!g541)));
	assign g540 = (((!sk[40]) & (!g101) & (g542)) + ((!sk[40]) & (!g101) & (g542)));
	assign g541 = (((g101) & (!sk[41]) & (g545)) + ((!g101) & (!sk[41]) & (g545)));
	assign g542 = (((!sk[42]) & (!g543) & (g544)) + ((sk[42]) & (!g543) & (!g544)));
	assign g543 = (((!e) & (!sk[43]) & (g547)) + ((!e) & (!sk[43]) & (g547)));
	assign g544 = (((e) & (!sk[44]) & (g548)) + ((!e) & (!sk[44]) & (g548)));
	assign g545 = (((!sk[45]) & (!e) & (g546)) + ((sk[45]) & (e) & (!g546)));
	assign g546 = (((e) & (!sk[46]) & (g549)) + ((!e) & (!sk[46]) & (g549)));
	assign g547 = (((!c) & (!sk[47]) & (d)) + ((!c) & (sk[47]) & (!d)) + ((!c) & (!sk[47]) & (d)));
	assign g548 = (((!sk[48]) & (!g81) & (!f) & (g455) & (!d)) + ((!sk[48]) & (!g81) & (!f) & (!g455) & (d)) + ((sk[48]) & (!g81) & (!f) & (!g455) & (!d)) + ((!sk[48]) & (g81) & (!f) & (!g455) & (d)) + ((!sk[48]) & (!g81) & (f) & (!g455) & (d)));
	assign g549 = (((!g81) & (!f) & (!sk[49]) & (g455) & (!d)) + ((!g81) & (!f) & (!sk[49]) & (!g455) & (d)) + ((!g81) & (!f) & (sk[49]) & (!g455) & (!d)) + ((g81) & (!f) & (!sk[49]) & (!g455) & (d)) + ((!g81) & (f) & (!sk[49]) & (!g455) & (d)));

endmodule