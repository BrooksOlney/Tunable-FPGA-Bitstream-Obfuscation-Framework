module misex3x6xv (a, b, c, d, e, f, g, h, i, j, k, l, m, n, r2, s2, p2, q2, t2, u2, j2, k2, h2, i2, n2, o2, l2, m2);

	input a;
	input b;
	input c;
	input d;
	input e;
	input f;
	input g;
	input h;
	input i;
	input j;
	input k;
	input l;
	input m;
	input n;
	output r2;
	output s2;
	output p2;
	output q2;
	output t2;
	output u2;
	output j2;
	output k2;
	output h2;
	output i2;
	output n2;
	output o2;
	output l2;
	output m2;

	wire [855 : 0] sk /* synthesis noprune */;

	lut_sub lut_3 ({sk[0], x5175x, x5098x, x5099x, x5135x, x5136x, x5137x}, r2);
	defparam lut_3.LUT_SIZE = 7;
	defparam lut_3.mask = 128'h5f5fffff5f5fffff7fffffffffffffff;

	lut_sub lut_10 ({sk[1], x5232x, x5233x, x5263x, x5267x, x7491x}, s2);
	defparam lut_10.LUT_SIZE = 6;
	defparam lut_10.mask = 64'h00ff00ffbfffffff;

	lut_sub lut_16 ({sk[2], x5307x, x5308x, x5327x, x5328x, x5329x, x5330x}, p2);
	defparam lut_16.LUT_SIZE = 7;
	defparam lut_16.mask = 128'h03133333777777777fffffffffffffff;

	lut_sub lut_23 ({sk[3], n_n1786, x5408x, x5409x, x5443x, x5444x, x5448x}, q2);
	defparam lut_23.LUT_SIZE = 7;
	defparam lut_23.mask = 128'h03133333777777777fffffffffffffff;

	lut_sub lut_30 ({sk[4], x5523x, x5466x, x5467x, n_n1425, x5517x, x5518x}, t2);
	defparam lut_30.LUT_SIZE = 7;
	defparam lut_30.mask = 128'h03133333777777777fffffffffffffff;

	lut_sub lut_37 ({sk[5], x5625x, x5621x, x5622x}, u2);
	defparam lut_37.LUT_SIZE = 4;
	defparam lut_37.mask = 16'h337f;

	lut_sub lut_41 ({sk[6], x5653x, x116x, x199x, x319x, x5648x}, j2);
	defparam lut_41.LUT_SIZE = 6;
	defparam lut_41.mask = 64'h5f7f5f7f7fffffff;

	lut_sub lut_47 ({sk[7], c, x5672x, x53x, x91x, x392x, x5667x}, k2);
	defparam lut_47.LUT_SIZE = 7;
	defparam lut_47.mask = 128'h5577ffffffffffff5f7fffff5f5fffff;

	lut_sub lut_52 ({sk[8], n_n1874, x5718x, x5719x, x5720x, x5721x, x5722x}, h2);
	defparam lut_52.LUT_SIZE = 7;
	defparam lut_52.mask = 128'h5577ffffffffffff7fffffffffffffff;

	lut_sub lut_59 ({sk[9], x5812x, x5807x, x5808x}, i2);
	defparam lut_59.LUT_SIZE = 4;
	defparam lut_59.mask = 16'h3f7f;

	lut_sub lut_63 ({sk[10], x5874x, x5848x, x5849x, x5850x, x5851x}, n2);
	defparam lut_63.LUT_SIZE = 6;
	defparam lut_63.mask = 64'h5f7f5f7f7fffffff;

	lut_sub lut_69 ({sk[11], n_n1653, x5936x, x5937x, x5938x}, o2);
	defparam lut_69.LUT_SIZE = 5;
	defparam lut_69.mask = 32'h5fff7fff;

	lut_sub lut_74 ({sk[12], n_n2020, n_n2019, x6303x, x6304x}, l2);
	defparam lut_74.LUT_SIZE = 5;
	defparam lut_74.mask = 32'h5fff7fff;

	lut_sub lut_79 ({sk[13], x199x, x157x, x267x, n_n1939, x6317x, x6322x}, m2);
	defparam lut_79.LUT_SIZE = 7;
	defparam lut_79.mask = 128'h5577ffffffffffff7fffffffffffffff;

	lut_sub lut_86 ({sk[14], x46x, x67x, x1126x, x5158x, x5170x, x5174x}, x5175x);
	defparam lut_86.LUT_SIZE = 7;
	defparam lut_86.mask = 128'h5577ffffffffffff7fff7fff7fffffff;

	lut_sub lut_92 ({sk[15], x187x, n_n703, x1208x, x5088x, n_n698, x5093x}, x5098x);
	defparam lut_92.LUT_SIZE = 7;
	defparam lut_92.mask = 128'h5577ffffffffffff55555fff77777fff;

	lut_sub lut_97 ({sk[16], n_n709, x417x, x1196x, x5090x, x5091x, x5092x}, x5099x);
	defparam lut_97.LUT_SIZE = 7;
	defparam lut_97.mask = 128'h5577ffffffffffff7fff7fff7fffffff;

	lut_sub lut_103 ({sk[17], n_n816, x315x, x302x, n_n825, x5121x, x5130x}, x5135x);
	defparam lut_103.LUT_SIZE = 7;
	defparam lut_103.mask = 128'h5577ffffffffffff777f777f777fffff;

	lut_sub lut_108 ({sk[18], n, x110x, x77x, x21x, x1161x, x5124x}, x5136x);
	defparam lut_108.LUT_SIZE = 7;
	defparam lut_108.mask = 128'h5577ffffffffffff777777ff77777fff;

	lut_sub lut_113 ({sk[19], x5117x, x5118x, x5119x, x5120x, x5133x}, x5137x);
	defparam lut_113.LUT_SIZE = 6;
	defparam lut_113.mask = 64'h5f7f5f7f7fffffff;

	lut_sub lut_119 ({sk[20], n, x377x, x115x, x21x, x5225x, x5228x}, x5232x);
	defparam lut_119.LUT_SIZE = 7;
	defparam lut_119.mask = 128'h5577ffffffffffff77777777777f7f7f;

	lut_sub lut_124 ({sk[21], x5221x, x5222x, x5226x, x5230x}, x5233x);
	defparam lut_124.LUT_SIZE = 5;
	defparam lut_124.mask = 32'h5fff7fff;

	lut_sub lut_129 ({sk[22], n_n904, x54x, x102x, x195x, x297x, x1049x}, x5263x);
	defparam lut_129.LUT_SIZE = 7;
	defparam lut_129.mask = 128'h5577ffffffffffff555577775fff7fff;

	lut_sub lut_134 ({sk[23], a, x171x, x138x, x1060x, x5260x, x5264x}, x5267x);
	defparam lut_134.LUT_SIZE = 7;
	defparam lut_134.mask = 128'h5577ffffffffffff7f7f7f7f7f7f7fff;

	lut_sub lut_139 ({sk[24], x5211x, x1047x, x1048x, x5209x, x5210x, x5256x}, x7491x);
	defparam lut_139.LUT_SIZE = 7;
	defparam lut_139.mask = 128'h5577ffffffffffff8000000000000000;

	lut_sub lut_141 ({sk[25], x125x, x265x, x5294x, x5295x, x5298x, x5299x}, x5307x);
	defparam lut_141.LUT_SIZE = 7;
	defparam lut_141.mask = 128'h5577ffffffffffff7fff7fff7fffffff;

	lut_sub lut_147 ({sk[26], x5291x, x5292x, x5296x, x5302x, x7490x}, x5308x);
	defparam lut_147.LUT_SIZE = 6;
	defparam lut_147.mask = 64'h5f7f5f7fbfffffff;

	lut_sub lut_153 ({sk[27], n_n920, n_n1193, x62x, x228x, x265x, x5324x}, x5327x);
	defparam lut_153.LUT_SIZE = 7;
	defparam lut_153.mask = 128'h5577ffffffffffff5577557755777f7f;

	lut_sub lut_158 ({sk[28], i, j, x58x, n_n1220, x82x, x240x}, x5328x);
	defparam lut_158.LUT_SIZE = 7;
	defparam lut_158.mask = 128'h5577ffffffffffff0000050500330537;

	lut_sub lut_161 ({sk[29], k, n_n1187, x83x, x82x, x265x, x51x}, x5329x);
	defparam lut_161.LUT_SIZE = 7;
	defparam lut_161.mask = 128'h5577ffffffffffff000011110000111f;

	lut_sub lut_164 ({sk[30], x125x, x228x, x5322x, x5325x}, x5330x);
	defparam lut_164.LUT_SIZE = 5;
	defparam lut_164.mask = 32'h5fff777f;

	lut_sub lut_168 ({sk[31], x5363x, x5364x, x5394x, x5395x, x5396x, x5397x}, n_n1786);
	defparam lut_168.LUT_SIZE = 7;
	defparam lut_168.mask = 128'h5577ffffffffffff7fffffffffffffff;

	lut_sub lut_175 ({sk[32], f, x15x, x194x, x142x, x5404x, x7489x}, x5408x);
	defparam lut_175.LUT_SIZE = 7;
	defparam lut_175.mask = 128'h5577ffffffffffffbbbbbbbbbbbbbbbf;

	lut_sub lut_179 ({sk[33], x54x, x99x, x106x, x142x}, x5409x);
	defparam lut_179.LUT_SIZE = 5;
	defparam lut_179.mask = 32'h5fff153f;

	lut_sub lut_184 ({sk[34], x54x, x62x, n_n1155, x5431x, x5432x, x5433x}, x5443x);
	defparam lut_184.LUT_SIZE = 7;
	defparam lut_184.mask = 128'h5577ffffffffffff7f7f7f7f7f7f7fff;

	lut_sub lut_189 ({sk[35], n_n1187, x51x, x291x, x380x, x906x, x5434x}, x5444x);
	defparam lut_189.LUT_SIZE = 7;
	defparam lut_189.mask = 128'h5577ffffffffffff777f777f777f7f7f;

	lut_sub lut_194 ({sk[36], x5429x, x5430x, x5437x, x5445x, x7488x}, x5448x);
	defparam lut_194.LUT_SIZE = 6;
	defparam lut_194.mask = 64'h5f7f5f7fbfffffff;

	lut_sub lut_200 ({sk[37], x5508x, x5509x, x5513x, x5515x, x7487x}, x5523x);
	defparam lut_200.LUT_SIZE = 6;
	defparam lut_200.mask = 64'h5f7f5f7fbfffffff;

	lut_sub lut_206 ({sk[38], b, x53x, x94x, x135x, x43x, x5462x}, x5466x);
	defparam lut_206.LUT_SIZE = 7;
	defparam lut_206.mask = 128'h5577ffffffffffff5577557755775f7f;

	lut_sub lut_210 ({sk[39], n_n730, n_n662, x94x, x126x, x874x, x5465x}, x5467x);
	defparam lut_210.LUT_SIZE = 7;
	defparam lut_210.mask = 128'h5577ffffffffffff77777f7f77ff7fff;

	lut_sub lut_215 ({sk[40], x102x, x138x, x390x, x43x, x5473x, x5474x}, n_n1425);
	defparam lut_215.LUT_SIZE = 7;
	defparam lut_215.mask = 128'h5577ffffffffffff777f7f7f7f7f7f7f;

	lut_sub lut_221 ({sk[41], a, x249x, x151x, x842x, x5506x, x7486x}, x5517x);
	defparam lut_221.LUT_SIZE = 7;
	defparam lut_221.mask = 128'h5577ffffffffffffbfbfbfbfbfbfbfff;

	lut_sub lut_226 ({sk[42], a, d, e, x102x, x390x, x5512x}, x5518x);
	defparam lut_226.LUT_SIZE = 7;
	defparam lut_226.mask = 128'h5577ffffffffffff5555555555557f55;

	lut_sub lut_230 ({sk[43], x5581x, x5582x, x5583x, x5584x, x5619x, x5620x}, x5625x);
	defparam lut_230.LUT_SIZE = 7;
	defparam lut_230.mask = 128'h5577ffffffffffff7fffffffffffffff;

	lut_sub lut_237 ({sk[44], n_n1187, x83x, x51x, x246x, x5612x, x5613x}, x5621x);
	defparam lut_237.LUT_SIZE = 7;
	defparam lut_237.mask = 128'h5577ffffffffffff77777777777777f7;

	lut_sub lut_241 ({sk[45], n_n1187, x148x, x83x, x82x, x99x, x246x}, x5622x);
	defparam lut_241.LUT_SIZE = 7;
	defparam lut_241.mask = 128'h5577ffffffffffff00003f0f11113f1f;

	lut_sub lut_245 ({sk[46], n_n1080, x382x, x5627x, n_n2499, x91x, x392x}, x5653x);
	defparam lut_245.LUT_SIZE = 7;
	defparam lut_245.mask = 128'h5577ffffffffffff3f3f3fff7f7f7fff;

	lut_sub lut_250 ({sk[47], k, x83x, n_n1104, x779x, n_n1204, n_n975}, x116x);
	defparam lut_250.LUT_SIZE = 7;
	defparam lut_250.mask = 128'h5577ffffffffffff0f0f0f1f0f0f0f0f;

	lut_sub lut_253 ({sk[48], h, i, j, n_n2602, n_n987, x370x}, x199x);
	defparam lut_253.LUT_SIZE = 7;
	defparam lut_253.mask = 128'h5577ffffffffffff0f0f0f1f0f0f0f0f;

	lut_sub lut_256 ({sk[49], n_n973, n_n1195, n_n1085, n_n982, x372x, x308x}, x319x);
	defparam lut_256.LUT_SIZE = 7;
	defparam lut_256.mask = 128'h5577ffffffffffff0003000300035557;

	lut_sub lut_259 ({sk[50], n_n1138, n_n1159, n_n978, x367x, x283x, x372x}, x5648x);
	defparam lut_259.LUT_SIZE = 7;
	defparam lut_259.mask = 128'h5577ffffffffffff0011001100110f1f;

	lut_sub lut_262 ({sk[51], x319x, x157x, x267x, x5666x}, x5672x);
	defparam lut_262.LUT_SIZE = 5;
	defparam lut_262.mask = 32'h5fff7fff;

	lut_sub lut_267 ({sk[52], d, e}, x53x);
	defparam lut_267.LUT_SIZE = 3;
	defparam lut_267.mask = 8'h54;

	lut_sub lut_269 ({sk[53], n_n1195, n_n987, n_n1085, x370x, n_n975, x308x}, x91x);
	defparam lut_269.LUT_SIZE = 7;
	defparam lut_269.mask = 128'h5577ffffffffffff0000000f1111111f;

	lut_sub lut_272 ({sk[54], i, j, k, l, n_n1165, n_n971}, x392x);
	defparam lut_272.LUT_SIZE = 7;
	defparam lut_272.mask = 128'h5577ffffffffffff0000000000000001;

	lut_sub lut_274 ({sk[55], i, n_n1080, n_n1190, n_n1202, n_n1039, n_n2493}, x5667x);
	defparam lut_274.LUT_SIZE = 7;
	defparam lut_274.mask = 128'h5577ffffffffffff5555555755555555;

	lut_sub lut_277 ({sk[56], x92x, x193x, x746x, x5684x, x5686x, x5687x}, n_n1874);
	defparam lut_277.LUT_SIZE = 7;
	defparam lut_277.mask = 128'h5577ffffffffffff7fff7fff7fffffff;

	lut_sub lut_283 ({sk[57], n_n949, x94x, x270x, x722x, x5711x}, x5718x);
	defparam lut_283.LUT_SIZE = 6;
	defparam lut_283.mask = 64'h5f7f5f7f7f7f7fff;

	lut_sub lut_288 ({sk[58], x57x, n_n949, x120x, x239x, x123x, x243x}, x5719x);
	defparam lut_288.LUT_SIZE = 7;
	defparam lut_288.mask = 128'h5577ffffffffffff00110f1f00000f0f;

	lut_sub lut_291 ({sk[59], x713x, x727x, x5706x, x5707x}, x5720x);
	defparam lut_291.LUT_SIZE = 5;
	defparam lut_291.mask = 32'h5fff7fff;

	lut_sub lut_296 ({sk[60], n_n876, n_n997, x182x, n_n864, x716x, x717x}, x5721x);
	defparam lut_296.LUT_SIZE = 7;
	defparam lut_296.mask = 128'h5577ffffffffffff777777ff777f77ff;

	lut_sub lut_301 ({sk[61], a, x249x, n_n997, x123x, x174x, x5710x}, x5722x);
	defparam lut_301.LUT_SIZE = 7;
	defparam lut_301.mask = 128'h5577ffffffffffff555f555f555f7f7f;

	lut_sub lut_306 ({sk[62], n_n1919, x5765x, x5766x, n_n1939, x5799x, x5806x}, x5812x);
	defparam lut_306.LUT_SIZE = 7;
	defparam lut_306.mask = 128'h5577ffffffffffff7fffffffffffffff;

	lut_sub lut_313 ({sk[63], a, x249x, x123x, x5794x, x5795x, x7482x}, x5807x);
	defparam lut_313.LUT_SIZE = 7;
	defparam lut_313.mask = 128'h5577ffffffffffffbfbfbfbfbfbfbfff;

	lut_sub lut_318 ({sk[64], x5731x, x5790x, x5791x, x5797x, x7481x}, x5808x);
	defparam lut_318.LUT_SIZE = 6;
	defparam lut_318.mask = 64'h5f7f5f7fbfffffff;

	lut_sub lut_324 ({sk[65], x5829x, x5870x, x5871x, x7480x}, x5874x);
	defparam lut_324.LUT_SIZE = 5;
	defparam lut_324.mask = 32'h5fffbfff;

	lut_sub lut_329 ({sk[66], x264x, x15x, n_n2953, x5841x, x5842x, x5843x}, x5848x);
	defparam lut_329.LUT_SIZE = 7;
	defparam lut_329.mask = 128'h5577ffffffffffff7fff7fff7fffffff;

	lut_sub lut_335 ({sk[67], n_n1187, x82x, x51x, x81x, x5831x, x5839x}, x5849x);
	defparam lut_335.LUT_SIZE = 7;
	defparam lut_335.mask = 128'h5577ffffffffffff00005555003f557f;

	lut_sub lut_339 ({sk[68], n_n1187, x82x, x51x, n_n605, x81x, x5831x}, x5850x);
	defparam lut_339.LUT_SIZE = 7;
	defparam lut_339.mask = 128'h5577ffffffffffff00007777000f777f;

	lut_sub lut_343 ({sk[69], x29x, x257x, x81x, x5831x, x5833x, x5847x}, x5851x);
	defparam lut_343.LUT_SIZE = 7;
	defparam lut_343.mask = 128'h5577ffffffffffff5777577757775fff;

	lut_sub lut_349 ({sk[70], x5903x, x5904x, x5905x, x5906x}, n_n1653);
	defparam lut_349.LUT_SIZE = 5;
	defparam lut_349.mask = 32'h5fff7fff;

	lut_sub lut_354 ({sk[71], k, n_n1187, x50x, x5924x, x5925x, x5926x}, x5936x);
	defparam lut_354.LUT_SIZE = 7;
	defparam lut_354.mask = 128'h5577ffffffffffff7f7f7f7f7f7f7fff;

	lut_sub lut_359 ({sk[72], x320x, x547x, x5919x, x5920x, x5921x, x5922x}, x5937x);
	defparam lut_359.LUT_SIZE = 7;
	defparam lut_359.mask = 128'h5577ffffffffffff7fffffffffffffff;

	lut_sub lut_366 ({sk[73], n_n1210, x235x, x548x, x555x, x556x, x5923x}, x5938x);
	defparam lut_366.LUT_SIZE = 7;
	defparam lut_366.mask = 128'h5577ffffffffffff7fff7fff7fffffff;

	lut_sub lut_372 ({sk[74], x6001x, x6002x, x6040x, x6041x, x6068x, x6069x}, n_n2020);
	defparam lut_372.LUT_SIZE = 7;
	defparam lut_372.mask = 128'h5577ffffffffffff7fffffffffffffff;

	lut_sub lut_379 ({sk[75], x6209x, x6210x, x6255x, x6256x, x6285x}, n_n2019);
	defparam lut_379.LUT_SIZE = 6;
	defparam lut_379.mask = 64'h5f7f5f7f7fffffff;

	lut_sub lut_385 ({sk[76], x6106x, x6093x, x6094x, x6095x, x6096x, x6301x}, x6303x);
	defparam lut_385.LUT_SIZE = 7;
	defparam lut_385.mask = 128'h5577ffffffffffff7fffffffffffffff;

	lut_sub lut_392 ({sk[77], n_n2060, x6139x, n_n2023, x7472x}, x6304x);
	defparam lut_392.LUT_SIZE = 5;
	defparam lut_392.mask = 32'h5fffbfff;

	lut_sub lut_397 ({sk[78], e, x112x, n_n978, x764x, n_n1264, n_n1253}, x157x);
	defparam lut_397.LUT_SIZE = 7;
	defparam lut_397.mask = 128'h5577ffffffffffff0f0f0f0f0f0f0f1f;

	lut_sub lut_400 ({sk[79], c, d, e, n_n1201, n_n2499, x141x}, x267x);
	defparam lut_400.LUT_SIZE = 7;
	defparam lut_400.mask = 128'h5577ffffffffffff3333333333333337;

	lut_sub lut_403 ({sk[80], x319x, x670x, x5771x, x5772x, x5773x}, n_n1939);
	defparam lut_403.LUT_SIZE = 6;
	defparam lut_403.mask = 64'h5f7f5f7f7fffffff;

	lut_sub lut_409 ({sk[81], f, n, x131x, n_n1118, x407x, x26x}, x6317x);
	defparam lut_409.LUT_SIZE = 7;
	defparam lut_409.mask = 128'h5577ffffffffffff5557555555555555;

	lut_sub lut_412 ({sk[82], n_n1028, x91x, x116x, x370x, x384x, x6316x}, x6322x);
	defparam lut_412.LUT_SIZE = 7;
	defparam lut_412.mask = 128'h5577ffffffffffff55ffffff57ffffff;

	lut_sub lut_417 ({sk[83], g, h, i, j, l}, x46x);
	defparam lut_417.LUT_SIZE = 6;
	defparam lut_417.mask = 64'h5f7f5f7f00440572;

	lut_sub lut_422 ({sk[84], a, b, c, d, e, n_n1187}, x67x);
	defparam lut_422.LUT_SIZE = 7;
	defparam lut_422.mask = 128'h5577ffffffffffff0000000000000414;

	lut_sub lut_425 ({sk[85], g, i, j, k, l, x67x}, x1126x);
	defparam lut_425.LUT_SIZE = 7;
	defparam lut_425.mask = 128'h5577ffffffffffff0000000000510010;

	lut_sub lut_429 ({sk[86], n_n1089, n_n842, n_n1161, n_n713, x75x, x84x}, x5158x);
	defparam lut_429.LUT_SIZE = 7;
	defparam lut_429.mask = 128'h5577ffffffffffff0003000300035557;

	lut_sub lut_432 ({sk[87], x110x, x172x, x5159x, x5160x, x5161x}, x5170x);
	defparam lut_432.LUT_SIZE = 6;
	defparam lut_432.mask = 64'h5f7f5f7f7f7f7fff;

	lut_sub lut_437 ({sk[88], b, x53x, x187x, x5157x, x5168x, x7496x}, x5174x);
	defparam lut_437.LUT_SIZE = 7;
	defparam lut_437.mask = 128'h5577ffffffffffff7f7f7f7f7f7f7fff;

	lut_sub lut_442 ({sk[89], x229x, n_n1165, n_n1229, x101x, n_n1069, x847x}, x5508x);
	defparam lut_442.LUT_SIZE = 7;
	defparam lut_442.mask = 128'h5577ffffffffffff5555555555555d55;

	lut_sub lut_445 ({sk[90], m, n, x101x, n_n1203, x184x, x49x}, x5509x);
	defparam lut_445.LUT_SIZE = 7;
	defparam lut_445.mask = 128'h5577ffffffffffff000f111100001111;

	lut_sub lut_448 ({sk[91], b, d, f, x46x, x120x, x846x}, x5513x);
	defparam lut_448.LUT_SIZE = 7;
	defparam lut_448.mask = 128'h5577ffffffffffff5555555755555555;

	lut_sub lut_451 ({sk[92], d, f, g, x38x, x74x, x92x}, x5515x);
	defparam lut_451.LUT_SIZE = 7;
	defparam lut_451.mask = 128'h5577ffffffffffff0505050705050505;

	lut_sub lut_454 ({sk[93], x112x, x256x, n_n730, x92x, x120x, x183x}, x7487x);
	defparam lut_454.LUT_SIZE = 7;
	defparam lut_454.mask = 128'h5577fffffffffffffffffcfcffeefcec;

	lut_sub lut_462 ({sk[94], x5560x, x5561x, x5574x}, x5581x);
	defparam lut_462.LUT_SIZE = 4;
	defparam lut_462.mask = 16'h3f7f;

	lut_sub lut_466 ({sk[95], x93x, n_n1210, x164x, x5564x, x5565x, x5566x}, x5582x);
	defparam lut_466.LUT_SIZE = 7;
	defparam lut_466.mask = 128'h5577ffffffffffff7f7f7f7f7f7f7fff;

	lut_sub lut_471 ({sk[96], n_n1201, x49x, x837x, x5526x, x5568x, x5577x}, x5583x);
	defparam lut_471.LUT_SIZE = 7;
	defparam lut_471.mask = 128'h5577ffffffffffff77ff77ff77ff7fff;

	lut_sub lut_476 ({sk[97], x5558x, x5559x, x5569x, x5570x, x5571x}, x5584x);
	defparam lut_476.LUT_SIZE = 6;
	defparam lut_476.mask = 64'h5f7f5f7f7fffffff;

	lut_sub lut_482 ({sk[98], x75x, x238x, x33x, x841x, x5557x, x5607x}, x5619x);
	defparam lut_482.LUT_SIZE = 7;
	defparam lut_482.mask = 128'h5577ffffffffffff555555ff7f7f7fff;

	lut_sub lut_487 ({sk[99], x5608x, x5609x, x5611x, x7485x}, x5620x);
	defparam lut_487.LUT_SIZE = 5;
	defparam lut_487.mask = 32'h5fffbfff;

	lut_sub lut_492 ({sk[100], c, d, e}, n_n1080);
	defparam lut_492.LUT_SIZE = 4;
	defparam lut_492.mask = 16'h3f80;

	lut_sub lut_494 ({sk[101], i, j, k, l, m, n}, x382x);
	defparam lut_494.LUT_SIZE = 7;
	defparam lut_494.mask = 128'h5577ffffffffffff0000000800000000;

	lut_sub lut_496 ({sk[102], c, d, e, f, g, h}, x5627x);
	defparam lut_496.LUT_SIZE = 7;
	defparam lut_496.mask = 128'h5577ffffffffffff0000000000002000;

	lut_sub lut_498 ({sk[103], c, x78x, x5632x, n_n992, n_n1222, n_n1260}, n_n2499);
	defparam lut_498.LUT_SIZE = 7;
	defparam lut_498.mask = 128'h5577ffffffffffff0000000000020000;

	lut_sub lut_500 ({sk[104], l, n_n2602, n_n987, n_n1210, n_n988, x283x}, x5666x);
	defparam lut_500.LUT_SIZE = 7;
	defparam lut_500.mask = 128'h5577ffffffffffff0000ffff0001ffff;

	lut_sub lut_503 ({sk[105], x223x, x55x, x18x, x388x, x5738x, x7484x}, n_n1919);
	defparam lut_503.LUT_SIZE = 7;
	defparam lut_503.mask = 128'h5577ffffffffffffbbbfbfbfbbffbfff;

	lut_sub lut_509 ({sk[106], x5755x, x5756x, x5762x}, x5765x);
	defparam lut_509.LUT_SIZE = 4;
	defparam lut_509.mask = 16'h3f7f;

	lut_sub lut_513 ({sk[107], x270x, x5754x, x5758x, x5759x, x7483x}, x5766x);
	defparam lut_513.LUT_SIZE = 6;
	defparam lut_513.mask = 64'h5f7f5f7fbfffffff;

	lut_sub lut_519 ({sk[108], n_n1082, x77x, x695x, n_n1253, x5788x, x5792x}, x5799x);
	defparam lut_519.LUT_SIZE = 7;
	defparam lut_519.mask = 128'h5577ffffffffffff777777ff77777fff;

	lut_sub lut_524 ({sk[109], n_n876, x123x, x174x, x243x, n_n872, x111x}, x5806x);
	defparam lut_524.LUT_SIZE = 7;
	defparam lut_524.mask = 128'h5577ffffffffffff0357575703ff57ff;

	lut_sub lut_529 ({sk[110], x320x, x5820x, x5821x, x5822x, x5823x}, x5829x);
	defparam lut_529.LUT_SIZE = 6;
	defparam lut_529.mask = 64'h5f7f5f7f7fffffff;

	lut_sub lut_535 ({sk[111], x5862x, x5863x, x5864x, x5865x}, x5870x);
	defparam lut_535.LUT_SIZE = 5;
	defparam lut_535.mask = 32'h5fff7fff;

	lut_sub lut_540 ({sk[112], k, n_n1165, n_n1264, x40x, x5270x, x52x}, x5871x);
	defparam lut_540.LUT_SIZE = 7;
	defparam lut_540.mask = 128'h5577ffffffffffff0303077703030707;

	lut_sub lut_545 ({sk[113], n_n1210, x208x, x351x, x211x, x5825x, x5861x}, x7480x);
	defparam lut_545.LUT_SIZE = 7;
	defparam lut_545.mask = 128'h5577ffffffffffff8800880080000000;

	lut_sub lut_548 ({sk[114], x113x, n_n992, x315x, x81x, x564x, x5893x}, x5903x);
	defparam lut_548.LUT_SIZE = 7;
	defparam lut_548.mask = 128'h5577ffffffffffff777f777f777f77ff;

	lut_sub lut_553 ({sk[115], h, j, k, l, x62x, x7479x}, x5904x);
	defparam lut_553.LUT_SIZE = 7;
	defparam lut_553.mask = 128'h5577ffffffffffffbbabbbaaaaabbbaa;

	lut_sub lut_558 ({sk[116], x5894x, x5895x, x5896x, x5897x}, x5905x);
	defparam lut_558.LUT_SIZE = 5;
	defparam lut_558.mask = 32'h5fff7fff;

	lut_sub lut_563 ({sk[117], h, j, k, l, n_n1187, x51x}, x5906x);
	defparam lut_563.LUT_SIZE = 7;
	defparam lut_563.mask = 128'h5577ffffffffffff1101110000011100;

	lut_sub lut_567 ({sk[118], g, h}, x114x);
	defparam lut_567.LUT_SIZE = 3;
	defparam lut_567.mask = 8'h58;

	lut_sub lut_569 ({sk[119], f, g, h}, n_n1089);
	defparam lut_569.LUT_SIZE = 4;
	defparam lut_569.mask = 16'h3f08;

	lut_sub lut_571 ({sk[120], c, d}, x171x);
	defparam lut_571.LUT_SIZE = 3;
	defparam lut_571.mask = 8'h54;

	lut_sub lut_573 ({sk[121], b, c, d}, n_n842);
	defparam lut_573.LUT_SIZE = 4;
	defparam lut_573.mask = 16'h3f04;

	lut_sub lut_575 ({sk[122], d, e}, x259x);
	defparam lut_575.LUT_SIZE = 3;
	defparam lut_575.mask = 8'h52;

	lut_sub lut_577 ({sk[123], b, d, e}, n_n840);
	defparam lut_577.LUT_SIZE = 4;
	defparam lut_577.mask = 16'h3f02;

	lut_sub lut_579 ({sk[124], e, g, h}, n_n1161);
	defparam lut_579.LUT_SIZE = 4;
	defparam lut_579.mask = 16'h3f20;

	lut_sub lut_581 ({sk[125], f, g}, x112x);
	defparam lut_581.LUT_SIZE = 3;
	defparam lut_581.mask = 8'h51;

	lut_sub lut_583 ({sk[126], f, g, h}, n_n1207);
	defparam lut_583.LUT_SIZE = 4;
	defparam lut_583.mask = 16'h3f02;

	lut_sub lut_585 ({sk[127], c, e}, x256x);
	defparam lut_585.LUT_SIZE = 3;
	defparam lut_585.mask = 8'h51;

	lut_sub lut_587 ({sk[128], b, c, e}, n_n711);
	defparam lut_587.LUT_SIZE = 4;
	defparam lut_587.mask = 16'h3f01;

	lut_sub lut_589 ({sk[129], c, d}, x249x);
	defparam lut_589.LUT_SIZE = 3;
	defparam lut_589.mask = 8'h52;

	lut_sub lut_591 ({sk[130], b, c, d}, n_n713);
	defparam lut_591.LUT_SIZE = 4;
	defparam lut_591.mask = 16'h3f02;

	lut_sub lut_593 ({sk[131], b, d, e}, n_n709);
	defparam lut_593.LUT_SIZE = 4;
	defparam lut_593.mask = 16'h3f04;

	lut_sub lut_595 ({sk[132], g, j, k}, n_n1188);
	defparam lut_595.LUT_SIZE = 4;
	defparam lut_595.mask = 16'h3f02;

	lut_sub lut_597 ({sk[133], e, f, h}, n_n886);
	defparam lut_597.LUT_SIZE = 4;
	defparam lut_597.mask = 16'h3f04;

	lut_sub lut_599 ({sk[134], a, b, c}, n_n920);
	defparam lut_599.LUT_SIZE = 4;
	defparam lut_599.mask = 16'h3f02;

	lut_sub lut_601 ({sk[135], m, n}, n_n1187);
	defparam lut_601.LUT_SIZE = 3;
	defparam lut_601.mask = 8'h52;

	lut_sub lut_603 ({sk[136], a, b, c, m, n}, x38x);
	defparam lut_603.LUT_SIZE = 6;
	defparam lut_603.mask = 64'h5f7f5f7f00000020;

	lut_sub lut_605 ({sk[137], m, n}, n_n1177);
	defparam lut_605.LUT_SIZE = 3;
	defparam lut_605.mask = 8'h54;

	lut_sub lut_607 ({sk[138], i, j, l}, n_n893);
	defparam lut_607.LUT_SIZE = 4;
	defparam lut_607.mask = 16'h3f04;

	lut_sub lut_609 ({sk[139], i, j, l, m, n}, x75x);
	defparam lut_609.LUT_SIZE = 6;
	defparam lut_609.mask = 64'h5f7f5f7f00000400;

	lut_sub lut_611 ({sk[140], i, k, m}, n_n1116);
	defparam lut_611.LUT_SIZE = 4;
	defparam lut_611.mask = 16'h3f02;

	lut_sub lut_613 ({sk[141], i, k, m, n}, x84x);
	defparam lut_613.LUT_SIZE = 5;
	defparam lut_613.mask = 32'h5fff0004;

	lut_sub lut_615 ({sk[142], e, f, g, h, n_n842, n_n713}, x110x);
	defparam lut_615.LUT_SIZE = 7;
	defparam lut_615.mask = 128'h5577ffffffffffff0005030700000303;

	lut_sub lut_619 ({sk[143], i, l, m, n}, x148x);
	defparam lut_619.LUT_SIZE = 5;
	defparam lut_619.mask = 32'h5fff0002;

	lut_sub lut_621 ({sk[144], a, b, c, d, e}, x153x);
	defparam lut_621.LUT_SIZE = 6;
	defparam lut_621.mask = 64'h5f7f5f7f00000026;

	lut_sub lut_624 ({sk[145], i, k, m, n}, x172x);
	defparam lut_624.LUT_SIZE = 5;
	defparam lut_624.mask = 32'h5fff0400;

	lut_sub lut_626 ({sk[146], e, f, g}, n_n1028);
	defparam lut_626.LUT_SIZE = 4;
	defparam lut_626.mask = 16'h3f80;

	lut_sub lut_628 ({sk[147], e, f, g}, x175x);
	defparam lut_628.LUT_SIZE = 4;
	defparam lut_628.mask = 16'h3fa0;

	lut_sub lut_631 ({sk[148], g, i, j, k, l, n_n1187}, x187x);
	defparam lut_631.LUT_SIZE = 7;
	defparam lut_631.mask = 128'h5577ffffffffffff0000000004510504;

	lut_sub lut_637 ({sk[149], b, c, d, e}, x202x);
	defparam lut_637.LUT_SIZE = 5;
	defparam lut_637.mask = 32'h5fff0074;

	lut_sub lut_640 ({sk[150], e, f, g}, n_n1252);
	defparam lut_640.LUT_SIZE = 4;
	defparam lut_640.mask = 16'h3f01;

	lut_sub lut_642 ({sk[151], e, f, g}, n_n940);
	defparam lut_642.LUT_SIZE = 4;
	defparam lut_642.mask = 16'h3f02;

	lut_sub lut_644 ({sk[152], e, f, g}, x229x);
	defparam lut_644.LUT_SIZE = 4;
	defparam lut_644.mask = 16'h3f03;

	lut_sub lut_647 ({sk[153], i, j, l}, n_n933);
	defparam lut_647.LUT_SIZE = 4;
	defparam lut_647.mask = 16'h3f10;

	lut_sub lut_649 ({sk[154], j, l, m, n}, x76x);
	defparam lut_649.LUT_SIZE = 5;
	defparam lut_649.mask = 32'h5fff0400;

	lut_sub lut_651 ({sk[155], f, h, i}, n_n1095);
	defparam lut_651.LUT_SIZE = 4;
	defparam lut_651.mask = 16'h3f04;

	lut_sub lut_653 ({sk[156], f, h, i, x76x}, x298x);
	defparam lut_653.LUT_SIZE = 5;
	defparam lut_653.mask = 32'h5fff0010;

	lut_sub lut_655 ({sk[157], h, k, m, n}, x190x);
	defparam lut_655.LUT_SIZE = 5;
	defparam lut_655.mask = 32'h5fff0002;

	lut_sub lut_657 ({sk[158], g, h, k, m, n}, x306x);
	defparam lut_657.LUT_SIZE = 6;
	defparam lut_657.mask = 64'h5f7f5f7f00020000;

	lut_sub lut_659 ({sk[159], b, e, f}, n_n703);
	defparam lut_659.LUT_SIZE = 4;
	defparam lut_659.mask = 16'h3f04;

	lut_sub lut_661 ({sk[160], b, e, f, g, h, i}, x374x);
	defparam lut_661.LUT_SIZE = 7;
	defparam lut_661.mask = 128'h5577ffffffffffff0000000000400000;

	lut_sub lut_663 ({sk[161], b, c, e, f, g, h}, x393x);
	defparam lut_663.LUT_SIZE = 7;
	defparam lut_663.mask = 128'h5577ffffffffffff00000000000000a0;

	lut_sub lut_666 ({sk[162], m, n}, n_n1165);
	defparam lut_666.LUT_SIZE = 3;
	defparam lut_666.mask = 8'h58;

	lut_sub lut_668 ({sk[163], a, c, d}, n_n904);
	defparam lut_668.LUT_SIZE = 4;
	defparam lut_668.mask = 16'h3f04;

	lut_sub lut_670 ({sk[164], e, f}, x189x);
	defparam lut_670.LUT_SIZE = 3;
	defparam lut_670.mask = 8'h54;

	lut_sub lut_672 ({sk[165], c, e, f}, n_n626);
	defparam lut_672.LUT_SIZE = 4;
	defparam lut_672.mask = 16'h3f04;

	lut_sub lut_674 ({sk[166], b, f}, x196x);
	defparam lut_674.LUT_SIZE = 3;
	defparam lut_674.mask = 8'h54;

	lut_sub lut_676 ({sk[167], b, c, f}, n_n671);
	defparam lut_676.LUT_SIZE = 4;
	defparam lut_676.mask = 16'h3f10;

	lut_sub lut_678 ({sk[168], c, d}, x57x);
	defparam lut_678.LUT_SIZE = 3;
	defparam lut_678.mask = 8'h5e;

	lut_sub lut_681 ({sk[169], c, d, e}, n_n1229);
	defparam lut_681.LUT_SIZE = 4;
	defparam lut_681.mask = 16'h3f01;

	lut_sub lut_683 ({sk[170], f, g, i}, n_n1193);
	defparam lut_683.LUT_SIZE = 4;
	defparam lut_683.mask = 16'h3f02;

	lut_sub lut_685 ({sk[171], h, i, j, k, l}, x181x);
	defparam lut_685.LUT_SIZE = 6;
	defparam lut_685.mask = 64'h5f7f5f7f0c555f0a;

	lut_sub lut_690 ({sk[172], e, f, g, m, n, n_n918}, x388x);
	defparam lut_690.LUT_SIZE = 7;
	defparam lut_690.mask = 128'h5577ffffffffffff0004000400000000;

	lut_sub lut_693 ({sk[173], e, f, g, x111x, x1114x, x1115x}, x1097x);
	defparam lut_693.LUT_SIZE = 7;
	defparam lut_693.mask = 128'h5577ffffffffffff0000000700000000;

	lut_sub lut_696 ({sk[174], n_n713, n_n1177, x101x, n_n1231, x111x, x7494x}, x5199x);
	defparam lut_696.LUT_SIZE = 7;
	defparam lut_696.mask = 128'h5577ffffffffffff222222222222222f;

	lut_sub lut_699 ({sk[175], d, e, g, x45x, n_n698, x111x}, x5200x);
	defparam lut_699.LUT_SIZE = 7;
	defparam lut_699.mask = 128'h5577ffffffffffff0000000000000007;

	lut_sub lut_702 ({sk[176], x75x, x393x, x1110x, x299x, x1114x, x1115x}, x5202x);
	defparam lut_702.LUT_SIZE = 7;
	defparam lut_702.mask = 128'h5577ffffffffffff0707070707ffffff;

	lut_sub lut_707 ({sk[177], x181x, x388x, x1097x, x5199x, x5200x, x5202x}, x5211x);
	defparam lut_707.LUT_SIZE = 7;
	defparam lut_707.mask = 128'h5577ffffffffffff7fff7fff7fffffff;

	lut_sub lut_713 ({sk[178], b, c, e, f, g, h}, x377x);
	defparam lut_713.LUT_SIZE = 7;
	defparam lut_713.mask = 128'h5577ffffffffffff0000000000000050;

	lut_sub lut_716 ({sk[179], b, c, d, e, f, h}, x115x);
	defparam lut_716.LUT_SIZE = 7;
	defparam lut_716.mask = 128'h5577ffffffffffff0000000000000410;

	lut_sub lut_719 ({sk[180], j, k, m}, x21x);
	defparam lut_719.LUT_SIZE = 4;
	defparam lut_719.mask = 16'h3f28;

	lut_sub lut_722 ({sk[181], c, d, f, n_n1166, n_n1204, x295x}, x5225x);
	defparam lut_722.LUT_SIZE = 7;
	defparam lut_722.mask = 128'h5577ffffffffffff0505050705050505;

	lut_sub lut_725 ({sk[182], x297x, n_n1220, n_n1191, x296x, x406x, x5219x}, x5228x);
	defparam lut_725.LUT_SIZE = 7;
	defparam lut_725.mask = 128'h5577ffffffffffff037703770377ffff;

	lut_sub lut_730 ({sk[183], d, n_n1095, n_n973, x78x, x387x, x296x}, x5221x);
	defparam lut_730.LUT_SIZE = 7;
	defparam lut_730.mask = 128'h5577ffffffffffff0000005530303075;

	lut_sub lut_733 ({sk[184], g, h, i, x76x, n_n626, n_n1210}, x5222x);
	defparam lut_733.LUT_SIZE = 7;
	defparam lut_733.mask = 128'h5577ffffffffffff0013110000000000;

	lut_sub lut_737 ({sk[185], a, b, c, d, e, x292x}, x5226x);
	defparam lut_737.LUT_SIZE = 7;
	defparam lut_737.mask = 128'h5577ffffffffffff0000010104000400;

	lut_sub lut_740 ({sk[186], a, x171x, x377x, x115x, x94x, x77x}, x5230x);
	defparam lut_740.LUT_SIZE = 7;
	defparam lut_740.mask = 128'h5577ffffffffffff0555055505553777;

	lut_sub lut_744 ({sk[187], k, l, m, n}, x22x);
	defparam lut_744.LUT_SIZE = 5;
	defparam lut_744.mask = 32'h5fff0020;

	lut_sub lut_746 ({sk[188], j, l, m}, n_n868);
	defparam lut_746.LUT_SIZE = 4;
	defparam lut_746.mask = 16'h3f04;

	lut_sub lut_748 ({sk[189], i, j, l, m}, x31x);
	defparam lut_748.LUT_SIZE = 5;
	defparam lut_748.mask = 32'h5fff1504;

	lut_sub lut_751 ({sk[190], j, k, l, m, n}, x45x);
	defparam lut_751.LUT_SIZE = 6;
	defparam lut_751.mask = 64'h5f7f5f7f00200200;

	lut_sub lut_754 ({sk[191], j, l, m, n}, x54x);
	defparam lut_754.LUT_SIZE = 5;
	defparam lut_754.mask = 32'h5fff0200;

	lut_sub lut_756 ({sk[192], h, k, l}, n_n235);
	defparam lut_756.LUT_SIZE = 4;
	defparam lut_756.mask = 16'h3f02;

	lut_sub lut_758 ({sk[193], h, i, j, k}, x65x);
	defparam lut_758.LUT_SIZE = 5;
	defparam lut_758.mask = 32'h5fff0576;

	lut_sub lut_763 ({sk[194], h, i, j, k, l}, x101x);
	defparam lut_763.LUT_SIZE = 6;
	defparam lut_763.mask = 64'h5f7f5f7f00333f3e;

	lut_sub lut_769 ({sk[195], f, g, h, n, x31x, x54x}, x5253x);
	defparam lut_769.LUT_SIZE = 7;
	defparam lut_769.mask = 128'h5577ffffffffffff0000000000550030;

	lut_sub lut_772 ({sk[196], i, l, m, n, n_n1207, x5253x}, x102x);
	defparam lut_772.LUT_SIZE = 7;
	defparam lut_772.mask = 128'h5577ffffffffffff5555555555555575;

	lut_sub lut_775 ({sk[197], f, g, j, k, l, n_n1187}, x264x);
	defparam lut_775.LUT_SIZE = 7;
	defparam lut_775.mask = 128'h5577ffffffffffff0000000000000400;

	lut_sub lut_777 ({sk[198], i, j, k, l, x112x, n_n1187}, x138x);
	defparam lut_777.LUT_SIZE = 7;
	defparam lut_777.mask = 128'h5577ffffffffffff0010000000110010;

	lut_sub lut_781 ({sk[199], g, h, k, l, m, n}, x1208x);
	defparam lut_781.LUT_SIZE = 7;
	defparam lut_781.mask = 128'h5577ffffffffffff0000004000000000;

	lut_sub lut_783 ({sk[200], g, h, j, k, m, n}, x5088x);
	defparam lut_783.LUT_SIZE = 7;
	defparam lut_783.mask = 128'h5577ffffffffffff0000044000000000;

	lut_sub lut_786 ({sk[201], k, l, m, n}, x58x);
	defparam lut_786.LUT_SIZE = 5;
	defparam lut_786.mask = 32'h5fff0200;

	lut_sub lut_788 ({sk[202], f, g, j, x58x}, x195x);
	defparam lut_788.LUT_SIZE = 5;
	defparam lut_788.mask = 32'h5fff0001;

	lut_sub lut_790 ({sk[203], c, d, e}, n_n973);
	defparam lut_790.LUT_SIZE = 4;
	defparam lut_790.mask = 16'h3f02;

	lut_sub lut_792 ({sk[204], b, c, d, e, f, h}, x1110x);
	defparam lut_792.LUT_SIZE = 7;
	defparam lut_792.mask = 128'h5577ffffffffffff0000000000000020;

	lut_sub lut_794 ({sk[205], a, c, d, e, g}, x258x);
	defparam lut_794.LUT_SIZE = 6;
	defparam lut_794.mask = 64'h5f7f5f7f00000400;

	lut_sub lut_796 ({sk[206], a, c, d, e, g, h}, x297x);
	defparam lut_796.LUT_SIZE = 7;
	defparam lut_796.mask = 128'h5577ffffffffffff0000000000400000;

	lut_sub lut_798 ({sk[207], n_n1193, n_n861, n_n876, n_n864, x14x, x16x}, x125x);
	defparam lut_798.LUT_SIZE = 7;
	defparam lut_798.mask = 128'h5577ffffffffffff000f333f555f777f;

	lut_sub lut_802 ({sk[208], j, k, m, n}, x265x);
	defparam lut_802.LUT_SIZE = 5;
	defparam lut_802.mask = 32'h5fff0020;

	lut_sub lut_804 ({sk[209], j, n_n709, n_n1210, x59x, x48x, x134x}, x5294x);
	defparam lut_804.LUT_SIZE = 7;
	defparam lut_804.mask = 128'h5577ffffffffffff0000000000110051;

	lut_sub lut_807 ({sk[210], j, n_n841, n_n1155, x59x, x192x, x304x}, x5295x);
	defparam lut_807.LUT_SIZE = 7;
	defparam lut_807.mask = 128'h5577ffffffffffff0000000003575757;

	lut_sub lut_811 ({sk[211], j, n_n841, n_n1155, n_n1210, x213x, x5293x}, x5298x);
	defparam lut_811.LUT_SIZE = 7;
	defparam lut_811.mask = 128'h5577ffffffffffff5555555555575757;

	lut_sub lut_815 ({sk[212], k, m, n, n_n1137, x176x, x213x}, x5299x);
	defparam lut_815.LUT_SIZE = 7;
	defparam lut_815.mask = 128'h5577ffffffffffff0037000000000000;

	lut_sub lut_818 ({sk[213], g, h, j, n_n1220, n_n698, n_n1171}, x5291x);
	defparam lut_818.LUT_SIZE = 7;
	defparam lut_818.mask = 128'h5577ffffffffffff0000000700000000;

	lut_sub lut_821 ({sk[214], e, x171x, x265x, n_n1137, n_n1171, n_n1202}, x5292x);
	defparam lut_821.LUT_SIZE = 7;
	defparam lut_821.mask = 128'h5577ffffffffffff0003050700030003;

	lut_sub lut_824 ({sk[215], g, h, j, n_n1036, x48x, x5290x}, x5296x);
	defparam lut_824.LUT_SIZE = 7;
	defparam lut_824.mask = 128'h5577ffffffffffff5555555755555555;

	lut_sub lut_827 ({sk[216], h, i, j, k, n_n1165, x52x}, x5302x);
	defparam lut_827.LUT_SIZE = 7;
	defparam lut_827.mask = 128'h5577ffffffffffff0000000100010000;

	lut_sub lut_830 ({sk[217], h, j, k, n_n1177, x59x, x218x}, x7490x);
	defparam lut_830.LUT_SIZE = 7;
	defparam lut_830.mask = 128'h5577fffffffffffffffffffeffffaafe;

	lut_sub lut_838 ({sk[218], i, j}, x83x);
	defparam lut_838.LUT_SIZE = 3;
	defparam lut_838.mask = 8'h51;

	lut_sub lut_840 ({sk[219], i, j, k}, n_n1217);
	defparam lut_840.LUT_SIZE = 4;
	defparam lut_840.mask = 16'h3f01;

	lut_sub lut_842 ({sk[220], f, g, h}, n_n1201);
	defparam lut_842.LUT_SIZE = 4;
	defparam lut_842.mask = 16'h3f01;

	lut_sub lut_844 ({sk[221], k, m, n}, n_n1220);
	defparam lut_844.LUT_SIZE = 4;
	defparam lut_844.mask = 16'h3f02;

	lut_sub lut_846 ({sk[222], b, c}, x396x);
	defparam lut_846.LUT_SIZE = 3;
	defparam lut_846.mask = 8'h52;

	lut_sub lut_848 ({sk[223], a, b, d}, n_n918);
	defparam lut_848.LUT_SIZE = 4;
	defparam lut_848.mask = 16'h3f01;

	lut_sub lut_850 ({sk[224], a, b, c}, n_n949);
	defparam lut_850.LUT_SIZE = 4;
	defparam lut_850.mask = 16'h3f04;

	lut_sub lut_852 ({sk[225], a, b, c, d}, x15x);
	defparam lut_852.LUT_SIZE = 5;
	defparam lut_852.mask = 32'h5fff0a30;

	lut_sub lut_855 ({sk[226], f, g, h}, n_n1195);
	defparam lut_855.LUT_SIZE = 4;
	defparam lut_855.mask = 16'h3f10;

	lut_sub lut_857 ({sk[227], a, b, d, m, n, n_n1195}, x219x);
	defparam lut_857.LUT_SIZE = 7;
	defparam lut_857.mask = 128'h5577ffffffffffff0000000000000004;

	lut_sub lut_859 ({sk[228], f, g, h, n_n920, n_n1187, n_n918}, x62x);
	defparam lut_859.LUT_SIZE = 7;
	defparam lut_859.mask = 128'h5577ffffffffffff0000001100000003;

	lut_sub lut_862 ({sk[229], a, c, d, e, g, h}, x299x);
	defparam lut_862.LUT_SIZE = 7;
	defparam lut_862.mask = 128'h5577ffffffffffff0000000000200000;

	lut_sub lut_864 ({sk[230], g, h}, x255x);
	defparam lut_864.LUT_SIZE = 3;
	defparam lut_864.mask = 8'h52;

	lut_sub lut_866 ({sk[231], a, c, d}, n_n876);
	defparam lut_866.LUT_SIZE = 4;
	defparam lut_866.mask = 16'h3f02;

	lut_sub lut_868 ({sk[232], a, c, d, e}, x14x);
	defparam lut_868.LUT_SIZE = 5;
	defparam lut_868.mask = 32'h5fff0045;

	lut_sub lut_871 ({sk[233], e, f, x299x, x255x, n_n876, x14x}, x64x);
	defparam lut_871.LUT_SIZE = 7;
	defparam lut_871.mask = 128'h5577ffffffffffff05ff00ff07ff03ff;

	lut_sub lut_875 ({sk[234], a, d, e}, n_n730);
	defparam lut_875.LUT_SIZE = 4;
	defparam lut_875.mask = 16'h3f02;

	lut_sub lut_877 ({sk[235], f, g, h, n_n904, x64x, n_n730}, x82x);
	defparam lut_877.LUT_SIZE = 7;
	defparam lut_877.mask = 128'h5577ffffffffffff3333333333337f33;

	lut_sub lut_881 ({sk[236], f, g, h, n_n920, n_n918, x15x}, x98x);
	defparam lut_881.LUT_SIZE = 7;
	defparam lut_881.mask = 128'h5577ffffffffffff0000330000005f00;

	lut_sub lut_885 ({sk[237], f, g, i}, n_n861);
	defparam lut_885.LUT_SIZE = 4;
	defparam lut_885.mask = 16'h3f20;

	lut_sub lut_887 ({sk[238], e, g, i}, n_n864);
	defparam lut_887.LUT_SIZE = 4;
	defparam lut_887.mask = 16'h3f02;

	lut_sub lut_889 ({sk[239], a, c, d, e}, x16x);
	defparam lut_889.LUT_SIZE = 5;
	defparam lut_889.mask = 32'h5fff0032;

	lut_sub lut_892 ({sk[240], j, l, m, n}, x228x);
	defparam lut_892.LUT_SIZE = 5;
	defparam lut_892.mask = 32'h5fff0002;

	lut_sub lut_894 ({sk[241], e, g, h}, n_n1148);
	defparam lut_894.LUT_SIZE = 4;
	defparam lut_894.mask = 16'h3f01;

	lut_sub lut_896 ({sk[242], a, c, d, e, n_n1201, n_n1196}, x32x);
	defparam lut_896.LUT_SIZE = 7;
	defparam lut_896.mask = 128'h5577ffffffffffff0000000000770030;

	lut_sub lut_900 ({sk[243], a, x249x, n_n1195, x14x, n_n1148, x32x}, x51x);
	defparam lut_900.LUT_SIZE = 7;
	defparam lut_900.mask = 128'h5577ffffffffffff555f555f555f777f;

	lut_sub lut_904 ({sk[244], a, c, d, e, x194x, n_n971}, x50x);
	defparam lut_904.LUT_SIZE = 7;
	defparam lut_904.mask = 128'h5577ffffffffffff0000000005000705;

	lut_sub lut_908 ({sk[245], f, g, h, x297x, x50x, x16x}, x99x);
	defparam lut_908.LUT_SIZE = 7;
	defparam lut_908.mask = 128'h5577ffffffffffff3f3f3f3f3f7f3f3f;

	lut_sub lut_912 ({sk[246], f, g, h, n_n920, n_n918}, x106x);
	defparam lut_912.LUT_SIZE = 6;
	defparam lut_912.mask = 64'h5f7f5f7f05000300;

	lut_sub lut_915 ({sk[247], g, h}, x194x);
	defparam lut_915.LUT_SIZE = 3;
	defparam lut_915.mask = 8'h54;

	lut_sub lut_917 ({sk[248], f, x297x, x106x, x194x, x50x, x16x}, x240x);
	defparam lut_917.LUT_SIZE = 7;
	defparam lut_917.mask = 128'h5577ffffffffffff33ffffff37ffffff;

	lut_sub lut_922 ({sk[249], a, b, e}, n_n698);
	defparam lut_922.LUT_SIZE = 4;
	defparam lut_922.mask = 16'h3f10;

	lut_sub lut_924 ({sk[250], g, h, i}, n_n841);
	defparam lut_924.LUT_SIZE = 4;
	defparam lut_924.mask = 16'h3f04;

	lut_sub lut_926 ({sk[251], g, h, j}, n_n1137);
	defparam lut_926.LUT_SIZE = 4;
	defparam lut_926.mask = 16'h3f01;

	lut_sub lut_928 ({sk[252], f, g, i, x228x, x265x}, x390x);
	defparam lut_928.LUT_SIZE = 6;
	defparam lut_928.mask = 64'h5f7f5f7f00000070;

	lut_sub lut_931 ({sk[253], f, g, h}, n_n1194);
	defparam lut_931.LUT_SIZE = 4;
	defparam lut_931.mask = 16'h3f04;

	lut_sub lut_933 ({sk[254], f, g, h, x15x}, x412x);
	defparam lut_933.LUT_SIZE = 5;
	defparam lut_933.mask = 32'h5fff0010;

	lut_sub lut_935 ({sk[255], f, g, i, x228x, x265x}, x417x);
	defparam lut_935.LUT_SIZE = 6;
	defparam lut_935.mask = 64'h5f7f5f7f00700000;

	lut_sub lut_938 ({sk[256], j, k, l}, n_n996);
	defparam lut_938.LUT_SIZE = 4;
	defparam lut_938.mask = 16'h3f10;

	lut_sub lut_940 ({sk[257], g, h}, x222x);
	defparam lut_940.LUT_SIZE = 3;
	defparam lut_940.mask = 8'h51;

	lut_sub lut_942 ({sk[258], g, h, i}, n_n1155);
	defparam lut_942.LUT_SIZE = 4;
	defparam lut_942.mask = 16'h3f02;

	lut_sub lut_944 ({sk[259], b, e, f}, n_n1171);
	defparam lut_944.LUT_SIZE = 4;
	defparam lut_944.mask = 16'h3f02;

	lut_sub lut_946 ({sk[260], a, b}, x78x);
	defparam lut_946.LUT_SIZE = 3;
	defparam lut_946.mask = 8'h5b;

	lut_sub lut_949 ({sk[261], j, k}, x245x);
	defparam lut_949.LUT_SIZE = 3;
	defparam lut_949.mask = 8'h52;

	lut_sub lut_951 ({sk[262], h, j, k}, n_n617);
	defparam lut_951.LUT_SIZE = 4;
	defparam lut_951.mask = 16'h3f02;

	lut_sub lut_953 ({sk[263], h, k}, x121x);
	defparam lut_953.LUT_SIZE = 3;
	defparam lut_953.mask = 8'h51;

	lut_sub lut_955 ({sk[264], f, g, i}, n_n857);
	defparam lut_955.LUT_SIZE = 4;
	defparam lut_955.mask = 16'h3f10;

	lut_sub lut_957 ({sk[265], g, h, i}, n_n821);
	defparam lut_957.LUT_SIZE = 4;
	defparam lut_957.mask = 16'h3f20;

	lut_sub lut_959 ({sk[266], c, d, e}, n_n700);
	defparam lut_959.LUT_SIZE = 4;
	defparam lut_959.mask = 16'h3f20;

	lut_sub lut_961 ({sk[267], h, i}, x314x);
	defparam lut_961.LUT_SIZE = 3;
	defparam lut_961.mask = 8'h52;

	lut_sub lut_963 ({sk[268], f, h, i}, n_n824);
	defparam lut_963.LUT_SIZE = 4;
	defparam lut_963.mask = 16'h3f02;

	lut_sub lut_965 ({sk[269], x76x, x235x, x5354x, x5355x}, x5363x);
	defparam lut_965.LUT_SIZE = 5;
	defparam lut_965.mask = 32'h5fff777f;

	lut_sub lut_969 ({sk[270], x968x, x5349x, x5356x, x5358x, x5359x}, x5364x);
	defparam lut_969.LUT_SIZE = 6;
	defparam lut_969.mask = 64'h5f7f5f7f7fffffff;

	lut_sub lut_975 ({sk[271], x380x, n_n978, x208x, n_n982, x176x, x5383x}, x5394x);
	defparam lut_975.LUT_SIZE = 7;
	defparam lut_975.mask = 128'h5577ffffffffffff575757ff57ff57ff;

	lut_sub lut_980 ({sk[272], x5379x, x5380x, x5384x, x5385x, x5386x}, x5395x);
	defparam lut_980.LUT_SIZE = 6;
	defparam lut_980.mask = 64'h5f7f5f7f7fffffff;

	lut_sub lut_986 ({sk[273], x961x, n_n1166, x52x, n_n1204, x303x, n_n670}, x5396x);
	defparam lut_986.LUT_SIZE = 7;
	defparam lut_986.mask = 128'h5577ffffffffffff0001000f1111ffff;

	lut_sub lut_991 ({sk[274], x374x, n_n978, x211x, x5377x, x954x, x5382x}, x5397x);
	defparam lut_991.LUT_SIZE = 7;
	defparam lut_991.mask = 128'h5577ffffffffffff77777fff7777ffff;

	lut_sub lut_997 ({sk[275], k, l, m, n}, x142x);
	defparam lut_997.LUT_SIZE = 5;
	defparam lut_997.mask = 32'h5fff0002;

	lut_sub lut_999 ({sk[276], n_n904, n_n698, n_n987, x247x, n_n694, x142x}, x5404x);
	defparam lut_999.LUT_SIZE = 7;
	defparam lut_999.mask = 128'h5577ffffffffffff000011110f001f11;

	lut_sub lut_1002 ({sk[277], x54x, x195x, n_n918, x412x, x29x, x247x}, x7489x);
	defparam lut_1002.LUT_SIZE = 7;
	defparam lut_1002.mask = 128'h5577ffffffffffffffaaccccf0a0c0c0;

	lut_sub lut_1013 ({sk[278], a, b, d, m, n}, x27x);
	defparam lut_1013.LUT_SIZE = 6;
	defparam lut_1013.mask = 64'h5f7f5f7f00000002;

	lut_sub lut_1015 ({sk[279], a, b, c, d}, x29x);
	defparam lut_1015.LUT_SIZE = 5;
	defparam lut_1015.mask = 32'h5fff0a3c;

	lut_sub lut_1019 ({sk[280], b, d, f}, n_n838);
	defparam lut_1019.LUT_SIZE = 4;
	defparam lut_1019.mask = 16'h3f01;

	lut_sub lut_1021 ({sk[281], b, d, e, f}, x30x);
	defparam lut_1021.LUT_SIZE = 5;
	defparam lut_1021.mask = 32'h5fff0045;

	lut_sub lut_1024 ({sk[282], c, d, e, f}, x34x);
	defparam lut_1024.LUT_SIZE = 5;
	defparam lut_1024.mask = 32'h5fff0554;

	lut_sub lut_1028 ({sk[283], a, c, d, m, n}, x129x);
	defparam lut_1028.LUT_SIZE = 6;
	defparam lut_1028.mask = 64'h5f7f5f7f00000200;

	lut_sub lut_1030 ({sk[284], j, k, l, m, n}, x133x);
	defparam lut_1030.LUT_SIZE = 6;
	defparam lut_1030.mask = 64'h5f7f5f7f00000004;

	lut_sub lut_1032 ({sk[285], c, f, g, l, m, n}, x961x);
	defparam lut_1032.LUT_SIZE = 7;
	defparam lut_1032.mask = 128'h5577ffffffffffff0000000000000400;

	lut_sub lut_1034 ({sk[286], f, g, h, i, j, l}, x921x);
	defparam lut_1034.LUT_SIZE = 7;
	defparam lut_1034.mask = 128'h5577ffffffffffff0000000000000100;

	lut_sub lut_1036 ({sk[287], b, c, e}, n_n1053);
	defparam lut_1036.LUT_SIZE = 4;
	defparam lut_1036.mask = 16'h3f20;

	lut_sub lut_1038 ({sk[288], b, c, d}, x36x);
	defparam lut_1038.LUT_SIZE = 4;
	defparam lut_1038.mask = 16'h3f06;

	lut_sub lut_1041 ({sk[289], b, c, d, e}, x210x);
	defparam lut_1041.LUT_SIZE = 5;
	defparam lut_1041.mask = 32'h5fff0a3c;

	lut_sub lut_1045 ({sk[290], a, c, d, e, g, i}, x87x);
	defparam lut_1045.LUT_SIZE = 7;
	defparam lut_1045.mask = 128'h5577ffffffffffff0000000000100100;

	lut_sub lut_1048 ({sk[291], f, g, i, x87x, x14x, x16x}, x238x);
	defparam lut_1048.LUT_SIZE = 7;
	defparam lut_1048.mask = 128'h5577ffffffffffff0f0f0f3f0f0f0f5f;

	lut_sub lut_1052 ({sk[292], f, g, h, m, n}, x257x);
	defparam lut_1052.LUT_SIZE = 6;
	defparam lut_1052.mask = 64'h5f7f5f7f00000020;

	lut_sub lut_1054 ({sk[293], f, g, h, m, n}, x147x);
	defparam lut_1054.LUT_SIZE = 6;
	defparam lut_1054.mask = 64'h5f7f5f7f00000002;

	lut_sub lut_1056 ({sk[294], f, g, h, m, n, x15x}, x291x);
	defparam lut_1056.LUT_SIZE = 7;
	defparam lut_1056.mask = 128'h5577ffffffffffff0000000000000004;

	lut_sub lut_1058 ({sk[295], b, d, e, f, h}, x309x);
	defparam lut_1058.LUT_SIZE = 6;
	defparam lut_1058.mask = 64'h5f7f5f7f00000400;

	lut_sub lut_1060 ({sk[296], g, h, i, x54x}, x380x);
	defparam lut_1060.LUT_SIZE = 5;
	defparam lut_1060.mask = 32'h5fff0004;

	lut_sub lut_1062 ({sk[297], j, k, l, m, n}, x415x);
	defparam lut_1062.LUT_SIZE = 6;
	defparam lut_1062.mask = 64'h5f7f5f7f00000008;

	lut_sub lut_1064 ({sk[298], c, d, e}, n_n1069);
	defparam lut_1064.LUT_SIZE = 4;
	defparam lut_1064.mask = 16'h3f40;

	lut_sub lut_1066 ({sk[299], f, g, h}, n_n1104);
	defparam lut_1066.LUT_SIZE = 4;
	defparam lut_1066.mask = 16'h3f20;

	lut_sub lut_1068 ({sk[300], c, e, f}, n_n1203);
	defparam lut_1068.LUT_SIZE = 4;
	defparam lut_1068.mask = 16'h3f02;

	lut_sub lut_1070 ({sk[301], h, i}, x132x);
	defparam lut_1070.LUT_SIZE = 3;
	defparam lut_1070.mask = 8'h54;

	lut_sub lut_1072 ({sk[302], h, i, j}, n_n1166);
	defparam lut_1072.LUT_SIZE = 4;
	defparam lut_1072.mask = 16'h3f20;

	lut_sub lut_1074 ({sk[303], f, g, h, k, l, n_n1187}, x94x);
	defparam lut_1074.LUT_SIZE = 7;
	defparam lut_1074.mask = 128'h5577ffffffffffff0000000000050004;

	lut_sub lut_1077 ({sk[304], g, h, j, k, l, n_n1177}, x135x);
	defparam lut_1077.LUT_SIZE = 7;
	defparam lut_1077.mask = 128'h5577ffffffffffff0000000000000454;

	lut_sub lut_1080 ({sk[305], a, b, d, e}, x43x);
	defparam lut_1080.LUT_SIZE = 5;
	defparam lut_1080.mask = 32'h5fff0d00;

	lut_sub lut_1083 ({sk[306], b, c, e, x184x, x77x, x117x}, x5462x);
	defparam lut_1083.LUT_SIZE = 7;
	defparam lut_1083.mask = 128'h5577ffffffffffff0303035703030303;

	lut_sub lut_1086 ({sk[307], f, h, i}, n_n662);
	defparam lut_1086.LUT_SIZE = 4;
	defparam lut_1086.mask = 16'h3f40;

	lut_sub lut_1088 ({sk[308], b, d, e, k, m, n}, x126x);
	defparam lut_1088.LUT_SIZE = 7;
	defparam lut_1088.mask = 128'h5577ffffffffffff0000000000040000;

	lut_sub lut_1090 ({sk[309], c, d, e, f, x132x, x296x}, x874x);
	defparam lut_1090.LUT_SIZE = 7;
	defparam lut_1090.mask = 128'h5577ffffffffffff0000000100010000;

	lut_sub lut_1093 ({sk[310], j, x309x, x77x, n_n1036, x5458x, x5460x}, x5465x);
	defparam lut_1093.LUT_SIZE = 7;
	defparam lut_1093.mask = 128'h5577ffffffffffff777777ff77777fff;

	lut_sub lut_1098 ({sk[311], n_n842, n_n1177, n_n1252, n_n235, x195x, x43x}, x5473x);
	defparam lut_1098.LUT_SIZE = 7;
	defparam lut_1098.mask = 128'h5577ffffffffffff111111111111111f;

	lut_sub lut_1101 ({sk[312], a, b, c, d, f, x44x}, x5474x);
	defparam lut_1101.LUT_SIZE = 7;
	defparam lut_1101.mask = 128'h5577ffffffffffff0000000001011000;

	lut_sub lut_1104 ({sk[313], i, j, k, l}, x39x);
	defparam lut_1104.LUT_SIZE = 5;
	defparam lut_1104.mask = 32'h5fff2532;

	lut_sub lut_1109 ({sk[314], i, j, k, l}, x74x);
	defparam lut_1109.LUT_SIZE = 5;
	defparam lut_1109.mask = 32'h5fff2d36;

	lut_sub lut_1116 ({sk[315], h, j}, x146x);
	defparam lut_1116.LUT_SIZE = 3;
	defparam lut_1116.mask = 8'h52;

	lut_sub lut_1118 ({sk[316], h, i, j, l}, x20x);
	defparam lut_1118.LUT_SIZE = 5;
	defparam lut_1118.mask = 32'h5fff0572;

	lut_sub lut_1122 ({sk[317], d, f, g, l, x146x, x20x}, x92x);
	defparam lut_1122.LUT_SIZE = 7;
	defparam lut_1122.mask = 128'h5577ffffffffffff0000035500000000;

	lut_sub lut_1125 ({sk[318], a, m, n}, x120x);
	defparam lut_1125.LUT_SIZE = 4;
	defparam lut_1125.mask = 16'h3f02;

	lut_sub lut_1127 ({sk[319], e, f, g, h, x190x, x22x}, x151x);
	defparam lut_1127.LUT_SIZE = 7;
	defparam lut_1127.mask = 128'h5577ffffffffffff0000000000003705;

	lut_sub lut_1130 ({sk[320], i, j, k, l}, x183x);
	defparam lut_1130.LUT_SIZE = 5;
	defparam lut_1130.mask = 32'h5fff2536;

	lut_sub lut_1136 ({sk[321], f, g, h}, n_n971);
	defparam lut_1136.LUT_SIZE = 4;
	defparam lut_1136.mask = 16'h3f40;

	lut_sub lut_1138 ({sk[322], b, c, d, e, n_n1195, n_n971}, x184x);
	defparam lut_1138.LUT_SIZE = 7;
	defparam lut_1138.mask = 128'h5577ffffffffffff0000000000330707;

	lut_sub lut_1142 ({sk[323], d, f, g, m, n, n_n920}, x223x);
	defparam lut_1142.LUT_SIZE = 7;
	defparam lut_1142.mask = 128'h5577ffffffffffff0000000400000000;

	lut_sub lut_1144 ({sk[324], f, g, h, i}, x230x);
	defparam lut_1144.LUT_SIZE = 5;
	defparam lut_1144.mask = 32'h5fff4404;

	lut_sub lut_1147 ({sk[325], f, g, i, x102x, x228x, x265x}, x239x);
	defparam lut_1147.LUT_SIZE = 7;
	defparam lut_1147.mask = 128'h5577ffffffffffff0f0f0f0f0f0f7f0f;

	lut_sub lut_1151 ({sk[326], i, j, k, m}, x49x);
	defparam lut_1151.LUT_SIZE = 5;
	defparam lut_1151.mask = 32'h5fff2a28;

	lut_sub lut_1155 ({sk[327], j, k, m, n}, x113x);
	defparam lut_1155.LUT_SIZE = 5;
	defparam lut_1155.mask = 32'h5fff0200;

	lut_sub lut_1157 ({sk[328], j, k, l, m, n}, x33x);
	defparam lut_1157.LUT_SIZE = 6;
	defparam lut_1157.mask = 64'h5f7f5f7f00220020;

	lut_sub lut_1160 ({sk[329], b, c, e, f}, x93x);
	defparam lut_1160.LUT_SIZE = 5;
	defparam lut_1160.mask = 32'h5fff0d22;

	lut_sub lut_1164 ({sk[330], f, g, h, n_n920, n_n918}, x156x);
	defparam lut_1164.LUT_SIZE = 6;
	defparam lut_1164.mask = 64'h5f7f5f7f00500030;

	lut_sub lut_1167 ({sk[331], f, g, i, n_n920, n_n918}, x203x);
	defparam lut_1167.LUT_SIZE = 6;
	defparam lut_1167.mask = 64'h5f7f5f7f00050003;

	lut_sub lut_1170 ({sk[332], b, d, e, f, g, h}, x841x);
	defparam lut_1170.LUT_SIZE = 7;
	defparam lut_1170.mask = 128'h5577ffffffffffff0000000000000200;

	lut_sub lut_1172 ({sk[333], b, c, d, e, g, h}, x5557x);
	defparam lut_1172.LUT_SIZE = 7;
	defparam lut_1172.mask = 128'h5577ffffffffffff0000000002022000;

	lut_sub lut_1175 ({sk[334], i, k}, x246x);
	defparam lut_1175.LUT_SIZE = 3;
	defparam lut_1175.mask = 8'h51;

	lut_sub lut_1177 ({sk[335], f, g, i}, n_n1228);
	defparam lut_1177.LUT_SIZE = 4;
	defparam lut_1177.mask = 16'h3f01;

	lut_sub lut_1179 ({sk[336], f, g, i, x15x}, x402x);
	defparam lut_1179.LUT_SIZE = 5;
	defparam lut_1179.mask = 32'h5fff0001;

	lut_sub lut_1181 ({sk[337], c, d}, x131x);
	defparam lut_1181.LUT_SIZE = 3;
	defparam lut_1181.mask = 8'h58;

	lut_sub lut_1183 ({sk[338], c, d, f}, n_n1138);
	defparam lut_1183.LUT_SIZE = 4;
	defparam lut_1183.mask = 16'h3f80;

	lut_sub lut_1185 ({sk[339], j, k, l}, n_n1159);
	defparam lut_1185.LUT_SIZE = 4;
	defparam lut_1185.mask = 16'h3f80;

	lut_sub lut_1187 ({sk[340], k, l, m, n}, n_n978);
	defparam lut_1187.LUT_SIZE = 5;
	defparam lut_1187.mask = 32'h5fff0004;

	lut_sub lut_1189 ({sk[341], d, f, j, l, m, n}, x5632x);
	defparam lut_1189.LUT_SIZE = 7;
	defparam lut_1189.mask = 128'h5577ffffffffffff0000000000000200;

	lut_sub lut_1191 ({sk[342], g, h, i}, n_n992);
	defparam lut_1191.LUT_SIZE = 4;
	defparam lut_1191.mask = 16'h3f01;

	lut_sub lut_1193 ({sk[343], k, m, n}, n_n1222);
	defparam lut_1193.LUT_SIZE = 4;
	defparam lut_1193.mask = 16'h3f20;

	lut_sub lut_1195 ({sk[344], d, e, f}, n_n1260);
	defparam lut_1195.LUT_SIZE = 4;
	defparam lut_1195.mask = 16'h3f01;

	lut_sub lut_1197 ({sk[345], e, f, g}, n_n987);
	defparam lut_1197.LUT_SIZE = 4;
	defparam lut_1197.mask = 16'h3f04;

	lut_sub lut_1199 ({sk[346], h, i, j}, n_n1085);
	defparam lut_1199.LUT_SIZE = 4;
	defparam lut_1199.mask = 16'h3f02;

	lut_sub lut_1201 ({sk[347], b, c, d, k, l, n_n1177}, x370x);
	defparam lut_1201.LUT_SIZE = 7;
	defparam lut_1201.mask = 128'h5577ffffffffffff0000001000000000;

	lut_sub lut_1203 ({sk[348], c, d, e}, n_n975);
	defparam lut_1203.LUT_SIZE = 4;
	defparam lut_1203.mask = 16'h3f10;

	lut_sub lut_1205 ({sk[349], i, j, k, l, m, n}, x308x);
	defparam lut_1205.LUT_SIZE = 7;
	defparam lut_1205.mask = 128'h5577ffffffffffff0000000008000000;

	lut_sub lut_1207 ({sk[350], g, h, i}, n_n1142);
	defparam lut_1207.LUT_SIZE = 4;
	defparam lut_1207.mask = 16'h3f10;

	lut_sub lut_1209 ({sk[351], a, b, c, m, n}, x193x);
	defparam lut_1209.LUT_SIZE = 6;
	defparam lut_1209.mask = 64'h5f7f5f7f00020000;

	lut_sub lut_1211 ({sk[352], d, l, x189x, x245x, n_n1142, x193x}, x779x);
	defparam lut_1211.LUT_SIZE = 7;
	defparam lut_1211.mask = 128'h5577ffffffffffff0000000000000001;

	lut_sub lut_1213 ({sk[353], l, m, n}, n_n1204);
	defparam lut_1213.LUT_SIZE = 4;
	defparam lut_1213.mask = 16'h3f08;

	lut_sub lut_1215 ({sk[354], c, f, g, h, x53x, x382x}, n_n2602);
	defparam lut_1215.LUT_SIZE = 7;
	defparam lut_1215.mask = 128'h5577ffffffffffff0000001000000000;

	lut_sub lut_1217 ({sk[355], k, l, m, n}, n_n982);
	defparam lut_1217.LUT_SIZE = 5;
	defparam lut_1217.mask = 32'h5fff0400;

	lut_sub lut_1219 ({sk[356], b, c, d, e, f, g}, x372x);
	defparam lut_1219.LUT_SIZE = 7;
	defparam lut_1219.mask = 128'h5577ffffffffffff0000000000000040;

	lut_sub lut_1221 ({sk[357], h, i, m, n}, x226x);
	defparam lut_1221.LUT_SIZE = 5;
	defparam lut_1221.mask = 32'h5fff8000;

	lut_sub lut_1223 ({sk[358], g, h, i, m, n}, x367x);
	defparam lut_1223.LUT_SIZE = 6;
	defparam lut_1223.mask = 64'h5f7f5f7f80000000;

	lut_sub lut_1225 ({sk[359], i, j, k, l, m, n}, x141x);
	defparam lut_1225.LUT_SIZE = 7;
	defparam lut_1225.mask = 128'h5577ffffffffffff0000000000000008;

	lut_sub lut_1227 ({sk[360], l, m, n}, n_n1190);
	defparam lut_1227.LUT_SIZE = 4;
	defparam lut_1227.mask = 16'h3f80;

	lut_sub lut_1229 ({sk[361], k, m, n}, n_n1202);
	defparam lut_1229.LUT_SIZE = 4;
	defparam lut_1229.mask = 16'h3f80;

	lut_sub lut_1231 ({sk[362], f, g, h}, n_n1039);
	defparam lut_1231.LUT_SIZE = 4;
	defparam lut_1231.mask = 16'h3f80;

	lut_sub lut_1233 ({sk[363], c, d, e, f, g, h}, x5657x);
	defparam lut_1233.LUT_SIZE = 7;
	defparam lut_1233.mask = 128'h5577ffffffffffff0000002000000000;

	lut_sub lut_1235 ({sk[364], d, e}, x90x);
	defparam lut_1235.LUT_SIZE = 3;
	defparam lut_1235.mask = 8'h51;

	lut_sub lut_1237 ({sk[365], c, f, g, h, x382x, x90x}, n_n2493);
	defparam lut_1237.LUT_SIZE = 7;
	defparam lut_1237.mask = 128'h5577ffffffffffff0010000000000000;

	lut_sub lut_1239 ({sk[366], a, b, c, m, n}, x145x);
	defparam lut_1239.LUT_SIZE = 6;
	defparam lut_1239.mask = 64'h5f7f5f7f00000002;

	lut_sub lut_1241 ({sk[367], j, k, l, n_n992, n_n1260, x145x}, x764x);
	defparam lut_1241.LUT_SIZE = 7;
	defparam lut_1241.mask = 128'h5577ffffffffffff0000000000000001;

	lut_sub lut_1243 ({sk[368], h, i, j}, n_n1264);
	defparam lut_1243.LUT_SIZE = 4;
	defparam lut_1243.mask = 16'h3f01;

	lut_sub lut_1245 ({sk[369], b, c, d}, n_n1253);
	defparam lut_1245.LUT_SIZE = 4;
	defparam lut_1245.mask = 16'h3f01;

	lut_sub lut_1247 ({sk[370], h, i}, x122x);
	defparam lut_1247.LUT_SIZE = 3;
	defparam lut_1247.mask = 8'h5e;

	lut_sub lut_1250 ({sk[371], a, c, e}, n_n761);
	defparam lut_1250.LUT_SIZE = 4;
	defparam lut_1250.mask = 16'h3f01;

	lut_sub lut_1252 ({sk[372], e, f, g}, n_n1231);
	defparam lut_1252.LUT_SIZE = 4;
	defparam lut_1252.mask = 16'h3f10;

	lut_sub lut_1254 ({sk[373], a, b, c}, n_n997);
	defparam lut_1254.LUT_SIZE = 4;
	defparam lut_1254.mask = 16'h3f10;

	lut_sub lut_1256 ({sk[374], a, c, d, n_n1187, n_n1231, x181x}, x746x);
	defparam lut_1256.LUT_SIZE = 7;
	defparam lut_1256.mask = 128'h5577ffffffffffff0000000000000001;

	lut_sub lut_1258 ({sk[375], f, g, h, n_n1069, x382x, x308x}, x5684x);
	defparam lut_1258.LUT_SIZE = 7;
	defparam lut_1258.mask = 128'h5577ffffffffffff0000000000000305;

	lut_sub lut_1261 ({sk[376], f, g, x46x, x57x, x74x, x145x}, x5686x);
	defparam lut_1261.LUT_SIZE = 7;
	defparam lut_1261.mask = 128'h5577ffffffffffff0050105000000000;

	lut_sub lut_1264 ({sk[377], g, x46x, x189x, x57x, x120x, x750x}, x5687x);
	defparam lut_1264.LUT_SIZE = 7;
	defparam lut_1264.mask = 128'h5577ffffffffffff5555557555555555;

	lut_sub lut_1267 ({sk[378], g, h, k, l, m, n}, x44x);
	defparam lut_1267.LUT_SIZE = 7;
	defparam lut_1267.mask = 128'h5577ffffffffffff0000002200000020;

	lut_sub lut_1270 ({sk[379], g, h, k, l, n_n1187, x189x}, x108x);
	defparam lut_1270.LUT_SIZE = 7;
	defparam lut_1270.mask = 128'h5577ffffffffffff0000001100000010;

	lut_sub lut_1273 ({sk[380], e, g, h, n, x31x}, x1116x);
	defparam lut_1273.LUT_SIZE = 6;
	defparam lut_1273.mask = 64'h5f7f5f7f00000004;

	lut_sub lut_1275 ({sk[381], e, g, h, x148x, x54x, x1116x}, x123x);
	defparam lut_1275.LUT_SIZE = 7;
	defparam lut_1275.mask = 128'h5577ffffffffffff5555555555775f55;

	lut_sub lut_1279 ({sk[382], e, g, h, k, m, n}, x387x);
	defparam lut_1279.LUT_SIZE = 7;
	defparam lut_1279.mask = 128'h5577ffffffffffff0000000000020000;

	lut_sub lut_1281 ({sk[383], e, g, h, k, l, n_n1187}, x174x);
	defparam lut_1281.LUT_SIZE = 7;
	defparam lut_1281.mask = 128'h5577ffffffffffff0000000000050004;

	lut_sub lut_1284 ({sk[384], e, g, i, x228x, x265x, x33x}, x182x);
	defparam lut_1284.LUT_SIZE = 7;
	defparam lut_1284.mask = 128'h5577ffffffffffff0000000000003f55;

	lut_sub lut_1288 ({sk[385], f, g, h, k, l, n_n1187}, x200x);
	defparam lut_1288.LUT_SIZE = 7;
	defparam lut_1288.mask = 128'h5577ffffffffffff0005000400000000;

	lut_sub lut_1291 ({sk[386], f, g, h, n}, x385x);
	defparam lut_1291.LUT_SIZE = 5;
	defparam lut_1291.mask = 32'h5fff0200;

	lut_sub lut_1293 ({sk[387], x148x, x31x, x54x, n_n1104, n_n971, x385x}, x243x);
	defparam lut_1293.LUT_SIZE = 7;
	defparam lut_1293.mask = 128'h5577ffffffffffff003355770f3f5f7f;

	lut_sub lut_1297 ({sk[388], k, l, m}, n_n1118);
	defparam lut_1297.LUT_SIZE = 4;
	defparam lut_1297.mask = 16'h3f80;

	lut_sub lut_1299 ({sk[389], g, j, k, l, m, n}, x247x);
	defparam lut_1299.LUT_SIZE = 7;
	defparam lut_1299.mask = 128'h5577ffffffffffff0000000000000200;

	lut_sub lut_1301 ({sk[390], e, g, i, x22x, n_n876, x247x}, x270x);
	defparam lut_1301.LUT_SIZE = 7;
	defparam lut_1301.mask = 128'h5577ffffffffffff0000000011111113;

	lut_sub lut_1304 ({sk[391], e, g, h}, n_n1082);
	defparam lut_1304.LUT_SIZE = 4;
	defparam lut_1304.mask = 16'h3f04;

	lut_sub lut_1306 ({sk[392], h, i}, x37x);
	defparam lut_1306.LUT_SIZE = 3;
	defparam lut_1306.mask = 8'h57;

	lut_sub lut_1309 ({sk[393], g, h, i}, x407x);
	defparam lut_1309.LUT_SIZE = 4;
	defparam lut_1309.mask = 16'h3f80;

	lut_sub lut_1311 ({sk[394], a, d, e}, n_n872);
	defparam lut_1311.LUT_SIZE = 4;
	defparam lut_1311.mask = 16'h3f04;

	lut_sub lut_1313 ({sk[395], i, j, k}, n_n977);
	defparam lut_1313.LUT_SIZE = 4;
	defparam lut_1313.mask = 16'h3f20;

	lut_sub lut_1315 ({sk[396], j, k, l}, x55x);
	defparam lut_1315.LUT_SIZE = 4;
	defparam lut_1315.mask = 16'h3f24;

	lut_sub lut_1318 ({sk[397], i, j, k, l}, x18x);
	defparam lut_1318.LUT_SIZE = 5;
	defparam lut_1318.mask = 32'h5fff0032;

	lut_sub lut_1321 ({sk[398], n_n1161, x75x, n_n940, x129x, n_n988, n_n942}, x5738x);
	defparam lut_1321.LUT_SIZE = 7;
	defparam lut_1321.mask = 128'h5577ffffffffffff0005000500053337;

	lut_sub lut_1324 ({sk[399], n_n1252, x129x, x74x, x223x, x55x, x20x}, x7484x);
	defparam lut_1324.LUT_SIZE = 7;
	defparam lut_1324.mask = 128'h5577fffffffffffffcfcfcfcfcfca800;

	lut_sub lut_1331 ({sk[400], k, m, n}, n_n1210);
	defparam lut_1331.LUT_SIZE = 4;
	defparam lut_1331.mask = 16'h3f04;

	lut_sub lut_1333 ({sk[401], e, g, h, x84x, n_n988, x77x}, x5755x);
	defparam lut_1333.LUT_SIZE = 7;
	defparam lut_1333.mask = 128'h5577ffffffffffff0000031100000000;

	lut_sub lut_1336 ({sk[402], n_n842, x76x, n_n841, n_n857, x33x, n_n872}, x5756x);
	defparam lut_1336.LUT_SIZE = 7;
	defparam lut_1336.mask = 128'h5577ffffffffffff01010101010101ff;

	lut_sub lut_1339 ({sk[403], n, x49x, n_n988, x695x, x696x, n_n1196}, x5762x);
	defparam lut_1339.LUT_SIZE = 7;
	defparam lut_1339.mask = 128'h5577ffffffffffff0000000000003f7f;

	lut_sub lut_1343 ({sk[404], a, x53x, n_n857, x113x, x414x, x247x}, x5754x);
	defparam lut_1343.LUT_SIZE = 7;
	defparam lut_1343.mask = 128'h5577ffffffffffff0303030303030357;

	lut_sub lut_1346 ({sk[405], b, c, d, e, x76x, n_n1095}, x5758x);
	defparam lut_1346.LUT_SIZE = 7;
	defparam lut_1346.mask = 128'h5577ffffffffffff0000001100100010;

	lut_sub lut_1349 ({sk[406], a, x249x, x228x, n_n864, x697x, x266x}, x5759x);
	defparam lut_1349.LUT_SIZE = 7;
	defparam lut_1349.mask = 128'h5577ffffffffffff113311331133153f;

	lut_sub lut_1354 ({sk[407], i, x114x, x84x, x298x, n_n838, x167x}, x7483x);
	defparam lut_1354.LUT_SIZE = 7;
	defparam lut_1354.mask = 128'h5577ffffffffffffffaaffaaffaafca8;

	lut_sub lut_1363 ({sk[408], e, f, g, n_n1253, x283x, x301x}, x670x);
	defparam lut_1363.LUT_SIZE = 7;
	defparam lut_1363.mask = 128'h5577ffffffffffff0000000000000001;

	lut_sub lut_1365 ({sk[409], h, x112x, n_n1069, n_n977, x302x, x308x}, x5771x);
	defparam lut_1365.LUT_SIZE = 7;
	defparam lut_1365.mask = 128'h5577ffffffffffff0000030300000055;

	lut_sub lut_1368 ({sk[410], l, x382x, x5627x, n_n1210, x283x, x372x}, x5772x);
	defparam lut_1368.LUT_SIZE = 7;
	defparam lut_1368.mask = 128'h5577ffffffffffff000000ff010101ff;

	lut_sub lut_1371 ({sk[411], n_n978, x382x, x5657x, n_n987, n_n988, x283x}, x5773x);
	defparam lut_1371.LUT_SIZE = 7;
	defparam lut_1371.mask = 128'h5577ffffffffffff000000ff010101ff;

	lut_sub lut_1374 ({sk[412], b, c, d}, n_n988);
	defparam lut_1374.LUT_SIZE = 4;
	defparam lut_1374.mask = 16'h3f10;

	lut_sub lut_1376 ({sk[413], k, l, m, n}, x77x);
	defparam lut_1376.LUT_SIZE = 5;
	defparam lut_1376.mask = 32'h5fff0040;

	lut_sub lut_1378 ({sk[414], f, h, i}, x59x);
	defparam lut_1378.LUT_SIZE = 4;
	defparam lut_1378.mask = 16'h3f06;

	lut_sub lut_1381 ({sk[415], f, h, i, j}, x89x);
	defparam lut_1381.LUT_SIZE = 5;
	defparam lut_1381.mask = 32'h5fff003e;

	lut_sub lut_1385 ({sk[416], a, b, c, m, n}, x111x);
	defparam lut_1385.LUT_SIZE = 6;
	defparam lut_1385.mask = 64'h5f7f5f7f00000200;

	lut_sub lut_1387 ({sk[417], f, h, k, l, m, n}, x893x);
	defparam lut_1387.LUT_SIZE = 7;
	defparam lut_1387.mask = 128'h5577ffffffffffff0000000000000040;

	lut_sub lut_1389 ({sk[418], f, h, j}, n_n823);
	defparam lut_1389.LUT_SIZE = 4;
	defparam lut_1389.mask = 16'h3f01;

	lut_sub lut_1391 ({sk[419], k, m, n, x893x, n_n823}, x117x);
	defparam lut_1391.LUT_SIZE = 6;
	defparam lut_1391.mask = 64'h5f7f5f7f37333333;

	lut_sub lut_1394 ({sk[420], a, d, e, f, g, i}, x697x);
	defparam lut_1394.LUT_SIZE = 7;
	defparam lut_1394.mask = 128'h5577ffffffffffff0000000000200000;

	lut_sub lut_1396 ({sk[421], b, d, e, f, g, h}, x695x);
	defparam lut_1396.LUT_SIZE = 7;
	defparam lut_1396.mask = 128'h5577ffffffffffff0000000000000010;

	lut_sub lut_1398 ({sk[422], b, c, d, e, g, h}, x696x);
	defparam lut_1398.LUT_SIZE = 7;
	defparam lut_1398.mask = 128'h5577ffffffffffff0000000000000004;

	lut_sub lut_1400 ({sk[423], g, h, j}, n_n820);
	defparam lut_1400.LUT_SIZE = 4;
	defparam lut_1400.mask = 16'h3f02;

	lut_sub lut_1402 ({sk[424], g, h, i, j}, x164x);
	defparam lut_1402.LUT_SIZE = 5;
	defparam lut_1402.mask = 32'h5fff003e;

	lut_sub lut_1406 ({sk[425], b, c, d, e, x114x, n_n1104}, x167x);
	defparam lut_1406.LUT_SIZE = 7;
	defparam lut_1406.mask = 128'h5577ffffffffffff0000000000050007;

	lut_sub lut_1409 ({sk[426], i, k}, x386x);
	defparam lut_1409.LUT_SIZE = 3;
	defparam lut_1409.mask = 8'h58;

	lut_sub lut_1411 ({sk[427], b, x53x, n_n1171, x70x, n_n992, x155x}, x320x);
	defparam lut_1411.LUT_SIZE = 7;
	defparam lut_1411.mask = 128'h5577ffffffffffff0507050705070707;

	lut_sub lut_1415 ({sk[428], n_n671, n_n700, n_n1264, n_n1036, n_n1227, x290x}, x5820x);
	defparam lut_1415.LUT_SIZE = 7;
	defparam lut_1415.mask = 128'h5577ffffffffffff00001111000f111f;

	lut_sub lut_1418 ({sk[429], k, n_n709, n_n1177, n_n1053, n_n820, x231x}, x5821x);
	defparam lut_1418.LUT_SIZE = 7;
	defparam lut_1418.mask = 128'h5577ffffffffffff0000000000030057;

	lut_sub lut_1421 ({sk[430], i, n_n840, x194x, n_n824, n_n1210, x48x}, x5822x);
	defparam lut_1421.LUT_SIZE = 7;
	defparam lut_1421.mask = 128'h5577ffffffffffff0011031300000303;

	lut_sub lut_1424 ({sk[431], g, j, k, x30x, x403x, x410x}, x5823x);
	defparam lut_1424.LUT_SIZE = 7;
	defparam lut_1424.mask = 128'h5577ffffffffffff0303030303570303;

	lut_sub lut_1427 ({sk[432], h, i, j, k}, x40x);
	defparam lut_1427.LUT_SIZE = 5;
	defparam lut_1427.mask = 32'h5fff0054;

	lut_sub lut_1430 ({sk[433], b, d, e, k, m, n}, x192x);
	defparam lut_1430.LUT_SIZE = 7;
	defparam lut_1430.mask = 128'h5577ffffffffffff0000000000000400;

	lut_sub lut_1432 ({sk[434], g, h, j, n_n703, n_n1171, n_n838}, x208x);
	defparam lut_1432.LUT_SIZE = 7;
	defparam lut_1432.mask = 128'h5577ffffffffffff00005f0000003300;

	lut_sub lut_1436 ({sk[435], b, c, f, g, m, n}, x5270x);
	defparam lut_1436.LUT_SIZE = 7;
	defparam lut_1436.mask = 128'h5577ffffffffffff0000004400000040;

	lut_sub lut_1439 ({sk[436], c, d, e, f, g}, x52x);
	defparam lut_1439.LUT_SIZE = 6;
	defparam lut_1439.mask = 64'h5f7f5f7f00333f3e;

	lut_sub lut_1445 ({sk[437], f, g}, x310x);
	defparam lut_1445.LUT_SIZE = 3;
	defparam lut_1445.mask = 8'h52;

	lut_sub lut_1447 ({sk[438], c, m, n, x196x, x52x, x310x}, x218x);
	defparam lut_1447.LUT_SIZE = 7;
	defparam lut_1447.mask = 128'h5577ffffffffffff33000000335f0000;

	lut_sub lut_1451 ({sk[439], j, k, m, n}, x70x);
	defparam lut_1451.LUT_SIZE = 5;
	defparam lut_1451.mask = 32'h5fff0040;

	lut_sub lut_1453 ({sk[440], g, j, k, l, m, n}, x266x);
	defparam lut_1453.LUT_SIZE = 7;
	defparam lut_1453.mask = 128'h5577ffffffffffff0000000000200000;

	lut_sub lut_1455 ({sk[441], k, m, n}, n_n1191);
	defparam lut_1455.LUT_SIZE = 4;
	defparam lut_1455.mask = 16'h3f08;

	lut_sub lut_1457 ({sk[442], c, d, e, k, m, n}, x304x);
	defparam lut_1457.LUT_SIZE = 7;
	defparam lut_1457.mask = 128'h5577ffffffffffff0000080000000000;

	lut_sub lut_1459 ({sk[443], a, c, d, e, g, i}, x414x);
	defparam lut_1459.LUT_SIZE = 7;
	defparam lut_1459.mask = 128'h5577ffffffffffff0000000000000100;

	lut_sub lut_1461 ({sk[444], n_n857, x113x, n_n1228, x14x, x414x, x16x}, x351x);
	defparam lut_1461.LUT_SIZE = 7;
	defparam lut_1461.mask = 128'h5577ffffffffffff0000337700003f7f;

	lut_sub lut_1465 ({sk[445], j, k, m}, n_n1227);
	defparam lut_1465.LUT_SIZE = 4;
	defparam lut_1465.mask = 16'h3f08;

	lut_sub lut_1467 ({sk[446], g, h, i, n, n_n1227}, x403x);
	defparam lut_1467.LUT_SIZE = 6;
	defparam lut_1467.mask = 64'h5f7f5f7f00010000;

	lut_sub lut_1469 ({sk[447], k, m, n}, n_n1036);
	defparam lut_1469.LUT_SIZE = 4;
	defparam lut_1469.mask = 16'h3f40;

	lut_sub lut_1471 ({sk[448], g, h, k}, n_n816);
	defparam lut_1471.LUT_SIZE = 4;
	defparam lut_1471.mask = 16'h3f10;

	lut_sub lut_1473 ({sk[449], b, c, d, e, f}, x48x);
	defparam lut_1473.LUT_SIZE = 6;
	defparam lut_1473.mask = 64'h5f7f5f7f00004577;

	lut_sub lut_1477 ({sk[450], g, h, i, n_n711, n_n1171, x30x}, x235x);
	defparam lut_1477.LUT_SIZE = 7;
	defparam lut_1477.mask = 128'h5577ffffffffffff005f000000330000;

	lut_sub lut_1481 ({sk[451], g, h, i, n}, x290x);
	defparam lut_1481.LUT_SIZE = 5;
	defparam lut_1481.mask = 32'h5fff0002;

	lut_sub lut_1483 ({sk[452], a, b, e, m, n}, x315x);
	defparam lut_1483.LUT_SIZE = 6;
	defparam lut_1483.mask = 64'h5f7f5f7f00020000;

	lut_sub lut_1485 ({sk[453], b, d, e, f, h, i}, x155x);
	defparam lut_1485.LUT_SIZE = 7;
	defparam lut_1485.mask = 128'h5577ffffffffffff0000000000100100;

	lut_sub lut_1488 ({sk[454], g, h, k, x171x, n_n1190, x529x}, x5950x);
	defparam lut_1488.LUT_SIZE = 7;
	defparam lut_1488.mask = 128'h5577ffffffffffff5755555555555555;

	lut_sub lut_1491 ({sk[455], c, d, g, h, n_n662, x282x}, x5951x);
	defparam lut_1491.LUT_SIZE = 7;
	defparam lut_1491.mask = 128'h5577ffffffffffff0000500011111111;

	lut_sub lut_1494 ({sk[456], d, n_n1165, n_n841, n_n1166, x268x, x282x}, x5952x);
	defparam lut_1494.LUT_SIZE = 7;
	defparam lut_1494.mask = 128'h5577ffffffffffff0055035700000303;

	lut_sub lut_1497 ({sk[457], k, n_n1161, n_n1165, x83x, n_n1159, n_n1160}, x5953x);
	defparam lut_1497.LUT_SIZE = 7;
	defparam lut_1497.mask = 128'h5577ffffffffffff0011001f00110011;

	lut_sub lut_1500 ({sk[458], x5950x, x5951x, x5952x, x5953x}, n_n2060);
	defparam lut_1500.LUT_SIZE = 5;
	defparam lut_1500.mask = 32'h5fff7fff;

	lut_sub lut_1505 ({sk[459], j, k, m, n}, x227x);
	defparam lut_1505.LUT_SIZE = 5;
	defparam lut_1505.mask = 32'h5fff0040;

	lut_sub lut_1507 ({sk[460], h, l, n_n1171, x103x, x144x, x227x}, x5968x);
	defparam lut_1507.LUT_SIZE = 7;
	defparam lut_1507.mask = 128'h5577ffffffffffff0357005503030000;

	lut_sub lut_1510 ({sk[461], b, f, n_n1161, x132x, x227x, x5968x}, x5970x);
	defparam lut_1510.LUT_SIZE = 7;
	defparam lut_1510.mask = 128'h5577ffffffffffff5577557757575555;

	lut_sub lut_1514 ({sk[462], x5989x, x5990x, x5991x, x5992x}, x6001x);
	defparam lut_1514.LUT_SIZE = 5;
	defparam lut_1514.mask = 32'h5fff7fff;

	lut_sub lut_1519 ({sk[463], x499x, x5986x, x5987x, x5988x, x5993x, x5995x}, x6002x);
	defparam lut_1519.LUT_SIZE = 7;
	defparam lut_1519.mask = 128'h5577ffffffffffff7fffffffffffffff;

	lut_sub lut_1526 ({sk[464], x6028x, x6029x, x6030x, x6031x}, x6040x);
	defparam lut_1526.LUT_SIZE = 5;
	defparam lut_1526.mask = 32'h5fff7fff;

	lut_sub lut_1531 ({sk[465], x6032x, x6033x, x6034x, x6035x}, x6041x);
	defparam lut_1531.LUT_SIZE = 5;
	defparam lut_1531.mask = 32'h5fff7fff;

	lut_sub lut_1536 ({sk[466], x462x, x464x, x6058x, x6059x}, x6068x);
	defparam lut_1536.LUT_SIZE = 5;
	defparam lut_1536.mask = 32'h5fff7fff;

	lut_sub lut_1541 ({sk[467], x461x, x6057x, x6060x, x6061x, x6062x}, x6069x);
	defparam lut_1541.LUT_SIZE = 6;
	defparam lut_1541.mask = 64'h5f7f5f7f7fffffff;

	lut_sub lut_1547 ({sk[468], c, f, x386x, x146x, n_n1204, x444x}, x6091x);
	defparam lut_1547.LUT_SIZE = 7;
	defparam lut_1547.mask = 128'h5577ffffffffffff5555555555555557;

	lut_sub lut_1550 ({sk[469], d, e, k, n_n1187, x145x, x447x}, x6092x);
	defparam lut_1550.LUT_SIZE = 7;
	defparam lut_1550.mask = 128'h5577ffffffffffff5755555555555555;

	lut_sub lut_1553 ({sk[470], c, f, g, h, x288x, x302x}, x6097x);
	defparam lut_1553.LUT_SIZE = 7;
	defparam lut_1553.mask = 128'h5577ffffffffffff0003000700030005;

	lut_sub lut_1557 ({sk[471], k, n_n1188, x83x, n_n1204, x262x, x158x}, x6098x);
	defparam lut_1557.LUT_SIZE = 7;
	defparam lut_1557.mask = 128'h5577ffffffffffff0000333300053337;

	lut_sub lut_1560 ({sk[472], h, j, x141x, n_n1260, n_n1091, x248x}, x6099x);
	defparam lut_1560.LUT_SIZE = 7;
	defparam lut_1560.mask = 128'h5577ffffffffffff5555000055d500c0;

	lut_sub lut_1563 ({sk[473], x6091x, x6092x, x6097x, x6098x, x6099x}, x6106x);
	defparam lut_1563.LUT_SIZE = 6;
	defparam lut_1563.mask = 64'h5f7f5f7f7fffffff;

	lut_sub lut_1569 ({sk[474], b, g, h, n_n1260, x145x, x288x}, x6130x);
	defparam lut_1569.LUT_SIZE = 7;
	defparam lut_1569.mask = 128'h5577ffffffffffff0303035503030300;

	lut_sub lut_1573 ({sk[475], d, e, x285x, x405x, x145x, x372x}, x6131x);
	defparam lut_1573.LUT_SIZE = 7;
	defparam lut_1573.mask = 128'h5577ffffffffffff0357005500550055;

	lut_sub lut_1576 ({sk[476], x314x, x144x, n_n1260, x145x, x288x, x372x}, x6132x);
	defparam lut_1576.LUT_SIZE = 7;
	defparam lut_1576.mask = 128'h5577ffffffffffff000c000c000c555d;

	lut_sub lut_1579 ({sk[477], l, n_n1177, n_n1116, n_n1118, x37x, x248x}, x6133x);
	defparam lut_1579.LUT_SIZE = 7;
	defparam lut_1579.mask = 128'h5577ffffffffffff5111511151115000;

	lut_sub lut_1583 ({sk[478], x6130x, x6131x, x6132x, x6133x}, x6139x);
	defparam lut_1583.LUT_SIZE = 5;
	defparam lut_1583.mask = 32'h5fff7fff;

	lut_sub lut_1588 ({sk[479], l, m, n}, n_n1219);
	defparam lut_1588.LUT_SIZE = 4;
	defparam lut_1588.mask = 16'h3f20;

	lut_sub lut_1590 ({sk[480], e, f, h}, n_n1160);
	defparam lut_1590.LUT_SIZE = 4;
	defparam lut_1590.mask = 16'h3f20;

	lut_sub lut_1592 ({sk[481], h, i, k, l, m, n}, x422x);
	defparam lut_1592.LUT_SIZE = 7;
	defparam lut_1592.mask = 128'h5577ffffffffffff0000800000000000;

	lut_sub lut_1594 ({sk[482], i, m, n, n_n1089, n_n1160, x422x}, x6149x);
	defparam lut_1594.LUT_SIZE = 7;
	defparam lut_1594.mask = 128'h5577ffffffffffff7f77555555555555;

	lut_sub lut_1599 ({sk[483], h, i, k, l, n_n1187, n_n1039}, x7474x);
	defparam lut_1599.LUT_SIZE = 7;
	defparam lut_1599.mask = 128'h5577ffffffffffffffffceeeffffeeee;

	lut_sub lut_1605 ({sk[484], h, k, l, m, n, n_n977}, x7497x);
	defparam lut_1605.LUT_SIZE = 7;
	defparam lut_1605.mask = 128'h5577ffffffffffffdfffffffffffffff;

	lut_sub lut_1621 ({sk[485], c, g, x226x, x7474x, x7497x}, x6150x);
	defparam lut_1621.LUT_SIZE = 6;
	defparam lut_1621.mask = 64'h5f7f5f7feeeeefee;

	lut_sub lut_1625 ({sk[486], c, e, f, l, n_n1165, x352x}, x6162x);
	defparam lut_1625.LUT_SIZE = 7;
	defparam lut_1625.mask = 128'h5577ffffffffffff5555555575555555;

	lut_sub lut_1628 ({sk[487], x57x, n_n1072, x68x, x204x, x286x}, x6163x);
	defparam lut_1628.LUT_SIZE = 6;
	defparam lut_1628.mask = 64'h5f7f5f7f000c555d;

	lut_sub lut_1631 ({sk[488], g, l, n_n1177, n_n1080, x103x, x356x}, x6166x);
	defparam lut_1631.LUT_SIZE = 7;
	defparam lut_1631.mask = 128'h5577ffffffffffff55775555555f555f;

	lut_sub lut_1635 ({sk[489], i, x114x, x131x, n_n1190, x404x, x6161x}, x6167x);
	defparam lut_1635.LUT_SIZE = 7;
	defparam lut_1635.mask = 128'h5577ffffffffffff55557777555f777f;

	lut_sub lut_1639 ({sk[490], f, j, n_n973, n_n1072, x161x, x399x}, x6168x);
	defparam lut_1639.LUT_SIZE = 7;
	defparam lut_1639.mask = 128'h5577ffffffffffff0303575703035703;

	lut_sub lut_1643 ({sk[491], k, m, n, n_n1028, n_n1072, x6164x}, x6170x);
	defparam lut_1643.LUT_SIZE = 7;
	defparam lut_1643.mask = 128'h5577ffffffffffff55575555555f5555;

	lut_sub lut_1647 ({sk[492], x6162x, x6163x, x6166x, x6167x, x6168x, x6170x}, n_n2023);
	defparam lut_1647.LUT_SIZE = 7;
	defparam lut_1647.mask = 128'h5577ffffffffffff7fffffffffffffff;

	lut_sub lut_1654 ({sk[493], k, n_n1177, n_n1028, x273x, x6199x, x6205x}, x6209x);
	defparam lut_1654.LUT_SIZE = 7;
	defparam lut_1654.mask = 128'h5577ffffffffffff7777777f777777ff;

	lut_sub lut_1659 ({sk[494], x335x, x6196x, x6203x, x6207x}, x6210x);
	defparam lut_1659.LUT_SIZE = 5;
	defparam lut_1659.mask = 32'h5fff7fff;

	lut_sub lut_1664 ({sk[495], x6244x, x6245x, x6246x, x6247x}, x6255x);
	defparam lut_1664.LUT_SIZE = 5;
	defparam lut_1664.mask = 32'h5fff7fff;

	lut_sub lut_1669 ({sk[496], n_n1072, x405x, x307x, x6243x, x6248x, x6249x}, x6256x);
	defparam lut_1669.LUT_SIZE = 7;
	defparam lut_1669.mask = 128'h5577ffffffffffff7fff7fff7fffffff;

	lut_sub lut_1675 ({sk[497], x6275x, x6276x, x6277x, x6278x, x6279x, x6280x}, x6285x);
	defparam lut_1675.LUT_SIZE = 7;
	defparam lut_1675.mask = 128'h5577ffffffffffff7fffffffffffffff;

	lut_sub lut_1682 ({sk[498], i, m, n}, x127x);
	defparam lut_1682.LUT_SIZE = 4;
	defparam lut_1682.mask = 16'h3f80;

	lut_sub lut_1684 ({sk[499], b, m, n}, x263x);
	defparam lut_1684.LUT_SIZE = 4;
	defparam lut_1684.mask = 16'h3f40;

	lut_sub lut_1686 ({sk[500], c, e, f}, n_n1167);
	defparam lut_1686.LUT_SIZE = 4;
	defparam lut_1686.mask = 16'h3f20;

	lut_sub lut_1688 ({sk[501], c, e, f}, x268x);
	defparam lut_1688.LUT_SIZE = 4;
	defparam lut_1688.mask = 16'h3f28;

	lut_sub lut_1691 ({sk[502], i, j, k, m, n}, x312x);
	defparam lut_1691.LUT_SIZE = 6;
	defparam lut_1691.mask = 64'h5f7f5f7f00002000;

	lut_sub lut_1693 ({sk[503], b, m, n}, x404x);
	defparam lut_1693.LUT_SIZE = 4;
	defparam lut_1693.mask = 16'h3f20;

	lut_sub lut_1695 ({sk[504], e, f}, x103x);
	defparam lut_1695.LUT_SIZE = 3;
	defparam lut_1695.mask = 8'h58;

	lut_sub lut_1697 ({sk[505], d, e, f}, n_n1072);
	defparam lut_1697.LUT_SIZE = 4;
	defparam lut_1697.mask = 16'h3f80;

	lut_sub lut_1699 ({sk[506], i, j}, x68x);
	defparam lut_1699.LUT_SIZE = 3;
	defparam lut_1699.mask = 8'h57;

	lut_sub lut_1702 ({sk[507], h, i, j}, x384x);
	defparam lut_1702.LUT_SIZE = 4;
	defparam lut_1702.mask = 16'h3f08;

	lut_sub lut_1704 ({sk[508], j, k, m, n}, x282x);
	defparam lut_1704.LUT_SIZE = 5;
	defparam lut_1704.mask = 32'h5fff0080;

	lut_sub lut_1706 ({sk[509], h, i, j, l}, x373x);
	defparam lut_1706.LUT_SIZE = 5;
	defparam lut_1706.mask = 32'h5fff4000;

	lut_sub lut_1708 ({sk[510], e, g, h}, n_n1196);
	defparam lut_1708.LUT_SIZE = 4;
	defparam lut_1708.mask = 16'h3f10;

	lut_sub lut_1710 ({sk[511], b, c, d, m, n}, x144x);
	defparam lut_1710.LUT_SIZE = 6;
	defparam lut_1710.mask = 64'h5f7f5f7f00000004;

	lut_sub lut_1712 ({sk[512], f, m, n}, x204x);
	defparam lut_1712.LUT_SIZE = 4;
	defparam lut_1712.mask = 16'h3fdf;

	lut_sub lut_1716 ({sk[513], b, j}, x273x);
	defparam lut_1716.LUT_SIZE = 3;
	defparam lut_1716.mask = 8'h57;

	lut_sub lut_1719 ({sk[514], b, e, f}, n_n1121);
	defparam lut_1719.LUT_SIZE = 4;
	defparam lut_1719.mask = 16'h3f20;

	lut_sub lut_1721 ({sk[515], j, k, m, n}, x221x);
	defparam lut_1721.LUT_SIZE = 5;
	defparam lut_1721.mask = 32'h5fff0400;

	lut_sub lut_1723 ({sk[516], h, i, j}, x234x);
	defparam lut_1723.LUT_SIZE = 4;
	defparam lut_1723.mask = 16'h3f7f;

	lut_sub lut_1727 ({sk[517], a, d, e, m, n}, x262x);
	defparam lut_1727.LUT_SIZE = 6;
	defparam lut_1727.mask = 64'h5f7f5f7f00200000;

	lut_sub lut_1729 ({sk[518], h, i, j}, x283x);
	defparam lut_1729.LUT_SIZE = 4;
	defparam lut_1729.mask = 16'h3f40;

	lut_sub lut_1731 ({sk[519], i, k, m, n}, x285x);
	defparam lut_1731.LUT_SIZE = 5;
	defparam lut_1731.mask = 32'h5fff4000;

	lut_sub lut_1733 ({sk[520], h, i, m, n}, x286x);
	defparam lut_1733.LUT_SIZE = 5;
	defparam lut_1733.mask = 32'h5fff4000;

	lut_sub lut_1735 ({sk[521], b, e, f, m, n}, x289x);
	defparam lut_1735.LUT_SIZE = 6;
	defparam lut_1735.mask = 64'h5f7f5f7f00400000;

	lut_sub lut_1737 ({sk[522], k, l, m, n}, x301x);
	defparam lut_1737.LUT_SIZE = 5;
	defparam lut_1737.mask = 32'h5fff4000;

	lut_sub lut_1739 ({sk[523], g, j, k, m, n}, x405x);
	defparam lut_1739.LUT_SIZE = 6;
	defparam lut_1739.mask = 64'h5f7f5f7f22020000;

	lut_sub lut_1742 ({sk[524], j, n_n1161, n_n886, x263x, x286x, x289x}, x5989x);
	defparam lut_1742.LUT_SIZE = 7;
	defparam lut_1742.mask = 128'h5577ffffffffffff0000030300550357;

	lut_sub lut_1745 ({sk[525], f, i, k, m, n, x262x}, x5990x);
	defparam lut_1745.LUT_SIZE = 7;
	defparam lut_1745.mask = 128'h5577ffffffffffff0400000004040004;

	lut_sub lut_1748 ({sk[526], b, x54x, x204x, n_n1121, n_n975, x234x}, x5991x);
	defparam lut_1748.LUT_SIZE = 7;
	defparam lut_1748.mask = 128'h5577ffffffffffff0300abaa03000300;

	lut_sub lut_1751 ({sk[527], b, f, h, x70x, x285x, x289x}, x5992x);
	defparam lut_1751.LUT_SIZE = 7;
	defparam lut_1751.mask = 128'h5577ffffffffffff11111f1111111111;

	lut_sub lut_1754 ({sk[528], h, i, j, n, n_n1227, x289x}, x499x);
	defparam lut_1754.LUT_SIZE = 7;
	defparam lut_1754.mask = 128'h5577ffffffffffff5400545400000000;

	lut_sub lut_1759 ({sk[529], j, m, n, x22x, n_n1171, x37x}, x5986x);
	defparam lut_1759.LUT_SIZE = 7;
	defparam lut_1759.mask = 128'h5577ffffffffffff002200000a2a0a0a;

	lut_sub lut_1762 ({sk[530], x58x, x146x, n_n1036, x263x, n_n1196, x234x}, x5987x);
	defparam lut_1762.LUT_SIZE = 7;
	defparam lut_1762.mask = 128'h5577ffffffffffff000000c0aaaaaaea;

	lut_sub lut_1765 ({sk[531], h, x196x, x54x, n_n1203, x301x, x5976x}, x5988x);
	defparam lut_1765.LUT_SIZE = 7;
	defparam lut_1765.mask = 128'h5577ffffffffffff0050337300500050;

	lut_sub lut_1768 ({sk[532], f, h, i, x221x, x262x, x289x}, x5993x);
	defparam lut_1768.LUT_SIZE = 7;
	defparam lut_1768.mask = 128'h5577ffffffffffff0505050505370505;

	lut_sub lut_1771 ({sk[533], a, e, f, g, x262x, x405x}, x5995x);
	defparam lut_1771.LUT_SIZE = 7;
	defparam lut_1771.mask = 128'h5577ffffffffffff5111111111111111;

	lut_sub lut_1774 ({sk[534], i, j, k}, n_n1133);
	defparam lut_1774.LUT_SIZE = 4;
	defparam lut_1774.mask = 16'h3f04;

	lut_sub lut_1776 ({sk[535], g, h, j}, n_n819);
	defparam lut_1776.LUT_SIZE = 4;
	defparam lut_1776.mask = 16'h3f20;

	lut_sub lut_1778 ({sk[536], g, i, k}, n_n1131);
	defparam lut_1778.LUT_SIZE = 4;
	defparam lut_1778.mask = 16'h3f01;

	lut_sub lut_1780 ({sk[537], c, d, e, f}, x79x);
	defparam lut_1780.LUT_SIZE = 5;
	defparam lut_1780.mask = 32'h5fff0c22;

	lut_sub lut_1783 ({sk[538], c, f, g, h}, x158x);
	defparam lut_1783.LUT_SIZE = 5;
	defparam lut_1783.mask = 32'h5fff1110;

	lut_sub lut_1786 ({sk[539], j, m, n}, x170x);
	defparam lut_1786.LUT_SIZE = 4;
	defparam lut_1786.mask = 16'h3f80;

	lut_sub lut_1788 ({sk[540], c, j, k, n_n1165, n_n1082, x488x}, x6028x);
	defparam lut_1788.LUT_SIZE = 7;
	defparam lut_1788.mask = 128'h5577ffffffffffff5555555557555555;

	lut_sub lut_1791 ({sk[541], h, x171x, n_n1202, n_n1222, x262x, n_n819}, x6029x);
	defparam lut_1791.LUT_SIZE = 7;
	defparam lut_1791.mask = 128'h5577ffffffffffff0303035700000055;

	lut_sub lut_1794 ({sk[542], x133x, n_n1159, x122x, n_n1260, x158x, x170x}, x6030x);
	defparam lut_1794.LUT_SIZE = 7;
	defparam lut_1794.mask = 128'h5577ffffffffffff00001111f000f111;

	lut_sub lut_1797 ({sk[543], h, i, x133x, n_n1195, x312x, n_n975}, x6031x);
	defparam lut_1797.LUT_SIZE = 7;
	defparam lut_1797.mask = 128'h5577ffffffffffff0303030303030357;

	lut_sub lut_1800 ({sk[544], e, g, h, i, x133x, x312x}, x6032x);
	defparam lut_1800.LUT_SIZE = 7;
	defparam lut_1800.mask = 128'h5577ffffffffffff0003000000030055;

	lut_sub lut_1803 ({sk[545], f, n_n861, n_n1080, n_n1133, x79x, x170x}, x6033x);
	defparam lut_1803.LUT_SIZE = 7;
	defparam lut_1803.mask = 128'h5577ffffffffffff0400440000004400;

	lut_sub lut_1806 ({sk[546], f, k, n_n1165, n_n1131, x79x, x486x}, x6034x);
	defparam lut_1806.LUT_SIZE = 7;
	defparam lut_1806.mask = 128'h5577ffffffffffff5555555d55555555;

	lut_sub lut_1809 ({sk[547], i, n_n1080, n_n1072, x170x, x7477x, x7478x}, x6035x);
	defparam lut_1809.LUT_SIZE = 7;
	defparam lut_1809.mask = 128'h5577ffffffffffffeeeeeeeeeeefeeee;

	lut_sub lut_1813 ({sk[548], f, g}, x287x);
	defparam lut_1813.LUT_SIZE = 3;
	defparam lut_1813.mask = 8'h58;

	lut_sub lut_1815 ({sk[549], c, f, g}, n_n1091);
	defparam lut_1815.LUT_SIZE = 4;
	defparam lut_1815.mask = 16'h3f80;

	lut_sub lut_1817 ({sk[550], k, m}, x303x);
	defparam lut_1817.LUT_SIZE = 3;
	defparam lut_1817.mask = 8'h52;

	lut_sub lut_1819 ({sk[551], c, f, g}, x95x);
	defparam lut_1819.LUT_SIZE = 4;
	defparam lut_1819.mask = 16'h3f5c;

	lut_sub lut_1822 ({sk[552], c, d, f}, x395x);
	defparam lut_1822.LUT_SIZE = 4;
	defparam lut_1822.mask = 16'h3fe0;

	lut_sub lut_1825 ({sk[553], g, i, j}, n_n529);
	defparam lut_1825.LUT_SIZE = 4;
	defparam lut_1825.mask = 16'h3f04;

	lut_sub lut_1827 ({sk[554], h, i, j}, n_n670);
	defparam lut_1827.LUT_SIZE = 4;
	defparam lut_1827.mask = 16'h3f04;

	lut_sub lut_1829 ({sk[555], l, m, n}, n_n1215);
	defparam lut_1829.LUT_SIZE = 4;
	defparam lut_1829.mask = 16'h3f02;

	lut_sub lut_1831 ({sk[556], k, l, m, n}, x96x);
	defparam lut_1831.LUT_SIZE = 5;
	defparam lut_1831.mask = 32'h5fff2202;

	lut_sub lut_1834 ({sk[557], g, h, i}, x134x);
	defparam lut_1834.LUT_SIZE = 4;
	defparam lut_1834.mask = 16'h3f60;

	lut_sub lut_1837 ({sk[558], b, d, e, f, h, j}, x176x);
	defparam lut_1837.LUT_SIZE = 7;
	defparam lut_1837.mask = 128'h5577ffffffffffff0000000000100100;

	lut_sub lut_1840 ({sk[559], b, c, d, e}, x47x);
	defparam lut_1840.LUT_SIZE = 5;
	defparam lut_1840.mask = 32'h5fff007c;

	lut_sub lut_1844 ({sk[560], b, c, d, e, f}, x213x);
	defparam lut_1844.LUT_SIZE = 6;
	defparam lut_1844.mask = 64'h5f7f5f7f00cc3ff2;

	lut_sub lut_1850 ({sk[561], g, i, j, k, m, n}, x1202x);
	defparam lut_1850.LUT_SIZE = 7;
	defparam lut_1850.mask = 128'h5577ffffffffffff0000000000000200;

	lut_sub lut_1852 ({sk[562], g, j, k, l, m, n}, x1203x);
	defparam lut_1852.LUT_SIZE = 7;
	defparam lut_1852.mask = 128'h5577ffffffffffff0000000000200000;

	lut_sub lut_1854 ({sk[563], b, g, h, j, x256x, x47x}, x211x);
	defparam lut_1854.LUT_SIZE = 7;
	defparam lut_1854.mask = 128'h5577ffffffffffff0000005000300050;

	lut_sub lut_1857 ({sk[564], f, h, j}, n_n1084);
	defparam lut_1857.LUT_SIZE = 4;
	defparam lut_1857.mask = 16'h3f20;

	lut_sub lut_1859 ({sk[565], f, h, i, j}, x231x);
	defparam lut_1859.LUT_SIZE = 5;
	defparam lut_1859.mask = 32'h5fff0e00;

	lut_sub lut_1862 ({sk[566], b, e, f, l, m, n}, x410x);
	defparam lut_1862.LUT_SIZE = 7;
	defparam lut_1862.mask = 128'h5577ffffffffffff0000000000002000;

	lut_sub lut_1864 ({sk[567], h, j, l}, n_n942);
	defparam lut_1864.LUT_SIZE = 4;
	defparam lut_1864.mask = 16'h3f04;

	lut_sub lut_1866 ({sk[568], e, f, g, m, n, n_n1253}, x248x);
	defparam lut_1866.LUT_SIZE = 7;
	defparam lut_1866.mask = 128'h5577ffffffffffff0000000000000010;

	lut_sub lut_1868 ({sk[569], i, j, k, l, m, n}, x288x);
	defparam lut_1868.LUT_SIZE = 7;
	defparam lut_1868.mask = 128'h5577ffffffffffff0000000000000002;

	lut_sub lut_1870 ({sk[570], c, d, e, l, m, n}, x302x);
	defparam lut_1870.LUT_SIZE = 7;
	defparam lut_1870.mask = 128'h5577ffffffffffff0000000000000080;

	lut_sub lut_1872 ({sk[571], j, k, l}, n_n605);
	defparam lut_1872.LUT_SIZE = 4;
	defparam lut_1872.mask = 16'h3f08;

	lut_sub lut_1874 ({sk[572], k, l, m, n, n_n698, n_n1137}, n_n2953);
	defparam lut_1874.LUT_SIZE = 7;
	defparam lut_1874.mask = 128'h5577ffffffffffff0010000000000000;

	lut_sub lut_1876 ({sk[573], g, h, i, j, x58x, x265x}, x81x);
	defparam lut_1876.LUT_SIZE = 7;
	defparam lut_1876.mask = 128'h5577ffffffffffff0000000000005703;

	lut_sub lut_1879 ({sk[574], g, h, i, j, x54x, x142x}, x5831x);
	defparam lut_1879.LUT_SIZE = 7;
	defparam lut_1879.mask = 128'h5577ffffffffffff0000000005003700;

	lut_sub lut_1882 ({sk[575], g, h, k}, n_n817);
	defparam lut_1882.LUT_SIZE = 4;
	defparam lut_1882.mask = 16'h3f01;

	lut_sub lut_1884 ({sk[576], k, l, m, n}, x161x);
	defparam lut_1884.LUT_SIZE = 5;
	defparam lut_1884.mask = 32'h5fff2220;

	lut_sub lut_1887 ({sk[577], g, k, m, n}, x399x);
	defparam lut_1887.LUT_SIZE = 5;
	defparam lut_1887.mask = 32'h5fff2000;

	lut_sub lut_1889 ({sk[578], e, f, g, m, n}, x416x);
	defparam lut_1889.LUT_SIZE = 6;
	defparam lut_1889.mask = 64'h5f7f5f7f40000000;

	lut_sub lut_1891 ({sk[579], a, c, d, e}, x369x);
	defparam lut_1891.LUT_SIZE = 5;
	defparam lut_1891.mask = 32'h5fff0004;

	lut_sub lut_1893 ({sk[580], g, h, i, n_n711, n_n1053, n_n978}, x5354x);
	defparam lut_1893.LUT_SIZE = 7;
	defparam lut_1893.mask = 128'h5577ffffffffffff0005000000110000;

	lut_sub lut_1896 ({sk[581], i, x114x, x195x, n_n730, n_n838, n_n978}, x5355x);
	defparam lut_1896.LUT_SIZE = 7;
	defparam lut_1896.mask = 128'h5577ffffffffffff000f000f000f111f;

	lut_sub lut_1899 ({sk[582], g, h, i, l, n_n1210, x47x}, x968x);
	defparam lut_1899.LUT_SIZE = 7;
	defparam lut_1899.mask = 128'h5577ffffffffffff0000000000010000;

	lut_sub lut_1901 ({sk[583], g, h, x228x, n_n1171, x247x, x369x}, x5349x);
	defparam lut_1901.LUT_SIZE = 7;
	defparam lut_1901.mask = 128'h5577ffffffffffff11111111111f1111;

	lut_sub lut_1904 ({sk[584], f, x76x, n_n841, x14x, x47x, x247x}, x5356x);
	defparam lut_1904.LUT_SIZE = 7;
	defparam lut_1904.mask = 128'h5577ffffffffffff0505053700000033;

	lut_sub lut_1907 ({sk[585], f, n_n840, n_n709, x76x, x132x, x5351x}, x5358x);
	defparam lut_1907.LUT_SIZE = 7;
	defparam lut_1907.mask = 128'h5577ffffffffffff5557555755555757;

	lut_sub lut_1911 ({sk[586], n_n1137, n_n1053, n_n978, n_n820, n_n982, x5353x}, x5359x);
	defparam lut_1911.LUT_SIZE = 7;
	defparam lut_1911.mask = 128'h5577ffffffffffff5555555f5555777f;

	lut_sub lut_1915 ({sk[587], d, e, g}, n_n919);
	defparam lut_1915.LUT_SIZE = 4;
	defparam lut_1915.mask = 16'h3f04;

	lut_sub lut_1917 ({sk[588], g, i, j}, n_n694);
	defparam lut_1917.LUT_SIZE = 4;
	defparam lut_1917.mask = 16'h3f02;

	lut_sub lut_1919 ({sk[589], e, l, m, n, n_n1171, x37x}, x6199x);
	defparam lut_1919.LUT_SIZE = 7;
	defparam lut_1919.mask = 128'h5577ffffffffffff0a00000002000000;

	lut_sub lut_1922 ({sk[590], x249x, x120x, x103x, x204x, x338x, x6198x}, x6205x);
	defparam lut_1922.LUT_SIZE = 7;
	defparam lut_1922.mask = 128'h5577ffffffffffff77f7777777777777;

	lut_sub lut_1926 ({sk[591], b, e, f, g, n_n1177, x37x}, x335x);
	defparam lut_1926.LUT_SIZE = 7;
	defparam lut_1926.mask = 128'h5577ffffffffffff2022002200000000;

	lut_sub lut_1929 ({sk[592], n_n1177, n_n973, n_n1171, n_n700, x287x, x336x}, x6196x);
	defparam lut_1929.LUT_SIZE = 7;
	defparam lut_1929.mask = 128'h5577ffffffffffff5555555575555555;

	lut_sub lut_1932 ({sk[593], n_n671, n_n700, x404x, n_n1121, n_n1260, x334x}, x6203x);
	defparam lut_1932.LUT_SIZE = 7;
	defparam lut_1932.mask = 128'h5577ffffffffffff55d5555555555555;

	lut_sub lut_1935 ({sk[594], d, i, n_n1177, n_n1028, n_n1121, x6202x}, x6207x);
	defparam lut_1935.LUT_SIZE = 7;
	defparam lut_1935.mask = 128'h5577ffffffffffff5577557f5555555f;

	lut_sub lut_1939 ({sk[595], c, e, f, g}, x35x);
	defparam lut_1939.LUT_SIZE = 5;
	defparam lut_1939.mask = 32'h5fff002e;

	lut_sub lut_1942 ({sk[596], c, e, f, m, n}, x418x);
	defparam lut_1942.LUT_SIZE = 6;
	defparam lut_1942.mask = 64'h5f7f5f7f00008000;

	lut_sub lut_1944 ({sk[597], i, j, n_n1165, n_n1072, n_n919, x418x}, x6244x);
	defparam lut_1944.LUT_SIZE = 7;
	defparam lut_1944.mask = 128'h5577ffffffffffff0005444500004444;

	lut_sub lut_1947 ({sk[598], e, f, g, i, x131x, x170x}, x6245x);
	defparam lut_1947.LUT_SIZE = 7;
	defparam lut_1947.mask = 128'h5577ffffffffffff0001111100010000;

	lut_sub lut_1950 ({sk[599], g, n_n1190, n_n1202, x127x, n_n1167, n_n1091}, x6246x);
	defparam lut_1950.LUT_SIZE = 7;
	defparam lut_1950.mask = 128'h5577ffffffffffff0050005000503373;

	lut_sub lut_1953 ({sk[600], c, d, e, n_n1177, x262x, x310x}, x6247x);
	defparam lut_1953.LUT_SIZE = 7;
	defparam lut_1953.mask = 128'h5577ffffffffffff0005330000000000;

	lut_sub lut_1956 ({sk[601], f, n_n857, x90x, x35x, x6217x, x6215x}, x307x);
	defparam lut_1956.LUT_SIZE = 7;
	defparam lut_1956.mask = 128'h5577ffffffffffff1010000010000000;

	lut_sub lut_1959 ({sk[602], a, n_n1187, x127x, n_n919, x6231x, x6234x}, x6243x);
	defparam lut_1959.LUT_SIZE = 7;
	defparam lut_1959.mask = 128'h5577ffffffffffff3000755530003000;

	lut_sub lut_1962 ({sk[603], j, n_n1165, n_n1219, x262x, x303x, x7476x}, x6248x);
	defparam lut_1962.LUT_SIZE = 7;
	defparam lut_1962.mask = 128'h5577ffffffffffff000f222f000f000f;

	lut_sub lut_1965 ({sk[604], m, n, x83x, x35x, x6229x, x325x}, x6249x);
	defparam lut_1965.LUT_SIZE = 7;
	defparam lut_1965.mask = 128'h5577ffffffffffff5575555555555555;

	lut_sub lut_1968 ({sk[605], g, h, j, k}, x216x);
	defparam lut_1968.LUT_SIZE = 5;
	defparam lut_1968.mask = 32'h5fff0d22;

	lut_sub lut_1972 ({sk[606], j, l, m, n}, x260x);
	defparam lut_1972.LUT_SIZE = 5;
	defparam lut_1972.mask = 32'h5fff0800;

	lut_sub lut_1974 ({sk[607], b, c, f, l, m, n}, x295x);
	defparam lut_1974.LUT_SIZE = 7;
	defparam lut_1974.mask = 128'h5577ffffffffffff0000000400000000;

	lut_sub lut_1976 ({sk[608], a, b, e, l, m, n}, x383x);
	defparam lut_1976.LUT_SIZE = 7;
	defparam lut_1976.mask = 128'h5577ffffffffffff0000000200000000;

	lut_sub lut_1978 ({sk[609], j, k, m, n}, x293x);
	defparam lut_1978.LUT_SIZE = 5;
	defparam lut_1978.mask = 32'h5fff0440;

	lut_sub lut_1981 ({sk[610], f, h, k}, n_n825);
	defparam lut_1981.LUT_SIZE = 4;
	defparam lut_1981.mask = 16'h3f10;

	lut_sub lut_1983 ({sk[611], h, i, j, l, m, n}, x296x);
	defparam lut_1983.LUT_SIZE = 7;
	defparam lut_1983.mask = 128'h5577ffffffffffff0000080000000000;

	lut_sub lut_1985 ({sk[612], c, d, e, f}, x109x);
	defparam lut_1985.LUT_SIZE = 5;
	defparam lut_1985.mask = 32'h5fff0d66;

	lut_sub lut_1990 ({sk[613], g, h, i, l, m, n}, x1114x);
	defparam lut_1990.LUT_SIZE = 7;
	defparam lut_1990.mask = 128'h5577ffffffffffff0000000000020200;

	lut_sub lut_1993 ({sk[614], g, h, j, l, m, n}, x1115x);
	defparam lut_1993.LUT_SIZE = 7;
	defparam lut_1993.mask = 128'h5577ffffffffffff0000000000000020;

	lut_sub lut_1995 ({sk[615], h, k, l, m, n}, x292x);
	defparam lut_1995.LUT_SIZE = 6;
	defparam lut_1995.mask = 64'h5f7f5f7f00000020;

	lut_sub lut_1997 ({sk[616], c, d, e, f, h, i}, x406x);
	defparam lut_1997.LUT_SIZE = 7;
	defparam lut_1997.mask = 128'h5577ffffffffffff0000000000000040;

	lut_sub lut_1999 ({sk[617], n_n703, x89x, x192x, n_n1219, x5079x, x5080x}, x5093x);
	defparam lut_1999.LUT_SIZE = 7;
	defparam lut_1999.mask = 128'h5577ffffffffffff030303ff575757ff;

	lut_sub lut_2003 ({sk[618], f, g, i, n_n709, x45x, x33x}, x1196x);
	defparam lut_2003.LUT_SIZE = 7;
	defparam lut_2003.mask = 128'h5577ffffffffffff0000030700000000;

	lut_sub lut_2006 ({sk[619], b, x259x, n_n1036, n_n823, x260x, x406x}, x5090x);
	defparam lut_2006.LUT_SIZE = 7;
	defparam lut_2006.mask = 128'h5577ffffffffffff111111111111111f;

	lut_sub lut_2009 ({sk[620], g, h, i, j, k, x383x}, x5091x);
	defparam lut_2009.LUT_SIZE = 7;
	defparam lut_2009.mask = 128'h5577ffffffffffff0000505004555504;

	lut_sub lut_2014 ({sk[621], k, n_n1177, x374x, n_n698, n_n1137, n_n1219}, x5092x);
	defparam lut_2014.LUT_SIZE = 7;
	defparam lut_2014.mask = 128'h5577ffffffffffff01010101010101ff;

	lut_sub lut_2017 ({sk[622], h, i, j, k, m, n}, x162x);
	defparam lut_2017.LUT_SIZE = 7;
	defparam lut_2017.mask = 128'h5577ffffffffffff0888088808880880;

	lut_sub lut_2022 ({sk[623], b, c, d, e, f, h}, x300x);
	defparam lut_2022.LUT_SIZE = 7;
	defparam lut_2022.mask = 128'h5577ffffffffffff0000000000000400;

	lut_sub lut_2024 ({sk[624], g, h, i, n_n996, n_n1072, x193x}, x26x);
	defparam lut_2024.LUT_SIZE = 7;
	defparam lut_2024.mask = 128'h5577ffffffffffff0000000001000000;

	lut_sub lut_2026 ({sk[625], i, j, k, n_n973, n_n971, n_n1204}, x42x);
	defparam lut_2026.LUT_SIZE = 7;
	defparam lut_2026.mask = 128'h5577ffffffffffff0100000000000000;

	lut_sub lut_2028 ({sk[626], g, h, i, j, k, m}, x253x);
	defparam lut_2028.LUT_SIZE = 7;
	defparam lut_2028.mask = 128'h5577ffffffffffff0000008000008000;

	lut_sub lut_2031 ({sk[627], c, d, e, f, g, j}, x6217x);
	defparam lut_2031.LUT_SIZE = 7;
	defparam lut_2031.mask = 128'h5577ffffffffffff3d3d0c3df0f0ccfd;

	lut_sub lut_2047 ({sk[628], e, f, g, i, m, n}, x6215x);
	defparam lut_2047.LUT_SIZE = 7;
	defparam lut_2047.mask = 128'h5577ffffffffffff0808000808080808;

	lut_sub lut_2051 ({sk[629], c, d, f, g, j}, x6229x);
	defparam lut_2051.LUT_SIZE = 6;
	defparam lut_2051.mask = 64'h5f7f5f7f3e00fefe;

	lut_sub lut_2059 ({sk[630], c, f, l, m, n}, x6231x);
	defparam lut_2059.LUT_SIZE = 6;
	defparam lut_2059.mask = 64'h5f7f5f7f80000000;

	lut_sub lut_2061 ({sk[631], e, f, h, i, j}, x6234x);
	defparam lut_2061.LUT_SIZE = 6;
	defparam lut_2061.mask = 64'h5f7f5f7f7f000000;

	lut_sub lut_2065 ({sk[632], a, e, f, k, l, n_n1187}, x325x);
	defparam lut_2065.LUT_SIZE = 7;
	defparam lut_2065.mask = 128'h5577ffffffffffff5400000000000000;

	lut_sub lut_2068 ({sk[633], b, f, l, n_n1177, x37x}, x334x);
	defparam lut_2068.LUT_SIZE = 6;
	defparam lut_2068.mask = 64'h5f7f5f7f00000002;

	lut_sub lut_2070 ({sk[634], b, e, f, g, l, n_n1177}, x336x);
	defparam lut_2070.LUT_SIZE = 7;
	defparam lut_2070.mask = 128'h5577ffffffffffff4000440000000000;

	lut_sub lut_2073 ({sk[635], g, h, i, j, m, n}, x338x);
	defparam lut_2073.LUT_SIZE = 7;
	defparam lut_2073.mask = 128'h5577ffffffffffff0000000080000000;

	lut_sub lut_2075 ({sk[636], h, i, k, l, m, n}, x340x);
	defparam lut_2075.LUT_SIZE = 7;
	defparam lut_2075.mask = 128'h5577ffffffffffff0040000000000000;

	lut_sub lut_2077 ({sk[637], c, d, h, i, m, n}, x348x);
	defparam lut_2077.LUT_SIZE = 7;
	defparam lut_2077.mask = 128'h5577ffffffffffff0000000080000000;

	lut_sub lut_2079 ({sk[638], c, d, f, g, m, n}, x352x);
	defparam lut_2079.LUT_SIZE = 7;
	defparam lut_2079.mask = 128'h5577ffffffffffff0080800000000000;

	lut_sub lut_2082 ({sk[639], c, d, f, g, m, n}, x356x);
	defparam lut_2082.LUT_SIZE = 7;
	defparam lut_2082.mask = 128'h5577ffffffffffff0000400000000000;

	lut_sub lut_2084 ({sk[640], e, f, h, i, j, x144x}, x432x);
	defparam lut_2084.LUT_SIZE = 7;
	defparam lut_2084.mask = 128'h5577ffffffffffff0111000000000000;

	lut_sub lut_2087 ({sk[641], c, d, e, n, n_n1228, n_n1227}, x434x);
	defparam lut_2087.LUT_SIZE = 7;
	defparam lut_2087.mask = 128'h5577ffffffffffff0000000000000010;

	lut_sub lut_2089 ({sk[642], b, c, d, e, l, x145x}, x444x);
	defparam lut_2089.LUT_SIZE = 7;
	defparam lut_2089.mask = 128'h5577ffffffffffff4040404040404000;

	lut_sub lut_2093 ({sk[643], h, i, m, n, x112x, n_n1229}, x447x);
	defparam lut_2093.LUT_SIZE = 7;
	defparam lut_2093.mask = 128'h5577ffffffffffff0000100000000000;

	lut_sub lut_2095 ({sk[644], h, k, m, n, n_n1203, x68x}, x449x);
	defparam lut_2095.LUT_SIZE = 7;
	defparam lut_2095.mask = 128'h5577ffffffffffff0000000020000000;

	lut_sub lut_2097 ({sk[645], d, f, x255x, n_n1203, n_n1227, n_n1204}, x461x);
	defparam lut_2097.LUT_SIZE = 7;
	defparam lut_2097.mask = 128'h5577ffffffffffff0040000000000000;

	lut_sub lut_2099 ({sk[646], c, d, f, i, x226x, x303x}, x462x);
	defparam lut_2099.LUT_SIZE = 7;
	defparam lut_2099.mask = 128'h5577ffffffffffff0000001000100010;

	lut_sub lut_2102 ({sk[647], c, f, g, h, n, n_n1227}, x464x);
	defparam lut_2102.LUT_SIZE = 7;
	defparam lut_2102.mask = 128'h5577ffffffffffff0000400040004000;

	lut_sub lut_2105 ({sk[648], c, e, f, n_n861, n_n1202}, x486x);
	defparam lut_2105.LUT_SIZE = 6;
	defparam lut_2105.mask = 64'h5f7f5f7f00111101;

	lut_sub lut_2110 ({sk[649], c, e, f, g, i, n_n1191}, x488x);
	defparam lut_2110.LUT_SIZE = 7;
	defparam lut_2110.mask = 128'h5577ffffffffffff0000000040000000;

	lut_sub lut_2112 ({sk[650], c, e, f, h, i, j}, x5976x);
	defparam lut_2112.LUT_SIZE = 7;
	defparam lut_2112.mask = 128'h5577ffffffffffff8080808000808080;

	lut_sub lut_2116 ({sk[651], e, f, m, n, x373x}, x529x);
	defparam lut_2116.LUT_SIZE = 6;
	defparam lut_2116.mask = 64'h5f7f5f7f00000400;

	lut_sub lut_2118 ({sk[652], g, h, i, k, n_n1177, x36x}, x539x);
	defparam lut_2118.LUT_SIZE = 7;
	defparam lut_2118.mask = 128'h5577ffffffffffff0000000000010000;

	lut_sub lut_2120 ({sk[653], h, i, k, m, n, x52x}, x547x);
	defparam lut_2120.LUT_SIZE = 7;
	defparam lut_2120.mask = 128'h5577ffffffffffff0000004000000000;

	lut_sub lut_2122 ({sk[654], j, k, m, n, x122x, x52x}, x548x);
	defparam lut_2122.LUT_SIZE = 7;
	defparam lut_2122.mask = 128'h5577ffffffffffff0000400000000000;

	lut_sub lut_2124 ({sk[655], c, n_n1203, n_n1202, n_n1264, n_n1036, x310x}, x555x);
	defparam lut_2124.LUT_SIZE = 7;
	defparam lut_2124.mask = 128'h5577ffffffffffff0000000f0105010f;

	lut_sub lut_2128 ({sk[656], f, g, h, n_n1220, n_n918, x29x}, x556x);
	defparam lut_2128.LUT_SIZE = 7;
	defparam lut_2128.mask = 128'h5577ffffffffffff0003000000050000;

	lut_sub lut_2131 ({sk[657], n_n1201, x146x, x48x, n_n1196, n_n1133, x293x}, x564x);
	defparam lut_2131.LUT_SIZE = 7;
	defparam lut_2131.mask = 128'h5577ffffffffffff0000001000000000;

	lut_sub lut_2133 ({sk[658], a, c, d, e, h, j}, x5880x);
	defparam lut_2133.LUT_SIZE = 7;
	defparam lut_2133.mask = 128'h5577ffffffffffff2222222220222020;

	lut_sub lut_2137 ({sk[659], f, g, h, i, n_n1187, n_n918}, x5833x);
	defparam lut_2137.LUT_SIZE = 7;
	defparam lut_2137.mask = 128'h5577ffffffffffff1111111111110100;

	lut_sub lut_2141 ({sk[660], i, k, m, n}, x5839x);
	defparam lut_2141.LUT_SIZE = 5;
	defparam lut_2141.mask = 32'h5fff0002;

	lut_sub lut_2143 ({sk[661], a, b, d, e, g, x190x}, x645x);
	defparam lut_2143.LUT_SIZE = 7;
	defparam lut_2143.mask = 128'h5577ffffffffffff0000000000000040;

	lut_sub lut_2145 ({sk[662], a, c, d, n_n1187, x417x, x182x}, x713x);
	defparam lut_2145.LUT_SIZE = 7;
	defparam lut_2145.mask = 128'h5577ffffffffffff0000000000000001;

	lut_sub lut_2147 ({sk[663], a, c, d, n_n1187, x183x, n_n1231}, x716x);
	defparam lut_2147.LUT_SIZE = 7;
	defparam lut_2147.mask = 128'h5577ffffffffffff0000000000000001;

	lut_sub lut_2149 ({sk[664], a, b, c, d, x44x, x174x}, x717x);
	defparam lut_2149.LUT_SIZE = 7;
	defparam lut_2149.mask = 128'h5577ffffffffffff0000000000000002;

	lut_sub lut_2151 ({sk[665], a, b, c, d, x108x}, x722x);
	defparam lut_2151.LUT_SIZE = 6;
	defparam lut_2151.mask = 64'h5f7f5f7f00040000;

	lut_sub lut_2153 ({sk[666], f, g, i, x45x, x33x, n_n761}, x727x);
	defparam lut_2153.LUT_SIZE = 7;
	defparam lut_2153.mask = 128'h5577ffffffffffff0000051500000000;

	lut_sub lut_2156 ({sk[667], d, f, g, n_n1187, x74x, n_n997}, x750x);
	defparam lut_2156.LUT_SIZE = 7;
	defparam lut_2156.mask = 128'h5577ffffffffffff0000000100000000;

	lut_sub lut_2158 ({sk[668], i, j, k, n_n1187, n_n1201, n_n698}, x785x);
	defparam lut_2158.LUT_SIZE = 7;
	defparam lut_2158.mask = 128'h5577ffffffffffff0000000000000100;

	lut_sub lut_2160 ({sk[669], f, g, h, n_n893, x148x, x29x}, x786x);
	defparam lut_2160.LUT_SIZE = 7;
	defparam lut_2160.mask = 128'h5577ffffffffffff0000000000010000;

	lut_sub lut_2162 ({sk[670], i, k, m, n, x15x, n_n1194}, x788x);
	defparam lut_2162.LUT_SIZE = 7;
	defparam lut_2162.mask = 128'h5577ffffffffffff0000000000000010;

	lut_sub lut_2164 ({sk[671], f, g, h, k, l, m}, x5530x);
	defparam lut_2164.LUT_SIZE = 7;
	defparam lut_2164.mask = 128'h5577ffffffffffff0000000000000008;

	lut_sub lut_2166 ({sk[672], b, c, e, g, h, x172x}, x813x);
	defparam lut_2166.LUT_SIZE = 7;
	defparam lut_2166.mask = 128'h5577ffffffffffff0000000000010000;

	lut_sub lut_2168 ({sk[673], f, l, x171x, n_n1165, n_n626, n_n817}, x829x);
	defparam lut_2168.LUT_SIZE = 7;
	defparam lut_2168.mask = 128'h5577ffffffffffff0101000001050000;

	lut_sub lut_2171 ({sk[674], g, h, i, l, n_n1187, n_n1171}, x837x);
	defparam lut_2171.LUT_SIZE = 7;
	defparam lut_2171.mask = 128'h5577ffffffffffff0000000000010000;

	lut_sub lut_2173 ({sk[675], b, f, x256x, x53x, x229x, x298x}, x842x);
	defparam lut_2173.LUT_SIZE = 7;
	defparam lut_2173.mask = 128'h5577ffffffffffff1100000010001000;

	lut_sub lut_2177 ({sk[676], b, d, f, g, x74x, x120x}, x845x);
	defparam lut_2177.LUT_SIZE = 7;
	defparam lut_2177.mask = 128'h5577ffffffffffff0000000100000000;

	lut_sub lut_2179 ({sk[677], f, g, n_n842, x46x, x75x, n_n1166}, x846x);
	defparam lut_2179.LUT_SIZE = 7;
	defparam lut_2179.mask = 128'h5577ffffffffffff0001000100010000;

	lut_sub lut_2182 ({sk[678], b, m, n, x171x, x229x, x101x}, x847x);
	defparam lut_2182.LUT_SIZE = 7;
	defparam lut_2182.mask = 128'h5577ffffffffffff0000000000010000;

	lut_sub lut_2184 ({sk[679], m, n, n_n996, x29x, x921x, n_n1228}, x905x);
	defparam lut_2184.LUT_SIZE = 7;
	defparam lut_2184.mask = 128'h5577ffffffffffff0000000003070000;

	lut_sub lut_2187 ({sk[680], g, h, i, n_n703, n_n838, x133x}, x906x);
	defparam lut_2187.LUT_SIZE = 7;
	defparam lut_2187.mask = 128'h5577ffffffffffff0000150000000000;

	lut_sub lut_2190 ({sk[681], b, d, e, f, h, j}, x5377x);
	defparam lut_2190.LUT_SIZE = 7;
	defparam lut_2190.mask = 128'h5577ffffffffffff0000000000000200;

	lut_sub lut_2192 ({sk[682], h, i, k, x961x, x52x, n_n1204}, x954x);
	defparam lut_2192.LUT_SIZE = 7;
	defparam lut_2192.mask = 128'h5577ffffffffffff0000001f00000000;

	lut_sub lut_2195 ({sk[683], i, n, x22x, x31x, x54x, x258x}, x1047x);
	defparam lut_2195.LUT_SIZE = 7;
	defparam lut_2195.mask = 128'h5577ffffffffffff0400000000000000;

	lut_sub lut_2197 ({sk[684], n, n_n904, n_n1193, x22x, x31x, x54x}, x1048x);
	defparam lut_2197.LUT_SIZE = 7;
	defparam lut_2197.mask = 128'h5577ffffffffffff0000002000000000;

	lut_sub lut_2199 ({sk[685], i, m, n, x101x, x258x}, x1049x);
	defparam lut_2199.LUT_SIZE = 6;
	defparam lut_2199.mask = 64'h5f7f5f7f00000010;

	lut_sub lut_2201 ({sk[686], c, e, f, x1208x, x5088x}, x1060x);
	defparam lut_2201.LUT_SIZE = 6;
	defparam lut_2201.mask = 64'h5f7f5f7f00000700;

	lut_sub lut_2204 ({sk[687], c, d, e, f, h, i}, x5219x);
	defparam lut_2204.LUT_SIZE = 7;
	defparam lut_2204.mask = 128'h5577ffffffffffff0000000000000400;

	lut_sub lut_2206 ({sk[688], e, f, g, n_n713, x75x, x20x}, x1091x);
	defparam lut_2206.LUT_SIZE = 7;
	defparam lut_2206.mask = 128'h5577ffffffffffff0000000100000000;

	lut_sub lut_2208 ({sk[689], e, f, g, h, k, x27x}, x1096x);
	defparam lut_2208.LUT_SIZE = 7;
	defparam lut_2208.mask = 128'h5577ffffffffffff0100010000000000;

	lut_sub lut_2211 ({sk[690], d, e, f, g, n_n920, x190x}, x1123x);
	defparam lut_2211.LUT_SIZE = 7;
	defparam lut_2211.mask = 128'h5577ffffffffffff0000001000000000;

	lut_sub lut_2213 ({sk[691], b, d, e, f, g, h}, x5104x);
	defparam lut_2213.LUT_SIZE = 7;
	defparam lut_2213.mask = 128'h5577ffffffffffff0000000000010000;

	lut_sub lut_2215 ({sk[692], b, d, e, h, x112x, x172x}, x1158x);
	defparam lut_2215.LUT_SIZE = 7;
	defparam lut_2215.mask = 128'h5577ffffffffffff0000000000010000;

	lut_sub lut_2217 ({sk[693], c, d, e, f, h}, x5107x);
	defparam lut_2217.LUT_SIZE = 6;
	defparam lut_2217.mask = 64'h5f7f5f7f00000004;

	lut_sub lut_2219 ({sk[694], c, d, f, x65x, x162x}, x1161x);
	defparam lut_2219.LUT_SIZE = 6;
	defparam lut_2219.mask = 64'h5f7f5f7f00000100;

	lut_sub lut_2221 ({sk[695], b, d, e, f, h, k}, x5079x);
	defparam lut_2221.LUT_SIZE = 7;
	defparam lut_2221.mask = 128'h5577ffffffffffff0000000000100000;

	lut_sub lut_2223 ({sk[696], g, h, i, k, m, n}, x5080x);
	defparam lut_2223.LUT_SIZE = 7;
	defparam lut_2223.mask = 128'h5577ffffffffffff0000040000000000;

	lut_sub lut_2225 ({sk[697], i, j, l, m, n_n709, x385x}, x5117x);
	defparam lut_2225.LUT_SIZE = 7;
	defparam lut_2225.mask = 128'h5577ffffffffffff0001010100000100;

	lut_sub lut_2228 ({sk[698], m, n, n_n626, n_n235, n_n617, x1158x}, x5118x);
	defparam lut_2228.LUT_SIZE = 7;
	defparam lut_2228.mask = 128'h5577ffffffffffff557f555555555555;

	lut_sub lut_2232 ({sk[699], f, n_n840, n_n709, n_n1201, x121x, x77x}, x5119x);
	defparam lut_2232.LUT_SIZE = 7;
	defparam lut_2232.mask = 128'h5577ffffffffffff0005000500051115;

	lut_sub lut_2235 ({sk[700], b, d, e, x54x, n_n1220, n_n971}, x5120x);
	defparam lut_2235.LUT_SIZE = 7;
	defparam lut_2235.mask = 128'h5577ffffffffffff0000000000150000;

	lut_sub lut_2238 ({sk[701], c, d, f, n_n235, n_n1191, x406x}, x5121x);
	defparam lut_2238.LUT_SIZE = 7;
	defparam lut_2238.mask = 128'h5577ffffffffffff1111111111131111;

	lut_sub lut_2241 ({sk[702], f, x249x, x172x, x377x, n_n1195, x296x}, x5124x);
	defparam lut_2241.LUT_SIZE = 7;
	defparam lut_2241.mask = 128'h5577ffffffffffff0003000300035557;

	lut_sub lut_2244 ({sk[703], x172x, n_n626, x65x, x296x, x162x, x300x}, x5130x);
	defparam lut_2244.LUT_SIZE = 7;
	defparam lut_2244.mask = 128'h5577ffffffffffff00000f3f55555f7f;

	lut_sub lut_2248 ({sk[704], x377x, x77x, x293x, x162x, x5104x, x5107x}, x5133x);
	defparam lut_2248.LUT_SIZE = 7;
	defparam lut_2248.mask = 128'h5577ffffffffffff0537053705ffffff;

	lut_sub lut_2253 ({sk[705], n_n711, n_n709, n_n1188, n_n886, x148x, x172x}, x5157x);
	defparam lut_2253.LUT_SIZE = 7;
	defparam lut_2253.mask = 128'h5577ffffffffffff0000003305050537;

	lut_sub lut_2256 ({sk[706], h, n_n713, x84x, x175x, x229x, x1123x}, x5159x);
	defparam lut_2256.LUT_SIZE = 7;
	defparam lut_2256.mask = 128'h5577ffffffffffff555555d555555555;

	lut_sub lut_2259 ({sk[707], n_n1207, x53x, x84x, x202x, x76x, n_n1095}, x5160x);
	defparam lut_2259.LUT_SIZE = 7;
	defparam lut_2259.mask = 128'h5577ffffffffffff01010000010f000f;

	lut_sub lut_2262 ({sk[708], i, k, m, n, n_n893, x393x}, x5161x);
	defparam lut_2262.LUT_SIZE = 7;
	defparam lut_2262.mask = 128'h5577ffffffffffff0100010001000500;

	lut_sub lut_2265 ({sk[709], x53x, x38x, x46x, x202x, x76x, n_n1095}, x5168x);
	defparam lut_2265.LUT_SIZE = 7;
	defparam lut_2265.mask = 128'h5577ffffffffffff00010001000100ff;

	lut_sub lut_2268 ({sk[710], n_n840, x153x, x187x, x298x, x306x, x374x}, x7496x);
	defparam lut_2268.LUT_SIZE = 7;
	defparam lut_2268.mask = 128'h5577ffffffffffff050537ff0f0f3fff;

	lut_sub lut_2281 ({sk[711], n_n1188, x27x, x90x, n_n819, n_n1215, x1091x}, x5197x);
	defparam lut_2281.LUT_SIZE = 7;
	defparam lut_2281.mask = 128'h5577ffffffffffff5555575555557755;

	lut_sub lut_2285 ({sk[712], d, e, f, g, x121x, n_n942}, x7494x);
	defparam lut_2285.LUT_SIZE = 7;
	defparam lut_2285.mask = 128'h5577ffffffffffffffafffffffafcfcf;

	lut_sub lut_2295 ({sk[713], e, f, g, x27x, x74x, x111x}, x5206x);
	defparam lut_2295.LUT_SIZE = 7;
	defparam lut_2295.mask = 128'h5577ffffffffffff0003001300000000;

	lut_sub lut_2299 ({sk[714], a, b, c, n_n1187, x182x, x90x}, x7493x);
	defparam lut_2299.LUT_SIZE = 7;
	defparam lut_2299.mask = 128'h5577ffffffffffffffffeeeefffeffff;

	lut_sub lut_2308 ({sk[715], n_n1187, n_n949, x108x, x1096x, x5197x, x7493x}, x5209x);
	defparam lut_2308.LUT_SIZE = 7;
	defparam lut_2308.mask = 128'h5577ffffffffffffbfbfbfbfbfbfbfff;

	lut_sub lut_2313 ({sk[716], a, b, x123x, x111x, x90x, x5206x}, x5210x);
	defparam lut_2313.LUT_SIZE = 7;
	defparam lut_2313.mask = 128'h5577ffffffffffff5557557755575557;

	lut_sub lut_2317 ({sk[717], f, h, m, n}, x5246x);
	defparam lut_2317.LUT_SIZE = 5;
	defparam lut_2317.mask = 32'h5fff0800;

	lut_sub lut_2319 ({sk[718], f, h, x31x, x45x, x54x, x258x}, x5256x);
	defparam lut_2319.LUT_SIZE = 7;
	defparam lut_2319.mask = 128'h5577ffffffffffff0505051505050505;

	lut_sub lut_2322 ({sk[719], x84x, x172x, x393x, x377x, x115x, x1110x}, x5260x);
	defparam lut_2322.LUT_SIZE = 7;
	defparam lut_2322.mask = 128'h5577ffffffffffff00003f3f55ff7fff;

	lut_sub lut_2327 ({sk[720], c, d, e, f, m, n}, x7492x);
	defparam lut_2327.LUT_SIZE = 7;
	defparam lut_2327.mask = 128'h5577fffffffffffffffff7f7fffff7ff;

	lut_sub lut_2333 ({sk[721], n_n1177, n_n671, n_n1229, x101x, x5246x, x7492x}, x5264x);
	defparam lut_2333.LUT_SIZE = 7;
	defparam lut_2333.mask = 128'h5577ffffffffffff0a0b0a0b0a0b0f0f;

	lut_sub lut_2337 ({sk[722], a, b, e, f, n_n529, x96x}, x5290x);
	defparam lut_2337.LUT_SIZE = 7;
	defparam lut_2337.mask = 128'h5577ffffffffffff0000001100000010;

	lut_sub lut_2340 ({sk[723], g, h, i, x58x, n_n698, n_n1171}, x5293x);
	defparam lut_2340.LUT_SIZE = 7;
	defparam lut_2340.mask = 128'h5577ffffffffffff0000000000070000;

	lut_sub lut_2343 ({sk[724], n_n1217, n_n1220, x265x, n_n698, n_n841, n_n1137}, x5319x);
	defparam lut_2343.LUT_SIZE = 7;
	defparam lut_2343.mask = 128'h5577ffffffffffff0005000500050307;

	lut_sub lut_2346 ({sk[725], j, n_n1201, n_n1220, x15x, x265x, n_n1194}, x5320x);
	defparam lut_2346.LUT_SIZE = 7;
	defparam lut_2346.mask = 128'h5577ffffffffffff0000030300050307;

	lut_sub lut_2349 ({sk[726], a, b, c, d, x390x, x417x}, x5322x);
	defparam lut_2349.LUT_SIZE = 7;
	defparam lut_2349.mask = 128'h5577ffffffffffff0000303000330505;

	lut_sub lut_2353 ({sk[727], i, x258x, x228x, x265x, x5319x, x5320x}, x5324x);
	defparam lut_2353.LUT_SIZE = 7;
	defparam lut_2353.mask = 128'h5577ffffffffffff77777fff77777777;

	lut_sub lut_2358 ({sk[728], i, j, k, n_n1187, x58x, x98x}, x5325x);
	defparam lut_2358.LUT_SIZE = 7;
	defparam lut_2358.mask = 128'h5577ffffffffffff0000000011111115;

	lut_sub lut_2361 ({sk[729], n_n709, x76x, n_n841, n_n1053, n_n662, n_n978}, x5351x);
	defparam lut_2361.LUT_SIZE = 7;
	defparam lut_2361.mask = 128'h5577ffffffffffff0000000f1111111f;

	lut_sub lut_2364 ({sk[730], b, x259x, n_n1095, n_n671, n_n978, n_n670}, x5353x);
	defparam lut_2364.LUT_SIZE = 7;
	defparam lut_2364.mask = 128'h5577ffffffffffff0101010101010133;

	lut_sub lut_2367 ({sk[731], g, k, n_n700, x132x, x146x, n_n1204}, x5379x);
	defparam lut_2367.LUT_SIZE = 7;
	defparam lut_2367.mask = 128'h5577ffffffffffff0000000000000015;

	lut_sub lut_2370 ({sk[732], n_n709, n_n1171, n_n978, n_n1084, n_n694, x142x}, x5380x);
	defparam lut_2370.LUT_SIZE = 7;
	defparam lut_2370.mask = 128'h5577ffffffffffff00001111000f111f;

	lut_sub lut_2373 ({sk[733], h, i, j, k, x295x}, x5382x);
	defparam lut_2373.LUT_SIZE = 6;
	defparam lut_2373.mask = 64'h5f7f5f7f00510404;

	lut_sub lut_2377 ({sk[734], j, n_n841, n_n1171, x121x, n_n978, x295x}, x5383x);
	defparam lut_2377.LUT_SIZE = 7;
	defparam lut_2377.mask = 128'h5577ffffffffffff0505053700000033;

	lut_sub lut_2380 ({sk[735], h, i, j, k, n_n711, x30x}, x7499x);
	defparam lut_2380.LUT_SIZE = 7;
	defparam lut_2380.mask = 128'h5577fffffffffffffffffdfdffdfffdf;

	lut_sub lut_2406 ({sk[736], l, n_n1187, n_n1171, n_n1036, x216x, x7499x}, x5384x);
	defparam lut_2406.LUT_SIZE = 7;
	defparam lut_2406.mask = 128'h5577ffffffffffff000000000a0a0a3b;

	lut_sub lut_2409 ({sk[737], g, h, j, x30x, n_n982, x47x}, x5385x);
	defparam lut_2409.LUT_SIZE = 7;
	defparam lut_2409.mask = 128'h5577ffffffffffff0000000300000011;

	lut_sub lut_2412 ({sk[738], c, d, e, l, n_n1137, n_n1202}, x7500x);
	defparam lut_2412.LUT_SIZE = 7;
	defparam lut_2412.mask = 128'h5577fffffffffffffffffeffffffffff;

	lut_sub lut_2427 ({sk[739], n_n841, n_n700, x216x, x260x, x383x, x7500x}, x5386x);
	defparam lut_2427.LUT_SIZE = 7;
	defparam lut_2427.mask = 128'h5577ffffffffffffaabbaabbaabbafbf;

	lut_sub lut_2431 ({sk[740], n_n711, n_n1155, n_n821, n_n700, x133x, x415x}, x5429x);
	defparam lut_2431.LUT_SIZE = 7;
	defparam lut_2431.mask = 128'h5577ffffffffffff0000050500330537;

	lut_sub lut_2434 ({sk[741], n_n996, n_n1155, n_n1171, n_n857, x27x, x133x}, x5430x);
	defparam lut_2434.LUT_SIZE = 7;
	defparam lut_2434.mask = 128'h5577ffffffffffff0000005503030357;

	lut_sub lut_2437 ({sk[742], x15x, x228x, n_n698, n_n730, x255x, x380x}, x5431x);
	defparam lut_2437.LUT_SIZE = 7;
	defparam lut_2437.mask = 128'h5577ffffffffffff0055035700550055;

	lut_sub lut_2440 ({sk[743], n_n709, n_n933, n_n821, n_n824, x133x, x309x}, x5432x);
	defparam lut_2440.LUT_SIZE = 7;
	defparam lut_2440.mask = 128'h5577ffffffffffff0000111103001311;

	lut_sub lut_2443 ({sk[744], m, n, n_n1207, n_n904, x228x, x29x}, x5433x);
	defparam lut_2443.LUT_SIZE = 7;
	defparam lut_2443.mask = 128'h5577ffffffffffff0000000000130000;

	lut_sub lut_2446 ({sk[745], x228x, n_n698, n_n1155, x133x, x210x, x257x}, x5434x);
	defparam lut_2446.LUT_SIZE = 7;
	defparam lut_2446.mask = 128'h5577ffffffffffff0003000300035557;

	lut_sub lut_2449 ({sk[746], f, x314x, x30x, x34x, x133x, x905x}, x5437x);
	defparam lut_2449.LUT_SIZE = 7;
	defparam lut_2449.mask = 128'h5577ffffffffffff5555555555555557;

	lut_sub lut_2452 ({sk[747], h, j, k, x961x, x52x, n_n1204}, x5445x);
	defparam lut_2452.LUT_SIZE = 7;
	defparam lut_2452.mask = 128'h5577ffffffffffff00000000001f1f00;

	lut_sub lut_2457 ({sk[748], m, n, x64x, x228x, n_n996, x238x}, x7488x);
	defparam lut_2457.LUT_SIZE = 7;
	defparam lut_2457.mask = 128'h5577fffffffffffffff0fff0eee0fff0;

	lut_sub lut_2466 ({sk[749], b, x53x, n_n1203, n_n1210, x231x, x296x}, x5458x);
	defparam lut_2466.LUT_SIZE = 7;
	defparam lut_2466.mask = 128'h5577ffffffffffff0055005500550357;

	lut_sub lut_2469 ({sk[750], b, x256x, x53x, n_n1210, x89x, x164x}, x5460x);
	defparam lut_2469.LUT_SIZE = 7;
	defparam lut_2469.mask = 128'h5577ffffffffffff0000030300050005;

	lut_sub lut_2472 ({sk[751], x256x, n_n709, x76x, n_n1095, x196x, x230x}, x5506x);
	defparam lut_2472.LUT_SIZE = 7;
	defparam lut_2472.mask = 128'h5577ffffffffffff0000005500030057;

	lut_sub lut_2475 ({sk[752], x112x, x256x, n_n1229, x74x, x120x, x845x}, x5512x);
	defparam lut_2475.LUT_SIZE = 7;
	defparam lut_2475.mask = 128'h5577ffffffffffff5555555555555755;

	lut_sub lut_2478 ({sk[753], b, x171x, x75x, x84x, x393x, n_n1104}, x7486x);
	defparam lut_2478.LUT_SIZE = 7;
	defparam lut_2478.mask = 128'h5577fffffffffffffcccfcccfcccf8c8;

	lut_sub lut_2484 ({sk[754], c, d, e, n}, x5526x);
	defparam lut_2484.LUT_SIZE = 5;
	defparam lut_2484.mask = 32'h5fff0020;

	lut_sub lut_2486 ({sk[755], c, n, n_n1207, x53x, n_n1116, x5530x}, x5558x);
	defparam lut_2486.LUT_SIZE = 7;
	defparam lut_2486.mask = 128'h5577ffffffffffff0000000005070000;

	lut_sub lut_2489 ({sk[756], g, i, j, x58x, n_n1171, x813x}, x5559x);
	defparam lut_2489.LUT_SIZE = 7;
	defparam lut_2489.mask = 128'h5577ffffffffffff5555555555555557;

	lut_sub lut_2492 ({sk[757], n_n868, x396x, n_n1171, x77x, x290x, n_n1148}, x5560x);
	defparam lut_2492.LUT_SIZE = 7;
	defparam lut_2492.mask = 128'h5577ffffffffffff0000050500330537;

	lut_sub lut_2495 ({sk[758], k, n_n1187, n_n698, n_n1171, n_n1142, n_n694}, x5561x);
	defparam lut_2495.LUT_SIZE = 7;
	defparam lut_2495.mask = 128'h5577ffffffffffff0000000000000777;

	lut_sub lut_2500 ({sk[759], g, h, i, x54x, n_n1171, x829x}, x5564x);
	defparam lut_2500.LUT_SIZE = 7;
	defparam lut_2500.mask = 128'h5577ffffffffffff5555555755555555;

	lut_sub lut_2503 ({sk[760], n_n698, n_n700, n_n1190, n_n1219, n_n1131, n_n817}, x5565x);
	defparam lut_2503.LUT_SIZE = 7;
	defparam lut_2503.mask = 128'h5577ffffffffffff0000005503030357;

	lut_sub lut_2506 ({sk[761], n_n698, n_n841, n_n1203, n_n1190, n_n1215, n_n817}, x5566x);
	defparam lut_2506.LUT_SIZE = 7;
	defparam lut_2506.mask = 128'h5577ffffffffffff0005000500053337;

	lut_sub lut_2509 ({sk[762], e, g, h, n_n713, x396x, x293x}, x5568x);
	defparam lut_2509.LUT_SIZE = 7;
	defparam lut_2509.mask = 128'h5577ffffffffffff0000000500000011;

	lut_sub lut_2512 ({sk[763], n_n840, n_n1201, n_n841, x260x, x293x, x109x}, x5569x);
	defparam lut_2512.LUT_SIZE = 7;
	defparam lut_2512.mask = 128'h5577ffffffffffff0005000500053337;

	lut_sub lut_2515 ({sk[764], g, h, i, j, n_n1191, x109x}, x5570x);
	defparam lut_2515.LUT_SIZE = 7;
	defparam lut_2515.mask = 128'h5577ffffffffffff0000000000111110;

	lut_sub lut_2519 ({sk[765], k, n_n1165, n_n1137, n_n1131, x410x, x109x}, x5571x);
	defparam lut_2519.LUT_SIZE = 7;
	defparam lut_2519.mask = 128'h5577ffffffffffff0303035703030303;

	lut_sub lut_2522 ({sk[766], n_n840, n_n713, x172x, n_n1201, x77x, n_n1196}, x5574x);
	defparam lut_2522.LUT_SIZE = 7;
	defparam lut_2522.mask = 128'h5577ffffffffffff00001155030f135f;

	lut_sub lut_2527 ({sk[767], n, n_n1116, x93x, x841x, x5557x, x135x}, x5577x);
	defparam lut_2527.LUT_SIZE = 7;
	defparam lut_2527.mask = 128'h5577ffffffffffff0055005500553f7f;

	lut_sub lut_2531 ({sk[768], c, n_n1207, x53x, n_n893, n_n1165, x785x}, x5607x);
	defparam lut_2531.LUT_SIZE = 7;
	defparam lut_2531.mask = 128'h5577ffffffffffff5555555555555557;

	lut_sub lut_2534 ({sk[769], i, j, k, x29x, x147x, x786x}, x5608x);
	defparam lut_2534.LUT_SIZE = 7;
	defparam lut_2534.mask = 128'h5577ffffffffffff5555555555555755;

	lut_sub lut_2537 ({sk[770], f, n_n893, x148x, n_n698, x194x, x788x}, x5609x);
	defparam lut_2537.LUT_SIZE = 7;
	defparam lut_2537.mask = 128'h5577ffffffffffff5555555555555557;

	lut_sub lut_2540 ({sk[771], m, n, n_n893, x148x, x106x, x246x}, x5611x);
	defparam lut_2540.LUT_SIZE = 7;
	defparam lut_2540.mask = 128'h5577ffffffffffff0003000311130003;

	lut_sub lut_2543 ({sk[772], g, x76x, x132x, x33x, x93x, x402x}, x5612x);
	defparam lut_2543.LUT_SIZE = 7;
	defparam lut_2543.mask = 128'h5577ffffffffffff0505050505050537;

	lut_sub lut_2546 ({sk[773], x148x, x22x, x113x, x156x, x203x}, x5613x);
	defparam lut_2546.LUT_SIZE = 6;
	defparam lut_2546.mask = 64'h5f7f5f7f05553777;

	lut_sub lut_2550 ({sk[774], n_n1207, x148x, x83x, x219x, x246x, x402x}, x7485x);
	defparam lut_2550.LUT_SIZE = 7;
	defparam lut_2550.mask = 128'h5577fffffffffffffff3fff3fff3aaa2;

	lut_sub lut_2560 ({sk[775], n, x415x, n_n1138, n_n1142, n_n1118, x407x}, x5706x);
	defparam lut_2560.LUT_SIZE = 7;
	defparam lut_2560.mask = 128'h5577ffffffffffff0011001f0000000f;

	lut_sub lut_2563 ({sk[776], a, b, c, x195x, n_n1220, n_n1082}, x5707x);
	defparam lut_2563.LUT_SIZE = 7;
	defparam lut_2563.mask = 128'h5577ffffffffffff00000011000f0000;

	lut_sub lut_2566 ({sk[777], a, b, c, e, g, x45x}, x7498x);
	defparam lut_2566.LUT_SIZE = 7;
	defparam lut_2566.mask = 128'h5577fffffffffffffffffffeffffffff;

	lut_sub lut_2581 ({sk[778], c, d, x120x, x387x, x200x, x7498x}, x5710x);
	defparam lut_2581.LUT_SIZE = 7;
	defparam lut_2581.mask = 128'h5577ffffffffffffaaaaaaaaaaaaaaab;

	lut_sub lut_2584 ({sk[779], a, b, c, d, e, x138x}, x5711x);
	defparam lut_2584.LUT_SIZE = 7;
	defparam lut_2584.mask = 128'h5577ffffffffffff0000000000550010;

	lut_sub lut_2587 ({sk[780], j, k, l, n_n1252, n_n987, x111x}, x5730x);
	defparam lut_2587.LUT_SIZE = 7;
	defparam lut_2587.mask = 128'h5577ffffffffffff0000050000150000;

	lut_sub lut_2591 ({sk[781], i, j, k, l, x223x, x388x}, x5731x);
	defparam lut_2591.LUT_SIZE = 7;
	defparam lut_2591.mask = 128'h5577ffffffffffff0000770700000000;

	lut_sub lut_2596 ({sk[782], i, k, n_n1080, n_n1190, n_n1039, x645x}, x5788x);
	defparam lut_2596.LUT_SIZE = 7;
	defparam lut_2596.mask = 128'h5577ffffffffffff5557555555555555;

	lut_sub lut_2599 ({sk[783], f, n_n920, x306x, n_n977, n_n987, x111x}, x5789x);
	defparam lut_2599.LUT_SIZE = 7;
	defparam lut_2599.mask = 128'h5577ffffffffffff01010101010101ff;

	lut_sub lut_2602 ({sk[784], n_n842, n_n1252, n_n838, n_n1210, x89x, x164x}, x5790x);
	defparam lut_2602.LUT_SIZE = 7;
	defparam lut_2602.mask = 128'h5577ffffffffffff0003000005070505;

	lut_sub lut_2605 ({sk[785], n_n1080, n_n971, x141x, n_n1210, n_n988, x89x}, x5791x);
	defparam lut_2605.LUT_SIZE = 7;
	defparam lut_2605.mask = 128'h5577ffffffffffff01010101010101ff;

	lut_sub lut_2608 ({sk[786], x75x, x265x, n_n876, n_n864, x697x, x167x}, x5792x);
	defparam lut_2608.LUT_SIZE = 7;
	defparam lut_2608.mask = 128'h5577ffffffffffff0000333f5555777f;

	lut_sub lut_2612 ({sk[787], n_n1252, n_n933, n_n977, x111x, x18x, x5789x}, x5794x);
	defparam lut_2612.LUT_SIZE = 7;
	defparam lut_2612.mask = 128'h5577ffffffffffff55555555575f5f5f;

	lut_sub lut_2617 ({sk[788], n_n1252, n_n838, x39x, n_n987, x111x, x117x}, x5795x);
	defparam lut_2617.LUT_SIZE = 7;
	defparam lut_2617.mask = 128'h5577ffffffffffff0003555700030003;

	lut_sub lut_2620 ({sk[789], n_n842, n_n988, x893x, x135x, n_n1036, n_n823}, x5797x);
	defparam lut_2620.LUT_SIZE = 7;
	defparam lut_2620.mask = 128'h5577ffffffffffff000011ff0f0f1fff;

	lut_sub lut_2624 ({sk[790], a, c, d, e, x151x, x200x}, x7482x);
	defparam lut_2624.LUT_SIZE = 7;
	defparam lut_2624.mask = 128'h5577fffffffffffffffffffffaccfaff;

	lut_sub lut_2634 ({sk[791], x259x, x38x, x46x, x27x, x92x, x5730x}, x7481x);
	defparam lut_2634.LUT_SIZE = 7;
	defparam lut_2634.mask = 128'h5577ffffffffffffaaaa8888aaa08880;

	lut_sub lut_2641 ({sk[792], n_n698, n_n1155, n_n1210, x213x, x1202x, x1203x}, x5825x);
	defparam lut_2641.LUT_SIZE = 7;
	defparam lut_2641.mask = 128'h5577ffffffffffff0000000f7777777f;

	lut_sub lut_2645 ({sk[793], k, n_n1207, n_n1187, n_n698, n_n841, x402x}, x5841x);
	defparam lut_2645.LUT_SIZE = 7;
	defparam lut_2645.mask = 128'h5577ffffffffffff0000000000030057;

	lut_sub lut_2648 ({sk[794], i, n_n1220, x29x, x147x, x156x, n_n605}, x5842x);
	defparam lut_2648.LUT_SIZE = 7;
	defparam lut_2648.mask = 128'h5577ffffffffffff0005000500053337;

	lut_sub lut_2651 ({sk[795], j, k, l, n_n1187, x219x, x402x}, x5843x);
	defparam lut_2651.LUT_SIZE = 7;
	defparam lut_2651.mask = 128'h5577ffffffffffff0000050533000000;

	lut_sub lut_2654 ({sk[796], n_n920, x15x, n_n698, x147x, x81x, x5831x}, x5847x);
	defparam lut_2654.LUT_SIZE = 7;
	defparam lut_2654.mask = 128'h5577ffffffffffff0077077707770777;

	lut_sub lut_2661 ({sk[797], g, h, i, j, n_n700, n_n1191}, x5860x);
	defparam lut_2661.LUT_SIZE = 7;
	defparam lut_2661.mask = 128'h5577ffffffffffff0000000000001110;

	lut_sub lut_2664 ({sk[798], f, h, j, n_n920, x264x, x192x}, x5861x);
	defparam lut_2664.LUT_SIZE = 7;
	defparam lut_2664.mask = 128'h5577ffffffffffff0303030303035703;

	lut_sub lut_2667 ({sk[799], i, x258x, x210x, x113x, x14x, x266x}, x5862x);
	defparam lut_2667.LUT_SIZE = 7;
	defparam lut_2667.mask = 128'h5577ffffffffffff0011001100110f1f;

	lut_sub lut_2670 ({sk[800], n_n711, n_n1142, n_n987, x14x, x70x, x266x}, x5863x);
	defparam lut_2670.LUT_SIZE = 7;
	defparam lut_2670.mask = 128'h5577ffffffffffff0005000500053337;

	lut_sub lut_2673 ({sk[801], n, x210x, x113x, x203x, n_n992, n_n1227}, x5864x);
	defparam lut_2673.LUT_SIZE = 7;
	defparam lut_2673.mask = 128'h5577ffffffffffff000f000f000f111f;

	lut_sub lut_2676 ({sk[802], n_n904, n_n918, n_n730, n_n987, x266x, x5860x}, x5865x);
	defparam lut_2676.LUT_SIZE = 7;
	defparam lut_2676.mask = 128'h5577ffffffffffff5555557775757577;

	lut_sub lut_2680 ({sk[803], x22x, n_n996, n_n1155, x14x, x315x, n_n1084}, x5893x);
	defparam lut_2680.LUT_SIZE = 7;
	defparam lut_2680.mask = 128'h5577ffffffffffff0000003305050537;

	lut_sub lut_2683 ({sk[804], f, n_n904, x22x, n_n730, x29x, x146x}, x5894x);
	defparam lut_2683.LUT_SIZE = 7;
	defparam lut_2683.mask = 128'h5577ffffffffffff0004000400040055;

	lut_sub lut_2686 ({sk[805], x22x, n_n918, n_n1053, n_n992, x293x, x5880x}, x5895x);
	defparam lut_2686.LUT_SIZE = 7;
	defparam lut_2686.mask = 128'h5577ffffffffffff0003000300035557;

	lut_sub lut_2689 ({sk[806], k, n_n920, x15x, n_n996, x147x, x146x}, x5896x);
	defparam lut_2689.LUT_SIZE = 7;
	defparam lut_2689.mask = 128'h5577ffffffffffff0023032300030303;

	lut_sub lut_2693 ({sk[807], f, x22x, x29x, x146x, n_n2953, x369x}, x5897x);
	defparam lut_2693.LUT_SIZE = 7;
	defparam lut_2693.mask = 128'h5577ffffffffffff333333333333373f;

	lut_sub lut_2697 ({sk[808], g, n_n1171, x122x, x221x, x47x, x155x}, x7479x);
	defparam lut_2697.LUT_SIZE = 7;
	defparam lut_2697.mask = 128'h5577fffffffffffffafafafaf8faf0fa;

	lut_sub lut_2702 ({sk[809], k, n_n1187, n_n730, n_n1053, n_n816, x539x}, x5919x);
	defparam lut_2702.LUT_SIZE = 7;
	defparam lut_2702.mask = 128'h5577ffffffffffff5555555555555575;

	lut_sub lut_2705 ({sk[810], h, i, j, k, n_n1177, n_n671}, x5920x);
	defparam lut_2705.LUT_SIZE = 7;
	defparam lut_2705.mask = 128'h5577ffffffffffff0000010100000010;

	lut_sub lut_2708 ({sk[811], c, x196x, n_n841, n_n1053, n_n1210, n_n1085}, x5921x);
	defparam lut_2708.LUT_SIZE = 7;
	defparam lut_2708.mask = 128'h5577ffffffffffff0003000300031113;

	lut_sub lut_2711 ({sk[812], k, n_n1187, n_n904, n_n698, n_n1194, n_n816}, x5922x);
	defparam lut_2711.LUT_SIZE = 7;
	defparam lut_2711.mask = 128'h5577ffffffffffff0000050500000537;

	lut_sub lut_2714 ({sk[813], h, j, k, n_n841, x304x, x315x}, x5923x);
	defparam lut_2714.LUT_SIZE = 7;
	defparam lut_2714.mask = 128'h5577ffffffffffff0303030303570303;

	lut_sub lut_2717 ({sk[814], e, x171x, x230x, x21x, x126x, x290x}, x5924x);
	defparam lut_2717.LUT_SIZE = 7;
	defparam lut_2717.mask = 128'h5577ffffffffffff0033053700330033;

	lut_sub lut_2720 ({sk[815], x34x, x230x, n_n1202, n_n1264, x192x, x48x}, x5925x);
	defparam lut_2720.LUT_SIZE = 7;
	defparam lut_2720.mask = 128'h5577ffffffffffff00001111000f111f;

	lut_sub lut_2723 ({sk[816], g, h, i, x36x, x70x, x48x}, x5926x);
	defparam lut_2723.LUT_SIZE = 7;
	defparam lut_2723.mask = 128'h5577ffffffffffff0000001100000003;

	lut_sub lut_2726 ({sk[817], e, h, i, j, k, x263x}, x7501x);
	defparam lut_2726.LUT_SIZE = 7;
	defparam lut_2726.mask = 128'h5577ffffffffffffffffffbfffffffff;

	lut_sub lut_2742 ({sk[818], d, f, m, n, x373x, x7501x}, x5965x);
	defparam lut_2742.LUT_SIZE = 7;
	defparam lut_2742.mask = 128'h5577ffffffffffffaaaaaaaaaabaaaaa;

	lut_sub lut_2745 ({sk[819], x222x, x78x, n_n1036, x312x, n_n1196, x273x}, x5966x);
	defparam lut_2745.LUT_SIZE = 7;
	defparam lut_2745.mask = 128'h5577ffffffffffff0022002200220f2f;

	lut_sub lut_2748 ({sk[820], c, g, h, j, n_n1165, n_n1159}, x7477x);
	defparam lut_2748.LUT_SIZE = 7;
	defparam lut_2748.mask = 128'h5577ffffffffffffffffffffffefffff;

	lut_sub lut_2764 ({sk[821], m, n, n_n1137, n_n700, n_n1203, n_n1195}, x7478x);
	defparam lut_2764.LUT_SIZE = 7;
	defparam lut_2764.mask = 128'h5577ffffffffffffffbfffffffffffff;

	lut_sub lut_2780 ({sk[822], f, h, i, n_n1165, n_n1203, n_n1227}, x6057x);
	defparam lut_2780.LUT_SIZE = 7;
	defparam lut_2780.mask = 128'h5577ffffffffffff0300000003550000;

	lut_sub lut_2783 ({sk[823], h, i, n_n1161, n_n1165, n_n857, x395x}, x6058x);
	defparam lut_2783.LUT_SIZE = 7;
	defparam lut_2783.mask = 128'h5577ffffffffffff0005040400000000;

	lut_sub lut_2786 ({sk[824], m, x255x, x367x, x386x, n_n1204, x95x}, x6059x);
	defparam lut_2786.LUT_SIZE = 7;
	defparam lut_2786.mask = 128'h5577ffffffffffff0022032300220022;

	lut_sub lut_2789 ({sk[825], h, n, x226x, n_n1190, n_n1118, x95x}, x6060x);
	defparam lut_2789.LUT_SIZE = 7;
	defparam lut_2789.mask = 128'h5577ffffffffffff1115000500050005;

	lut_sub lut_2792 ({sk[826], c, d, e, x132x, x367x, x70x}, x6061x);
	defparam lut_2792.LUT_SIZE = 7;
	defparam lut_2792.mask = 128'h5577ffffffffffff0500373305000500;

	lut_sub lut_2795 ({sk[827], h, n, n_n1161, x189x, n_n1227, x285x}, x6062x);
	defparam lut_2795.LUT_SIZE = 7;
	defparam lut_2795.mask = 128'h5577ffffffffffff0055035700550055;

	lut_sub lut_2798 ({sk[828], i, j, n_n1210, x103x, n_n1253, x449x}, x6093x);
	defparam lut_2798.LUT_SIZE = 7;
	defparam lut_2798.mask = 128'h5577ffffffffffff5557555555575557;

	lut_sub lut_2802 ({sk[829], f, n_n1188, n_n1193, x120x, x373x, x302x}, x6094x);
	defparam lut_2802.LUT_SIZE = 7;
	defparam lut_2802.mask = 128'h5577ffffffffffff0357030300550000;

	lut_sub lut_2805 ({sk[830], x189x, x194x, n_n1138, x141x, n_n1253, x145x}, x6095x);
	defparam lut_2805.LUT_SIZE = 7;
	defparam lut_2805.mask = 128'h5577ffffffffffff00000f0044444f44;

	lut_sub lut_2808 ({sk[831], i, j, l, x112x, n_n1165, n_n1229}, x6096x);
	defparam lut_2808.LUT_SIZE = 7;
	defparam lut_2808.mask = 128'h5577ffffffffffff0001000101010000;

	lut_sub lut_2811 ({sk[832], l, n_n1177, x196x, n_n1217, n_n1264, x432x}, x6128x);
	defparam lut_2811.LUT_SIZE = 7;
	defparam lut_2811.mask = 128'h5577ffffffffffff5555555555555557;

	lut_sub lut_2814 ({sk[833], e, f, h, j, x144x, x434x}, x6129x);
	defparam lut_2814.LUT_SIZE = 7;
	defparam lut_2814.mask = 128'h5577ffffffffffff7555555555555555;

	lut_sub lut_2817 ({sk[834], a, d, e, f, g, h}, x7473x);
	defparam lut_2817.LUT_SIZE = 7;
	defparam lut_2817.mask = 128'h5577fffffffffffffefefefefefefeff;

	lut_sub lut_2822 ({sk[835], h, i, n_n1252, x144x, x288x, x7473x}, x6134x);
	defparam lut_2822.LUT_SIZE = 7;
	defparam lut_2822.mask = 128'h5577ffffffffffff2222222f22222222;

	lut_sub lut_2825 ({sk[836], e, g, j, x131x, x204x, x286x}, x6161x);
	defparam lut_2825.LUT_SIZE = 7;
	defparam lut_2825.mask = 128'h5577ffffffffffff5d5d5d0c55555500;

	lut_sub lut_2829 ({sk[837], c, d, n_n1190, x68x, x287x, x416x}, x6164x);
	defparam lut_2829.LUT_SIZE = 7;
	defparam lut_2829.mask = 128'h5577ffffffffffff05cd050505050505;

	lut_sub lut_2832 ({sk[838], a, b, g, j, n_n1222, x340x}, x6198x);
	defparam lut_2832.LUT_SIZE = 7;
	defparam lut_2832.mask = 128'h5577ffffffffffff5755555557555755;

	lut_sub lut_2836 ({sk[839], x120x, n_n1039, x407x, n_n1191, n_n1072, x348x}, x6202x);
	defparam lut_2836.LUT_SIZE = 7;
	defparam lut_2836.mask = 128'h5577ffffffffffff555f555f777fffff;

	lut_sub lut_2841 ({sk[840], c, d, e, f, g, i}, x7476x);
	defparam lut_2841.LUT_SIZE = 7;
	defparam lut_2841.mask = 128'h5577ffffffffffffbebebfbfffffffff;

	lut_sub lut_2861 ({sk[841], f, g, j, x131x, x127x, x253x}, x6275x);
	defparam lut_2861.LUT_SIZE = 7;
	defparam lut_2861.mask = 128'h5577ffffffffffff5555575755555755;

	lut_sub lut_2865 ({sk[842], n, x114x, n_n1118, x146x, x127x, n_n1091}, x6276x);
	defparam lut_2865.LUT_SIZE = 7;
	defparam lut_2865.mask = 128'h5577ffffffffffff000c00ae000c000c;

	lut_sub lut_2868 ({sk[843], x114x, n_n1080, n_n1082, x146x, n_n1036, x127x}, x6277x);
	defparam lut_2868.LUT_SIZE = 7;
	defparam lut_2868.mask = 128'h5577ffffffffffff0003555700030003;

	lut_sub lut_2871 ({sk[844], h, n_n1194, n_n1202, x127x, n_n1167, n_n819}, x6278x);
	defparam lut_2871.LUT_SIZE = 7;
	defparam lut_2871.mask = 128'h5577ffffffffffff0000005503030357;

	lut_sub lut_2874 ({sk[845], g, h, x189x, n_n1202, n_n694, x418x}, x6279x);
	defparam lut_2874.LUT_SIZE = 7;
	defparam lut_2874.mask = 128'h5577ffffffffffff5555000300000003;

	lut_sub lut_2877 ({sk[846], c, d, f, g, h, i}, x7475x);
	defparam lut_2877.LUT_SIZE = 7;
	defparam lut_2877.mask = 128'h5577ffffffffffffcaf0caffffffffff;

	lut_sub lut_2889 ({sk[847], g, n_n1202, n_n1118, x127x, x395x, x7475x}, x6280x);
	defparam lut_2889.LUT_SIZE = 7;
	defparam lut_2889.mask = 128'h5577ffffffffffff03000b0a00000a0a;

	lut_sub lut_2892 ({sk[848], k, m, n, x114x, x57x, x146x}, x6292x);
	defparam lut_2892.LUT_SIZE = 7;
	defparam lut_2892.mask = 128'h5577ffffffffffff00110f0000000f00;

	lut_sub lut_2895 ({sk[849], f, x131x, n_n1202, x146x, n_n1036, x268x}, x6294x);
	defparam lut_2895.LUT_SIZE = 7;
	defparam lut_2895.mask = 128'h5577ffffffffffff000a0000030b0303;

	lut_sub lut_2898 ({sk[850], c, d, i, n_n1165, x222x, x312x}, x6295x);
	defparam lut_2898.LUT_SIZE = 7;
	defparam lut_2898.mask = 128'h5577ffffffffffff1311111111110000;

	lut_sub lut_2902 ({sk[851], j, k, l, m, n, x6292x}, x6296x);
	defparam lut_2902.LUT_SIZE = 7;
	defparam lut_2902.mask = 128'h5577ffffffffffff5d55555555555555;

	lut_sub lut_2905 ({sk[852], a, b, c, m, n, x6294x}, x6297x);
	defparam lut_2905.LUT_SIZE = 7;
	defparam lut_2905.mask = 128'h5577ffffffffffff7d5d555575555555;

	lut_sub lut_2909 ({sk[853], x6149x, x6150x, x6295x, x6296x, x6297x}, x6301x);
	defparam lut_2909.LUT_SIZE = 6;
	defparam lut_2909.mask = 64'h5f7f5f7f7fffffff;

	lut_sub lut_2915 ({sk[854], x5970x, x5965x, x5966x, x6128x, x6129x, x6134x}, x7472x);
	defparam lut_2915.LUT_SIZE = 7;
	defparam lut_2915.mask = 128'h5577ffffffffffff8000000000000000;

	lut_sub lut_2917 ({sk[855], c, d, f, x415x, n_n1142, x42x}, x6316x);
	defparam lut_2917.LUT_SIZE = 7;
	defparam lut_2917.mask = 128'h5577ffffffffffff5755555555555555;


endmodule