module spla (
	i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, 
	i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, i_14_, i_15_, o_0_, o_1_, 
	o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, 
	o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_, o_21_, 
	o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_, o_31_, 
	o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_, o_41_, 
	o_42_, o_43_, o_44_, o_45_);

input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_, i_11_, i_12_, i_13_, i_14_, i_15_;

output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_, o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_, o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_, o_41_, o_42_, o_43_, o_44_, o_45_;

wire n3, n7, n14, n13, n11, n15, n20, n19, n23, n27, n32, n29, n35, n33, n37, n38, n36, n39, n40, n42, n43, n44, n46, n47, n48, n49, n41, n51, n52, n53, n50, n55, n56, n54, n57, n58, n59, n60, n61, n65, n66, n67, n68, n69, n70, n62, n72, n73, n71, n74, n75, n76, n77, n78, n79, n80, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n95, n97, n98, n99, n101, n93, n102, n103, n104, n105, n106, n108, n110, n112, n113, n114, n115, n116, n117, n118, n119, n111, n121, n122, n123, n124, n120, n125, n126, n127, n129, n128, n130, n134, n135, n136, n133, n139, n143, n140, n144, n147, n151, n150, n156, n154, n160, n157, n161, n166, n167, n164, n165, n163, n169, n170, n171, n172, n173, n174, n168, n176, n177, n178, n179, n175, n182, n180, n181, n184, n185, n187, n183, n192, n188, n193, n198, n197, n203, n204, n205, n206, n207, n208, n209, n210, n202, n212, n211, n216, n217, n215, n214, n221, n219, n220, n218, n223, n222, n229, n225, n233, n230, n237, n236, n234, n239, n240, n238, n243, n244, n245, n246, n247, n248, n249, n250, n242, n251, n254, n255, n256, n257, n258, n259, n260, n261, n253, n263, n262, n265, n266, n264, n268, n269, n270, n271, n272, n273, n274, n275, n267, n277, n276, n280, n281, n282, n283, n284, n285, n286, n287, n279, n289, n290, n291, n292, n293, n294, n295, n296, n288, n298, n299, n300, n301, n302, n303, n304, n305, n297, n307, n308, n306, n312, n313, n310, n317, n315, n316, n314, n319, n318, n321, n322, n323, n324, n325, n326, n327, n328, n320, n330, n329, n333, n331, n337, n338, n335, n334, n340, n341, n339, n343, n342, n347, n344, n350, n349, n348, n351, n356, n354, n357, n358, n359, n360, n361, n362, n363, n364, n367, n368, n366, n365, n371, n372, n370, n369, n375, n376, n374, n373, n378, n379, n377, n382, n383, n381, n380, n385, n386, n384, n389, n390, n388, n387, n392, n391, n394, n395, n396, n397, n398, n399, n393, n401, n400, n404, n405, n406, n407, n408, n409, n410, n411, n403, n412, n415, n416, n417, n418, n419, n420, n421, n422, n414, n425, n424, n423, n428, n429, n427, n426, n432, n431, n430, n435, n436, n434, n433, n439, n437, n442, n443, n441, n440, n445, n446, n444, n448, n449, n447, n451, n452, n450, n454, n453, n456, n455, n458, n459, n460, n457, n462, n464, n461, n466, n465, n468, n467, n470, n471, n472, n469, n473, n476, n482, n479, n486, n483, n487, n490, n491, n492, n493, n494, n495, n496, n497, n489, n499, n500, n498, n503, n504, n505, n506, n509, n507, n508, n511, n510, n514, n513, n512, n517, n515, n520, n519, n525, n524, n522, n526, n527, n531, n530, n533, n538, n537, n536, n539, n541, n540, n544, n545, n546, n547, n548, n549, n543, n552, n553, n550, n555, n554, n559, n560, n561, n562, n563, n564, n557, n565, n570, n567, n572, n571, n574, n573, n577, n578, n575, n580, n581, n582, n583, n584, n585, n586, n587, n579, n588, n591, n592, n590, n589, n594, n595, n596, n597, n598, n599, n600, n601, n593, n602, n603, n604, n605, n609, n608, n606, n611, n612, n610, n614, n613, n615, n617, n616, n619, n618, n620, n623, n624, n622, n621, n626, n625, n628, n627, n631, n632, n630, n629, n635, n636, n634, n633, n639, n640, n638, n637, n642, n643, n641, n647, n645, n646, n644, n649, n648, n652, n651, n650, n654, n656, n657, n658, n653, n660, n661, n662, n663, n664, n665, n659, n667, n666, n669, n670, n668, n673, n671, n675, n674, n677, n678, n679, n680, n676, n681, n683, n686, n692, n688, n693, n699, n696, n701, n702, n700, n703, n707, n706, n709, n710, n711, n712, n713, n714, n715, n716, n708, n718, n717, n719, n723, n722, n721, n725, n726, n727, n724, n732, n728, n734, n733, n736, n737, n738, n739, n740, n741, n742, n743, n735, n745, n746, n744, n748, n749, n750, n751, n747, n753, n754, n755, n756, n757, n752, n759, n761, n762, n758, n765, n763, n767, n768, n769, n770, n772, n773, n771, n774, n776, n778, n775, n782, n783, n780, n781, n779, n785, n784, n786, n790, n789, n794, n793, n791, n796, n795, n799, n798, n800, n801, n804, n803, n802, n806, n807, n805, n809, n810, n811, n812, n808, n814, n815, n816, n817, n819, n813, n821, n822, n820, n824, n823, n828, n826, n827, n825, n829, n831, n832, n833, n834, n835, n836, n837, n838, n830, n839, n842, n840, n845, n846, n844, n843, n848, n847, n849, n855, n854, n852, n856, n858, n861, n864, n863, n865, n867, n868, n869, n870, n871, n872, n873, n874, n866, n876, n877, n875, n881, n878, n885, n883, n882, n888, n887, n886, n892, n893, n890, n891, n889, n895, n896, n897, n898, n894, n900, n901, n902, n903, n904, n905, n906, n907, n899, n908, n909, n911, n912, n913, n914, n915, n910, n917, n916, n919, n920, n918, n922, n921, n924, n925, n926, n927, n928, n929, n930, n923, n932, n933, n931, n935, n934, n938, n937, n941, n940, n939, n943, n944, n945, n946, n947, n948, n949, n942, n950, n952, n953, n954, n955, n956, n957, n958, n960, n961, n959, n963, n962, n966, n967, n964, n968, n970, n975, n973, n976, n977, n981, n982, n983, n984, n985, n986, n987, n988, n980, n990, n992, n993, n989, n995, n994, n997, n998, n996, n999, n1002, n1004, n1007, n1009, n1008, n1011, n1010, n1012, n1014, n1016, n1017, n1018, n1019, n1020, n1021, n1023, n1024, n1025, n1026, n1027, n1028, n1032, n1033, n1034, n1038, n1039, n1040, n1041, n1042, n1043, n1045, n1051, n1050, n1056, n1054, n1060, n1057, n1058, n1062, n1063, n1064, n1065, n1066, n1061, n1068, n1069, n1070, n1071, n1067, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1081, n1082, n1083, n1080, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1084, n1094, n1095, n1096, n1097, n1098, n1099, n1093, n1102, n1100, n1105, n1103, n1108, n1109, n1110, n1107, n1111, n1112, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1116, n1124, n1126, n1127, n1128, n1125, n1130, n1129, n1131, n1138, n1135, n1140, n1139, n1143, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1145, n1154, n1155, n1157, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1178, n1180, n1182, n1184, n1189, n1190, n1191, n1194, n1195, n1198, n1200, n1202, n1203, n1204, n1206, n1205, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1222, n1223, n1224, n1226, n1227, n1228, n1229, n1230, n1231, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1252, n1253, n1254, n1255, n1256, n1257, n1259, n1260, n1261, n1258, n1263, n1264, n1262, n1265, n1267, n1268, n1269, n1270, n1271, n1272, n1274, n1275, n1277, n1276, n1278, n1279, n1280, n1281, n1282, n1283, n1285, n1286, n1287, n1284, n1288, n1289, n1290, n1292, n1293, n1294, n1295, n1291, n1297, n1298, n1299, n1300, n1301, n1302, n1296, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1303, n1311, n1312, n1313, n1314, n1315, n1316, n1318, n1317, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1327, n1328, n1326, n1329, n1330, n1331, n1332, n1333, n1334, n1336, n1337, n1338, n1335, n1339, n1340, n1341, n1342, n1344, n1345, n1346, n1343, n1347, n1349, n1350, n1351, n1352, n1348, n1353, n1354, n1355, n1356, n1358, n1359, n1360, n1357, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1370, n1371, n1372, n1373, n1374, n1375, n1369, n1376, n1377, n1379, n1380, n1381, n1382, n1378, n1383, n1384, n1385, n1386, n1388, n1389, n1391, n1392, n1393, n1394, n1395, n1390, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1427, n1428, n1429, n1430, n1431, n1426, n1433, n1434, n1435, n1436, n1437, n1438, n1432, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1439, n1448, n1449, n1450, n1451, n1452, n1453, n1447, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1472, n1473, n1474, n1475, n1471, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1476, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1485, n1494, n1495, n1497, n1498, n1499, n1500, n1502, n1503, n1501, n1505, n1506, n1504, n1507, n1508, n1509, n1510, n1511, n1512, n1514, n1515, n1516, n1517, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1535, n1534, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1537, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1554, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1608, n1607, n1610, n1611, n1609, n1613, n1614, n1615, n1616, n1617, n1618, n1612, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1627, n1635, n1636, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1646, n1647, n1648, n1649, n1645, n1655, n1656, n1650, n1657, n1658, n1660, n1661, n1662, n1659, n1663, n1664, n1666, n1668, n1669, n1670, n1667, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1681, n1682, n1683, n1680, n1685, n1686, n1687, n1688, n1684, n1690, n1691, n1692, n1693, n1694, n1689, n1696, n1697, n1698, n1699, n1700, n1701, n1695, n1703, n1702, n1704, n1705, n1706, n1707, n1708, n1709, n1711, n1712, n1713, n1714, n1715, n1716, n1710, n1718, n1719, n1720, n1717, n1722, n1723, n1721, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1724, n1733, n1735, n1734, n1736, n1738, n1739, n1741, n1743, n1744, n1740, n1745, n1746, n1747, n1749, n1750, n1751, n1752, n1753, n1754, n1748, n1756, n1757, n1759, n1760, n1761, n1763, n1764, n1765, n1766, n1767, n1768, n1762, n1770, n1771, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1795, n1796, n1797, n1798, n1799, n1800, n1794, n1802, n1803, n1804, n1805, n1806, n1807, n1801, n1809, n1811, n1812, n1813, n1808, n1816, n1817, n1814, n1819, n1820, n1821, n1822, n1823, n1824, n1818, n1825, n1828, n1829, n1830, n1831, n1832, n1833, n1826, n1835, n1836, n1837, n1834, n1840, n1842, n1843, n1844, n1845, n1846, n1848, n1847, n1849, n1850, n1851, n1852, n1853, n1856, n1857, n1858, n1859, n1854, n1861, n1862, n1863, n1864, n1860, n1868, n1869, n1870, n1865, n1871, n1872, n1873, n1874, n1875, n1876, n1878, n1879, n1880, n1881, n1882, n1883, n1877, n1887, n1884, n1888, n1891, n1892, n1893, n1894, n1895, n1896, n1890, n1898, n1899, n1901, n1902, n1903, n1905, n1906, n1907, n1908, n1910, n1911, n1912, n1913, n1914, n1909, n1915, n1917, n1918, n1919, n1916, n1920, n1921, n1923, n1924, n1925, n1927, n1929, n1931, n1932, n1933, n1934, n1935, n1928, n1936, n1937, n1938, n1939, n1940, n1941, n1945, n1946, n1947, n1948, n1950, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1951, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1970, n1971, n1972, n1969, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1985, n1986, n1987, n1988, n1989, n1990, n1984, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2004, n2003, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2046, n2047, n2048, n2045, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2061, n2062, n2063, n2064, n2065, n2066, n2060, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2076, n2075, n2077, n2078, n2080, n2079, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2090, n2089, n2092, n2091, n2093, n2094, n2095, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2110, n2111, n2112, n2109, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2131, n2130, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2147, n2148, n2149, n2146, n2151, n2152, n2150, n2153, n2155, n2156, n2154, n2158, n2157, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2168, n2169, n2167, n2170, n2171, n2172, n2173, n2177, n2178, n2176, n2179, n2182, n2181, n2183, n2184, n2186, n2185, n2189, n2190, n2191, n2192, n2193, n2194, n2196, n2195, n2197, n2198, n2199, n2200, n2201, n2203, n2202, n2205, n2206, n2204, n2207, n2209, n2211, n2212, n2213, n2214, n2216, n2217, n2218, n2219, n2221, n2223, n2225, n2228, n2227, n2229, n2230, n2231, n2233, n2232, n2235, n2234, n2237, n2236, n2239, n2240, n2238, n2242, n2241, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2254, n2255, n2256, n2257, n2258, n2259, n2261, n2260, n2262, n2265, n2266, n2268, n2269, n2270, n2272, n2271, n2273, n2275, n2278, n2277, n2279, n2283, n2285, n2284, n2287, n2286, n2288, n2290, n2289, n2292, n2291, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2301, n2302, n2303, n2304, n2305, n2306, n2308, n2307, n2309, n2311, n2312, n2314, n2313, n2315, n2316, n2317, n2319, n2318, n2320, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2336, n2337, n2338, n2340, n2341, n2342, n2343, n2344, n2345, n2347, n2348, n2349, n2351, n2352, n2353, n2354, n2355, n2356, n2358, n2357, n2359, n2360, n2361, n2362, n2363, n2364, n2366, n2367, n2368, n2369, n2375, n2374, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2385, n2387, n2388, n2389, n2390, n2392, n2391, n2393, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2406, n2405, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2431, n2433, n2432, n2436, n2438, n2439, n2441, n2440, n2442, n2446, n2448, n2447, n2449, n2450, n2452, n2454, n2453, n2455, n2456, n2458, n2457, n2460, n2461, n2462, n2463, n2465, n2467, n2468, n2472, n2474, n2475, n2476, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2489, n2488, n2490, n2491, n2492, n2494, n2495, n2496, n2497, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518;

assign o_0_ = ( (~ n139) ) ;
 assign o_1_ = ( (~ n39) ) ;
 assign o_2_ = ( n106  &  (~ n1057)  &  (~ n1180) ) | ( n106  &  (~ n1167)  &  (~ n1180) ) ;
 assign o_3_ = ( (~ n133) ) ;
 assign o_4_ = ( (~ n130) ) ;
 assign o_5_ = ( (~ n557) ) ;
 assign o_6_ = ( (~ n128) ) ;
 assign o_7_ = ( (~ n489) ) ;
 assign o_8_ = ( (~ i_0_)  &  (~ i_1_)  &  i_3_ ) ;
 assign o_9_ = ( (~ n127) ) ;
 assign o_10_ = ( (~ n126) ) ;
 assign o_11_ = ( (~ n125) ) ;
 assign o_12_ = ( (~ n1145) ) ;
 assign o_13_ = ( (~ n120) ) ;
 assign o_14_ = ( (~ n1107) ) ;
 assign o_15_ = ( (~ n1093) ) ;
 assign o_16_ = ( (~ n111) ) ;
 assign o_17_ = ( (~ n1084) ) ;
 assign o_18_ = ( (~ n110) ) ;
 assign o_19_ = ( i_3_  &  (~ i_4_)  &  i_5_  &  n106  &  (~ n1167) ) ;
 assign o_20_ = ( n106  &  n108  &  (~ n1167) ) ;
 assign o_21_ = ( n103 ) | ( n104 ) | ( n105 ) ;
 assign o_22_ = ( (~ n102) ) ;
 assign o_23_ = ( (~ n93) ) ;
 assign o_24_ = ( n90  &  (~ n1178) ) ;
 assign o_25_ = ( n90  &  n91 ) ;
 assign o_26_ = ( n80 ) | ( n85 ) | ( n89 ) | ( n75 ) ;
 assign o_27_ = ( n79 ) | ( n86 ) | ( (~ n95) ) | ( (~ n2457) ) ;
 assign o_28_ = ( n85 ) | ( n86 ) | ( n87 ) | ( n88 ) ;
 assign o_29_ = ( n79 ) | ( n80 ) | ( n82 ) | ( n83 ) | ( n84 ) | ( (~ n95) ) ;
 assign o_30_ = ( (~ n71) ) | ( n74 ) | ( n75 ) | ( n76 ) | ( n77 ) | ( n78 ) ;
 assign o_31_ = ( n1012 ) | ( n1014 ) | ( (~ n1736) ) | ( (~ n2452) ) ;
 assign o_32_ = ( (~ n1010) ) ;
 assign o_33_ = ( (~ n1008) ) ;
 assign o_34_ = ( (~ n71) ) ;
 assign o_35_ = ( (~ n62) ) ;
 assign o_36_ = ( (~ n980) ) ;
 assign o_37_ = ( (~ n61) ) ;
 assign o_38_ = ( (~ n910) ) ;
 assign o_39_ = ( (~ n813) ) ;
 assign o_40_ = ( (~ n60) ) ;
 assign o_41_ = ( n57  &  n58  &  n59 ) ;
 assign o_42_ = ( (~ n54) ) ;
 assign o_43_ = ( (~ n50) ) ;
 assign o_44_ = ( (~ n41) ) ;
 assign o_45_ = ( (~ n40) ) ;
 assign n3 = ( (~ n441)  &  (~ n472) ) | ( (~ n441)  &  (~ n1705) ) ;
 assign n7 = ( (~ n313)  &  (~ n458) ) | ( (~ n313)  &  (~ n1214) ) ;
 assign n14 = ( n552  &  n1210 ) ;
 assign n13 = ( (~ n812) ) | ( (~ n1339) ) ;
 assign n11 = ( n14  &  n13 ) | ( n14  &  (~ n434) ) ;
 assign n15 = ( (~ n827)  &  (~ n887) ) | ( (~ n827)  &  (~ n890) ) ;
 assign n20 = ( n156 ) | ( (~ n219) ) ;
 assign n19 = ( n20  &  (~ n374) ) | ( (~ n374)  &  (~ n810) ) ;
 assign n23 = ( (~ n164)  &  (~ n343) ) | ( (~ n164)  &  (~ n638) ) ;
 assign n27 = ( n14  &  (~ n1214) ) | ( n14  &  (~ n1318) ) ;
 assign n32 = ( (~ n1578) ) | ( (~ n1588) ) ;
 assign n29 = ( n32  &  (~ n374) ) | ( (~ n374)  &  (~ n1262) ) | ( (~ n374)  &  (~ n1343) ) ;
 assign n35 = ( n356 ) | ( (~ n998) ) ;
 assign n33 = ( n35  &  (~ n827) ) | ( (~ n827)  &  (~ n1081) ) ;
 assign n37 = ( n1180 ) | ( (~ n1639) ) ;
 assign n38 = ( i_7_ ) | ( i_6_ ) ;
 assign n36 = ( n37 ) | ( n38 ) ;
 assign n39 = ( (~ n59)  &  n1060 ) | ( n1060  &  n1057 ) | ( n1060  &  n1058 ) ;
 assign n40 = ( n498  &  n675  &  n673 ) | ( n498  &  n675  &  n674 ) ;
 assign n42 = ( n735  &  n752  &  n767  &  n721  &  n724  &  n768  &  n769  &  n770 ) ;
 assign n43 = ( n377  &  (~ n719)  &  n1781  &  n1782  &  n1783  &  n1785  &  n1786  &  n1787 ) ;
 assign n44 = ( n1788  &  n1789  &  n1790  &  n1791  &  n1792  &  n1793  &  n717 ) ;
 assign n46 = ( n298  &  n1777  &  n1778  &  n1779  &  n774  &  n1780 ) ;
 assign n47 = ( n2351  &  n374 ) | ( n2351  &  n1082  &  n1677 ) ;
 assign n48 = ( n1801  &  n1808  &  n1794  &  n708  &  n1814  &  n676  &  n1818 ) ;
 assign n49 = ( (~ n19)  &  (~ n29)  &  n111  &  n2344  &  n2345  &  n2347  &  n2348  &  n2349 ) ;
 assign n41 = ( n42  &  n43  &  n44  &  n46  &  n47  &  n48  &  n49  &  (~ n775) ) ;
 assign n51 = ( (~ n150)  &  n779  &  (~ n791)  &  (~ n795)  &  n1834  &  n1840  &  n1842  &  n1843 ) ;
 assign n52 = ( (~ n401) ) | ( n1226 ) ;
 assign n53 = ( (~ n401) ) | ( n1315 ) ;
 assign n50 = ( n42  &  n51  &  n52  &  n53 ) ;
 assign n55 = ( n121  &  n182  &  n180 ) | ( n121  &  n182  &  n181 ) ;
 assign n56 = ( n122  &  n454  &  n453 ) | ( n122  &  n454  &  n181 ) ;
 assign n54 = ( n55  &  n56 ) ;
 assign n57 = ( (~ i_9_)  &  (~ i_10_)  &  (~ i_11_) ) ;
 assign n58 = ( (~ i_8_)  &  n1230 ) ;
 assign n59 = ( (~ n1180)  &  n1844 ) ;
 assign n60 = ( n799  &  n504  &  n798 ) | ( n799  &  n504  &  n570 ) ;
 assign n61 = ( n724  &  n952  &  n953  &  n954  &  n955  &  n956  &  n957  &  n958 ) ;
 assign n65 = ( n427  &  (~ n1002) ) | ( n773  &  n997  &  (~ n1002) ) ;
 assign n66 = ( n2446  &  n994 ) | ( n2446  &  n780 ) ;
 assign n67 = ( n2447  &  n2449  &  n772 ) | ( n2447  &  n2449  &  n374 ) ;
 assign n68 = ( n329  &  n387  &  n1609  &  n268  &  n1432  &  n1471 ) ;
 assign n69 = ( n830  &  n1909  &  n1928  &  n650  &  n579  &  n1740 ) ;
 assign n70 = ( (~ n33)  &  (~ n999)  &  n1374  &  n2018  &  n2058  &  n2071  &  n2440  &  n2442 ) ;
 assign n62 = ( n65  &  n66  &  n67  &  n68  &  n69  &  n70  &  (~ n1004)  &  (~ n1007) ) ;
 assign n72 = ( n1169  &  n1170  &  n1171  &  n1172  &  n1173  &  n1174  &  n1175  &  n1176 ) ;
 assign n73 = ( n666  &  n659 ) ;
 assign n71 = ( n72  &  n73 ) ;
 assign n74 = ( (~ n511)  &  (~ n1946) ) ;
 assign n75 = ( n1023 ) | ( n1024 ) | ( n1025 ) | ( n1026 ) | ( n1027 ) | ( n1028 ) | ( (~ n2453) ) ;
 assign n76 = ( n1016 ) | ( n1017 ) | ( n1018 ) | ( n1019 ) | ( n1020 ) | ( n1021 ) | ( (~ n2455) ) ;
 assign n77 = ( (~ n500)  &  (~ n511) ) ;
 assign n78 = ( (~ n511)  &  n1657 ) ;
 assign n79 = ( n1941 ) | ( n1945 ) | ( n1646 ) ;
 assign n80 = ( n1647 ) | ( n1034 ) | ( n1939 ) | ( n1660 ) ;
 assign n82 = ( (~ n500)  &  (~ n1329) ) ;
 assign n83 = ( (~ n1329)  &  n1657 ) ;
 assign n84 = ( (~ n1329)  &  (~ n1946) ) ;
 assign n85 = ( (~ n36) ) | ( n1045 ) | ( n1648 ) | ( n1661 ) | ( n1848 ) | ( n1940 ) | ( n1947 ) | ( n1948 ) ;
 assign n86 = ( n1038 ) | ( n1039 ) | ( n1040 ) | ( n1041 ) | ( n1042 ) | ( n1043 ) | ( (~ n2456) ) ;
 assign n87 = ( (~ n499)  &  n1657 ) ;
 assign n88 = ( (~ n499)  &  (~ n500) ) | ( (~ n499)  &  (~ n1946) ) ;
 assign n89 = ( n108  &  (~ n1635)  &  (~ n2458) ) ;
 assign n90 = ( n108  &  (~ n1635) ) | ( n161  &  (~ n1635) ) ;
 assign n91 = ( (~ i_6_)  &  i_7_ ) ;
 assign n95 = ( n503  &  n1032 ) | ( n503  &  n1033 ) ;
 assign n97 = ( n802  &  n265 ) | ( n802  &  n500 ) ;
 assign n98 = ( n509  &  n500 ) | ( n509  &  n507  &  n508 ) ;
 assign n99 = ( (~ n1645)  &  (~ n1659) ) ;
 assign n101 = ( n37  &  (~ n1017) ) ;
 assign n93 = ( n95  &  n97  &  n98  &  n99  &  n101  &  (~ n105)  &  (~ n1050)  &  (~ n1847) ) ;
 assign n102 = ( n505  &  (~ n1051)  &  n1056 ) | ( n505  &  n1056  &  n1054 ) ;
 assign n103 = ( n552  &  n553  &  (~ n670) ) ;
 assign n104 = ( n553  &  (~ n670)  &  (~ n1228) ) ;
 assign n105 = ( n1939 ) | ( n1026 ) | ( n1940 ) | ( n1941 ) | ( n1018 ) | ( n1040 ) ;
 assign n106 = ( (~ n1058)  &  n1844 ) ;
 assign n108 = ( i_3_  &  i_4_  &  (~ i_5_) ) ;
 assign n110 = ( n916  &  n1072  &  n1073  &  n1074  &  n1075  &  n1076  &  n1077  &  n1078 ) ;
 assign n112 = ( n701 ) | ( n1470 ) ;
 assign n113 = ( n537 ) | ( n701 ) ;
 assign n114 = ( (~ n35) ) | ( n701 ) ;
 assign n115 = ( n1377 ) | ( n701 ) ;
 assign n116 = ( n701 ) | ( n1425 ) ;
 assign n117 = ( n701 ) | ( n524 ) ;
 assign n118 = ( n701 ) | ( n1456 ) ;
 assign n119 = ( n1748  &  n952  &  n1762  &  n1421  &  n2004  &  n700 ) ;
 assign n111 = ( n112  &  n113  &  n114  &  n115  &  n116  &  n117  &  n118  &  n119 ) ;
 assign n121 = ( n1253  &  n1254  &  n1255 ) ;
 assign n122 = ( n1595  &  n450  &  n1596  &  n1597 ) ;
 assign n123 = ( n602  &  n603  &  n604  &  n605 ) ;
 assign n124 = ( n1898  &  n609  &  n589 ) ;
 assign n120 = ( n121  &  n122  &  n123  &  n124  &  n73 ) ;
 assign n125 = ( n136  &  n800  &  (~ n1847) ) | ( n136  &  n801  &  (~ n1847) ) ;
 assign n126 = ( n403  &  n242  &  n1161  &  n1162  &  n1163  &  n1164  &  n1165  &  n1166 ) ;
 assign n127 = ( n357  &  n358  &  n359  &  n360  &  n361  &  n362  &  n363  &  n364 ) ;
 assign n129 = ( n503  &  n504  &  n505  &  n506  &  n498 ) ;
 assign n128 = ( n37  &  n98  &  n129 ) ;
 assign n130 = ( n99  &  (~ n1644)  &  (~ n1664) ) ;
 assign n134 = ( n98  &  n800 ) | ( n98  &  n801 ) ;
 assign n135 = ( n37  &  (~ n1847) ) ;
 assign n136 = ( n805  &  n802  &  n799  &  n1056 ) ;
 assign n133 = ( n134  &  n135  &  n129  &  n136 ) ;
 assign n139 = ( (~ n59)  &  (~ n1639) ) | ( n1058  &  (~ n1639) ) | ( n1167  &  (~ n1639) ) ;
 assign n143 = ( n1208  &  n1210 ) ;
 assign n140 = ( n143  &  (~ n1229) ) | ( n143  &  (~ n1248) ) ;
 assign n144 = ( (~ n313)  &  (~ n748) ) | ( (~ n313)  &  (~ n1770) ) ;
 assign n147 = ( (~ n441)  &  (~ n1323) ) | ( (~ n441)  &  (~ n1339) ) ;
 assign n151 = ( n1184  &  n58 ) ;
 assign n150 = ( n151  &  (~ n1376) ) | ( (~ n780)  &  (~ n1376) ) ;
 assign n156 = ( (~ n812) ) | ( (~ n1063) ) ;
 assign n154 = ( n156  &  (~ n164) ) | ( (~ n164)  &  (~ n572) ) ;
 assign n160 = ( n1210  &  n58 ) ;
 assign n157 = ( n160  &  (~ n812) ) | ( n160  &  (~ n1239) ) ;
 assign n161 = ( i_5_  &  i_4_  &  i_3_ ) ;
 assign n166 = ( n164 ) | ( n1220 ) ;
 assign n167 = ( n164 ) | ( n1219 ) ;
 assign n164 = ( (~ n552) ) | ( (~ n1200) ) ;
 assign n165 = ( n1194 ) | ( n1195 ) ;
 assign n163 = ( n166  &  n167  &  n164 ) | ( n166  &  n167  &  n165 ) ;
 assign n169 = ( n1313  &  n1319 ) ;
 assign n170 = ( n1229  &  n178 ) ;
 assign n171 = ( n315  &  n340 ) ;
 assign n172 = ( n1190 ) | ( n1203 ) ;
 assign n173 = ( n1203 ) | ( n1218 ) ;
 assign n174 = ( n864  &  n176 ) ;
 assign n168 = ( n169  &  n170  &  n171  &  n172  &  n173  &  n174 ) ;
 assign n176 = ( n1218 ) | ( n1282 ) ;
 assign n177 = ( n1218 ) | ( n1278 ) ;
 assign n178 = ( n1194 ) | ( n1218 ) ;
 assign n179 = ( n1212 ) | ( n1234 ) ;
 assign n175 = ( n176  &  n173  &  n177  &  n178  &  n179 ) ;
 assign n182 = ( n1898  &  n2196  &  n2195 ) | ( n1898  &  n2196  &  n215 ) ;
 assign n180 = ( (~ i_9_) ) | ( (~ i_10_) ) | ( i_11_ ) ;
 assign n181 = ( n1057 ) | ( (~ n1250) ) ;
 assign n184 = ( n1167 ) | ( (~ n1184) ) ;
 assign n185 = ( n1190 ) | ( n1213 ) ;
 assign n187 = ( n1213 ) | ( n1218 ) ;
 assign n183 = ( (~ n143)  &  n184 ) | ( (~ n143)  &  n185 ) | ( n184  &  n187 ) | ( n185  &  n187 ) ;
 assign n192 = ( n388  &  n427 ) ;
 assign n188 = ( n192  &  (~ n198)  &  (~ n347)  &  (~ n848) ) ;
 assign n193 = ( (~ n751)  &  (~ n1268) ) | ( (~ n1063)  &  (~ n1268) ) ;
 assign n198 = ( (~ n313) ) | ( (~ n827) ) ;
 assign n197 = ( n198  &  (~ n1064) ) | ( (~ n462)  &  (~ n1064) ) | ( (~ n1064)  &  (~ n1281) ) ;
 assign n203 = ( (~ n193)  &  n1279 ) | ( (~ n193)  &  n811  &  n1241 ) ;
 assign n204 = ( (~ n154)  &  (~ n237) ) | ( (~ n154)  &  n1220  &  n1262 ) ;
 assign n205 = ( n177  &  (~ n197)  &  n2209 ) | ( (~ n197)  &  n2178  &  n2209 ) ;
 assign n206 = ( n1925  &  n967  &  n933  &  n445  &  n592  &  n1668  &  n643  &  n640 ) ;
 assign n207 = ( n663  &  n183  &  n2216  &  n2217  &  n2214  &  n2213  &  n2212  &  n2211 ) ;
 assign n208 = ( n429  &  n382  &  n822  &  n877  &  n893  &  n1869  &  n442  &  n636 ) ;
 assign n209 = ( n647  &  n436  &  n632  &  n2207  &  n371  &  n367  &  n1833  &  n1832 ) ;
 assign n210 = ( n1778  &  n386  &  n379  &  n376  &  n1760  &  n742  &  n2202  &  n2204 ) ;
 assign n202 = ( n203  &  n204  &  n205  &  n206  &  n207  &  n208  &  n209  &  n210 ) ;
 assign n212 = ( n1231 ) | ( (~ n1250) ) ;
 assign n211 = ( (~ n57) ) | ( n212 ) ;
 assign n216 = ( n452 ) | ( n212 ) ;
 assign n217 = ( n1243 ) | ( n212 ) ;
 assign n215 = ( i_9_ ) | ( (~ i_10_) ) | ( i_11_ ) ;
 assign n214 = ( n216  &  n217  &  n215 ) | ( n216  &  n217  &  n212 ) ;
 assign n221 = ( n164 ) | ( n1332 ) ;
 assign n219 = ( n1339  &  n1340  &  n1341 ) ;
 assign n220 = ( n1238 ) | ( n1311 ) ;
 assign n218 = ( n221  &  n164 ) | ( n221  &  n219  &  n220 ) ;
 assign n223 = ( n531 ) | ( (~ n827) ) ;
 assign n222 = ( n223  &  (~ n1325) ) | ( (~ n462)  &  (~ n1325) ) ;
 assign n229 = ( n160 ) | ( (~ n427) ) ;
 assign n225 = ( n229  &  (~ n864) ) | ( n229  &  (~ n1319) ) | ( n229  &  (~ n1347) ) ;
 assign n233 = ( (~ n343) ) | ( (~ n1423) ) ;
 assign n230 = ( (~ n219)  &  (~ n1268) ) | ( n233  &  (~ n1268) ) | ( (~ n1268)  &  (~ n1326) ) ;
 assign n237 = ( (~ n184) ) | ( (~ n374) ) ;
 assign n236 = ( (~ n165) ) | ( (~ n1469) ) ;
 assign n234 = ( n237  &  n236 ) | ( n237  &  (~ n1317) ) | ( n237  &  (~ n1343) ) ;
 assign n239 = ( (~ n184) ) | ( n855 ) ;
 assign n240 = ( (~ n313) ) | ( (~ n427) ) | ( (~ n462) ) ;
 assign n238 = ( n223  &  (~ n1315) ) | ( n239  &  (~ n1315) ) | ( n240  &  (~ n1315) ) ;
 assign n243 = ( (~ n225)  &  n1312 ) | ( (~ n225)  &  n441  &  n1271 ) ;
 assign n244 = ( (~ n222)  &  n2173 ) | ( (~ n222)  &  n646  &  n1322 ) ;
 assign n245 = ( (~ n230)  &  n1333  &  n2176 ) | ( (~ n230)  &  n2176  &  n2179 ) ;
 assign n246 = ( n1921  &  n2172  &  n960  &  n966  &  n1172  &  n932  &  n591  &  n642 ) ;
 assign n247 = ( (~ n234)  &  (~ n238)  &  n2181  &  n2183  &  n2184  &  n2185 ) ;
 assign n248 = ( n432  &  n639  &  n428  &  n425  &  n383  &  n821  &  n876  &  n892 ) ;
 assign n249 = ( n1870  &  n635  &  n435  &  n631  &  n372  &  n368  &  n1830  &  n2171 ) ;
 assign n250 = ( n378  &  n375  &  n1761  &  n1718  &  n1723  &  n2170  &  n2166  &  n2167 ) ;
 assign n242 = ( n243  &  n244  &  n245  &  n246  &  n247  &  n248  &  n249  &  n250 ) ;
 assign n251 = ( n177 ) | ( (~ n392) ) ;
 assign n254 = ( n427 ) | ( n1267 ) ;
 assign n255 = ( n173 ) | ( (~ n855) ) ;
 assign n256 = ( n427 ) | ( n517 ) ;
 assign n257 = ( n427 ) | ( n1263 ) ;
 assign n258 = ( n177 ) | ( (~ n975) ) ;
 assign n259 = ( n1752  &  n594  &  n1873  &  n580  &  n1698  &  n1711 ) ;
 assign n260 = ( (~ n150)  &  n660  &  n1378  &  n1390  &  n1766  &  n1831  &  n2157  &  n2159 ) ;
 assign n261 = ( n741  &  n2153  &  n1836  &  n1862  &  n1849  &  n2150  &  n2146  &  n2145 ) ;
 assign n253 = ( n254  &  n255  &  n256  &  n257  &  n258  &  n259  &  n260  &  n261 ) ;
 assign n263 = ( n374  &  n388 ) ;
 assign n262 = ( n179 ) | ( n263 ) ;
 assign n265 = ( n1191 ) | ( n1223 ) ;
 assign n266 = ( n1191 ) | ( n1240 ) ;
 assign n264 = ( n265  &  n266 ) ;
 assign n268 = ( n1419  &  n1420  &  n113  &  n1421  &  n262  &  n1422 ) ;
 assign n269 = ( n1413  &  n1414  &  n1415  &  n1416  &  n1417  &  n1418 ) ;
 assign n270 = ( n1405  &  n1406  &  n1407  &  n1408  &  n1409  &  n1410  &  n1411  &  n1412 ) ;
 assign n271 = ( n1398  &  n1399  &  n1400  &  n1401  &  n1402  &  n1403  &  n1404 ) ;
 assign n272 = ( (~ n151)  &  n2136  &  n2137 ) | ( n179  &  n2136  &  n2137 ) ;
 assign n273 = ( n1927  &  n1901  &  n1691  &  n1767  &  n1828  &  n1903  &  n1856  &  n2135 ) ;
 assign n274 = ( n598  &  n1715  &  n1753  &  n1905  &  n846  &  n2134 ) ;
 assign n275 = ( n1819  &  n1728  &  n2132  &  n2133  &  n1796  &  n2130 ) ;
 assign n267 = ( n268  &  n269  &  n270  &  n271  &  n272  &  n273  &  n274  &  n275 ) ;
 assign n277 = ( n1195 ) | ( n1282 ) ;
 assign n276 = ( (~ n160) ) | ( n277 ) ;
 assign n280 = ( n427 ) | ( n277 ) ;
 assign n281 = ( (~ n855) ) | ( n864 ) ;
 assign n282 = ( n427 ) | ( n458 ) ;
 assign n283 = ( n427 ) | ( n1344 ) ;
 assign n284 = ( (~ n975) ) | ( n1342 ) ;
 assign n285 = ( n1697  &  n1861  &  n583  &  n597  &  n1716 ) ;
 assign n286 = ( n1920  &  n2118  &  n1859  &  n2116  &  n1447  &  n1439  &  n2117  &  n1432 ) ;
 assign n287 = ( n2114  &  n2115  &  n1850  &  n816  &  n817  &  n2113  &  n2109 ) ;
 assign n279 = ( n280  &  n281  &  n282  &  n283  &  n284  &  n285  &  n286  &  n287 ) ;
 assign n289 = ( n1463  &  n1464  &  n1465  &  n1466  &  n1467  &  n1468 ) ;
 assign n290 = ( n1457  &  n1458  &  n1459  &  n1460  &  n1461  &  n1462 ) ;
 assign n291 = ( (~ n855)  &  n2097 ) | ( n1033  &  n2097 ) ;
 assign n292 = ( (~ n151)  &  n388 ) | ( (~ n151)  &  n749 ) | ( n388  &  n1347 ) | ( n749  &  n1347 ) ;
 assign n293 = ( n2095  &  n184 ) | ( n2095  &  n1127 ) ;
 assign n294 = ( n1829  &  n2094  &  n1764  &  n1857  &  n1768  &  n2093 ) ;
 assign n295 = ( n1754  &  n1750  &  n845  &  n1675  &  n1906  &  n599  &  n585  &  n2091 ) ;
 assign n296 = ( n712  &  n1795  &  n1802  &  n1812  &  n1792  &  n2089 ) ;
 assign n288 = ( n289  &  n290  &  n291  &  n292  &  n293  &  n294  &  n295  &  n296 ) ;
 assign n298 = ( n184 ) | ( n1328 ) ;
 assign n299 = ( n184 ) | ( n1206 ) ;
 assign n300 = ( n1219 ) | ( n374 ) ;
 assign n301 = ( n184 ) | ( n1340 ) ;
 assign n302 = ( n184 ) | ( n1247 ) ;
 assign n303 = ( n1823  &  n1822  &  n1744  &  n1726  &  n1727  &  n740 ) ;
 assign n304 = ( n1699  &  n1811  &  n1700  &  n582  &  n1706  &  n2077  &  n1789  &  n2075 ) ;
 assign n305 = ( n2084  &  n1693  &  n1763  &  n2081  &  n1476  &  n1471  &  n2083  &  n2079 ) ;
 assign n297 = ( n298  &  n299  &  n300  &  n301  &  n302  &  n303  &  n304  &  n305 ) ;
 assign n307 = ( n1190 ) | ( n1211 ) ;
 assign n308 = ( n1211 ) | ( n1218 ) ;
 assign n306 = ( n307  &  n308  &  (~ n935) ) ;
 assign n312 = ( n1329  &  n811 ) ;
 assign n313 = ( (~ n552) ) | ( (~ n1184) ) ;
 assign n310 = ( n306  &  n312 ) | ( n306  &  n313 ) | ( n312  &  (~ n401) ) | ( n313  &  (~ n401) ) ;
 assign n317 = ( n313 ) | ( n1239 ) ;
 assign n315 = ( n1323  &  n1239 ) ;
 assign n316 = ( n646  &  n1241 ) ;
 assign n314 = ( n317  &  (~ n401) ) | ( n317  &  n315  &  n316 ) ;
 assign n319 = ( (~ n922)  &  n1248 ) ;
 assign n318 = ( n319 ) | ( (~ n392) ) ;
 assign n321 = ( n164 ) | ( n1455 ) ;
 assign n322 = ( n374 ) | ( n1456 ) ;
 assign n323 = ( n313 ) | ( n1455 ) ;
 assign n324 = ( n313 ) | ( n749 ) ;
 assign n325 = ( n164 ) | ( n1347 ) ;
 assign n326 = ( n441 ) | ( n1455 ) ;
 assign n327 = ( n1277 ) | ( n1456 ) ;
 assign n328 = ( n118  &  n1840  &  n2005  &  n2006  &  n2003  &  n2007 ) ;
 assign n320 = ( n321  &  n322  &  n323  &  n324  &  n325  &  n326  &  n327  &  n328 ) ;
 assign n330 = ( n164  &  (~ n356) ) | ( n164  &  n388 ) | ( (~ n356)  &  n1071 ) | ( n388  &  n1071 ) ;
 assign n329 = ( n330  &  n320 ) ;
 assign n333 = ( (~ n1057)  &  n1210 ) ;
 assign n331 = ( n333  &  (~ n1347) ) | ( n333  &  (~ n1456) ) ;
 assign n337 = ( (~ n14) ) | ( n811 ) ;
 assign n338 = ( n2518 ) | ( n164 ) ;
 assign n335 = ( (~ n922)  &  n1330 ) ;
 assign n334 = ( (~ n14)  &  n337  &  n338 ) | ( n337  &  n338  &  n335 ) ;
 assign n340 = ( n307  &  n308 ) ;
 assign n341 = ( (~ n356)  &  n1396  &  n1511 ) ;
 assign n339 = ( n340  &  n172  &  n341 ) ;
 assign n343 = ( n499  &  n1330 ) ;
 assign n342 = ( n343  &  (~ n935) ) ;
 assign n347 = ( (~ n184) ) | ( n333 ) ;
 assign n344 = ( (~ n174)  &  n347 ) | ( (~ n340)  &  n347 ) ;
 assign n350 = ( n143 ) | ( n14 ) ;
 assign n349 = ( (~ n308) ) | ( (~ n1397) ) ;
 assign n348 = ( n350  &  n349 ) | ( n350  &  n13 ) ;
 assign n351 = ( n237  &  (~ n1066) ) | ( n237  &  (~ n1245) ) ;
 assign n356 = ( (~ n1376) ) | ( (~ n1424) ) ;
 assign n354 = ( n333  &  n356 ) | ( n333  &  (~ n651) ) ;
 assign n357 = ( n184  &  (~ n198) ) | ( n184  &  (~ n233) ) | ( (~ n198)  &  n1738 ) | ( (~ n233)  &  n1738 ) ;
 assign n358 = ( n263  &  (~ n356) ) | ( (~ n356)  &  n657 ) | ( n263  &  n701 ) | ( n657  &  n701 ) ;
 assign n359 = ( n315  &  n319 ) | ( n374  &  n319 ) | ( n315  &  n827 ) | ( n374  &  n827 ) ;
 assign n360 = ( n1265  &  n1937 ) | ( n762  &  n1937 ) | ( n1265  &  n1277 ) | ( n762  &  n1277 ) ;
 assign n361 = ( n390  &  n329  &  n1170  &  n334  &  n2245  &  n2244 ) ;
 assign n362 = ( n253  &  n267  &  n279  &  n288  &  n202  &  n242  &  n163  &  n2246 ) ;
 assign n363 = ( n2241  &  n2243  &  n2238  &  n2236  &  n2234  &  n2232  &  n2231  &  n2230 ) ;
 assign n364 = ( (~ n140)  &  n2218  &  n2219  &  n2221  &  n2223  &  n2225  &  n2227  &  n2229 ) ;
 assign n367 = ( n164 ) | ( n1235 ) ;
 assign n368 = ( n164 ) | ( n172 ) ;
 assign n366 = ( n1191 ) | ( n1203 ) ;
 assign n365 = ( n367  &  n368  &  n164 ) | ( n367  &  n368  &  n366 ) ;
 assign n371 = ( n164 ) | ( n1236 ) ;
 assign n372 = ( n164 ) | ( n1319 ) ;
 assign n370 = ( n1191 ) | ( n1194 ) ;
 assign n369 = ( n371  &  n372  &  n164 ) | ( n371  &  n372  &  n370 ) ;
 assign n375 = ( n374 ) | ( n172 ) ;
 assign n376 = ( n374 ) | ( n173 ) ;
 assign n374 = ( (~ n1184) ) | ( n1228 ) ;
 assign n373 = ( n375  &  n376  &  n374 ) | ( n375  &  n376  &  n366 ) ;
 assign n378 = ( n374 ) | ( n1319 ) ;
 assign n379 = ( n374 ) | ( n178 ) ;
 assign n377 = ( n378  &  n379  &  n374 ) | ( n378  &  n379  &  n370 ) ;
 assign n382 = ( n164 ) | ( n1248 ) ;
 assign n383 = ( n164 ) | ( n1313 ) ;
 assign n381 = ( n1191 ) | ( n1215 ) ;
 assign n380 = ( n382  &  n383  &  n164 ) | ( n382  &  n383  &  n381 ) ;
 assign n385 = ( n374 ) | ( n1313 ) ;
 assign n386 = ( n374 ) | ( n1229 ) ;
 assign n384 = ( n385  &  n386  &  n374 ) | ( n385  &  n386  &  n381 ) ;
 assign n389 = ( n313 ) | ( n1376 ) ;
 assign n390 = ( n1522  &  n1523  &  n1095  &  n1524  &  n115  &  n1525 ) ;
 assign n388 = ( (~ n1200) ) | ( n1228 ) ;
 assign n387 = ( n389  &  n390  &  n388 ) | ( n389  &  n390  &  n176 ) ;
 assign n392 = ( (~ n313) ) | ( n401 ) ;
 assign n391 = ( n392  &  (~ n1248) ) | ( (~ n827)  &  (~ n1248) ) ;
 assign n394 = ( n1546  &  n1547  &  n1548  &  n1549  &  n1550  &  n1551  &  n1552  &  n1553 ) ;
 assign n395 = ( (~ n531)  &  n1485  &  n2269 ) | ( n1236  &  n1485  &  n2269 ) ;
 assign n396 = ( n184  &  (~ n848) ) | ( n184  &  n1263 ) | ( (~ n848)  &  n1267 ) | ( n1263  &  n1267 ) ;
 assign n397 = ( n2266  &  n1581 ) | ( n1376  &  n1581 ) | ( n2266  &  n308 ) | ( n1376  &  n308 ) ;
 assign n398 = ( n176  &  n2268 ) | ( (~ n531)  &  n1581  &  n2268 ) ;
 assign n399 = ( (~ n391)  &  n1239 ) | ( (~ n392)  &  (~ n391)  &  n1579 ) ;
 assign n393 = ( n253  &  n394  &  n387  &  n395  &  n396  &  n397  &  n398  &  n399 ) ;
 assign n401 = ( n1184  &  n1208 ) ;
 assign n400 = ( n401  &  (~ n1323) ) | ( (~ n1323)  &  (~ n1579) ) ;
 assign n404 = ( n441 ) | ( n1423 ) ;
 assign n405 = ( n441 ) | ( n1334 ) ;
 assign n406 = ( (~ n400)  &  n864 ) | ( (~ n400)  &  n1581  &  n1582 ) ;
 assign n407 = ( n172  &  (~ n541) ) | ( n172  &  n1425 ) | ( (~ n541)  &  n2265 ) | ( n1425  &  n2265 ) ;
 assign n408 = ( n1641 ) | ( n1423 ) ;
 assign n409 = ( n1581  &  n1583 ) | ( n307  &  n1583 ) | ( n1581  &  n1334 ) | ( n307  &  n1334 ) ;
 assign n410 = ( n2266  &  n2242 ) | ( n1424  &  n2242 ) | ( n2266  &  n1344 ) | ( n1424  &  n1344 ) ;
 assign n411 = ( (~ n143)  &  n279  &  n1169 ) | ( n279  &  n1169  &  n1339 ) ;
 assign n403 = ( n404  &  n405  &  n406  &  n407  &  n408  &  n409  &  n410  &  n411 ) ;
 assign n412 = ( n333  &  (~ n638) ) | ( n333  &  (~ n1587) ) ;
 assign n415 = ( n441 ) | ( n634 ) ;
 assign n416 = ( n441 ) | ( n1585 ) ;
 assign n417 = ( n441 ) | ( n630 ) ;
 assign n418 = ( (~ n14) ) | ( n634 ) ;
 assign n419 = ( (~ n143)  &  n2260 ) | ( n434  &  n634  &  n2260 ) ;
 assign n420 = ( (~ n350)  &  n701 ) | ( n645  &  n701 ) | ( (~ n350)  &  n1587 ) | ( n645  &  n1587 ) ;
 assign n421 = ( (~ n412)  &  n1589  &  n1590  &  n1591  &  n1592  &  n1594 ) ;
 assign n422 = ( (~ n692)  &  n2262 ) | ( n1602  &  n2262 ) ;
 assign n414 = ( n415  &  n416  &  n417  &  n418  &  n419  &  n420  &  n421  &  n422 ) ;
 assign n425 = ( (~ n160) ) | ( n172 ) ;
 assign n424 = ( n366  &  n173 ) ;
 assign n423 = ( (~ n160)  &  n425 ) | ( n425  &  n424 ) ;
 assign n428 = ( n427 ) | ( n1313 ) ;
 assign n429 = ( n1229 ) | ( n427 ) ;
 assign n427 = ( (~ n1210) ) | ( n1231 ) ;
 assign n426 = ( n428  &  n429  &  n427 ) | ( n428  &  n429  &  n381 ) ;
 assign n432 = ( (~ n160) ) | ( n1313 ) ;
 assign n431 = ( n381  &  n1229 ) ;
 assign n430 = ( (~ n160)  &  n432 ) | ( n432  &  n431 ) ;
 assign n435 = ( n427 ) | ( n1323 ) ;
 assign n436 = ( n427 ) | ( n1239 ) ;
 assign n434 = ( n1191 ) | ( n1238 ) ;
 assign n433 = ( n435  &  n436  &  n427 ) | ( n435  &  n436  &  n434 ) ;
 assign n439 = ( (~ n174) ) | ( (~ n456) ) ;
 assign n437 = ( n160  &  n439 ) | ( n160  &  (~ n460) ) ;
 assign n442 = ( n441 ) | ( n1235 ) ;
 assign n443 = ( n441 ) | ( n172 ) ;
 assign n441 = ( (~ n1210) ) | ( n1224 ) ;
 assign n440 = ( n442  &  n443  &  n441 ) | ( n442  &  n443  &  n366 ) ;
 assign n445 = ( n441 ) | ( n1248 ) ;
 assign n446 = ( n441 ) | ( n1313 ) ;
 assign n444 = ( n445  &  n446  &  n441 ) | ( n445  &  n446  &  n381 ) ;
 assign n448 = ( (~ n1140)  &  n2251 ) | ( n998  &  n1130  &  n2251 ) ;
 assign n449 = ( (~ n333) ) | ( n748 ) ;
 assign n447 = ( n440  &  n444  &  n448  &  n449 ) ;
 assign n451 = ( (~ n1208) ) | ( (~ n1250) ) ;
 assign n452 = ( i_9_ ) | ( i_10_ ) | ( (~ i_11_) ) ;
 assign n450 = ( n451 ) | ( n452 ) ;
 assign n454 = ( n2250  &  n2195 ) | ( n2250  &  n452 ) ;
 assign n453 = ( (~ i_9_) ) | ( i_10_ ) | ( (~ i_11_) ) ;
 assign n456 = ( n1191 ) | ( n1282 ) ;
 assign n455 = ( n456 ) | ( n313 ) ;
 assign n458 = ( n1195 ) | ( n1211 ) ;
 assign n459 = ( n1585  &  n1587  &  n590  &  n1601  &  n1602 ) ;
 assign n460 = ( n1217 ) | ( n1282 ) ;
 assign n457 = ( n165  &  n277  &  n458  &  n459  &  n460 ) ;
 assign n462 = ( n164  &  n263 ) ;
 assign n464 = ( (~ n392)  &  (~ n855) ) ;
 assign n461 = ( n462  &  n464  &  (~ n1138) ) ;
 assign n466 = ( n1194 ) | ( n1217 ) ;
 assign n465 = ( n466  &  n460  &  n370  &  n456 ) ;
 assign n468 = ( (~ n143) ) | ( n2513 ) ;
 assign n467 = ( (~ n143)  &  n468 ) | ( n466  &  n468 ) ;
 assign n470 = ( n1217 ) | ( n1238 ) ;
 assign n471 = ( n1217 ) | ( n1278 ) ;
 assign n472 = ( n1211 ) | ( n1217 ) ;
 assign n469 = ( n470  &  n471  &  n472 ) ;
 assign n473 = ( (~ n308)  &  n350 ) | ( n350  &  (~ n470) ) ;
 assign n476 = ( (~ n366)  &  (~ n827) ) | ( (~ n517)  &  (~ n827) ) ;
 assign n482 = ( (~ n388) ) | ( (~ n891) ) ;
 assign n479 = ( n482  &  (~ n1235) ) | ( n482  &  (~ n1248) ) | ( n482  &  (~ n1578) ) ;
 assign n486 = ( n482 ) | ( (~ n1268) ) ;
 assign n483 = ( n486  &  (~ n517) ) | ( n486  &  (~ n1334) ) | ( n486  &  (~ n1423) ) ;
 assign n487 = ( (~ n434)  &  (~ n462) ) | ( (~ n456)  &  (~ n462) ) | ( (~ n462)  &  (~ n812) ) ;
 assign n490 = ( (~ n237)  &  n366 ) | ( n366  &  n1578 ) | ( (~ n237)  &  n1580 ) | ( n1578  &  n1580 ) ;
 assign n491 = ( n1271  &  n1269 ) | ( n457  &  n1269 ) | ( n1271  &  n456 ) | ( n457  &  n456 ) ;
 assign n492 = ( n1604  &  n1967 ) | ( n471  &  n1967 ) | ( n1604  &  n517 ) | ( n471  &  n517 ) ;
 assign n493 = ( n2283  &  n2177 ) | ( n1600  &  n2177 ) | ( n2283  &  n748 ) | ( n1600  &  n748 ) ;
 assign n494 = ( (~ n479)  &  (~ n483)  &  (~ n487)  &  n2275  &  n2277  &  n2279 ) ;
 assign n495 = ( n1692  &  n1670  &  n941  &  n1852  &  n2273  &  n2271 ) ;
 assign n496 = ( n888  &  n1851  &  n1785  &  n1765  &  n1759  &  n1751  &  n2270  &  n1719 ) ;
 assign n497 = ( n2294  &  n2293  &  n2296  &  n2291  &  n2289  &  n2288  &  n2298  &  n2297 ) ;
 assign n489 = ( n490  &  n491  &  n492  &  n493  &  n494  &  n495  &  n496  &  n497 ) ;
 assign n499 = ( n1215 ) | ( n1316 ) ;
 assign n500 = ( (~ n1208) ) | ( n1636 ) ;
 assign n498 = ( (~ n77)  &  (~ n82)  &  n499 ) | ( (~ n77)  &  (~ n82)  &  n500 ) ;
 assign n503 = ( n1033 ) | ( n500 ) ;
 assign n504 = ( n1638 ) | ( n1058 ) ;
 assign n505 = ( n1638 ) | ( n670 ) ;
 assign n506 = ( n1638  &  n265 ) | ( n807  &  n265 ) | ( n1638  &  n500 ) | ( n807  &  n500 ) ;
 assign n509 = ( (~ n1230) ) | ( n1636 ) ;
 assign n507 = ( n657  &  n1346 ) ;
 assign n508 = ( n1127  &  n1066 ) ;
 assign n511 = ( n1191 ) | ( n1216 ) ;
 assign n510 = ( (~ n14)  &  n337 ) | ( n337  &  n511 ) ;
 assign n514 = ( (~ n14) ) | ( n1330 ) ;
 assign n513 = ( (~ n349)  &  n1509 ) ;
 assign n512 = ( (~ n143)  &  n510  &  n514 ) | ( n510  &  n514  &  n513 ) ;
 assign n517 = ( n1213 ) | ( n1217 ) ;
 assign n515 = ( (~ n14)  &  (~ n27) ) | ( (~ n27)  &  (~ n349)  &  n517 ) ;
 assign n520 = ( n1190 ) | ( n1216 ) ;
 assign n519 = ( (~ n143)  &  (~ n140)  &  n515 ) | ( (~ n140)  &  n515  &  n520 ) ;
 assign n525 = ( n1563  &  n1564  &  n1565  &  n1566  &  n1567  &  n1568  &  n1569  &  n1570 ) ;
 assign n524 = ( n1212 ) | ( n1321 ) ;
 assign n522 = ( (~ n333)  &  n525 ) | ( n525  &  n524 ) ;
 assign n526 = ( (~ n164)  &  (~ n1318) ) | ( n401  &  (~ n1318) ) ;
 assign n527 = ( n14  &  (~ n520) ) | ( (~ n520)  &  (~ n1641) ) ;
 assign n531 = ( (~ n1057)  &  n1200 ) ;
 assign n530 = ( n392  &  (~ n1219) ) | ( n531  &  (~ n1219) ) ;
 assign n533 = ( (~ n164)  &  (~ n1470) ) | ( (~ n1277)  &  (~ n1470) ) ;
 assign n538 = ( n1571  &  n1572  &  n1573  &  n832  &  n1574  &  n1575  &  n1576  &  n1577 ) ;
 assign n537 = ( n1191 ) | ( n1234 ) ;
 assign n536 = ( (~ n333)  &  n538 ) | ( n538  &  n537 ) ;
 assign n539 = ( (~ n160)  &  n263 ) ;
 assign n541 = ( (~ n164) ) | ( n229 ) ;
 assign n540 = ( (~ n537)  &  n541 ) | ( (~ n537)  &  (~ n1277) ) ;
 assign n544 = ( n313  &  (~ n401) ) | ( (~ n401)  &  n811 ) | ( n313  &  n1241 ) | ( n811  &  n1241 ) ;
 assign n545 = ( (~ n160)  &  n374 ) | ( (~ n160)  &  n1066 ) | ( n374  &  n1233 ) | ( n1066  &  n1233 ) ;
 assign n546 = ( n265  &  (~ n392) ) | ( (~ n392)  &  (~ n848) ) | ( n265  &  n1220 ) | ( (~ n848)  &  n1220 ) ;
 assign n547 = ( n539  &  n1583 ) | ( n1245  &  n1583 ) | ( n539  &  n1128 ) | ( n1245  &  n1128 ) ;
 assign n548 = ( n511  &  (~ n540) ) | ( (~ n143)  &  (~ n540)  &  n1641 ) ;
 assign n549 = ( n1506  &  n166  &  n2299 ) ;
 assign n543 = ( n536  &  n267  &  n544  &  n545  &  n546  &  n547  &  n548  &  n549 ) ;
 assign n552 = ( i_8_  &  (~ n1178) ) ;
 assign n553 = ( n1198  &  (~ n1635) ) ;
 assign n550 = ( n552  &  n553  &  (~ n807) ) ;
 assign n555 = ( n1208  &  n553 ) ;
 assign n554 = ( n555  &  (~ n673) ) ;
 assign n559 = ( n202  &  n393  &  n827 ) | ( n202  &  n393  &  n176 ) ;
 assign n560 = ( n512  &  n519  &  n1650  &  n543 ) ;
 assign n561 = ( (~ n401)  &  (~ n531) ) | ( n517  &  (~ n531) ) | ( (~ n401)  &  n1220 ) | ( n517  &  n1220 ) ;
 assign n562 = ( (~ n14)  &  n1340 ) | ( n812  &  n1340 ) | ( (~ n14)  &  n2292 ) | ( n812  &  n2292 ) ;
 assign n563 = ( n2318  &  n2320  &  n2173 ) | ( n2318  &  n2320  &  n1233 ) ;
 assign n564 = ( n2307  &  n2317  &  n2309  &  n2306  &  n2305  &  n2316  &  n2315  &  n2313 ) ;
 assign n557 = ( n559  &  n560  &  n561  &  n562  &  n563  &  n564  &  (~ n1644)  &  (~ n1645) ) ;
 assign n565 = ( n553  &  (~ n807)  &  (~ n1228) ) ;
 assign n570 = ( n1167 ) | ( (~ n1733) ) ;
 assign n567 = ( n570  &  (~ n1208) ) | ( n570  &  (~ n1733) ) ;
 assign n572 = ( n1218 ) | ( n1240 ) ;
 assign n571 = ( n470  &  n572 ) ;
 assign n574 = ( n1189 ) | ( n1316 ) ;
 assign n573 = ( (~ n333)  &  n441 ) | ( n441  &  n571 ) | ( (~ n333)  &  n574 ) | ( n571  &  n574 ) ;
 assign n577 = ( (~ n333) ) | ( n1267 ) ;
 assign n578 = ( n1706  &  n1707  &  n417  &  n1708  &  n1709 ) ;
 assign n575 = ( (~ n333)  &  n577  &  n578 ) | ( (~ n439)  &  n577  &  n578 ) ;
 assign n580 = ( n441 ) | ( n1267 ) ;
 assign n581 = ( n441 ) | ( n864 ) ;
 assign n582 = ( n441 ) | ( n1246 ) ;
 assign n583 = ( n441 ) | ( n277 ) ;
 assign n584 = ( n441 ) | ( n1245 ) ;
 assign n585 = ( n441 ) | ( n749 ) ;
 assign n586 = ( n441 ) | ( n750 ) ;
 assign n587 = ( n416  &  n441 ) | ( n416  &  n456 ) ;
 assign n579 = ( n580  &  n581  &  n582  &  n583  &  n584  &  n585  &  n586  &  n587 ) ;
 assign n588 = ( (~ n333) ) | ( n366 ) ;
 assign n591 = ( (~ n160) ) | ( n1315 ) ;
 assign n592 = ( (~ n160) ) | ( n1226 ) ;
 assign n590 = ( n1215 ) | ( n1217 ) ;
 assign n589 = ( (~ n160)  &  n591  &  n592 ) | ( n591  &  n592  &  n590 ) ;
 assign n594 = ( n441 ) | ( n1236 ) ;
 assign n595 = ( n441 ) | ( n1319 ) ;
 assign n596 = ( n1219 ) | ( n441 ) ;
 assign n597 = ( n165 ) | ( n441 ) ;
 assign n598 = ( n1220 ) | ( n441 ) ;
 assign n599 = ( n441 ) | ( n1454 ) ;
 assign n600 = ( n441 ) | ( n1469 ) ;
 assign n601 = ( n415  &  n441 ) | ( n415  &  n370 ) ;
 assign n593 = ( n594  &  n595  &  n596  &  n597  &  n598  &  n599  &  n600  &  n601 ) ;
 assign n602 = ( n427 ) | ( n187 ) ;
 assign n603 = ( n427 ) | ( n617 ) ;
 assign n604 = ( n427 ) | ( n1331 ) ;
 assign n605 = ( (~ n160)  &  (~ n229) ) | ( (~ n160)  &  n773 ) | ( (~ n229)  &  n1705 ) | ( n773  &  n1705 ) ;
 assign n609 = ( (~ n160) ) | ( n617 ) ;
 assign n608 = ( n1244 ) | ( n1316 ) ;
 assign n606 = ( n609  &  n608 ) | ( n609  &  (~ n1140) ) ;
 assign n611 = ( (~ n356)  &  n370  &  n381  &  n619 ) ;
 assign n612 = ( n460  &  n1704 ) ;
 assign n610 = ( n611  &  n340  &  n612 ) ;
 assign n614 = ( n1240 ) | ( n1316 ) ;
 assign n613 = ( n220  &  n614 ) ;
 assign n615 = ( (~ n333)  &  n441 ) | ( (~ n333)  &  n470 ) | ( n441  &  n613 ) | ( n470  &  n613 ) ;
 assign n617 = ( n1216 ) | ( n1316 ) ;
 assign n616 = ( n617 ) | ( n441 ) ;
 assign n619 = ( n1204 ) | ( n1316 ) ;
 assign n618 = ( (~ n160) ) | ( n619 ) ;
 assign n620 = ( (~ n160) ) | ( n608 ) ;
 assign n623 = ( n2511 ) | ( n427 ) ;
 assign n624 = ( n2084  &  n2118  &  n2094 ) ;
 assign n622 = ( n781  &  n1508 ) ;
 assign n621 = ( (~ n160)  &  n623  &  n624 ) | ( n623  &  n624  &  n622 ) ;
 assign n626 = ( n634  &  n1242  &  n1324 ) ;
 assign n625 = ( n427 ) | ( n626 ) ;
 assign n628 = ( n1586  &  n761 ) ;
 assign n627 = ( n427 ) | ( n628 ) ;
 assign n631 = ( (~ n160) ) | ( n1322 ) ;
 assign n632 = ( (~ n160) ) | ( n1237 ) ;
 assign n630 = ( n1195 ) | ( n1204 ) ;
 assign n629 = ( (~ n160)  &  n631  &  n632 ) | ( n631  &  n632  &  n630 ) ;
 assign n635 = ( (~ n160) ) | ( n1324 ) ;
 assign n636 = ( (~ n160) ) | ( n1242 ) ;
 assign n634 = ( n1189 ) | ( n1195 ) ;
 assign n633 = ( (~ n160)  &  n635  &  n636 ) | ( n635  &  n636  &  n634 ) ;
 assign n639 = ( n427 ) | ( n1329 ) ;
 assign n640 = ( n427 ) | ( n811 ) ;
 assign n638 = ( n1195 ) | ( n1216 ) ;
 assign n637 = ( n639  &  n640  &  n427 ) | ( n639  &  n640  &  n638 ) ;
 assign n642 = ( (~ n160) ) | ( n1329 ) ;
 assign n643 = ( (~ n160) ) | ( n811 ) ;
 assign n641 = ( (~ n160)  &  n642  &  n643 ) | ( n638  &  n642  &  n643 ) ;
 assign n647 = ( n427 ) | ( n1241 ) ;
 assign n645 = ( n1195 ) | ( n1240 ) ;
 assign n646 = ( n1240 ) | ( n1311 ) ;
 assign n644 = ( n647  &  n427 ) | ( n647  &  n645  &  n646 ) ;
 assign n649 = ( n1585  &  n1396  &  n1455 ) ;
 assign n648 = ( n427 ) | ( n649 ) ;
 assign n652 = ( n1672  &  n280  &  n254  &  n1673  &  n1674  &  n1675  &  n648 ) ;
 assign n651 = ( n537  &  n1425  &  n524 ) ;
 assign n650 = ( n652  &  n651 ) | ( n652  &  n427 ) ;
 assign n654 = ( n1678  &  n824  &  n1082  &  n1068  &  n1081 ) ;
 assign n656 = ( n466  &  n1676 ) ;
 assign n657 = ( n1213 ) | ( n1311 ) ;
 assign n658 = ( n1245  &  n1246 ) ;
 assign n653 = ( (~ n356)  &  n614  &  n654  &  n656  &  n657  &  n658 ) ;
 assign n660 = ( (~ n157)  &  n868  &  n1383  &  n1384  &  n1385  &  n1386  &  n1388  &  n1389 ) ;
 assign n661 = ( n1353  &  n1354  &  n1355  &  n1356  &  n1335 ) ;
 assign n662 = ( (~ n160)  &  n427 ) | ( n427  &  n653 ) | ( (~ n160)  &  n1677 ) | ( n653  &  n1677 ) ;
 assign n663 = ( n1288  &  n1289  &  n867  &  n1290  &  n1258 ) ;
 assign n664 = ( n1524  &  n2331  &  n2005  &  n2332  &  n1918  &  n2333 ) ;
 assign n665 = ( n1689  &  n1684  &  n1695  &  n1702  &  n621  &  n2334 ) ;
 assign n659 = ( n660  &  n661  &  n270  &  n662  &  n663  &  n664  &  n665 ) ;
 assign n667 = ( n1069 ) | ( n427 ) ;
 assign n666 = ( (~ n160)  &  n667 ) | ( n574  &  n667 ) ;
 assign n669 = ( n1226  &  n590 ) ;
 assign n670 = ( n1213 ) | ( n1316 ) ;
 assign n668 = ( (~ n333)  &  n441 ) | ( n441  &  n669 ) | ( (~ n333)  &  n670 ) | ( n669  &  n670 ) ;
 assign n673 = ( n511  &  n499  &  n1329 ) ;
 assign n671 = ( (~ n555) ) | ( n673 ) ;
 assign n675 = ( n72  &  n659  &  n666  &  n671  &  (~ n1663)  &  n1736 ) ;
 assign n674 = ( n801  &  n1734 ) ;
 assign n677 = ( n374 ) | ( n1256 ) ;
 assign n678 = ( n374 ) | ( n619 ) ;
 assign n679 = ( n374 ) | ( n1332 ) ;
 assign n680 = ( n184  &  (~ n237) ) | ( n184  &  n992 ) | ( (~ n237)  &  n1704 ) | ( n992  &  n1704 ) ;
 assign n676 = ( n677  &  n678  &  n679  &  n680 ) ;
 assign n681 = ( (~ n374)  &  (~ n649) ) | ( (~ n374)  &  (~ n1245) ) | ( (~ n374)  &  (~ n1325) ) ;
 assign n683 = ( (~ n174)  &  (~ n184) ) | ( (~ n184)  &  (~ n1739) ) ;
 assign n686 = ( (~ n237) ) | ( n456 ) ;
 assign n692 = ( (~ n1057)  &  n1184 ) ;
 assign n688 = ( n692  &  (~ n1344) ) | ( n692  &  (~ n1746) ) | ( n692  &  (~ n2336) ) ;
 assign n693 = ( n692  &  (~ n917) ) | ( n692  &  (~ n1586) ) ;
 assign n699 = ( (~ n614) ) | ( (~ n1063) ) | ( (~ n1339) ) ;
 assign n696 = ( n692  &  n699 ) | ( n692  &  (~ n1666) ) | ( n692  &  (~ n1747) ) ;
 assign n701 = ( (~ n1184) ) | ( n1224 ) ;
 assign n702 = ( n1587  &  n997 ) ;
 assign n700 = ( n701 ) | ( n702 ) ;
 assign n703 = ( (~ n184)  &  (~ n707) ) | ( (~ n184)  &  (~ n1226) ) ;
 assign n707 = ( n617  &  n1315 ) ;
 assign n706 = ( n374 ) | ( n707 ) ;
 assign n709 = ( n184 ) | ( n1319 ) ;
 assign n710 = ( n178 ) | ( n184 ) ;
 assign n711 = ( n184 ) | ( n1236 ) ;
 assign n712 = ( n184 ) | ( n1454 ) ;
 assign n713 = ( n1219 ) | ( n184 ) ;
 assign n714 = ( n184 ) | ( n1320 ) ;
 assign n715 = ( n1227 ) | ( n184 ) ;
 assign n716 = ( n2343  &  n1220 ) | ( n2343  &  n184 ) ;
 assign n708 = ( n709  &  n710  &  n711  &  n712  &  n713  &  n714  &  n715  &  n716 ) ;
 assign n718 = ( n1191 ) | ( n1211 ) ;
 assign n717 = ( n718 ) | ( n374 ) ;
 assign n719 = ( n236  &  (~ n374) ) | ( (~ n374)  &  (~ n1220) ) ;
 assign n723 = ( n172 ) | ( (~ n401) ) ;
 assign n722 = ( n366  &  n630  &  n887 ) ;
 assign n721 = ( (~ n401)  &  n723 ) | ( n723  &  n722 ) ;
 assign n725 = ( n313 ) | ( n1331 ) ;
 assign n726 = ( n313 ) | ( n187 ) ;
 assign n727 = ( (~ n392)  &  (~ n401) ) | ( (~ n401)  &  n773 ) | ( (~ n392)  &  n1083 ) | ( n773  &  n1083 ) ;
 assign n724 = ( n725  &  n726  &  n727 ) ;
 assign n732 = ( n58  &  n1250 ) ;
 assign n728 = ( (~ n180)  &  n732 ) | ( (~ n453)  &  n732 ) | ( n732  &  (~ n1222) ) ;
 assign n734 = ( n638  &  n634 ) ;
 assign n733 = ( (~ n392) ) | ( n734 ) ;
 assign n736 = ( n313 ) | ( n1236 ) ;
 assign n737 = ( n313 ) | ( n1319 ) ;
 assign n738 = ( n2509 ) | ( n313 ) ;
 assign n739 = ( n313 ) | ( n1454 ) ;
 assign n740 = ( n313 ) | ( n1469 ) ;
 assign n741 = ( n313 ) | ( n178 ) ;
 assign n742 = ( n313 ) | ( n1227 ) ;
 assign n743 = ( n2169  &  n313 ) | ( n2169  &  n370  &  n466 ) ;
 assign n735 = ( n736  &  n737  &  n738  &  n739  &  n740  &  n741  &  n742  &  n743 ) ;
 assign n745 = ( n277  &  n1585  &  n658 ) ;
 assign n746 = ( n1322  &  n1237 ) ;
 assign n744 = ( n722  &  n745  &  n746  &  n456 ) ;
 assign n748 = ( n1203 ) | ( n1217 ) ;
 assign n749 = ( n1282 ) | ( n1316 ) ;
 assign n750 = ( n1212 ) | ( n1282 ) ;
 assign n751 = ( n1267  &  n658 ) ;
 assign n747 = ( n277  &  (~ n439)  &  n649  &  n748  &  n749  &  n750  &  n751 ) ;
 assign n753 = ( n313 ) | ( n1396 ) ;
 assign n754 = ( n173 ) | ( (~ n401) ) ;
 assign n755 = ( n313  &  (~ n401) ) | ( (~ n401)  &  n744 ) | ( n313  &  n747 ) | ( n744  &  n747 ) ;
 assign n756 = ( (~ n392) ) | ( n842 ) ;
 assign n757 = ( n1474  &  n2011  &  n324  &  n2010  &  n2112  &  n1433 ) ;
 assign n752 = ( n323  &  n753  &  n754  &  n755  &  n756  &  n757 ) ;
 assign n759 = ( n574  &  n466 ) ;
 assign n761 = ( n657  &  n1397 ) ;
 assign n762 = ( n517  &  n1214 ) ;
 assign n758 = ( (~ n20)  &  (~ n356)  &  n370  &  n614  &  n617  &  n759  &  n761  &  n762 ) ;
 assign n765 = ( n1314  &  n1070 ) ;
 assign n763 = ( (~ n233)  &  n381  &  n654  &  n765  &  (~ n963) ) ;
 assign n767 = ( (~ n728)  &  n733  &  n1773  &  n1774 ) ;
 assign n768 = ( n1117  &  n1476  &  n1534  &  n269  &  n1390  &  n1447 ) ;
 assign n769 = ( n2341  &  n2342  &  n313 ) | ( n2341  &  n2342  &  n614 ) ;
 assign n770 = ( (~ n144)  &  n2168  &  n2206  &  n2337  &  n2338  &  n2340 ) ;
 assign n772 = ( n1066  &  n1317  &  n1705 ) ;
 assign n773 = ( n670  &  n472 ) ;
 assign n771 = ( n772  &  n773  &  n590  &  n614 ) ;
 assign n774 = ( n366 ) | ( n184 ) ;
 assign n776 = ( (~ n316) ) | ( (~ n340) ) | ( (~ n654) ) ;
 assign n778 = ( (~ n1127) ) | ( (~ n1343) ) | ( (~ n1578) ) ;
 assign n775 = ( (~ n184)  &  n776 ) | ( (~ n184)  &  n778 ) | ( (~ n184)  &  (~ n1062) ) ;
 assign n782 = ( n780 ) | ( n1033 ) ;
 assign n783 = ( n780 ) | ( n1233 ) ;
 assign n780 = ( (~ n1184) ) | ( n1231 ) ;
 assign n781 = ( n1195 ) | ( n1223 ) ;
 assign n779 = ( n782  &  n783  &  n780 ) | ( n782  &  n783  &  n781 ) ;
 assign n785 = ( n1588  &  n1342 ) ;
 assign n784 = ( n780 ) | ( n785 ) ;
 assign n786 = ( n151  &  (~ n781) ) | ( n151  &  (~ n1343) ) | ( n151  &  (~ n1825) ) ;
 assign n790 = ( n471  &  n765 ) ;
 assign n789 = ( n780 ) | ( n790 ) ;
 assign n794 = ( n151 ) | ( (~ n780) ) ;
 assign n793 = ( (~ n998) ) | ( (~ n1587) ) ;
 assign n791 = ( n794  &  n793 ) | ( n794  &  (~ n1424) ) ;
 assign n796 = ( (~ n179) ) | ( (~ n1347) ) ;
 assign n795 = ( n151  &  n796 ) | ( n151  &  (~ n997) ) ;
 assign n799 = ( n1058 ) | ( n806 ) ;
 assign n798 = ( n800  &  n1845 ) ;
 assign n800 = ( n1033  &  n673 ) ;
 assign n801 = ( n1167 ) | ( n1636 ) ;
 assign n804 = ( (~ n91) ) | ( n1636 ) ;
 assign n803 = ( n265  &  n507 ) ;
 assign n802 = ( n804  &  n801 ) | ( n804  &  n803  &  n508 ) ;
 assign n806 = ( n1228 ) | ( n1636 ) ;
 assign n807 = ( n1223 ) | ( n1316 ) ;
 assign n805 = ( n806 ) | ( n807 ) ;
 assign n809 = ( n1330  &  n1339 ) ;
 assign n810 = ( n434  &  n315 ) ;
 assign n811 = ( n1212 ) | ( n1216 ) ;
 assign n812 = ( n1217 ) | ( n1240 ) ;
 assign n808 = ( n809  &  n810  &  n187  &  n466  &  n811  &  n511  &  n812  &  n634 ) ;
 assign n814 = ( n1849  &  n1850  &  n418  &  n1851  &  n1852 ) ;
 assign n815 = ( (~ n14)  &  n1284  &  n1378 ) | ( n520  &  n1284  &  n1378 ) ;
 assign n816 = ( (~ n143) ) | ( n1319 ) ;
 assign n817 = ( (~ n14) ) | ( n1323 ) ;
 assign n819 = ( (~ n143)  &  n468  &  n2352 ) | ( n468  &  n808  &  n2352 ) ;
 assign n813 = ( (~ n11)  &  n512  &  n519  &  n814  &  n815  &  n816  &  n817  &  n819 ) ;
 assign n821 = ( n219 ) | ( n388 ) ;
 assign n822 = ( (~ n156) ) | ( n388 ) ;
 assign n820 = ( n821  &  n822  &  n810 ) | ( n821  &  n822  &  n388 ) ;
 assign n824 = ( n645  &  n434 ) ;
 assign n823 = ( n164 ) | ( n824 ) ;
 assign n828 = ( n649 ) | ( n827 ) ;
 assign n826 = ( n1245  &  n1738 ) ;
 assign n827 = ( (~ n1200) ) | ( n1224 ) ;
 assign n825 = ( n828  &  n826 ) | ( n828  &  n827 ) ;
 assign n829 = ( n608 ) | ( n441 ) ;
 assign n831 = ( n441 ) | ( n646 ) ;
 assign n832 = ( n441 ) | ( n1241 ) ;
 assign n833 = ( (~ n14)  &  (~ n147) ) | ( (~ n147)  &  n1747 ) ;
 assign n834 = ( n2379  &  n427 ) | ( n2379  &  n470 ) ;
 assign n835 = ( n1854  &  n953  &  n820  &  n644  &  n1607  &  n2380 ) ;
 assign n836 = ( (~ n19)  &  n1408  &  n1442  &  n1591  &  n2037  &  n2163  &  n2348  &  n2378 ) ;
 assign n837 = ( n1953  &  n1362  &  n2193  &  n2249  &  n2189  &  n920  &  n1364  &  n2377 ) ;
 assign n838 = ( n1483  &  n2143  &  n2105  &  n2323  &  n2106  &  n2126  &  n1484  &  n2376 ) ;
 assign n830 = ( n831  &  n832  &  n833  &  n834  &  n835  &  n836  &  n837  &  n838 ) ;
 assign n839 = ( n439  &  n531 ) | ( n531  &  (~ n1739) ) ;
 assign n842 = ( n608  &  n612 ) ;
 assign n840 = ( (~ n223)  &  n619 ) | ( (~ n223)  &  n827 ) | ( n619  &  n842 ) | ( n827  &  n842 ) ;
 assign n845 = ( n164 ) | ( n1322 ) ;
 assign n846 = ( n164 ) | ( n1237 ) ;
 assign n844 = ( n630  &  n1326 ) ;
 assign n843 = ( n845  &  n846  &  n844 ) | ( n845  &  n846  &  n164 ) ;
 assign n848 = ( (~ n164) ) | ( n855 ) ;
 assign n847 = ( (~ n456)  &  n848 ) | ( (~ n460)  &  n848 ) ;
 assign n849 = ( (~ n164)  &  (~ n1520) ) | ( (~ n164)  &  (~ n1585) ) ;
 assign n855 = ( n1200  &  n1208 ) ;
 assign n854 = ( (~ n649) ) | ( (~ n1704) ) ;
 assign n852 = ( (~ n608)  &  n855 ) | ( (~ n751)  &  n855 ) | ( n855  &  n854 ) ;
 assign n856 = ( n439  &  (~ n891) ) | ( (~ n649)  &  (~ n891) ) ;
 assign n858 = ( (~ n388)  &  n439 ) | ( (~ n388)  &  (~ n619) ) ;
 assign n861 = ( (~ n482) ) | ( n842 ) ;
 assign n864 = ( n1190 ) | ( n1282 ) ;
 assign n863 = ( n460  &  n277  &  n658  &  n864  &  n176  &  n456 ) ;
 assign n865 = ( (~ n164)  &  (~ n608) ) | ( n333  &  (~ n608) ) ;
 assign n867 = ( (~ n160) ) | ( n1256 ) ;
 assign n868 = ( (~ n160) ) | ( n1235 ) ;
 assign n869 = ( n1770 ) | ( n441 ) ;
 assign n870 = ( n427 ) | ( (~ n439) ) ;
 assign n871 = ( (~ n865)  &  n1332 ) | ( (~ n333)  &  n441  &  (~ n865) ) ;
 assign n872 = ( (~ n1140)  &  n1355 ) | ( n460  &  n1256  &  n1355 ) ;
 assign n873 = ( n2329  &  n1463  &  n2034  &  n2138  &  n1918  &  n1261  &  n1260  &  n1259 ) ;
 assign n874 = ( n1075  &  n1865  &  n676  &  n1814  &  n840  &  n1877  &  n1884  &  n2374 ) ;
 assign n866 = ( n867  &  n868  &  n869  &  n870  &  n871  &  n872  &  n873  &  n874 ) ;
 assign n876 = ( n1512 ) | ( n388 ) ;
 assign n877 = ( n1514 ) | ( n388 ) ;
 assign n875 = ( n876  &  n877  &  n626 ) | ( n876  &  n877  &  n388 ) ;
 assign n881 = ( (~ n1454) ) | ( (~ n1469) ) ;
 assign n878 = ( (~ n164)  &  (~ n634) ) | ( (~ n164)  &  (~ n656) ) | ( (~ n164)  &  n881 ) ;
 assign n885 = ( (~ n531) ) | ( n626 ) ;
 assign n883 = ( n1512  &  n1514 ) ;
 assign n882 = ( (~ n531)  &  n885 ) | ( n885  &  n883 ) ;
 assign n888 = ( (~ n531) ) | ( n890 ) ;
 assign n887 = ( n1235  &  n1326  &  n1771 ) ;
 assign n886 = ( (~ n531)  &  n888 ) | ( n888  &  n887 ) ;
 assign n892 = ( n2515 ) | ( n891 ) ;
 assign n893 = ( n2514 ) | ( n891 ) ;
 assign n890 = ( n172  &  n424 ) ;
 assign n891 = ( n1167 ) | ( (~ n1200) ) ;
 assign n889 = ( n892  &  n893  &  n890 ) | ( n892  &  n893  &  n891 ) ;
 assign n895 = ( n629  &  n2357  &  n184 ) | ( n629  &  n2357  &  n1312 ) ;
 assign n896 = ( n2063  &  n2257  &  n1996  &  n2356  &  n1963  &  n2043  &  n1962  &  n2355 ) ;
 assign n897 = ( n1995  &  n2053  &  n1460  &  n1400  &  n2354  &  n1956  &  n1086  &  n1954 ) ;
 assign n898 = ( n1773  &  n2340  &  n1528  &  n2124  &  n2170  &  n2203  &  n2353  &  n2035 ) ;
 assign n894 = ( n886  &  n889  &  n46  &  n721  &  n895  &  n896  &  n897  &  n898 ) ;
 assign n900 = ( n184  &  n759 ) | ( (~ n236)  &  n759 ) | ( n184  &  n1516 ) | ( (~ n236)  &  n1516 ) ;
 assign n901 = ( n2362  &  n2363 ) | ( n370  &  n2363 ) | ( n2362  &  n453 ) | ( n370  &  n453 ) ;
 assign n902 = ( (~ n531)  &  n1283 ) | ( n1102  &  n1283 ) | ( (~ n531)  &  n1676 ) | ( n1102  &  n1676 ) ;
 assign n903 = ( n634  &  n2256 ) | ( (~ n143)  &  n1265  &  n2256 ) ;
 assign n904 = ( n894  &  n708  &  n882  &  n633  &  n467  &  n2364 ) ;
 assign n905 = ( n1572  &  n1565  &  n1981  &  n1632  &  n1566  &  n2022  &  n1998  &  n2361 ) ;
 assign n906 = ( n1467  &  n1556  &  n1440  &  n1405  &  n2000  &  n2068  &  n1617  &  n2360 ) ;
 assign n907 = ( n2206  &  n2014  &  n1417  &  n1530  &  n1595  &  n2168  &  n1382  &  n2359 ) ;
 assign n899 = ( n900  &  n901  &  n902  &  n903  &  n904  &  n905  &  n906  &  n907 ) ;
 assign n908 = ( (~ n219)  &  (~ n1268) ) | ( (~ n1063)  &  (~ n1268) ) ;
 assign n909 = ( n13  &  n143 ) | ( n143  &  (~ n810) ) | ( n143  &  (~ n1747) ) ;
 assign n911 = ( (~ n333)  &  n2389 ) | ( n434  &  n2389 ) ;
 assign n912 = ( n866  &  n1890  &  n830  &  n1794  &  n1748  &  n899 ) ;
 assign n913 = ( n2385  &  n2388  &  n1923 ) | ( n2385  &  n2388  &  n990 ) ;
 assign n914 = ( (~ n157)  &  (~ n908)  &  n2019  &  n2059  &  n2073  &  n2164 ) ;
 assign n915 = ( n1398  &  n1550  &  n1462  &  n2025  &  n1952  &  n1427  &  n2381  &  n2383 ) ;
 assign n910 = ( n615  &  n314  &  n573  &  n911  &  n912  &  n913  &  n914  &  n915 ) ;
 assign n917 = ( n1705  &  n773 ) ;
 assign n916 = ( n164  &  (~ n848) ) | ( n617  &  (~ n848) ) | ( n164  &  n917 ) | ( n617  &  n917 ) ;
 assign n919 = ( (~ n531) ) | ( n2517 ) ;
 assign n920 = ( n2358 ) | ( n827 ) ;
 assign n918 = ( (~ n233)  &  n919  &  n920 ) | ( (~ n531)  &  n919  &  n920 ) ;
 assign n922 = ( (~ n511) ) | ( (~ n520) ) ;
 assign n921 = ( n233  &  n855 ) | ( (~ n638)  &  n855 ) | ( n855  &  n922 ) ;
 assign n924 = ( (~ n143)  &  (~ n333) ) | ( (~ n143)  &  n638 ) | ( (~ n333)  &  n811 ) | ( n638  &  n811 ) ;
 assign n925 = ( (~ n401)  &  n590 ) | ( (~ n401)  &  (~ n1138) ) | ( n590  &  n2410 ) | ( (~ n1138)  &  n2410 ) ;
 assign n926 = ( n2362  &  n2363 ) | ( n381  &  n2363 ) | ( n2362  &  n180 ) | ( n381  &  n180 ) ;
 assign n927 = ( n1076  &  n124  &  n918  &  n641  &  n365  &  n1808 ) ;
 assign n928 = ( n2031  &  n1431  &  n1172  &  n2409  &  n1304  &  n1959  &  n1373  &  n2407 ) ;
 assign n929 = ( n1621  &  n1858  &  n2024  &  n1287  &  n1299  &  n1297  &  n1546  &  n2405 ) ;
 assign n930 = ( n1391  &  n1994  &  n2062  &  n1987  &  n2123  &  n2104  &  n2015  &  n2404 ) ;
 assign n923 = ( n924  &  n430  &  n925  &  n926  &  n927  &  n928  &  n929  &  n930 ) ;
 assign n932 = ( n388 ) | ( (~ n935) ) ;
 assign n933 = ( n762 ) | ( n388 ) ;
 assign n931 = ( n932  &  n933  &  n628 ) | ( n932  &  n933  &  n388 ) ;
 assign n935 = ( (~ n1127) ) | ( (~ n1317) ) ;
 assign n934 = ( (~ n164)  &  n935 ) | ( (~ n164)  &  (~ n1678) ) ;
 assign n938 = ( n1224 ) | ( (~ n1250) ) ;
 assign n937 = ( n212  &  n938 ) ;
 assign n941 = ( n2516 ) | ( n827 ) ;
 assign n940 = ( (~ n233)  &  n319 ) ;
 assign n939 = ( n941  &  n940 ) | ( n941  &  n827 ) ;
 assign n943 = ( n2517 ) | ( n388 ) ;
 assign n944 = ( (~ n233) ) | ( n388 ) ;
 assign n945 = ( n388 ) | ( n617 ) ;
 assign n946 = ( n2395  &  n1087  &  n1069 ) | ( n2395  &  n1087  &  n164 ) ;
 assign n947 = ( n1613  &  n1380  &  n2199  &  n2002  &  n2069  &  n1379 ) ;
 assign n948 = ( n426  &  n334  &  n444  &  n2396  &  n1501  &  n939  &  n1801  &  n2397 ) ;
 assign n949 = ( n2001  &  n1564  &  n2259  &  n2088  &  n2044  &  n667  &  n2393  &  n2391 ) ;
 assign n942 = ( n943  &  n944  &  n945  &  n946  &  n947  &  n948  &  n949 ) ;
 assign n950 = ( (~ n184)  &  (~ n517) ) | ( (~ n184)  &  (~ n1127) ) ;
 assign n952 = ( (~ n693)  &  n1756  &  n1757  &  n1759  &  n1760  &  n1761 ) ;
 assign n953 = ( n829  &  n825  &  n217  &  n1853 ) ;
 assign n954 = ( n123  &  n668  &  n310  &  n183 ) ;
 assign n955 = ( n923  &  n1909  &  n916  &  n866  &  n894  &  n942 ) ;
 assign n956 = ( n2420  &  n2421  &  n2419  &  n2418  &  n2417  &  n2422  &  n2415  &  n2414 ) ;
 assign n957 = ( n1409  &  n2038  &  n1370  &  n1307  &  n2074  &  n1443  &  n1495  &  n2413 ) ;
 assign n958 = ( n2412  &  n1365  &  n2190  &  n1619  &  n1428  &  n1549  &  n221  &  n2411 ) ;
 assign n960 = ( n1343 ) | ( n891 ) ;
 assign n961 = ( n2511 ) | ( n388 ) ;
 assign n959 = ( n960  &  n961  &  n622 ) | ( n960  &  n961  &  n891 ) ;
 assign n963 = ( (~ n781) ) | ( (~ n1588) ) ;
 assign n962 = ( (~ n164)  &  n963 ) | ( (~ n164)  &  (~ n1262) ) ;
 assign n966 = ( n1343 ) | ( n388 ) ;
 assign n967 = ( n1262 ) | ( n388 ) ;
 assign n964 = ( (~ n32)  &  n966  &  n967 ) | ( n388  &  n966  &  n967 ) ;
 assign n968 = ( (~ n164)  &  (~ n807) ) | ( (~ n164)  &  (~ n1070) ) ;
 assign n970 = ( (~ n313)  &  (~ n2423) ) | ( (~ n313)  &  (~ n2424) ) ;
 assign n975 = ( n1200  &  n58 ) ;
 assign n973 = ( n975  &  (~ n1343) ) | ( n975  &  (~ n1588) ) | ( n975  &  (~ n1746) ) ;
 assign n976 = ( n590  &  n748  &  n781  &  n177 ) ;
 assign n977 = ( n333  &  (~ n471) ) | ( (~ n471)  &  (~ n1923) ) ;
 assign n981 = ( n1270  &  n1265 ) | ( n1745  &  n1265 ) | ( n1270  &  n1588 ) | ( n1745  &  n1588 ) ;
 assign n982 = ( n1343 ) | ( n184 ) ;
 assign n983 = ( (~ n32)  &  (~ n333) ) | ( (~ n32)  &  n669 ) | ( (~ n333)  &  n1580 ) | ( n669  &  n1580 ) ;
 assign n984 = ( (~ n239)  &  (~ n401) ) | ( (~ n239)  &  n976 ) | ( (~ n401)  &  n1775 ) | ( n976  &  n1775 ) ;
 assign n985 = ( (~ n977)  &  n1305  &  n1349  &  n1356  &  n1494  &  n2072  &  n2255 ) ;
 assign n986 = ( n923  &  n899  &  n1860  &  n1826  &  n1928  &  n1098  &  n959  &  n2438 ) ;
 assign n987 = ( n1386  &  n1631  &  n1429  &  n2032  &  n1407  &  n2039  &  n1290  &  n2432 ) ;
 assign n988 = ( n1415  &  n1477  &  n1393  &  n1451  &  n1478  &  n1452  &  n2012  &  n2431 ) ;
 assign n980 = ( n981  &  n982  &  n983  &  n984  &  n985  &  n986  &  n987  &  n988 ) ;
 assign n990 = ( n614  &  n470 ) ;
 assign n992 = ( n608  &  n460 ) ;
 assign n993 = ( n471  &  n997 ) ;
 assign n989 = ( n456  &  n773  &  (~ n793)  &  n990  &  n992  &  n993 ) ;
 assign n995 = ( n1058  &  n1600 ) ;
 assign n994 = ( (~ n356)  &  n790  &  (~ n793)  &  n995 ) ;
 assign n997 = ( n1257  &  n1333  &  n995 ) ;
 assign n998 = ( n1191 ) | ( n1321 ) ;
 assign n996 = ( n997  &  n670  &  n470  &  n998 ) ;
 assign n999 = ( n198  &  (~ n842) ) | ( n198  &  (~ n1936) ) ;
 assign n1002 = ( (~ n388)  &  (~ n864) ) | ( (~ n388)  &  (~ n1704) ) ;
 assign n1004 = ( (~ n313)  &  (~ n654) ) | ( (~ n313)  &  (~ n745) ) | ( (~ n313)  &  (~ n1239) ) ;
 assign n1007 = ( (~ n164)  &  (~ n1325) ) | ( (~ n164)  &  (~ n1585) ) | ( (~ n164)  &  (~ n1705) ) ;
 assign n1009 = ( n503  &  n798 ) | ( n503  &  n1735 ) ;
 assign n1008 = ( n97  &  (~ n105)  &  n134  &  n135  &  n498  &  n1009 ) ;
 assign n1011 = ( n567  &  (~ n1017)  &  n2450 ) | ( n798  &  (~ n1017)  &  n2450 ) ;
 assign n1010 = ( n675  &  n99  &  n1011 ) ;
 assign n1012 = ( n1230  &  n553 ) ;
 assign n1014 = ( n91  &  n553 ) ;
 assign n1016 = ( n1230  &  n1658 ) ;
 assign n1017 = ( n1230  &  n1642 ) ;
 assign n1018 = ( (~ n265)  &  n1938 ) ;
 assign n1019 = ( n1230  &  n1846 ) ;
 assign n1020 = ( (~ n265)  &  n555 ) ;
 assign n1021 = ( (~ n265)  &  n1657 ) ;
 assign n1023 = ( (~ n1066)  &  n1657 ) ;
 assign n1024 = ( (~ n1178)  &  n1658 ) ;
 assign n1025 = ( (~ n1178)  &  n1642 ) ;
 assign n1026 = ( (~ n1066)  &  n1938 ) ;
 assign n1027 = ( n555  &  (~ n1066) ) ;
 assign n1028 = ( (~ n1178)  &  n1846 ) ;
 assign n1032 = ( n674  &  (~ n1051) ) ;
 assign n1033 = ( n1223 ) | ( n1311 ) ;
 assign n1034 = ( (~ n657)  &  (~ n2454) ) ;
 assign n1038 = ( n91  &  n1658 ) ;
 assign n1039 = ( n91  &  n1642 ) ;
 assign n1040 = ( (~ n1346)  &  n1938 ) ;
 assign n1041 = ( n91  &  n1846 ) ;
 assign n1042 = ( n555  &  (~ n1346) ) ;
 assign n1043 = ( (~ n1346)  &  n1657 ) ;
 assign n1045 = ( (~ n1127)  &  (~ n2454) ) ;
 assign n1051 = ( n58  &  n1733 ) ;
 assign n1050 = ( n1051  &  (~ n1845) ) | ( (~ n1734)  &  (~ n1845) ) ;
 assign n1056 = ( n670 ) | ( n806 ) ;
 assign n1054 = ( n1033  &  n1845 ) ;
 assign n1060 = ( i_0_  &  n2507 ) | ( (~ i_2_)  &  n2507 ) ;
 assign n1057 = ( i_8_ ) | ( (~ n91) ) ;
 assign n1058 = ( n1234 ) | ( n1316 ) ;
 assign n1062 = ( n765  &  n761  &  n611  &  n759  &  n1775  &  n1776 ) ;
 assign n1063 = ( n266  &  n1247 ) ;
 assign n1064 = ( n1204 ) | ( n1218 ) ;
 assign n1065 = ( n634  &  n1454 ) ;
 assign n1066 = ( n1191 ) | ( n1213 ) ;
 assign n1061 = ( n1062  &  n654  &  n219  &  n1063  &  n617  &  n1064  &  n1065  &  n1066 ) ;
 assign n1068 = ( n807  &  n1677 ) ;
 assign n1069 = ( n1315  &  n669 ) ;
 assign n1070 = ( n1218 ) | ( n1223 ) ;
 assign n1071 = ( n1470  &  n1456  &  n651 ) ;
 assign n1067 = ( n608  &  (~ n793)  &  n1068  &  n1069  &  n1070  &  n1071 ) ;
 assign n1072 = ( (~ n934)  &  n1902  &  n1903  &  n1905  &  n1906  &  n1907 ) ;
 assign n1073 = ( (~ n962)  &  n1920  &  n1921 ) ;
 assign n1074 = ( n163  &  n369  &  (~ n878)  &  n1888 ) ;
 assign n1075 = ( n281  &  n1871  &  n1872  &  n1873  &  n1473  &  n1874  &  n1875  &  n1876 ) ;
 assign n1076 = ( (~ n921)  &  n1608  &  n1899  &  n1901 ) ;
 assign n1077 = ( n380  &  n394  &  n1854  &  n1426  &  n271  &  n290 ) ;
 assign n1078 = ( (~ n23)  &  n338  &  n1348  &  n2207  &  n2354  &  n2460  &  n2461  &  n2462 ) ;
 assign n1079 = ( (~ n531) ) | ( n574 ) ;
 assign n1081 = ( n1377  &  n1071 ) ;
 assign n1082 = ( n998  &  (~ n1105)  &  n1666 ) ;
 assign n1083 = ( n590  &  n1705 ) ;
 assign n1080 = ( (~ n20)  &  (~ n356)  &  n656  &  n707  &  n1081  &  n1082  &  n1083 ) ;
 assign n1085 = ( n622 ) | ( n827 ) ;
 assign n1086 = ( (~ n531) ) | ( n2358 ) ;
 assign n1087 = ( n1069 ) | ( n827 ) ;
 assign n1088 = ( (~ n33)  &  (~ n223) ) | ( (~ n33)  &  n1068  &  n1936 ) ;
 assign n1089 = ( n1619  &  n1620  &  n1621  &  n1622  &  n1623  &  n1624  &  n1625  &  n1626 ) ;
 assign n1090 = ( n1361  &  n1362  &  n1363  &  n1364  &  n1365  &  n1366  &  n1367  &  n1368 ) ;
 assign n1091 = ( (~ n531)  &  n1296 ) | ( n1080  &  n1296 ) ;
 assign n1092 = ( n1951  &  n939  &  n918  &  n882  &  n886  &  n1884  &  n840  &  n825 ) ;
 assign n1084 = ( n1085  &  n1086  &  n1087  &  n1088  &  n1089  &  n1090  &  n1091  &  n1092 ) ;
 assign n1094 = ( n1277 ) | ( n1424 ) ;
 assign n1095 = ( n1376 ) | ( n1277 ) ;
 assign n1096 = ( n1277 ) | ( n1425 ) ;
 assign n1097 = ( n1277 ) | ( n524 ) ;
 assign n1098 = ( n258  &  n284  &  (~ n973)  &  n1924  &  n1925  &  n1927 ) ;
 assign n1099 = ( n2006  &  n1419  &  n2448 ) | ( n2006  &  n1419  &  n1277 ) ;
 assign n1093 = ( n1094  &  n1095  &  n1096  &  n327  &  n1097  &  n1098  &  n51  &  n1099 ) ;
 assign n1102 = ( n574  &  n656 ) ;
 assign n1100 = ( (~ n32)  &  n315  &  n617  &  n761  &  (~ n776)  &  n1083  &  n1102 ) ;
 assign n1105 = ( n796 ) | ( (~ n1587) ) ;
 assign n1103 = ( (~ n388)  &  (~ n998) ) | ( (~ n388)  &  (~ n1068) ) | ( (~ n388)  &  n1105 ) ;
 assign n1108 = ( n1959  &  n945  &  n1960  &  n943  &  n1961  &  n1962  &  n1963  &  n1964 ) ;
 assign n1109 = ( n820  &  n1612  &  n1865 ) ;
 assign n1110 = ( n2356  &  n1879  &  n1853  &  n2395  &  n2426  &  n1369  &  n1303  &  n2465 ) ;
 assign n1107 = ( n1108  &  n959  &  n964  &  n931  &  n889  &  n875  &  n1109  &  n1110 ) ;
 assign n1111 = ( n827  &  n184 ) ;
 assign n1112 = ( (~ n427)  &  (~ n1324) ) | ( (~ n427)  &  (~ n1455) ) ;
 assign n1117 = ( n1526  &  n1527  &  n1528  &  n1529  &  n1530  &  n1531  &  n1532  &  n1533 ) ;
 assign n1118 = ( (~ n331)  &  n831  &  n1494  &  n1495  &  n1497  &  n1498  &  n1499  &  n1500 ) ;
 assign n1119 = ( n320  &  (~ n531) ) | ( n320  &  n1454 ) ;
 assign n1120 = ( n313  &  (~ n401) ) | ( n313  &  n646 ) | ( (~ n401)  &  n1329 ) | ( n646  &  n1329 ) ;
 assign n1121 = ( n1111  &  n1583 ) | ( n749  &  n1583 ) | ( n1111  &  n1126 ) | ( n749  &  n1126 ) ;
 assign n1122 = ( n164  &  (~ n1112) ) | ( (~ n1112)  &  n1127  &  n1456 ) ;
 assign n1123 = ( (~ n160)  &  n2467 ) | ( n1033  &  n2467 ) ;
 assign n1116 = ( n1117  &  n1118  &  n288  &  n1119  &  n1120  &  n1121  &  n1122  &  n1123 ) ;
 assign n1124 = ( (~ n160)  &  n184  &  (~ n392)  &  (~ n848)  &  (~ n1140) ) ;
 assign n1126 = ( n499  &  n1327 ) ;
 assign n1127 = ( n1211 ) | ( n1316 ) ;
 assign n1128 = ( n1191 ) | ( n1204 ) ;
 assign n1125 = ( n1126  &  n1127  &  n511  &  n1128 ) ;
 assign n1130 = ( n1588  &  n434  &  n718 ) ;
 assign n1129 = ( n1130  &  n670  &  n614  &  n807 ) ;
 assign n1131 = ( (~ n266)  &  (~ n2292) ) | ( (~ n1341)  &  (~ n2292) ) ;
 assign n1138 = ( (~ n184) ) | ( (~ n891) ) ;
 assign n1135 = ( (~ n316)  &  n1138 ) | ( n1138  &  (~ n1508) ) ;
 assign n1140 = ( n333 ) | ( (~ n441) ) ;
 assign n1139 = ( (~ n574)  &  n1140 ) | ( (~ n574)  &  (~ n1516) ) ;
 assign n1143 = ( (~ n184)  &  (~ n1397) ) | ( n350  &  (~ n1397) ) | ( n482  &  (~ n1397) ) ;
 assign n1146 = ( n617  &  (~ n1139) ) | ( (~ n237)  &  (~ n1139)  &  n1281 ) ;
 assign n1147 = ( (~ n1135)  &  n1274 ) | ( n456  &  (~ n1135)  &  n1965 ) ;
 assign n1148 = ( n1809  &  n2468  &  n2278 ) | ( n1809  &  n2468  &  n1129 ) ;
 assign n1149 = ( n2476  &  n2475  &  n2474  &  n2472 ) ;
 assign n1150 = ( n1793  &  n1804  &  n1173  &  n1703  &  n919  &  n2343  &  n2348  &  n1783 ) ;
 assign n1151 = ( n1779  &  n1888  &  n885  &  n828  &  n2338  &  n1782  &  n1338  &  n1261 ) ;
 assign n1152 = ( n1916  &  n767  &  n606  &  n1680  &  n1108  &  n1951  &  n1116  &  n2488 ) ;
 assign n1153 = ( n2485  &  n2484  &  n2483  &  n2482  &  n2481  &  n2480  &  n2479  &  n2478 ) ;
 assign n1145 = ( n1146  &  n1147  &  n1148  &  n1149  &  n1150  &  n1151  &  n1152  &  n1153 ) ;
 assign n1154 = ( n143  &  (~ n520) ) | ( n486  &  (~ n520) ) ;
 assign n1155 = ( (~ n164)  &  (~ n165) ) | ( (~ n165)  &  (~ n313) ) | ( (~ n165)  &  (~ n1268) ) ;
 assign n1157 = ( (~ n172)  &  n531 ) | ( n531  &  (~ n749) ) | ( n531  &  (~ n1469) ) ;
 assign n1161 = ( n2506  &  n827 ) | ( n2506  &  n864 ) ;
 assign n1162 = ( n1116  &  n1650  &  (~ n1659)  &  (~ n1664) ) ;
 assign n1163 = ( n1268  &  n1279 ) | ( n1334  &  n1279 ) | ( n1268  &  n1324 ) | ( n1334  &  n1324 ) ;
 assign n1164 = ( (~ n229)  &  n2505 ) | ( n1342  &  n2505 ) ;
 assign n1165 = ( n2503  &  n2504  &  n2173 ) | ( n2503  &  n2504  &  n1033 ) ;
 assign n1166 = ( n2502  &  n2501  &  n2500  &  n2497  &  n2496  &  n2495  &  n2492  &  n2491 ) ;
 assign n1167 = ( i_8_ ) | ( n38 ) ;
 assign n1169 = ( n1537  &  n1584 ) ;
 assign n1170 = ( n1521  &  n1485  &  n1118  &  n1501  &  n1504 ) ;
 assign n1171 = ( (~ n333)  &  n2327 ) | ( n574  &  n917  &  n2327 ) ;
 assign n1172 = ( (~ n333) ) | ( n1315 ) ;
 assign n1173 = ( (~ n333) ) | ( n617 ) ;
 assign n1174 = ( (~ n333)  &  n993 ) | ( n610  &  n993 ) | ( (~ n333)  &  (~ n1140) ) | ( n610  &  (~ n1140) ) ;
 assign n1175 = ( (~ n3)  &  n2170  &  n2203  &  n2322  &  n2323  &  n2324  &  n2325  &  n2326 ) ;
 assign n1176 = ( n589  &  n593  &  n123  &  n1721  &  n575  &  n1724  &  n573  &  n2328 ) ;
 assign n1178 = ( (~ i_6_) ) | ( i_7_ ) ;
 assign n1180 = ( i_3_ ) | ( i_4_ ) | ( (~ i_5_) ) ;
 assign n1182 = ( (~ i_0_)  &  (~ i_1_)  &  (~ i_2_) ) ;
 assign n1184 = ( (~ n1180)  &  n1182 ) ;
 assign n1189 = ( i_15_ ) | ( n453 ) ;
 assign n1190 = ( i_12_ ) | ( (~ i_13_) ) | ( (~ i_14_) ) ;
 assign n1191 = ( i_12_ ) | ( i_13_ ) | ( (~ i_14_) ) ;
 assign n1194 = ( (~ i_15_) ) | ( n453 ) ;
 assign n1195 = ( (~ i_12_) ) | ( (~ i_13_) ) | ( i_14_ ) ;
 assign n1198 = ( (~ i_3_)  &  i_4_  &  (~ i_5_) ) ;
 assign n1200 = ( n1182  &  n1198 ) ;
 assign n1202 = ( (~ i_9_) ) | ( (~ i_10_) ) | ( (~ i_11_) ) ;
 assign n1203 = ( (~ i_15_) ) | ( n1202 ) ;
 assign n1204 = ( i_15_ ) | ( n1202 ) ;
 assign n1206 = ( n1190 ) | ( n1204 ) ;
 assign n1205 = ( n1128  &  n1206 ) ;
 assign n1208 = ( (~ i_8_)  &  (~ n1178) ) ;
 assign n1209 = ( (~ i_3_)  &  i_4_  &  i_5_ ) ;
 assign n1210 = ( n1182  &  n1209 ) ;
 assign n1211 = ( (~ i_15_) ) | ( n215 ) ;
 assign n1212 = ( (~ i_12_) ) | ( i_13_ ) | ( i_14_ ) ;
 assign n1213 = ( i_15_ ) | ( n215 ) ;
 assign n1214 = ( n1066  &  n185 ) ;
 assign n1215 = ( (~ i_15_) ) | ( n180 ) ;
 assign n1216 = ( i_15_ ) | ( n180 ) ;
 assign n1217 = ( (~ i_12_) ) | ( (~ i_13_) ) | ( (~ i_14_) ) ;
 assign n1218 = ( (~ i_12_) ) | ( i_13_ ) | ( (~ i_14_) ) ;
 assign n1219 = ( n1189 ) | ( n1190 ) ;
 assign n1220 = ( n1189 ) | ( n1191 ) ;
 assign n1222 = ( (~ i_9_) ) | ( i_10_ ) | ( i_11_ ) ;
 assign n1223 = ( i_15_ ) | ( n1222 ) ;
 assign n1224 = ( (~ i_8_) ) | ( (~ n91) ) ;
 assign n1226 = ( n1216 ) | ( n1218 ) ;
 assign n1227 = ( n1189 ) | ( n1218 ) ;
 assign n1228 = ( (~ i_8_) ) | ( n38 ) ;
 assign n1229 = ( n1215 ) | ( n1218 ) ;
 assign n1230 = ( i_6_  &  i_7_ ) ;
 assign n1231 = ( (~ i_8_) ) | ( (~ n1230) ) ;
 assign n1233 = ( n1212 ) | ( n1223 ) ;
 assign n1234 = ( i_15_ ) | ( (~ n57) ) ;
 assign n1235 = ( n1204 ) | ( n1217 ) ;
 assign n1236 = ( n1189 ) | ( n1217 ) ;
 assign n1237 = ( n1204 ) | ( n1212 ) ;
 assign n1238 = ( (~ i_15_) ) | ( n452 ) ;
 assign n1239 = ( n1218 ) | ( n1238 ) ;
 assign n1240 = ( i_15_ ) | ( n452 ) ;
 assign n1241 = ( n1212 ) | ( n1240 ) ;
 assign n1242 = ( n1189 ) | ( n1212 ) ;
 assign n1243 = ( i_9_ ) | ( (~ i_10_) ) | ( (~ i_11_) ) ;
 assign n1244 = ( i_15_ ) | ( n1243 ) ;
 assign n1245 = ( n1191 ) | ( n1244 ) ;
 assign n1246 = ( n1190 ) | ( n1244 ) ;
 assign n1247 = ( n1190 ) | ( n1240 ) ;
 assign n1248 = ( n1216 ) | ( n1217 ) ;
 assign n1249 = ( (~ i_3_)  &  (~ i_4_)  &  (~ i_5_) ) ;
 assign n1250 = ( n1182  &  n1249 ) ;
 assign n1252 = ( (~ n552) ) | ( (~ n1250) ) ;
 assign n1253 = ( n180 ) | ( n1252 ) ;
 assign n1254 = ( n215 ) | ( n451 ) ;
 assign n1255 = ( n215 ) | ( n1252 ) ;
 assign n1256 = ( n1218 ) | ( n1244 ) ;
 assign n1257 = ( n1218 ) | ( n1234 ) ;
 assign n1259 = ( n1235 ) | ( n427 ) ;
 assign n1260 = ( n427 ) | ( n1206 ) ;
 assign n1261 = ( n427 ) | ( n1128 ) ;
 assign n1258 = ( n1259  &  n1260  &  n1261 ) ;
 assign n1263 = ( n1217 ) | ( n1223 ) ;
 assign n1264 = ( n1190 ) | ( n1223 ) ;
 assign n1262 = ( n1263  &  n1264  &  n265 ) ;
 assign n1265 = ( (~ n401)  &  (~ n855) ) ;
 assign n1267 = ( n1217 ) | ( n1244 ) ;
 assign n1268 = ( (~ n531)  &  n1265 ) ;
 assign n1269 = ( (~ n1138)  &  n1268 ) ;
 assign n1270 = ( (~ n198)  &  n1269 ) ;
 assign n1271 = ( n462  &  n1270 ) ;
 assign n1272 = ( (~ n229)  &  (~ n1140) ) ;
 assign n1274 = ( n1271  &  n1272 ) ;
 assign n1275 = ( n701  &  n1274 ) ;
 assign n1277 = ( (~ n1200) ) | ( n1231 ) ;
 assign n1276 = ( n1277  &  n1275 ) ;
 assign n1278 = ( (~ i_15_) ) | ( n1222 ) ;
 assign n1279 = ( (~ n223)  &  n263  &  (~ n1138) ) ;
 assign n1280 = ( n891  &  n1268 ) ;
 assign n1281 = ( n441  &  n1280 ) ;
 assign n1282 = ( (~ i_15_) ) | ( n1243 ) ;
 assign n1283 = ( (~ n160)  &  n891 ) ;
 assign n1285 = ( (~ n14) ) | ( n1226 ) ;
 assign n1286 = ( (~ n14) ) | ( n187 ) ;
 assign n1287 = ( (~ n143) ) | ( n1226 ) ;
 assign n1284 = ( n1285  &  n1286  &  n1287 ) ;
 assign n1288 = ( n1227 ) | ( n427 ) ;
 assign n1289 = ( n1064 ) | ( n427 ) ;
 assign n1290 = ( (~ n160) ) | ( n1070 ) ;
 assign n1292 = ( n1937 ) | ( n780 ) ;
 assign n1293 = ( n780 ) | ( n1257 ) ;
 assign n1294 = ( n164 ) | ( n1256 ) ;
 assign n1295 = ( n427 ) | ( n1256 ) ;
 assign n1291 = ( n1292  &  n1293  &  n677  &  n726  &  n1294  &  n1295  &  n602 ) ;
 assign n1297 = ( n319 ) | ( (~ n531) ) ;
 assign n1298 = ( n187 ) | ( n827 ) ;
 assign n1299 = ( (~ n531) ) | ( n1226 ) ;
 assign n1300 = ( n1262 ) | ( n827 ) ;
 assign n1301 = ( (~ n531) ) | ( n1262 ) ;
 assign n1302 = ( n2189  &  n2190  &  n2191  &  n2192  &  n2193  &  n2194 ) ;
 assign n1296 = ( n1297  &  n1298  &  n1299  &  n1300  &  n1301  &  n1302 ) ;
 assign n1304 = ( n1226 ) | ( n891 ) ;
 assign n1305 = ( n1262 ) | ( n891 ) ;
 assign n1306 = ( n1937 ) | ( n388 ) ;
 assign n1307 = ( n762 ) | ( n891 ) ;
 assign n1308 = ( n319 ) | ( n891 ) ;
 assign n1309 = ( n388 ) | ( n187 ) ;
 assign n1310 = ( n2197  &  n2198  &  n2199  &  n1880  &  n2200  &  n2201 ) ;
 assign n1303 = ( n1304  &  n1305  &  n1306  &  n1307  &  n1308  &  n1309  &  n1310 ) ;
 assign n1311 = ( i_12_ ) | ( (~ i_13_) ) | ( i_14_ ) ;
 assign n1312 = ( n1203 ) | ( n1311 ) ;
 assign n1313 = ( n1190 ) | ( n1215 ) ;
 assign n1314 = ( n1278 ) | ( n1311 ) ;
 assign n1315 = ( n1215 ) | ( n1311 ) ;
 assign n1316 = ( i_12_ ) | ( i_14_ ) | ( i_13_ ) ;
 assign n1318 = ( n1211 ) | ( n1212 ) ;
 assign n1317 = ( n1318  &  n458 ) ;
 assign n1319 = ( n1190 ) | ( n1194 ) ;
 assign n1320 = ( n1194 ) | ( n1311 ) ;
 assign n1321 = ( (~ i_15_) ) | ( (~ n57) ) ;
 assign n1322 = ( n1204 ) | ( n1311 ) ;
 assign n1323 = ( n1190 ) | ( n1238 ) ;
 assign n1324 = ( n1189 ) | ( n1311 ) ;
 assign n1325 = ( n750  &  n277 ) ;
 assign n1327 = ( n1203 ) | ( n1316 ) ;
 assign n1328 = ( n1203 ) | ( n1212 ) ;
 assign n1326 = ( n1327  &  n1328 ) ;
 assign n1329 = ( n1216 ) | ( n1311 ) ;
 assign n1330 = ( n1212 ) | ( n1215 ) ;
 assign n1331 = ( n1211 ) | ( n1311 ) ;
 assign n1332 = ( n1282 ) | ( n1311 ) ;
 assign n1333 = ( n1311 ) | ( n1321 ) ;
 assign n1334 = ( n1195 ) | ( n1203 ) ;
 assign n1336 = ( n427 ) | ( n1334 ) ;
 assign n1337 = ( n427 ) | ( n1328 ) ;
 assign n1338 = ( n427 ) | ( n1327 ) ;
 assign n1335 = ( n1336  &  n1337  &  n1338 ) ;
 assign n1339 = ( n1195 ) | ( n1238 ) ;
 assign n1340 = ( n1212 ) | ( n1238 ) ;
 assign n1341 = ( n1238 ) | ( n1316 ) ;
 assign n1342 = ( n1190 ) | ( n1278 ) ;
 assign n1344 = ( n1195 ) | ( n1278 ) ;
 assign n1345 = ( n1212 ) | ( n1278 ) ;
 assign n1346 = ( n1278 ) | ( n1316 ) ;
 assign n1343 = ( n1344  &  n1345  &  n1346 ) ;
 assign n1347 = ( n1234 ) | ( n1311 ) ;
 assign n1349 = ( (~ n855) ) | ( n1343 ) ;
 assign n1350 = ( (~ n855) ) | ( (~ n935) ) ;
 assign n1351 = ( (~ n855) ) | ( n1320 ) ;
 assign n1352 = ( n164 ) | ( n1314 ) ;
 assign n1348 = ( n1349  &  n1350  &  n1351  &  n1352 ) ;
 assign n1353 = ( n427 ) | ( n1320 ) ;
 assign n1354 = ( n427 ) | ( n1312 ) ;
 assign n1355 = ( (~ n160) ) | ( n1332 ) ;
 assign n1356 = ( (~ n160) ) | ( n1314 ) ;
 assign n1358 = ( n1966 ) | ( n780 ) ;
 assign n1359 = ( n780 ) | ( n1333 ) ;
 assign n1360 = ( n427 ) | ( n1332 ) ;
 assign n1357 = ( n1358  &  n1359  &  n679  &  n725  &  n1360  &  n604  &  n211 ) ;
 assign n1361 = ( n1512 ) | ( n827 ) ;
 assign n1362 = ( n219 ) | ( n827 ) ;
 assign n1363 = ( n827 ) | ( n1320 ) ;
 assign n1364 = ( n827 ) | ( n220 ) ;
 assign n1365 = ( (~ n531) ) | ( (~ n935) ) ;
 assign n1366 = ( n827 ) | ( (~ n935) ) ;
 assign n1367 = ( n827 ) | ( n1331 ) ;
 assign n1368 = ( n2160  &  n2161 ) ;
 assign n1370 = ( n891 ) | ( (~ n935) ) ;
 assign n1371 = ( (~ n233) ) | ( n891 ) ;
 assign n1372 = ( n388 ) | ( n1331 ) ;
 assign n1373 = ( n891 ) | ( n1315 ) ;
 assign n1374 = ( n1966 ) | ( n388 ) ;
 assign n1375 = ( n2162  &  n2163  &  n944  &  n1878  &  n2164  &  n2165 ) ;
 assign n1369 = ( n1370  &  n1371  &  n1372  &  n1373  &  n1374  &  n1375 ) ;
 assign n1376 = ( n1218 ) | ( n1321 ) ;
 assign n1377 = ( n1217 ) | ( n1234 ) ;
 assign n1379 = ( (~ n14) ) | ( n1229 ) ;
 assign n1380 = ( (~ n14) ) | ( n1248 ) ;
 assign n1381 = ( (~ n14) ) | ( n1239 ) ;
 assign n1382 = ( (~ n143) ) | ( n178 ) ;
 assign n1378 = ( n1379  &  n1380  &  n1381  &  n1382 ) ;
 assign n1383 = ( (~ n160) ) | ( n308 ) ;
 assign n1384 = ( (~ n160) ) | ( n517 ) ;
 assign n1385 = ( (~ n160) ) | ( n1248 ) ;
 assign n1386 = ( (~ n160) ) | ( n1263 ) ;
 assign n1388 = ( n427 ) | ( n1248 ) ;
 assign n1389 = ( n2138  &  n2139  &  n2140 ) ;
 assign n1391 = ( (~ n401) ) | ( n1229 ) ;
 assign n1392 = ( n313 ) | ( n1263 ) ;
 assign n1393 = ( (~ n401) ) | ( n1263 ) ;
 assign n1394 = ( n313 ) | ( n1229 ) ;
 assign n1395 = ( n2141  &  n2142  &  n1910  &  n1881  &  n2143  &  n2144 ) ;
 assign n1390 = ( n1391  &  n1392  &  n1393  &  n1394  &  n251  &  n1395 ) ;
 assign n1396 = ( n1212 ) | ( n1244 ) ;
 assign n1397 = ( n1212 ) | ( n1213 ) ;
 assign n1398 = ( (~ n855) ) | ( n1241 ) ;
 assign n1399 = ( (~ n855) ) | ( n1242 ) ;
 assign n1400 = ( (~ n855) ) | ( n1237 ) ;
 assign n1401 = ( n164 ) | ( n1242 ) ;
 assign n1402 = ( n164 ) | ( n811 ) ;
 assign n1403 = ( n164 ) | ( n1233 ) ;
 assign n1404 = ( (~ n855) ) | ( n1220 ) ;
 assign n1405 = ( (~ n160) ) | ( n1220 ) ;
 assign n1406 = ( (~ n160) ) | ( n1397 ) ;
 assign n1407 = ( (~ n160) ) | ( n265 ) ;
 assign n1408 = ( n427 ) | ( n266 ) ;
 assign n1409 = ( (~ n160) ) | ( n1066 ) ;
 assign n1410 = ( (~ n160) ) | ( n511 ) ;
 assign n1411 = ( (~ n160) ) | ( n1241 ) ;
 assign n1412 = ( n2119  &  n2120  &  n2121 ) ;
 assign n1413 = ( n313 ) | ( n265 ) ;
 assign n1414 = ( n313 ) | ( n1233 ) ;
 assign n1415 = ( n265 ) | ( (~ n401) ) ;
 assign n1416 = ( (~ n401) ) | ( n1233 ) ;
 assign n1417 = ( (~ n401) ) | ( n1242 ) ;
 assign n1418 = ( n2122  &  n1911  &  n2123  &  n2124  &  n2125  &  n2126 ) ;
 assign n1419 = ( n179 ) | ( n1277 ) ;
 assign n1420 = ( n780 ) | ( n179 ) ;
 assign n1421 = ( n179 ) | ( n701 ) ;
 assign n1422 = ( n1871  &  n2127  &  n2128  &  n753  &  n2129  &  n1874 ) ;
 assign n1423 = ( n1195 ) | ( n1215 ) ;
 assign n1424 = ( n1190 ) | ( n1321 ) ;
 assign n1425 = ( n1195 ) | ( n1321 ) ;
 assign n1427 = ( (~ n855) ) | ( n1323 ) ;
 assign n1428 = ( n307 ) | ( (~ n855) ) ;
 assign n1429 = ( (~ n855) ) | ( n1342 ) ;
 assign n1430 = ( (~ n855) ) | ( n1319 ) ;
 assign n1431 = ( (~ n855) ) | ( n1313 ) ;
 assign n1426 = ( n1427  &  n1428  &  n1429  &  n1430  &  n1431 ) ;
 assign n1433 = ( n313 ) | ( n864 ) ;
 assign n1434 = ( n374 ) | ( n864 ) ;
 assign n1435 = ( n374 ) | ( n1424 ) ;
 assign n1436 = ( n374 ) | ( n1425 ) ;
 assign n1437 = ( n164 ) | ( n864 ) ;
 assign n1438 = ( n1096  &  n116  &  n2098  &  n1094 ) ;
 assign n1432 = ( n1433  &  n1434  &  n1435  &  n1436  &  n1437  &  n1438 ) ;
 assign n1440 = ( (~ n160) ) | ( n165 ) ;
 assign n1441 = ( (~ n160) ) | ( n307 ) ;
 assign n1442 = ( n427 ) | ( n1339 ) ;
 assign n1443 = ( (~ n160) ) | ( n458 ) ;
 assign n1444 = ( (~ n160) ) | ( n1423 ) ;
 assign n1445 = ( (~ n160) ) | ( n1323 ) ;
 assign n1446 = ( n2099  &  n2100  &  n2101 ) ;
 assign n1439 = ( n1440  &  n1441  &  n1442  &  n1443  &  n276  &  n1444  &  n1445  &  n1446 ) ;
 assign n1448 = ( n313 ) | ( n1342 ) ;
 assign n1449 = ( n313 ) | ( n1344 ) ;
 assign n1450 = ( n313 ) | ( n1424 ) ;
 assign n1451 = ( (~ n401) ) | ( n1342 ) ;
 assign n1452 = ( (~ n401) ) | ( n1344 ) ;
 assign n1453 = ( n2102  &  n2103  &  n2104  &  n2105  &  n2106  &  n2107 ) ;
 assign n1447 = ( n1448  &  n1449  &  n1450  &  n1451  &  n1452  &  n1453 ) ;
 assign n1454 = ( n1194 ) | ( n1316 ) ;
 assign n1455 = ( n1244 ) | ( n1311 ) ;
 assign n1456 = ( n1316 ) | ( n1321 ) ;
 assign n1457 = ( (~ n855) ) | ( n1324 ) ;
 assign n1458 = ( n164 ) | ( n1329 ) ;
 assign n1459 = ( n164 ) | ( n1033 ) ;
 assign n1460 = ( (~ n855) ) | ( n1322 ) ;
 assign n1461 = ( n164 ) | ( n1324 ) ;
 assign n1462 = ( n646 ) | ( (~ n855) ) ;
 assign n1463 = ( (~ n160) ) | ( n749 ) ;
 assign n1464 = ( (~ n160) ) | ( n1341 ) ;
 assign n1465 = ( (~ n160) ) | ( n646 ) ;
 assign n1466 = ( n427 ) | ( n1341 ) ;
 assign n1467 = ( (~ n160) ) | ( n1454 ) ;
 assign n1468 = ( n2085  &  n2086  &  n2087  &  n2088 ) ;
 assign n1469 = ( n1194 ) | ( n1212 ) ;
 assign n1470 = ( n1190 ) | ( n1234 ) ;
 assign n1472 = ( n374 ) | ( n524 ) ;
 assign n1473 = ( n164 ) | ( n1246 ) ;
 assign n1474 = ( n313 ) | ( n750 ) ;
 assign n1475 = ( n374 ) | ( n1470 ) ;
 assign n1471 = ( n1472  &  n1473  &  n1474  &  n1475  &  n1097  &  n112  &  n117 ) ;
 assign n1477 = ( (~ n401) ) | ( n1264 ) ;
 assign n1478 = ( (~ n401) ) | ( n1345 ) ;
 assign n1479 = ( n313 ) | ( n1264 ) ;
 assign n1480 = ( n313 ) | ( n1345 ) ;
 assign n1481 = ( (~ n401) ) | ( n1469 ) ;
 assign n1482 = ( n313 ) | ( n1318 ) ;
 assign n1483 = ( n313 ) | ( n1247 ) ;
 assign n1484 = ( n313 ) | ( n1340 ) ;
 assign n1476 = ( n1477  &  n1478  &  n1479  &  n1480  &  n1481  &  n1482  &  n1483  &  n1484 ) ;
 assign n1486 = ( n441 ) | ( n1229 ) ;
 assign n1487 = ( (~ n333) ) | ( n517 ) ;
 assign n1488 = ( n441 ) | ( n308 ) ;
 assign n1489 = ( (~ n333) ) | ( n1229 ) ;
 assign n1490 = ( (~ n333) ) | ( n1248 ) ;
 assign n1491 = ( n1980  &  n1981  &  n1982 ) ;
 assign n1492 = ( (~ n333)  &  n1983 ) | ( n177  &  n1377  &  n1983 ) ;
 assign n1493 = ( n1973  &  n1974  &  n1975  &  n1976  &  n1977  &  n1978  &  n1979  &  n1969 ) ;
 assign n1485 = ( n1486  &  n1487  &  n1488  &  n1489  &  n1490  &  n1491  &  n1492  &  n1493 ) ;
 assign n1494 = ( (~ n333) ) | ( n1033 ) ;
 assign n1495 = ( (~ n333) ) | ( n657 ) ;
 assign n1497 = ( n441 ) | ( n1347 ) ;
 assign n1498 = ( n441 ) | ( n1127 ) ;
 assign n1499 = ( n1997  &  n1998  &  n1999  &  n2000  &  n2001  &  n2002 ) ;
 assign n1500 = ( n1991  &  n1992  &  n1993  &  n1994  &  n1995  &  n1996  &  n1984 ) ;
 assign n1502 = ( n441 ) | ( n520 ) ;
 assign n1503 = ( n441 ) | ( n511 ) ;
 assign n1501 = ( n1502  &  n1503  &  n404 ) ;
 assign n1505 = ( n441 ) | ( n1206 ) ;
 assign n1506 = ( n441 ) | ( n1128 ) ;
 assign n1504 = ( n1505  &  n1506  &  n405 ) ;
 assign n1507 = ( n1397  &  n1242 ) ;
 assign n1508 = ( n1033  &  n1233 ) ;
 assign n1509 = ( n1318  &  n762 ) ;
 assign n1510 = ( n388  &  n1270 ) ;
 assign n1511 = ( n657  &  n1455 ) ;
 assign n1512 = ( (~ n236)  &  n1454 ) ;
 assign n1514 = ( n1236  &  n1219  &  n1220 ) ;
 assign n1515 = ( (~ n1138)  &  n1265 ) ;
 assign n1516 = ( (~ n160)  &  n1515 ) ;
 assign n1517 = ( n374  &  (~ n531)  &  (~ n692)  &  (~ n1140) ) ;
 assign n1519 = ( n313  &  n1516 ) ;
 assign n1520 = ( n749  &  n1325 ) ;
 assign n1521 = ( (~ n333) ) | ( n2518 ) ;
 assign n1522 = ( n164 ) | ( n176 ) ;
 assign n1523 = ( n164 ) | ( n1267 ) ;
 assign n1524 = ( n427 ) | ( n1377 ) ;
 assign n1525 = ( n1816  &  n2008  &  n2009  &  n1730  &  n2010  &  n2011 ) ;
 assign n1526 = ( n313 ) | ( n1341 ) ;
 assign n1527 = ( n313 ) | ( n646 ) ;
 assign n1528 = ( (~ n401) ) | ( n1322 ) ;
 assign n1529 = ( n313 ) | ( n1324 ) ;
 assign n1530 = ( (~ n401) ) | ( n1454 ) ;
 assign n1531 = ( n313 ) | ( n1127 ) ;
 assign n1532 = ( n313 ) | ( n657 ) ;
 assign n1533 = ( n2012  &  n2013  &  n2014  &  n2015  &  n2016  &  n2017 ) ;
 assign n1535 = ( (~ n401) ) | ( n2509 ) ;
 assign n1534 = ( (~ n7)  &  n310  &  n314  &  n318  &  n389  &  n1535 ) ;
 assign n1538 = ( (~ n333) ) | ( n1344 ) ;
 assign n1539 = ( (~ n333) ) | ( n1323 ) ;
 assign n1540 = ( n441 ) | ( n1344 ) ;
 assign n1541 = ( n441 ) | ( n1424 ) ;
 assign n1542 = ( (~ n333) ) | ( n1319 ) ;
 assign n1543 = ( (~ n333) ) | ( n458 ) ;
 assign n1544 = ( n441 ) | ( n307 ) ;
 assign n1545 = ( (~ n147)  &  n2018  &  n2019  &  n2021  &  n2022  &  n2023 ) ;
 assign n1537 = ( n1538  &  n1539  &  n1540  &  n1541  &  n1542  &  n1543  &  n1544  &  n1545 ) ;
 assign n1546 = ( (~ n855) ) | ( n1229 ) ;
 assign n1547 = ( n164 ) | ( n177 ) ;
 assign n1548 = ( n164 ) | ( n1229 ) ;
 assign n1549 = ( n308 ) | ( (~ n855) ) ;
 assign n1550 = ( n812 ) | ( (~ n855) ) ;
 assign n1551 = ( n164 ) | ( n1239 ) ;
 assign n1552 = ( n2024  &  n1892  &  n2025 ) ;
 assign n1553 = ( n2026  &  n2027  &  n2028  &  n2029  &  n2030  &  n2031  &  n2032  &  n2033 ) ;
 assign n1555 = ( (~ n160) ) | ( n1219 ) ;
 assign n1556 = ( (~ n160) ) | ( n1469 ) ;
 assign n1557 = ( (~ n160) ) | ( n1247 ) ;
 assign n1558 = ( n427 ) | ( n1340 ) ;
 assign n1559 = ( n427 ) | ( n1330 ) ;
 assign n1560 = ( (~ n160) ) | ( n1330 ) ;
 assign n1561 = ( n2034  &  n2035  &  n2036 ) ;
 assign n1562 = ( n2037  &  n2038  &  n2039  &  n2040  &  n2041  &  n2042  &  n2043  &  n2044 ) ;
 assign n1554 = ( n1555  &  n1556  &  n1557  &  n1558  &  n1559  &  n1560  &  n1561  &  n1562 ) ;
 assign n1563 = ( (~ n333) ) | ( n1340 ) ;
 assign n1564 = ( n441 ) | ( n1330 ) ;
 assign n1565 = ( (~ n333) ) | ( n1219 ) ;
 assign n1566 = ( (~ n333) ) | ( n1469 ) ;
 assign n1567 = ( n441 ) | ( n524 ) ;
 assign n1568 = ( n2056  &  n2057  &  n2058 ) ;
 assign n1569 = ( (~ n333)  &  n2059 ) | ( n1470  &  n2059 ) ;
 assign n1570 = ( n2049  &  n2050  &  n2051  &  n2052  &  n2053  &  n2054  &  n2055  &  n2045 ) ;
 assign n1571 = ( n441 ) | ( n1233 ) ;
 assign n1572 = ( (~ n333) ) | ( n1220 ) ;
 assign n1573 = ( n441 ) | ( n179 ) ;
 assign n1574 = ( n441 ) | ( n1066 ) ;
 assign n1575 = ( n2071  &  n2072  &  n2073 ) ;
 assign n1576 = ( n179  &  n2074 ) | ( (~ n333)  &  n2074 ) ;
 assign n1577 = ( n1893  &  n2067  &  n2068  &  n2069  &  n2070  &  n2060 ) ;
 assign n1578 = ( n1342  &  n177 ) ;
 assign n1579 = ( (~ n143)  &  n263  &  n891 ) ;
 assign n1580 = ( (~ n333)  &  (~ n1138) ) ;
 assign n1581 = ( (~ n401)  &  n1580 ) ;
 assign n1582 = ( n388  &  (~ n531) ) ;
 assign n1583 = ( n164  &  (~ n198) ) ;
 assign n1584 = ( (~ n333)  &  (~ n1140) ) | ( (~ n333)  &  n1342 ) | ( (~ n1140)  &  n1425 ) | ( n1342  &  n1425 ) ;
 assign n1585 = ( n1195 ) | ( n1244 ) ;
 assign n1586 = ( n1195 ) | ( n1213 ) ;
 assign n1587 = ( n1195 ) | ( n1234 ) ;
 assign n1588 = ( n1191 ) | ( n1278 ) ;
 assign n1589 = ( n441 ) | ( n781 ) ;
 assign n1590 = ( n441 ) | ( n1587 ) ;
 assign n1591 = ( n441 ) | ( n645 ) ;
 assign n1592 = ( n441 ) | ( n1586 ) ;
 assign n1594 = ( n2254  &  n2255  &  n2256  &  n2257  &  n2258  &  n2259 ) ;
 assign n1595 = ( n453 ) | ( n451 ) ;
 assign n1596 = ( n453 ) | ( n1252 ) ;
 assign n1597 = ( n452 ) | ( n1252 ) ;
 assign n1598 = ( (~ n531)  &  n1519 ) ;
 assign n1599 = ( n164  &  n1519 ) ;
 assign n1600 = ( n1217 ) | ( n1321 ) ;
 assign n1601 = ( n630  &  n734 ) ;
 assign n1602 = ( n781  &  n645  &  n1586 ) ;
 assign n1603 = ( (~ n848)  &  n1279 ) ;
 assign n1604 = ( (~ n794)  &  (~ n975) ) ;
 assign n1608 = ( n164 ) | ( n748 ) ;
 assign n1607 = ( (~ n11)  &  n623  &  n961  &  n1608 ) ;
 assign n1610 = ( n427 ) | ( n460 ) ;
 assign n1611 = ( (~ n439) ) | ( n827 ) ;
 assign n1609 = ( n1610  &  n455  &  n114  &  n1611 ) ;
 assign n1613 = ( n2516 ) | ( n388 ) ;
 assign n1614 = ( n1908 ) | ( n388 ) ;
 assign n1615 = ( n2516 ) | ( n891 ) ;
 assign n1616 = ( n890 ) | ( n388 ) ;
 assign n1617 = ( n2511 ) | ( n891 ) ;
 assign n1618 = ( n388 ) | ( n466 ) ;
 assign n1612 = ( n1613  &  n1614  &  n1615  &  n1616  &  n1617  &  n1618 ) ;
 assign n1619 = ( (~ n531) ) | ( n1908 ) ;
 assign n1620 = ( n1908 ) | ( n827 ) ;
 assign n1621 = ( (~ n531) ) | ( n2516 ) ;
 assign n1622 = ( (~ n32) ) | ( n827 ) ;
 assign n1623 = ( (~ n32) ) | ( (~ n531) ) ;
 assign n1624 = ( (~ n531) ) | ( n2511 ) ;
 assign n1625 = ( n827 ) | ( n466 ) ;
 assign n1626 = ( n2247  &  n2248  &  n2249 ) ;
 assign n1628 = ( n427 ) | ( n466 ) ;
 assign n1629 = ( n427 ) | ( n748 ) ;
 assign n1630 = ( n890 ) | ( n427 ) ;
 assign n1631 = ( (~ n32) ) | ( (~ n160) ) ;
 assign n1632 = ( (~ n160) ) | ( n2511 ) ;
 assign n1633 = ( (~ n35) ) | ( n427 ) ;
 assign n1634 = ( n423  &  n426  &  n430  &  n433  &  (~ n437)  &  n2252 ) ;
 assign n1627 = ( n1628  &  n1629  &  n1630  &  n870  &  n1631  &  n1632  &  n1633  &  n1634 ) ;
 assign n1635 = ( i_0_ ) | ( (~ i_1_) ) | ( i_2_ ) ;
 assign n1636 = ( (~ n1249) ) | ( n1635 ) ;
 assign n1638 = ( (~ n552) ) | ( n1636 ) ;
 assign n1639 = ( i_0_  &  (~ i_1_) ) ;
 assign n1640 = ( n1330  &  n1328 ) ;
 assign n1641 = ( (~ n333)  &  n1583 ) ;
 assign n1642 = ( n1209  &  n1639 ) ;
 assign n1643 = ( (~ n223)  &  (~ n692) ) ;
 assign n1644 = ( n550 ) | ( n554 ) | ( n1017 ) | ( n103 ) ;
 assign n1646 = ( n555  &  (~ n1033) ) ;
 assign n1647 = ( n555  &  (~ n657) ) ;
 assign n1648 = ( n555  &  (~ n1127) ) ;
 assign n1649 = ( n1039 ) | ( n1025 ) | ( n1947 ) ;
 assign n1645 = ( n1027 ) | ( n1646 ) | ( n1647 ) | ( n1042 ) | ( n1648 ) | ( n1012 ) | ( n1020 ) | ( n1649 ) ;
 assign n1655 = ( n1502  &  n1583 ) | ( n1502  &  n1640  &  n1206 ) ;
 assign n1656 = ( n522  &  n297  &  n1554  &  n2303  &  n2302  &  n2301 ) ;
 assign n1650 = ( n167  &  (~ n526)  &  (~ n527)  &  (~ n530)  &  (~ n533)  &  n1505  &  n1655  &  n1656 ) ;
 assign n1657 = ( n553  &  (~ n1167) ) ;
 assign n1658 = ( n1198  &  n1639 ) ;
 assign n1660 = ( (~ n657)  &  n1657 ) ;
 assign n1661 = ( (~ n1127)  &  n1657 ) ;
 assign n1662 = ( n1948 ) | ( n1945 ) | ( n1021 ) | ( n1016 ) | ( n1038 ) | ( n1024 ) ;
 assign n1659 = ( n1043 ) | ( n1660 ) | ( n1023 ) | ( n1661 ) | ( n1014 ) | ( n1662 ) ;
 assign n1663 = ( n83 ) | ( n78 ) | ( n87 ) ;
 assign n1664 = ( n104 ) | ( n565 ) | ( n1663 ) ;
 assign n1666 = ( n220  &  n572 ) ;
 assign n1668 = ( (~ n160) ) | ( n1064 ) ;
 assign n1669 = ( (~ n160) ) | ( n1312 ) ;
 assign n1670 = ( (~ n160) ) | ( n748 ) ;
 assign n1667 = ( n1668  &  n618  &  n1669  &  n1670 ) ;
 assign n1672 = ( n427 ) | ( n1245 ) ;
 assign n1673 = ( n427 ) | ( n1246 ) ;
 assign n1674 = ( n427 ) | ( n750 ) ;
 assign n1675 = ( n427 ) | ( n749 ) ;
 assign n1676 = ( n1320  &  n1227 ) ;
 assign n1677 = ( n470  &  n993 ) ;
 assign n1678 = ( n1586  &  n718 ) ;
 assign n1681 = ( n427 ) | ( (~ n1105) ) ;
 assign n1682 = ( n427 ) | ( n619 ) ;
 assign n1683 = ( n2329  &  n2330 ) ;
 assign n1680 = ( n633  &  n629  &  n641  &  n637  &  n1681  &  n644  &  n1682  &  n1683 ) ;
 assign n1685 = ( n427 ) | ( n1066 ) ;
 assign n1686 = ( n427 ) | ( n185 ) ;
 assign n1687 = ( n427 ) | ( n1318 ) ;
 assign n1688 = ( n427 ) | ( n1127 ) ;
 assign n1684 = ( n1685  &  n282  &  n256  &  n1686  &  n1687  &  n1688  &  n627 ) ;
 assign n1690 = ( n427 ) | ( n1264 ) ;
 assign n1691 = ( n427 ) | ( n265 ) ;
 assign n1692 = ( (~ n32) ) | ( n427 ) ;
 assign n1693 = ( n427 ) | ( n1345 ) ;
 assign n1694 = ( n427 ) | ( n1346 ) ;
 assign n1689 = ( n1690  &  n1691  &  n1692  &  n257  &  n283  &  n1693  &  n1694 ) ;
 assign n1696 = ( n1220 ) | ( n427 ) ;
 assign n1697 = ( n165 ) | ( n427 ) ;
 assign n1698 = ( n1236 ) | ( n427 ) ;
 assign n1699 = ( n1219 ) | ( n427 ) ;
 assign n1700 = ( n427 ) | ( n1469 ) ;
 assign n1701 = ( n427 ) | ( n1454 ) ;
 assign n1695 = ( n1696  &  n1697  &  n1698  &  n1699  &  n1700  &  n1701  &  n625 ) ;
 assign n1703 = ( n427 ) | ( n608 ) ;
 assign n1702 = ( n1703  &  n620  &  n1667  &  n1610  &  n1295  &  n1360 ) ;
 assign n1704 = ( n1332  &  n1256 ) ;
 assign n1705 = ( n1331  &  n187 ) ;
 assign n1706 = ( n441 ) | ( n1328 ) ;
 assign n1707 = ( n441 ) | ( n1327 ) ;
 assign n1708 = ( n441 ) | ( n1237 ) ;
 assign n1709 = ( n441 ) | ( n1322 ) ;
 assign n1711 = ( (~ n333) ) | ( n1235 ) ;
 assign n1712 = ( (~ n333) ) | ( n1206 ) ;
 assign n1713 = ( n173 ) | ( (~ n333) ) ;
 assign n1714 = ( n172 ) | ( (~ n333) ) ;
 assign n1715 = ( (~ n333) ) | ( n1128 ) ;
 assign n1716 = ( (~ n333) ) | ( n1334 ) ;
 assign n1710 = ( n1711  &  n1712  &  n1713  &  n1714  &  n1715  &  n1716  &  n588 ) ;
 assign n1718 = ( n441 ) | ( n1315 ) ;
 assign n1719 = ( n441 ) | ( n590 ) ;
 assign n1720 = ( n441 ) | ( n1226 ) ;
 assign n1717 = ( n1718  &  n616  &  n1719  &  n1720 ) ;
 assign n1722 = ( n441 ) | ( n1070 ) ;
 assign n1723 = ( n441 ) | ( n1314 ) ;
 assign n1721 = ( n1722  &  n1723  &  n869 ) ;
 assign n1725 = ( n277 ) | ( (~ n333) ) ;
 assign n1726 = ( (~ n333) ) | ( n750 ) ;
 assign n1727 = ( (~ n333) ) | ( n1246 ) ;
 assign n1728 = ( (~ n333) ) | ( n1245 ) ;
 assign n1729 = ( (~ n333) ) | ( n749 ) ;
 assign n1730 = ( n441 ) | ( n176 ) ;
 assign n1731 = ( (~ n333) ) | ( n1396 ) ;
 assign n1732 = ( n326  &  n1710  &  n579  &  n2092  &  n2261  &  n2127 ) ;
 assign n1724 = ( n1725  &  n1726  &  n1727  &  n1728  &  n1729  &  n1730  &  n1731  &  n1732 ) ;
 assign n1733 = ( n1209  &  (~ n1635) ) ;
 assign n1735 = ( n1180 ) | ( (~ n1208) ) | ( n1635 ) ;
 assign n1734 = ( n1735  &  n567 ) ;
 assign n1736 = ( n38 ) | ( (~ n161) ) | ( n1635 ) ;
 assign n1738 = ( n1267  &  n1246  &  n1520 ) ;
 assign n1739 = ( n649  &  n826 ) ;
 assign n1741 = ( n374 ) | ( n749 ) ;
 assign n1743 = ( n374 ) | ( n1267 ) ;
 assign n1744 = ( n374 ) | ( n1246 ) ;
 assign n1740 = ( (~ n681)  &  n1741  &  n1743  &  n1744 ) ;
 assign n1745 = ( n807  &  n765 ) ;
 assign n1746 = ( n781  &  n471  &  n1745 ) ;
 assign n1747 = ( n470  &  n645 ) ;
 assign n1749 = ( (~ n692) ) | ( n1340 ) ;
 assign n1750 = ( (~ n692) ) | ( n1341 ) ;
 assign n1751 = ( (~ n692) ) | ( n810 ) ;
 assign n1752 = ( (~ n692) ) | ( n812 ) ;
 assign n1753 = ( (~ n692) ) | ( n1241 ) ;
 assign n1754 = ( n646 ) | ( (~ n692) ) ;
 assign n1748 = ( (~ n696)  &  n1749  &  n1750  &  n1751  &  n1752  &  n1753  &  n1754 ) ;
 assign n1756 = ( (~ n692) ) | ( n1397 ) ;
 assign n1757 = ( n657 ) | ( (~ n692) ) ;
 assign n1759 = ( (~ n692) ) | ( n1908 ) ;
 assign n1760 = ( (~ n692) ) | ( n762 ) ;
 assign n1761 = ( (~ n692) ) | ( (~ n935) ) ;
 assign n1763 = ( (~ n692) ) | ( n1345 ) ;
 assign n1764 = ( (~ n692) ) | ( n1346 ) ;
 assign n1765 = ( (~ n32) ) | ( (~ n692) ) ;
 assign n1766 = ( (~ n692) ) | ( n1263 ) ;
 assign n1767 = ( (~ n692) ) | ( n1233 ) ;
 assign n1768 = ( (~ n692) ) | ( n1033 ) ;
 assign n1762 = ( (~ n688)  &  n1763  &  n1764  &  n1765  &  n1766  &  n1767  &  n1768 ) ;
 assign n1770 = ( n1064  &  n1312  &  n619 ) ;
 assign n1771 = ( n1334  &  n1205 ) ;
 assign n1773 = ( (~ n732) ) | ( n1202 ) ;
 assign n1774 = ( n313 ) | ( n574 ) ;
 assign n1775 = ( n1262  &  n622 ) ;
 assign n1776 = ( n185  &  (~ n236)  &  n517  &  n748  &  n1312  &  n1588 ) ;
 assign n1777 = ( n184 ) | ( n1327 ) ;
 assign n1778 = ( n1064 ) | ( n184 ) ;
 assign n1779 = ( n1915 ) | ( n184 ) ;
 assign n1780 = ( n299  &  n2132  &  n2110  &  n2148  &  n2111  &  n2147 ) ;
 assign n1781 = ( n374 ) | ( n1320 ) ;
 assign n1782 = ( n374 ) | ( n574 ) ;
 assign n1783 = ( n626 ) | ( n374 ) ;
 assign n1785 = ( n374 ) | ( n466 ) ;
 assign n1786 = ( n1227 ) | ( n374 ) ;
 assign n1787 = ( n2149  &  n300  &  n2090 ) ;
 assign n1788 = ( n374 ) | ( n517 ) ;
 assign n1789 = ( n374 ) | ( n185 ) ;
 assign n1790 = ( n374 ) | ( n308 ) ;
 assign n1791 = ( n374 ) | ( n307 ) ;
 assign n1792 = ( n374 ) | ( n1127 ) ;
 assign n1793 = ( n628 ) | ( n374 ) ;
 assign n1795 = ( n184 ) | ( n1341 ) ;
 assign n1796 = ( n184 ) | ( n266 ) ;
 assign n1797 = ( n184 ) | ( n1339 ) ;
 assign n1798 = ( n184 ) | ( n812 ) ;
 assign n1799 = ( n184 ) | ( n1239 ) ;
 assign n1800 = ( n184 ) | ( n1323 ) ;
 assign n1794 = ( n301  &  n1795  &  n1796  &  n1797  &  n1798  &  n302  &  n1799  &  n1800 ) ;
 assign n1802 = ( n374 ) | ( n499 ) ;
 assign n1803 = ( n1226 ) | ( n374 ) ;
 assign n1804 = ( n2517 ) | ( n374 ) ;
 assign n1805 = ( n374 ) | ( n1423 ) ;
 assign n1806 = ( n374 ) | ( n1330 ) ;
 assign n1807 = ( n2152  &  n2076  &  n2133 ) ;
 assign n1801 = ( n1802  &  n1803  &  n1804  &  n706  &  n384  &  n1805  &  n1806  &  n1807 ) ;
 assign n1809 = ( n2517 ) | ( n184 ) ;
 assign n1811 = ( n184 ) | ( n1330 ) ;
 assign n1812 = ( n184 ) | ( n499 ) ;
 assign n1813 = ( n2077  &  n2131  &  n2114  &  n2151  &  n2115  &  n2153 ) ;
 assign n1808 = ( n52  &  n53  &  (~ n703)  &  n1809  &  n1811  &  n1812  &  n1813 ) ;
 assign n1816 = ( n374 ) | ( n176 ) ;
 assign n1817 = ( n1915 ) | ( n374 ) ;
 assign n1814 = ( (~ n683)  &  n686  &  n1434  &  n1740  &  n1816  &  n1817 ) ;
 assign n1819 = ( n374 ) | ( n1128 ) ;
 assign n1820 = ( n374 ) | ( n1334 ) ;
 assign n1821 = ( n374 ) | ( n1235 ) ;
 assign n1822 = ( n374 ) | ( n1206 ) ;
 assign n1823 = ( n374 ) | ( n1328 ) ;
 assign n1824 = ( n374 ) | ( n1327 ) ;
 assign n1818 = ( n1819  &  n1820  &  n1821  &  n1822  &  n1823  &  n1824  &  n373 ) ;
 assign n1825 = ( n471  &  n807  &  n785 ) ;
 assign n1828 = ( (~ n151) ) | ( n1233 ) ;
 assign n1829 = ( (~ n151) ) | ( n1033 ) ;
 assign n1830 = ( (~ n151) ) | ( n1314 ) ;
 assign n1831 = ( (~ n151) ) | ( n177 ) ;
 assign n1832 = ( (~ n151) ) | ( n1262 ) ;
 assign n1833 = ( (~ n151) ) | ( n1070 ) ;
 assign n1826 = ( (~ n786)  &  n789  &  n1828  &  n1829  &  n1830  &  n1831  &  n1832  &  n1833 ) ;
 assign n1835 = ( n1343 ) | ( n780 ) ;
 assign n1836 = ( n780 ) | ( n177 ) ;
 assign n1837 = ( n1262 ) | ( n780 ) ;
 assign n1834 = ( n1835  &  n784  &  n1836  &  n1837 ) ;
 assign n1840 = ( n780 ) | ( n1347 ) ;
 assign n1842 = ( n1826  &  n995 ) | ( n1826  &  n780 ) ;
 assign n1843 = ( n1359  &  n1420  &  n1917  &  n1293  &  n1292  &  n1358  &  n2205  &  n2171 ) ;
 assign n1844 = ( i_0_  &  i_1_  &  (~ i_2_) ) ;
 assign n1845 = ( n508  &  n803 ) ;
 assign n1846 = ( n1249  &  n1639 ) ;
 assign n1848 = ( (~ n38)  &  n1846 ) ;
 assign n1847 = ( n1028 ) | ( n1848 ) | ( n1019 ) | ( n1041 ) ;
 assign n1849 = ( (~ n14) ) | ( n178 ) ;
 assign n1850 = ( (~ n14) ) | ( n1319 ) ;
 assign n1851 = ( (~ n14) ) | ( n466 ) ;
 assign n1852 = ( (~ n14) ) | ( n2513 ) ;
 assign n1853 = ( n1739 ) | ( n388 ) ;
 assign n1856 = ( n164 ) | ( n1241 ) ;
 assign n1857 = ( n164 ) | ( n646 ) ;
 assign n1858 = ( n1771 ) | ( n164 ) ;
 assign n1859 = ( n164 ) | ( n1323 ) ;
 assign n1854 = ( (~ n154)  &  n218  &  n365  &  n823  &  n1856  &  n1857  &  n1858  &  n1859 ) ;
 assign n1861 = ( n172 ) | ( (~ n855) ) ;
 assign n1862 = ( (~ n855) ) | ( n1235 ) ;
 assign n1863 = ( (~ n855) ) | ( n1771 ) ;
 assign n1864 = ( n255  &  n366 ) | ( n255  &  (~ n855) ) ;
 assign n1860 = ( n1861  &  n1862  &  n1863  &  n1864 ) ;
 assign n1868 = ( n1915 ) | ( n388 ) ;
 assign n1869 = ( n751 ) | ( n891 ) ;
 assign n1870 = ( n1520 ) | ( n891 ) ;
 assign n1865 = ( (~ n856)  &  (~ n858)  &  n861  &  n1868  &  n1869  &  n1870 ) ;
 assign n1871 = ( n164 ) | ( n1396 ) ;
 assign n1872 = ( n1770 ) | ( n164 ) ;
 assign n1873 = ( n176 ) | ( (~ n855) ) ;
 assign n1874 = ( n164 ) | ( n1245 ) ;
 assign n1875 = ( n1522  &  n1437  &  n1523 ) ;
 assign n1876 = ( n321  &  n843  &  (~ n847)  &  (~ n849)  &  (~ n852)  &  n1294  &  n1860  &  n2172 ) ;
 assign n1878 = ( n2515 ) | ( n388 ) ;
 assign n1879 = ( n2358 ) | ( n388 ) ;
 assign n1880 = ( n2514 ) | ( n388 ) ;
 assign n1881 = ( n313 ) | ( n173 ) ;
 assign n1882 = ( n1630  &  n1970  &  n2251 ) ;
 assign n1883 = ( (~ n144)  &  n440  &  n1289  &  n1354  &  n1504  &  n1682  &  n1818  &  n2345 ) ;
 assign n1877 = ( n1878  &  n1879  &  n1616  &  n1880  &  n1881  &  n1629  &  n1882  &  n1883 ) ;
 assign n1887 = ( n1915 ) | ( n827 ) ;
 assign n1884 = ( (~ n15)  &  (~ n839)  &  n1611  &  n1887 ) ;
 assign n1888 = ( n164 ) | ( n574 ) ;
 assign n1891 = ( n827 ) | ( n574 ) ;
 assign n1892 = ( n164 ) | ( n178 ) ;
 assign n1893 = ( n441 ) | ( n1242 ) ;
 assign n1894 = ( n2197  &  n2162  &  n1991  &  n1618 ) ;
 assign n1895 = ( n1074  &  n875  &  n43  &  n814  &  n593  &  n735  &  n1695  &  n2369 ) ;
 assign n1896 = ( n2194  &  n1363  &  n1955  &  n1625  &  n2192  &  n1361  &  n2368  &  n2367 ) ;
 assign n1890 = ( n1891  &  n1892  &  n1401  &  n1461  &  n1893  &  n1894  &  n1895  &  n1896 ) ;
 assign n1898 = ( n180 ) | ( n451 ) ;
 assign n1899 = ( (~ n855) ) | ( n1329 ) ;
 assign n1901 = ( n811 ) | ( (~ n855) ) ;
 assign n1902 = ( n164 ) | ( n185 ) ;
 assign n1903 = ( n164 ) | ( n1066 ) ;
 assign n1905 = ( n164 ) | ( n1397 ) ;
 assign n1906 = ( n164 ) | ( n657 ) ;
 assign n1907 = ( n164 ) | ( n307 ) ;
 assign n1908 = ( n718  &  n340 ) ;
 assign n1910 = ( n313 ) | ( n517 ) ;
 assign n1911 = ( n313 ) | ( n1397 ) ;
 assign n1912 = ( (~ n3)  &  n1488  &  n1544  &  n1986  &  n2103  &  n2142 ) ;
 assign n1913 = ( n1366  &  n2399  &  n1298  &  n1367  &  n2070  &  n1620  &  n2191  &  n2398 ) ;
 assign n1914 = ( n515  &  n1684  &  n44  &  n1072  &  n931  &  n2402  &  n2403  &  n2401 ) ;
 assign n1909 = ( (~ n7)  &  n1482  &  n1531  &  n1910  &  n1911  &  n1912  &  n1913  &  n1914 ) ;
 assign n1915 = ( n630  &  n746 ) ;
 assign n1917 = ( n780 ) | ( n807 ) ;
 assign n1918 = ( n1915 ) | ( n427 ) ;
 assign n1919 = ( n2426  &  n2349  &  n1085  &  n2331  &  n779  &  n2425 ) ;
 assign n1916 = ( n1917  &  n1887  &  n1918  &  n678  &  n1868  &  n1817  &  n603  &  n1919 ) ;
 assign n1920 = ( n164 ) | ( n1342 ) ;
 assign n1921 = ( n1343 ) | ( n164 ) ;
 assign n1923 = ( (~ n160)  &  n1271 ) ;
 assign n1924 = ( (~ n975) ) | ( n1033 ) ;
 assign n1925 = ( (~ n975) ) | ( n1262 ) ;
 assign n1927 = ( (~ n975) ) | ( n1233 ) ;
 assign n1929 = ( n1745  &  n427 ) | ( n388  &  n427 ) | ( n1745  &  n471 ) | ( n388  &  n471 ) ;
 assign n1931 = ( n441  &  (~ n968) ) | ( n574  &  (~ n968)  &  n1825 ) ;
 assign n1932 = ( (~ n29)  &  n1352  &  n1403  &  n1459  &  n1571  &  n1589  &  n1997 ) ;
 assign n1933 = ( n1721  &  n1834  &  n843  &  n1335  &  n1689  &  n578 ) ;
 assign n1934 = ( n1916  &  n964  &  n1073  &  n1877  &  n1890  &  n942 ) ;
 assign n1935 = ( (~ n15)  &  n1300  &  n1547  &  n1622  &  n1872  &  n2160  &  n2428  &  n2429 ) ;
 assign n1928 = ( (~ n970)  &  n1258  &  n1929  &  n1931  &  n1932  &  n1933  &  n1934  &  n1935 ) ;
 assign n1936 = ( n614  &  n765  &  n773 ) ;
 assign n1937 = ( n1377  &  n1470  &  n537 ) ;
 assign n1938 = ( n58  &  (~ n1180)  &  (~ n1635) ) ;
 assign n1939 = ( (~ n657)  &  n1938 ) ;
 assign n1940 = ( (~ n1127)  &  n1938 ) ;
 assign n1941 = ( (~ n1033)  &  n1938 ) ;
 assign n1945 = ( (~ n1033)  &  n1657 ) ;
 assign n1946 = ( (~ n555)  &  n674 ) ;
 assign n1947 = ( (~ n38)  &  n1642 ) ;
 assign n1948 = ( (~ n38)  &  n1658 ) ;
 assign n1950 = ( (~ n91)  &  (~ n1230) ) ;
 assign n1952 = ( (~ n531) ) | ( n2512 ) ;
 assign n1953 = ( n2512 ) | ( n827 ) ;
 assign n1954 = ( (~ n531) ) | ( n1915 ) ;
 assign n1955 = ( n626 ) | ( n827 ) ;
 assign n1956 = ( (~ n531) ) | ( n619 ) ;
 assign n1957 = ( n2517 ) | ( n827 ) ;
 assign n1958 = ( n2433  &  n2441  &  n1079  &  n2412  &  n2399  &  n2392 ) ;
 assign n1951 = ( n1952  &  n1953  &  n1954  &  n1955  &  n1956  &  n1891  &  n1957  &  n1958 ) ;
 assign n1959 = ( n2517 ) | ( n891 ) ;
 assign n1960 = ( n388 ) | ( n574 ) ;
 assign n1961 = ( n626 ) | ( n891 ) ;
 assign n1962 = ( n891 ) | ( n619 ) ;
 assign n1963 = ( n1915 ) | ( n891 ) ;
 assign n1964 = ( n2512 ) | ( n388 ) ;
 assign n1965 = ( n366  &  n370  &  n381 ) ;
 assign n1966 = ( n1425  &  n524  &  n1456 ) ;
 assign n1967 = ( (~ n350)  &  (~ n692) ) ;
 assign n1970 = ( n441 ) | ( n173 ) ;
 assign n1971 = ( n441 ) | ( n177 ) ;
 assign n1972 = ( n441 ) | ( n1263 ) ;
 assign n1969 = ( n1970  &  n1971  &  n1972 ) ;
 assign n1973 = ( n441 ) | ( n178 ) ;
 assign n1974 = ( (~ n333) ) | ( n1239 ) ;
 assign n1975 = ( n441 ) | ( n1239 ) ;
 assign n1976 = ( n441 ) | ( n812 ) ;
 assign n1977 = ( n178 ) | ( (~ n333) ) ;
 assign n1978 = ( n441 ) | ( n1376 ) ;
 assign n1979 = ( (~ n333) ) | ( n1263 ) ;
 assign n1980 = ( (~ n333) ) | ( n812 ) ;
 assign n1981 = ( (~ n333) ) | ( n1236 ) ;
 assign n1982 = ( n441 ) | ( n1377 ) ;
 assign n1983 = ( n441 ) | ( n517 ) ;
 assign n1985 = ( (~ n333) ) | ( n1127 ) ;
 assign n1986 = ( n441 ) | ( n657 ) ;
 assign n1987 = ( (~ n333) ) | ( n499 ) ;
 assign n1988 = ( n441 ) | ( n1346 ) ;
 assign n1989 = ( (~ n333) ) | ( n1346 ) ;
 assign n1990 = ( n441 ) | ( n1341 ) ;
 assign n1984 = ( n1985  &  n1986  &  n1987  &  n1988  &  n1989  &  n1990 ) ;
 assign n1991 = ( n441 ) | ( n1324 ) ;
 assign n1992 = ( (~ n333) ) | ( n1341 ) ;
 assign n1993 = ( (~ n333) ) | ( n646 ) ;
 assign n1994 = ( (~ n333) ) | ( n1329 ) ;
 assign n1995 = ( (~ n333) ) | ( n1327 ) ;
 assign n1996 = ( (~ n333) ) | ( n1322 ) ;
 assign n1997 = ( n441 ) | ( n1033 ) ;
 assign n1998 = ( (~ n333) ) | ( n1454 ) ;
 assign n1999 = ( n441 ) | ( n1456 ) ;
 assign n2000 = ( (~ n333) ) | ( n1324 ) ;
 assign n2001 = ( n441 ) | ( n499 ) ;
 assign n2002 = ( n441 ) | ( n1329 ) ;
 assign n2004 = ( n1347 ) | ( n701 ) ;
 assign n2003 = ( n2004  &  n263 ) | ( n2004  &  n1347 ) ;
 assign n2005 = ( n427 ) | ( n1456 ) ;
 assign n2006 = ( n1347 ) | ( n1277 ) ;
 assign n2007 = ( n164 ) | ( n749 ) ;
 assign n2008 = ( n374 ) | ( n1376 ) ;
 assign n2009 = ( n374 ) | ( n1377 ) ;
 assign n2010 = ( n313 ) | ( n176 ) ;
 assign n2011 = ( n313 ) | ( n1267 ) ;
 assign n2012 = ( (~ n401) ) | ( n1346 ) ;
 assign n2013 = ( (~ n401) ) | ( n1033 ) ;
 assign n2014 = ( (~ n401) ) | ( n1324 ) ;
 assign n2015 = ( (~ n401) ) | ( n1329 ) ;
 assign n2016 = ( n313 ) | ( n1346 ) ;
 assign n2017 = ( n313 ) | ( n1033 ) ;
 assign n2018 = ( n441 ) | ( n1425 ) ;
 assign n2019 = ( (~ n333) ) | ( n1339 ) ;
 assign n2021 = ( (~ n333) ) | ( n1313 ) ;
 assign n2022 = ( n165 ) | ( (~ n333) ) ;
 assign n2023 = ( n441 ) | ( n458 ) ;
 assign n2024 = ( n164 ) | ( n173 ) ;
 assign n2025 = ( (~ n855) ) | ( n1239 ) ;
 assign n2026 = ( n164 ) | ( n308 ) ;
 assign n2027 = ( n164 ) | ( n517 ) ;
 assign n2028 = ( n164 ) | ( n1376 ) ;
 assign n2029 = ( n164 ) | ( n1377 ) ;
 assign n2030 = ( (~ n855) ) | ( n1236 ) ;
 assign n2031 = ( (~ n855) ) | ( n1248 ) ;
 assign n2032 = ( n177 ) | ( (~ n855) ) ;
 assign n2033 = ( n178 ) | ( (~ n855) ) ;
 assign n2034 = ( (~ n160) ) | ( n750 ) ;
 assign n2035 = ( (~ n160) ) | ( n1328 ) ;
 assign n2036 = ( (~ n160) ) | ( n1340 ) ;
 assign n2037 = ( n427 ) | ( n1247 ) ;
 assign n2038 = ( (~ n160) ) | ( n185 ) ;
 assign n2039 = ( (~ n160) ) | ( n1264 ) ;
 assign n2040 = ( n427 ) | ( n1470 ) ;
 assign n2041 = ( (~ n160) ) | ( n1318 ) ;
 assign n2042 = ( (~ n160) ) | ( n520 ) ;
 assign n2043 = ( (~ n160) ) | ( n1206 ) ;
 assign n2044 = ( n427 ) | ( n520 ) ;
 assign n2046 = ( n441 ) | ( n1264 ) ;
 assign n2047 = ( n441 ) | ( n1345 ) ;
 assign n2048 = ( (~ n333) ) | ( n1264 ) ;
 assign n2045 = ( n2046  &  n2047  &  n2048 ) ;
 assign n2049 = ( n441 ) | ( n1340 ) ;
 assign n2050 = ( n185 ) | ( (~ n333) ) ;
 assign n2051 = ( (~ n333) ) | ( n1318 ) ;
 assign n2052 = ( (~ n333) ) | ( n1330 ) ;
 assign n2053 = ( (~ n333) ) | ( n1328 ) ;
 assign n2054 = ( (~ n333) ) | ( n1345 ) ;
 assign n2055 = ( n441 ) | ( n1247 ) ;
 assign n2056 = ( n441 ) | ( n185 ) ;
 assign n2057 = ( n441 ) | ( n1318 ) ;
 assign n2058 = ( n441 ) | ( n1470 ) ;
 assign n2059 = ( (~ n333) ) | ( n1247 ) ;
 assign n2061 = ( (~ n333) ) | ( n1066 ) ;
 assign n2062 = ( (~ n333) ) | ( n811 ) ;
 assign n2063 = ( (~ n333) ) | ( n1237 ) ;
 assign n2064 = ( n441 ) | ( n265 ) ;
 assign n2065 = ( n265 ) | ( (~ n333) ) ;
 assign n2066 = ( n441 ) | ( n266 ) ;
 assign n2060 = ( n2061  &  n2062  &  n2063  &  n2064  &  n2065  &  n2066 ) ;
 assign n2067 = ( (~ n333) ) | ( n1241 ) ;
 assign n2068 = ( (~ n333) ) | ( n1242 ) ;
 assign n2069 = ( n441 ) | ( n811 ) ;
 assign n2070 = ( n441 ) | ( n1397 ) ;
 assign n2071 = ( n441 ) | ( n537 ) ;
 assign n2072 = ( (~ n333) ) | ( n1233 ) ;
 assign n2073 = ( n266 ) | ( (~ n333) ) ;
 assign n2074 = ( (~ n333) ) | ( n1397 ) ;
 assign n2076 = ( n374 ) | ( n520 ) ;
 assign n2075 = ( n2076  &  n713  &  n1806 ) ;
 assign n2077 = ( n184 ) | ( n520 ) ;
 assign n2078 = ( n1749  &  n600  &  n1673  &  n1712  &  n586  &  n596 ) ;
 assign n2080 = ( (~ n855) ) | ( n1219 ) ;
 assign n2079 = ( n1686  &  n1674  &  n1687  &  n1690  &  n2080  &  n2078 ) ;
 assign n2081 = ( (~ n692)  &  n1902 ) | ( n1247  &  n1264  &  n1902 ) ;
 assign n2082 = ( (~ n160)  &  (~ n848) ) | ( (~ n160)  &  n1469 ) | ( (~ n848)  &  n1470 ) | ( n1469  &  n1470 ) ;
 assign n2083 = ( (~ n401)  &  n2082 ) | ( n750  &  n2082 ) ;
 assign n2084 = ( (~ n160) ) | ( n1345 ) ;
 assign n2085 = ( (~ n160) ) | ( n1127 ) ;
 assign n2086 = ( (~ n160) ) | ( n499 ) ;
 assign n2087 = ( (~ n160) ) | ( n1327 ) ;
 assign n2088 = ( n427 ) | ( n499 ) ;
 assign n2090 = ( n374 ) | ( n1454 ) ;
 assign n2089 = ( n1777  &  n1741  &  n2090  &  n739  &  n1729  &  n1824 ) ;
 assign n2092 = ( (~ n333) ) | ( n1455 ) ;
 assign n2091 = ( n1707  &  n1701  &  n2092 ) ;
 assign n2093 = ( n1924  &  n1899  &  n1694  &  n1709  &  n1688  &  n1757 ) ;
 assign n2094 = ( (~ n160) ) | ( n1346 ) ;
 assign n2095 = ( n263  &  (~ n848) ) | ( n263  &  n1454 ) | ( (~ n848)  &  n1455 ) | ( n1454  &  n1455 ) ;
 assign n2097 = ( (~ n160)  &  n313 ) | ( (~ n160)  &  n1322 ) | ( n313  &  n1456 ) | ( n1322  &  n1456 ) ;
 assign n2098 = ( n164 ) | ( n1424 ) ;
 assign n2099 = ( (~ n160) ) | ( n1334 ) ;
 assign n2100 = ( (~ n160) ) | ( n1339 ) ;
 assign n2101 = ( n427 ) | ( n1423 ) ;
 assign n2102 = ( n313 ) | ( n1313 ) ;
 assign n2103 = ( n313 ) | ( n307 ) ;
 assign n2104 = ( (~ n401) ) | ( n1313 ) ;
 assign n2105 = ( n313 ) | ( n1323 ) ;
 assign n2106 = ( n313 ) | ( n1339 ) ;
 assign n2107 = ( (~ n401) ) | ( n1319 ) ;
 assign n2108 = ( n581  &  n1725  &  n1714 ) ;
 assign n2110 = ( n184 ) | ( n1334 ) ;
 assign n2111 = ( n184 ) | ( n172 ) ;
 assign n2112 = ( n313 ) | ( n172 ) ;
 assign n2109 = ( n737  &  n723  &  n1820  &  n2110  &  n2111  &  n2112  &  n595  &  n2108 ) ;
 assign n2113 = ( n1797  &  n1800  &  n709  &  n1791  &  n1805 ) ;
 assign n2114 = ( n184 ) | ( n1423 ) ;
 assign n2115 = ( n184 ) | ( n1313 ) ;
 assign n2116 = ( (~ n794)  &  n1907 ) | ( n1342  &  n1424  &  n1907 ) ;
 assign n2117 = ( (~ n692)  &  n1426 ) | ( n1339  &  n1344  &  n1426 ) ;
 assign n2118 = ( (~ n160) ) | ( n1344 ) ;
 assign n2119 = ( (~ n160) ) | ( n1128 ) ;
 assign n2120 = ( (~ n160) ) | ( n266 ) ;
 assign n2121 = ( n427 ) | ( n511 ) ;
 assign n2122 = ( n313 ) | ( n1241 ) ;
 assign n2123 = ( (~ n401) ) | ( n811 ) ;
 assign n2124 = ( (~ n401) ) | ( n1237 ) ;
 assign n2125 = ( n313 ) | ( n1242 ) ;
 assign n2126 = ( n313 ) | ( n266 ) ;
 assign n2127 = ( n441 ) | ( n1396 ) ;
 assign n2128 = ( n164 ) | ( n179 ) ;
 assign n2129 = ( n374 ) | ( n537 ) ;
 assign n2131 = ( n184 ) | ( n511 ) ;
 assign n2130 = ( n584  &  n1731  &  n1696  &  n2131 ) ;
 assign n2132 = ( n184 ) | ( n1128 ) ;
 assign n2133 = ( n374 ) | ( n511 ) ;
 assign n2134 = ( n1756  &  n1708  &  n1685  &  n1672 ) ;
 assign n2135 = ( n264  &  n1265 ) | ( (~ n692)  &  n1265 ) | ( n264  &  n1397 ) | ( (~ n692)  &  n1397 ) ;
 assign n2136 = ( (~ n143)  &  n263 ) | ( n263  &  n811 ) | ( (~ n143)  &  n1396 ) | ( n811  &  n1396 ) ;
 assign n2137 = ( n313  &  (~ n855) ) | ( n313  &  n1233 ) | ( (~ n855)  &  n1237 ) | ( n1233  &  n1237 ) ;
 assign n2138 = ( (~ n160) ) | ( n1267 ) ;
 assign n2139 = ( n427 ) | ( n812 ) ;
 assign n2140 = ( (~ n160) ) | ( n1236 ) ;
 assign n2141 = ( (~ n401) ) | ( n1236 ) ;
 assign n2142 = ( n313 ) | ( n308 ) ;
 assign n2143 = ( n313 ) | ( n812 ) ;
 assign n2144 = ( n178 ) | ( (~ n401) ) ;
 assign n2145 = ( n1821  &  n736  &  n1743  &  n1713  &  n577  &  n754 ) ;
 assign n2147 = ( n184 ) | ( n1235 ) ;
 assign n2148 = ( n173 ) | ( n184 ) ;
 assign n2149 = ( n374 ) | ( n1236 ) ;
 assign n2146 = ( n2147  &  n2148  &  n2149  &  n1798  &  n1799 ) ;
 assign n2151 = ( n1229 ) | ( n184 ) ;
 assign n2152 = ( n374 ) | ( n1248 ) ;
 assign n2150 = ( n1788  &  n1790  &  n2151  &  n711  &  n710  &  n2152 ) ;
 assign n2153 = ( n184 ) | ( n1248 ) ;
 assign n2155 = ( (~ n223)  &  (~ n392) ) ;
 assign n2156 = ( n388  &  n827 ) ;
 assign n2154 = ( n2155  &  n2156 ) | ( n1235  &  n2156 ) | ( n2155  &  n1267 ) | ( n1235  &  n1267 ) ;
 assign n2158 = ( (~ n401)  &  (~ n531) ) ;
 assign n2157 = ( n2154  &  n2158 ) | ( n2154  &  n812 ) ;
 assign n2159 = ( (~ n160)  &  n184 ) | ( (~ n160)  &  n517 ) | ( n184  &  n1377 ) | ( n517  &  n1377 ) ;
 assign n2160 = ( n1343 ) | ( n827 ) ;
 assign n2161 = ( (~ n531) ) | ( n1343 ) ;
 assign n2162 = ( n388 ) | ( n1320 ) ;
 assign n2163 = ( n388 ) | ( n220 ) ;
 assign n2164 = ( n219 ) | ( n891 ) ;
 assign n2165 = ( n1512 ) | ( n891 ) ;
 assign n2166 = ( n443  &  n1669  &  n446 ) ;
 assign n2168 = ( (~ n401) ) | ( n1320 ) ;
 assign n2169 = ( n313 ) | ( n1320 ) ;
 assign n2167 = ( n782  &  n1835  &  n53  &  n2168  &  n2169  &  n714  &  n1781  &  n385 ) ;
 assign n2170 = ( (~ n333) ) | ( n1312 ) ;
 assign n2171 = ( (~ n151) ) | ( n1966 ) ;
 assign n2172 = ( (~ n855) ) | ( n1520 ) ;
 assign n2173 = ( n427  &  n1279 ) ;
 assign n2177 = ( n263  &  n1270 ) ;
 assign n2178 = ( (~ n692)  &  n1279 ) ;
 assign n2176 = ( n2177  &  n2178 ) | ( n1314  &  n2178 ) | ( n2177  &  n1342 ) | ( n1314  &  n1342 ) ;
 assign n2179 = ( (~ n151)  &  n1276 ) ;
 assign n2182 = ( n164  &  (~ n531)  &  (~ n1140)  &  n1283 ) ;
 assign n2181 = ( n165  &  n1320 ) | ( (~ n350)  &  n1320 ) | ( n165  &  n2182 ) | ( (~ n350)  &  n2182 ) ;
 assign n2183 = ( n219  &  n277 ) | ( n277  &  n374 ) | ( n219  &  (~ n392) ) | ( n374  &  (~ n392) ) ;
 assign n2184 = ( n1279  &  n1270 ) | ( n1329  &  n1270 ) | ( n1279  &  n1347 ) | ( n1329  &  n1347 ) ;
 assign n2186 = ( (~ n401) ) | ( n749 ) ;
 assign n2185 = ( n1369  &  n1090  &  n1357  &  n661  &  n214  &  n1348  &  n218  &  n2186 ) ;
 assign n2189 = ( n572 ) | ( n827 ) ;
 assign n2190 = ( (~ n531) ) | ( n762 ) ;
 assign n2191 = ( n762 ) | ( n827 ) ;
 assign n2192 = ( n1514 ) | ( n827 ) ;
 assign n2193 = ( (~ n156) ) | ( n827 ) ;
 assign n2194 = ( n1227 ) | ( n827 ) ;
 assign n2196 = ( n180 ) | ( n938 ) ;
 assign n2195 = ( n181  &  n938 ) ;
 assign n2197 = ( n1227 ) | ( n388 ) ;
 assign n2198 = ( n388 ) | ( n572 ) ;
 assign n2199 = ( n319 ) | ( n388 ) ;
 assign n2200 = ( (~ n156) ) | ( n891 ) ;
 assign n2201 = ( n1514 ) | ( n891 ) ;
 assign n2203 = ( (~ n333) ) | ( n1064 ) ;
 assign n2202 = ( n1722  &  n2203  &  n1720 ) ;
 assign n2205 = ( (~ n151) ) | ( n1937 ) ;
 assign n2206 = ( (~ n401) ) | ( n1227 ) ;
 assign n2204 = ( n2205  &  n783  &  n1837  &  n52  &  n2206  &  n1803  &  n715  &  n1786 ) ;
 assign n2207 = ( (~ n855) ) | ( n1227 ) ;
 assign n2209 = ( n188  &  n2179 ) | ( n1226  &  n2179 ) | ( n188  &  n1257 ) | ( n1226  &  n1257 ) ;
 assign n2211 = ( n175  &  n1237 ) | ( (~ n229)  &  n1237 ) | ( n175  &  n2173 ) | ( (~ n229)  &  n2173 ) ;
 assign n2212 = ( (~ n198)  &  n1227 ) | ( n658  &  n1227 ) | ( (~ n198)  &  n2182 ) | ( n658  &  n2182 ) ;
 assign n2213 = ( (~ n350)  &  n1070 ) | ( n1070  &  n1236 ) | ( (~ n350)  &  n1271 ) | ( n1236  &  n1271 ) ;
 assign n2214 = ( (~ n156)  &  n179 ) | ( n179  &  n374 ) | ( (~ n156)  &  n1270 ) | ( n374  &  n1270 ) ;
 assign n2216 = ( (~ n160)  &  n1284 ) | ( n1229  &  n1284 ) ;
 assign n2217 = ( n1303  &  n55  &  n1296  &  n1291 ) ;
 assign n2218 = ( (~ n27)  &  n738  &  n1858  &  n1863 ) ;
 assign n2219 = ( (~ n344)  &  n2173 ) | ( (~ n344)  &  n1324  &  n1507 ) ;
 assign n2221 = ( (~ n229)  &  (~ n348) ) | ( (~ n348)  &  n651  &  n1508 ) ;
 assign n2223 = ( (~ n143)  &  (~ n351) ) | ( n315  &  (~ n351)  &  n1509 ) ;
 assign n2225 = ( (~ n354)  &  (~ n855) ) | ( n165  &  (~ n354)  &  (~ n922) ) ;
 assign n2228 = ( (~ n1140)  &  n1510 ) ;
 assign n2227 = ( n342  &  n1704 ) | ( n164  &  n1704 ) | ( n342  &  n2228 ) | ( n164  &  n2228 ) ;
 assign n2229 = ( (~ n143) ) | ( n335 ) ;
 assign n2230 = ( n171  &  n339 ) | ( n171  &  n427 ) | ( n339  &  (~ n692) ) | ( n427  &  (~ n692) ) ;
 assign n2231 = ( (~ n531)  &  n1771 ) | ( n883  &  n1771 ) | ( (~ n531)  &  n2155 ) | ( n883  &  n2155 ) ;
 assign n2233 = ( (~ n160)  &  n388 ) ;
 assign n2232 = ( n658  &  n1270 ) | ( n2233  &  n1270 ) | ( n658  &  n1081 ) | ( n2233  &  n1081 ) ;
 assign n2235 = ( (~ n223)  &  n1516 ) ;
 assign n2234 = ( n1279  &  n341 ) | ( n1508  &  n341 ) | ( n1279  &  n2235 ) | ( n1508  &  n2235 ) ;
 assign n2237 = ( (~ n223)  &  (~ n482) ) ;
 assign n2236 = ( n174  &  n168 ) | ( n168  &  (~ n401) ) | ( n174  &  n2237 ) | ( (~ n401)  &  n2237 ) ;
 assign n2239 = ( n164  &  n1516  &  n1517 ) ;
 assign n2240 = ( n427  &  n1517  &  n1519 ) ;
 assign n2238 = ( n1705  &  n1666 ) | ( n2239  &  n1666 ) | ( n1705  &  n2240 ) | ( n2239  &  n2240 ) ;
 assign n2242 = ( (~ n151)  &  (~ n975) ) ;
 assign n2241 = ( n1343  &  n1583 ) | ( n2242  &  n1583 ) | ( n1343  &  n1326 ) | ( n2242  &  n1326 ) ;
 assign n2243 = ( n765 ) | ( n2319 ) ;
 assign n2244 = ( (~ n223)  &  (~ n848) ) | ( n749  &  (~ n848) ) | ( (~ n223)  &  n1262 ) | ( n749  &  n1262 ) ;
 assign n2245 = ( (~ n14)  &  n1272 ) | ( n517  &  n1272 ) | ( (~ n14)  &  n1342 ) | ( n517  &  n1342 ) ;
 assign n2246 = ( n297  &  n538  &  n525  &  n1554  &  n394  &  n1537  &  n1534  &  n1117 ) ;
 assign n2247 = ( n2511 ) | ( n827 ) ;
 assign n2248 = ( (~ n531) ) | ( n810 ) ;
 assign n2249 = ( n810 ) | ( n827 ) ;
 assign n2250 = ( n453 ) | ( n938 ) ;
 assign n2251 = ( n441 ) | ( n748 ) ;
 assign n2252 = ( n1908 ) | ( n427 ) ;
 assign n2254 = ( (~ n333) ) | ( n1586 ) ;
 assign n2255 = ( (~ n333) ) | ( n781 ) ;
 assign n2256 = ( (~ n333) ) | ( n634 ) ;
 assign n2257 = ( (~ n333) ) | ( n630 ) ;
 assign n2258 = ( (~ n333) ) | ( n645 ) ;
 assign n2259 = ( n441 ) | ( n638 ) ;
 assign n2261 = ( (~ n333) ) | ( n1585 ) ;
 assign n2260 = ( (~ n793)  &  n2261 ) | ( (~ n794)  &  n1277  &  n2261 ) ;
 assign n2262 = ( n1604  &  n2242 ) | ( n1588  &  n2242 ) | ( n1604  &  n781 ) | ( n1588  &  n781 ) ;
 assign n2265 = ( n891  &  n827 ) ;
 assign n2266 = ( (~ n223)  &  (~ n333)  &  n388 ) ;
 assign n2268 = ( n2265 ) | ( n173 ) ;
 assign n2269 = ( (~ n143)  &  n1277 ) | ( n812  &  n1277 ) | ( (~ n143)  &  n1377 ) | ( n812  &  n1377 ) ;
 assign n2270 = ( n1336  &  n1259 ) ;
 assign n2272 = ( (~ n794)  &  n1510 ) ;
 assign n2271 = ( (~ n140)  &  n2272 ) | ( (~ n140)  &  n1377  &  n1425 ) ;
 assign n2273 = ( n466  &  (~ n473) ) | ( n164  &  (~ n473)  &  n1598 ) ;
 assign n2275 = ( (~ n476)  &  n718 ) | ( n374  &  (~ n476)  &  n1599 ) ;
 assign n2278 = ( (~ n692)  &  n1274 ) ;
 assign n2277 = ( n1965  &  n2278 ) | ( n464  &  n2278 ) | ( n1965  &  n469 ) | ( n464  &  n469 ) ;
 assign n2279 = ( n461  &  n465 ) | ( n461  &  (~ n1140) ) | ( n465  &  n1588 ) | ( (~ n1140)  &  n1588 ) ;
 assign n2283 = ( (~ n794)  &  n1276 ) ;
 assign n2285 = ( (~ n482)  &  n827 ) ;
 assign n2284 = ( n2285  &  n2265 ) | ( n1236  &  n2265 ) | ( n2285  &  n812 ) | ( n1236  &  n812 ) ;
 assign n2287 = ( n780  &  n1603 ) ;
 assign n2286 = ( n1923  &  n2287 ) | ( n998  &  n2287 ) | ( n1923  &  n1344 ) | ( n998  &  n1344 ) ;
 assign n2288 = ( n2284  &  n2286  &  n1280 ) | ( n2284  &  n2286  &  n1267 ) ;
 assign n2290 = ( n1279  &  n1604 ) ;
 assign n2289 = ( (~ n347)  &  n1263 ) | ( n381  &  n1263 ) | ( (~ n347)  &  n2290 ) | ( n381  &  n2290 ) ;
 assign n2292 = ( n827  &  n462  &  n1280 ) ;
 assign n2291 = ( (~ n229)  &  n1339 ) | ( n459  &  n1339 ) | ( (~ n229)  &  n2292 ) | ( n459  &  n2292 ) ;
 assign n2293 = ( (~ n356)  &  n434 ) | ( n434  &  n1516 ) | ( (~ n356)  &  n1519 ) | ( n1516  &  n1519 ) ;
 assign n2294 = ( n184  &  n458 ) | ( n370  &  n458 ) | ( n184  &  (~ n692) ) | ( n370  &  (~ n692) ) ;
 assign n2295 = ( (~ n333)  &  n780 ) | ( n590  &  n780 ) | ( (~ n333)  &  n781 ) | ( n590  &  n781 ) ;
 assign n2296 = ( n467  &  (~ n531)  &  n2295 ) | ( n467  &  n1248  &  n2295 ) ;
 assign n2297 = ( n414  &  n1627  &  n447  &  n56  &  n1089  &  n1612  &  n1609  &  n1607 ) ;
 assign n2298 = ( n365  &  n369  &  n373  &  n377  &  n380  &  n384  &  n393  &  n403 ) ;
 assign n2299 = ( n1503  &  n427 ) | ( n1503  &  n1507  &  n1396 ) ;
 assign n2301 = ( n524  &  n1246 ) | ( (~ n541)  &  n1246 ) | ( n524  &  n2233 ) | ( (~ n541)  &  n2233 ) ;
 assign n2302 = ( (~ n848)  &  n1345 ) | ( n1264  &  n1345 ) | ( (~ n848)  &  n2242 ) | ( n1264  &  n2242 ) ;
 assign n2303 = ( (~ n143) ) | ( n1330 ) ;
 assign n2304 = ( n1337  &  n1279 ) | ( n1337  &  n1507  &  n1469 ) ;
 assign n2305 = ( n2304  &  n184 ) | ( n2304  &  n658  &  n1066 ) ;
 assign n2306 = ( n170  &  n1603 ) | ( n2237  &  n1603 ) | ( n170  &  n750 ) | ( n2237  &  n750 ) ;
 assign n2308 = ( n192  &  n1643 ) ;
 assign n2307 = ( n2308  &  n2228 ) | ( n308  &  n2228 ) | ( n2308  &  n1256 ) | ( n308  &  n1256 ) ;
 assign n2309 = ( n173  &  (~ n486) ) | ( (~ n486)  &  n1582 ) | ( n173  &  n1640 ) | ( n1582  &  n1640 ) ;
 assign n2311 = ( (~ n855)  &  n1318 ) | ( n1318  &  n1509 ) | ( (~ n855)  &  n2178 ) | ( n1509  &  n2178 ) ;
 assign n2312 = ( (~ n392)  &  n1396 ) | ( n1214  &  n1396 ) | ( (~ n392)  &  n2235 ) | ( n1214  &  n2235 ) ;
 assign n2314 = ( n427  &  n701  &  n1516 ) ;
 assign n2313 = ( n2311  &  n2312  &  n2314 ) | ( n2311  &  n2312  &  n1376 ) ;
 assign n2315 = ( n1643  &  n2239 ) | ( n1239  &  n2239 ) | ( n1643  &  n187 ) | ( n1239  &  n187 ) ;
 assign n2316 = ( n2287  &  n2240 ) | ( n1345  &  n2240 ) | ( n2287  &  n572 ) | ( n1345  &  n572 ) ;
 assign n2317 = ( n1205 ) | ( n1268 ) ;
 assign n2319 = ( (~ n333)  &  n427  &  (~ n692)  &  n780  &  (~ n975) ) ;
 assign n2318 = ( (~ n922)  &  n1070 ) | ( n1070  &  n1265 ) | ( (~ n922)  &  n2319 ) | ( n1265  &  n2319 ) ;
 assign n2320 = ( n2272  &  n1270 ) | ( n524  &  n1270 ) | ( n2272  &  n1937 ) | ( n524  &  n1937 ) ;
 assign n2322 = ( (~ n333) ) | ( n656 ) ;
 assign n2323 = ( n2508 ) | ( n441 ) ;
 assign n2324 = ( n656 ) | ( n441 ) ;
 assign n2325 = ( (~ n333) ) | ( n1745 ) ;
 assign n2326 = ( n612 ) | ( n441 ) ;
 assign n2327 = ( n441 ) | ( n807 ) ;
 assign n2328 = ( n606  &  n615  &  n1717  &  n668  &  n536  &  n522  &  n447  &  n421 ) ;
 assign n2329 = ( (~ n160) ) | ( n649 ) ;
 assign n2330 = ( n427 ) | ( n574 ) ;
 assign n2331 = ( n622 ) | ( n427 ) ;
 assign n2332 = ( n1745 ) | ( n427 ) ;
 assign n2333 = ( n2508 ) | ( n427 ) ;
 assign n2334 = ( n650  &  n1627  &  n1680  &  n289  &  n1439  &  n1554 ) ;
 assign n2336 = ( n1264  &  n265 ) ;
 assign n2337 = ( n1069 ) | ( n313 ) ;
 assign n2338 = ( n313 ) | ( n617 ) ;
 assign n2340 = ( (~ n401) ) | ( n1770 ) ;
 assign n2341 = ( (~ n392)  &  (~ n401) ) | ( (~ n392)  &  n758 ) | ( (~ n401)  &  n763 ) | ( n758  &  n763 ) ;
 assign n2342 = ( (~ n57)  &  n214 ) | ( n212  &  n214 ) ;
 assign n2343 = ( n626 ) | ( n184 ) ;
 assign n2344 = ( n1472  &  n322  &  n2129  &  n1436  &  n2009  &  n1475  &  n2008  &  n1435 ) ;
 assign n2345 = ( n2358 ) | ( n374 ) ;
 assign n2347 = ( n1745 ) | ( n374 ) ;
 assign n2348 = ( n2512 ) | ( n374 ) ;
 assign n2349 = ( n622 ) | ( n374 ) ;
 assign n2351 = ( (~ n237) ) | ( n771 ) ;
 assign n2352 = ( (~ n350) ) | ( n1747 ) ;
 assign n2353 = ( n2099  &  n2119 ) ;
 assign n2354 = ( n844 ) | ( (~ n855) ) ;
 assign n2355 = ( n619  &  n2087 ) | ( (~ n347)  &  (~ n855)  &  n2087 ) ;
 assign n2356 = ( n2358 ) | ( n891 ) ;
 assign n2358 = ( n748  &  n1064  &  n1312 ) ;
 assign n2357 = ( (~ n347)  &  (~ n855) ) | ( n748  &  (~ n855) ) | ( (~ n347)  &  n2358 ) | ( n748  &  n2358 ) ;
 assign n2359 = ( n1481  &  n1535  &  n2141  &  n2107  &  n2144  &  n2322  &  n1542  &  n1977 ) ;
 assign n2360 = ( n1555  &  n2140  &  n1351  &  n2207  &  n1457  &  n1399  &  n1624  &  n816 ) ;
 assign n2361 = ( n1404  &  n2080  &  n2030  &  n1430  &  n2033  &  n1961  &  n2165  &  n2201 ) ;
 assign n2362 = ( (~ n347)  &  n1265 ) ;
 assign n2363 = ( n181  &  (~ n732) ) ;
 assign n2364 = ( (~ n333)  &  (~ n855) ) | ( n574  &  (~ n855) ) | ( (~ n333)  &  n1512 ) | ( n574  &  n1512 ) ;
 assign n2366 = ( n1628  &  n1288 ) ;
 assign n2367 = ( n1529  &  n1774  &  n2324  &  n2125  &  n2330  &  n1973  &  n1353  &  n2366 ) ;
 assign n2368 = ( n2250  &  n1596  &  n2247 ) ;
 assign n2369 = ( n1960  &  n313 ) | ( n1960  &  n634 ) ;
 assign n2375 = ( (~ n160) ) | ( n863 ) ;
 assign n2374 = ( n752  &  n575  &  n1724  &  n1702  &  n652  &  n423  &  n1335  &  n2375 ) ;
 assign n2376 = ( n2055  &  n1976  &  n1975  &  n2333  &  n2049  &  n2066  &  n1990 ) ;
 assign n2377 = ( n216  &  n1527  &  n2122  &  n1526  &  n1381  &  n1597  &  n817 ) ;
 assign n2378 = ( n1558  &  n2139  &  n1551  &  n2024  &  n1964  &  n1466  &  n2198 ) ;
 assign n2379 = ( n1666  &  n441 ) | ( n374  &  n441 ) | ( n1666  &  n434 ) | ( n374  &  n434 ) ;
 assign n2380 = ( n433  &  n452 ) | ( n433  &  n938 ) ;
 assign n2381 = ( n1539  &  n1974  &  n2248  &  n2100  &  n2120  &  n2036 ) ;
 assign n2382 = ( n1465  &  n1411  &  n1980  &  n1557  &  n1445  &  n1464 ) ;
 assign n2383 = ( n1993  &  n2067  &  n2200  &  n1992  &  n1563  &  n2258  &  n2382 ) ;
 assign n2385 = ( n452  &  (~ n909) ) | ( n181  &  n451  &  (~ n909) ) ;
 assign n2387 = ( n2158  &  n1519 ) | ( n812  &  n1519 ) | ( n2158  &  n824 ) | ( n812  &  n824 ) ;
 assign n2388 = ( n2387  &  n1666 ) | ( n2387  &  n1598 ) ;
 assign n2389 = ( n315  &  n316 ) | ( n316  &  n891 ) | ( n315  &  (~ n1138) ) | ( n891  &  (~ n1138) ) ;
 assign n2390 = ( n2102  &  n1486  &  n1394  &  n2101  &  n2121  &  n1559 ) ;
 assign n2392 = ( n827 ) | ( n617 ) ;
 assign n2391 = ( n1957  &  n1285  &  n2392  &  n2196  &  n2338  &  n1253  &  n2390 ) ;
 assign n2393 = ( (~ n23)  &  n1388  &  n1402  &  n1458  &  n1548  &  n2337 ) ;
 assign n2395 = ( n1069 ) | ( n388 ) ;
 assign n2396 = ( n374  &  n313 ) | ( n590  &  n313 ) | ( n374  &  n381 ) | ( n590  &  n381 ) ;
 assign n2397 = ( n637  &  n380  &  n1717 ) ;
 assign n2398 = ( n1532  &  n1255  &  n1286 ) ;
 assign n2399 = ( n628 ) | ( n827 ) ;
 assign n2400 = ( n1614  &  n1309  &  n1372 ) ;
 assign n2401 = ( n2252  &  n1983  &  n2056  &  n1574  &  n2023  &  n2026  &  n2027  &  n2400 ) ;
 assign n2402 = ( n2057  &  n1498  &  n1592 ) ;
 assign n2403 = ( n937  &  n441 ) | ( n215  &  n441 ) | ( n937  &  n718 ) | ( n215  &  n718 ) ;
 assign n2404 = ( n1489  &  n1560  &  n1444  &  n1410  &  n1490  &  n2021  &  n2052 ) ;
 assign n2406 = ( (~ n855) ) | ( n1069 ) ;
 assign n2405 = ( n1521  &  n2086  &  n1173  &  n1385  &  n2406  &  n2042 ) ;
 assign n2407 = ( n1371  &  n1308  &  n1615  &  n2229 ) ;
 assign n2408 = ( (~ n140)  &  n617 ) | ( (~ n140)  &  n891  &  n1265 ) ;
 assign n2409 = ( (~ n531)  &  n2408 ) | ( n590  &  n707  &  n2408 ) ;
 assign n2410 = ( n638  &  n940 ) ;
 assign n2411 = ( n1543  &  n2061  &  n2050  &  n1487  &  n1985  &  n2051  &  n1254 ) ;
 assign n2412 = ( (~ n531) ) | ( n628 ) ;
 assign n2413 = ( n2041  &  n1384  &  n1441  &  n1383  &  n1406  &  n2085  &  n2254 ) ;
 assign n2414 = ( n1350  &  n1705 ) | ( (~ n531)  &  n891  &  n1350 ) ;
 assign n2415 = ( (~ n333)  &  (~ n950) ) | ( n917  &  (~ n950)  &  n1908 ) ;
 assign n2417 = ( n1519  &  n1515 ) | ( n1678  &  n1515 ) | ( n1519  &  n1397 ) | ( n1678  &  n1397 ) ;
 assign n2418 = ( (~ n143)  &  (~ n237) ) | ( (~ n237)  &  n513 ) | ( (~ n143)  &  n772 ) | ( n513  &  n772 ) ;
 assign n2419 = ( n1265  &  n1279 ) | ( n762  &  n1279 ) | ( n1265  &  n773 ) | ( n762  &  n773 ) ;
 assign n2420 = ( n340  &  n657 ) | ( n657  &  (~ n1138) ) | ( n340  &  n1516 ) | ( (~ n1138)  &  n1516 ) ;
 assign n2421 = ( n215 ) | ( n181 ) ;
 assign n2422 = ( n2410 ) | ( n313 ) ;
 assign n2423 = ( n520  &  n1423  &  n1330  &  n366  &  n177  &  n1248 ) ;
 assign n2424 = ( n638  &  n673  &  n811  &  n887  &  (~ n963)  &  n1915 ) ;
 assign n2425 = ( n2156  &  n164 ) | ( n619  &  n164 ) | ( n2156  &  n617 ) | ( n619  &  n617 ) ;
 assign n2426 = ( n622 ) | ( n388 ) ;
 assign n2427 = ( n1448  &  n1392  &  n1479  &  n1988  &  n2112  &  n2347 ) ;
 assign n2428 = ( n1972  &  n2046  &  n2332  &  n1971  &  n2064  &  n1540  &  n2047  &  n2427 ) ;
 assign n2429 = ( n2016  &  n1414  &  n2017  &  n1413  &  n1449  &  n1480 ) ;
 assign n2431 = ( n754  &  n2325  &  n1989  &  n2054  &  n1538  &  n2065  &  n2048  &  n1979 ) ;
 assign n2433 = ( (~ n531) ) | ( n622 ) ;
 assign n2432 = ( n1623  &  n868  &  n2013  &  n1416  &  n2161  &  n1301  &  n2433 ) ;
 assign n2436 = ( (~ n160)  &  (~ n732) ) | ( (~ n732)  &  n807 ) | ( (~ n160)  &  n1222 ) | ( n807  &  n1222 ) ;
 assign n2438 = ( n1710  &  n621  &  n1762  &  n1667  &  n423  &  n2436 ) ;
 assign n2439 = ( n2040  &  n1681  &  n1982  &  n2028  &  n2029  &  n1633 ) ;
 assign n2441 = ( n827 ) | ( (~ n1105) ) ;
 assign n2440 = ( n1541  &  n2326  &  n870  &  n1978  &  n1450  &  n1703  &  n2441  &  n2439 ) ;
 assign n2442 = ( n1573  &  n1497  &  n1306  &  n1567  &  n1999  &  n1590 ) ;
 assign n2446 = ( n996  &  n702 ) | ( n441  &  n702 ) | ( n996  &  n701 ) | ( n441  &  n701 ) ;
 assign n2448 = ( (~ n793)  &  n997  &  n1937 ) ;
 assign n2447 = ( n2448  &  n462 ) | ( n1277  &  n462 ) | ( n2448  &  n989 ) | ( n1277  &  n989 ) ;
 assign n2449 = ( n1291  &  n1357  &  n1068 ) | ( n1291  &  n1357  &  n827 ) ;
 assign n2450 = ( (~ n1051) ) | ( n1054 ) ;
 assign n2452 = ( (~ n90)  &  n1636 ) | ( (~ n1230)  &  n1636 ) | ( (~ n90)  &  n1950 ) | ( (~ n1230)  &  n1950 ) ;
 assign n2454 = ( n500  &  n1032 ) ;
 assign n2453 = ( n1178  &  n2454 ) | ( n37  &  n2454 ) | ( n1178  &  n1066 ) | ( n37  &  n1066 ) ;
 assign n2455 = ( n37  &  n265 ) | ( n265  &  (~ n1230) ) | ( n37  &  n2454 ) | ( (~ n1230)  &  n2454 ) ;
 assign n2456 = ( n37  &  n1346 ) | ( (~ n91)  &  n1346 ) | ( n37  &  n2454 ) | ( (~ n91)  &  n2454 ) ;
 assign n2458 = ( n1178  &  n1950 ) ;
 assign n2457 = ( (~ n76)  &  (~ n161) ) | ( (~ n76)  &  n1635 ) | ( (~ n76)  &  n2458 ) ;
 assign n2460 = ( n2080  &  n2406  &  n2098 ) ;
 assign n2461 = ( n325  &  n2128  &  n1067 ) | ( n325  &  n2128  &  n164 ) ;
 assign n2462 = ( n614  &  (~ n855) ) | ( (~ n848)  &  (~ n855) ) | ( n614  &  n1061 ) | ( (~ n848)  &  n1061 ) ;
 assign n2463 = ( (~ n482)  &  (~ n1103) ) | ( (~ n356)  &  (~ n1103)  &  n1936 ) ;
 assign n2465 = ( n2463  &  n1100 ) | ( n2463  &  n891 ) ;
 assign n2467 = ( n2242  &  n192 ) | ( n1346  &  n192 ) | ( n2242  &  n657 ) | ( n1346  &  n657 ) ;
 assign n2468 = ( (~ n1131)  &  n2272 ) | ( n537  &  (~ n1131)  &  n1456 ) ;
 assign n2472 = ( n1066  &  (~ n1143) ) | ( (~ n350)  &  (~ n1143)  &  n1510 ) ;
 assign n2474 = ( n1275  &  n2283 ) | ( n998  &  n2283 ) | ( n1275  &  n1058 ) | ( n998  &  n1058 ) ;
 assign n2475 = ( (~ n486)  &  n1599 ) | ( n1125  &  n1599 ) | ( (~ n486)  &  n1602 ) | ( n1125  &  n1602 ) ;
 assign n2476 = ( (~ n240)  &  n619 ) | ( (~ n240)  &  n1124 ) | ( n619  &  n1585 ) | ( n1124  &  n1585 ) ;
 assign n2478 = ( n649  &  (~ n848) ) | ( (~ n848)  &  n1269 ) | ( n649  &  n1601 ) | ( n1269  &  n1601 ) ;
 assign n2479 = ( (~ n1105)  &  n1454 ) | ( n1454  &  n1598 ) | ( (~ n1105)  &  n2285 ) | ( n1598  &  n2285 ) ;
 assign n2480 = ( n508  &  n749 ) | ( (~ n692)  &  n749 ) | ( n508  &  n1280 ) | ( (~ n692)  &  n1280 ) ;
 assign n2481 = ( n1923  &  n2287 ) | ( n608  &  n2287 ) | ( n1923  &  n1346 ) | ( n608  &  n1346 ) ;
 assign n2482 = ( n2290  &  n2242 ) | ( n265  &  n2242 ) | ( n2290  &  n807 ) | ( n265  &  n807 ) ;
 assign n2483 = ( n192  &  n626 ) | ( n1586  &  n626 ) | ( n192  &  n388 ) | ( n1586  &  n388 ) ;
 assign n2484 = ( (~ n350)  &  (~ n392) ) | ( n370  &  (~ n392) ) | ( (~ n350)  &  n630 ) | ( n370  &  n630 ) ;
 assign n2485 = ( n462  &  n1279 ) | ( n1587  &  n1279 ) | ( n462  &  n1220 ) | ( n1587  &  n1220 ) ;
 assign n2486 = ( n1516  &  n1270 ) | ( n657  &  n1270 ) | ( n1516  &  n1245 ) | ( n657  &  n1245 ) ;
 assign n2487 = ( (~ n14)  &  n427 ) | ( n427  &  n434 ) | ( (~ n14)  &  n634 ) | ( n434  &  n634 ) ;
 assign n2489 = ( n827 ) | ( n1127 ) ;
 assign n2488 = ( n543  &  n510  &  n414  &  n2489  &  n2487  &  n2486 ) ;
 assign n2490 = ( n1260  &  n1270 ) | ( n1260  &  n1966  &  n1246 ) ;
 assign n2491 = ( n458  &  n2490 ) | ( n164  &  (~ n392)  &  n2490 ) ;
 assign n2492 = ( n185  &  (~ n1154) ) | ( (~ n1154)  &  n1510  &  n1967 ) ;
 assign n2494 = ( (~ n14)  &  n169 ) | ( n169  &  n809 ) | ( (~ n14)  &  n2237 ) | ( n809  &  n2237 ) ;
 assign n2495 = ( n2494  &  n1511 ) | ( n2494  &  n2235 ) ;
 assign n2496 = ( n2308  &  n2228 ) | ( n307  &  n2228 ) | ( n2308  &  n1332 ) | ( n307  &  n1332 ) ;
 assign n2497 = ( (~ n1155)  &  (~ n1157)  &  n1219 ) | ( (~ n1155)  &  (~ n1157)  &  n2285 ) ;
 assign n2500 = ( n2314  &  n1643 ) | ( n1424  &  n1643 ) | ( n2314  &  n1323 ) | ( n1424  &  n1323 ) ;
 assign n2501 = ( n2239  &  n2290 ) | ( n1331  &  n2290 ) | ( n2239  &  n1264 ) | ( n1331  &  n1264 ) ;
 assign n2502 = ( n2240  &  n192 ) | ( n220  &  n192 ) | ( n2240  &  n172 ) | ( n220  &  n172 ) ;
 assign n2503 = ( n2319  &  n1325 ) | ( n1314  &  n1325 ) | ( n2319  &  n184 ) | ( n1314  &  n184 ) ;
 assign n2504 = ( (~ n486)  &  n1470 ) | ( n1206  &  n1470 ) | ( (~ n486)  &  n2272 ) | ( n1206  &  n2272 ) ;
 assign n2505 = ( (~ n350)  &  n1247 ) | ( n1247  &  n1318 ) | ( (~ n350)  &  n2292 ) | ( n1318  &  n2292 ) ;
 assign n2506 = ( n374  &  (~ n401) ) | ( (~ n401)  &  n657 ) | ( n374  &  n1127 ) | ( n657  &  n1127 ) ;
 assign n2507 = ( (~ i_0_) ) | ( i_1_ ) | ( i_2_ ) ;
 assign n2508 = ( n614  &  n1666 ) ;
 assign n2509 = ( n1219  &  n1220  &  n165 ) ;
 assign n2511 = ( n178  &  n1319  &  n370 ) ;
 assign n2512 = ( n645  &  n316 ) ;
 assign n2513 = ( n370  &  n1236  &  n165 ) ;
 assign n2514 = ( n1235  &  n1205 ) ;
 assign n2515 = ( n1334  &  n1326 ) ;
 assign n2516 = ( n1313  &  n431 ) ;
 assign n2517 = ( n638  &  n312 ) ;
 assign n2518 = ( (~ n922)  &  n1423 ) ;


endmodule

