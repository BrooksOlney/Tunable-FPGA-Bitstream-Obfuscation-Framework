module ex5p (
	i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, 
	o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, 
	o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, 
	o_20_, o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, 
	o_30_, o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, 
	o_40_, o_41_, o_42_, o_43_, o_44_, o_45_, o_46_, o_47_, o_48_, o_49_, 
	o_50_, o_51_, o_52_, o_53_, o_54_, o_55_, o_56_, o_57_, o_58_, o_59_, 
	o_60_, o_61_, o_62_);

input i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_;

output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_, o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_, o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_, o_41_, o_42_, o_43_, o_44_, o_45_, o_46_, o_47_, o_48_, o_49_, o_50_, o_51_, o_52_, o_53_, o_54_, o_55_, o_56_, o_57_, o_58_, o_59_, o_60_, o_61_, o_62_;

wire n2, n3, n1, n5, n6, n4, n8, n9, n7, n11, n12, n10, n14, n15, n13, n17, n18, n16, n20, n19, n23, n24, n22, n26, n25, n29, n30, n31, n32, n33, n28, n35, n36, n37, n38, n39, n40, n41, n42, n34, n44, n45, n46, n47, n48, n49, n50, n51, n43, n53, n54, n55, n56, n57, n58, n52, n60, n61, n62, n63, n64, n65, n66, n59, n68, n69, n70, n71, n72, n73, n74, n67, n76, n77, n78, n79, n80, n81, n82, n83, n75, n85, n86, n87, n88, n89, n84, n91, n92, n93, n94, n95, n90, n97, n98, n99, n100, n101, n96, n103, n104, n105, n106, n107, n102, n109, n108, n111, n112, n113, n114, n110, n116, n117, n118, n119, n120, n121, n115, n123, n124, n125, n126, n122, n128, n127, n130, n131, n132, n133, n129, n135, n136, n137, n134, n139, n140, n141, n142, n143, n138, n145, n144, n147, n148, n149, n150, n151, n152, n153, n146, n155, n156, n157, n158, n159, n160, n154, n162, n163, n164, n165, n161, n167, n168, n169, n170, n171, n172, n166, n174, n175, n176, n177, n173, n179, n180, n181, n182, n183, n178, n185, n186, n187, n188, n189, n190, n184, n192, n193, n194, n195, n196, n197, n191, n199, n200, n201, n198, n203, n204, n205, n202, n207, n208, n209, n206, n211, n212, n213, n210, n215, n216, n214, n218, n219, n220, n221, n217, n223, n222, n225, n226, n224, n228, n229, n230, n227, n232, n233, n234, n231, n237, n235, n242, n240, n241, n239, n245, n244, n243, n246, n248, n247, n250, n249, n251, n253, n254, n252, n257, n258, n256, n260, n259, n261, n262, n265, n266, n264, n267, n268, n272, n270, n273, n274, n275, n276, n279, n278, n277, n280, n281, n284, n285, n283, n282, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n297, n296, n298, n299, n301, n300, n303, n304, n302, n306, n305, n309, n310, n312, n316, n317, n319, n320, n321, n322, n323, n324, n325, n327, n328, n329, n331, n332, n333, n334, n330, n335, n337, n336, n339, n340, n342, n341, n343, n344, n345, n346, n347, n348, n349, n351, n350, n353, n352, n355, n356, n357, n354, n359, n358, n361, n360, n362, n364, n365, n363, n366, n368, n367, n369, n371, n370, n372, n373, n374, n376, n375, n377, n380, n381, n379, n383, n384, n382, n386, n385, n388, n387, n390, n389, n391, n392, n393, n395, n396, n394, n397, n398, n399, n400, n401, n402, n403, n404, n405, n408, n406, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n422, n421, n423, n425, n424, n426, n428, n429, n427, n430, n432, n433, n431, n434, n436, n435, n437, n438, n440, n441, n439, n442, n443, n445, n446, n447, n444, n448, n449, n450, n451, n452, n454, n453, n455, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485;

assign o_0_ = ( (~ n231) ) ;
 assign o_1_ = ( (~ n227) ) ;
 assign o_2_ = ( (~ n278) ) ;
 assign o_3_ = ( (~ n241) ) ;
 assign o_4_ = ( (~ n334) ) ;
 assign o_5_ = ( (~ n224) ) ;
 assign o_6_ = ( (~ n1) ) ;
 assign o_7_ = ( (~ n50) ) ;
 assign o_8_ = ( (~ n335) ) ;
 assign o_9_ = ( (~ n376) ) ;
 assign o_10_ = ( (~ n4) ) ;
 assign o_11_ = ( (~ n49) ) ;
 assign o_12_ = ( (~ n258) ) ;
 assign o_13_ = ( (~ n356) ) ;
 assign o_14_ = ( (~ n392) ) ;
 assign o_15_ = ( (~ n6) ) ;
 assign o_16_ = ( (~ n284) ) ;
 assign o_17_ = ( (~ n222) ) ;
 assign o_18_ = ( (~ n297) ) ;
 assign o_19_ = ( (~ n295) ) ;
 assign o_20_ = ( (~ n7) ) ;
 assign o_21_ = ( (~ n10) ) ;
 assign o_22_ = ( (~ n13) ) ;
 assign o_23_ = ( (~ n217) ) ;
 assign o_24_ = ( (~ n390) ) ;
 assign o_25_ = ( (~ n70) ) ;
 assign o_26_ = ( (~ n16) ) ;
 assign o_27_ = ( (~ n130) ) ;
 assign o_28_ = ( (~ n443) ) ;
 assign o_29_ = ( (~ n391) ) ;
 assign o_30_ = ( (~ n18) ) ;
 assign o_31_ = ( (~ n214) ) ;
 assign o_32_ = ( (~ n210) ) ;
 assign o_33_ = ( (~ n206) ) ;
 assign o_34_ = ( (~ n202) ) ;
 assign o_35_ = ( (~ n198) ) ;
 assign o_36_ = ( (~ n191) ) ;
 assign o_37_ = ( (~ n184) ) ;
 assign o_38_ = ( (~ n178) ) ;
 assign o_39_ = ( (~ n173) ) ;
 assign o_40_ = ( (~ n166) ) ;
 assign o_41_ = ( (~ n161) ) ;
 assign o_42_ = ( (~ n154) ) ;
 assign o_43_ = ( (~ n146) ) ;
 assign o_44_ = ( (~ n144) ) ;
 assign o_45_ = ( (~ n138) ) ;
 assign o_46_ = ( (~ n134) ) ;
 assign o_47_ = ( (~ n129) ) ;
 assign o_48_ = ( (~ n127) ) ;
 assign o_49_ = ( (~ n122) ) ;
 assign o_50_ = ( (~ n115) ) ;
 assign o_51_ = ( (~ n110) ) ;
 assign o_52_ = ( (~ n102) ) ;
 assign o_53_ = ( (~ n96) ) ;
 assign o_54_ = ( (~ n90) ) ;
 assign o_55_ = ( (~ n84) ) ;
 assign o_56_ = ( (~ n75) ) ;
 assign o_57_ = ( (~ n67) ) ;
 assign o_58_ = ( (~ n59) ) ;
 assign o_59_ = ( (~ n52) ) ;
 assign o_60_ = ( (~ n43) ) ;
 assign o_61_ = ( (~ n34) ) ;
 assign o_62_ = ( (~ n28) ) ;
 assign n2 = ( n24 ) | ( n321 ) ;
 assign n3 = ( n24 ) | ( n323 ) ;
 assign n1 = ( n2  &  n3 ) ;
 assign n5 = ( n317 ) | ( n209 ) ;
 assign n6 = ( n328 ) | ( n209 ) ;
 assign n4 = ( n5  &  n6 ) ;
 assign n8 = ( n346 ) | ( n20 ) ;
 assign n9 = ( n347 ) | ( n20 ) ;
 assign n7 = ( n8  &  n9 ) ;
 assign n11 = ( n321 ) | ( n20 ) ;
 assign n12 = ( n323 ) | ( n20 ) ;
 assign n10 = ( n11  &  n12 ) ;
 assign n14 = ( n312 ) | ( n20 ) ;
 assign n15 = ( n329 ) | ( n20 ) ;
 assign n13 = ( n14  &  n15 ) ;
 assign n17 = ( n312 ) | ( n244 ) ;
 assign n18 = ( n312 ) | ( n240 ) ;
 assign n16 = ( n17  &  n18 ) ;
 assign n20 = ( (~ i_0_) ) | ( i_1_ ) | ( i_2_ ) ;
 assign n19 = ( n20 ) | ( (~ n253) ) ;
 assign n23 = ( (~ i_3_) ) | ( (~ i_4_) ) | ( (~ i_5_) ) ;
 assign n24 = ( i_0_ ) | ( i_1_ ) | ( (~ i_2_) ) ;
 assign n22 = ( n23 ) | ( n24 ) ;
 assign n26 = ( i_0_ ) | ( i_1_ ) | ( i_2_ ) ;
 assign n25 = ( n26 ) | ( (~ n237) ) ;
 assign n29 = ( n244  &  n208 ) ;
 assign n30 = ( n399  &  n389  &  n233 ) ;
 assign n31 = ( n400  &  n209  &  n139  &  n65  &  n379 ) ;
 assign n32 = ( n49  &  n341  &  n285  &  n345  &  n243 ) ;
 assign n33 = ( n18  &  n401  &  n402  &  n46  &  n336 ) ;
 assign n28 = ( n29  &  n30  &  n31  &  n32  &  n33 ) ;
 assign n35 = ( n273  &  n419  &  n421 ) ;
 assign n36 = ( n409  &  n410 ) ;
 assign n37 = ( n287  &  n387 ) ;
 assign n38 = ( n390  &  n233 ) ;
 assign n39 = ( n334  &  n443 ) ;
 assign n40 = ( n245  &  n442  &  n50 ) ;
 assign n41 = ( n124  &  n113  &  n275 ) ;
 assign n42 = ( n403  &  n62  &  n439 ) ;
 assign n34 = ( n35  &  n36  &  n37  &  n38  &  n39  &  n40  &  n41  &  n42 ) ;
 assign n44 = ( n78  &  n179  &  n450  &  n297  &  n124  &  n403 ) ;
 assign n45 = ( n282  &  n444  &  n62  &  n35  &  n342  &  n345  &  n18  &  n401 ) ;
 assign n46 = ( n335  &  n330 ) ;
 assign n47 = ( n232  &  n440  &  n336 ) ;
 assign n48 = ( n240 ) | ( n346 ) ;
 assign n49 = ( n317 ) | ( n283 ) ;
 assign n50 = ( n317 ) | ( n140 ) ;
 assign n51 = ( n240 ) | ( n347 ) ;
 assign n43 = ( n44  &  n45  &  n46  &  n47  &  n48  &  n49  &  n50  &  n51 ) ;
 assign n53 = ( n26  &  n286  &  n287 ) | ( (~ n254)  &  n286  &  n287 ) ;
 assign n54 = ( n436  &  n168 ) ;
 assign n55 = ( n293  &  n109 ) | ( n293  &  n283 ) ;
 assign n56 = ( n457  &  n458  &  n180  &  n215  &  n39  &  n204  &  n125  &  n33 ) ;
 assign n57 = ( n135  &  n461  &  n40  &  n73 ) ;
 assign n58 = ( (~ n252)  &  n260  &  n270  &  n285  &  n368  &  n370  &  n377  &  n482 ) ;
 assign n52 = ( n53  &  n54  &  n55  &  n56  &  n57  &  n58 ) ;
 assign n60 = ( n8  &  n167  &  (~ n235)  &  n289  &  n330  &  n418  &  n463  &  n464 ) ;
 assign n61 = ( (~ n252)  &  n375  &  n377 ) ;
 assign n62 = ( n280  &  n437  &  n277  &  n10  &  n438  &  n435 ) ;
 assign n63 = ( n450  &  n142 ) ;
 assign n64 = ( n297  &  n369  &  n370 ) ;
 assign n65 = ( n362  &  n363  &  n358  &  n360 ) ;
 assign n66 = ( n221  &  n25  &  n23 ) | ( n221  &  n25  &  n26 ) ;
 assign n59 = ( n60  &  n61  &  n62  &  n63  &  n64  &  n65  &  n6  &  n66 ) ;
 assign n68 = ( n355  &  n353 ) ;
 assign n69 = ( n18  &  n423 ) ;
 assign n70 = ( n140 ) | ( n325 ) ;
 assign n71 = ( n131  &  n356  &  n267 ) ;
 assign n72 = ( n98  &  n209  &  n289 ) | ( n98  &  (~ n254)  &  n289 ) ;
 assign n73 = ( n49  &  n460 ) ;
 assign n74 = ( n91  &  n85  &  n296  &  n55  &  n298  &  n170 ) ;
 assign n67 = ( n68  &  n69  &  n70  &  n71  &  n36  &  n72  &  n73  &  n74 ) ;
 assign n76 = ( n466  &  n467  &  n439  &  n39 ) ;
 assign n77 = ( n180  &  n465 ) ;
 assign n78 = ( n379  &  n449 ) ;
 assign n79 = ( (~ n268)  &  n376  &  n468 ) ;
 assign n80 = ( n17  &  n250  &  n241  &  n294  &  n176 ) ;
 assign n81 = ( n385  &  n450 ) ;
 assign n82 = ( n50  &  n403 ) ;
 assign n83 = ( n98  &  n41  &  n350  &  n66  &  n482  &  n248  &  n422  &  n356 ) ;
 assign n75 = ( n76  &  n77  &  n78  &  n79  &  n80  &  n81  &  n82  &  n83 ) ;
 assign n85 = ( n450  &  n53 ) ;
 assign n86 = ( (~ n235)  &  n330  &  n425 ) ;
 assign n87 = ( n422  &  n145  &  n4  &  n7 ) ;
 assign n88 = ( n458  &  n459  &  n54  &  n469  &  n207  &  n470 ) ;
 assign n89 = ( n22  &  n41  &  n303  &  n70 ) ;
 assign n84 = ( n85  &  n86  &  n50  &  n36  &  n87  &  n88  &  n89 ) ;
 assign n91 = ( n272  &  n50  &  n29 ) ;
 assign n92 = ( n359  &  n117 ) ;
 assign n93 = ( n404  &  n218  &  n380 ) ;
 assign n94 = ( n357  &  n355 ) ;
 assign n95 = ( n460  &  n463  &  n362  &  n424  &  n25  &  n341  &  n422  &  n353 ) ;
 assign n90 = ( n79  &  n89  &  n63  &  n91  &  n92  &  n93  &  n94  &  n95 ) ;
 assign n97 = ( n333  &  n335 ) ;
 assign n98 = ( n411  &  n412 ) ;
 assign n99 = ( n14  &  n413  &  n414  &  n415  &  n416 ) ;
 assign n100 = ( n265  &  n266  &  n264 ) | ( n265  &  n266  &  n209 ) ;
 assign n101 = ( n361  &  n471  &  n425  &  n5  &  n9  &  n422 ) ;
 assign n96 = ( n44  &  n88  &  n97  &  n98  &  n99  &  n100  &  n101 ) ;
 assign n103 = ( n221  &  n85 ) ;
 assign n104 = ( n124  &  n380  &  n447  &  n395  &  n132  &  n162  &  n300 ) ;
 assign n105 = ( n260  &  n376 ) ;
 assign n106 = ( n257  &  n258  &  n244 ) | ( n257  &  n258  &  n256 ) ;
 assign n107 = ( n396  &  n436 ) ;
 assign n102 = ( n103  &  n104  &  n94  &  n105  &  n106  &  n56  &  n32  &  n107 ) ;
 assign n109 = ( (~ n253)  &  (~ n254) ) ;
 assign n108 = ( n24 ) | ( n109 ) ;
 assign n111 = ( n125  &  n108  &  n261  &  n260  &  n472  &  n376 ) ;
 assign n112 = ( n372  &  n373 ) ;
 assign n113 = ( n297  &  n366 ) ;
 assign n114 = ( n124  &  n380  &  n337 ) ;
 assign n110 = ( n45  &  n82  &  n97  &  n103  &  n111  &  n112  &  n113  &  n114 ) ;
 assign n116 = ( n444  &  n73 ) ;
 assign n117 = ( n285  &  n283 ) | ( (~ n253)  &  (~ n254)  &  n285 ) ;
 assign n118 = ( n70  &  n368  &  n371 ) ;
 assign n119 = ( n428  &  n426 ) ;
 assign n120 = ( n410  &  n62  &  n287  &  n385  &  n38  &  n158  &  n163 ) ;
 assign n121 = ( n421  &  n430  &  n431  &  n360  &  n251  &  n419 ) ;
 assign n115 = ( n116  &  n117  &  n118  &  n119  &  n120  &  n121 ) ;
 assign n123 = ( n158  &  n118  &  n212  &  n474  &  n136 ) ;
 assign n124 = ( n24 ) | ( n329 ) ;
 assign n125 = ( n24 ) | ( n325 ) ;
 assign n126 = ( n220  &  n25  &  n221  &  n405 ) ;
 assign n122 = ( n63  &  n105  &  n123  &  n124  &  n125  &  n126 ) ;
 assign n128 = ( n124  &  n111  &  n3  &  n2 ) ;
 assign n127 = ( n128  &  n123  &  n112  &  n30 ) ;
 assign n130 = ( n325 ) | ( n209 ) ;
 assign n131 = ( n312 ) | ( n209 ) ;
 assign n132 = ( n302  &  n151  &  n118 ) ;
 assign n133 = ( n292  &  n94  &  n264 ) | ( n292  &  n94  &  n140 ) ;
 assign n129 = ( n130  &  n60  &  n4  &  n131  &  n132  &  n120  &  n133 ) ;
 assign n135 = ( n297  &  n22  &  n353  &  n70 ) ;
 assign n136 = ( n80  &  n473  &  n215  &  n77 ) ;
 assign n137 = ( n66  &  n379  &  n30  &  n272  &  n50  &  n400 ) ;
 assign n134 = ( n135  &  n61  &  n76  &  n133  &  n136  &  n137 ) ;
 assign n139 = ( n64  &  n66  &  (~ n252)  &  n375  &  n377 ) ;
 assign n140 = ( i_0_ ) | ( (~ i_1_) ) | ( i_2_ ) ;
 assign n141 = ( n130  &  n131 ) ;
 assign n142 = ( n386  &  n200  &  n295  &  n286  &  n383  &  n384 ) ;
 assign n143 = ( n465  &  n76  &  n80 ) ;
 assign n138 = ( n139  &  n38  &  n140  &  n141  &  n142  &  n87  &  n143 ) ;
 assign n145 = ( n416  &  n455  &  n14  &  n415 ) ;
 assign n144 = ( n81  &  n143  &  n31  &  n145 ) ;
 assign n147 = ( n5  &  n98  &  (~ n268)  &  (~ n290)  &  n366  &  n416  &  n453 ) ;
 assign n148 = ( n66  &  n200  &  n330  &  n305  &  n124  &  n376  &  n476  &  n477 ) ;
 assign n149 = ( n367  &  n233  &  n371  &  n388 ) ;
 assign n150 = ( n50  &  n140 ) | ( n50  &  n225 ) ;
 assign n151 = ( n361  &  n471  &  n353  &  n272 ) ;
 assign n152 = ( n168  &  n292  &  n92 ) ;
 assign n153 = ( n394  &  n280  &  n382  &  n393  &  n243  &  n247  &  n49  &  n483 ) ;
 assign n146 = ( n147  &  n148  &  n119  &  n149  &  n150  &  n151  &  n152  &  n153 ) ;
 assign n155 = ( n360  &  n267  &  n356  &  n250 ) ;
 assign n156 = ( n288  &  n298  &  n478  &  n6  &  n12  &  n98 ) ;
 assign n157 = ( n49  &  n441 ) ;
 assign n158 = ( n296  &  n113 ) ;
 assign n159 = ( n294  &  n295  &  n467 ) ;
 assign n160 = ( n435  &  n281  &  n282  &  n450  &  n457  &  n286  &  n251  &  n484 ) ;
 assign n154 = ( n155  &  n156  &  n118  &  n148  &  n157  &  n158  &  n159  &  n160 ) ;
 assign n162 = ( n20  &  n158  &  n277 ) | ( n158  &  (~ n237)  &  n277 ) ;
 assign n163 = ( n196  &  n300  &  n128 ) ;
 assign n164 = ( n473  &  n474  &  n215  &  n118 ) ;
 assign n165 = ( n434  &  n280  &  n444  &  n427  &  n430  &  n431 ) ;
 assign n161 = ( n162  &  n163  &  n164  &  n63  &  n77  &  n93  &  n165 ) ;
 assign n167 = ( n341  &  n116  &  n117 ) ;
 assign n168 = ( n279  &  n434 ) ;
 assign n169 = ( n226  &  n437  &  n451 ) ;
 assign n170 = ( n124  &  n275  &  n430 ) ;
 assign n171 = ( n280  &  n188  &  n354  &  n423  &  n361  &  n352  &  n359  &  n283 ) ;
 assign n172 = ( n366  &  n286  &  n19  &  n209  &  n251  &  n200  &  n409 ) ;
 assign n166 = ( n145  &  n167  &  n168  &  n169  &  n170  &  n149  &  n171  &  n172 ) ;
 assign n174 = ( n461  &  n55  &  n469  &  n475  &  n185  &  n37  &  n73  &  n479 ) ;
 assign n175 = ( n19  &  n417 ) ;
 assign n176 = ( n226  &  n451  &  n54 ) ;
 assign n177 = ( n7  &  n10  &  n64  &  n131  &  (~ n254)  &  n355 ) ;
 assign n173 = ( n147  &  n155  &  n174  &  n175  &  n176  &  n128  &  n177 ) ;
 assign n179 = ( n66  &  n375  &  n448 ) ;
 assign n180 = ( n7  &  n145  &  (~ n290) ) ;
 assign n181 = ( n17  &  n168  &  n294 ) ;
 assign n182 = ( n15  &  n241  &  n393 ) ;
 assign n183 = ( n197  &  n387  &  n233 ) ;
 assign n178 = ( n179  &  n180  &  n76  &  n164  &  n181  &  n182  &  n78  &  n183 ) ;
 assign n185 = ( n463  &  n464  &  n342  &  n336 ) ;
 assign n186 = ( n332  &  n398  &  n343 ) ;
 assign n187 = ( n331  &  n397  &  n1  &  n10  &  n412  &  n381  &  n344 ) ;
 assign n188 = ( n411  &  n362  &  n363 ) ;
 assign n189 = ( n280  &  n449  &  n466  &  n100  &  n418  &  n239 ) ;
 assign n190 = ( n429  &  n443  &  n15  &  n333  &  n396  &  n438  &  n452  &  n485 ) ;
 assign n184 = ( n185  &  n186  &  n187  &  n81  &  n104  &  n188  &  n189  &  n190 ) ;
 assign n192 = ( n360  &  n437  &  n212  &  n188  &  n181  &  n356  &  n355  &  n480 ) ;
 assign n193 = ( n14  &  n478 ) ;
 assign n194 = ( (~ n254)  &  n260  &  n376  &  n417  &  n436  &  n448 ) ;
 assign n195 = ( n226  &  n392 ) ;
 assign n196 = ( n112  &  n126 ) ;
 assign n197 = ( n366  &  n124 ) ;
 assign n191 = ( n192  &  n193  &  n63  &  n194  &  n195  &  n196  &  n197  &  n64 ) ;
 assign n199 = ( n20  &  n195  &  n223 ) | ( n195  &  n223  &  (~ n253) ) ;
 assign n200 = ( n400  &  n381 ) ;
 assign n201 = ( n417  &  n371  &  n369 ) ;
 assign n198 = ( n113  &  n163  &  n192  &  n193  &  n199  &  n200  &  n81  &  n201 ) ;
 assign n203 = ( n11  &  n20 ) | ( n11  &  (~ n254) ) ;
 assign n204 = ( n140  &  n291  &  n292 ) | ( (~ n237)  &  n291  &  n292 ) ;
 assign n205 = ( n403  &  n273  &  n113  &  n50  &  n124  &  n393 ) ;
 assign n202 = ( n156  &  n174  &  n194  &  n168  &  n203  &  n204  &  n205 ) ;
 assign n207 = ( n460  &  n466  &  n157 ) ;
 assign n208 = ( n20  &  n394  &  n182  &  n279  &  n397  &  n398 ) ;
 assign n209 = ( i_0_ ) | ( (~ i_1_) ) | ( (~ i_2_) ) ;
 assign n206 = ( n86  &  n171  &  n81  &  n207  &  n208  &  n78  &  n209  &  n139 ) ;
 assign n211 = ( n437  &  n181  &  n199 ) ;
 assign n212 = ( n76  &  n93 ) ;
 assign n213 = ( n50  &  n366 ) ;
 assign n210 = ( n149  &  n211  &  n128  &  n212  &  n196  &  n142  &  n35  &  n213 ) ;
 assign n215 = ( n72  &  n288  &  n453 ) ;
 assign n216 = ( n99  &  n175  &  n200  &  n233  &  (~ n290)  &  n389  &  n409 ) ;
 assign n214 = ( n215  &  n76  &  n41  &  n204  &  n94  &  n132  &  n211  &  n216 ) ;
 assign n218 = ( n26 ) | ( n241 ) ;
 assign n219 = ( n404  &  n405 ) ;
 assign n220 = ( n23 ) | ( n26 ) ;
 assign n221 = ( n328 ) | ( n26 ) ;
 assign n217 = ( n218  &  n219  &  n220  &  n221 ) ;
 assign n223 = ( n20 ) | ( (~ n237) ) ;
 assign n222 = ( n19  &  n223 ) ;
 assign n225 = ( n316 ) | ( n324 ) ;
 assign n226 = ( n324 ) | ( n327 ) ;
 assign n224 = ( n225  &  n226 ) ;
 assign n228 = ( n26 ) | ( n346 ) ;
 assign n229 = ( n372  &  n400  &  n48  &  n440  &  n186  &  n272  &  n371  &  n481 ) ;
 assign n230 = ( n320 ) | ( (~ n237)  &  (~ n253) ) ;
 assign n227 = ( n11  &  n228  &  n2  &  n8  &  n229  &  n230 ) ;
 assign n232 = ( n283 ) | ( n347 ) ;
 assign n233 = ( n228  &  n391 ) ;
 assign n234 = ( n353  &  n368  &  n373  &  n7  &  n395  &  n349 ) ;
 assign n231 = ( n51  &  n232  &  n233  &  n187  &  n229  &  n234 ) ;
 assign n237 = ( i_3_  &  i_4_  &  (~ i_5_) ) ;
 assign n235 = ( (~ n23)  &  (~ n240) ) | ( n237  &  (~ n240) ) ;
 assign n242 = ( n240 ) | ( n226  &  n250 ) ;
 assign n240 = ( (~ i_0_) ) | ( (~ i_1_) ) | ( (~ i_2_) ) ;
 assign n241 = ( n320 ) | ( n327 ) ;
 assign n239 = ( n242  &  n240 ) | ( n242  &  n241 ) ;
 assign n245 = ( n328 ) | ( n244 ) ;
 assign n244 = ( (~ i_0_) ) | ( i_1_ ) | ( (~ i_2_) ) ;
 assign n243 = ( n245  &  n244 ) | ( n23  &  (~ n237)  &  n245 ) ;
 assign n246 = ( n209 ) | ( n109 ) ;
 assign n248 = ( n348  &  n349 ) ;
 assign n247 = ( n248  &  n140 ) | ( n248  &  n23 ) ;
 assign n250 = ( n322 ) | ( n327 ) ;
 assign n249 = ( n140 ) | ( n226  &  n250 ) ;
 assign n251 = ( n50  &  n140 ) | ( n50  &  (~ n253) ) ;
 assign n253 = ( (~ i_3_)  &  i_4_  &  (~ i_5_) ) ;
 assign n254 = ( (~ i_3_)  &  i_4_  &  i_5_ ) ;
 assign n252 = ( (~ n24)  &  n253 ) | ( (~ n24)  &  n254 ) ;
 assign n257 = ( n244 ) | ( n225 ) ;
 assign n258 = ( n317 ) | ( n244 ) ;
 assign n256 = ( n316 ) | ( n322 ) ;
 assign n260 = ( n24 ) | ( n317 ) ;
 assign n259 = ( n24  &  n260 ) | ( (~ n253)  &  n260 ) ;
 assign n261 = ( n24 ) | ( n225  &  n256 ) ;
 assign n262 = ( (~ n23)  &  (~ n26) ) | ( (~ n26)  &  n237 ) ;
 assign n265 = ( n250 ) | ( n209 ) ;
 assign n266 = ( n8  &  n6  &  n454 ) ;
 assign n264 = ( n23  &  (~ n237) ) ;
 assign n267 = ( n130  &  n248  &  n264 ) | ( n130  &  n248  &  n140 ) ;
 assign n268 = ( (~ n209)  &  n253 ) | ( (~ n209)  &  n254 ) ;
 assign n272 = ( n140 ) | ( n321 ) ;
 assign n270 = ( n140  &  n272 ) | ( (~ n254)  &  n272 ) ;
 assign n273 = ( n68  &  n140  &  n270 ) | ( n68  &  (~ n253)  &  n270 ) ;
 assign n274 = ( n24 ) | ( (~ n254) ) ;
 assign n275 = ( n1  &  n109 ) | ( n1  &  n24 ) ;
 assign n276 = ( n240 ) | ( n225  &  n256 ) ;
 assign n279 = ( n325 ) | ( n244 ) ;
 assign n278 = ( n316 ) | ( n320 ) ;
 assign n277 = ( n17  &  n279  &  n244 ) | ( n17  &  n279  &  n278 ) ;
 assign n280 = ( n106  &  n109 ) | ( n106  &  n244 ) ;
 assign n281 = ( n245  &  n264 ) | ( n245  &  n244 ) ;
 assign n284 = ( n283 ) | ( n328 ) ;
 assign n285 = ( n343  &  n344 ) ;
 assign n283 = ( (~ i_0_) ) | ( (~ i_1_) ) | ( i_2_ ) ;
 assign n282 = ( n284  &  n285  &  n264 ) | ( n284  &  n285  &  n283 ) ;
 assign n286 = ( n317 ) | ( n26 ) ;
 assign n287 = ( n26 ) | ( (~ n253) ) ;
 assign n288 = ( n5  &  n209 ) | ( n5  &  (~ n253) ) ;
 assign n289 = ( n265  &  n452  &  n422 ) ;
 assign n290 = ( (~ n23)  &  (~ n209) ) | ( (~ n209)  &  n237 ) ;
 assign n291 = ( n141  &  n247 ) ;
 assign n292 = ( n356  &  n249 ) ;
 assign n293 = ( n284  &  n339  &  n340 ) ;
 assign n294 = ( n244  &  n258 ) | ( (~ n253)  &  n258 ) ;
 assign n295 = ( n26  &  n287 ) | ( (~ n254)  &  n287 ) ;
 assign n297 = ( n24 ) | ( (~ n237) ) ;
 assign n296 = ( n297  &  n24 ) | ( n297  &  n23 ) ;
 assign n298 = ( n209 ) | ( n109  &  n264 ) ;
 assign n299 = ( n244 ) | ( n264 ) ;
 assign n301 = ( n24 ) | ( n226  &  n250 ) ;
 assign n300 = ( n301  &  n24 ) | ( n301  &  n241 ) ;
 assign n303 = ( n312 ) | ( n140 ) ;
 assign n304 = ( n140 ) | ( n256  &  n278 ) ;
 assign n302 = ( n150  &  n303  &  n304 ) ;
 assign n306 = ( n283 ) | ( n312  &  n325 ) ;
 assign n305 = ( n256  &  n225  &  n306 ) ;
 assign n309 = ( i_3_ ) | ( i_4_ ) | ( i_5_ ) ;
 assign n310 = ( (~ i_6_) ) | ( (~ i_7_) ) ;
 assign n312 = ( n309 ) | ( n310 ) ;
 assign n316 = ( i_3_ ) | ( i_4_ ) | ( (~ i_5_) ) ;
 assign n317 = ( n310 ) | ( n316 ) ;
 assign n319 = ( (~ i_3_) ) | ( i_4_ ) | ( i_5_ ) ;
 assign n320 = ( i_6_ ) | ( i_7_ ) ;
 assign n321 = ( n319 ) | ( n320 ) ;
 assign n322 = ( i_6_ ) | ( (~ i_7_) ) ;
 assign n323 = ( n319 ) | ( n322 ) ;
 assign n324 = ( (~ i_6_) ) | ( i_7_ ) ;
 assign n325 = ( n309 ) | ( n324 ) ;
 assign n327 = ( (~ i_3_) ) | ( i_4_ ) | ( (~ i_5_) ) ;
 assign n328 = ( n310 ) | ( n327 ) ;
 assign n329 = ( n310 ) | ( n319 ) ;
 assign n331 = ( n240 ) | ( n323 ) ;
 assign n332 = ( n240 ) | ( n321 ) ;
 assign n333 = ( n240 ) | ( n329 ) ;
 assign n334 = ( n319 ) | ( n324 ) ;
 assign n330 = ( n331  &  n332  &  n333  &  n334 ) ;
 assign n335 = ( n317 ) | ( n240 ) ;
 assign n337 = ( n240 ) | ( n328 ) ;
 assign n336 = ( (~ n235)  &  n337 ) ;
 assign n339 = ( n283 ) | ( n226 ) ;
 assign n340 = ( n283 ) | ( n250 ) ;
 assign n342 = ( n283 ) | ( n329 ) ;
 assign n341 = ( n342  &  n293 ) ;
 assign n343 = ( n321 ) | ( n283 ) ;
 assign n344 = ( n323 ) | ( n283 ) ;
 assign n345 = ( n278  &  n305 ) ;
 assign n346 = ( n309 ) | ( n320 ) ;
 assign n347 = ( n309 ) | ( n322 ) ;
 assign n348 = ( n209 ) | ( n346 ) ;
 assign n349 = ( n209 ) | ( n347 ) ;
 assign n351 = ( n278 ) | ( n209 ) ;
 assign n350 = ( n351  &  n141 ) ;
 assign n353 = ( n140 ) | ( n323 ) ;
 assign n352 = ( n353  &  n272 ) ;
 assign n355 = ( n140 ) | ( n329 ) ;
 assign n356 = ( n140 ) | ( n328 ) ;
 assign n357 = ( n140 ) | ( n241 ) ;
 assign n354 = ( n355  &  n249  &  n356  &  n357 ) ;
 assign n359 = ( n140 ) | ( (~ n237) ) ;
 assign n358 = ( n359  &  n354 ) ;
 assign n361 = ( n140 ) | ( (~ n254) ) ;
 assign n360 = ( n361  &  n352 ) ;
 assign n362 = ( n247  &  n350 ) ;
 assign n364 = ( n256 ) | ( n209 ) ;
 assign n365 = ( n225 ) | ( n209 ) ;
 assign n363 = ( n364  &  n246  &  n5  &  n365 ) ;
 assign n366 = ( n24 ) | ( n328 ) ;
 assign n368 = ( n140 ) | ( n347 ) ;
 assign n367 = ( n303  &  n70  &  n368 ) ;
 assign n369 = ( n367  &  n251 ) ;
 assign n371 = ( n140 ) | ( n346 ) ;
 assign n370 = ( n371  &  n22 ) ;
 assign n372 = ( n24 ) | ( n346 ) ;
 assign n373 = ( n24 ) | ( n347 ) ;
 assign n374 = ( n125  &  n112 ) ;
 assign n376 = ( n312 ) | ( n24 ) ;
 assign n375 = ( n260  &  n376  &  n374 ) ;
 assign n377 = ( n1  &  n197 ) ;
 assign n380 = ( n329 ) | ( n26 ) ;
 assign n381 = ( n323 ) | ( n26 ) ;
 assign n379 = ( n380  &  n381 ) ;
 assign n383 = ( n225 ) | ( n26 ) ;
 assign n384 = ( n256 ) | ( n26 ) ;
 assign n382 = ( n286  &  n383  &  n384 ) ;
 assign n386 = ( n278 ) | ( n26 ) ;
 assign n385 = ( n386  &  n382 ) ;
 assign n388 = ( n312 ) | ( n26 ) ;
 assign n387 = ( n388  &  n385 ) ;
 assign n390 = ( n325 ) | ( n26 ) ;
 assign n389 = ( n287  &  n390  &  n387 ) ;
 assign n391 = ( n26 ) | ( n347 ) ;
 assign n392 = ( n328 ) | ( n20 ) ;
 assign n393 = ( n250  &  n195 ) ;
 assign n395 = ( n323 ) | ( n244 ) ;
 assign n396 = ( n321 ) | ( n244 ) ;
 assign n394 = ( n395  &  n396 ) ;
 assign n397 = ( n244 ) | ( n347 ) ;
 assign n398 = ( n244 ) | ( n346 ) ;
 assign n399 = ( n26 ) | ( (~ n254) ) ;
 assign n400 = ( n321 ) | ( n26 ) ;
 assign n401 = ( n240 ) | ( n325 ) ;
 assign n402 = ( n264 ) | ( n283 ) ;
 assign n403 = ( n371  &  n22  &  n367 ) ;
 assign n404 = ( n250 ) | ( n26 ) ;
 assign n405 = ( n226 ) | ( n26 ) ;
 assign n408 = ( n472  &  n376  &  n125 ) ;
 assign n406 = ( n219  &  n221  &  n259  &  n261  &  (~ n262)  &  n372  &  n373  &  n408 ) ;
 assign n409 = ( n380  &  n406 ) ;
 assign n410 = ( n399  &  n200 ) ;
 assign n411 = ( n321 ) | ( n209 ) ;
 assign n412 = ( n323 ) | ( n209 ) ;
 assign n413 = ( n225 ) | ( n20 ) ;
 assign n414 = ( n256 ) | ( n20 ) ;
 assign n415 = ( n278 ) | ( n20 ) ;
 assign n416 = ( n325 ) | ( n20 ) ;
 assign n417 = ( n317 ) | ( n20 ) ;
 assign n418 = ( n9  &  n99  &  n175 ) ;
 assign n419 = ( n5  &  n71  &  (~ n268) ) ;
 assign n422 = ( n329 ) | ( n209 ) ;
 assign n421 = ( n100  &  n418  &  n422  &  n98 ) ;
 assign n423 = ( n401  &  n51  &  n48 ) ;
 assign n425 = ( n109 ) | ( n240 ) ;
 assign n424 = ( n425  &  n330  &  n336  &  n276  &  n239 ) ;
 assign n426 = ( n284  &  n339 ) ;
 assign n428 = ( (~ n237) ) | ( n283 ) ;
 assign n429 = ( n283 ) | ( n241 ) ;
 assign n427 = ( n428  &  n285  &  n426  &  n340  &  n429  &  n342 ) ;
 assign n430 = ( n335  &  n424 ) ;
 assign n432 = ( n240 ) | ( n278 ) ;
 assign n433 = ( n23 ) | ( n283 ) ;
 assign n431 = ( n432  &  n433  &  n69 ) ;
 assign n434 = ( n398  &  n397 ) ;
 assign n436 = ( n23 ) | ( n20 ) ;
 assign n435 = ( n195  &  n434  &  n223  &  n436 ) ;
 assign n437 = ( n15  &  n250  &  n241 ) ;
 assign n438 = ( n20 ) | ( (~ n254) ) ;
 assign n440 = ( n283 ) | ( n346 ) ;
 assign n441 = ( n109 ) | ( n283 ) ;
 assign n439 = ( n430  &  n431  &  n345  &  n427  &  n440  &  n441  &  n49  &  n232 ) ;
 assign n442 = ( n244 ) | ( (~ n254) ) ;
 assign n443 = ( n329 ) | ( n244 ) ;
 assign n445 = ( n226 ) | ( n244 ) ;
 assign n446 = ( n250 ) | ( n244 ) ;
 assign n447 = ( n244 ) | ( n241 ) ;
 assign n444 = ( n394  &  n39  &  n281  &  n445  &  n446  &  n447 ) ;
 assign n448 = ( n1  &  (~ n252) ) ;
 assign n449 = ( n400  &  n399  &  n287 ) ;
 assign n450 = ( n388  &  n38 ) ;
 assign n451 = ( n392  &  n223 ) ;
 assign n452 = ( n209 ) | ( n241 ) ;
 assign n454 = ( n226 ) | ( n209 ) ;
 assign n453 = ( n6  &  n454 ) ;
 assign n455 = ( n417  &  n413  &  n414 ) ;
 assign n457 = ( n19  &  n203 ) ;
 assign n458 = ( n12  &  n169 ) ;
 assign n459 = ( n17  &  n294 ) ;
 assign n460 = ( n232  &  n440  &  n345 ) ;
 assign n461 = ( n196  &  n459  &  n410  &  n38 ) ;
 assign n462 = ( n335  &  n425  &  n276 ) ;
 assign n463 = ( n402  &  n69 ) ;
 assign n464 = ( n432  &  n462 ) ;
 assign n465 = ( n19  &  n203  &  n12  &  n15 ) ;
 assign n466 = ( n446  &  n299  &  n245  &  n445 ) ;
 assign n467 = ( n395  &  n396  &  n442 ) ;
 assign n468 = ( n220  &  n374 ) ;
 assign n469 = ( n39  &  n467 ) ;
 assign n470 = ( n354  &  n423  &  n457  &  n18  &  n341  &  n141 ) ;
 assign n471 = ( n140 ) | ( (~ n253) ) ;
 assign n472 = ( n24 ) | ( n278 ) ;
 assign n473 = ( n351  &  n291  &  n365  &  n364 ) ;
 assign n474 = ( n302  &  n151  &  n133 ) ;
 assign n475 = ( n422  &  n380 ) ;
 assign n476 = ( n342  &  n131  &  n355 ) ;
 assign n477 = ( n468  &  n475  &  n455  &  n462  &  n423  &  n47  &  n259  &  n275 ) ;
 assign n478 = ( n7  &  n416 ) ;
 assign n479 = ( n330  &  n285  &  n243 ) ;
 assign n480 = ( n10  &  n209  &  n359 ) ;
 assign n481 = ( n396  &  n411  &  n348 ) ;
 assign n482 = ( n109 ) | ( n140 ) ;
 assign n483 = ( n433  &  n130 ) ;
 assign n484 = ( n16  &  n279  &  n303 ) ;
 assign n485 = ( n293  &  n358  &  n406  &  n422  &  n218  &  n274 ) ;


endmodule

