module _salsaa_qmap_o (input reset, input clk, input data_req, input start, input [255:0] key, input [63:0] nonce, output data_valid, output reg [31:0] data);



	wire g65, g64, g7197, g88, g7198, g111, g7199, g134, g7200, g157, g7201;
	wire g180, g7202, g203, g7203, g226, g7204, g249, g7205, g272, g7206, g295;
	wire g7207, g318, g7208, g341, g7209, g364, g7210, g387, g7211, g410, g7212;
	wire g433, g7213, g456, g7214, g479, g7215, g502, g7216, g525, g7217, g548;
	wire g7218, g571, g7219, g594, g7220, g617, g7221, g640, g7222, g663, g7223;
	wire g686, g7224, g709, g7225, g732, g7226, g755, g7227, g778, g7228, g37;
	wire g797, g796, g7229, g799, g7230, g44, g49, g54, g59, g825, g7231;
	wire g826, g7232, g7233, g62, g832, g829, g7234, g70, g75, g80, g85;
	wire g86, g865, g7235, g93, g98, g103, g108, g109, g899, g7236, g116;
	wire g121, g126, g131, g132, g932, g7237, g139, g144, g149, g154, g155;
	wire g966, g7238, g162, g167, g172, g177, g178, g999, g7239, g185, g190;
	wire g195, g200, g201, g1033, g7240, g208, g213, g218, g223, g224, g1066;
	wire g7241, g231, g236, g241, g246, g247, g1100, g7242, g254, g259, g264;
	wire g269, g270, g1133, g7243, g277, g282, g287, g292, g293, g1167, g7244;
	wire g300, g305, g310, g315, g316, g1204, g7245, g323, g328, g333, g338;
	wire g339, g1237, g7246, g346, g351, g356, g361, g362, g1271, g7247, g369;
	wire g374, g379, g384, g385, g1305, g7248, g392, g397, g402, g407, g408;
	wire g1338, g7249, g415, g420, g425, g430, g431, g1374, g7250, g438, g443;
	wire g448, g453, g454, g1407, g7251, g461, g466, g471, g476, g477, g1441;
	wire g7252, g484, g489, g494, g499, g500, g1475, g7253, g507, g512, g517;
	wire g522, g523, g1508, g7254, g530, g535, g540, g545, g546, g1545, g7255;
	wire g553, g558, g563, g568, g569, g1578, g7256, g576, g581, g586, g591;
	wire g592, g1612, g7257, g599, g604, g609, g614, g615, g1645, g7258, g622;
	wire g627, g632, g637, g638, g1679, g7259, g645, g650, g655, g660, g661;
	wire g1712, g7260, g668, g673, g678, g683, g684, g1746, g7261, g691, g696;
	wire g701, g706, g707, g1782, g7262, g714, g719, g724, g729, g730, g1815;
	wire g7263, g737, g742, g747, g752, g753, g1849, g7264, g760, g765, g770;
	wire g775, g776, g1882, g7265, g780, g781, g782, g783, g784, g785, g786;
	wire g787, g788, g789, g1885, g7266, g791, g1887, g7267, g793, g1889, g7268;
	wire g795, g798, g1891, g7269, g801, g1893, g7270, g803, g1895, g7271, g805;
	wire g1897, g7272, g807, g1899, g7273, g809, g1901, g7274, g811, g1903, g7275;
	wire g813, g1905, g7276, g815, g1907, g7277, g817, g1909, g7278, g819, g1911;
	wire g7279, g821, g1913, g7280, g823, g824, g1938, g1937, g7281, g2017, g7190;
	wire g7282, g833, g2021, g7283, g835, g2023, g7284, g837, g2024, g7285, g839;
	wire g2025, g7286, g841, g2027, g7287, g843, g2029, g7288, g845, g2031, g7289;
	wire g847, g2033, g7290, g849, g2035, g7291, g851, g2037, g7292, g853, g2039;
	wire g7293, g855, g2040, g7294, g857, g2042, g7295, g859, g2044, g7296, g861;
	wire g2046, g7297, g863, g7184, g7298, g866, g2054, g7299, g868, g2057, g7300;
	wire g870, g2059, g7301, g872, g2061, g7302, g874, g2064, g7303, g876, g2067;
	wire g7304, g878, g2070, g7305, g880, g2073, g7306, g882, g2076, g7307, g884;
	wire g2079, g7308, g886, g2082, g7309, g888, g2084, g7310, g890, g2087, g7311;
	wire g892, g2090, g7312, g894, g2093, g7313, g896, g7177, g7314, g898, g900;
	wire g2103, g7315, g902, g2105, g7316, g904, g2106, g7317, g906, g2107, g7318;
	wire g908, g2109, g7319, g910, g2111, g7320, g912, g2113, g7321, g914, g2115;
	wire g7322, g916, g2117, g7323, g918, g2119, g7324, g920, g2121, g7325, g922;
	wire g2122, g7326, g924, g2124, g7327, g926, g2126, g7328, g928, g2128, g7329;
	wire g930, g7171, g7330, g933, g2136, g7331, g935, g2139, g7332, g937, g2141;
	wire g7333, g939, g2143, g7334, g941, g2146, g7335, g943, g2149, g7336, g945;
	wire g2152, g7337, g947, g2155, g7338, g949, g2158, g7339, g951, g2161, g7340;
	wire g953, g2164, g7341, g955, g2166, g7342, g957, g2169, g7343, g959, g2172;
	wire g7344, g961, g2175, g7345, g963, g7165, g7346, g965, g967, g2183, g7347;
	wire g969, g2185, g7348, g971, g2186, g7349, g973, g2187, g7350, g975, g2189;
	wire g7351, g977, g2191, g7352, g979, g2193, g7353, g981, g2195, g7354, g983;
	wire g2197, g7355, g985, g2199, g7356, g987, g2201, g7357, g989, g2202, g7358;
	wire g991, g2204, g7359, g993, g2206, g7360, g995, g2208, g7361, g997, g7158;
	wire g7362, g1000, g2216, g7363, g1002, g2219, g7364, g1004, g2221, g7365, g1006;
	wire g2223, g7366, g1008, g2226, g7367, g1010, g2229, g7368, g1012, g2232, g7369;
	wire g1014, g2235, g7370, g1016, g2238, g7371, g1018, g2241, g7372, g1020, g2244;
	wire g7373, g1022, g2246, g7374, g1024, g2249, g7375, g1026, g2252, g7376, g1028;
	wire g2255, g7377, g1030, g2265, g7378, g1032, g1034, g2266, g7379, g1036, g2268;
	wire g7380, g1038, g2269, g7381, g1040, g2270, g7382, g1042, g2272, g7383, g1044;
	wire g2274, g7384, g1046, g2276, g7385, g1048, g2278, g7386, g1050, g2280, g7387;
	wire g1052, g2282, g7388, g1054, g2284, g7389, g1056, g2285, g7390, g1058, g2287;
	wire g7391, g1060, g2289, g7392, g1062, g2291, g7393, g1064, g2301, g7394, g1067;
	wire g2303, g7395, g1069, g2306, g7396, g1071, g2308, g7397, g1073, g2310, g7398;
	wire g1075, g2313, g7399, g1077, g2316, g7400, g1079, g2319, g7401, g1081, g2322;
	wire g7402, g1083, g2325, g7403, g1085, g2328, g7404, g1087, g2331, g7405, g1089;
	wire g2333, g7406, g1091, g2336, g7407, g1093, g2339, g7408, g1095, g2342, g7409;
	wire g1097, g7152, g7410, g1099, g1101, g2349, g7411, g1103, g2351, g7412, g1105;
	wire g2352, g7413, g1107, g2353, g7414, g1109, g2355, g7415, g1111, g2357, g7416;
	wire g1113, g2359, g7417, g1115, g2361, g7418, g1117, g2363, g7419, g1119, g2365;
	wire g7420, g1121, g2367, g7421, g1123, g2368, g7422, g1125, g2370, g7423, g1127;
	wire g2372, g7424, g1129, g2374, g7425, g1131, g7146, g7426, g1134, g2382, g7427;
	wire g1136, g2385, g7428, g1138, g2387, g7429, g1140, g2389, g7430, g1142, g2392;
	wire g7431, g1144, g2395, g7432, g1146, g2398, g7433, g1148, g2401, g7434, g1150;
	wire g2404, g7435, g1152, g2407, g7436, g1154, g2410, g7437, g1156, g2412, g7438;
	wire g1158, g2415, g7439, g1160, g2418, g7440, g1162, g2421, g7441, g1164, g7140;
	wire g7442, g1166, g1168, g2433, g7443, g1170, g2439, g7444, g1172, g2444, g7445;
	wire g1174, g2449, g7446, g1176, g2455, g7447, g1178, g2461, g7448, g1180, g2467;
	wire g7449, g1182, g2473, g7450, g1184, g2479, g7451, g1186, g2485, g7452, g1188;
	wire g2491, g7453, g1190, g2496, g7454, g1192, g2502, g7455, g1194, g2508, g7456;
	wire g1196, g2514, g7457, g1198, g2521, g7458, g1200, g1201, g1202, g1203, g1205;
	wire g2522, g7459, g1207, g2524, g7460, g1209, g2525, g7461, g1211, g2526, g7462;
	wire g1213, g2528, g7463, g1215, g2530, g7464, g1217, g2532, g7465, g1219, g2534;
	wire g7466, g1221, g2536, g7467, g1223, g2538, g7468, g1225, g2540, g7469, g1227;
	wire g2541, g7470, g1229, g2543, g7471, g1231, g2545, g7472, g1233, g2547, g7473;
	wire g1235, g7133, g7474, g1238, g2558, g7475, g1240, g2561, g7476, g1242, g2563;
	wire g7477, g1244, g2565, g7478, g1246, g2568, g7479, g1248, g2571, g7480, g1250;
	wire g2574, g7481, g1252, g2577, g7482, g1254, g2580, g7483, g1256, g2583, g7484;
	wire g1258, g2586, g7485, g1260, g2588, g7486, g1262, g2591, g7487, g1264, g2594;
	wire g7488, g1266, g2597, g7489, g1268, g2604, g7490, g1270, g1272, g2606, g7491;
	wire g1274, g2609, g7492, g1276, g2611, g7493, g1278, g2613, g7494, g1280, g2616;
	wire g7495, g1282, g2619, g7496, g1284, g2622, g7497, g1286, g2625, g7498, g1288;
	wire g2628, g7499, g1290, g2631, g7500, g1292, g2634, g7501, g1294, g2636, g7502;
	wire g1296, g2639, g7503, g1298, g2642, g7504, g1300, g2645, g7505, g1302, g7126;
	wire g7506, g1304, g1306, g2652, g7507, g1308, g2654, g7508, g1310, g2655, g7509;
	wire g1312, g2656, g7510, g1314, g2658, g7511, g1316, g2660, g7512, g1318, g2662;
	wire g7513, g1320, g2664, g7514, g1322, g2666, g7515, g1324, g2668, g7516, g1326;
	wire g2670, g7517, g1328, g2671, g7518, g1330, g2673, g7519, g1332, g2675, g7520;
	wire g1334, g2677, g7521, g1336, g2685, g7522, g1339, g2689, g7523, g1341, g2694;
	wire g7524, g1343, g2698, g7525, g1345, g2702, g7526, g1347, g2707, g7527, g1349;
	wire g2712, g7528, g1351, g2717, g7529, g1353, g2722, g7530, g1355, g2727, g7531;
	wire g1357, g2732, g7532, g1359, g2737, g7533, g1361, g2741, g7534, g1363, g2746;
	wire g7535, g1365, g2751, g7536, g1367, g2756, g7537, g1369, g2762, g7538, g5721;
	wire g5722, g1371, g1372, g1373, g1375, g2763, g7539, g1377, g2765, g7540, g1379;
	wire g2766, g7541, g1381, g2767, g7542, g1383, g2769, g7543, g1385, g2771, g7544;
	wire g1387, g2773, g7545, g1389, g2775, g7546, g1391, g2777, g7547, g1393, g2779;
	wire g7548, g1395, g2781, g7549, g1397, g2782, g7550, g1399, g2784, g7551, g1401;
	wire g2786, g7552, g1403, g2788, g7553, g1405, g7120, g7554, g1408, g2796, g7555;
	wire g1410, g2799, g7556, g1412, g2801, g7557, g1414, g2803, g7558, g1416, g2806;
	wire g7559, g1418, g2809, g7560, g1420, g2812, g7561, g1422, g2815, g7562, g1424;
	wire g2818, g7563, g1426, g2821, g7564, g1428, g2824, g7565, g1430, g2826, g7566;
	wire g1432, g2829, g7567, g1434, g2832, g7568, g1436, g2835, g7569, g1438, g7114;
	wire g7570, g1440, g1442, g2837, g7571, g1444, g2840, g7572, g1446, g2842, g7573;
	wire g1448, g2844, g7574, g1450, g2847, g7575, g1452, g2850, g7576, g1454, g2853;
	wire g7577, g1456, g2856, g7578, g1458, g2859, g7579, g1460, g2862, g7580, g1462;
	wire g2865, g7581, g1464, g2867, g7582, g1466, g2870, g7583, g1468, g2873, g7584;
	wire g1470, g2876, g7585, g1472, g2879, g7586, g1474, g1476, g2880, g7587, g1478;
	wire g2882, g7588, g1480, g2883, g7589, g1482, g2884, g7590, g1484, g2886, g7591;
	wire g1486, g2888, g7592, g1488, g2890, g7593, g1490, g2892, g7594, g1492, g2894;
	wire g7595, g1494, g2896, g7596, g1496, g2898, g7597, g1498, g2899, g7598, g1500;
	wire g2901, g7599, g1502, g2903, g7600, g1504, g2905, g7601, g1506, g2910, g7602;
	wire g1509, g2915, g7603, g1511, g2921, g7604, g1513, g2926, g7605, g1515, g2931;
	wire g7606, g1517, g2937, g7607, g1519, g2943, g7608, g1521, g2949, g7609, g1523;
	wire g2955, g7610, g1525, g2961, g7611, g1527, g2967, g7612, g1529, g2973, g7613;
	wire g1531, g2978, g7614, g1533, g2984, g7615, g1535, g2990, g7616, g1537, g2996;
	wire g7617, g1539, g7107, g7618, g1541, g1542, g1543, g1544, g1546, g2998, g7619;
	wire g1548, g3000, g7620, g1550, g3001, g7621, g1552, g3002, g7622, g1554, g3004;
	wire g7623, g1556, g3006, g7624, g1558, g3008, g7625, g1560, g3010, g7626, g1562;
	wire g3012, g7627, g1564, g3014, g7628, g1566, g3016, g7629, g1568, g3017, g7630;
	wire g1570, g3019, g7631, g1572, g3021, g7632, g1574, g3023, g7633, g1576, g3028;
	wire g7634, g1579, g3030, g7635, g1581, g3033, g7636, g1583, g3035, g7637, g1585;
	wire g3037, g7638, g1587, g3040, g7639, g1589, g3043, g7640, g1591, g3046, g7641;
	wire g1593, g3049, g7642, g1595, g3052, g7643, g1597, g3055, g7644, g1599, g3058;
	wire g7645, g1601, g3060, g7646, g1603, g3063, g7647, g1605, g3066, g7648, g1607;
	wire g3069, g7649, g1609, g3072, g7650, g1611, g1613, g3073, g7651, g1615, g3075;
	wire g7652, g1617, g3076, g7653, g1619, g3077, g7654, g1621, g3079, g7655, g1623;
	wire g3081, g7656, g1625, g3083, g7657, g1627, g3085, g7658, g1629, g3087, g7659;
	wire g1631, g3089, g7660, g1633, g3091, g7661, g1635, g3092, g7662, g1637, g3094;
	wire g7663, g1639, g3096, g7664, g1641, g3098, g7665, g1643, g3103, g7666, g1646;
	wire g3105, g7667, g1648, g3108, g7668, g1650, g3110, g7669, g1652, g3112, g7670;
	wire g1654, g3115, g7671, g1656, g3118, g7672, g1658, g3121, g7673, g1660, g3124;
	wire g7674, g1662, g3127, g7675, g1664, g3130, g7676, g1666, g3133, g7677, g1668;
	wire g3135, g7678, g1670, g3138, g7679, g1672, g3141, g7680, g1674, g3144, g7681;
	wire g1676, g3147, g7682, g1678, g1680, g3148, g7683, g1682, g3150, g7684, g1684;
	wire g3151, g7685, g1686, g3152, g7686, g1688, g3154, g7687, g1690, g3156, g7688;
	wire g1692, g3158, g7689, g1694, g3160, g7690, g1696, g3162, g7691, g1698, g3164;
	wire g7692, g1700, g3166, g7693, g1702, g3167, g7694, g1704, g3169, g7695, g1706;
	wire g3171, g7696, g1708, g3173, g7697, g1710, g7101, g7698, g1713, g3176, g7699;
	wire g1715, g3179, g7700, g1717, g3181, g7701, g1719, g3183, g7702, g1721, g3186;
	wire g7703, g1723, g3189, g7704, g1725, g3192, g7705, g1727, g3195, g7706, g1729;
	wire g3198, g7707, g1731, g3201, g7708, g1733, g3204, g7709, g1735, g3206, g7710;
	wire g1737, g3209, g7711, g1739, g3212, g7712, g1741, g3215, g7713, g1743, g7095;
	wire g7714, g1745, g1747, g3221, g7715, g1749, g3226, g7716, g1751, g3230, g7717;
	wire g1753, g3234, g7718, g1755, g3239, g7719, g1757, g3244, g7720, g1759, g3249;
	wire g7721, g1761, g3254, g7722, g1763, g3259, g7723, g1765, g3264, g7724, g1767;
	wire g3269, g7725, g1769, g3273, g7726, g1771, g3278, g7727, g1773, g3283, g7728;
	wire g1775, g3288, g7729, g1777, g7089, g7730, g1779, g1780, g1781, g1783, g3290;
	wire g7731, g1785, g3292, g7732, g1787, g3293, g7733, g1789, g3294, g7734, g1791;
	wire g3296, g7735, g1793, g3298, g7736, g1795, g3300, g7737, g1797, g3302, g7738;
	wire g1799, g3304, g7739, g1801, g3306, g7740, g1803, g3308, g7741, g1805, g3309;
	wire g7742, g1807, g3311, g7743, g1809, g3313, g7744, g1811, g3315, g7745, g1813;
	wire g3320, g7746, g5648, g1816, g3322, g7747, g1818, g3325, g7748, g1820, g3327;
	wire g7749, g1822, g3329, g7750, g1824, g3332, g7751, g1826, g3335, g7752, g1828;
	wire g3338, g7753, g1830, g3341, g7754, g1832, g3344, g7755, g1834, g3347, g7756;
	wire g1836, g3350, g7757, g1838, g3352, g7758, g1840, g3355, g7759, g1842, g3358;
	wire g7760, g1844, g3361, g7761, g1846, g3364, g7762, g1848, g1850, g3365, g7763;
	wire g1852, g3367, g7764, g1854, g3368, g7765, g1856, g3369, g7766, g1858, g3371;
	wire g7767, g1860, g3373, g7768, g1862, g3375, g7769, g1864, g3377, g7770, g1866;
	wire g3379, g7771, g1868, g3381, g7772, g1870, g3383, g7773, g1872, g3384, g7774;
	wire g1874, g3386, g7775, g1876, g3388, g7776, g1878, g3390, g7777, g1880, g7083;
	wire g7778, g1883, g3429, g3428, g7779, g3464, g3462, g7780, g3499, g3498, g7781;
	wire g3534, g7782, g7053, g7783, g3587, g7784, g3620, g7785, g3653, g7786, g3688;
	wire g7787, g7012, g7788, g3744, g7789, g3777, g7790, g3810, g7791, g3845, g7792;
	wire g6982, g7793, g3869, g3868, g7794, g3872, g7795, g3873, g7796, g3874, g7797;
	wire g3875, g7798, g3876, g7799, g3877, g7800, g1921, g3878, g7801, g1923, g3880;
	wire g3879, g7802, g3881, g7803, g3884, g7804, g3885, g7805, g3886, g7806, g3887;
	wire g7807, g1930, g3888, g7808, g3889, g7809, g1933, g1934, g3890, g7810, g1936;
	wire g3895, g7811, g3901, g7812, g3904, g7813, g3911, g7814, g1943, g3920, g7815;
	wire g3924, g7816, g3929, g7817, g3933, g7818, g3938, g7819, g3941, g7820, g1950;
	wire g1951, g1952, g3944, g7821, g3947, g7822, g3950, g7823, g6971, g7824, g1957;
	wire g3957, g7825, g3961, g7826, g3963, g7827, g3967, g7828, g3970, g7829, g3973;
	wire g7830, g1964, g1965, g1966, g3978, g7831, g3981, g7832, g3984, g7833, g6961;
	wire g7834, g1971, g3989, g7835, g3992, g7836, g1974, g3995, g7837, g3997, g7838;
	wire g4001, g7839, g4007, g7840, g4011, g7841, g4018, g7842, g1981, g4028, g7843;
	wire g4032, g7844, g4037, g7845, g4041, g7846, g4047, g7847, g4050, g7848, g1988;
	wire g1989, g1990, g4054, g7849, g4057, g7850, g4061, g7851, g6926, g7852, g1995;
	wire g4069, g7853, g4073, g7854, g4076, g7855, g4080, g7856, g2000, g4084, g7857;
	wire g4087, g7858, g4092, g7859, g4095, g7860, g4099, g7861, g6916, g7862, g2007;
	wire g2008, g2009, g2010, g4105, g7863, g4108, g7864, g4111, g7865, g4113, g7866;
	wire g2015, g2016, g2018, g2019, g2020, g4119, g7867, g6887, g7868, g4128, g7869;
	wire g4134, g7870, g4140, g7871, g4146, g7872, g6880, g7873, g4153, g7874, g4159;
	wire g7875, g4164, g7876, g6874, g7877, g4171, g7878, g4174, g7879, g2049, g2050;
	wire g4178, g7880, g4181, g7881, g2053, g4188, g7882, g2056, g2058, g2060, g6855;
	wire g7883, g2063, g4200, g7884, g2066, g4207, g7885, g2069, g4214, g7886, g2072;
	wire g4222, g7887, g2075, g6848, g7888, g2078, g4229, g7889, g2081, g2083, g4236;
	wire g7890, g2086, g4239, g7891, g2089, g6841, g7892, g2092, g2094, g2095, g2096;
	wire g2097, g4246, g7893, g4250, g7894, g4253, g7895, g4257, g7896, g2102, g4261;
	wire g7897, g6824, g7898, g4268, g7899, g4272, g7900, g4276, g7901, g4280, g7902;
	wire g6817, g7903, g4291, g7904, g4295, g7905, g4304, g7906, g6811, g7907, g4309;
	wire g7908, g4312, g7909, g2131, g2132, g4316, g7910, g4319, g7911, g2135, g4323;
	wire g7912, g2138, g2140, g2142, g6782, g7913, g2145, g4330, g7914, g2148, g4334;
	wire g7915, g2151, g4338, g7916, g2154, g4343, g7917, g2157, g6776, g7918, g2160;
	wire g4351, g7919, g2163, g2165, g4355, g7920, g2168, g4360, g7921, g2171, g6769;
	wire g7922, g2174, g2176, g4368, g7923, g4372, g7924, g2179, g4378, g7925, g4382;
	wire g7926, g2182, g4385, g7927, g6762, g7928, g4391, g7929, g4394, g7930, g4397;
	wire g7931, g4400, g7932, g6755, g7933, g4407, g7934, g4410, g7935, g4415, g7936;
	wire g6748, g7937, g2209, g4420, g7938, g4424, g7939, g4427, g7940, g4431, g7941;
	wire g2214, g2215, g4434, g7942, g2218, g2220, g2222, g4439, g7943, g2225, g4442;
	wire g7944, g2228, g4445, g7945, g2231, g4448, g7946, g2234, g4452, g7947, g2237;
	wire g4457, g7948, g2240, g4460, g7949, g2243, g2245, g4463, g7950, g2248, g4466;
	wire g7951, g2251, g4471, g7952, g2254, g4476, g7953, g4479, g7954, g2258, g2259;
	wire g2260, g2261, g4483, g7955, g4486, g7956, g2264, g6713, g7957, g4496, g7958;
	wire g6702, g7959, g6691, g7960, g6680, g7961, g6669, g7962, g4519, g7963, g4522;
	wire g7964, g6658, g7965, g4529, g7966, g4535, g7967, g2292, g2293, g2294, g4538;
	wire g7968, g4542, g7969, g2297, g4546, g7970, g4550, g7971, g2300, g2302, g4554;
	wire g7972, g2305, g2307, g2309, g6651, g7973, g2312, g4560, g7974, g2315, g4564;
	wire g7975, g2318, g4568, g7976, g2321, g4573, g7977, g2324, g6645, g7978, g2327;
	wire g4578, g7979, g2330, g2332, g4582, g7980, g2335, g4585, g7981, g2338, g6638;
	wire g7982, g2341, g4590, g7983, g4593, g7984, g2345, g2346, g4597, g7985, g4600;
	wire g7986, g4604, g7987, g6610, g7988, g4611, g7989, g4615, g7990, g4619, g7991;
	wire g4623, g7992, g6604, g7993, g4627, g7994, g4631, g7995, g4633, g7996, g6598;
	wire g7997, g2375, g4640, g7998, g4644, g7999, g4650, g8000, g4654, g8001, g2380;
	wire g2381, g4657, g8002, g2384, g2386, g2388, g6591, g8003, g2391, g4663, g8004;
	wire g2394, g4666, g8005, g2397, g4669, g8006, g2400, g4673, g8007, g2403, g6584;
	wire g8008, g2406, g4679, g8009, g2409, g2411, g4682, g8010, g2414, g4685, g8011;
	wire g2417, g6577, g8012, g2420, g2422, g4691, g8013, g4694, g8014, g2425, g4697;
	wire g8015, g4700, g8016, g2428, g2429, g2430, g2431, g2432, g4703, g8017, g2435;
	wire g2436, g2437, g2438, g2440, g2441, g2442, g2443, g2445, g2446, g2447, g2448;
	wire g4706, g8018, g2451, g2452, g2453, g2454, g4710, g8019, g2457, g2458, g2459;
	wire g2460, g4713, g8020, g2463, g2464, g2465, g2466, g4716, g8021, g2469, g2470;
	wire g2471, g2472, g4719, g8022, g2475, g2476, g2477, g2478, g4722, g8023, g2481;
	wire g2482, g2483, g2484, g4727, g8024, g2487, g2488, g2489, g2490, g2492, g2493;
	wire g2494, g2495, g4730, g8025, g2498, g2499, g2500, g2501, g4735, g8026, g2504;
	wire g2505, g2506, g2507, g4738, g8027, g2510, g2511, g2512, g2513, g4743, g8028;
	wire g4746, g8029, g2517, g4750, g8030, g4753, g8031, g2520, g6521, g8032, g6515;
	wire g8033, g6505, g8034, g6495, g8035, g6485, g8036, g6475, g8037, g6469, g8038;
	wire g4767, g8039, g6459, g8040, g4770, g8041, g6453, g8042, g2548, g2549, g2550;
	wire g4778, g8043, g4782, g8044, g2553, g5723, g5724, g2554, g4785, g8045, g4789;
	wire g8046, g2557, g4792, g8047, g2560, g2562, g2564, g4795, g8048, g2567, g4799;
	wire g8049, g2570, g4802, g8050, g2573, g4805, g8051, g2576, g4808, g8052, g2579;
	wire g4811, g8053, g2582, g4816, g8054, g2585, g2587, g4819, g8055, g2590, g4824;
	wire g8056, g2593, g4827, g8057, g2596, g4830, g8058, g4832, g8059, g2600, g4836;
	wire g8060, g4838, g8061, g2603, g2605, g4840, g8062, g2608, g2610, g2612, g6403;
	wire g8063, g2615, g4844, g8064, g2618, g4846, g8065, g2621, g4848, g8066, g2624;
	wire g4851, g8067, g2627, g6352, g8068, g2630, g4856, g8069, g2633, g2635, g4858;
	wire g8070, g2638, g4861, g8071, g2641, g6334, g8072, g2644, g2646, g4868, g8073;
	wire g4872, g8074, g4878, g8075, g4882, g8076, g5684, g2651, g4885, g8077, g4889;
	wire g8078, g4893, g8079, g4896, g8080, g4899, g8081, g4902, g8082, g4906, g8083;
	wire g4911, g8084, g4914, g8085, g4919, g8086, g4923, g8087, g4926, g8088, g4929;
	wire g8089, g2680, g2681, g2682, g4932, g8090, g4935, g8091, g5688, g5689, g5690;
	wire g5735, g5736, g2686, g2687, g2688, g4939, g8092, g5747, g5748, g2691, g2692;
	wire g2693, g5759, g5760, g2695, g2696, g2697, g5726, g5727, g2699, g2700, g2701;
	wire g4943, g8093, g5738, g5739, g2704, g2705, g2706, g4947, g8094, g5750, g5751;
	wire g2709, g2710, g2711, g4951, g8095, g5762, g5763, g2714, g2715, g2716, g4955;
	wire g8096, g5729, g5730, g2719, g2720, g2721, g4960, g8097, g5741, g5742, g2724;
	wire g2725, g2726, g4964, g8098, g5753, g5754, g2729, g2730, g2731, g4967, g8099;
	wire g5765, g5766, g2734, g2735, g2736, g5732, g5733, g2738, g2739, g2740, g4971;
	wire g8100, g5744, g5745, g2743, g2744, g2745, g4974, g8101, g5756, g5757, g2748;
	wire g2749, g2750, g4978, g8102, g5768, g5769, g2753, g2754, g2755, g2757, g4981;
	wire g8103, g4984, g8104, g4988, g8105, g4991, g8106, g5692, g5693, g4994, g8107;
	wire g6266, g8108, g5000, g8109, g5003, g8110, g5006, g8111, g5009, g8112, g6216;
	wire g8113, g5014, g8114, g5017, g8115, g5020, g8116, g6199, g8117, g5027, g8118;
	wire g5030, g8119, g2791, g2792, g5034, g8120, g5037, g8121, g2795, g5041, g8122;
	wire g2798, g2800, g2802, g6193, g8123, g2805, g5045, g8124, g2808, g5049, g8125;
	wire g2811, g5053, g8126, g2814, g5058, g8127, g2817, g6187, g8128, g2820, g5063;
	wire g8129, g2823, g2825, g5067, g8130, g2828, g5072, g8131, g2831, g6181, g8132;
	wire g2834, g2836, g5076, g8133, g2839, g2841, g2843, g5079, g8134, g2846, g5084;
	wire g8135, g2849, g5088, g8136, g2852, g5092, g8137, g2855, g5096, g8138, g2858;
	wire g5099, g8139, g2861, g5102, g8140, g2864, g2866, g5106, g8141, g2869, g5109;
	wire g8142, g2872, g5112, g8143, g2875, g2877, g2878, g5115, g8144, g5120, g8145;
	wire g5123, g8146, g5126, g8147, g5129, g8148, g5133, g8149, g5138, g8150, g5143;
	wire g8151, g5146, g8152, g5151, g8153, g5156, g8154, g2906, g2907, g2908, g2909;
	wire g2911, g2912, g2913, g2914, g5160, g8155, g2917, g2918, g2919, g2920, g2922;
	wire g2923, g2924, g2925, g2927, g2928, g2929, g2930, g6174, g8156, g2933, g2934;
	wire g2935, g2936, g5166, g8157, g2939, g2940, g2941, g2942, g5170, g8158, g2945;
	wire g2946, g2947, g2948, g5174, g8159, g2951, g2952, g2953, g2954, g5178, g8160;
	wire g2957, g2958, g2959, g2960, g6167, g8161, g2963, g2964, g2965, g2966, g5182;
	wire g8162, g2969, g2970, g2971, g2972, g2974, g2975, g2976, g2977, g5186, g8163;
	wire g2980, g2981, g2982, g2983, g5189, g8164, g2986, g2987, g2988, g2989, g6160;
	wire g8165, g2992, g2993, g2994, g2995, g2997, g5193, g8166, g5198, g8167, g5201;
	wire g8168, g5204, g8169, g5207, g8170, g5211, g8171, g5216, g8172, g5219, g8173;
	wire g5222, g8174, g5225, g8175, g5230, g8176, g3024, g3025, g3026, g3027, g3029;
	wire g5234, g8177, g3032, g3034, g3036, g5237, g8178, g3039, g5242, g8179, g3042;
	wire g5246, g8180, g3045, g5250, g8181, g3048, g5254, g8182, g3051, g5257, g8183;
	wire g3054, g5262, g8184, g3057, g3059, g5266, g8185, g3062, g5271, g8186, g3065;
	wire g5274, g8187, g3068, g3070, g3071, g5277, g8188, g5282, g8189, g5285, g8190;
	wire g5288, g8191, g5291, g8192, g5295, g8193, g5300, g8194, g5303, g8195, g5306;
	wire g8196, g5309, g8197, g5314, g8198, g3099, g3100, g3101, g3102, g3104, g5317;
	wire g8199, g3107, g3109, g3111, g5320, g8200, g3114, g5324, g8201, g3117, g5327;
	wire g8202, g3120, g5330, g8203, g3123, g5333, g8204, g3126, g5336, g8205, g3129;
	wire g5341, g8206, g3132, g3134, g5344, g8207, g3137, g5349, g8208, g3140, g5352;
	wire g8209, g3143, g3145, g3146, g5356, g8210, g6022, g8211, g5361, g8212, g5365;
	wire g8213, g5369, g8214, g5374, g8215, g6016, g8216, g5378, g8217, g5382, g8218;
	wire g5385, g8219, g6010, g8220, g3174, g3175, g5388, g8221, g3178, g3180, g3182;
	wire g5992, g8222, g3185, g5394, g8223, g3188, g5396, g8224, g3191, g5398, g8225;
	wire g3194, g5400, g8226, g3197, g5953, g8227, g3200, g5405, g8228, g3203, g3205;
	wire g5407, g8229, g3208, g5410, g8230, g3211, g5935, g8231, g3214, g3216, g3217;
	wire g3218, g3219, g3220, g5416, g8232, g3223, g3224, g3225, g3227, g3228, g3229;
	wire g3231, g3232, g3233, g5928, g8233, g3236, g3237, g3238, g5421, g8234, g3241;
	wire g3242, g3243, g5425, g8235, g3246, g3247, g3248, g5429, g8236, g3251, g3252;
	wire g3253, g5435, g8237, g3256, g3257, g3258, g5921, g8238, g3261, g3262, g3263;
	wire g5441, g8239, g3266, g3267, g3268, g3270, g3271, g3272, g5445, g8240, g3275;
	wire g3276, g3277, g5450, g8241, g3280, g3281, g3282, g5915, g8242, g3285, g3286;
	wire g3287, g3289, g5649, g5454, g8243, g5650, g5651, g5652, g5459, g8244, g5653;
	wire g5464, g8245, g5654, g5467, g8246, g5655, g5470, g8247, g5656, g5473, g8248;
	wire g5657, g5478, g8249, g5658, g5481, g8250, g5659, g5660, g5484, g8251, g5661;
	wire g5487, g8252, g5662, g5492, g8253, g5663, g3316, g3317, g3318, g3319, g3321;
	wire g5495, g8254, g3324, g3326, g3328, g5498, g8255, g3331, g5501, g8256, g3334;
	wire g5504, g8257, g3337, g5507, g8258, g3340, g5511, g8259, g3343, g5514, g8260;
	wire g3346, g5517, g8261, g3349, g3351, g5520, g8262, g3354, g5523, g8263, g3357;
	wire g5526, g8264, g3360, g3362, g3363, g5529, g8265, g5844, g8266, g5534, g8267;
	wire g5537, g8268, g5540, g8269, g5543, g8270, g5838, g8271, g5549, g8272, g5552;
	wire g8273, g5557, g8274, g5832, g8275, g3391, g3392, g3393, g3394, g3395, g3396;
	wire g3397, g3398, g3399, g3400, g3401, g3402, g3403, g3404, g3405, g3406, g3407;
	wire g3408, g3409, g3410, g3411, g3412, g3413, g3414, g5794, g5795, g3415, g3416;
	wire g3417, g3418, g3419, g3420, g3421, g3422, g3423, g3424, g3425, g3426, g5560;
	wire g5559, g8276, g3430, g3431, g3432, g3433, g3434, g3435, g3436, g3437, g3438;
	wire g3439, g3440, g3441, g3442, g3443, g3444, g3445, g3446, g3447, g3448, g3449;
	wire g3450, g3451, g3452, g5797, g5798, g3453, g3454, g3455, g3456, g3457, g3458;
	wire g3459, g3460, g3461, g7070, g3463, g3465, g3466, g3467, g3468, g3469, g3470;
	wire g3471, g3472, g3473, g3474, g3475, g3476, g3477, g3478, g3479, g3480, g3481;
	wire g3482, g3483, g3484, g3485, g3486, g3487, g3488, g3489, g3490, g3491, g3492;
	wire g3493, g3494, g3495, g3496, g3497, g7059, g3500, g3501, g3502, g3503, g3504;
	wire g5791, g5792, g3505, g3506, g3507, g3508, g3509, g3510, g3511, g3512, g3513;
	wire g3514, g3515, g3516, g3517, g3518, g3519, g3520, g3521, g3522, g3523, g3524;
	wire g3525, g5815, g5816, g3526, g3527, g3528, g3529, g3530, g3531, g3532, g3533;
	wire g3535, g3536, g3537, g3538, g3539, g5830, g5831, g3540, g3541, g3542, g3543;
	wire g3544, g3545, g3546, g3547, g3548, g3549, g3550, g3551, g3552, g3553, g3554;
	wire g3555, g3556, g3557, g3558, g3559, g5788, g5789, g3560, g3561, g3562, g3563;
	wire g3564, g3565, g3566, g3567, g3568, g3569, g3570, g3571, g3572, g3573, g3574;
	wire g3575, g3576, g3577, g3578, g3579, g3580, g3581, g3582, g3583, g3584, g3585;
	wire g3586, g7042, g3588, g3589, g3590, g3591, g3592, g3593, g3594, g3595, g3596;
	wire g3597, g3598, g3599, g3600, g3601, g3602, g3603, g3604, g3605, g3606, g3607;
	wire g3608, g3609, g3610, g5800, g5801, g3611, g3612, g3613, g3614, g3615, g3616;
	wire g3617, g3618, g3619, g7029, g3621, g3622, g3623, g3624, g3625, g3626, g3627;
	wire g3628, g3629, g5803, g5804, g3630, g3631, g3632, g3633, g3634, g3635, g3636;
	wire g3637, g3638, g3639, g3640, g3641, g3642, g3643, g3644, g3645, g3646, g3647;
	wire g3648, g3649, g3650, g3651, g3652, g7018, g3654, g3655, g3656, g3657, g3658;
	wire g3659, g3660, g3661, g3662, g3663, g3664, g3665, g3666, g3667, g3668, g3669;
	wire g3670, g3671, g3672, g3673, g3674, g3675, g3676, g3677, g5806, g5807, g3678;
	wire g3679, g3680, g3681, g3682, g3683, g3684, g3685, g3686, g5569, g8277, g3689;
	wire g3690, g3691, g3692, g3693, g3694, g3695, g3696, g3697, g3698, g3699, g3700;
	wire g3701, g3702, g3703, g3704, g3705, g3706, g3707, g3708, g3709, g3710, g3711;
	wire g3712, g3713, g3714, g3715, g3716, g3717, g3718, g5818, g5819, g3719, g3720;
	wire g3721, g3722, g3723, g3724, g3725, g3726, g3727, g3728, g3729, g3730, g3731;
	wire g3732, g3733, g3734, g3735, g5821, g5822, g3736, g3737, g3738, g3739, g3740;
	wire g3741, g3742, g3743, g3745, g3746, g3747, g3748, g3749, g3750, g3751, g3752;
	wire g3753, g3754, g3755, g3756, g3757, g3758, g3759, g3760, g3761, g3762, g3763;
	wire g3764, g3765, g3766, g3767, g5809, g5810, g3768, g3769, g3770, g3771, g3772;
	wire g3773, g3774, g3775, g3776, g6999, g3778, g3779, g3780, g3781, g3782, g3783;
	wire g3784, g3785, g3786, g5812, g5813, g3787, g3788, g3789, g3790, g3791, g3792;
	wire g3793, g3794, g3795, g3796, g3797, g3798, g3799, g3800, g3801, g3802, g3803;
	wire g3804, g3805, g3806, g3807, g3808, g3809, g6988, g3811, g3812, g3813, g3814;
	wire g3815, g3816, g3817, g3818, g3819, g5824, g5825, g3820, g3821, g3822, g3823;
	wire g3824, g3825, g3826, g3827, g3828, g3829, g3830, g3831, g3832, g3833, g3834;
	wire g3835, g3836, g5827, g5828, g3837, g3838, g3839, g3840, g3841, g3842, g3843;
	wire g3844, g3846, g3847, g3848, g3849, g3850, g3851, g3852, g3853, g3854, g3855;
	wire g3856, g3857, g3858, g3859, g3860, g3861, g3862, g3863, g3864, g3865, g3866;
	wire g3867, g3870, g3871, g3882, g3883, g3891, g3892, g3893, g3894, g3896, g3897;
	wire g3898, g3899, g3900, g3902, g3903, g3905, g3906, g3907, g3908, g3909, g3910;
	wire g3912, g3913, g3914, g3915, g3916, g3917, g3918, g3919, g3921, g3922, g3923;
	wire g3925, g3926, g3927, g3928, g3930, g3931, g3932, g3934, g3935, g3936, g3937;
	wire g3939, g3940, g5665, g3942, g3943, g3945, g3946, g3948, g3949, g5672, g3951;
	wire g3952, g3953, g3954, g3955, g3956, g3958, g3959, g3960, g3962, g3964, g3965;
	wire g3966, g3968, g3969, g3971, g3972, g3974, g3975, g3976, g3977, g3979, g3980;
	wire g5677, g3982, g3983, g3985, g3986, g3987, g3988, g3990, g3991, g3993, g3994;
	wire g3996, g6950, g3998, g3999, g5570, g8278, g6937, g4002, g4003, g4004, g4005;
	wire g4006, g4008, g4009, g5571, g8279, g4012, g4013, g4014, g4015, g4016, g4017;
	wire g4019, g4020, g4021, g4022, g4023, g4024, g4025, g4026, g5572, g8280, g4029;
	wire g4030, g4031, g4033, g4034, g4035, g5573, g8281, g4038, g4039, g4040, g4042;
	wire g4043, g4044, g4045, g5574, g8282, g5776, g5777, g4048, g4049, g5670, g4051;
	wire g4052, g5575, g8283, g4055, g4056, g4058, g4059, g5576, g8284, g5673, g4062;
	wire g4063, g4064, g4065, g4066, g4067, g5577, g8285, g4070, g4071, g4072, g4074;
	wire g5578, g8286, g4077, g4078, g4079, g4081, g4082, g5579, g8287, g4085, g4086;
	wire g4088, g4089, g4090, g5580, g8288, g4093, g4094, g5682, g4096, g4097, g5581;
	wire g8289, g4100, g4101, g4102, g4103, g5582, g8290, g4106, g4107, g4109, g5584;
	wire g8291, g6905, g4112, g6894, g4114, g4115, g4116, g4117, g4118, g4120, g4121;
	wire g4122, g4123, g4124, g4125, g4126, g5585, g8292, g4129, g4130, g4131, g4132;
	wire g4133, g4135, g4136, g4137, g4138, g4139, g4141, g4142, g4143, g4144, g4145;
	wire g4147, g4148, g4149, g4150, g4151, g4152, g4154, g4155, g4156, g4157, g4158;
	wire g4160, g4161, g4162, g4163, g4165, g4166, g4167, g4168, g4169, g4170, g4172;
	wire g4173, g4175, g4176, g5586, g8293, g6861, g4179, g4180, g4182, g4183, g4184;
	wire g4185, g4186, g4187, g4189, g4190, g4191, g4192, g4193, g4194, g4195, g4196;
	wire g4197, g4198, g4199, g4201, g4202, g4203, g4204, g4205, g4206, g4208, g4209;
	wire g4210, g4211, g4212, g4213, g4215, g4216, g4217, g4218, g4219, g4220, g5587;
	wire g8294, g5771, g5772, g4223, g4224, g4225, g4226, g4227, g4228, g4230, g4231;
	wire g4232, g4233, g4234, g4235, g4237, g4238, g5774, g5775, g4240, g4241, g4242;
	wire g4243, g4244, g4245, g4247, g4248, g4249, g4251, g5588, g8295, g6830, g4254;
	wire g4255, g4256, g4258, g4259, g4260, g4262, g4263, g4264, g4265, g4266, g5589;
	wire g8296, g4269, g4270, g4271, g4273, g4274, g4275, g4277, g4278, g4279, g4281;
	wire g4282, g4283, g4284, g4285, g4286, g4287, g4288, g4289, g4290, g4292, g4293;
	wire g4294, g4296, g4297, g4298, g4299, g4300, g4301, g4302, g4303, g4305, g4306;
	wire g4307, g4308, g4310, g4311, g6800, g4313, g4314, g5591, g8297, g4317, g4318;
	wire g6789, g4320, g4321, g4322, g4324, g4325, g4326, g4327, g4328, g4329, g4331;
	wire g4332, g4333, g4335, g4336, g4337, g4339, g4340, g4341, g5593, g8298, g4344;
	wire g4345, g4346, g4347, g4348, g4349, g4350, g4352, g4353, g4354, g4356, g4357;
	wire g4358, g4359, g4361, g4362, g4363, g4364, g4365, g4366, g4367, g4369, g4370;
	wire g4371, g4373, g4374, g4375, g4376, g5594, g8299, g4379, g4380, g4381, g4383;
	wire g4384, g5664, g4386, g4387, g4388, g4389, g5595, g8300, g5666, g4392, g4393;
	wire g5667, g4395, g4396, g5668, g4398, g4399, g5669, g4401, g4402, g4403, g4404;
	wire g4405, g4406, g4408, g4409, g5671, g4411, g4412, g4413, g4414, g4416, g4417;
	wire g4418, g4419, g4421, g4422, g4423, g4425, g5596, g8301, g6737, g4428, g4429;
	wire g4430, g4432, g4433, g4435, g5778, g5779, g5780, g4436, g4437, g4438, g4440;
	wire g4441, g4443, g4444, g4446, g4447, g4449, g4450, g5598, g8302, g4453, g5781;
	wire g5782, g5783, g4454, g4455, g4456, g4458, g4459, g4461, g4462, g4464, g4465;
	wire g4467, g5784, g5785, g5786, g4468, g4469, g4470, g4472, g4473, g4474, g4475;
	wire g4477, g4478, g4480, g4481, g5599, g8303, g6724, g4484, g4485, g4487, g4488;
	wire g4489, g4490, g4491, g4492, g4493, g4494, g4495, g4497, g4498, g4499, g4500;
	wire g5600, g8304, g4502, g4503, g4504, g4505, g4506, g4507, g4508, g4509, g4510;
	wire g4511, g4512, g4513, g4514, g4515, g4516, g4517, g4518, g4520, g4521, g5674;
	wire g4523, g4524, g4525, g4526, g4527, g4528, g5675, g4530, g4531, g4532, g4533;
	wire g4534, g4536, g4537, g4539, g4540, g4541, g4543, g4544, g5601, g8305, g4547;
	wire g4548, g4549, g4551, g4552, g4553, g4555, g4556, g4557, g4558, g4559, g4561;
	wire g4562, g4563, g4565, g4566, g4567, g4569, g4570, g4571, g5602, g8306, g4574;
	wire g4575, g4576, g4577, g4579, g4580, g4581, g4583, g4584, g4586, g4587, g4588;
	wire g4589, g4591, g4592, g6627, g4594, g4595, g5603, g8307, g4598, g4599, g6616;
	wire g4601, g4602, g4603, g4605, g4606, g4607, g4608, g4609, g5605, g8308, g4612;
	wire g4613, g4614, g4616, g4617, g4618, g4620, g4621, g4622, g4624, g4625, g4626;
	wire g4628, g4629, g4630, g4632, g4634, g4635, g4636, g4637, g4638, g4639, g4641;
	wire g4642, g4643, g4645, g4646, g4647, g4648, g5607, g8309, g4651, g4652, g4653;
	wire g4655, g4656, g4658, g4659, g4660, g4661, g4662, g4664, g4665, g4667, g4668;
	wire g4670, g4671, g5608, g8310, g4674, g4675, g4676, g4677, g4678, g4680, g4681;
	wire g4683, g4684, g4686, g4687, g4688, g4689, g4690, g4692, g4693, g6566, g4695;
	wire g5609, g8311, g6555, g4698, g4699, g6544, g4701, g4702, g5676, g4704, g4705;
	wire g4707, g4708, g5610, g8312, g5678, g4711, g4712, g5679, g4714, g4715, g5680;
	wire g4717, g4718, g5681, g4720, g4721, g4723, g4724, g4725, g4726, g4728, g4729;
	wire g5683, g4731, g4732, g4733, g4734, g4736, g4737, g4739, g4740, g4741, g4742;
	wire g4744, g4745, g4747, g4748, g5611, g8313, g6531, g4751, g4752, g4754, g4755;
	wire g4756, g4757, g4758, g5613, g8314, g4760, g4761, g4762, g4763, g4764, g4765;
	wire g4766, g4768, g4769, g4771, g4772, g4773, g4774, g4775, g4776, g4777, g4779;
	wire g4780, g4781, g4783, g5614, g8315, g6442, g4786, g4787, g4788, g4790, g4791;
	wire g4793, g4794, g4796, g4797, g5615, g8316, g4800, g4801, g4803, g4804, g4806;
	wire g4807, g4809, g4810, g4812, g4813, g4814, g4815, g4817, g4818, g4820, g4821;
	wire g4822, g4823, g4825, g4826, g4828, g4829, g4831, g6431, g4833, g4834, g5617;
	wire g8317, g4837, g6420, g4839, g6409, g4841, g5685, g4842, g4843, g6392, g4845;
	wire g6381, g4847, g6370, g4849, g5619, g8318, g6359, g4852, g5686, g4853, g4854;
	wire g4855, g4857, g6341, g4859, g4860, g4862, g5687, g4863, g4864, g4865, g4866;
	wire g4867, g4869, g4870, g4871, g4873, g4874, g4875, g4876, g5620, g8319, g4879;
	wire g4880, g4881, g4883, g4884, g4886, g4887, g4888, g5710, g5711, g4890, g4891;
	wire g5622, g8320, g4894, g4895, g4897, g4898, g4900, g4901, g4903, g4904, g4905;
	wire g5712, g5713, g4907, g4908, g4909, g4910, g4912, g4913, g4915, g4916, g4917;
	wire g4918, g4920, g4921, g4922, g5714, g5715, g4924, g4925, g4927, g4928, g6297;
	wire g4930, g5624, g8321, g6323, g4933, g4934, g6310, g4936, g4937, g4938, g4940;
	wire g5717, g4941, g4942, g4944, g4945, g4946, g4948, g4949, g4950, g4952, g4953;
	wire g4954, g4956, g4957, g4958, g5625, g8322, g4961, g5718, g4962, g4963, g4965;
	wire g4966, g4968, g4969, g4970, g4972, g4973, g4975, g5719, g4976, g4977, g4979;
	wire g4980, g4982, g4983, g4985, g4986, g5626, g8323, g6284, g4989, g4990, g4992;
	wire g4993, g6273, g4995, g4996, g4997, g4998, g5627, g8324, g6255, g5001, g5002;
	wire g6244, g5004, g5005, g6233, g5007, g5008, g6222, g5010, g5011, g5012, g5013;
	wire g5015, g5016, g6205, g5018, g5019, g5021, g5022, g5023, g5024, g5025, g5026;
	wire g5028, g5029, g5031, g5032, g5628, g8325, g5035, g5036, g5038, g5039, g5040;
	wire g5042, g5043, g5044, g5046, g5047, g5048, g5050, g5051, g5052, g5054, g5055;
	wire g5056, g5629, g8326, g5059, g5060, g5061, g5062, g5064, g5065, g5066, g5068;
	wire g5069, g5070, g5071, g5073, g5074, g5075, g5077, g5078, g5080, g5081, g5082;
	wire g5631, g8327, g5085, g5086, g5087, g5089, g5090, g5091, g5093, g5094, g5095;
	wire g5097, g5098, g5100, g5101, g5103, g5104, g5105, g5107, g5108, g5110, g5111;
	wire g5113, g5114, g5116, g5117, g5118, g5119, g5121, g5122, g5124, g5125, g5127;
	wire g5128, g5130, g5131, g5632, g8328, g5134, g5135, g5136, g5137, g5139, g5140;
	wire g5141, g5142, g5144, g5145, g5147, g5148, g5149, g5150, g5152, g5153, g5154;
	wire g5155, g5157, g5158, g5159, g5161, g5162, g5163, g5164, g5634, g8329, g5167;
	wire g5168, g5169, g5171, g5172, g5173, g5175, g5176, g5177, g5179, g5180, g5181;
	wire g5183, g5184, g5185, g5187, g5188, g5190, g5191, g5192, g6149, g5194, g5195;
	wire g5196, g5197, g5199, g5200, g6138, g5202, g5203, g6127, g5205, g5206, g6116;
	wire g5208, g5209, g5635, g8330, g6105, g5212, g5213, g5214, g5215, g5217, g5218;
	wire g5220, g5221, g6094, g5223, g5224, g5226, g5227, g5228, g5229, g5231, g5232;
	wire g5233, g5235, g5236, g5238, g5239, g5240, g5636, g8331, g5243, g5244, g5245;
	wire g5247, g5248, g5249, g5251, g5252, g5253, g5255, g5256, g5258, g5259, g5260;
	wire g5261, g5263, g5264, g5265, g5267, g5268, g5269, g5270, g5272, g5273, g5275;
	wire g5276, g6083, g5278, g5279, g5280, g5281, g5283, g5284, g6072, g5286, g5287;
	wire g6061, g5289, g5290, g6050, g5292, g5293, g5638, g8332, g6039, g5296, g5297;
	wire g5298, g5299, g5301, g5302, g5304, g5305, g6028, g5307, g5308, g5310, g5311;
	wire g5312, g5313, g5315, g5316, g5318, g5319, g5321, g5322, g5639, g8333, g5325;
	wire g5326, g5328, g5329, g5331, g5332, g5334, g5335, g5337, g5338, g5339, g5340;
	wire g5342, g5343, g5345, g5346, g5347, g5348, g5350, g5351, g5353, g5354, g5355;
	wire g5357, g5358, g5359, g5360, g5362, g5363, g5364, g5366, g5367, g5368, g5370;
	wire g5371, g5372, g5640, g8334, g5375, g5376, g5377, g5379, g5380, g5381, g5383;
	wire g5384, g5386, g5387, g5999, g5389, g5390, g5391, g5392, g5642, g8335, g5395;
	wire g5981, g5397, g5970, g5399, g5959, g5401, g5402, g5403, g5404, g5406, g5942;
	wire g5408, g5409, g5411, g5412, g5413, g5414, g5415, g5417, g5418, g5419, g5420;
	wire g5422, g5423, g5424, g5426, g5427, g5428, g5430, g5431, g5432, g5433, g5643;
	wire g8336, g5436, g5437, g5438, g5439, g5440, g5442, g5443, g5444, g5446, g5447;
	wire g5448, g5449, g5451, g5452, g5453, g5902, g5455, g5456, g5457, g5458, g5460;
	wire g5461, g5462, g5645, g8337, g5465, g5466, g5889, g5468, g5469, g5876, g5471;
	wire g5472, g5863, g5474, g5475, g5476, g5477, g5479, g5480, g5482, g5483, g5850;
	wire g5485, g5486, g5488, g5489, g5490, g5491, g5493, g5494, g5496, g5497, g5499;
	wire g5500, g5502, g5503, g5505, g5506, g5508, g5509, g5646, g8338, g5512, g5513;
	wire g5515, g5516, g5518, g5519, g5521, g5522, g5524, g5525, g5527, g5528, g5530;
	wire g5531, g5532, g5647, g8339, g5535, g5536, g5538, g5539, g5541, g5542, g5544;
	wire g5545, g5546, g5547, g5548, g5550, g5551, g5553, g5554, g5555, g5556, g5558;
	wire g5561, g5562, g5716, g5563, g5564, g5565, g5566, g5567, g5568, g5583, g5590;
	wire g5592, g5597, g5604, g5606, g5612, g5616, g5618, g5621, g5623, g5630, g5633;
	wire g5637, g5641, g5644, g5691, g5694, g5695, g5696, g5697, g5698, g5699, g5700;
	wire g5701, g5702, g5703, g5704, g5705, g5706, g5707, g5708, g5709, g5720, g5725;
	wire g5728, g5731, g5734, g5737, g5740, g5743, g5746, g5749, g5752, g5755, g5758;
	wire g5761, g5764, g5767, g5770, g5773, g5787, g5790, g5793, g5796, g5799, g5802;
	wire g5805, g5808, g5811, g5814, g5817, g5820, g5823, g5826, g5829, g5833, g5834;
	wire g5835, g5836, g5837, g5839, g5840, g5841, g5842, g5843, g5845, g5846, g5847;
	wire g5848, g5849, g5851, g5852, g5853, g5856, g5854, g5855, g5859, g5860, g5857;
	wire g5858, g5861, g5862, g5864, g5865, g5866, g5869, g5867, g5868, g5872, g5873;
	wire g5870, g5871, g5874, g5875, g5877, g5878, g5879, g5882, g5880, g5881, g5885;
	wire g5886, g5883, g5884, g5887, g5888, g5890, g5891, g5892, g5895, g5893, g5894;
	wire g5898, g5899, g5896, g5897, g5900, g5901, g5903, g5904, g5905, g5908, g5906;
	wire g5907, g5911, g5912, g5909, g5910, g5913, g5914, g5916, g5917, g5918, g5919;
	wire g5920, g5922, g5923, g5924, g5925, g5926, g5927, g5929, g5930, g5931, g5932;
	wire g5933, g5934, g5936, g5937, g5938, g5939, g5940, g5941, g5943, g5944, g5945;
	wire g5948, g5946, g5947, g5951, g5949, g5950, g5952, g5954, g5955, g5956, g5957;
	wire g5958, g5960, g5961, g5962, g5965, g5963, g5964, g5968, g5966, g5967, g5969;
	wire g5971, g5972, g5973, g5976, g5974, g5975, g5979, g5977, g5978, g5980, g5982;
	wire g5983, g5984, g5987, g5985, g5986, g5990, g5988, g5989, g5991, g5993, g5994;
	wire g5995, g5996, g5997, g5998, g6000, g6001, g6002, g6005, g6003, g6004, g6008;
	wire g6006, g6007, g6009, g6011, g6012, g6013, g6014, g6015, g6017, g6018, g6019;
	wire g6020, g6021, g6023, g6024, g6025, g6026, g6027, g6029, g6030, g6031, g6034;
	wire g6032, g6033, g6037, g6035, g6036, g6038, g6040, g6041, g6042, g6045, g6043;
	wire g6044, g6048, g6046, g6047, g6049, g6051, g6052, g6053, g6056, g6054, g6055;
	wire g6059, g6057, g6058, g6060, g6062, g6063, g6064, g6067, g6065, g6066, g6070;
	wire g6068, g6069, g6071, g6073, g6074, g6075, g6078, g6076, g6077, g6081, g6079;
	wire g6080, g6082, g6084, g6085, g6086, g6089, g6087, g6088, g6092, g6090, g6091;
	wire g6093, g6095, g6096, g6097, g6100, g6098, g6099, g6103, g6101, g6102, g6104;
	wire g6106, g6107, g6108, g6111, g6109, g6110, g6114, g6112, g6113, g6115, g6117;
	wire g6118, g6119, g6122, g6120, g6121, g6125, g6123, g6124, g6126, g6128, g6129;
	wire g6130, g6133, g6131, g6132, g6136, g6134, g6135, g6137, g6139, g6140, g6141;
	wire g6144, g6142, g6143, g6147, g6145, g6146, g6148, g6150, g6151, g6152, g6155;
	wire g6153, g6154, g6158, g6156, g6157, g6159, g6161, g6162, g6163, g6164, g6165;
	wire g6166, g6168, g6169, g6170, g6171, g6172, g6173, g6175, g6176, g6177, g6178;
	wire g6179, g6180, g6182, g6183, g6184, g6185, g6186, g6188, g6189, g6190, g6191;
	wire g6192, g6194, g6195, g6196, g6197, g6198, g6200, g6201, g6202, g6203, g6204;
	wire g6206, g6207, g6208, g6211, g6209, g6210, g6214, g6212, g6213, g6215, g6217;
	wire g6218, g6219, g6220, g6221, g6223, g6224, g6225, g6228, g6226, g6227, g6231;
	wire g6229, g6230, g6232, g6234, g6235, g6236, g6239, g6237, g6238, g6242, g6240;
	wire g6241, g6243, g6245, g6246, g6247, g6250, g6248, g6249, g6253, g6251, g6252;
	wire g6254, g6256, g6257, g6258, g6261, g6259, g6260, g6264, g6262, g6263, g6265;
	wire g6267, g6268, g6269, g6270, g6271, g6272, g6274, g6275, g6276, g6279, g6277;
	wire g6278, g6282, g6280, g6281, g6283, g6285, g6286, g6287, g6290, g6288, g6289;
	wire g6293, g6294, g6291, g6292, g6295, g6296, g6298, g6299, g6300, g6303, g6301;
	wire g6302, g6306, g6307, g6304, g6305, g6308, g6309, g6311, g6312, g6313, g6316;
	wire g6314, g6315, g6319, g6320, g6317, g6318, g6321, g6322, g6324, g6325, g6326;
	wire g6329, g6327, g6328, g6332, g6330, g6331, g6333, g6335, g6336, g6337, g6338;
	wire g6339, g6340, g6342, g6343, g6344, g6347, g6345, g6346, g6350, g6348, g6349;
	wire g6351, g6353, g6354, g6355, g6356, g6357, g6358, g6360, g6361, g6362, g6365;
	wire g6363, g6364, g6368, g6366, g6367, g6369, g6371, g6372, g6373, g6376, g6374;
	wire g6375, g6379, g6377, g6378, g6380, g6382, g6383, g6384, g6387, g6385, g6386;
	wire g6390, g6388, g6389, g6391, g6393, g6394, g6395, g6398, g6396, g6397, g6401;
	wire g6399, g6400, g6402, g6404, g6405, g6406, g6407, g6408, g6410, g6411, g6412;
	wire g6415, g6413, g6414, g6418, g6416, g6417, g6419, g6421, g6422, g6423, g6426;
	wire g6424, g6425, g6429, g6427, g6428, g6430, g6432, g6433, g6434, g6437, g6435;
	wire g6436, g6440, g6438, g6439, g6441, g6443, g6444, g6445, g6448, g6446, g6447;
	wire g6451, g6449, g6450, g6452, g6454, g6455, g6456, g6457, g6458, g6460, g6461;
	wire g6462, g6465, g6463, g6464, g6468, g6466, g6467, g6470, g6471, g6472, g6473;
	wire g6474, g6476, g6477, g6478, g6481, g6479, g6480, g6482, g6483, g6484, g6486;
	wire g6487, g6488, g6491, g6489, g6490, g6494, g6492, g6493, g6496, g6497, g6498;
	wire g6501, g6499, g6500, g6502, g6503, g6504, g6506, g6507, g6508, g6511, g6509;
	wire g6510, g6514, g6512, g6513, g6516, g6517, g6518, g6519, g6520, g6522, g6523;
	wire g6524, g6527, g6525, g6526, g6528, g6529, g6530, g6532, g6533, g6534, g6537;
	wire g6535, g6536, g6540, g6541, g6538, g6539, g6542, g6543, g6545, g6546, g6547;
	wire g6550, g6548, g6549, g6553, g6551, g6552, g6554, g6556, g6557, g6558, g6561;
	wire g6559, g6560, g6564, g6562, g6563, g6565, g6567, g6568, g6569, g6572, g6570;
	wire g6571, g6575, g6573, g6574, g6576, g6578, g6579, g6580, g6581, g6582, g6583;
	wire g6585, g6586, g6587, g6588, g6589, g6590, g6592, g6593, g6594, g6595, g6596;
	wire g6597, g6599, g6600, g6601, g6602, g6603, g6605, g6606, g6607, g6608, g6609;
	wire g6611, g6612, g6613, g6614, g6615, g6617, g6618, g6619, g6622, g6620, g6621;
	wire g6625, g6623, g6624, g6626, g6628, g6629, g6630, g6633, g6631, g6632, g6636;
	wire g6634, g6635, g6637, g6639, g6640, g6641, g6642, g6643, g6644, g6646, g6647;
	wire g6648, g6649, g6650, g6652, g6653, g6654, g6655, g6656, g6657, g6659, g6660;
	wire g6661, g6664, g6662, g6663, g6665, g6666, g6667, g6668, g6670, g6671, g6672;
	wire g6675, g6673, g6674, g6676, g6677, g6678, g6679, g6681, g6682, g6683, g6686;
	wire g6684, g6685, g6687, g6688, g6689, g6690, g6692, g6693, g6694, g6697, g6695;
	wire g6696, g6698, g6699, g6700, g6701, g6703, g6704, g6705, g6708, g6706, g6707;
	wire g6709, g6710, g6711, g6712, g6714, g6715, g6716, g6719, g6717, g6718, g6720;
	wire g6721, g6722, g6723, g6725, g6726, g6727, g6730, g6728, g6729, g6733, g6734;
	wire g6731, g6732, g6735, g6736, g6738, g6739, g6740, g6743, g6741, g6742, g6746;
	wire g6744, g6745, g6747, g6749, g6750, g6751, g6752, g6753, g6754, g6756, g6757;
	wire g6758, g6759, g6760, g6761, g6763, g6764, g6765, g6766, g6767, g6768, g6770;
	wire g6771, g6772, g6773, g6774, g6775, g6777, g6778, g6779, g6780, g6781, g6783;
	wire g6784, g6785, g6786, g6787, g6788, g6790, g6791, g6792, g6795, g6793, g6794;
	wire g6798, g6796, g6797, g6799, g6801, g6802, g6803, g6806, g6804, g6805, g6809;
	wire g6807, g6808, g6810, g6812, g6813, g6814, g6815, g6816, g6818, g6819, g6820;
	wire g6821, g6822, g6823, g6825, g6826, g6827, g6828, g6829, g6831, g6832, g6833;
	wire g6836, g6834, g6835, g6839, g6837, g6838, g6840, g6842, g6843, g6844, g6845;
	wire g6846, g6847, g6849, g6850, g6851, g6852, g6853, g6854, g6856, g6857, g6858;
	wire g6859, g6860, g6862, g6863, g6864, g6867, g6865, g6866, g6870, g6871, g6868;
	wire g6869, g6872, g6873, g6875, g6876, g6877, g6878, g6879, g6881, g6882, g6883;
	wire g6884, g6885, g6886, g6888, g6889, g6890, g6891, g6892, g6893, g6895, g6896;
	wire g6897, g6900, g6898, g6899, g6903, g6901, g6902, g6904, g6906, g6907, g6908;
	wire g6911, g6909, g6910, g6914, g6912, g6913, g6915, g6917, g6918, g6919, g6922;
	wire g6920, g6921, g6925, g6923, g6924, g6927, g6928, g6929, g6932, g6930, g6931;
	wire g6933, g6934, g6935, g6936, g6938, g6939, g6940, g6943, g6941, g6942, g6946;
	wire g6947, g6944, g6945, g6948, g6949, g6951, g6952, g6953, g6956, g6954, g6955;
	wire g6959, g6957, g6958, g6960, g6962, g6963, g6964, g6967, g6965, g6966, g6968;
	wire g6969, g6970, g6972, g6973, g6974, g6977, g6975, g6976, g6978, g6979, g6980;
	wire g6981, g6983, g6984, g6985, g6986, g6987, g6989, g6990, g6991, g6994, g6992;
	wire g6993, g6997, g6995, g6996, g6998, g7000, g7001, g7002, g7005, g7003, g7004;
	wire g7008, g7009, g7006, g7007, g7010, g7011, g7013, g7014, g7015, g7016, g7017;
	wire g7019, g7020, g7021, g7024, g7022, g7023, g7027, g7025, g7026, g7028, g7030;
	wire g7031, g7032, g7035, g7033, g7034, g7038, g7039, g7036, g7037, g7040, g7041;
	wire g7043, g7044, g7045, g7048, g7046, g7047, g7051, g7049, g7050, g7052, g7054;
	wire g7055, g7056, g7057, g7058, g7060, g7061, g7062, g7065, g7063, g7064, g7068;
	wire g7066, g7067, g7069, g7071, g7072, g7073, g7076, g7074, g7075, g7079, g7080;
	wire g7077, g7078, g7081, g7082, g7084, g7085, g7086, g7087, g7088, g7090, g7091;
	wire g7092, g7093, g7094, g7096, g7097, g7098, g7099, g7100, g7102, g7103, g7104;
	wire g7105, g7106, g7108, g7109, g7110, g7111, g7112, g7113, g7115, g7116, g7117;
	wire g7118, g7119, g7121, g7122, g7123, g7124, g7125, g7127, g7128, g7129, g7130;
	wire g7131, g7132, g7134, g7135, g7136, g7137, g7138, g7139, g7141, g7142, g7143;
	wire g7144, g7145, g7147, g7148, g7149, g7150, g7151, g7153, g7154, g7155, g7156;
	wire g7157, g7159, g7160, g7161, g7162, g7163, g7164, g7166, g7167, g7168, g7169;
	wire g7170, g7172, g7173, g7174, g7175, g7176, g7178, g7179, g7180, g7181, g7182;
	wire g7183, g7185, g7186, g7187, g7188, g7189, g7191, g7192, g7193, g7194, g7195;
	wire g7196;


	reg g1, g34, g35, g36, g38, g39, g40, g41, g42;
	reg g43, g45, g46, g47, g48, g50, g51, g52, g53;
	reg g55, g56, g57, g58, g60, g61, g63, g66, g67;
	reg g68, g69, g71, g72, g73, g74, g76, g77, g78;
	reg g79, g81, g82, g83, g84, g87, g89, g90, g91;
	reg g92, g94, g95, g96, g97, g99, g100, g101, g102;
	reg g104, g105, g106, g107, g110, g112, g113, g114, g115;
	reg g117, g118, g119, g120, g122, g123, g124, g125, g127;
	reg g128, g129, g130, g133, g135, g136, g137, g138, g140;
	reg g141, g142, g143, g145, g146, g147, g148, g150, g151;
	reg g152, g153, g156, g158, g159, g160, g161, g163, g164;
	reg g165, g166, g168, g169, g170, g171, g173, g174, g175;
	reg g176, g179, g181, g182, g183, g184, g186, g187, g188;
	reg g189, g191, g192, g193, g194, g196, g197, g198, g199;
	reg g202, g204, g205, g206, g207, g209, g210, g211, g212;
	reg g214, g215, g216, g217, g219, g220, g221, g222, g225;
	reg g227, g228, g229, g230, g232, g233, g234, g235, g237;
	reg g238, g239, g240, g242, g243, g244, g245, g248, g250;
	reg g251, g252, g253, g255, g256, g257, g258, g260, g261;
	reg g262, g263, g265, g266, g267, g268, g271, g273, g274;
	reg g275, g276, g278, g279, g280, g281, g283, g284, g285;
	reg g286, g288, g289, g290, g291, g294, g296, g297, g298;
	reg g299, g301, g302, g303, g304, g306, g307, g308, g309;
	reg g311, g312, g313, g314, g317, g319, g320, g321, g322;
	reg g324, g325, g326, g327, g329, g330, g331, g332, g334;
	reg g335, g336, g337, g340, g342, g343, g344, g345, g347;
	reg g348, g349, g350, g352, g353, g354, g355, g357, g358;
	reg g359, g360, g363, g365, g366, g367, g368, g370, g371;
	reg g372, g373, g375, g376, g377, g378, g380, g381, g382;
	reg g383, g386, g388, g389, g390, g391, g393, g394, g395;
	reg g396, g398, g399, g400, g401, g403, g404, g405, g406;
	reg g409, g411, g412, g413, g414, g416, g417, g418, g419;
	reg g421, g422, g423, g424, g426, g427, g428, g429, g432;
	reg g434, g435, g436, g437, g439, g440, g441, g442, g444;
	reg g445, g446, g447, g449, g450, g451, g452, g455, g457;
	reg g458, g459, g460, g462, g463, g464, g465, g467, g468;
	reg g469, g470, g472, g473, g474, g475, g478, g480, g481;
	reg g482, g483, g485, g486, g487, g488, g490, g491, g492;
	reg g493, g495, g496, g497, g498, g501, g503, g504, g505;
	reg g506, g508, g509, g510, g511, g513, g514, g515, g516;
	reg g518, g519, g520, g521, g524, g526, g527, g528, g529;
	reg g531, g532, g533, g534, g536, g537, g538, g539, g541;
	reg g542, g543, g544, g547, g549, g550, g551, g552, g554;
	reg g555, g556, g557, g559, g560, g561, g562, g564, g565;
	reg g566, g567, g570, g572, g573, g574, g575, g577, g578;
	reg g579, g580, g582, g583, g584, g585, g587, g588, g589;
	reg g590, g593, g595, g596, g597, g598, g600, g601, g602;
	reg g603, g605, g606, g607, g608, g610, g611, g612, g613;
	reg g616, g618, g619, g620, g621, g623, g624, g625, g626;
	reg g628, g629, g630, g631, g633, g634, g635, g636, g639;
	reg g641, g642, g643, g644, g646, g647, g648, g649, g651;
	reg g652, g653, g654, g656, g657, g658, g659, g662, g664;
	reg g665, g666, g667, g669, g670, g671, g672, g674, g675;
	reg g676, g677, g679, g680, g681, g682, g685, g687, g688;
	reg g689, g690, g692, g693, g694, g695, g697, g698, g699;
	reg g700, g702, g703, g704, g705, g708, g710, g711, g712;
	reg g713, g715, g716, g717, g718, g720, g721, g722, g723;
	reg g725, g726, g727, g728, g731, g733, g734, g735, g736;
	reg g738, g739, g740, g741, g743, g744, g745, g746, g748;
	reg g749, g750, g751, g754, g756, g757, g758, g759, g761;
	reg g762, g763, g764, g766, g767, g768, g769, g771, g772;
	reg g773, g774, g777, g779, g790, g792, g794, g800, g802;
	reg g804, g806, g808, g810, g812, g814, g816, g818, g820;
	reg g822, g827, g828, g830, g831, g834, g836, g838, g840;
	reg g842, g844, g846, g848, g850, g852, g854, g856, g858;
	reg g860, g862, g864, g867, g869, g871, g873, g875, g877;
	reg g879, g881, g883, g885, g887, g889, g891, g893, g895;
	reg g897, g901, g903, g905, g907, g909, g911, g913, g915;
	reg g917, g919, g921, g923, g925, g927, g929, g931, g934;
	reg g936, g938, g940, g942, g944, g946, g948, g950, g952;
	reg g954, g956, g958, g960, g962, g964, g968, g970, g972;
	reg g974, g976, g978, g980, g982, g984, g986, g988, g990;
	reg g992, g994, g996, g998, g1001, g1003, g1005, g1007, g1009;
	reg g1011, g1013, g1015, g1017, g1019, g1021, g1023, g1025, g1027;
	reg g1029, g1031, g1035, g1037, g1039, g1041, g1043, g1045, g1047;
	reg g1049, g1051, g1053, g1055, g1057, g1059, g1061, g1063, g1065;
	reg g1068, g1070, g1072, g1074, g1076, g1078, g1080, g1082, g1084;
	reg g1086, g1088, g1090, g1092, g1094, g1096, g1098, g1102, g1104;
	reg g1106, g1108, g1110, g1112, g1114, g1116, g1118, g1120, g1122;
	reg g1124, g1126, g1128, g1130, g1132, g1135, g1137, g1139, g1141;
	reg g1143, g1145, g1147, g1149, g1151, g1153, g1155, g1157, g1159;
	reg g1161, g1163, g1165, g1169, g1171, g1173, g1175, g1177, g1179;
	reg g1181, g1183, g1185, g1187, g1189, g1191, g1193, g1195, g1197;
	reg g1199, g1206, g1208, g1210, g1212, g1214, g1216, g1218, g1220;
	reg g1222, g1224, g1226, g1228, g1230, g1232, g1234, g1236, g1239;
	reg g1241, g1243, g1245, g1247, g1249, g1251, g1253, g1255, g1257;
	reg g1259, g1261, g1263, g1265, g1267, g1269, g1273, g1275, g1277;
	reg g1279, g1281, g1283, g1285, g1287, g1289, g1291, g1293, g1295;
	reg g1297, g1299, g1301, g1303, g1307, g1309, g1311, g1313, g1315;
	reg g1317, g1319, g1321, g1323, g1325, g1327, g1329, g1331, g1333;
	reg g1335, g1337, g1340, g1342, g1344, g1346, g1348, g1350, g1352;
	reg g1354, g1356, g1358, g1360, g1362, g1364, g1366, g1368, g1370;
	reg g1376, g1378, g1380, g1382, g1384, g1386, g1388, g1390, g1392;
	reg g1394, g1396, g1398, g1400, g1402, g1404, g1406, g1409, g1411;
	reg g1413, g1415, g1417, g1419, g1421, g1423, g1425, g1427, g1429;
	reg g1431, g1433, g1435, g1437, g1439, g1443, g1445, g1447, g1449;
	reg g1451, g1453, g1455, g1457, g1459, g1461, g1463, g1465, g1467;
	reg g1469, g1471, g1473, g1477, g1479, g1481, g1483, g1485, g1487;
	reg g1489, g1491, g1493, g1495, g1497, g1499, g1501, g1503, g1505;
	reg g1507, g1510, g1512, g1514, g1516, g1518, g1520, g1522, g1524;
	reg g1526, g1528, g1530, g1532, g1534, g1536, g1538, g1540, g1547;
	reg g1549, g1551, g1553, g1555, g1557, g1559, g1561, g1563, g1565;
	reg g1567, g1569, g1571, g1573, g1575, g1577, g1580, g1582, g1584;
	reg g1586, g1588, g1590, g1592, g1594, g1596, g1598, g1600, g1602;
	reg g1604, g1606, g1608, g1610, g1614, g1616, g1618, g1620, g1622;
	reg g1624, g1626, g1628, g1630, g1632, g1634, g1636, g1638, g1640;
	reg g1642, g1644, g1647, g1649, g1651, g1653, g1655, g1657, g1659;
	reg g1661, g1663, g1665, g1667, g1669, g1671, g1673, g1675, g1677;
	reg g1681, g1683, g1685, g1687, g1689, g1691, g1693, g1695, g1697;
	reg g1699, g1701, g1703, g1705, g1707, g1709, g1711, g1714, g1716;
	reg g1718, g1720, g1722, g1724, g1726, g1728, g1730, g1732, g1734;
	reg g1736, g1738, g1740, g1742, g1744, g1748, g1750, g1752, g1754;
	reg g1756, g1758, g1760, g1762, g1764, g1766, g1768, g1770, g1772;
	reg g1774, g1776, g1778, g1784, g1786, g1788, g1790, g1792, g1794;
	reg g1796, g1798, g1800, g1802, g1804, g1806, g1808, g1810, g1812;
	reg g1814, g1817, g1819, g1821, g1823, g1825, g1827, g1829, g1831;
	reg g1833, g1835, g1837, g1839, g1841, g1843, g1845, g1847, g1851;
	reg g1853, g1855, g1857, g1859, g1861, g1863, g1865, g1867, g1869;
	reg g1871, g1873, g1875, g1877, g1879, g1881, g1884, g1886, g1888;
	reg g1890, g1892, g1894, g1896, g1898, g1900, g1902, g1904, g1906;
	reg g1908, g1910, g1912, g1914, g1915, g1916, g1917, g1918, g1919;
	reg g1920, g1922, g1924, g1925, g1926, g1927, g1928, g1929, g1931;
	reg g1932, g1935, g1939, g1940, g1941, g1942, g1944, g1945, g1946;
	reg g1947, g1948, g1949, g1953, g1954, g1955, g1956, g1958, g1959;
	reg g1960, g1961, g1962, g1963, g1967, g1968, g1969, g1970, g1972;
	reg g1973, g1975, g1976, g1977, g1978, g1979, g1980, g1982, g1983;
	reg g1984, g1985, g1986, g1987, g1991, g1992, g1993, g1994, g1996;
	reg g1997, g1998, g1999, g2001, g2002, g2003, g2004, g2005, g2006;
	reg g2011, g2012, g2013, g2014, g2022, g2026, g2028, g2030, g2032;
	reg g2034, g2036, g2038, g2041, g2043, g2045, g2047, g2048, g2051;
	reg g2052, g2055, g2062, g2065, g2068, g2071, g2074, g2077, g2080;
	reg g2085, g2088, g2091, g2098, g2099, g2100, g2101, g2104, g2108;
	reg g2110, g2112, g2114, g2116, g2118, g2120, g2123, g2125, g2127;
	reg g2129, g2130, g2133, g2134, g2137, g2144, g2147, g2150, g2153;
	reg g2156, g2159, g2162, g2167, g2170, g2173, g2177, g2178, g2180;
	reg g2181, g2184, g2188, g2190, g2192, g2194, g2196, g2198, g2200;
	reg g2203, g2205, g2207, g2210, g2211, g2212, g2213, g2217, g2224;
	reg g2227, g2230, g2233, g2236, g2239, g2242, g2247, g2250, g2253;
	reg g2256, g2257, g2262, g2263, g2267, g2271, g2273, g2275, g2277;
	reg g2279, g2281, g2283, g2286, g2288, g2290, g2295, g2296, g2298;
	reg g2299, g2304, g2311, g2314, g2317, g2320, g2323, g2326, g2329;
	reg g2334, g2337, g2340, g2343, g2344, g2347, g2348, g2350, g2354;
	reg g2356, g2358, g2360, g2362, g2364, g2366, g2369, g2371, g2373;
	reg g2376, g2377, g2378, g2379, g2383, g2390, g2393, g2396, g2399;
	reg g2402, g2405, g2408, g2413, g2416, g2419, g2423, g2424, g2426;
	reg g2427, g2434, g2450, g2456, g2462, g2468, g2474, g2480, g2486;
	reg g2497, g2503, g2509, g2515, g2516, g2518, g2519, g2523, g2527;
	reg g2529, g2531, g2533, g2535, g2537, g2539, g2542, g2544, g2546;
	reg g2551, g2552, g2555, g2556, g2559, g2566, g2569, g2572, g2575;
	reg g2578, g2581, g2584, g2589, g2592, g2595, g2598, g2599, g2601;
	reg g2602, g2607, g2614, g2617, g2620, g2623, g2626, g2629, g2632;
	reg g2637, g2640, g2643, g2647, g2648, g2649, g2650, g2653, g2657;
	reg g2659, g2661, g2663, g2665, g2667, g2669, g2672, g2674, g2676;
	reg g2678, g2679, g2683, g2684, g2690, g2703, g2708, g2713, g2718;
	reg g2723, g2728, g2733, g2742, g2747, g2752, g2758, g2759, g2760;
	reg g2761, g2764, g2768, g2770, g2772, g2774, g2776, g2778, g2780;
	reg g2783, g2785, g2787, g2789, g2790, g2793, g2794, g2797, g2804;
	reg g2807, g2810, g2813, g2816, g2819, g2822, g2827, g2830, g2833;
	reg g2838, g2845, g2848, g2851, g2854, g2857, g2860, g2863, g2868;
	reg g2871, g2874, g2881, g2885, g2887, g2889, g2891, g2893, g2895;
	reg g2897, g2900, g2902, g2904, g2916, g2932, g2938, g2944, g2950;
	reg g2956, g2962, g2968, g2979, g2985, g2991, g2999, g3003, g3005;
	reg g3007, g3009, g3011, g3013, g3015, g3018, g3020, g3022, g3031;
	reg g3038, g3041, g3044, g3047, g3050, g3053, g3056, g3061, g3064;
	reg g3067, g3074, g3078, g3080, g3082, g3084, g3086, g3088, g3090;
	reg g3093, g3095, g3097, g3106, g3113, g3116, g3119, g3122, g3125;
	reg g3128, g3131, g3136, g3139, g3142, g3149, g3153, g3155, g3157;
	reg g3159, g3161, g3163, g3165, g3168, g3170, g3172, g3177, g3184;
	reg g3187, g3190, g3193, g3196, g3199, g3202, g3207, g3210, g3213;
	reg g3222, g3235, g3240, g3245, g3250, g3255, g3260, g3265, g3274;
	reg g3279, g3284, g3291, g3295, g3297, g3299, g3301, g3303, g3305;
	reg g3307, g3310, g3312, g3314, g3323, g3330, g3333, g3336, g3339;
	reg g3342, g3345, g3348, g3353, g3356, g3359, g3366, g3370, g3372;
	reg g3374, g3376, g3378, g3380, g3382, g3385, g3387, g3389, g3427;
	reg g3687, g4000, g4010, g4027, g4036, g4046, g4053, g4060, g4068;
	reg g4075, g4083, g4091, g4098, g4104, g4110, g4127, g4177, g4221;
	reg g4252, g4267, g4315, g4342, g4377, g4390, g4426, g4451, g4482;
	reg g4501, g4545, g4572, g4596, g4610, g4649, g4672, g4696, g4709;
	reg g4749, g4759, g4784, g4798, g4835, g4850, g4877, g4892, g4931;
	reg g4959, g4987, g4999, g5033, g5057, g5083, g5132, g5165, g5210;
	reg g5241, g5294, g5323, g5373, g5393, g5434, g5463, g5510, g5533;
	always @ (posedge clk) begin g1 <= g37; end
	always @ (posedge clk) begin data[0] <= g7197; end
	always @ (posedge clk) begin data[1] <= g7198; end
	always @ (posedge clk) begin data[2] <= g7199; end
	always @ (posedge clk) begin data[3] <= g7200; end
	always @ (posedge clk) begin data[4] <= g7201; end
	always @ (posedge clk) begin data[5] <= g7202; end
	always @ (posedge clk) begin data[6] <= g7203; end
	always @ (posedge clk) begin data[7] <= g7204; end
	always @ (posedge clk) begin data[8] <= g7205; end
	always @ (posedge clk) begin data[9] <= g7206; end
	always @ (posedge clk) begin data[10] <= g7207; end
	always @ (posedge clk) begin data[11] <= g7208; end
	always @ (posedge clk) begin data[12] <= g7209; end
	always @ (posedge clk) begin data[13] <= g7210; end
	always @ (posedge clk) begin data[14] <= g7211; end
	always @ (posedge clk) begin data[15] <= g7212; end
	always @ (posedge clk) begin data[16] <= g7213; end
	always @ (posedge clk) begin data[17] <= g7214; end
	always @ (posedge clk) begin data[18] <= g7215; end
	always @ (posedge clk) begin data[19] <= g7216; end
	always @ (posedge clk) begin data[20] <= g7217; end
	always @ (posedge clk) begin data[21] <= g7218; end
	always @ (posedge clk) begin data[22] <= g7219; end
	always @ (posedge clk) begin data[23] <= g7220; end
	always @ (posedge clk) begin data[24] <= g7221; end
	always @ (posedge clk) begin data[25] <= g7222; end
	always @ (posedge clk) begin data[26] <= g7223; end
	always @ (posedge clk) begin data[27] <= g7224; end
	always @ (posedge clk) begin data[28] <= g7225; end
	always @ (posedge clk) begin data[29] <= g7226; end
	always @ (posedge clk) begin data[30] <= g7227; end
	always @ (posedge clk) begin data[31] <= g7228; end
	always @ (posedge clk) begin g34 <= g783; end
	always @ (posedge clk) begin g35 <= g784; end
	always @ (posedge clk) begin g36 <= g788; end
	always @ (posedge clk) begin g38 <= g789; end
	always @ (posedge clk) begin g39 <= g791; end
	always @ (posedge clk) begin g40 <= g793; end
	always @ (posedge clk) begin g41 <= g795; end
	always @ (posedge clk) begin g42 <= g7229; end
	always @ (posedge clk) begin g43 <= g7230; end
	always @ (posedge clk) begin g45 <= g801; end
	always @ (posedge clk) begin g46 <= g803; end
	always @ (posedge clk) begin g47 <= g805; end
	always @ (posedge clk) begin g48 <= g807; end
	always @ (posedge clk) begin g50 <= g809; end
	always @ (posedge clk) begin g51 <= g811; end
	always @ (posedge clk) begin g52 <= g813; end
	always @ (posedge clk) begin g53 <= g815; end
	always @ (posedge clk) begin g55 <= g817; end
	always @ (posedge clk) begin g56 <= g819; end
	always @ (posedge clk) begin g57 <= g821; end
	always @ (posedge clk) begin g58 <= g823; end
	always @ (posedge clk) begin g60 <= g7231; end
	always @ (posedge clk) begin g61 <= g7233; end
	always @ (posedge clk) begin g63 <= g7234; end
	always @ (posedge clk) begin g66 <= g833; end
	always @ (posedge clk) begin g67 <= g835; end
	always @ (posedge clk) begin g68 <= g837; end
	always @ (posedge clk) begin g69 <= g839; end
	always @ (posedge clk) begin g71 <= g841; end
	always @ (posedge clk) begin g72 <= g843; end
	always @ (posedge clk) begin g73 <= g845; end
	always @ (posedge clk) begin g74 <= g847; end
	always @ (posedge clk) begin g76 <= g849; end
	always @ (posedge clk) begin g77 <= g851; end
	always @ (posedge clk) begin g78 <= g853; end
	always @ (posedge clk) begin g79 <= g855; end
	always @ (posedge clk) begin g81 <= g857; end
	always @ (posedge clk) begin g82 <= g859; end
	always @ (posedge clk) begin g83 <= g861; end
	always @ (posedge clk) begin g84 <= g863; end
	always @ (posedge clk) begin g87 <= g7235; end
	always @ (posedge clk) begin g89 <= g866; end
	always @ (posedge clk) begin g90 <= g868; end
	always @ (posedge clk) begin g91 <= g870; end
	always @ (posedge clk) begin g92 <= g872; end
	always @ (posedge clk) begin g94 <= g874; end
	always @ (posedge clk) begin g95 <= g876; end
	always @ (posedge clk) begin g96 <= g878; end
	always @ (posedge clk) begin g97 <= g880; end
	always @ (posedge clk) begin g99 <= g882; end
	always @ (posedge clk) begin g100 <= g884; end
	always @ (posedge clk) begin g101 <= g886; end
	always @ (posedge clk) begin g102 <= g888; end
	always @ (posedge clk) begin g104 <= g890; end
	always @ (posedge clk) begin g105 <= g892; end
	always @ (posedge clk) begin g106 <= g894; end
	always @ (posedge clk) begin g107 <= g896; end
	always @ (posedge clk) begin g110 <= g7236; end
	always @ (posedge clk) begin g112 <= g900; end
	always @ (posedge clk) begin g113 <= g902; end
	always @ (posedge clk) begin g114 <= g904; end
	always @ (posedge clk) begin g115 <= g906; end
	always @ (posedge clk) begin g117 <= g908; end
	always @ (posedge clk) begin g118 <= g910; end
	always @ (posedge clk) begin g119 <= g912; end
	always @ (posedge clk) begin g120 <= g914; end
	always @ (posedge clk) begin g122 <= g916; end
	always @ (posedge clk) begin g123 <= g918; end
	always @ (posedge clk) begin g124 <= g920; end
	always @ (posedge clk) begin g125 <= g922; end
	always @ (posedge clk) begin g127 <= g924; end
	always @ (posedge clk) begin g128 <= g926; end
	always @ (posedge clk) begin g129 <= g928; end
	always @ (posedge clk) begin g130 <= g930; end
	always @ (posedge clk) begin g133 <= g7237; end
	always @ (posedge clk) begin g135 <= g933; end
	always @ (posedge clk) begin g136 <= g935; end
	always @ (posedge clk) begin g137 <= g937; end
	always @ (posedge clk) begin g138 <= g939; end
	always @ (posedge clk) begin g140 <= g941; end
	always @ (posedge clk) begin g141 <= g943; end
	always @ (posedge clk) begin g142 <= g945; end
	always @ (posedge clk) begin g143 <= g947; end
	always @ (posedge clk) begin g145 <= g949; end
	always @ (posedge clk) begin g146 <= g951; end
	always @ (posedge clk) begin g147 <= g953; end
	always @ (posedge clk) begin g148 <= g955; end
	always @ (posedge clk) begin g150 <= g957; end
	always @ (posedge clk) begin g151 <= g959; end
	always @ (posedge clk) begin g152 <= g961; end
	always @ (posedge clk) begin g153 <= g963; end
	always @ (posedge clk) begin g156 <= g7238; end
	always @ (posedge clk) begin g158 <= g967; end
	always @ (posedge clk) begin g159 <= g969; end
	always @ (posedge clk) begin g160 <= g971; end
	always @ (posedge clk) begin g161 <= g973; end
	always @ (posedge clk) begin g163 <= g975; end
	always @ (posedge clk) begin g164 <= g977; end
	always @ (posedge clk) begin g165 <= g979; end
	always @ (posedge clk) begin g166 <= g981; end
	always @ (posedge clk) begin g168 <= g983; end
	always @ (posedge clk) begin g169 <= g985; end
	always @ (posedge clk) begin g170 <= g987; end
	always @ (posedge clk) begin g171 <= g989; end
	always @ (posedge clk) begin g173 <= g991; end
	always @ (posedge clk) begin g174 <= g993; end
	always @ (posedge clk) begin g175 <= g995; end
	always @ (posedge clk) begin g176 <= g997; end
	always @ (posedge clk) begin g179 <= g7239; end
	always @ (posedge clk) begin g181 <= g1000; end
	always @ (posedge clk) begin g182 <= g1002; end
	always @ (posedge clk) begin g183 <= g1004; end
	always @ (posedge clk) begin g184 <= g1006; end
	always @ (posedge clk) begin g186 <= g1008; end
	always @ (posedge clk) begin g187 <= g1010; end
	always @ (posedge clk) begin g188 <= g1012; end
	always @ (posedge clk) begin g189 <= g1014; end
	always @ (posedge clk) begin g191 <= g1016; end
	always @ (posedge clk) begin g192 <= g1018; end
	always @ (posedge clk) begin g193 <= g1020; end
	always @ (posedge clk) begin g194 <= g1022; end
	always @ (posedge clk) begin g196 <= g1024; end
	always @ (posedge clk) begin g197 <= g1026; end
	always @ (posedge clk) begin g198 <= g1028; end
	always @ (posedge clk) begin g199 <= g1030; end
	always @ (posedge clk) begin g202 <= g7240; end
	always @ (posedge clk) begin g204 <= g1034; end
	always @ (posedge clk) begin g205 <= g1036; end
	always @ (posedge clk) begin g206 <= g1038; end
	always @ (posedge clk) begin g207 <= g1040; end
	always @ (posedge clk) begin g209 <= g1042; end
	always @ (posedge clk) begin g210 <= g1044; end
	always @ (posedge clk) begin g211 <= g1046; end
	always @ (posedge clk) begin g212 <= g1048; end
	always @ (posedge clk) begin g214 <= g1050; end
	always @ (posedge clk) begin g215 <= g1052; end
	always @ (posedge clk) begin g216 <= g1054; end
	always @ (posedge clk) begin g217 <= g1056; end
	always @ (posedge clk) begin g219 <= g1058; end
	always @ (posedge clk) begin g220 <= g1060; end
	always @ (posedge clk) begin g221 <= g1062; end
	always @ (posedge clk) begin g222 <= g1064; end
	always @ (posedge clk) begin g225 <= g7241; end
	always @ (posedge clk) begin g227 <= g1067; end
	always @ (posedge clk) begin g228 <= g1069; end
	always @ (posedge clk) begin g229 <= g1071; end
	always @ (posedge clk) begin g230 <= g1073; end
	always @ (posedge clk) begin g232 <= g1075; end
	always @ (posedge clk) begin g233 <= g1077; end
	always @ (posedge clk) begin g234 <= g1079; end
	always @ (posedge clk) begin g235 <= g1081; end
	always @ (posedge clk) begin g237 <= g1083; end
	always @ (posedge clk) begin g238 <= g1085; end
	always @ (posedge clk) begin g239 <= g1087; end
	always @ (posedge clk) begin g240 <= g1089; end
	always @ (posedge clk) begin g242 <= g1091; end
	always @ (posedge clk) begin g243 <= g1093; end
	always @ (posedge clk) begin g244 <= g1095; end
	always @ (posedge clk) begin g245 <= g1097; end
	always @ (posedge clk) begin g248 <= g7242; end
	always @ (posedge clk) begin g250 <= g1101; end
	always @ (posedge clk) begin g251 <= g1103; end
	always @ (posedge clk) begin g252 <= g1105; end
	always @ (posedge clk) begin g253 <= g1107; end
	always @ (posedge clk) begin g255 <= g1109; end
	always @ (posedge clk) begin g256 <= g1111; end
	always @ (posedge clk) begin g257 <= g1113; end
	always @ (posedge clk) begin g258 <= g1115; end
	always @ (posedge clk) begin g260 <= g1117; end
	always @ (posedge clk) begin g261 <= g1119; end
	always @ (posedge clk) begin g262 <= g1121; end
	always @ (posedge clk) begin g263 <= g1123; end
	always @ (posedge clk) begin g265 <= g1125; end
	always @ (posedge clk) begin g266 <= g1127; end
	always @ (posedge clk) begin g267 <= g1129; end
	always @ (posedge clk) begin g268 <= g1131; end
	always @ (posedge clk) begin g271 <= g7243; end
	always @ (posedge clk) begin g273 <= g1134; end
	always @ (posedge clk) begin g274 <= g1136; end
	always @ (posedge clk) begin g275 <= g1138; end
	always @ (posedge clk) begin g276 <= g1140; end
	always @ (posedge clk) begin g278 <= g1142; end
	always @ (posedge clk) begin g279 <= g1144; end
	always @ (posedge clk) begin g280 <= g1146; end
	always @ (posedge clk) begin g281 <= g1148; end
	always @ (posedge clk) begin g283 <= g1150; end
	always @ (posedge clk) begin g284 <= g1152; end
	always @ (posedge clk) begin g285 <= g1154; end
	always @ (posedge clk) begin g286 <= g1156; end
	always @ (posedge clk) begin g288 <= g1158; end
	always @ (posedge clk) begin g289 <= g1160; end
	always @ (posedge clk) begin g290 <= g1162; end
	always @ (posedge clk) begin g291 <= g1164; end
	always @ (posedge clk) begin g294 <= g7244; end
	always @ (posedge clk) begin g296 <= g1168; end
	always @ (posedge clk) begin g297 <= g1170; end
	always @ (posedge clk) begin g298 <= g1172; end
	always @ (posedge clk) begin g299 <= g1174; end
	always @ (posedge clk) begin g301 <= g1176; end
	always @ (posedge clk) begin g302 <= g1178; end
	always @ (posedge clk) begin g303 <= g1180; end
	always @ (posedge clk) begin g304 <= g1182; end
	always @ (posedge clk) begin g306 <= g1184; end
	always @ (posedge clk) begin g307 <= g1186; end
	always @ (posedge clk) begin g308 <= g1188; end
	always @ (posedge clk) begin g309 <= g1190; end
	always @ (posedge clk) begin g311 <= g1192; end
	always @ (posedge clk) begin g312 <= g1194; end
	always @ (posedge clk) begin g313 <= g1196; end
	always @ (posedge clk) begin g314 <= g1198; end
	always @ (posedge clk) begin g317 <= g7245; end
	always @ (posedge clk) begin g319 <= g1205; end
	always @ (posedge clk) begin g320 <= g1207; end
	always @ (posedge clk) begin g321 <= g1209; end
	always @ (posedge clk) begin g322 <= g1211; end
	always @ (posedge clk) begin g324 <= g1213; end
	always @ (posedge clk) begin g325 <= g1215; end
	always @ (posedge clk) begin g326 <= g1217; end
	always @ (posedge clk) begin g327 <= g1219; end
	always @ (posedge clk) begin g329 <= g1221; end
	always @ (posedge clk) begin g330 <= g1223; end
	always @ (posedge clk) begin g331 <= g1225; end
	always @ (posedge clk) begin g332 <= g1227; end
	always @ (posedge clk) begin g334 <= g1229; end
	always @ (posedge clk) begin g335 <= g1231; end
	always @ (posedge clk) begin g336 <= g1233; end
	always @ (posedge clk) begin g337 <= g1235; end
	always @ (posedge clk) begin g340 <= g7246; end
	always @ (posedge clk) begin g342 <= g1238; end
	always @ (posedge clk) begin g343 <= g1240; end
	always @ (posedge clk) begin g344 <= g1242; end
	always @ (posedge clk) begin g345 <= g1244; end
	always @ (posedge clk) begin g347 <= g1246; end
	always @ (posedge clk) begin g348 <= g1248; end
	always @ (posedge clk) begin g349 <= g1250; end
	always @ (posedge clk) begin g350 <= g1252; end
	always @ (posedge clk) begin g352 <= g1254; end
	always @ (posedge clk) begin g353 <= g1256; end
	always @ (posedge clk) begin g354 <= g1258; end
	always @ (posedge clk) begin g355 <= g1260; end
	always @ (posedge clk) begin g357 <= g1262; end
	always @ (posedge clk) begin g358 <= g1264; end
	always @ (posedge clk) begin g359 <= g1266; end
	always @ (posedge clk) begin g360 <= g1268; end
	always @ (posedge clk) begin g363 <= g7247; end
	always @ (posedge clk) begin g365 <= g1272; end
	always @ (posedge clk) begin g366 <= g1274; end
	always @ (posedge clk) begin g367 <= g1276; end
	always @ (posedge clk) begin g368 <= g1278; end
	always @ (posedge clk) begin g370 <= g1280; end
	always @ (posedge clk) begin g371 <= g1282; end
	always @ (posedge clk) begin g372 <= g1284; end
	always @ (posedge clk) begin g373 <= g1286; end
	always @ (posedge clk) begin g375 <= g1288; end
	always @ (posedge clk) begin g376 <= g1290; end
	always @ (posedge clk) begin g377 <= g1292; end
	always @ (posedge clk) begin g378 <= g1294; end
	always @ (posedge clk) begin g380 <= g1296; end
	always @ (posedge clk) begin g381 <= g1298; end
	always @ (posedge clk) begin g382 <= g1300; end
	always @ (posedge clk) begin g383 <= g1302; end
	always @ (posedge clk) begin g386 <= g7248; end
	always @ (posedge clk) begin g388 <= g1306; end
	always @ (posedge clk) begin g389 <= g1308; end
	always @ (posedge clk) begin g390 <= g1310; end
	always @ (posedge clk) begin g391 <= g1312; end
	always @ (posedge clk) begin g393 <= g1314; end
	always @ (posedge clk) begin g394 <= g1316; end
	always @ (posedge clk) begin g395 <= g1318; end
	always @ (posedge clk) begin g396 <= g1320; end
	always @ (posedge clk) begin g398 <= g1322; end
	always @ (posedge clk) begin g399 <= g1324; end
	always @ (posedge clk) begin g400 <= g1326; end
	always @ (posedge clk) begin g401 <= g1328; end
	always @ (posedge clk) begin g403 <= g1330; end
	always @ (posedge clk) begin g404 <= g1332; end
	always @ (posedge clk) begin g405 <= g1334; end
	always @ (posedge clk) begin g406 <= g1336; end
	always @ (posedge clk) begin g409 <= g7249; end
	always @ (posedge clk) begin g411 <= g1339; end
	always @ (posedge clk) begin g412 <= g1341; end
	always @ (posedge clk) begin g413 <= g1343; end
	always @ (posedge clk) begin g414 <= g1345; end
	always @ (posedge clk) begin g416 <= g1347; end
	always @ (posedge clk) begin g417 <= g1349; end
	always @ (posedge clk) begin g418 <= g1351; end
	always @ (posedge clk) begin g419 <= g1353; end
	always @ (posedge clk) begin g421 <= g1355; end
	always @ (posedge clk) begin g422 <= g1357; end
	always @ (posedge clk) begin g423 <= g1359; end
	always @ (posedge clk) begin g424 <= g1361; end
	always @ (posedge clk) begin g426 <= g1363; end
	always @ (posedge clk) begin g427 <= g1365; end
	always @ (posedge clk) begin g428 <= g1367; end
	always @ (posedge clk) begin g429 <= g1369; end
	always @ (posedge clk) begin g432 <= g7250; end
	always @ (posedge clk) begin g434 <= g1375; end
	always @ (posedge clk) begin g435 <= g1377; end
	always @ (posedge clk) begin g436 <= g1379; end
	always @ (posedge clk) begin g437 <= g1381; end
	always @ (posedge clk) begin g439 <= g1383; end
	always @ (posedge clk) begin g440 <= g1385; end
	always @ (posedge clk) begin g441 <= g1387; end
	always @ (posedge clk) begin g442 <= g1389; end
	always @ (posedge clk) begin g444 <= g1391; end
	always @ (posedge clk) begin g445 <= g1393; end
	always @ (posedge clk) begin g446 <= g1395; end
	always @ (posedge clk) begin g447 <= g1397; end
	always @ (posedge clk) begin g449 <= g1399; end
	always @ (posedge clk) begin g450 <= g1401; end
	always @ (posedge clk) begin g451 <= g1403; end
	always @ (posedge clk) begin g452 <= g1405; end
	always @ (posedge clk) begin g455 <= g7251; end
	always @ (posedge clk) begin g457 <= g1408; end
	always @ (posedge clk) begin g458 <= g1410; end
	always @ (posedge clk) begin g459 <= g1412; end
	always @ (posedge clk) begin g460 <= g1414; end
	always @ (posedge clk) begin g462 <= g1416; end
	always @ (posedge clk) begin g463 <= g1418; end
	always @ (posedge clk) begin g464 <= g1420; end
	always @ (posedge clk) begin g465 <= g1422; end
	always @ (posedge clk) begin g467 <= g1424; end
	always @ (posedge clk) begin g468 <= g1426; end
	always @ (posedge clk) begin g469 <= g1428; end
	always @ (posedge clk) begin g470 <= g1430; end
	always @ (posedge clk) begin g472 <= g1432; end
	always @ (posedge clk) begin g473 <= g1434; end
	always @ (posedge clk) begin g474 <= g1436; end
	always @ (posedge clk) begin g475 <= g1438; end
	always @ (posedge clk) begin g478 <= g7252; end
	always @ (posedge clk) begin g480 <= g1442; end
	always @ (posedge clk) begin g481 <= g1444; end
	always @ (posedge clk) begin g482 <= g1446; end
	always @ (posedge clk) begin g483 <= g1448; end
	always @ (posedge clk) begin g485 <= g1450; end
	always @ (posedge clk) begin g486 <= g1452; end
	always @ (posedge clk) begin g487 <= g1454; end
	always @ (posedge clk) begin g488 <= g1456; end
	always @ (posedge clk) begin g490 <= g1458; end
	always @ (posedge clk) begin g491 <= g1460; end
	always @ (posedge clk) begin g492 <= g1462; end
	always @ (posedge clk) begin g493 <= g1464; end
	always @ (posedge clk) begin g495 <= g1466; end
	always @ (posedge clk) begin g496 <= g1468; end
	always @ (posedge clk) begin g497 <= g1470; end
	always @ (posedge clk) begin g498 <= g1472; end
	always @ (posedge clk) begin g501 <= g7253; end
	always @ (posedge clk) begin g503 <= g1476; end
	always @ (posedge clk) begin g504 <= g1478; end
	always @ (posedge clk) begin g505 <= g1480; end
	always @ (posedge clk) begin g506 <= g1482; end
	always @ (posedge clk) begin g508 <= g1484; end
	always @ (posedge clk) begin g509 <= g1486; end
	always @ (posedge clk) begin g510 <= g1488; end
	always @ (posedge clk) begin g511 <= g1490; end
	always @ (posedge clk) begin g513 <= g1492; end
	always @ (posedge clk) begin g514 <= g1494; end
	always @ (posedge clk) begin g515 <= g1496; end
	always @ (posedge clk) begin g516 <= g1498; end
	always @ (posedge clk) begin g518 <= g1500; end
	always @ (posedge clk) begin g519 <= g1502; end
	always @ (posedge clk) begin g520 <= g1504; end
	always @ (posedge clk) begin g521 <= g1506; end
	always @ (posedge clk) begin g524 <= g7254; end
	always @ (posedge clk) begin g526 <= g1509; end
	always @ (posedge clk) begin g527 <= g1511; end
	always @ (posedge clk) begin g528 <= g1513; end
	always @ (posedge clk) begin g529 <= g1515; end
	always @ (posedge clk) begin g531 <= g1517; end
	always @ (posedge clk) begin g532 <= g1519; end
	always @ (posedge clk) begin g533 <= g1521; end
	always @ (posedge clk) begin g534 <= g1523; end
	always @ (posedge clk) begin g536 <= g1525; end
	always @ (posedge clk) begin g537 <= g1527; end
	always @ (posedge clk) begin g538 <= g1529; end
	always @ (posedge clk) begin g539 <= g1531; end
	always @ (posedge clk) begin g541 <= g1533; end
	always @ (posedge clk) begin g542 <= g1535; end
	always @ (posedge clk) begin g543 <= g1537; end
	always @ (posedge clk) begin g544 <= g1539; end
	always @ (posedge clk) begin g547 <= g7255; end
	always @ (posedge clk) begin g549 <= g1546; end
	always @ (posedge clk) begin g550 <= g1548; end
	always @ (posedge clk) begin g551 <= g1550; end
	always @ (posedge clk) begin g552 <= g1552; end
	always @ (posedge clk) begin g554 <= g1554; end
	always @ (posedge clk) begin g555 <= g1556; end
	always @ (posedge clk) begin g556 <= g1558; end
	always @ (posedge clk) begin g557 <= g1560; end
	always @ (posedge clk) begin g559 <= g1562; end
	always @ (posedge clk) begin g560 <= g1564; end
	always @ (posedge clk) begin g561 <= g1566; end
	always @ (posedge clk) begin g562 <= g1568; end
	always @ (posedge clk) begin g564 <= g1570; end
	always @ (posedge clk) begin g565 <= g1572; end
	always @ (posedge clk) begin g566 <= g1574; end
	always @ (posedge clk) begin g567 <= g1576; end
	always @ (posedge clk) begin g570 <= g7256; end
	always @ (posedge clk) begin g572 <= g1579; end
	always @ (posedge clk) begin g573 <= g1581; end
	always @ (posedge clk) begin g574 <= g1583; end
	always @ (posedge clk) begin g575 <= g1585; end
	always @ (posedge clk) begin g577 <= g1587; end
	always @ (posedge clk) begin g578 <= g1589; end
	always @ (posedge clk) begin g579 <= g1591; end
	always @ (posedge clk) begin g580 <= g1593; end
	always @ (posedge clk) begin g582 <= g1595; end
	always @ (posedge clk) begin g583 <= g1597; end
	always @ (posedge clk) begin g584 <= g1599; end
	always @ (posedge clk) begin g585 <= g1601; end
	always @ (posedge clk) begin g587 <= g1603; end
	always @ (posedge clk) begin g588 <= g1605; end
	always @ (posedge clk) begin g589 <= g1607; end
	always @ (posedge clk) begin g590 <= g1609; end
	always @ (posedge clk) begin g593 <= g7257; end
	always @ (posedge clk) begin g595 <= g1613; end
	always @ (posedge clk) begin g596 <= g1615; end
	always @ (posedge clk) begin g597 <= g1617; end
	always @ (posedge clk) begin g598 <= g1619; end
	always @ (posedge clk) begin g600 <= g1621; end
	always @ (posedge clk) begin g601 <= g1623; end
	always @ (posedge clk) begin g602 <= g1625; end
	always @ (posedge clk) begin g603 <= g1627; end
	always @ (posedge clk) begin g605 <= g1629; end
	always @ (posedge clk) begin g606 <= g1631; end
	always @ (posedge clk) begin g607 <= g1633; end
	always @ (posedge clk) begin g608 <= g1635; end
	always @ (posedge clk) begin g610 <= g1637; end
	always @ (posedge clk) begin g611 <= g1639; end
	always @ (posedge clk) begin g612 <= g1641; end
	always @ (posedge clk) begin g613 <= g1643; end
	always @ (posedge clk) begin g616 <= g7258; end
	always @ (posedge clk) begin g618 <= g1646; end
	always @ (posedge clk) begin g619 <= g1648; end
	always @ (posedge clk) begin g620 <= g1650; end
	always @ (posedge clk) begin g621 <= g1652; end
	always @ (posedge clk) begin g623 <= g1654; end
	always @ (posedge clk) begin g624 <= g1656; end
	always @ (posedge clk) begin g625 <= g1658; end
	always @ (posedge clk) begin g626 <= g1660; end
	always @ (posedge clk) begin g628 <= g1662; end
	always @ (posedge clk) begin g629 <= g1664; end
	always @ (posedge clk) begin g630 <= g1666; end
	always @ (posedge clk) begin g631 <= g1668; end
	always @ (posedge clk) begin g633 <= g1670; end
	always @ (posedge clk) begin g634 <= g1672; end
	always @ (posedge clk) begin g635 <= g1674; end
	always @ (posedge clk) begin g636 <= g1676; end
	always @ (posedge clk) begin g639 <= g7259; end
	always @ (posedge clk) begin g641 <= g1680; end
	always @ (posedge clk) begin g642 <= g1682; end
	always @ (posedge clk) begin g643 <= g1684; end
	always @ (posedge clk) begin g644 <= g1686; end
	always @ (posedge clk) begin g646 <= g1688; end
	always @ (posedge clk) begin g647 <= g1690; end
	always @ (posedge clk) begin g648 <= g1692; end
	always @ (posedge clk) begin g649 <= g1694; end
	always @ (posedge clk) begin g651 <= g1696; end
	always @ (posedge clk) begin g652 <= g1698; end
	always @ (posedge clk) begin g653 <= g1700; end
	always @ (posedge clk) begin g654 <= g1702; end
	always @ (posedge clk) begin g656 <= g1704; end
	always @ (posedge clk) begin g657 <= g1706; end
	always @ (posedge clk) begin g658 <= g1708; end
	always @ (posedge clk) begin g659 <= g1710; end
	always @ (posedge clk) begin g662 <= g7260; end
	always @ (posedge clk) begin g664 <= g1713; end
	always @ (posedge clk) begin g665 <= g1715; end
	always @ (posedge clk) begin g666 <= g1717; end
	always @ (posedge clk) begin g667 <= g1719; end
	always @ (posedge clk) begin g669 <= g1721; end
	always @ (posedge clk) begin g670 <= g1723; end
	always @ (posedge clk) begin g671 <= g1725; end
	always @ (posedge clk) begin g672 <= g1727; end
	always @ (posedge clk) begin g674 <= g1729; end
	always @ (posedge clk) begin g675 <= g1731; end
	always @ (posedge clk) begin g676 <= g1733; end
	always @ (posedge clk) begin g677 <= g1735; end
	always @ (posedge clk) begin g679 <= g1737; end
	always @ (posedge clk) begin g680 <= g1739; end
	always @ (posedge clk) begin g681 <= g1741; end
	always @ (posedge clk) begin g682 <= g1743; end
	always @ (posedge clk) begin g685 <= g7261; end
	always @ (posedge clk) begin g687 <= g1747; end
	always @ (posedge clk) begin g688 <= g1749; end
	always @ (posedge clk) begin g689 <= g1751; end
	always @ (posedge clk) begin g690 <= g1753; end
	always @ (posedge clk) begin g692 <= g1755; end
	always @ (posedge clk) begin g693 <= g1757; end
	always @ (posedge clk) begin g694 <= g1759; end
	always @ (posedge clk) begin g695 <= g1761; end
	always @ (posedge clk) begin g697 <= g1763; end
	always @ (posedge clk) begin g698 <= g1765; end
	always @ (posedge clk) begin g699 <= g1767; end
	always @ (posedge clk) begin g700 <= g1769; end
	always @ (posedge clk) begin g702 <= g1771; end
	always @ (posedge clk) begin g703 <= g1773; end
	always @ (posedge clk) begin g704 <= g1775; end
	always @ (posedge clk) begin g705 <= g1777; end
	always @ (posedge clk) begin g708 <= g7262; end
	always @ (posedge clk) begin g710 <= g1783; end
	always @ (posedge clk) begin g711 <= g1785; end
	always @ (posedge clk) begin g712 <= g1787; end
	always @ (posedge clk) begin g713 <= g1789; end
	always @ (posedge clk) begin g715 <= g1791; end
	always @ (posedge clk) begin g716 <= g1793; end
	always @ (posedge clk) begin g717 <= g1795; end
	always @ (posedge clk) begin g718 <= g1797; end
	always @ (posedge clk) begin g720 <= g1799; end
	always @ (posedge clk) begin g721 <= g1801; end
	always @ (posedge clk) begin g722 <= g1803; end
	always @ (posedge clk) begin g723 <= g1805; end
	always @ (posedge clk) begin g725 <= g1807; end
	always @ (posedge clk) begin g726 <= g1809; end
	always @ (posedge clk) begin g727 <= g1811; end
	always @ (posedge clk) begin g728 <= g1813; end
	always @ (posedge clk) begin g731 <= g7263; end
	always @ (posedge clk) begin g733 <= g1816; end
	always @ (posedge clk) begin g734 <= g1818; end
	always @ (posedge clk) begin g735 <= g1820; end
	always @ (posedge clk) begin g736 <= g1822; end
	always @ (posedge clk) begin g738 <= g1824; end
	always @ (posedge clk) begin g739 <= g1826; end
	always @ (posedge clk) begin g740 <= g1828; end
	always @ (posedge clk) begin g741 <= g1830; end
	always @ (posedge clk) begin g743 <= g1832; end
	always @ (posedge clk) begin g744 <= g1834; end
	always @ (posedge clk) begin g745 <= g1836; end
	always @ (posedge clk) begin g746 <= g1838; end
	always @ (posedge clk) begin g748 <= g1840; end
	always @ (posedge clk) begin g749 <= g1842; end
	always @ (posedge clk) begin g750 <= g1844; end
	always @ (posedge clk) begin g751 <= g1846; end
	always @ (posedge clk) begin g754 <= g7264; end
	always @ (posedge clk) begin g756 <= g1850; end
	always @ (posedge clk) begin g757 <= g1852; end
	always @ (posedge clk) begin g758 <= g1854; end
	always @ (posedge clk) begin g759 <= g1856; end
	always @ (posedge clk) begin g761 <= g1858; end
	always @ (posedge clk) begin g762 <= g1860; end
	always @ (posedge clk) begin g763 <= g1862; end
	always @ (posedge clk) begin g764 <= g1864; end
	always @ (posedge clk) begin g766 <= g1866; end
	always @ (posedge clk) begin g767 <= g1868; end
	always @ (posedge clk) begin g768 <= g1870; end
	always @ (posedge clk) begin g769 <= g1872; end
	always @ (posedge clk) begin g771 <= g1874; end
	always @ (posedge clk) begin g772 <= g1876; end
	always @ (posedge clk) begin g773 <= g1878; end
	always @ (posedge clk) begin g774 <= g1880; end
	always @ (posedge clk) begin g777 <= g7265; end
	always @ (posedge clk) begin g779 <= g1883; end
	always @ (posedge clk) begin g790 <= g7266; end
	always @ (posedge clk) begin g792 <= g7267; end
	always @ (posedge clk) begin g794 <= g7268; end
	always @ (posedge clk) begin g800 <= g7269; end
	always @ (posedge clk) begin g802 <= g7270; end
	always @ (posedge clk) begin g804 <= g7271; end
	always @ (posedge clk) begin g806 <= g7272; end
	always @ (posedge clk) begin g808 <= g7273; end
	always @ (posedge clk) begin g810 <= g7274; end
	always @ (posedge clk) begin g812 <= g7275; end
	always @ (posedge clk) begin g814 <= g7276; end
	always @ (posedge clk) begin g816 <= g7277; end
	always @ (posedge clk) begin g818 <= g7278; end
	always @ (posedge clk) begin g820 <= g7279; end
	always @ (posedge clk) begin g822 <= g7280; end
	always @ (posedge clk) begin g827 <= g7281; end
	always @ (posedge clk) begin g828 <= g7282; end
	always @ (posedge clk) begin g830 <= g2018; end
	always @ (posedge clk) begin g831 <= g2020; end
	always @ (posedge clk) begin g834 <= g7283; end
	always @ (posedge clk) begin g836 <= g7284; end
	always @ (posedge clk) begin g838 <= g7285; end
	always @ (posedge clk) begin g840 <= g7286; end
	always @ (posedge clk) begin g842 <= g7287; end
	always @ (posedge clk) begin g844 <= g7288; end
	always @ (posedge clk) begin g846 <= g7289; end
	always @ (posedge clk) begin g848 <= g7290; end
	always @ (posedge clk) begin g850 <= g7291; end
	always @ (posedge clk) begin g852 <= g7292; end
	always @ (posedge clk) begin g854 <= g7293; end
	always @ (posedge clk) begin g856 <= g7294; end
	always @ (posedge clk) begin g858 <= g7295; end
	always @ (posedge clk) begin g860 <= g7296; end
	always @ (posedge clk) begin g862 <= g7297; end
	always @ (posedge clk) begin g864 <= g7298; end
	always @ (posedge clk) begin g867 <= g7299; end
	always @ (posedge clk) begin g869 <= g7300; end
	always @ (posedge clk) begin g871 <= g7301; end
	always @ (posedge clk) begin g873 <= g7302; end
	always @ (posedge clk) begin g875 <= g7303; end
	always @ (posedge clk) begin g877 <= g7304; end
	always @ (posedge clk) begin g879 <= g7305; end
	always @ (posedge clk) begin g881 <= g7306; end
	always @ (posedge clk) begin g883 <= g7307; end
	always @ (posedge clk) begin g885 <= g7308; end
	always @ (posedge clk) begin g887 <= g7309; end
	always @ (posedge clk) begin g889 <= g7310; end
	always @ (posedge clk) begin g891 <= g7311; end
	always @ (posedge clk) begin g893 <= g7312; end
	always @ (posedge clk) begin g895 <= g7313; end
	always @ (posedge clk) begin g897 <= g7314; end
	always @ (posedge clk) begin g901 <= g7315; end
	always @ (posedge clk) begin g903 <= g7316; end
	always @ (posedge clk) begin g905 <= g7317; end
	always @ (posedge clk) begin g907 <= g7318; end
	always @ (posedge clk) begin g909 <= g7319; end
	always @ (posedge clk) begin g911 <= g7320; end
	always @ (posedge clk) begin g913 <= g7321; end
	always @ (posedge clk) begin g915 <= g7322; end
	always @ (posedge clk) begin g917 <= g7323; end
	always @ (posedge clk) begin g919 <= g7324; end
	always @ (posedge clk) begin g921 <= g7325; end
	always @ (posedge clk) begin g923 <= g7326; end
	always @ (posedge clk) begin g925 <= g7327; end
	always @ (posedge clk) begin g927 <= g7328; end
	always @ (posedge clk) begin g929 <= g7329; end
	always @ (posedge clk) begin g931 <= g7330; end
	always @ (posedge clk) begin g934 <= g7331; end
	always @ (posedge clk) begin g936 <= g7332; end
	always @ (posedge clk) begin g938 <= g7333; end
	always @ (posedge clk) begin g940 <= g7334; end
	always @ (posedge clk) begin g942 <= g7335; end
	always @ (posedge clk) begin g944 <= g7336; end
	always @ (posedge clk) begin g946 <= g7337; end
	always @ (posedge clk) begin g948 <= g7338; end
	always @ (posedge clk) begin g950 <= g7339; end
	always @ (posedge clk) begin g952 <= g7340; end
	always @ (posedge clk) begin g954 <= g7341; end
	always @ (posedge clk) begin g956 <= g7342; end
	always @ (posedge clk) begin g958 <= g7343; end
	always @ (posedge clk) begin g960 <= g7344; end
	always @ (posedge clk) begin g962 <= g7345; end
	always @ (posedge clk) begin g964 <= g7346; end
	always @ (posedge clk) begin g968 <= g7347; end
	always @ (posedge clk) begin g970 <= g7348; end
	always @ (posedge clk) begin g972 <= g7349; end
	always @ (posedge clk) begin g974 <= g7350; end
	always @ (posedge clk) begin g976 <= g7351; end
	always @ (posedge clk) begin g978 <= g7352; end
	always @ (posedge clk) begin g980 <= g7353; end
	always @ (posedge clk) begin g982 <= g7354; end
	always @ (posedge clk) begin g984 <= g7355; end
	always @ (posedge clk) begin g986 <= g7356; end
	always @ (posedge clk) begin g988 <= g7357; end
	always @ (posedge clk) begin g990 <= g7358; end
	always @ (posedge clk) begin g992 <= g7359; end
	always @ (posedge clk) begin g994 <= g7360; end
	always @ (posedge clk) begin g996 <= g7361; end
	always @ (posedge clk) begin g998 <= g7362; end
	always @ (posedge clk) begin g1001 <= g7363; end
	always @ (posedge clk) begin g1003 <= g7364; end
	always @ (posedge clk) begin g1005 <= g7365; end
	always @ (posedge clk) begin g1007 <= g7366; end
	always @ (posedge clk) begin g1009 <= g7367; end
	always @ (posedge clk) begin g1011 <= g7368; end
	always @ (posedge clk) begin g1013 <= g7369; end
	always @ (posedge clk) begin g1015 <= g7370; end
	always @ (posedge clk) begin g1017 <= g7371; end
	always @ (posedge clk) begin g1019 <= g7372; end
	always @ (posedge clk) begin g1021 <= g7373; end
	always @ (posedge clk) begin g1023 <= g7374; end
	always @ (posedge clk) begin g1025 <= g7375; end
	always @ (posedge clk) begin g1027 <= g7376; end
	always @ (posedge clk) begin g1029 <= g7377; end
	always @ (posedge clk) begin g1031 <= g7378; end
	always @ (posedge clk) begin g1035 <= g7379; end
	always @ (posedge clk) begin g1037 <= g7380; end
	always @ (posedge clk) begin g1039 <= g7381; end
	always @ (posedge clk) begin g1041 <= g7382; end
	always @ (posedge clk) begin g1043 <= g7383; end
	always @ (posedge clk) begin g1045 <= g7384; end
	always @ (posedge clk) begin g1047 <= g7385; end
	always @ (posedge clk) begin g1049 <= g7386; end
	always @ (posedge clk) begin g1051 <= g7387; end
	always @ (posedge clk) begin g1053 <= g7388; end
	always @ (posedge clk) begin g1055 <= g7389; end
	always @ (posedge clk) begin g1057 <= g7390; end
	always @ (posedge clk) begin g1059 <= g7391; end
	always @ (posedge clk) begin g1061 <= g7392; end
	always @ (posedge clk) begin g1063 <= g7393; end
	always @ (posedge clk) begin g1065 <= g7394; end
	always @ (posedge clk) begin g1068 <= g7395; end
	always @ (posedge clk) begin g1070 <= g7396; end
	always @ (posedge clk) begin g1072 <= g7397; end
	always @ (posedge clk) begin g1074 <= g7398; end
	always @ (posedge clk) begin g1076 <= g7399; end
	always @ (posedge clk) begin g1078 <= g7400; end
	always @ (posedge clk) begin g1080 <= g7401; end
	always @ (posedge clk) begin g1082 <= g7402; end
	always @ (posedge clk) begin g1084 <= g7403; end
	always @ (posedge clk) begin g1086 <= g7404; end
	always @ (posedge clk) begin g1088 <= g7405; end
	always @ (posedge clk) begin g1090 <= g7406; end
	always @ (posedge clk) begin g1092 <= g7407; end
	always @ (posedge clk) begin g1094 <= g7408; end
	always @ (posedge clk) begin g1096 <= g7409; end
	always @ (posedge clk) begin g1098 <= g7410; end
	always @ (posedge clk) begin g1102 <= g7411; end
	always @ (posedge clk) begin g1104 <= g7412; end
	always @ (posedge clk) begin g1106 <= g7413; end
	always @ (posedge clk) begin g1108 <= g7414; end
	always @ (posedge clk) begin g1110 <= g7415; end
	always @ (posedge clk) begin g1112 <= g7416; end
	always @ (posedge clk) begin g1114 <= g7417; end
	always @ (posedge clk) begin g1116 <= g7418; end
	always @ (posedge clk) begin g1118 <= g7419; end
	always @ (posedge clk) begin g1120 <= g7420; end
	always @ (posedge clk) begin g1122 <= g7421; end
	always @ (posedge clk) begin g1124 <= g7422; end
	always @ (posedge clk) begin g1126 <= g7423; end
	always @ (posedge clk) begin g1128 <= g7424; end
	always @ (posedge clk) begin g1130 <= g7425; end
	always @ (posedge clk) begin g1132 <= g7426; end
	always @ (posedge clk) begin g1135 <= g7427; end
	always @ (posedge clk) begin g1137 <= g7428; end
	always @ (posedge clk) begin g1139 <= g7429; end
	always @ (posedge clk) begin g1141 <= g7430; end
	always @ (posedge clk) begin g1143 <= g7431; end
	always @ (posedge clk) begin g1145 <= g7432; end
	always @ (posedge clk) begin g1147 <= g7433; end
	always @ (posedge clk) begin g1149 <= g7434; end
	always @ (posedge clk) begin g1151 <= g7435; end
	always @ (posedge clk) begin g1153 <= g7436; end
	always @ (posedge clk) begin g1155 <= g7437; end
	always @ (posedge clk) begin g1157 <= g7438; end
	always @ (posedge clk) begin g1159 <= g7439; end
	always @ (posedge clk) begin g1161 <= g7440; end
	always @ (posedge clk) begin g1163 <= g7441; end
	always @ (posedge clk) begin g1165 <= g7442; end
	always @ (posedge clk) begin g1169 <= g7443; end
	always @ (posedge clk) begin g1171 <= g7444; end
	always @ (posedge clk) begin g1173 <= g7445; end
	always @ (posedge clk) begin g1175 <= g7446; end
	always @ (posedge clk) begin g1177 <= g7447; end
	always @ (posedge clk) begin g1179 <= g7448; end
	always @ (posedge clk) begin g1181 <= g7449; end
	always @ (posedge clk) begin g1183 <= g7450; end
	always @ (posedge clk) begin g1185 <= g7451; end
	always @ (posedge clk) begin g1187 <= g7452; end
	always @ (posedge clk) begin g1189 <= g7453; end
	always @ (posedge clk) begin g1191 <= g7454; end
	always @ (posedge clk) begin g1193 <= g7455; end
	always @ (posedge clk) begin g1195 <= g7456; end
	always @ (posedge clk) begin g1197 <= g7457; end
	always @ (posedge clk) begin g1199 <= g7458; end
	always @ (posedge clk) begin g1206 <= g7459; end
	always @ (posedge clk) begin g1208 <= g7460; end
	always @ (posedge clk) begin g1210 <= g7461; end
	always @ (posedge clk) begin g1212 <= g7462; end
	always @ (posedge clk) begin g1214 <= g7463; end
	always @ (posedge clk) begin g1216 <= g7464; end
	always @ (posedge clk) begin g1218 <= g7465; end
	always @ (posedge clk) begin g1220 <= g7466; end
	always @ (posedge clk) begin g1222 <= g7467; end
	always @ (posedge clk) begin g1224 <= g7468; end
	always @ (posedge clk) begin g1226 <= g7469; end
	always @ (posedge clk) begin g1228 <= g7470; end
	always @ (posedge clk) begin g1230 <= g7471; end
	always @ (posedge clk) begin g1232 <= g7472; end
	always @ (posedge clk) begin g1234 <= g7473; end
	always @ (posedge clk) begin g1236 <= g7474; end
	always @ (posedge clk) begin g1239 <= g7475; end
	always @ (posedge clk) begin g1241 <= g7476; end
	always @ (posedge clk) begin g1243 <= g7477; end
	always @ (posedge clk) begin g1245 <= g7478; end
	always @ (posedge clk) begin g1247 <= g7479; end
	always @ (posedge clk) begin g1249 <= g7480; end
	always @ (posedge clk) begin g1251 <= g7481; end
	always @ (posedge clk) begin g1253 <= g7482; end
	always @ (posedge clk) begin g1255 <= g7483; end
	always @ (posedge clk) begin g1257 <= g7484; end
	always @ (posedge clk) begin g1259 <= g7485; end
	always @ (posedge clk) begin g1261 <= g7486; end
	always @ (posedge clk) begin g1263 <= g7487; end
	always @ (posedge clk) begin g1265 <= g7488; end
	always @ (posedge clk) begin g1267 <= g7489; end
	always @ (posedge clk) begin g1269 <= g7490; end
	always @ (posedge clk) begin g1273 <= g7491; end
	always @ (posedge clk) begin g1275 <= g7492; end
	always @ (posedge clk) begin g1277 <= g7493; end
	always @ (posedge clk) begin g1279 <= g7494; end
	always @ (posedge clk) begin g1281 <= g7495; end
	always @ (posedge clk) begin g1283 <= g7496; end
	always @ (posedge clk) begin g1285 <= g7497; end
	always @ (posedge clk) begin g1287 <= g7498; end
	always @ (posedge clk) begin g1289 <= g7499; end
	always @ (posedge clk) begin g1291 <= g7500; end
	always @ (posedge clk) begin g1293 <= g7501; end
	always @ (posedge clk) begin g1295 <= g7502; end
	always @ (posedge clk) begin g1297 <= g7503; end
	always @ (posedge clk) begin g1299 <= g7504; end
	always @ (posedge clk) begin g1301 <= g7505; end
	always @ (posedge clk) begin g1303 <= g7506; end
	always @ (posedge clk) begin g1307 <= g7507; end
	always @ (posedge clk) begin g1309 <= g7508; end
	always @ (posedge clk) begin g1311 <= g7509; end
	always @ (posedge clk) begin g1313 <= g7510; end
	always @ (posedge clk) begin g1315 <= g7511; end
	always @ (posedge clk) begin g1317 <= g7512; end
	always @ (posedge clk) begin g1319 <= g7513; end
	always @ (posedge clk) begin g1321 <= g7514; end
	always @ (posedge clk) begin g1323 <= g7515; end
	always @ (posedge clk) begin g1325 <= g7516; end
	always @ (posedge clk) begin g1327 <= g7517; end
	always @ (posedge clk) begin g1329 <= g7518; end
	always @ (posedge clk) begin g1331 <= g7519; end
	always @ (posedge clk) begin g1333 <= g7520; end
	always @ (posedge clk) begin g1335 <= g7521; end
	always @ (posedge clk) begin g1337 <= g7522; end
	always @ (posedge clk) begin g1340 <= g7523; end
	always @ (posedge clk) begin g1342 <= g7524; end
	always @ (posedge clk) begin g1344 <= g7525; end
	always @ (posedge clk) begin g1346 <= g7526; end
	always @ (posedge clk) begin g1348 <= g7527; end
	always @ (posedge clk) begin g1350 <= g7528; end
	always @ (posedge clk) begin g1352 <= g7529; end
	always @ (posedge clk) begin g1354 <= g7530; end
	always @ (posedge clk) begin g1356 <= g7531; end
	always @ (posedge clk) begin g1358 <= g7532; end
	always @ (posedge clk) begin g1360 <= g7533; end
	always @ (posedge clk) begin g1362 <= g7534; end
	always @ (posedge clk) begin g1364 <= g7535; end
	always @ (posedge clk) begin g1366 <= g7536; end
	always @ (posedge clk) begin g1368 <= g7537; end
	always @ (posedge clk) begin g1370 <= g7538; end
	always @ (posedge clk) begin g1376 <= g7539; end
	always @ (posedge clk) begin g1378 <= g7540; end
	always @ (posedge clk) begin g1380 <= g7541; end
	always @ (posedge clk) begin g1382 <= g7542; end
	always @ (posedge clk) begin g1384 <= g7543; end
	always @ (posedge clk) begin g1386 <= g7544; end
	always @ (posedge clk) begin g1388 <= g7545; end
	always @ (posedge clk) begin g1390 <= g7546; end
	always @ (posedge clk) begin g1392 <= g7547; end
	always @ (posedge clk) begin g1394 <= g7548; end
	always @ (posedge clk) begin g1396 <= g7549; end
	always @ (posedge clk) begin g1398 <= g7550; end
	always @ (posedge clk) begin g1400 <= g7551; end
	always @ (posedge clk) begin g1402 <= g7552; end
	always @ (posedge clk) begin g1404 <= g7553; end
	always @ (posedge clk) begin g1406 <= g7554; end
	always @ (posedge clk) begin g1409 <= g7555; end
	always @ (posedge clk) begin g1411 <= g7556; end
	always @ (posedge clk) begin g1413 <= g7557; end
	always @ (posedge clk) begin g1415 <= g7558; end
	always @ (posedge clk) begin g1417 <= g7559; end
	always @ (posedge clk) begin g1419 <= g7560; end
	always @ (posedge clk) begin g1421 <= g7561; end
	always @ (posedge clk) begin g1423 <= g7562; end
	always @ (posedge clk) begin g1425 <= g7563; end
	always @ (posedge clk) begin g1427 <= g7564; end
	always @ (posedge clk) begin g1429 <= g7565; end
	always @ (posedge clk) begin g1431 <= g7566; end
	always @ (posedge clk) begin g1433 <= g7567; end
	always @ (posedge clk) begin g1435 <= g7568; end
	always @ (posedge clk) begin g1437 <= g7569; end
	always @ (posedge clk) begin g1439 <= g7570; end
	always @ (posedge clk) begin g1443 <= g7571; end
	always @ (posedge clk) begin g1445 <= g7572; end
	always @ (posedge clk) begin g1447 <= g7573; end
	always @ (posedge clk) begin g1449 <= g7574; end
	always @ (posedge clk) begin g1451 <= g7575; end
	always @ (posedge clk) begin g1453 <= g7576; end
	always @ (posedge clk) begin g1455 <= g7577; end
	always @ (posedge clk) begin g1457 <= g7578; end
	always @ (posedge clk) begin g1459 <= g7579; end
	always @ (posedge clk) begin g1461 <= g7580; end
	always @ (posedge clk) begin g1463 <= g7581; end
	always @ (posedge clk) begin g1465 <= g7582; end
	always @ (posedge clk) begin g1467 <= g7583; end
	always @ (posedge clk) begin g1469 <= g7584; end
	always @ (posedge clk) begin g1471 <= g7585; end
	always @ (posedge clk) begin g1473 <= g7586; end
	always @ (posedge clk) begin g1477 <= g7587; end
	always @ (posedge clk) begin g1479 <= g7588; end
	always @ (posedge clk) begin g1481 <= g7589; end
	always @ (posedge clk) begin g1483 <= g7590; end
	always @ (posedge clk) begin g1485 <= g7591; end
	always @ (posedge clk) begin g1487 <= g7592; end
	always @ (posedge clk) begin g1489 <= g7593; end
	always @ (posedge clk) begin g1491 <= g7594; end
	always @ (posedge clk) begin g1493 <= g7595; end
	always @ (posedge clk) begin g1495 <= g7596; end
	always @ (posedge clk) begin g1497 <= g7597; end
	always @ (posedge clk) begin g1499 <= g7598; end
	always @ (posedge clk) begin g1501 <= g7599; end
	always @ (posedge clk) begin g1503 <= g7600; end
	always @ (posedge clk) begin g1505 <= g7601; end
	always @ (posedge clk) begin g1507 <= g7602; end
	always @ (posedge clk) begin g1510 <= g7603; end
	always @ (posedge clk) begin g1512 <= g7604; end
	always @ (posedge clk) begin g1514 <= g7605; end
	always @ (posedge clk) begin g1516 <= g7606; end
	always @ (posedge clk) begin g1518 <= g7607; end
	always @ (posedge clk) begin g1520 <= g7608; end
	always @ (posedge clk) begin g1522 <= g7609; end
	always @ (posedge clk) begin g1524 <= g7610; end
	always @ (posedge clk) begin g1526 <= g7611; end
	always @ (posedge clk) begin g1528 <= g7612; end
	always @ (posedge clk) begin g1530 <= g7613; end
	always @ (posedge clk) begin g1532 <= g7614; end
	always @ (posedge clk) begin g1534 <= g7615; end
	always @ (posedge clk) begin g1536 <= g7616; end
	always @ (posedge clk) begin g1538 <= g7617; end
	always @ (posedge clk) begin g1540 <= g7618; end
	always @ (posedge clk) begin g1547 <= g7619; end
	always @ (posedge clk) begin g1549 <= g7620; end
	always @ (posedge clk) begin g1551 <= g7621; end
	always @ (posedge clk) begin g1553 <= g7622; end
	always @ (posedge clk) begin g1555 <= g7623; end
	always @ (posedge clk) begin g1557 <= g7624; end
	always @ (posedge clk) begin g1559 <= g7625; end
	always @ (posedge clk) begin g1561 <= g7626; end
	always @ (posedge clk) begin g1563 <= g7627; end
	always @ (posedge clk) begin g1565 <= g7628; end
	always @ (posedge clk) begin g1567 <= g7629; end
	always @ (posedge clk) begin g1569 <= g7630; end
	always @ (posedge clk) begin g1571 <= g7631; end
	always @ (posedge clk) begin g1573 <= g7632; end
	always @ (posedge clk) begin g1575 <= g7633; end
	always @ (posedge clk) begin g1577 <= g7634; end
	always @ (posedge clk) begin g1580 <= g7635; end
	always @ (posedge clk) begin g1582 <= g7636; end
	always @ (posedge clk) begin g1584 <= g7637; end
	always @ (posedge clk) begin g1586 <= g7638; end
	always @ (posedge clk) begin g1588 <= g7639; end
	always @ (posedge clk) begin g1590 <= g7640; end
	always @ (posedge clk) begin g1592 <= g7641; end
	always @ (posedge clk) begin g1594 <= g7642; end
	always @ (posedge clk) begin g1596 <= g7643; end
	always @ (posedge clk) begin g1598 <= g7644; end
	always @ (posedge clk) begin g1600 <= g7645; end
	always @ (posedge clk) begin g1602 <= g7646; end
	always @ (posedge clk) begin g1604 <= g7647; end
	always @ (posedge clk) begin g1606 <= g7648; end
	always @ (posedge clk) begin g1608 <= g7649; end
	always @ (posedge clk) begin g1610 <= g7650; end
	always @ (posedge clk) begin g1614 <= g7651; end
	always @ (posedge clk) begin g1616 <= g7652; end
	always @ (posedge clk) begin g1618 <= g7653; end
	always @ (posedge clk) begin g1620 <= g7654; end
	always @ (posedge clk) begin g1622 <= g7655; end
	always @ (posedge clk) begin g1624 <= g7656; end
	always @ (posedge clk) begin g1626 <= g7657; end
	always @ (posedge clk) begin g1628 <= g7658; end
	always @ (posedge clk) begin g1630 <= g7659; end
	always @ (posedge clk) begin g1632 <= g7660; end
	always @ (posedge clk) begin g1634 <= g7661; end
	always @ (posedge clk) begin g1636 <= g7662; end
	always @ (posedge clk) begin g1638 <= g7663; end
	always @ (posedge clk) begin g1640 <= g7664; end
	always @ (posedge clk) begin g1642 <= g7665; end
	always @ (posedge clk) begin g1644 <= g7666; end
	always @ (posedge clk) begin g1647 <= g7667; end
	always @ (posedge clk) begin g1649 <= g7668; end
	always @ (posedge clk) begin g1651 <= g7669; end
	always @ (posedge clk) begin g1653 <= g7670; end
	always @ (posedge clk) begin g1655 <= g7671; end
	always @ (posedge clk) begin g1657 <= g7672; end
	always @ (posedge clk) begin g1659 <= g7673; end
	always @ (posedge clk) begin g1661 <= g7674; end
	always @ (posedge clk) begin g1663 <= g7675; end
	always @ (posedge clk) begin g1665 <= g7676; end
	always @ (posedge clk) begin g1667 <= g7677; end
	always @ (posedge clk) begin g1669 <= g7678; end
	always @ (posedge clk) begin g1671 <= g7679; end
	always @ (posedge clk) begin g1673 <= g7680; end
	always @ (posedge clk) begin g1675 <= g7681; end
	always @ (posedge clk) begin g1677 <= g7682; end
	always @ (posedge clk) begin g1681 <= g7683; end
	always @ (posedge clk) begin g1683 <= g7684; end
	always @ (posedge clk) begin g1685 <= g7685; end
	always @ (posedge clk) begin g1687 <= g7686; end
	always @ (posedge clk) begin g1689 <= g7687; end
	always @ (posedge clk) begin g1691 <= g7688; end
	always @ (posedge clk) begin g1693 <= g7689; end
	always @ (posedge clk) begin g1695 <= g7690; end
	always @ (posedge clk) begin g1697 <= g7691; end
	always @ (posedge clk) begin g1699 <= g7692; end
	always @ (posedge clk) begin g1701 <= g7693; end
	always @ (posedge clk) begin g1703 <= g7694; end
	always @ (posedge clk) begin g1705 <= g7695; end
	always @ (posedge clk) begin g1707 <= g7696; end
	always @ (posedge clk) begin g1709 <= g7697; end
	always @ (posedge clk) begin g1711 <= g7698; end
	always @ (posedge clk) begin g1714 <= g7699; end
	always @ (posedge clk) begin g1716 <= g7700; end
	always @ (posedge clk) begin g1718 <= g7701; end
	always @ (posedge clk) begin g1720 <= g7702; end
	always @ (posedge clk) begin g1722 <= g7703; end
	always @ (posedge clk) begin g1724 <= g7704; end
	always @ (posedge clk) begin g1726 <= g7705; end
	always @ (posedge clk) begin g1728 <= g7706; end
	always @ (posedge clk) begin g1730 <= g7707; end
	always @ (posedge clk) begin g1732 <= g7708; end
	always @ (posedge clk) begin g1734 <= g7709; end
	always @ (posedge clk) begin g1736 <= g7710; end
	always @ (posedge clk) begin g1738 <= g7711; end
	always @ (posedge clk) begin g1740 <= g7712; end
	always @ (posedge clk) begin g1742 <= g7713; end
	always @ (posedge clk) begin g1744 <= g7714; end
	always @ (posedge clk) begin g1748 <= g7715; end
	always @ (posedge clk) begin g1750 <= g7716; end
	always @ (posedge clk) begin g1752 <= g7717; end
	always @ (posedge clk) begin g1754 <= g7718; end
	always @ (posedge clk) begin g1756 <= g7719; end
	always @ (posedge clk) begin g1758 <= g7720; end
	always @ (posedge clk) begin g1760 <= g7721; end
	always @ (posedge clk) begin g1762 <= g7722; end
	always @ (posedge clk) begin g1764 <= g7723; end
	always @ (posedge clk) begin g1766 <= g7724; end
	always @ (posedge clk) begin g1768 <= g7725; end
	always @ (posedge clk) begin g1770 <= g7726; end
	always @ (posedge clk) begin g1772 <= g7727; end
	always @ (posedge clk) begin g1774 <= g7728; end
	always @ (posedge clk) begin g1776 <= g7729; end
	always @ (posedge clk) begin g1778 <= g7730; end
	always @ (posedge clk) begin g1784 <= g7731; end
	always @ (posedge clk) begin g1786 <= g7732; end
	always @ (posedge clk) begin g1788 <= g7733; end
	always @ (posedge clk) begin g1790 <= g7734; end
	always @ (posedge clk) begin g1792 <= g7735; end
	always @ (posedge clk) begin g1794 <= g7736; end
	always @ (posedge clk) begin g1796 <= g7737; end
	always @ (posedge clk) begin g1798 <= g7738; end
	always @ (posedge clk) begin g1800 <= g7739; end
	always @ (posedge clk) begin g1802 <= g7740; end
	always @ (posedge clk) begin g1804 <= g7741; end
	always @ (posedge clk) begin g1806 <= g7742; end
	always @ (posedge clk) begin g1808 <= g7743; end
	always @ (posedge clk) begin g1810 <= g7744; end
	always @ (posedge clk) begin g1812 <= g7745; end
	always @ (posedge clk) begin g1814 <= g7746; end
	always @ (posedge clk) begin g1817 <= g7747; end
	always @ (posedge clk) begin g1819 <= g7748; end
	always @ (posedge clk) begin g1821 <= g7749; end
	always @ (posedge clk) begin g1823 <= g7750; end
	always @ (posedge clk) begin g1825 <= g7751; end
	always @ (posedge clk) begin g1827 <= g7752; end
	always @ (posedge clk) begin g1829 <= g7753; end
	always @ (posedge clk) begin g1831 <= g7754; end
	always @ (posedge clk) begin g1833 <= g7755; end
	always @ (posedge clk) begin g1835 <= g7756; end
	always @ (posedge clk) begin g1837 <= g7757; end
	always @ (posedge clk) begin g1839 <= g7758; end
	always @ (posedge clk) begin g1841 <= g7759; end
	always @ (posedge clk) begin g1843 <= g7760; end
	always @ (posedge clk) begin g1845 <= g7761; end
	always @ (posedge clk) begin g1847 <= g7762; end
	always @ (posedge clk) begin g1851 <= g7763; end
	always @ (posedge clk) begin g1853 <= g7764; end
	always @ (posedge clk) begin g1855 <= g7765; end
	always @ (posedge clk) begin g1857 <= g7766; end
	always @ (posedge clk) begin g1859 <= g7767; end
	always @ (posedge clk) begin g1861 <= g7768; end
	always @ (posedge clk) begin g1863 <= g7769; end
	always @ (posedge clk) begin g1865 <= g7770; end
	always @ (posedge clk) begin g1867 <= g7771; end
	always @ (posedge clk) begin g1869 <= g7772; end
	always @ (posedge clk) begin g1871 <= g7773; end
	always @ (posedge clk) begin g1873 <= g7774; end
	always @ (posedge clk) begin g1875 <= g7775; end
	always @ (posedge clk) begin g1877 <= g7776; end
	always @ (posedge clk) begin g1879 <= g7777; end
	always @ (posedge clk) begin g1881 <= g7778; end
	always @ (posedge clk) begin g1884 <= g7779; end
	always @ (posedge clk) begin g1886 <= g7780; end
	always @ (posedge clk) begin g1888 <= g7781; end
	always @ (posedge clk) begin g1890 <= g7782; end
	always @ (posedge clk) begin g1892 <= g7783; end
	always @ (posedge clk) begin g1894 <= g7784; end
	always @ (posedge clk) begin g1896 <= g7785; end
	always @ (posedge clk) begin g1898 <= g7786; end
	always @ (posedge clk) begin g1900 <= g7787; end
	always @ (posedge clk) begin g1902 <= g7788; end
	always @ (posedge clk) begin g1904 <= g7789; end
	always @ (posedge clk) begin g1906 <= g7790; end
	always @ (posedge clk) begin g1908 <= g7791; end
	always @ (posedge clk) begin g1910 <= g7792; end
	always @ (posedge clk) begin g1912 <= g7793; end
	always @ (posedge clk) begin g1914 <= g7794; end
	always @ (posedge clk) begin g1915 <= g7795; end
	always @ (posedge clk) begin g1916 <= g7796; end
	always @ (posedge clk) begin g1917 <= g7797; end
	always @ (posedge clk) begin g1918 <= g7798; end
	always @ (posedge clk) begin g1919 <= g7799; end
	always @ (posedge clk) begin g1920 <= g7800; end
	always @ (posedge clk) begin g1922 <= g7801; end
	always @ (posedge clk) begin g1924 <= g7802; end
	always @ (posedge clk) begin g1925 <= g7803; end
	always @ (posedge clk) begin g1926 <= g7804; end
	always @ (posedge clk) begin g1927 <= g7805; end
	always @ (posedge clk) begin g1928 <= g7806; end
	always @ (posedge clk) begin g1929 <= g7807; end
	always @ (posedge clk) begin g1931 <= g7808; end
	always @ (posedge clk) begin g1932 <= g7809; end
	always @ (posedge clk) begin g1935 <= g7810; end
	always @ (posedge clk) begin g1939 <= g7811; end
	always @ (posedge clk) begin g1940 <= g7812; end
	always @ (posedge clk) begin g1941 <= g7813; end
	always @ (posedge clk) begin g1942 <= g7814; end
	always @ (posedge clk) begin g1944 <= g7815; end
	always @ (posedge clk) begin g1945 <= g7816; end
	always @ (posedge clk) begin g1946 <= g7817; end
	always @ (posedge clk) begin g1947 <= g7818; end
	always @ (posedge clk) begin g1948 <= g7819; end
	always @ (posedge clk) begin g1949 <= g7820; end
	always @ (posedge clk) begin g1953 <= g7821; end
	always @ (posedge clk) begin g1954 <= g7822; end
	always @ (posedge clk) begin g1955 <= g7823; end
	always @ (posedge clk) begin g1956 <= g7824; end
	always @ (posedge clk) begin g1958 <= g7825; end
	always @ (posedge clk) begin g1959 <= g7826; end
	always @ (posedge clk) begin g1960 <= g7827; end
	always @ (posedge clk) begin g1961 <= g7828; end
	always @ (posedge clk) begin g1962 <= g7829; end
	always @ (posedge clk) begin g1963 <= g7830; end
	always @ (posedge clk) begin g1967 <= g7831; end
	always @ (posedge clk) begin g1968 <= g7832; end
	always @ (posedge clk) begin g1969 <= g7833; end
	always @ (posedge clk) begin g1970 <= g7834; end
	always @ (posedge clk) begin g1972 <= g7835; end
	always @ (posedge clk) begin g1973 <= g7836; end
	always @ (posedge clk) begin g1975 <= g7837; end
	always @ (posedge clk) begin g1976 <= g7838; end
	always @ (posedge clk) begin g1977 <= g7839; end
	always @ (posedge clk) begin g1978 <= g7840; end
	always @ (posedge clk) begin g1979 <= g7841; end
	always @ (posedge clk) begin g1980 <= g7842; end
	always @ (posedge clk) begin g1982 <= g7843; end
	always @ (posedge clk) begin g1983 <= g7844; end
	always @ (posedge clk) begin g1984 <= g7845; end
	always @ (posedge clk) begin g1985 <= g7846; end
	always @ (posedge clk) begin g1986 <= g7847; end
	always @ (posedge clk) begin g1987 <= g7848; end
	always @ (posedge clk) begin g1991 <= g7849; end
	always @ (posedge clk) begin g1992 <= g7850; end
	always @ (posedge clk) begin g1993 <= g7851; end
	always @ (posedge clk) begin g1994 <= g7852; end
	always @ (posedge clk) begin g1996 <= g7853; end
	always @ (posedge clk) begin g1997 <= g7854; end
	always @ (posedge clk) begin g1998 <= g7855; end
	always @ (posedge clk) begin g1999 <= g7856; end
	always @ (posedge clk) begin g2001 <= g7857; end
	always @ (posedge clk) begin g2002 <= g7858; end
	always @ (posedge clk) begin g2003 <= g7859; end
	always @ (posedge clk) begin g2004 <= g7860; end
	always @ (posedge clk) begin g2005 <= g7861; end
	always @ (posedge clk) begin g2006 <= g7862; end
	always @ (posedge clk) begin g2011 <= g7863; end
	always @ (posedge clk) begin g2012 <= g7864; end
	always @ (posedge clk) begin g2013 <= g7865; end
	always @ (posedge clk) begin g2014 <= g7866; end
	always @ (posedge clk) begin g2022 <= g7867; end
	always @ (posedge clk) begin g2026 <= g7868; end
	always @ (posedge clk) begin g2028 <= g7869; end
	always @ (posedge clk) begin g2030 <= g7870; end
	always @ (posedge clk) begin g2032 <= g7871; end
	always @ (posedge clk) begin g2034 <= g7872; end
	always @ (posedge clk) begin g2036 <= g7873; end
	always @ (posedge clk) begin g2038 <= g7874; end
	always @ (posedge clk) begin g2041 <= g7875; end
	always @ (posedge clk) begin g2043 <= g7876; end
	always @ (posedge clk) begin g2045 <= g7877; end
	always @ (posedge clk) begin g2047 <= g7878; end
	always @ (posedge clk) begin g2048 <= g7879; end
	always @ (posedge clk) begin g2051 <= g7880; end
	always @ (posedge clk) begin g2052 <= g7881; end
	always @ (posedge clk) begin g2055 <= g7882; end
	always @ (posedge clk) begin g2062 <= g7883; end
	always @ (posedge clk) begin g2065 <= g7884; end
	always @ (posedge clk) begin g2068 <= g7885; end
	always @ (posedge clk) begin g2071 <= g7886; end
	always @ (posedge clk) begin g2074 <= g7887; end
	always @ (posedge clk) begin g2077 <= g7888; end
	always @ (posedge clk) begin g2080 <= g7889; end
	always @ (posedge clk) begin g2085 <= g7890; end
	always @ (posedge clk) begin g2088 <= g7891; end
	always @ (posedge clk) begin g2091 <= g7892; end
	always @ (posedge clk) begin g2098 <= g7893; end
	always @ (posedge clk) begin g2099 <= g7894; end
	always @ (posedge clk) begin g2100 <= g7895; end
	always @ (posedge clk) begin g2101 <= g7896; end
	always @ (posedge clk) begin g2104 <= g7897; end
	always @ (posedge clk) begin g2108 <= g7898; end
	always @ (posedge clk) begin g2110 <= g7899; end
	always @ (posedge clk) begin g2112 <= g7900; end
	always @ (posedge clk) begin g2114 <= g7901; end
	always @ (posedge clk) begin g2116 <= g7902; end
	always @ (posedge clk) begin g2118 <= g7903; end
	always @ (posedge clk) begin g2120 <= g7904; end
	always @ (posedge clk) begin g2123 <= g7905; end
	always @ (posedge clk) begin g2125 <= g7906; end
	always @ (posedge clk) begin g2127 <= g7907; end
	always @ (posedge clk) begin g2129 <= g7908; end
	always @ (posedge clk) begin g2130 <= g7909; end
	always @ (posedge clk) begin g2133 <= g7910; end
	always @ (posedge clk) begin g2134 <= g7911; end
	always @ (posedge clk) begin g2137 <= g7912; end
	always @ (posedge clk) begin g2144 <= g7913; end
	always @ (posedge clk) begin g2147 <= g7914; end
	always @ (posedge clk) begin g2150 <= g7915; end
	always @ (posedge clk) begin g2153 <= g7916; end
	always @ (posedge clk) begin g2156 <= g7917; end
	always @ (posedge clk) begin g2159 <= g7918; end
	always @ (posedge clk) begin g2162 <= g7919; end
	always @ (posedge clk) begin g2167 <= g7920; end
	always @ (posedge clk) begin g2170 <= g7921; end
	always @ (posedge clk) begin g2173 <= g7922; end
	always @ (posedge clk) begin g2177 <= g7923; end
	always @ (posedge clk) begin g2178 <= g7924; end
	always @ (posedge clk) begin g2180 <= g7925; end
	always @ (posedge clk) begin g2181 <= g7926; end
	always @ (posedge clk) begin g2184 <= g7927; end
	always @ (posedge clk) begin g2188 <= g7928; end
	always @ (posedge clk) begin g2190 <= g7929; end
	always @ (posedge clk) begin g2192 <= g7930; end
	always @ (posedge clk) begin g2194 <= g7931; end
	always @ (posedge clk) begin g2196 <= g7932; end
	always @ (posedge clk) begin g2198 <= g7933; end
	always @ (posedge clk) begin g2200 <= g7934; end
	always @ (posedge clk) begin g2203 <= g7935; end
	always @ (posedge clk) begin g2205 <= g7936; end
	always @ (posedge clk) begin g2207 <= g7937; end
	always @ (posedge clk) begin g2210 <= g7938; end
	always @ (posedge clk) begin g2211 <= g7939; end
	always @ (posedge clk) begin g2212 <= g7940; end
	always @ (posedge clk) begin g2213 <= g7941; end
	always @ (posedge clk) begin g2217 <= g7942; end
	always @ (posedge clk) begin g2224 <= g7943; end
	always @ (posedge clk) begin g2227 <= g7944; end
	always @ (posedge clk) begin g2230 <= g7945; end
	always @ (posedge clk) begin g2233 <= g7946; end
	always @ (posedge clk) begin g2236 <= g7947; end
	always @ (posedge clk) begin g2239 <= g7948; end
	always @ (posedge clk) begin g2242 <= g7949; end
	always @ (posedge clk) begin g2247 <= g7950; end
	always @ (posedge clk) begin g2250 <= g7951; end
	always @ (posedge clk) begin g2253 <= g7952; end
	always @ (posedge clk) begin g2256 <= g7953; end
	always @ (posedge clk) begin g2257 <= g7954; end
	always @ (posedge clk) begin g2262 <= g7955; end
	always @ (posedge clk) begin g2263 <= g7956; end
	always @ (posedge clk) begin g2267 <= g7957; end
	always @ (posedge clk) begin g2271 <= g7958; end
	always @ (posedge clk) begin g2273 <= g7959; end
	always @ (posedge clk) begin g2275 <= g7960; end
	always @ (posedge clk) begin g2277 <= g7961; end
	always @ (posedge clk) begin g2279 <= g7962; end
	always @ (posedge clk) begin g2281 <= g7963; end
	always @ (posedge clk) begin g2283 <= g7964; end
	always @ (posedge clk) begin g2286 <= g7965; end
	always @ (posedge clk) begin g2288 <= g7966; end
	always @ (posedge clk) begin g2290 <= g7967; end
	always @ (posedge clk) begin g2295 <= g7968; end
	always @ (posedge clk) begin g2296 <= g7969; end
	always @ (posedge clk) begin g2298 <= g7970; end
	always @ (posedge clk) begin g2299 <= g7971; end
	always @ (posedge clk) begin g2304 <= g7972; end
	always @ (posedge clk) begin g2311 <= g7973; end
	always @ (posedge clk) begin g2314 <= g7974; end
	always @ (posedge clk) begin g2317 <= g7975; end
	always @ (posedge clk) begin g2320 <= g7976; end
	always @ (posedge clk) begin g2323 <= g7977; end
	always @ (posedge clk) begin g2326 <= g7978; end
	always @ (posedge clk) begin g2329 <= g7979; end
	always @ (posedge clk) begin g2334 <= g7980; end
	always @ (posedge clk) begin g2337 <= g7981; end
	always @ (posedge clk) begin g2340 <= g7982; end
	always @ (posedge clk) begin g2343 <= g7983; end
	always @ (posedge clk) begin g2344 <= g7984; end
	always @ (posedge clk) begin g2347 <= g7985; end
	always @ (posedge clk) begin g2348 <= g7986; end
	always @ (posedge clk) begin g2350 <= g7987; end
	always @ (posedge clk) begin g2354 <= g7988; end
	always @ (posedge clk) begin g2356 <= g7989; end
	always @ (posedge clk) begin g2358 <= g7990; end
	always @ (posedge clk) begin g2360 <= g7991; end
	always @ (posedge clk) begin g2362 <= g7992; end
	always @ (posedge clk) begin g2364 <= g7993; end
	always @ (posedge clk) begin g2366 <= g7994; end
	always @ (posedge clk) begin g2369 <= g7995; end
	always @ (posedge clk) begin g2371 <= g7996; end
	always @ (posedge clk) begin g2373 <= g7997; end
	always @ (posedge clk) begin g2376 <= g7998; end
	always @ (posedge clk) begin g2377 <= g7999; end
	always @ (posedge clk) begin g2378 <= g8000; end
	always @ (posedge clk) begin g2379 <= g8001; end
	always @ (posedge clk) begin g2383 <= g8002; end
	always @ (posedge clk) begin g2390 <= g8003; end
	always @ (posedge clk) begin g2393 <= g8004; end
	always @ (posedge clk) begin g2396 <= g8005; end
	always @ (posedge clk) begin g2399 <= g8006; end
	always @ (posedge clk) begin g2402 <= g8007; end
	always @ (posedge clk) begin g2405 <= g8008; end
	always @ (posedge clk) begin g2408 <= g8009; end
	always @ (posedge clk) begin g2413 <= g8010; end
	always @ (posedge clk) begin g2416 <= g8011; end
	always @ (posedge clk) begin g2419 <= g8012; end
	always @ (posedge clk) begin g2423 <= g8013; end
	always @ (posedge clk) begin g2424 <= g8014; end
	always @ (posedge clk) begin g2426 <= g8015; end
	always @ (posedge clk) begin g2427 <= g8016; end
	always @ (posedge clk) begin g2434 <= g8017; end
	always @ (posedge clk) begin g2450 <= g8018; end
	always @ (posedge clk) begin g2456 <= g8019; end
	always @ (posedge clk) begin g2462 <= g8020; end
	always @ (posedge clk) begin g2468 <= g8021; end
	always @ (posedge clk) begin g2474 <= g8022; end
	always @ (posedge clk) begin g2480 <= g8023; end
	always @ (posedge clk) begin g2486 <= g8024; end
	always @ (posedge clk) begin g2497 <= g8025; end
	always @ (posedge clk) begin g2503 <= g8026; end
	always @ (posedge clk) begin g2509 <= g8027; end
	always @ (posedge clk) begin g2515 <= g8028; end
	always @ (posedge clk) begin g2516 <= g8029; end
	always @ (posedge clk) begin g2518 <= g8030; end
	always @ (posedge clk) begin g2519 <= g8031; end
	always @ (posedge clk) begin g2523 <= g8032; end
	always @ (posedge clk) begin g2527 <= g8033; end
	always @ (posedge clk) begin g2529 <= g8034; end
	always @ (posedge clk) begin g2531 <= g8035; end
	always @ (posedge clk) begin g2533 <= g8036; end
	always @ (posedge clk) begin g2535 <= g8037; end
	always @ (posedge clk) begin g2537 <= g8038; end
	always @ (posedge clk) begin g2539 <= g8039; end
	always @ (posedge clk) begin g2542 <= g8040; end
	always @ (posedge clk) begin g2544 <= g8041; end
	always @ (posedge clk) begin g2546 <= g8042; end
	always @ (posedge clk) begin g2551 <= g8043; end
	always @ (posedge clk) begin g2552 <= g8044; end
	always @ (posedge clk) begin g2555 <= g8045; end
	always @ (posedge clk) begin g2556 <= g8046; end
	always @ (posedge clk) begin g2559 <= g8047; end
	always @ (posedge clk) begin g2566 <= g8048; end
	always @ (posedge clk) begin g2569 <= g8049; end
	always @ (posedge clk) begin g2572 <= g8050; end
	always @ (posedge clk) begin g2575 <= g8051; end
	always @ (posedge clk) begin g2578 <= g8052; end
	always @ (posedge clk) begin g2581 <= g8053; end
	always @ (posedge clk) begin g2584 <= g8054; end
	always @ (posedge clk) begin g2589 <= g8055; end
	always @ (posedge clk) begin g2592 <= g8056; end
	always @ (posedge clk) begin g2595 <= g8057; end
	always @ (posedge clk) begin g2598 <= g8058; end
	always @ (posedge clk) begin g2599 <= g8059; end
	always @ (posedge clk) begin g2601 <= g8060; end
	always @ (posedge clk) begin g2602 <= g8061; end
	always @ (posedge clk) begin g2607 <= g8062; end
	always @ (posedge clk) begin g2614 <= g8063; end
	always @ (posedge clk) begin g2617 <= g8064; end
	always @ (posedge clk) begin g2620 <= g8065; end
	always @ (posedge clk) begin g2623 <= g8066; end
	always @ (posedge clk) begin g2626 <= g8067; end
	always @ (posedge clk) begin g2629 <= g8068; end
	always @ (posedge clk) begin g2632 <= g8069; end
	always @ (posedge clk) begin g2637 <= g8070; end
	always @ (posedge clk) begin g2640 <= g8071; end
	always @ (posedge clk) begin g2643 <= g8072; end
	always @ (posedge clk) begin g2647 <= g8073; end
	always @ (posedge clk) begin g2648 <= g8074; end
	always @ (posedge clk) begin g2649 <= g8075; end
	always @ (posedge clk) begin g2650 <= g8076; end
	always @ (posedge clk) begin g2653 <= g8077; end
	always @ (posedge clk) begin g2657 <= g8078; end
	always @ (posedge clk) begin g2659 <= g8079; end
	always @ (posedge clk) begin g2661 <= g8080; end
	always @ (posedge clk) begin g2663 <= g8081; end
	always @ (posedge clk) begin g2665 <= g8082; end
	always @ (posedge clk) begin g2667 <= g8083; end
	always @ (posedge clk) begin g2669 <= g8084; end
	always @ (posedge clk) begin g2672 <= g8085; end
	always @ (posedge clk) begin g2674 <= g8086; end
	always @ (posedge clk) begin g2676 <= g8087; end
	always @ (posedge clk) begin g2678 <= g8088; end
	always @ (posedge clk) begin g2679 <= g8089; end
	always @ (posedge clk) begin g2683 <= g8090; end
	always @ (posedge clk) begin g2684 <= g8091; end
	always @ (posedge clk) begin g2690 <= g8092; end
	always @ (posedge clk) begin g2703 <= g8093; end
	always @ (posedge clk) begin g2708 <= g8094; end
	always @ (posedge clk) begin g2713 <= g8095; end
	always @ (posedge clk) begin g2718 <= g8096; end
	always @ (posedge clk) begin g2723 <= g8097; end
	always @ (posedge clk) begin g2728 <= g8098; end
	always @ (posedge clk) begin g2733 <= g8099; end
	always @ (posedge clk) begin g2742 <= g8100; end
	always @ (posedge clk) begin g2747 <= g8101; end
	always @ (posedge clk) begin g2752 <= g8102; end
	always @ (posedge clk) begin g2758 <= g8103; end
	always @ (posedge clk) begin g2759 <= g8104; end
	always @ (posedge clk) begin g2760 <= g8105; end
	always @ (posedge clk) begin g2761 <= g8106; end
	always @ (posedge clk) begin g2764 <= g8107; end
	always @ (posedge clk) begin g2768 <= g8108; end
	always @ (posedge clk) begin g2770 <= g8109; end
	always @ (posedge clk) begin g2772 <= g8110; end
	always @ (posedge clk) begin g2774 <= g8111; end
	always @ (posedge clk) begin g2776 <= g8112; end
	always @ (posedge clk) begin g2778 <= g8113; end
	always @ (posedge clk) begin g2780 <= g8114; end
	always @ (posedge clk) begin g2783 <= g8115; end
	always @ (posedge clk) begin g2785 <= g8116; end
	always @ (posedge clk) begin g2787 <= g8117; end
	always @ (posedge clk) begin g2789 <= g8118; end
	always @ (posedge clk) begin g2790 <= g8119; end
	always @ (posedge clk) begin g2793 <= g8120; end
	always @ (posedge clk) begin g2794 <= g8121; end
	always @ (posedge clk) begin g2797 <= g8122; end
	always @ (posedge clk) begin g2804 <= g8123; end
	always @ (posedge clk) begin g2807 <= g8124; end
	always @ (posedge clk) begin g2810 <= g8125; end
	always @ (posedge clk) begin g2813 <= g8126; end
	always @ (posedge clk) begin g2816 <= g8127; end
	always @ (posedge clk) begin g2819 <= g8128; end
	always @ (posedge clk) begin g2822 <= g8129; end
	always @ (posedge clk) begin g2827 <= g8130; end
	always @ (posedge clk) begin g2830 <= g8131; end
	always @ (posedge clk) begin g2833 <= g8132; end
	always @ (posedge clk) begin g2838 <= g8133; end
	always @ (posedge clk) begin g2845 <= g8134; end
	always @ (posedge clk) begin g2848 <= g8135; end
	always @ (posedge clk) begin g2851 <= g8136; end
	always @ (posedge clk) begin g2854 <= g8137; end
	always @ (posedge clk) begin g2857 <= g8138; end
	always @ (posedge clk) begin g2860 <= g8139; end
	always @ (posedge clk) begin g2863 <= g8140; end
	always @ (posedge clk) begin g2868 <= g8141; end
	always @ (posedge clk) begin g2871 <= g8142; end
	always @ (posedge clk) begin g2874 <= g8143; end
	always @ (posedge clk) begin g2881 <= g8144; end
	always @ (posedge clk) begin g2885 <= g8145; end
	always @ (posedge clk) begin g2887 <= g8146; end
	always @ (posedge clk) begin g2889 <= g8147; end
	always @ (posedge clk) begin g2891 <= g8148; end
	always @ (posedge clk) begin g2893 <= g8149; end
	always @ (posedge clk) begin g2895 <= g8150; end
	always @ (posedge clk) begin g2897 <= g8151; end
	always @ (posedge clk) begin g2900 <= g8152; end
	always @ (posedge clk) begin g2902 <= g8153; end
	always @ (posedge clk) begin g2904 <= g8154; end
	always @ (posedge clk) begin g2916 <= g8155; end
	always @ (posedge clk) begin g2932 <= g8156; end
	always @ (posedge clk) begin g2938 <= g8157; end
	always @ (posedge clk) begin g2944 <= g8158; end
	always @ (posedge clk) begin g2950 <= g8159; end
	always @ (posedge clk) begin g2956 <= g8160; end
	always @ (posedge clk) begin g2962 <= g8161; end
	always @ (posedge clk) begin g2968 <= g8162; end
	always @ (posedge clk) begin g2979 <= g8163; end
	always @ (posedge clk) begin g2985 <= g8164; end
	always @ (posedge clk) begin g2991 <= g8165; end
	always @ (posedge clk) begin g2999 <= g8166; end
	always @ (posedge clk) begin g3003 <= g8167; end
	always @ (posedge clk) begin g3005 <= g8168; end
	always @ (posedge clk) begin g3007 <= g8169; end
	always @ (posedge clk) begin g3009 <= g8170; end
	always @ (posedge clk) begin g3011 <= g8171; end
	always @ (posedge clk) begin g3013 <= g8172; end
	always @ (posedge clk) begin g3015 <= g8173; end
	always @ (posedge clk) begin g3018 <= g8174; end
	always @ (posedge clk) begin g3020 <= g8175; end
	always @ (posedge clk) begin g3022 <= g8176; end
	always @ (posedge clk) begin g3031 <= g8177; end
	always @ (posedge clk) begin g3038 <= g8178; end
	always @ (posedge clk) begin g3041 <= g8179; end
	always @ (posedge clk) begin g3044 <= g8180; end
	always @ (posedge clk) begin g3047 <= g8181; end
	always @ (posedge clk) begin g3050 <= g8182; end
	always @ (posedge clk) begin g3053 <= g8183; end
	always @ (posedge clk) begin g3056 <= g8184; end
	always @ (posedge clk) begin g3061 <= g8185; end
	always @ (posedge clk) begin g3064 <= g8186; end
	always @ (posedge clk) begin g3067 <= g8187; end
	always @ (posedge clk) begin g3074 <= g8188; end
	always @ (posedge clk) begin g3078 <= g8189; end
	always @ (posedge clk) begin g3080 <= g8190; end
	always @ (posedge clk) begin g3082 <= g8191; end
	always @ (posedge clk) begin g3084 <= g8192; end
	always @ (posedge clk) begin g3086 <= g8193; end
	always @ (posedge clk) begin g3088 <= g8194; end
	always @ (posedge clk) begin g3090 <= g8195; end
	always @ (posedge clk) begin g3093 <= g8196; end
	always @ (posedge clk) begin g3095 <= g8197; end
	always @ (posedge clk) begin g3097 <= g8198; end
	always @ (posedge clk) begin g3106 <= g8199; end
	always @ (posedge clk) begin g3113 <= g8200; end
	always @ (posedge clk) begin g3116 <= g8201; end
	always @ (posedge clk) begin g3119 <= g8202; end
	always @ (posedge clk) begin g3122 <= g8203; end
	always @ (posedge clk) begin g3125 <= g8204; end
	always @ (posedge clk) begin g3128 <= g8205; end
	always @ (posedge clk) begin g3131 <= g8206; end
	always @ (posedge clk) begin g3136 <= g8207; end
	always @ (posedge clk) begin g3139 <= g8208; end
	always @ (posedge clk) begin g3142 <= g8209; end
	always @ (posedge clk) begin g3149 <= g8210; end
	always @ (posedge clk) begin g3153 <= g8211; end
	always @ (posedge clk) begin g3155 <= g8212; end
	always @ (posedge clk) begin g3157 <= g8213; end
	always @ (posedge clk) begin g3159 <= g8214; end
	always @ (posedge clk) begin g3161 <= g8215; end
	always @ (posedge clk) begin g3163 <= g8216; end
	always @ (posedge clk) begin g3165 <= g8217; end
	always @ (posedge clk) begin g3168 <= g8218; end
	always @ (posedge clk) begin g3170 <= g8219; end
	always @ (posedge clk) begin g3172 <= g8220; end
	always @ (posedge clk) begin g3177 <= g8221; end
	always @ (posedge clk) begin g3184 <= g8222; end
	always @ (posedge clk) begin g3187 <= g8223; end
	always @ (posedge clk) begin g3190 <= g8224; end
	always @ (posedge clk) begin g3193 <= g8225; end
	always @ (posedge clk) begin g3196 <= g8226; end
	always @ (posedge clk) begin g3199 <= g8227; end
	always @ (posedge clk) begin g3202 <= g8228; end
	always @ (posedge clk) begin g3207 <= g8229; end
	always @ (posedge clk) begin g3210 <= g8230; end
	always @ (posedge clk) begin g3213 <= g8231; end
	always @ (posedge clk) begin g3222 <= g8232; end
	always @ (posedge clk) begin g3235 <= g8233; end
	always @ (posedge clk) begin g3240 <= g8234; end
	always @ (posedge clk) begin g3245 <= g8235; end
	always @ (posedge clk) begin g3250 <= g8236; end
	always @ (posedge clk) begin g3255 <= g8237; end
	always @ (posedge clk) begin g3260 <= g8238; end
	always @ (posedge clk) begin g3265 <= g8239; end
	always @ (posedge clk) begin g3274 <= g8240; end
	always @ (posedge clk) begin g3279 <= g8241; end
	always @ (posedge clk) begin g3284 <= g8242; end
	always @ (posedge clk) begin g3291 <= g8243; end
	always @ (posedge clk) begin g3295 <= g8244; end
	always @ (posedge clk) begin g3297 <= g8245; end
	always @ (posedge clk) begin g3299 <= g8246; end
	always @ (posedge clk) begin g3301 <= g8247; end
	always @ (posedge clk) begin g3303 <= g8248; end
	always @ (posedge clk) begin g3305 <= g8249; end
	always @ (posedge clk) begin g3307 <= g8250; end
	always @ (posedge clk) begin g3310 <= g8251; end
	always @ (posedge clk) begin g3312 <= g8252; end
	always @ (posedge clk) begin g3314 <= g8253; end
	always @ (posedge clk) begin g3323 <= g8254; end
	always @ (posedge clk) begin g3330 <= g8255; end
	always @ (posedge clk) begin g3333 <= g8256; end
	always @ (posedge clk) begin g3336 <= g8257; end
	always @ (posedge clk) begin g3339 <= g8258; end
	always @ (posedge clk) begin g3342 <= g8259; end
	always @ (posedge clk) begin g3345 <= g8260; end
	always @ (posedge clk) begin g3348 <= g8261; end
	always @ (posedge clk) begin g3353 <= g8262; end
	always @ (posedge clk) begin g3356 <= g8263; end
	always @ (posedge clk) begin g3359 <= g8264; end
	always @ (posedge clk) begin g3366 <= g8265; end
	always @ (posedge clk) begin g3370 <= g8266; end
	always @ (posedge clk) begin g3372 <= g8267; end
	always @ (posedge clk) begin g3374 <= g8268; end
	always @ (posedge clk) begin g3376 <= g8269; end
	always @ (posedge clk) begin g3378 <= g8270; end
	always @ (posedge clk) begin g3380 <= g8271; end
	always @ (posedge clk) begin g3382 <= g8272; end
	always @ (posedge clk) begin g3385 <= g8273; end
	always @ (posedge clk) begin g3387 <= g8274; end
	always @ (posedge clk) begin g3389 <= g8275; end
	always @ (posedge clk) begin g3427 <= g8276; end
	always @ (posedge clk) begin g3687 <= g8277; end
	always @ (posedge clk) begin g4000 <= g8278; end
	always @ (posedge clk) begin g4010 <= g8279; end
	always @ (posedge clk) begin g4027 <= g8280; end
	always @ (posedge clk) begin g4036 <= g8281; end
	always @ (posedge clk) begin g4046 <= g8282; end
	always @ (posedge clk) begin g4053 <= g8283; end
	always @ (posedge clk) begin g4060 <= g8284; end
	always @ (posedge clk) begin g4068 <= g8285; end
	always @ (posedge clk) begin g4075 <= g8286; end
	always @ (posedge clk) begin g4083 <= g8287; end
	always @ (posedge clk) begin g4091 <= g8288; end
	always @ (posedge clk) begin g4098 <= g8289; end
	always @ (posedge clk) begin g4104 <= g8290; end
	always @ (posedge clk) begin g4110 <= g8291; end
	always @ (posedge clk) begin g4127 <= g8292; end
	always @ (posedge clk) begin g4177 <= g8293; end
	always @ (posedge clk) begin g4221 <= g8294; end
	always @ (posedge clk) begin g4252 <= g8295; end
	always @ (posedge clk) begin g4267 <= g8296; end
	always @ (posedge clk) begin g4315 <= g8297; end
	always @ (posedge clk) begin g4342 <= g8298; end
	always @ (posedge clk) begin g4377 <= g8299; end
	always @ (posedge clk) begin g4390 <= g8300; end
	always @ (posedge clk) begin g4426 <= g8301; end
	always @ (posedge clk) begin g4451 <= g8302; end
	always @ (posedge clk) begin g4482 <= g8303; end
	always @ (posedge clk) begin g4501 <= g8304; end
	always @ (posedge clk) begin g4545 <= g8305; end
	always @ (posedge clk) begin g4572 <= g8306; end
	always @ (posedge clk) begin g4596 <= g8307; end
	always @ (posedge clk) begin g4610 <= g8308; end
	always @ (posedge clk) begin g4649 <= g8309; end
	always @ (posedge clk) begin g4672 <= g8310; end
	always @ (posedge clk) begin g4696 <= g8311; end
	always @ (posedge clk) begin g4709 <= g8312; end
	always @ (posedge clk) begin g4749 <= g8313; end
	always @ (posedge clk) begin g4759 <= g8314; end
	always @ (posedge clk) begin g4784 <= g8315; end
	always @ (posedge clk) begin g4798 <= g8316; end
	always @ (posedge clk) begin g4835 <= g8317; end
	always @ (posedge clk) begin g4850 <= g8318; end
	always @ (posedge clk) begin g4877 <= g8319; end
	always @ (posedge clk) begin g4892 <= g8320; end
	always @ (posedge clk) begin g4931 <= g8321; end
	always @ (posedge clk) begin g4959 <= g8322; end
	always @ (posedge clk) begin g4987 <= g8323; end
	always @ (posedge clk) begin g4999 <= g8324; end
	always @ (posedge clk) begin g5033 <= g8325; end
	always @ (posedge clk) begin g5057 <= g8326; end
	always @ (posedge clk) begin g5083 <= g8327; end
	always @ (posedge clk) begin g5132 <= g8328; end
	always @ (posedge clk) begin g5165 <= g8329; end
	always @ (posedge clk) begin g5210 <= g8330; end
	always @ (posedge clk) begin g5241 <= g8331; end
	always @ (posedge clk) begin g5294 <= g8332; end
	always @ (posedge clk) begin g5323 <= g8333; end
	always @ (posedge clk) begin g5373 <= g8334; end
	always @ (posedge clk) begin g5393 <= g8335; end
	always @ (posedge clk) begin g5434 <= g8336; end
	always @ (posedge clk) begin g5463 <= g8337; end
	always @ (posedge clk) begin g5510 <= g8338; end
	always @ (posedge clk) begin g5533 <= g8339; end

	assign data_valid = (((g1)));
	assign g7197 = (((!g65) & (g64) & (!data[0])) + ((!g65) & (g64) & (data[0])) + ((g65) & (!g64) & (data[0])) + ((g65) & (g64) & (data[0])));
	assign g7198 = (((!g65) & (g88) & (!data[1])) + ((!g65) & (g88) & (data[1])) + ((g65) & (!g88) & (data[1])) + ((g65) & (g88) & (data[1])));
	assign g7199 = (((!g65) & (g111) & (!data[2])) + ((!g65) & (g111) & (data[2])) + ((g65) & (!g111) & (data[2])) + ((g65) & (g111) & (data[2])));
	assign g7200 = (((!g65) & (g134) & (!data[3])) + ((!g65) & (g134) & (data[3])) + ((g65) & (!g134) & (data[3])) + ((g65) & (g134) & (data[3])));
	assign g7201 = (((!g65) & (g157) & (!data[4])) + ((!g65) & (g157) & (data[4])) + ((g65) & (!g157) & (data[4])) + ((g65) & (g157) & (data[4])));
	assign g7202 = (((!g65) & (g180) & (!data[5])) + ((!g65) & (g180) & (data[5])) + ((g65) & (!g180) & (data[5])) + ((g65) & (g180) & (data[5])));
	assign g7203 = (((!g65) & (g203) & (!data[6])) + ((!g65) & (g203) & (data[6])) + ((g65) & (!g203) & (data[6])) + ((g65) & (g203) & (data[6])));
	assign g7204 = (((!g65) & (g226) & (!data[7])) + ((!g65) & (g226) & (data[7])) + ((g65) & (!g226) & (data[7])) + ((g65) & (g226) & (data[7])));
	assign g7205 = (((!g65) & (g249) & (!data[8])) + ((!g65) & (g249) & (data[8])) + ((g65) & (!g249) & (data[8])) + ((g65) & (g249) & (data[8])));
	assign g7206 = (((!g65) & (g272) & (!data[9])) + ((!g65) & (g272) & (data[9])) + ((g65) & (!g272) & (data[9])) + ((g65) & (g272) & (data[9])));
	assign g7207 = (((!g65) & (g295) & (!data[10])) + ((!g65) & (g295) & (data[10])) + ((g65) & (!g295) & (data[10])) + ((g65) & (g295) & (data[10])));
	assign g7208 = (((!g65) & (g318) & (!data[11])) + ((!g65) & (g318) & (data[11])) + ((g65) & (!g318) & (data[11])) + ((g65) & (g318) & (data[11])));
	assign g7209 = (((!g65) & (g341) & (!data[12])) + ((!g65) & (g341) & (data[12])) + ((g65) & (!g341) & (data[12])) + ((g65) & (g341) & (data[12])));
	assign g7210 = (((!g65) & (g364) & (!data[13])) + ((!g65) & (g364) & (data[13])) + ((g65) & (!g364) & (data[13])) + ((g65) & (g364) & (data[13])));
	assign g7211 = (((!g65) & (g387) & (!data[14])) + ((!g65) & (g387) & (data[14])) + ((g65) & (!g387) & (data[14])) + ((g65) & (g387) & (data[14])));
	assign g7212 = (((!g65) & (g410) & (!data[15])) + ((!g65) & (g410) & (data[15])) + ((g65) & (!g410) & (data[15])) + ((g65) & (g410) & (data[15])));
	assign g7213 = (((!g65) & (g433) & (!data[16])) + ((!g65) & (g433) & (data[16])) + ((g65) & (!g433) & (data[16])) + ((g65) & (g433) & (data[16])));
	assign g7214 = (((!g65) & (g456) & (!data[17])) + ((!g65) & (g456) & (data[17])) + ((g65) & (!g456) & (data[17])) + ((g65) & (g456) & (data[17])));
	assign g7215 = (((!g65) & (g479) & (!data[18])) + ((!g65) & (g479) & (data[18])) + ((g65) & (!g479) & (data[18])) + ((g65) & (g479) & (data[18])));
	assign g7216 = (((!g65) & (g502) & (!data[19])) + ((!g65) & (g502) & (data[19])) + ((g65) & (!g502) & (data[19])) + ((g65) & (g502) & (data[19])));
	assign g7217 = (((!g65) & (g525) & (!data[20])) + ((!g65) & (g525) & (data[20])) + ((g65) & (!g525) & (data[20])) + ((g65) & (g525) & (data[20])));
	assign g7218 = (((!g65) & (g548) & (!data[21])) + ((!g65) & (g548) & (data[21])) + ((g65) & (!g548) & (data[21])) + ((g65) & (g548) & (data[21])));
	assign g7219 = (((!g65) & (g571) & (!data[22])) + ((!g65) & (g571) & (data[22])) + ((g65) & (!g571) & (data[22])) + ((g65) & (g571) & (data[22])));
	assign g7220 = (((!g65) & (g594) & (!data[23])) + ((!g65) & (g594) & (data[23])) + ((g65) & (!g594) & (data[23])) + ((g65) & (g594) & (data[23])));
	assign g7221 = (((!g65) & (g617) & (!data[24])) + ((!g65) & (g617) & (data[24])) + ((g65) & (!g617) & (data[24])) + ((g65) & (g617) & (data[24])));
	assign g7222 = (((!g65) & (g640) & (!data[25])) + ((!g65) & (g640) & (data[25])) + ((g65) & (!g640) & (data[25])) + ((g65) & (g640) & (data[25])));
	assign g7223 = (((!g65) & (g663) & (!data[26])) + ((!g65) & (g663) & (data[26])) + ((g65) & (!g663) & (data[26])) + ((g65) & (g663) & (data[26])));
	assign g7224 = (((!g65) & (g686) & (!data[27])) + ((!g65) & (g686) & (data[27])) + ((g65) & (!g686) & (data[27])) + ((g65) & (g686) & (data[27])));
	assign g7225 = (((!g65) & (g709) & (!data[28])) + ((!g65) & (g709) & (data[28])) + ((g65) & (!g709) & (data[28])) + ((g65) & (g709) & (data[28])));
	assign g7226 = (((!g65) & (g732) & (!data[29])) + ((!g65) & (g732) & (data[29])) + ((g65) & (!g732) & (data[29])) + ((g65) & (g732) & (data[29])));
	assign g7227 = (((!g65) & (g755) & (!data[30])) + ((!g65) & (g755) & (data[30])) + ((g65) & (!g755) & (data[30])) + ((g65) & (g755) & (data[30])));
	assign g7228 = (((!g65) & (g778) & (!data[31])) + ((!g65) & (g778) & (data[31])) + ((g65) & (!g778) & (data[31])) + ((g65) & (g778) & (data[31])));
	assign g37 = (((!g34) & (g35) & (!g1) & (g36) & (!reset)) + ((!g34) & (g35) & (g1) & (g36) & (!reset)) + ((g34) & (!g35) & (!g1) & (g36) & (!reset)) + ((g34) & (!g35) & (g1) & (g36) & (!reset)) + ((g34) & (g35) & (g1) & (g36) & (!reset)));
	assign g7229 = (((!g797) & (g796) & (!g42)) + ((!g797) & (g796) & (g42)) + ((g797) & (!g796) & (g42)) + ((g797) & (g796) & (g42)));
	assign g7230 = (((!g797) & (g799) & (!g43)) + ((!g797) & (g799) & (g43)) + ((g797) & (!g799) & (g43)) + ((g797) & (g799) & (g43)));
	assign g44 = (((!g38) & (!g39) & (!g40) & (g41) & (g42) & (g43)) + ((!g38) & (!g39) & (g40) & (!g41) & (!g42) & (g43)) + ((!g38) & (!g39) & (g40) & (g41) & (!g42) & (g43)) + ((!g38) & (!g39) & (g40) & (g41) & (g42) & (g43)) + ((!g38) & (g39) & (!g40) & (!g41) & (g42) & (!g43)) + ((!g38) & (g39) & (!g40) & (g41) & (g42) & (!g43)) + ((!g38) & (g39) & (!g40) & (g41) & (g42) & (g43)) + ((!g38) & (g39) & (g40) & (!g41) & (!g42) & (g43)) + ((!g38) & (g39) & (g40) & (!g41) & (g42) & (!g43)) + ((!g38) & (g39) & (g40) & (g41) & (!g42) & (g43)) + ((!g38) & (g39) & (g40) & (g41) & (g42) & (!g43)) + ((!g38) & (g39) & (g40) & (g41) & (g42) & (g43)) + ((g38) & (!g39) & (!g40) & (!g41) & (!g42) & (!g43)) + ((g38) & (!g39) & (!g40) & (g41) & (!g42) & (!g43)) + ((g38) & (!g39) & (!g40) & (g41) & (g42) & (g43)) + ((g38) & (!g39) & (g40) & (!g41) & (!g42) & (!g43)) + ((g38) & (!g39) & (g40) & (!g41) & (!g42) & (g43)) + ((g38) & (!g39) & (g40) & (g41) & (!g42) & (!g43)) + ((g38) & (!g39) & (g40) & (g41) & (!g42) & (g43)) + ((g38) & (!g39) & (g40) & (g41) & (g42) & (g43)) + ((g38) & (g39) & (!g40) & (!g41) & (!g42) & (!g43)) + ((g38) & (g39) & (!g40) & (!g41) & (g42) & (!g43)) + ((g38) & (g39) & (!g40) & (g41) & (!g42) & (!g43)) + ((g38) & (g39) & (!g40) & (g41) & (g42) & (!g43)) + ((g38) & (g39) & (!g40) & (g41) & (g42) & (g43)) + ((g38) & (g39) & (g40) & (!g41) & (!g42) & (!g43)) + ((g38) & (g39) & (g40) & (!g41) & (!g42) & (g43)) + ((g38) & (g39) & (g40) & (!g41) & (g42) & (!g43)) + ((g38) & (g39) & (g40) & (g41) & (!g42) & (!g43)) + ((g38) & (g39) & (g40) & (g41) & (!g42) & (g43)) + ((g38) & (g39) & (g40) & (g41) & (g42) & (!g43)) + ((g38) & (g39) & (g40) & (g41) & (g42) & (g43)));
	assign g49 = (((!g45) & (!g46) & (!g47) & (g48) & (g42) & (g43)) + ((!g45) & (!g46) & (g47) & (!g48) & (!g42) & (g43)) + ((!g45) & (!g46) & (g47) & (g48) & (!g42) & (g43)) + ((!g45) & (!g46) & (g47) & (g48) & (g42) & (g43)) + ((!g45) & (g46) & (!g47) & (!g48) & (g42) & (!g43)) + ((!g45) & (g46) & (!g47) & (g48) & (g42) & (!g43)) + ((!g45) & (g46) & (!g47) & (g48) & (g42) & (g43)) + ((!g45) & (g46) & (g47) & (!g48) & (!g42) & (g43)) + ((!g45) & (g46) & (g47) & (!g48) & (g42) & (!g43)) + ((!g45) & (g46) & (g47) & (g48) & (!g42) & (g43)) + ((!g45) & (g46) & (g47) & (g48) & (g42) & (!g43)) + ((!g45) & (g46) & (g47) & (g48) & (g42) & (g43)) + ((g45) & (!g46) & (!g47) & (!g48) & (!g42) & (!g43)) + ((g45) & (!g46) & (!g47) & (g48) & (!g42) & (!g43)) + ((g45) & (!g46) & (!g47) & (g48) & (g42) & (g43)) + ((g45) & (!g46) & (g47) & (!g48) & (!g42) & (!g43)) + ((g45) & (!g46) & (g47) & (!g48) & (!g42) & (g43)) + ((g45) & (!g46) & (g47) & (g48) & (!g42) & (!g43)) + ((g45) & (!g46) & (g47) & (g48) & (!g42) & (g43)) + ((g45) & (!g46) & (g47) & (g48) & (g42) & (g43)) + ((g45) & (g46) & (!g47) & (!g48) & (!g42) & (!g43)) + ((g45) & (g46) & (!g47) & (!g48) & (g42) & (!g43)) + ((g45) & (g46) & (!g47) & (g48) & (!g42) & (!g43)) + ((g45) & (g46) & (!g47) & (g48) & (g42) & (!g43)) + ((g45) & (g46) & (!g47) & (g48) & (g42) & (g43)) + ((g45) & (g46) & (g47) & (!g48) & (!g42) & (!g43)) + ((g45) & (g46) & (g47) & (!g48) & (!g42) & (g43)) + ((g45) & (g46) & (g47) & (!g48) & (g42) & (!g43)) + ((g45) & (g46) & (g47) & (g48) & (!g42) & (!g43)) + ((g45) & (g46) & (g47) & (g48) & (!g42) & (g43)) + ((g45) & (g46) & (g47) & (g48) & (g42) & (!g43)) + ((g45) & (g46) & (g47) & (g48) & (g42) & (g43)));
	assign g54 = (((!g50) & (!g51) & (!g52) & (g53) & (g42) & (g43)) + ((!g50) & (!g51) & (g52) & (!g53) & (!g42) & (g43)) + ((!g50) & (!g51) & (g52) & (g53) & (!g42) & (g43)) + ((!g50) & (!g51) & (g52) & (g53) & (g42) & (g43)) + ((!g50) & (g51) & (!g52) & (!g53) & (g42) & (!g43)) + ((!g50) & (g51) & (!g52) & (g53) & (g42) & (!g43)) + ((!g50) & (g51) & (!g52) & (g53) & (g42) & (g43)) + ((!g50) & (g51) & (g52) & (!g53) & (!g42) & (g43)) + ((!g50) & (g51) & (g52) & (!g53) & (g42) & (!g43)) + ((!g50) & (g51) & (g52) & (g53) & (!g42) & (g43)) + ((!g50) & (g51) & (g52) & (g53) & (g42) & (!g43)) + ((!g50) & (g51) & (g52) & (g53) & (g42) & (g43)) + ((g50) & (!g51) & (!g52) & (!g53) & (!g42) & (!g43)) + ((g50) & (!g51) & (!g52) & (g53) & (!g42) & (!g43)) + ((g50) & (!g51) & (!g52) & (g53) & (g42) & (g43)) + ((g50) & (!g51) & (g52) & (!g53) & (!g42) & (!g43)) + ((g50) & (!g51) & (g52) & (!g53) & (!g42) & (g43)) + ((g50) & (!g51) & (g52) & (g53) & (!g42) & (!g43)) + ((g50) & (!g51) & (g52) & (g53) & (!g42) & (g43)) + ((g50) & (!g51) & (g52) & (g53) & (g42) & (g43)) + ((g50) & (g51) & (!g52) & (!g53) & (!g42) & (!g43)) + ((g50) & (g51) & (!g52) & (!g53) & (g42) & (!g43)) + ((g50) & (g51) & (!g52) & (g53) & (!g42) & (!g43)) + ((g50) & (g51) & (!g52) & (g53) & (g42) & (!g43)) + ((g50) & (g51) & (!g52) & (g53) & (g42) & (g43)) + ((g50) & (g51) & (g52) & (!g53) & (!g42) & (!g43)) + ((g50) & (g51) & (g52) & (!g53) & (!g42) & (g43)) + ((g50) & (g51) & (g52) & (!g53) & (g42) & (!g43)) + ((g50) & (g51) & (g52) & (g53) & (!g42) & (!g43)) + ((g50) & (g51) & (g52) & (g53) & (!g42) & (g43)) + ((g50) & (g51) & (g52) & (g53) & (g42) & (!g43)) + ((g50) & (g51) & (g52) & (g53) & (g42) & (g43)));
	assign g59 = (((!g55) & (!g56) & (!g57) & (g58) & (g42) & (g43)) + ((!g55) & (!g56) & (g57) & (!g58) & (!g42) & (g43)) + ((!g55) & (!g56) & (g57) & (g58) & (!g42) & (g43)) + ((!g55) & (!g56) & (g57) & (g58) & (g42) & (g43)) + ((!g55) & (g56) & (!g57) & (!g58) & (g42) & (!g43)) + ((!g55) & (g56) & (!g57) & (g58) & (g42) & (!g43)) + ((!g55) & (g56) & (!g57) & (g58) & (g42) & (g43)) + ((!g55) & (g56) & (g57) & (!g58) & (!g42) & (g43)) + ((!g55) & (g56) & (g57) & (!g58) & (g42) & (!g43)) + ((!g55) & (g56) & (g57) & (g58) & (!g42) & (g43)) + ((!g55) & (g56) & (g57) & (g58) & (g42) & (!g43)) + ((!g55) & (g56) & (g57) & (g58) & (g42) & (g43)) + ((g55) & (!g56) & (!g57) & (!g58) & (!g42) & (!g43)) + ((g55) & (!g56) & (!g57) & (g58) & (!g42) & (!g43)) + ((g55) & (!g56) & (!g57) & (g58) & (g42) & (g43)) + ((g55) & (!g56) & (g57) & (!g58) & (!g42) & (!g43)) + ((g55) & (!g56) & (g57) & (!g58) & (!g42) & (g43)) + ((g55) & (!g56) & (g57) & (g58) & (!g42) & (!g43)) + ((g55) & (!g56) & (g57) & (g58) & (!g42) & (g43)) + ((g55) & (!g56) & (g57) & (g58) & (g42) & (g43)) + ((g55) & (g56) & (!g57) & (!g58) & (!g42) & (!g43)) + ((g55) & (g56) & (!g57) & (!g58) & (g42) & (!g43)) + ((g55) & (g56) & (!g57) & (g58) & (!g42) & (!g43)) + ((g55) & (g56) & (!g57) & (g58) & (g42) & (!g43)) + ((g55) & (g56) & (!g57) & (g58) & (g42) & (g43)) + ((g55) & (g56) & (g57) & (!g58) & (!g42) & (!g43)) + ((g55) & (g56) & (g57) & (!g58) & (!g42) & (g43)) + ((g55) & (g56) & (g57) & (!g58) & (g42) & (!g43)) + ((g55) & (g56) & (g57) & (g58) & (!g42) & (!g43)) + ((g55) & (g56) & (g57) & (g58) & (!g42) & (g43)) + ((g55) & (g56) & (g57) & (g58) & (g42) & (!g43)) + ((g55) & (g56) & (g57) & (g58) & (g42) & (g43)));
	assign g7231 = (((!g797) & (g825) & (!g60)) + ((!g797) & (g825) & (g60)) + ((g797) & (!g825) & (g60)) + ((g797) & (g825) & (g60)));
	assign g7232 = (((!g826)));
	assign g7233 = (((!g797) & (g7232) & (!g61)) + ((!g797) & (g7232) & (g61)) + ((g797) & (!g7232) & (g61)) + ((g797) & (g7232) & (g61)));
	assign g62 = (((!g44) & (!g49) & (!g54) & (g59) & (g60) & (g61)) + ((!g44) & (!g49) & (g54) & (!g59) & (!g60) & (g61)) + ((!g44) & (!g49) & (g54) & (g59) & (!g60) & (g61)) + ((!g44) & (!g49) & (g54) & (g59) & (g60) & (g61)) + ((!g44) & (g49) & (!g54) & (!g59) & (g60) & (!g61)) + ((!g44) & (g49) & (!g54) & (g59) & (g60) & (!g61)) + ((!g44) & (g49) & (!g54) & (g59) & (g60) & (g61)) + ((!g44) & (g49) & (g54) & (!g59) & (!g60) & (g61)) + ((!g44) & (g49) & (g54) & (!g59) & (g60) & (!g61)) + ((!g44) & (g49) & (g54) & (g59) & (!g60) & (g61)) + ((!g44) & (g49) & (g54) & (g59) & (g60) & (!g61)) + ((!g44) & (g49) & (g54) & (g59) & (g60) & (g61)) + ((g44) & (!g49) & (!g54) & (!g59) & (!g60) & (!g61)) + ((g44) & (!g49) & (!g54) & (g59) & (!g60) & (!g61)) + ((g44) & (!g49) & (!g54) & (g59) & (g60) & (g61)) + ((g44) & (!g49) & (g54) & (!g59) & (!g60) & (!g61)) + ((g44) & (!g49) & (g54) & (!g59) & (!g60) & (g61)) + ((g44) & (!g49) & (g54) & (g59) & (!g60) & (!g61)) + ((g44) & (!g49) & (g54) & (g59) & (!g60) & (g61)) + ((g44) & (!g49) & (g54) & (g59) & (g60) & (g61)) + ((g44) & (g49) & (!g54) & (!g59) & (!g60) & (!g61)) + ((g44) & (g49) & (!g54) & (!g59) & (g60) & (!g61)) + ((g44) & (g49) & (!g54) & (g59) & (!g60) & (!g61)) + ((g44) & (g49) & (!g54) & (g59) & (g60) & (!g61)) + ((g44) & (g49) & (!g54) & (g59) & (g60) & (g61)) + ((g44) & (g49) & (g54) & (!g59) & (!g60) & (!g61)) + ((g44) & (g49) & (g54) & (!g59) & (!g60) & (g61)) + ((g44) & (g49) & (g54) & (!g59) & (g60) & (!g61)) + ((g44) & (g49) & (g54) & (g59) & (!g60) & (!g61)) + ((g44) & (g49) & (g54) & (g59) & (!g60) & (g61)) + ((g44) & (g49) & (g54) & (g59) & (g60) & (!g61)) + ((g44) & (g49) & (g54) & (g59) & (g60) & (g61)));
	assign g7234 = (((!g832) & (g829) & (!g63)) + ((!g832) & (g829) & (g63)) + ((g832) & (!g829) & (g63)) + ((g832) & (g829) & (g63)));
	assign g64 = (((!g34) & (!reset) & (!g62) & (g63)) + ((!g34) & (!reset) & (g62) & (g63)) + ((g34) & (!reset) & (g62) & (!g63)) + ((g34) & (!reset) & (g62) & (g63)));
	assign g65 = (((!g34) & (!g35) & (!g36) & (!reset)) + ((!g34) & (!g35) & (g36) & (!reset)) + ((!g34) & (g35) & (!g36) & (!reset)) + ((g34) & (!g35) & (!g36) & (!reset)) + ((g34) & (g35) & (!g36) & (!reset)) + ((g34) & (g35) & (g36) & (!reset)));
	assign g70 = (((!g66) & (!g67) & (!g68) & (g69) & (g60) & (g61)) + ((!g66) & (!g67) & (g68) & (!g69) & (!g60) & (g61)) + ((!g66) & (!g67) & (g68) & (g69) & (!g60) & (g61)) + ((!g66) & (!g67) & (g68) & (g69) & (g60) & (g61)) + ((!g66) & (g67) & (!g68) & (!g69) & (g60) & (!g61)) + ((!g66) & (g67) & (!g68) & (g69) & (g60) & (!g61)) + ((!g66) & (g67) & (!g68) & (g69) & (g60) & (g61)) + ((!g66) & (g67) & (g68) & (!g69) & (!g60) & (g61)) + ((!g66) & (g67) & (g68) & (!g69) & (g60) & (!g61)) + ((!g66) & (g67) & (g68) & (g69) & (!g60) & (g61)) + ((!g66) & (g67) & (g68) & (g69) & (g60) & (!g61)) + ((!g66) & (g67) & (g68) & (g69) & (g60) & (g61)) + ((g66) & (!g67) & (!g68) & (!g69) & (!g60) & (!g61)) + ((g66) & (!g67) & (!g68) & (g69) & (!g60) & (!g61)) + ((g66) & (!g67) & (!g68) & (g69) & (g60) & (g61)) + ((g66) & (!g67) & (g68) & (!g69) & (!g60) & (!g61)) + ((g66) & (!g67) & (g68) & (!g69) & (!g60) & (g61)) + ((g66) & (!g67) & (g68) & (g69) & (!g60) & (!g61)) + ((g66) & (!g67) & (g68) & (g69) & (!g60) & (g61)) + ((g66) & (!g67) & (g68) & (g69) & (g60) & (g61)) + ((g66) & (g67) & (!g68) & (!g69) & (!g60) & (!g61)) + ((g66) & (g67) & (!g68) & (!g69) & (g60) & (!g61)) + ((g66) & (g67) & (!g68) & (g69) & (!g60) & (!g61)) + ((g66) & (g67) & (!g68) & (g69) & (g60) & (!g61)) + ((g66) & (g67) & (!g68) & (g69) & (g60) & (g61)) + ((g66) & (g67) & (g68) & (!g69) & (!g60) & (!g61)) + ((g66) & (g67) & (g68) & (!g69) & (!g60) & (g61)) + ((g66) & (g67) & (g68) & (!g69) & (g60) & (!g61)) + ((g66) & (g67) & (g68) & (g69) & (!g60) & (!g61)) + ((g66) & (g67) & (g68) & (g69) & (!g60) & (g61)) + ((g66) & (g67) & (g68) & (g69) & (g60) & (!g61)) + ((g66) & (g67) & (g68) & (g69) & (g60) & (g61)));
	assign g75 = (((!g71) & (!g72) & (!g73) & (g74) & (g60) & (g61)) + ((!g71) & (!g72) & (g73) & (!g74) & (!g60) & (g61)) + ((!g71) & (!g72) & (g73) & (g74) & (!g60) & (g61)) + ((!g71) & (!g72) & (g73) & (g74) & (g60) & (g61)) + ((!g71) & (g72) & (!g73) & (!g74) & (g60) & (!g61)) + ((!g71) & (g72) & (!g73) & (g74) & (g60) & (!g61)) + ((!g71) & (g72) & (!g73) & (g74) & (g60) & (g61)) + ((!g71) & (g72) & (g73) & (!g74) & (!g60) & (g61)) + ((!g71) & (g72) & (g73) & (!g74) & (g60) & (!g61)) + ((!g71) & (g72) & (g73) & (g74) & (!g60) & (g61)) + ((!g71) & (g72) & (g73) & (g74) & (g60) & (!g61)) + ((!g71) & (g72) & (g73) & (g74) & (g60) & (g61)) + ((g71) & (!g72) & (!g73) & (!g74) & (!g60) & (!g61)) + ((g71) & (!g72) & (!g73) & (g74) & (!g60) & (!g61)) + ((g71) & (!g72) & (!g73) & (g74) & (g60) & (g61)) + ((g71) & (!g72) & (g73) & (!g74) & (!g60) & (!g61)) + ((g71) & (!g72) & (g73) & (!g74) & (!g60) & (g61)) + ((g71) & (!g72) & (g73) & (g74) & (!g60) & (!g61)) + ((g71) & (!g72) & (g73) & (g74) & (!g60) & (g61)) + ((g71) & (!g72) & (g73) & (g74) & (g60) & (g61)) + ((g71) & (g72) & (!g73) & (!g74) & (!g60) & (!g61)) + ((g71) & (g72) & (!g73) & (!g74) & (g60) & (!g61)) + ((g71) & (g72) & (!g73) & (g74) & (!g60) & (!g61)) + ((g71) & (g72) & (!g73) & (g74) & (g60) & (!g61)) + ((g71) & (g72) & (!g73) & (g74) & (g60) & (g61)) + ((g71) & (g72) & (g73) & (!g74) & (!g60) & (!g61)) + ((g71) & (g72) & (g73) & (!g74) & (!g60) & (g61)) + ((g71) & (g72) & (g73) & (!g74) & (g60) & (!g61)) + ((g71) & (g72) & (g73) & (g74) & (!g60) & (!g61)) + ((g71) & (g72) & (g73) & (g74) & (!g60) & (g61)) + ((g71) & (g72) & (g73) & (g74) & (g60) & (!g61)) + ((g71) & (g72) & (g73) & (g74) & (g60) & (g61)));
	assign g80 = (((!g76) & (!g77) & (!g78) & (g79) & (g60) & (g61)) + ((!g76) & (!g77) & (g78) & (!g79) & (!g60) & (g61)) + ((!g76) & (!g77) & (g78) & (g79) & (!g60) & (g61)) + ((!g76) & (!g77) & (g78) & (g79) & (g60) & (g61)) + ((!g76) & (g77) & (!g78) & (!g79) & (g60) & (!g61)) + ((!g76) & (g77) & (!g78) & (g79) & (g60) & (!g61)) + ((!g76) & (g77) & (!g78) & (g79) & (g60) & (g61)) + ((!g76) & (g77) & (g78) & (!g79) & (!g60) & (g61)) + ((!g76) & (g77) & (g78) & (!g79) & (g60) & (!g61)) + ((!g76) & (g77) & (g78) & (g79) & (!g60) & (g61)) + ((!g76) & (g77) & (g78) & (g79) & (g60) & (!g61)) + ((!g76) & (g77) & (g78) & (g79) & (g60) & (g61)) + ((g76) & (!g77) & (!g78) & (!g79) & (!g60) & (!g61)) + ((g76) & (!g77) & (!g78) & (g79) & (!g60) & (!g61)) + ((g76) & (!g77) & (!g78) & (g79) & (g60) & (g61)) + ((g76) & (!g77) & (g78) & (!g79) & (!g60) & (!g61)) + ((g76) & (!g77) & (g78) & (!g79) & (!g60) & (g61)) + ((g76) & (!g77) & (g78) & (g79) & (!g60) & (!g61)) + ((g76) & (!g77) & (g78) & (g79) & (!g60) & (g61)) + ((g76) & (!g77) & (g78) & (g79) & (g60) & (g61)) + ((g76) & (g77) & (!g78) & (!g79) & (!g60) & (!g61)) + ((g76) & (g77) & (!g78) & (!g79) & (g60) & (!g61)) + ((g76) & (g77) & (!g78) & (g79) & (!g60) & (!g61)) + ((g76) & (g77) & (!g78) & (g79) & (g60) & (!g61)) + ((g76) & (g77) & (!g78) & (g79) & (g60) & (g61)) + ((g76) & (g77) & (g78) & (!g79) & (!g60) & (!g61)) + ((g76) & (g77) & (g78) & (!g79) & (!g60) & (g61)) + ((g76) & (g77) & (g78) & (!g79) & (g60) & (!g61)) + ((g76) & (g77) & (g78) & (g79) & (!g60) & (!g61)) + ((g76) & (g77) & (g78) & (g79) & (!g60) & (g61)) + ((g76) & (g77) & (g78) & (g79) & (g60) & (!g61)) + ((g76) & (g77) & (g78) & (g79) & (g60) & (g61)));
	assign g85 = (((!g81) & (!g82) & (!g83) & (g84) & (g60) & (g61)) + ((!g81) & (!g82) & (g83) & (!g84) & (!g60) & (g61)) + ((!g81) & (!g82) & (g83) & (g84) & (!g60) & (g61)) + ((!g81) & (!g82) & (g83) & (g84) & (g60) & (g61)) + ((!g81) & (g82) & (!g83) & (!g84) & (g60) & (!g61)) + ((!g81) & (g82) & (!g83) & (g84) & (g60) & (!g61)) + ((!g81) & (g82) & (!g83) & (g84) & (g60) & (g61)) + ((!g81) & (g82) & (g83) & (!g84) & (!g60) & (g61)) + ((!g81) & (g82) & (g83) & (!g84) & (g60) & (!g61)) + ((!g81) & (g82) & (g83) & (g84) & (!g60) & (g61)) + ((!g81) & (g82) & (g83) & (g84) & (g60) & (!g61)) + ((!g81) & (g82) & (g83) & (g84) & (g60) & (g61)) + ((g81) & (!g82) & (!g83) & (!g84) & (!g60) & (!g61)) + ((g81) & (!g82) & (!g83) & (g84) & (!g60) & (!g61)) + ((g81) & (!g82) & (!g83) & (g84) & (g60) & (g61)) + ((g81) & (!g82) & (g83) & (!g84) & (!g60) & (!g61)) + ((g81) & (!g82) & (g83) & (!g84) & (!g60) & (g61)) + ((g81) & (!g82) & (g83) & (g84) & (!g60) & (!g61)) + ((g81) & (!g82) & (g83) & (g84) & (!g60) & (g61)) + ((g81) & (!g82) & (g83) & (g84) & (g60) & (g61)) + ((g81) & (g82) & (!g83) & (!g84) & (!g60) & (!g61)) + ((g81) & (g82) & (!g83) & (!g84) & (g60) & (!g61)) + ((g81) & (g82) & (!g83) & (g84) & (!g60) & (!g61)) + ((g81) & (g82) & (!g83) & (g84) & (g60) & (!g61)) + ((g81) & (g82) & (!g83) & (g84) & (g60) & (g61)) + ((g81) & (g82) & (g83) & (!g84) & (!g60) & (!g61)) + ((g81) & (g82) & (g83) & (!g84) & (!g60) & (g61)) + ((g81) & (g82) & (g83) & (!g84) & (g60) & (!g61)) + ((g81) & (g82) & (g83) & (g84) & (!g60) & (!g61)) + ((g81) & (g82) & (g83) & (g84) & (!g60) & (g61)) + ((g81) & (g82) & (g83) & (g84) & (g60) & (!g61)) + ((g81) & (g82) & (g83) & (g84) & (g60) & (g61)));
	assign g86 = (((!g70) & (!g75) & (!g80) & (g85) & (g42) & (g43)) + ((!g70) & (!g75) & (g80) & (!g85) & (!g42) & (g43)) + ((!g70) & (!g75) & (g80) & (g85) & (!g42) & (g43)) + ((!g70) & (!g75) & (g80) & (g85) & (g42) & (g43)) + ((!g70) & (g75) & (!g80) & (!g85) & (g42) & (!g43)) + ((!g70) & (g75) & (!g80) & (g85) & (g42) & (!g43)) + ((!g70) & (g75) & (!g80) & (g85) & (g42) & (g43)) + ((!g70) & (g75) & (g80) & (!g85) & (!g42) & (g43)) + ((!g70) & (g75) & (g80) & (!g85) & (g42) & (!g43)) + ((!g70) & (g75) & (g80) & (g85) & (!g42) & (g43)) + ((!g70) & (g75) & (g80) & (g85) & (g42) & (!g43)) + ((!g70) & (g75) & (g80) & (g85) & (g42) & (g43)) + ((g70) & (!g75) & (!g80) & (!g85) & (!g42) & (!g43)) + ((g70) & (!g75) & (!g80) & (g85) & (!g42) & (!g43)) + ((g70) & (!g75) & (!g80) & (g85) & (g42) & (g43)) + ((g70) & (!g75) & (g80) & (!g85) & (!g42) & (!g43)) + ((g70) & (!g75) & (g80) & (!g85) & (!g42) & (g43)) + ((g70) & (!g75) & (g80) & (g85) & (!g42) & (!g43)) + ((g70) & (!g75) & (g80) & (g85) & (!g42) & (g43)) + ((g70) & (!g75) & (g80) & (g85) & (g42) & (g43)) + ((g70) & (g75) & (!g80) & (!g85) & (!g42) & (!g43)) + ((g70) & (g75) & (!g80) & (!g85) & (g42) & (!g43)) + ((g70) & (g75) & (!g80) & (g85) & (!g42) & (!g43)) + ((g70) & (g75) & (!g80) & (g85) & (g42) & (!g43)) + ((g70) & (g75) & (!g80) & (g85) & (g42) & (g43)) + ((g70) & (g75) & (g80) & (!g85) & (!g42) & (!g43)) + ((g70) & (g75) & (g80) & (!g85) & (!g42) & (g43)) + ((g70) & (g75) & (g80) & (!g85) & (g42) & (!g43)) + ((g70) & (g75) & (g80) & (g85) & (!g42) & (!g43)) + ((g70) & (g75) & (g80) & (g85) & (!g42) & (g43)) + ((g70) & (g75) & (g80) & (g85) & (g42) & (!g43)) + ((g70) & (g75) & (g80) & (g85) & (g42) & (g43)));
	assign g7235 = (((!g832) & (g865) & (!g87)) + ((!g832) & (g865) & (g87)) + ((g832) & (!g865) & (g87)) + ((g832) & (g865) & (g87)));
	assign g88 = (((!g34) & (!reset) & (!g86) & (g87)) + ((!g34) & (!reset) & (g86) & (g87)) + ((g34) & (!reset) & (g86) & (!g87)) + ((g34) & (!reset) & (g86) & (g87)));
	assign g93 = (((!g89) & (!g90) & (!g91) & (g92) & (g42) & (g43)) + ((!g89) & (!g90) & (g91) & (!g92) & (!g42) & (g43)) + ((!g89) & (!g90) & (g91) & (g92) & (!g42) & (g43)) + ((!g89) & (!g90) & (g91) & (g92) & (g42) & (g43)) + ((!g89) & (g90) & (!g91) & (!g92) & (g42) & (!g43)) + ((!g89) & (g90) & (!g91) & (g92) & (g42) & (!g43)) + ((!g89) & (g90) & (!g91) & (g92) & (g42) & (g43)) + ((!g89) & (g90) & (g91) & (!g92) & (!g42) & (g43)) + ((!g89) & (g90) & (g91) & (!g92) & (g42) & (!g43)) + ((!g89) & (g90) & (g91) & (g92) & (!g42) & (g43)) + ((!g89) & (g90) & (g91) & (g92) & (g42) & (!g43)) + ((!g89) & (g90) & (g91) & (g92) & (g42) & (g43)) + ((g89) & (!g90) & (!g91) & (!g92) & (!g42) & (!g43)) + ((g89) & (!g90) & (!g91) & (g92) & (!g42) & (!g43)) + ((g89) & (!g90) & (!g91) & (g92) & (g42) & (g43)) + ((g89) & (!g90) & (g91) & (!g92) & (!g42) & (!g43)) + ((g89) & (!g90) & (g91) & (!g92) & (!g42) & (g43)) + ((g89) & (!g90) & (g91) & (g92) & (!g42) & (!g43)) + ((g89) & (!g90) & (g91) & (g92) & (!g42) & (g43)) + ((g89) & (!g90) & (g91) & (g92) & (g42) & (g43)) + ((g89) & (g90) & (!g91) & (!g92) & (!g42) & (!g43)) + ((g89) & (g90) & (!g91) & (!g92) & (g42) & (!g43)) + ((g89) & (g90) & (!g91) & (g92) & (!g42) & (!g43)) + ((g89) & (g90) & (!g91) & (g92) & (g42) & (!g43)) + ((g89) & (g90) & (!g91) & (g92) & (g42) & (g43)) + ((g89) & (g90) & (g91) & (!g92) & (!g42) & (!g43)) + ((g89) & (g90) & (g91) & (!g92) & (!g42) & (g43)) + ((g89) & (g90) & (g91) & (!g92) & (g42) & (!g43)) + ((g89) & (g90) & (g91) & (g92) & (!g42) & (!g43)) + ((g89) & (g90) & (g91) & (g92) & (!g42) & (g43)) + ((g89) & (g90) & (g91) & (g92) & (g42) & (!g43)) + ((g89) & (g90) & (g91) & (g92) & (g42) & (g43)));
	assign g98 = (((!g94) & (!g95) & (!g96) & (g97) & (g42) & (g43)) + ((!g94) & (!g95) & (g96) & (!g97) & (!g42) & (g43)) + ((!g94) & (!g95) & (g96) & (g97) & (!g42) & (g43)) + ((!g94) & (!g95) & (g96) & (g97) & (g42) & (g43)) + ((!g94) & (g95) & (!g96) & (!g97) & (g42) & (!g43)) + ((!g94) & (g95) & (!g96) & (g97) & (g42) & (!g43)) + ((!g94) & (g95) & (!g96) & (g97) & (g42) & (g43)) + ((!g94) & (g95) & (g96) & (!g97) & (!g42) & (g43)) + ((!g94) & (g95) & (g96) & (!g97) & (g42) & (!g43)) + ((!g94) & (g95) & (g96) & (g97) & (!g42) & (g43)) + ((!g94) & (g95) & (g96) & (g97) & (g42) & (!g43)) + ((!g94) & (g95) & (g96) & (g97) & (g42) & (g43)) + ((g94) & (!g95) & (!g96) & (!g97) & (!g42) & (!g43)) + ((g94) & (!g95) & (!g96) & (g97) & (!g42) & (!g43)) + ((g94) & (!g95) & (!g96) & (g97) & (g42) & (g43)) + ((g94) & (!g95) & (g96) & (!g97) & (!g42) & (!g43)) + ((g94) & (!g95) & (g96) & (!g97) & (!g42) & (g43)) + ((g94) & (!g95) & (g96) & (g97) & (!g42) & (!g43)) + ((g94) & (!g95) & (g96) & (g97) & (!g42) & (g43)) + ((g94) & (!g95) & (g96) & (g97) & (g42) & (g43)) + ((g94) & (g95) & (!g96) & (!g97) & (!g42) & (!g43)) + ((g94) & (g95) & (!g96) & (!g97) & (g42) & (!g43)) + ((g94) & (g95) & (!g96) & (g97) & (!g42) & (!g43)) + ((g94) & (g95) & (!g96) & (g97) & (g42) & (!g43)) + ((g94) & (g95) & (!g96) & (g97) & (g42) & (g43)) + ((g94) & (g95) & (g96) & (!g97) & (!g42) & (!g43)) + ((g94) & (g95) & (g96) & (!g97) & (!g42) & (g43)) + ((g94) & (g95) & (g96) & (!g97) & (g42) & (!g43)) + ((g94) & (g95) & (g96) & (g97) & (!g42) & (!g43)) + ((g94) & (g95) & (g96) & (g97) & (!g42) & (g43)) + ((g94) & (g95) & (g96) & (g97) & (g42) & (!g43)) + ((g94) & (g95) & (g96) & (g97) & (g42) & (g43)));
	assign g103 = (((!g99) & (!g100) & (!g101) & (g102) & (g42) & (g43)) + ((!g99) & (!g100) & (g101) & (!g102) & (!g42) & (g43)) + ((!g99) & (!g100) & (g101) & (g102) & (!g42) & (g43)) + ((!g99) & (!g100) & (g101) & (g102) & (g42) & (g43)) + ((!g99) & (g100) & (!g101) & (!g102) & (g42) & (!g43)) + ((!g99) & (g100) & (!g101) & (g102) & (g42) & (!g43)) + ((!g99) & (g100) & (!g101) & (g102) & (g42) & (g43)) + ((!g99) & (g100) & (g101) & (!g102) & (!g42) & (g43)) + ((!g99) & (g100) & (g101) & (!g102) & (g42) & (!g43)) + ((!g99) & (g100) & (g101) & (g102) & (!g42) & (g43)) + ((!g99) & (g100) & (g101) & (g102) & (g42) & (!g43)) + ((!g99) & (g100) & (g101) & (g102) & (g42) & (g43)) + ((g99) & (!g100) & (!g101) & (!g102) & (!g42) & (!g43)) + ((g99) & (!g100) & (!g101) & (g102) & (!g42) & (!g43)) + ((g99) & (!g100) & (!g101) & (g102) & (g42) & (g43)) + ((g99) & (!g100) & (g101) & (!g102) & (!g42) & (!g43)) + ((g99) & (!g100) & (g101) & (!g102) & (!g42) & (g43)) + ((g99) & (!g100) & (g101) & (g102) & (!g42) & (!g43)) + ((g99) & (!g100) & (g101) & (g102) & (!g42) & (g43)) + ((g99) & (!g100) & (g101) & (g102) & (g42) & (g43)) + ((g99) & (g100) & (!g101) & (!g102) & (!g42) & (!g43)) + ((g99) & (g100) & (!g101) & (!g102) & (g42) & (!g43)) + ((g99) & (g100) & (!g101) & (g102) & (!g42) & (!g43)) + ((g99) & (g100) & (!g101) & (g102) & (g42) & (!g43)) + ((g99) & (g100) & (!g101) & (g102) & (g42) & (g43)) + ((g99) & (g100) & (g101) & (!g102) & (!g42) & (!g43)) + ((g99) & (g100) & (g101) & (!g102) & (!g42) & (g43)) + ((g99) & (g100) & (g101) & (!g102) & (g42) & (!g43)) + ((g99) & (g100) & (g101) & (g102) & (!g42) & (!g43)) + ((g99) & (g100) & (g101) & (g102) & (!g42) & (g43)) + ((g99) & (g100) & (g101) & (g102) & (g42) & (!g43)) + ((g99) & (g100) & (g101) & (g102) & (g42) & (g43)));
	assign g108 = (((!g104) & (!g105) & (!g106) & (g107) & (g42) & (g43)) + ((!g104) & (!g105) & (g106) & (!g107) & (!g42) & (g43)) + ((!g104) & (!g105) & (g106) & (g107) & (!g42) & (g43)) + ((!g104) & (!g105) & (g106) & (g107) & (g42) & (g43)) + ((!g104) & (g105) & (!g106) & (!g107) & (g42) & (!g43)) + ((!g104) & (g105) & (!g106) & (g107) & (g42) & (!g43)) + ((!g104) & (g105) & (!g106) & (g107) & (g42) & (g43)) + ((!g104) & (g105) & (g106) & (!g107) & (!g42) & (g43)) + ((!g104) & (g105) & (g106) & (!g107) & (g42) & (!g43)) + ((!g104) & (g105) & (g106) & (g107) & (!g42) & (g43)) + ((!g104) & (g105) & (g106) & (g107) & (g42) & (!g43)) + ((!g104) & (g105) & (g106) & (g107) & (g42) & (g43)) + ((g104) & (!g105) & (!g106) & (!g107) & (!g42) & (!g43)) + ((g104) & (!g105) & (!g106) & (g107) & (!g42) & (!g43)) + ((g104) & (!g105) & (!g106) & (g107) & (g42) & (g43)) + ((g104) & (!g105) & (g106) & (!g107) & (!g42) & (!g43)) + ((g104) & (!g105) & (g106) & (!g107) & (!g42) & (g43)) + ((g104) & (!g105) & (g106) & (g107) & (!g42) & (!g43)) + ((g104) & (!g105) & (g106) & (g107) & (!g42) & (g43)) + ((g104) & (!g105) & (g106) & (g107) & (g42) & (g43)) + ((g104) & (g105) & (!g106) & (!g107) & (!g42) & (!g43)) + ((g104) & (g105) & (!g106) & (!g107) & (g42) & (!g43)) + ((g104) & (g105) & (!g106) & (g107) & (!g42) & (!g43)) + ((g104) & (g105) & (!g106) & (g107) & (g42) & (!g43)) + ((g104) & (g105) & (!g106) & (g107) & (g42) & (g43)) + ((g104) & (g105) & (g106) & (!g107) & (!g42) & (!g43)) + ((g104) & (g105) & (g106) & (!g107) & (!g42) & (g43)) + ((g104) & (g105) & (g106) & (!g107) & (g42) & (!g43)) + ((g104) & (g105) & (g106) & (g107) & (!g42) & (!g43)) + ((g104) & (g105) & (g106) & (g107) & (!g42) & (g43)) + ((g104) & (g105) & (g106) & (g107) & (g42) & (!g43)) + ((g104) & (g105) & (g106) & (g107) & (g42) & (g43)));
	assign g109 = (((!g93) & (!g98) & (!g103) & (g108) & (g60) & (g61)) + ((!g93) & (!g98) & (g103) & (!g108) & (!g60) & (g61)) + ((!g93) & (!g98) & (g103) & (g108) & (!g60) & (g61)) + ((!g93) & (!g98) & (g103) & (g108) & (g60) & (g61)) + ((!g93) & (g98) & (!g103) & (!g108) & (g60) & (!g61)) + ((!g93) & (g98) & (!g103) & (g108) & (g60) & (!g61)) + ((!g93) & (g98) & (!g103) & (g108) & (g60) & (g61)) + ((!g93) & (g98) & (g103) & (!g108) & (!g60) & (g61)) + ((!g93) & (g98) & (g103) & (!g108) & (g60) & (!g61)) + ((!g93) & (g98) & (g103) & (g108) & (!g60) & (g61)) + ((!g93) & (g98) & (g103) & (g108) & (g60) & (!g61)) + ((!g93) & (g98) & (g103) & (g108) & (g60) & (g61)) + ((g93) & (!g98) & (!g103) & (!g108) & (!g60) & (!g61)) + ((g93) & (!g98) & (!g103) & (g108) & (!g60) & (!g61)) + ((g93) & (!g98) & (!g103) & (g108) & (g60) & (g61)) + ((g93) & (!g98) & (g103) & (!g108) & (!g60) & (!g61)) + ((g93) & (!g98) & (g103) & (!g108) & (!g60) & (g61)) + ((g93) & (!g98) & (g103) & (g108) & (!g60) & (!g61)) + ((g93) & (!g98) & (g103) & (g108) & (!g60) & (g61)) + ((g93) & (!g98) & (g103) & (g108) & (g60) & (g61)) + ((g93) & (g98) & (!g103) & (!g108) & (!g60) & (!g61)) + ((g93) & (g98) & (!g103) & (!g108) & (g60) & (!g61)) + ((g93) & (g98) & (!g103) & (g108) & (!g60) & (!g61)) + ((g93) & (g98) & (!g103) & (g108) & (g60) & (!g61)) + ((g93) & (g98) & (!g103) & (g108) & (g60) & (g61)) + ((g93) & (g98) & (g103) & (!g108) & (!g60) & (!g61)) + ((g93) & (g98) & (g103) & (!g108) & (!g60) & (g61)) + ((g93) & (g98) & (g103) & (!g108) & (g60) & (!g61)) + ((g93) & (g98) & (g103) & (g108) & (!g60) & (!g61)) + ((g93) & (g98) & (g103) & (g108) & (!g60) & (g61)) + ((g93) & (g98) & (g103) & (g108) & (g60) & (!g61)) + ((g93) & (g98) & (g103) & (g108) & (g60) & (g61)));
	assign g7236 = (((!g832) & (g899) & (!g110)) + ((!g832) & (g899) & (g110)) + ((g832) & (!g899) & (g110)) + ((g832) & (g899) & (g110)));
	assign g111 = (((!g34) & (!reset) & (!g109) & (g110)) + ((!g34) & (!reset) & (g109) & (g110)) + ((g34) & (!reset) & (g109) & (!g110)) + ((g34) & (!reset) & (g109) & (g110)));
	assign g116 = (((!g112) & (!g113) & (!g114) & (g115) & (g60) & (g61)) + ((!g112) & (!g113) & (g114) & (!g115) & (!g60) & (g61)) + ((!g112) & (!g113) & (g114) & (g115) & (!g60) & (g61)) + ((!g112) & (!g113) & (g114) & (g115) & (g60) & (g61)) + ((!g112) & (g113) & (!g114) & (!g115) & (g60) & (!g61)) + ((!g112) & (g113) & (!g114) & (g115) & (g60) & (!g61)) + ((!g112) & (g113) & (!g114) & (g115) & (g60) & (g61)) + ((!g112) & (g113) & (g114) & (!g115) & (!g60) & (g61)) + ((!g112) & (g113) & (g114) & (!g115) & (g60) & (!g61)) + ((!g112) & (g113) & (g114) & (g115) & (!g60) & (g61)) + ((!g112) & (g113) & (g114) & (g115) & (g60) & (!g61)) + ((!g112) & (g113) & (g114) & (g115) & (g60) & (g61)) + ((g112) & (!g113) & (!g114) & (!g115) & (!g60) & (!g61)) + ((g112) & (!g113) & (!g114) & (g115) & (!g60) & (!g61)) + ((g112) & (!g113) & (!g114) & (g115) & (g60) & (g61)) + ((g112) & (!g113) & (g114) & (!g115) & (!g60) & (!g61)) + ((g112) & (!g113) & (g114) & (!g115) & (!g60) & (g61)) + ((g112) & (!g113) & (g114) & (g115) & (!g60) & (!g61)) + ((g112) & (!g113) & (g114) & (g115) & (!g60) & (g61)) + ((g112) & (!g113) & (g114) & (g115) & (g60) & (g61)) + ((g112) & (g113) & (!g114) & (!g115) & (!g60) & (!g61)) + ((g112) & (g113) & (!g114) & (!g115) & (g60) & (!g61)) + ((g112) & (g113) & (!g114) & (g115) & (!g60) & (!g61)) + ((g112) & (g113) & (!g114) & (g115) & (g60) & (!g61)) + ((g112) & (g113) & (!g114) & (g115) & (g60) & (g61)) + ((g112) & (g113) & (g114) & (!g115) & (!g60) & (!g61)) + ((g112) & (g113) & (g114) & (!g115) & (!g60) & (g61)) + ((g112) & (g113) & (g114) & (!g115) & (g60) & (!g61)) + ((g112) & (g113) & (g114) & (g115) & (!g60) & (!g61)) + ((g112) & (g113) & (g114) & (g115) & (!g60) & (g61)) + ((g112) & (g113) & (g114) & (g115) & (g60) & (!g61)) + ((g112) & (g113) & (g114) & (g115) & (g60) & (g61)));
	assign g121 = (((!g117) & (!g118) & (!g119) & (g120) & (g60) & (g61)) + ((!g117) & (!g118) & (g119) & (!g120) & (!g60) & (g61)) + ((!g117) & (!g118) & (g119) & (g120) & (!g60) & (g61)) + ((!g117) & (!g118) & (g119) & (g120) & (g60) & (g61)) + ((!g117) & (g118) & (!g119) & (!g120) & (g60) & (!g61)) + ((!g117) & (g118) & (!g119) & (g120) & (g60) & (!g61)) + ((!g117) & (g118) & (!g119) & (g120) & (g60) & (g61)) + ((!g117) & (g118) & (g119) & (!g120) & (!g60) & (g61)) + ((!g117) & (g118) & (g119) & (!g120) & (g60) & (!g61)) + ((!g117) & (g118) & (g119) & (g120) & (!g60) & (g61)) + ((!g117) & (g118) & (g119) & (g120) & (g60) & (!g61)) + ((!g117) & (g118) & (g119) & (g120) & (g60) & (g61)) + ((g117) & (!g118) & (!g119) & (!g120) & (!g60) & (!g61)) + ((g117) & (!g118) & (!g119) & (g120) & (!g60) & (!g61)) + ((g117) & (!g118) & (!g119) & (g120) & (g60) & (g61)) + ((g117) & (!g118) & (g119) & (!g120) & (!g60) & (!g61)) + ((g117) & (!g118) & (g119) & (!g120) & (!g60) & (g61)) + ((g117) & (!g118) & (g119) & (g120) & (!g60) & (!g61)) + ((g117) & (!g118) & (g119) & (g120) & (!g60) & (g61)) + ((g117) & (!g118) & (g119) & (g120) & (g60) & (g61)) + ((g117) & (g118) & (!g119) & (!g120) & (!g60) & (!g61)) + ((g117) & (g118) & (!g119) & (!g120) & (g60) & (!g61)) + ((g117) & (g118) & (!g119) & (g120) & (!g60) & (!g61)) + ((g117) & (g118) & (!g119) & (g120) & (g60) & (!g61)) + ((g117) & (g118) & (!g119) & (g120) & (g60) & (g61)) + ((g117) & (g118) & (g119) & (!g120) & (!g60) & (!g61)) + ((g117) & (g118) & (g119) & (!g120) & (!g60) & (g61)) + ((g117) & (g118) & (g119) & (!g120) & (g60) & (!g61)) + ((g117) & (g118) & (g119) & (g120) & (!g60) & (!g61)) + ((g117) & (g118) & (g119) & (g120) & (!g60) & (g61)) + ((g117) & (g118) & (g119) & (g120) & (g60) & (!g61)) + ((g117) & (g118) & (g119) & (g120) & (g60) & (g61)));
	assign g126 = (((!g122) & (!g123) & (!g124) & (g125) & (g60) & (g61)) + ((!g122) & (!g123) & (g124) & (!g125) & (!g60) & (g61)) + ((!g122) & (!g123) & (g124) & (g125) & (!g60) & (g61)) + ((!g122) & (!g123) & (g124) & (g125) & (g60) & (g61)) + ((!g122) & (g123) & (!g124) & (!g125) & (g60) & (!g61)) + ((!g122) & (g123) & (!g124) & (g125) & (g60) & (!g61)) + ((!g122) & (g123) & (!g124) & (g125) & (g60) & (g61)) + ((!g122) & (g123) & (g124) & (!g125) & (!g60) & (g61)) + ((!g122) & (g123) & (g124) & (!g125) & (g60) & (!g61)) + ((!g122) & (g123) & (g124) & (g125) & (!g60) & (g61)) + ((!g122) & (g123) & (g124) & (g125) & (g60) & (!g61)) + ((!g122) & (g123) & (g124) & (g125) & (g60) & (g61)) + ((g122) & (!g123) & (!g124) & (!g125) & (!g60) & (!g61)) + ((g122) & (!g123) & (!g124) & (g125) & (!g60) & (!g61)) + ((g122) & (!g123) & (!g124) & (g125) & (g60) & (g61)) + ((g122) & (!g123) & (g124) & (!g125) & (!g60) & (!g61)) + ((g122) & (!g123) & (g124) & (!g125) & (!g60) & (g61)) + ((g122) & (!g123) & (g124) & (g125) & (!g60) & (!g61)) + ((g122) & (!g123) & (g124) & (g125) & (!g60) & (g61)) + ((g122) & (!g123) & (g124) & (g125) & (g60) & (g61)) + ((g122) & (g123) & (!g124) & (!g125) & (!g60) & (!g61)) + ((g122) & (g123) & (!g124) & (!g125) & (g60) & (!g61)) + ((g122) & (g123) & (!g124) & (g125) & (!g60) & (!g61)) + ((g122) & (g123) & (!g124) & (g125) & (g60) & (!g61)) + ((g122) & (g123) & (!g124) & (g125) & (g60) & (g61)) + ((g122) & (g123) & (g124) & (!g125) & (!g60) & (!g61)) + ((g122) & (g123) & (g124) & (!g125) & (!g60) & (g61)) + ((g122) & (g123) & (g124) & (!g125) & (g60) & (!g61)) + ((g122) & (g123) & (g124) & (g125) & (!g60) & (!g61)) + ((g122) & (g123) & (g124) & (g125) & (!g60) & (g61)) + ((g122) & (g123) & (g124) & (g125) & (g60) & (!g61)) + ((g122) & (g123) & (g124) & (g125) & (g60) & (g61)));
	assign g131 = (((!g127) & (!g128) & (!g129) & (g130) & (g60) & (g61)) + ((!g127) & (!g128) & (g129) & (!g130) & (!g60) & (g61)) + ((!g127) & (!g128) & (g129) & (g130) & (!g60) & (g61)) + ((!g127) & (!g128) & (g129) & (g130) & (g60) & (g61)) + ((!g127) & (g128) & (!g129) & (!g130) & (g60) & (!g61)) + ((!g127) & (g128) & (!g129) & (g130) & (g60) & (!g61)) + ((!g127) & (g128) & (!g129) & (g130) & (g60) & (g61)) + ((!g127) & (g128) & (g129) & (!g130) & (!g60) & (g61)) + ((!g127) & (g128) & (g129) & (!g130) & (g60) & (!g61)) + ((!g127) & (g128) & (g129) & (g130) & (!g60) & (g61)) + ((!g127) & (g128) & (g129) & (g130) & (g60) & (!g61)) + ((!g127) & (g128) & (g129) & (g130) & (g60) & (g61)) + ((g127) & (!g128) & (!g129) & (!g130) & (!g60) & (!g61)) + ((g127) & (!g128) & (!g129) & (g130) & (!g60) & (!g61)) + ((g127) & (!g128) & (!g129) & (g130) & (g60) & (g61)) + ((g127) & (!g128) & (g129) & (!g130) & (!g60) & (!g61)) + ((g127) & (!g128) & (g129) & (!g130) & (!g60) & (g61)) + ((g127) & (!g128) & (g129) & (g130) & (!g60) & (!g61)) + ((g127) & (!g128) & (g129) & (g130) & (!g60) & (g61)) + ((g127) & (!g128) & (g129) & (g130) & (g60) & (g61)) + ((g127) & (g128) & (!g129) & (!g130) & (!g60) & (!g61)) + ((g127) & (g128) & (!g129) & (!g130) & (g60) & (!g61)) + ((g127) & (g128) & (!g129) & (g130) & (!g60) & (!g61)) + ((g127) & (g128) & (!g129) & (g130) & (g60) & (!g61)) + ((g127) & (g128) & (!g129) & (g130) & (g60) & (g61)) + ((g127) & (g128) & (g129) & (!g130) & (!g60) & (!g61)) + ((g127) & (g128) & (g129) & (!g130) & (!g60) & (g61)) + ((g127) & (g128) & (g129) & (!g130) & (g60) & (!g61)) + ((g127) & (g128) & (g129) & (g130) & (!g60) & (!g61)) + ((g127) & (g128) & (g129) & (g130) & (!g60) & (g61)) + ((g127) & (g128) & (g129) & (g130) & (g60) & (!g61)) + ((g127) & (g128) & (g129) & (g130) & (g60) & (g61)));
	assign g132 = (((!g116) & (!g121) & (!g126) & (g131) & (g42) & (g43)) + ((!g116) & (!g121) & (g126) & (!g131) & (!g42) & (g43)) + ((!g116) & (!g121) & (g126) & (g131) & (!g42) & (g43)) + ((!g116) & (!g121) & (g126) & (g131) & (g42) & (g43)) + ((!g116) & (g121) & (!g126) & (!g131) & (g42) & (!g43)) + ((!g116) & (g121) & (!g126) & (g131) & (g42) & (!g43)) + ((!g116) & (g121) & (!g126) & (g131) & (g42) & (g43)) + ((!g116) & (g121) & (g126) & (!g131) & (!g42) & (g43)) + ((!g116) & (g121) & (g126) & (!g131) & (g42) & (!g43)) + ((!g116) & (g121) & (g126) & (g131) & (!g42) & (g43)) + ((!g116) & (g121) & (g126) & (g131) & (g42) & (!g43)) + ((!g116) & (g121) & (g126) & (g131) & (g42) & (g43)) + ((g116) & (!g121) & (!g126) & (!g131) & (!g42) & (!g43)) + ((g116) & (!g121) & (!g126) & (g131) & (!g42) & (!g43)) + ((g116) & (!g121) & (!g126) & (g131) & (g42) & (g43)) + ((g116) & (!g121) & (g126) & (!g131) & (!g42) & (!g43)) + ((g116) & (!g121) & (g126) & (!g131) & (!g42) & (g43)) + ((g116) & (!g121) & (g126) & (g131) & (!g42) & (!g43)) + ((g116) & (!g121) & (g126) & (g131) & (!g42) & (g43)) + ((g116) & (!g121) & (g126) & (g131) & (g42) & (g43)) + ((g116) & (g121) & (!g126) & (!g131) & (!g42) & (!g43)) + ((g116) & (g121) & (!g126) & (!g131) & (g42) & (!g43)) + ((g116) & (g121) & (!g126) & (g131) & (!g42) & (!g43)) + ((g116) & (g121) & (!g126) & (g131) & (g42) & (!g43)) + ((g116) & (g121) & (!g126) & (g131) & (g42) & (g43)) + ((g116) & (g121) & (g126) & (!g131) & (!g42) & (!g43)) + ((g116) & (g121) & (g126) & (!g131) & (!g42) & (g43)) + ((g116) & (g121) & (g126) & (!g131) & (g42) & (!g43)) + ((g116) & (g121) & (g126) & (g131) & (!g42) & (!g43)) + ((g116) & (g121) & (g126) & (g131) & (!g42) & (g43)) + ((g116) & (g121) & (g126) & (g131) & (g42) & (!g43)) + ((g116) & (g121) & (g126) & (g131) & (g42) & (g43)));
	assign g7237 = (((!g832) & (g932) & (!g133)) + ((!g832) & (g932) & (g133)) + ((g832) & (!g932) & (g133)) + ((g832) & (g932) & (g133)));
	assign g134 = (((!g34) & (!reset) & (!g132) & (g133)) + ((!g34) & (!reset) & (g132) & (g133)) + ((g34) & (!reset) & (g132) & (!g133)) + ((g34) & (!reset) & (g132) & (g133)));
	assign g139 = (((!g135) & (!g136) & (!g137) & (g138) & (g42) & (g43)) + ((!g135) & (!g136) & (g137) & (!g138) & (!g42) & (g43)) + ((!g135) & (!g136) & (g137) & (g138) & (!g42) & (g43)) + ((!g135) & (!g136) & (g137) & (g138) & (g42) & (g43)) + ((!g135) & (g136) & (!g137) & (!g138) & (g42) & (!g43)) + ((!g135) & (g136) & (!g137) & (g138) & (g42) & (!g43)) + ((!g135) & (g136) & (!g137) & (g138) & (g42) & (g43)) + ((!g135) & (g136) & (g137) & (!g138) & (!g42) & (g43)) + ((!g135) & (g136) & (g137) & (!g138) & (g42) & (!g43)) + ((!g135) & (g136) & (g137) & (g138) & (!g42) & (g43)) + ((!g135) & (g136) & (g137) & (g138) & (g42) & (!g43)) + ((!g135) & (g136) & (g137) & (g138) & (g42) & (g43)) + ((g135) & (!g136) & (!g137) & (!g138) & (!g42) & (!g43)) + ((g135) & (!g136) & (!g137) & (g138) & (!g42) & (!g43)) + ((g135) & (!g136) & (!g137) & (g138) & (g42) & (g43)) + ((g135) & (!g136) & (g137) & (!g138) & (!g42) & (!g43)) + ((g135) & (!g136) & (g137) & (!g138) & (!g42) & (g43)) + ((g135) & (!g136) & (g137) & (g138) & (!g42) & (!g43)) + ((g135) & (!g136) & (g137) & (g138) & (!g42) & (g43)) + ((g135) & (!g136) & (g137) & (g138) & (g42) & (g43)) + ((g135) & (g136) & (!g137) & (!g138) & (!g42) & (!g43)) + ((g135) & (g136) & (!g137) & (!g138) & (g42) & (!g43)) + ((g135) & (g136) & (!g137) & (g138) & (!g42) & (!g43)) + ((g135) & (g136) & (!g137) & (g138) & (g42) & (!g43)) + ((g135) & (g136) & (!g137) & (g138) & (g42) & (g43)) + ((g135) & (g136) & (g137) & (!g138) & (!g42) & (!g43)) + ((g135) & (g136) & (g137) & (!g138) & (!g42) & (g43)) + ((g135) & (g136) & (g137) & (!g138) & (g42) & (!g43)) + ((g135) & (g136) & (g137) & (g138) & (!g42) & (!g43)) + ((g135) & (g136) & (g137) & (g138) & (!g42) & (g43)) + ((g135) & (g136) & (g137) & (g138) & (g42) & (!g43)) + ((g135) & (g136) & (g137) & (g138) & (g42) & (g43)));
	assign g144 = (((!g140) & (!g141) & (!g142) & (g143) & (g42) & (g43)) + ((!g140) & (!g141) & (g142) & (!g143) & (!g42) & (g43)) + ((!g140) & (!g141) & (g142) & (g143) & (!g42) & (g43)) + ((!g140) & (!g141) & (g142) & (g143) & (g42) & (g43)) + ((!g140) & (g141) & (!g142) & (!g143) & (g42) & (!g43)) + ((!g140) & (g141) & (!g142) & (g143) & (g42) & (!g43)) + ((!g140) & (g141) & (!g142) & (g143) & (g42) & (g43)) + ((!g140) & (g141) & (g142) & (!g143) & (!g42) & (g43)) + ((!g140) & (g141) & (g142) & (!g143) & (g42) & (!g43)) + ((!g140) & (g141) & (g142) & (g143) & (!g42) & (g43)) + ((!g140) & (g141) & (g142) & (g143) & (g42) & (!g43)) + ((!g140) & (g141) & (g142) & (g143) & (g42) & (g43)) + ((g140) & (!g141) & (!g142) & (!g143) & (!g42) & (!g43)) + ((g140) & (!g141) & (!g142) & (g143) & (!g42) & (!g43)) + ((g140) & (!g141) & (!g142) & (g143) & (g42) & (g43)) + ((g140) & (!g141) & (g142) & (!g143) & (!g42) & (!g43)) + ((g140) & (!g141) & (g142) & (!g143) & (!g42) & (g43)) + ((g140) & (!g141) & (g142) & (g143) & (!g42) & (!g43)) + ((g140) & (!g141) & (g142) & (g143) & (!g42) & (g43)) + ((g140) & (!g141) & (g142) & (g143) & (g42) & (g43)) + ((g140) & (g141) & (!g142) & (!g143) & (!g42) & (!g43)) + ((g140) & (g141) & (!g142) & (!g143) & (g42) & (!g43)) + ((g140) & (g141) & (!g142) & (g143) & (!g42) & (!g43)) + ((g140) & (g141) & (!g142) & (g143) & (g42) & (!g43)) + ((g140) & (g141) & (!g142) & (g143) & (g42) & (g43)) + ((g140) & (g141) & (g142) & (!g143) & (!g42) & (!g43)) + ((g140) & (g141) & (g142) & (!g143) & (!g42) & (g43)) + ((g140) & (g141) & (g142) & (!g143) & (g42) & (!g43)) + ((g140) & (g141) & (g142) & (g143) & (!g42) & (!g43)) + ((g140) & (g141) & (g142) & (g143) & (!g42) & (g43)) + ((g140) & (g141) & (g142) & (g143) & (g42) & (!g43)) + ((g140) & (g141) & (g142) & (g143) & (g42) & (g43)));
	assign g149 = (((!g145) & (!g146) & (!g147) & (g148) & (g42) & (g43)) + ((!g145) & (!g146) & (g147) & (!g148) & (!g42) & (g43)) + ((!g145) & (!g146) & (g147) & (g148) & (!g42) & (g43)) + ((!g145) & (!g146) & (g147) & (g148) & (g42) & (g43)) + ((!g145) & (g146) & (!g147) & (!g148) & (g42) & (!g43)) + ((!g145) & (g146) & (!g147) & (g148) & (g42) & (!g43)) + ((!g145) & (g146) & (!g147) & (g148) & (g42) & (g43)) + ((!g145) & (g146) & (g147) & (!g148) & (!g42) & (g43)) + ((!g145) & (g146) & (g147) & (!g148) & (g42) & (!g43)) + ((!g145) & (g146) & (g147) & (g148) & (!g42) & (g43)) + ((!g145) & (g146) & (g147) & (g148) & (g42) & (!g43)) + ((!g145) & (g146) & (g147) & (g148) & (g42) & (g43)) + ((g145) & (!g146) & (!g147) & (!g148) & (!g42) & (!g43)) + ((g145) & (!g146) & (!g147) & (g148) & (!g42) & (!g43)) + ((g145) & (!g146) & (!g147) & (g148) & (g42) & (g43)) + ((g145) & (!g146) & (g147) & (!g148) & (!g42) & (!g43)) + ((g145) & (!g146) & (g147) & (!g148) & (!g42) & (g43)) + ((g145) & (!g146) & (g147) & (g148) & (!g42) & (!g43)) + ((g145) & (!g146) & (g147) & (g148) & (!g42) & (g43)) + ((g145) & (!g146) & (g147) & (g148) & (g42) & (g43)) + ((g145) & (g146) & (!g147) & (!g148) & (!g42) & (!g43)) + ((g145) & (g146) & (!g147) & (!g148) & (g42) & (!g43)) + ((g145) & (g146) & (!g147) & (g148) & (!g42) & (!g43)) + ((g145) & (g146) & (!g147) & (g148) & (g42) & (!g43)) + ((g145) & (g146) & (!g147) & (g148) & (g42) & (g43)) + ((g145) & (g146) & (g147) & (!g148) & (!g42) & (!g43)) + ((g145) & (g146) & (g147) & (!g148) & (!g42) & (g43)) + ((g145) & (g146) & (g147) & (!g148) & (g42) & (!g43)) + ((g145) & (g146) & (g147) & (g148) & (!g42) & (!g43)) + ((g145) & (g146) & (g147) & (g148) & (!g42) & (g43)) + ((g145) & (g146) & (g147) & (g148) & (g42) & (!g43)) + ((g145) & (g146) & (g147) & (g148) & (g42) & (g43)));
	assign g154 = (((!g150) & (!g151) & (!g152) & (g153) & (g42) & (g43)) + ((!g150) & (!g151) & (g152) & (!g153) & (!g42) & (g43)) + ((!g150) & (!g151) & (g152) & (g153) & (!g42) & (g43)) + ((!g150) & (!g151) & (g152) & (g153) & (g42) & (g43)) + ((!g150) & (g151) & (!g152) & (!g153) & (g42) & (!g43)) + ((!g150) & (g151) & (!g152) & (g153) & (g42) & (!g43)) + ((!g150) & (g151) & (!g152) & (g153) & (g42) & (g43)) + ((!g150) & (g151) & (g152) & (!g153) & (!g42) & (g43)) + ((!g150) & (g151) & (g152) & (!g153) & (g42) & (!g43)) + ((!g150) & (g151) & (g152) & (g153) & (!g42) & (g43)) + ((!g150) & (g151) & (g152) & (g153) & (g42) & (!g43)) + ((!g150) & (g151) & (g152) & (g153) & (g42) & (g43)) + ((g150) & (!g151) & (!g152) & (!g153) & (!g42) & (!g43)) + ((g150) & (!g151) & (!g152) & (g153) & (!g42) & (!g43)) + ((g150) & (!g151) & (!g152) & (g153) & (g42) & (g43)) + ((g150) & (!g151) & (g152) & (!g153) & (!g42) & (!g43)) + ((g150) & (!g151) & (g152) & (!g153) & (!g42) & (g43)) + ((g150) & (!g151) & (g152) & (g153) & (!g42) & (!g43)) + ((g150) & (!g151) & (g152) & (g153) & (!g42) & (g43)) + ((g150) & (!g151) & (g152) & (g153) & (g42) & (g43)) + ((g150) & (g151) & (!g152) & (!g153) & (!g42) & (!g43)) + ((g150) & (g151) & (!g152) & (!g153) & (g42) & (!g43)) + ((g150) & (g151) & (!g152) & (g153) & (!g42) & (!g43)) + ((g150) & (g151) & (!g152) & (g153) & (g42) & (!g43)) + ((g150) & (g151) & (!g152) & (g153) & (g42) & (g43)) + ((g150) & (g151) & (g152) & (!g153) & (!g42) & (!g43)) + ((g150) & (g151) & (g152) & (!g153) & (!g42) & (g43)) + ((g150) & (g151) & (g152) & (!g153) & (g42) & (!g43)) + ((g150) & (g151) & (g152) & (g153) & (!g42) & (!g43)) + ((g150) & (g151) & (g152) & (g153) & (!g42) & (g43)) + ((g150) & (g151) & (g152) & (g153) & (g42) & (!g43)) + ((g150) & (g151) & (g152) & (g153) & (g42) & (g43)));
	assign g155 = (((!g139) & (!g144) & (!g149) & (g154) & (g60) & (g61)) + ((!g139) & (!g144) & (g149) & (!g154) & (!g60) & (g61)) + ((!g139) & (!g144) & (g149) & (g154) & (!g60) & (g61)) + ((!g139) & (!g144) & (g149) & (g154) & (g60) & (g61)) + ((!g139) & (g144) & (!g149) & (!g154) & (g60) & (!g61)) + ((!g139) & (g144) & (!g149) & (g154) & (g60) & (!g61)) + ((!g139) & (g144) & (!g149) & (g154) & (g60) & (g61)) + ((!g139) & (g144) & (g149) & (!g154) & (!g60) & (g61)) + ((!g139) & (g144) & (g149) & (!g154) & (g60) & (!g61)) + ((!g139) & (g144) & (g149) & (g154) & (!g60) & (g61)) + ((!g139) & (g144) & (g149) & (g154) & (g60) & (!g61)) + ((!g139) & (g144) & (g149) & (g154) & (g60) & (g61)) + ((g139) & (!g144) & (!g149) & (!g154) & (!g60) & (!g61)) + ((g139) & (!g144) & (!g149) & (g154) & (!g60) & (!g61)) + ((g139) & (!g144) & (!g149) & (g154) & (g60) & (g61)) + ((g139) & (!g144) & (g149) & (!g154) & (!g60) & (!g61)) + ((g139) & (!g144) & (g149) & (!g154) & (!g60) & (g61)) + ((g139) & (!g144) & (g149) & (g154) & (!g60) & (!g61)) + ((g139) & (!g144) & (g149) & (g154) & (!g60) & (g61)) + ((g139) & (!g144) & (g149) & (g154) & (g60) & (g61)) + ((g139) & (g144) & (!g149) & (!g154) & (!g60) & (!g61)) + ((g139) & (g144) & (!g149) & (!g154) & (g60) & (!g61)) + ((g139) & (g144) & (!g149) & (g154) & (!g60) & (!g61)) + ((g139) & (g144) & (!g149) & (g154) & (g60) & (!g61)) + ((g139) & (g144) & (!g149) & (g154) & (g60) & (g61)) + ((g139) & (g144) & (g149) & (!g154) & (!g60) & (!g61)) + ((g139) & (g144) & (g149) & (!g154) & (!g60) & (g61)) + ((g139) & (g144) & (g149) & (!g154) & (g60) & (!g61)) + ((g139) & (g144) & (g149) & (g154) & (!g60) & (!g61)) + ((g139) & (g144) & (g149) & (g154) & (!g60) & (g61)) + ((g139) & (g144) & (g149) & (g154) & (g60) & (!g61)) + ((g139) & (g144) & (g149) & (g154) & (g60) & (g61)));
	assign g7238 = (((!g832) & (g966) & (!g156)) + ((!g832) & (g966) & (g156)) + ((g832) & (!g966) & (g156)) + ((g832) & (g966) & (g156)));
	assign g157 = (((!g34) & (!reset) & (!g155) & (g156)) + ((!g34) & (!reset) & (g155) & (g156)) + ((g34) & (!reset) & (g155) & (!g156)) + ((g34) & (!reset) & (g155) & (g156)));
	assign g162 = (((!g158) & (!g159) & (!g160) & (g161) & (g60) & (g61)) + ((!g158) & (!g159) & (g160) & (!g161) & (!g60) & (g61)) + ((!g158) & (!g159) & (g160) & (g161) & (!g60) & (g61)) + ((!g158) & (!g159) & (g160) & (g161) & (g60) & (g61)) + ((!g158) & (g159) & (!g160) & (!g161) & (g60) & (!g61)) + ((!g158) & (g159) & (!g160) & (g161) & (g60) & (!g61)) + ((!g158) & (g159) & (!g160) & (g161) & (g60) & (g61)) + ((!g158) & (g159) & (g160) & (!g161) & (!g60) & (g61)) + ((!g158) & (g159) & (g160) & (!g161) & (g60) & (!g61)) + ((!g158) & (g159) & (g160) & (g161) & (!g60) & (g61)) + ((!g158) & (g159) & (g160) & (g161) & (g60) & (!g61)) + ((!g158) & (g159) & (g160) & (g161) & (g60) & (g61)) + ((g158) & (!g159) & (!g160) & (!g161) & (!g60) & (!g61)) + ((g158) & (!g159) & (!g160) & (g161) & (!g60) & (!g61)) + ((g158) & (!g159) & (!g160) & (g161) & (g60) & (g61)) + ((g158) & (!g159) & (g160) & (!g161) & (!g60) & (!g61)) + ((g158) & (!g159) & (g160) & (!g161) & (!g60) & (g61)) + ((g158) & (!g159) & (g160) & (g161) & (!g60) & (!g61)) + ((g158) & (!g159) & (g160) & (g161) & (!g60) & (g61)) + ((g158) & (!g159) & (g160) & (g161) & (g60) & (g61)) + ((g158) & (g159) & (!g160) & (!g161) & (!g60) & (!g61)) + ((g158) & (g159) & (!g160) & (!g161) & (g60) & (!g61)) + ((g158) & (g159) & (!g160) & (g161) & (!g60) & (!g61)) + ((g158) & (g159) & (!g160) & (g161) & (g60) & (!g61)) + ((g158) & (g159) & (!g160) & (g161) & (g60) & (g61)) + ((g158) & (g159) & (g160) & (!g161) & (!g60) & (!g61)) + ((g158) & (g159) & (g160) & (!g161) & (!g60) & (g61)) + ((g158) & (g159) & (g160) & (!g161) & (g60) & (!g61)) + ((g158) & (g159) & (g160) & (g161) & (!g60) & (!g61)) + ((g158) & (g159) & (g160) & (g161) & (!g60) & (g61)) + ((g158) & (g159) & (g160) & (g161) & (g60) & (!g61)) + ((g158) & (g159) & (g160) & (g161) & (g60) & (g61)));
	assign g167 = (((!g163) & (!g164) & (!g165) & (g166) & (g60) & (g61)) + ((!g163) & (!g164) & (g165) & (!g166) & (!g60) & (g61)) + ((!g163) & (!g164) & (g165) & (g166) & (!g60) & (g61)) + ((!g163) & (!g164) & (g165) & (g166) & (g60) & (g61)) + ((!g163) & (g164) & (!g165) & (!g166) & (g60) & (!g61)) + ((!g163) & (g164) & (!g165) & (g166) & (g60) & (!g61)) + ((!g163) & (g164) & (!g165) & (g166) & (g60) & (g61)) + ((!g163) & (g164) & (g165) & (!g166) & (!g60) & (g61)) + ((!g163) & (g164) & (g165) & (!g166) & (g60) & (!g61)) + ((!g163) & (g164) & (g165) & (g166) & (!g60) & (g61)) + ((!g163) & (g164) & (g165) & (g166) & (g60) & (!g61)) + ((!g163) & (g164) & (g165) & (g166) & (g60) & (g61)) + ((g163) & (!g164) & (!g165) & (!g166) & (!g60) & (!g61)) + ((g163) & (!g164) & (!g165) & (g166) & (!g60) & (!g61)) + ((g163) & (!g164) & (!g165) & (g166) & (g60) & (g61)) + ((g163) & (!g164) & (g165) & (!g166) & (!g60) & (!g61)) + ((g163) & (!g164) & (g165) & (!g166) & (!g60) & (g61)) + ((g163) & (!g164) & (g165) & (g166) & (!g60) & (!g61)) + ((g163) & (!g164) & (g165) & (g166) & (!g60) & (g61)) + ((g163) & (!g164) & (g165) & (g166) & (g60) & (g61)) + ((g163) & (g164) & (!g165) & (!g166) & (!g60) & (!g61)) + ((g163) & (g164) & (!g165) & (!g166) & (g60) & (!g61)) + ((g163) & (g164) & (!g165) & (g166) & (!g60) & (!g61)) + ((g163) & (g164) & (!g165) & (g166) & (g60) & (!g61)) + ((g163) & (g164) & (!g165) & (g166) & (g60) & (g61)) + ((g163) & (g164) & (g165) & (!g166) & (!g60) & (!g61)) + ((g163) & (g164) & (g165) & (!g166) & (!g60) & (g61)) + ((g163) & (g164) & (g165) & (!g166) & (g60) & (!g61)) + ((g163) & (g164) & (g165) & (g166) & (!g60) & (!g61)) + ((g163) & (g164) & (g165) & (g166) & (!g60) & (g61)) + ((g163) & (g164) & (g165) & (g166) & (g60) & (!g61)) + ((g163) & (g164) & (g165) & (g166) & (g60) & (g61)));
	assign g172 = (((!g168) & (!g169) & (!g170) & (g171) & (g60) & (g61)) + ((!g168) & (!g169) & (g170) & (!g171) & (!g60) & (g61)) + ((!g168) & (!g169) & (g170) & (g171) & (!g60) & (g61)) + ((!g168) & (!g169) & (g170) & (g171) & (g60) & (g61)) + ((!g168) & (g169) & (!g170) & (!g171) & (g60) & (!g61)) + ((!g168) & (g169) & (!g170) & (g171) & (g60) & (!g61)) + ((!g168) & (g169) & (!g170) & (g171) & (g60) & (g61)) + ((!g168) & (g169) & (g170) & (!g171) & (!g60) & (g61)) + ((!g168) & (g169) & (g170) & (!g171) & (g60) & (!g61)) + ((!g168) & (g169) & (g170) & (g171) & (!g60) & (g61)) + ((!g168) & (g169) & (g170) & (g171) & (g60) & (!g61)) + ((!g168) & (g169) & (g170) & (g171) & (g60) & (g61)) + ((g168) & (!g169) & (!g170) & (!g171) & (!g60) & (!g61)) + ((g168) & (!g169) & (!g170) & (g171) & (!g60) & (!g61)) + ((g168) & (!g169) & (!g170) & (g171) & (g60) & (g61)) + ((g168) & (!g169) & (g170) & (!g171) & (!g60) & (!g61)) + ((g168) & (!g169) & (g170) & (!g171) & (!g60) & (g61)) + ((g168) & (!g169) & (g170) & (g171) & (!g60) & (!g61)) + ((g168) & (!g169) & (g170) & (g171) & (!g60) & (g61)) + ((g168) & (!g169) & (g170) & (g171) & (g60) & (g61)) + ((g168) & (g169) & (!g170) & (!g171) & (!g60) & (!g61)) + ((g168) & (g169) & (!g170) & (!g171) & (g60) & (!g61)) + ((g168) & (g169) & (!g170) & (g171) & (!g60) & (!g61)) + ((g168) & (g169) & (!g170) & (g171) & (g60) & (!g61)) + ((g168) & (g169) & (!g170) & (g171) & (g60) & (g61)) + ((g168) & (g169) & (g170) & (!g171) & (!g60) & (!g61)) + ((g168) & (g169) & (g170) & (!g171) & (!g60) & (g61)) + ((g168) & (g169) & (g170) & (!g171) & (g60) & (!g61)) + ((g168) & (g169) & (g170) & (g171) & (!g60) & (!g61)) + ((g168) & (g169) & (g170) & (g171) & (!g60) & (g61)) + ((g168) & (g169) & (g170) & (g171) & (g60) & (!g61)) + ((g168) & (g169) & (g170) & (g171) & (g60) & (g61)));
	assign g177 = (((!g173) & (!g174) & (!g175) & (g176) & (g60) & (g61)) + ((!g173) & (!g174) & (g175) & (!g176) & (!g60) & (g61)) + ((!g173) & (!g174) & (g175) & (g176) & (!g60) & (g61)) + ((!g173) & (!g174) & (g175) & (g176) & (g60) & (g61)) + ((!g173) & (g174) & (!g175) & (!g176) & (g60) & (!g61)) + ((!g173) & (g174) & (!g175) & (g176) & (g60) & (!g61)) + ((!g173) & (g174) & (!g175) & (g176) & (g60) & (g61)) + ((!g173) & (g174) & (g175) & (!g176) & (!g60) & (g61)) + ((!g173) & (g174) & (g175) & (!g176) & (g60) & (!g61)) + ((!g173) & (g174) & (g175) & (g176) & (!g60) & (g61)) + ((!g173) & (g174) & (g175) & (g176) & (g60) & (!g61)) + ((!g173) & (g174) & (g175) & (g176) & (g60) & (g61)) + ((g173) & (!g174) & (!g175) & (!g176) & (!g60) & (!g61)) + ((g173) & (!g174) & (!g175) & (g176) & (!g60) & (!g61)) + ((g173) & (!g174) & (!g175) & (g176) & (g60) & (g61)) + ((g173) & (!g174) & (g175) & (!g176) & (!g60) & (!g61)) + ((g173) & (!g174) & (g175) & (!g176) & (!g60) & (g61)) + ((g173) & (!g174) & (g175) & (g176) & (!g60) & (!g61)) + ((g173) & (!g174) & (g175) & (g176) & (!g60) & (g61)) + ((g173) & (!g174) & (g175) & (g176) & (g60) & (g61)) + ((g173) & (g174) & (!g175) & (!g176) & (!g60) & (!g61)) + ((g173) & (g174) & (!g175) & (!g176) & (g60) & (!g61)) + ((g173) & (g174) & (!g175) & (g176) & (!g60) & (!g61)) + ((g173) & (g174) & (!g175) & (g176) & (g60) & (!g61)) + ((g173) & (g174) & (!g175) & (g176) & (g60) & (g61)) + ((g173) & (g174) & (g175) & (!g176) & (!g60) & (!g61)) + ((g173) & (g174) & (g175) & (!g176) & (!g60) & (g61)) + ((g173) & (g174) & (g175) & (!g176) & (g60) & (!g61)) + ((g173) & (g174) & (g175) & (g176) & (!g60) & (!g61)) + ((g173) & (g174) & (g175) & (g176) & (!g60) & (g61)) + ((g173) & (g174) & (g175) & (g176) & (g60) & (!g61)) + ((g173) & (g174) & (g175) & (g176) & (g60) & (g61)));
	assign g178 = (((!g162) & (!g167) & (!g172) & (g177) & (g42) & (g43)) + ((!g162) & (!g167) & (g172) & (!g177) & (!g42) & (g43)) + ((!g162) & (!g167) & (g172) & (g177) & (!g42) & (g43)) + ((!g162) & (!g167) & (g172) & (g177) & (g42) & (g43)) + ((!g162) & (g167) & (!g172) & (!g177) & (g42) & (!g43)) + ((!g162) & (g167) & (!g172) & (g177) & (g42) & (!g43)) + ((!g162) & (g167) & (!g172) & (g177) & (g42) & (g43)) + ((!g162) & (g167) & (g172) & (!g177) & (!g42) & (g43)) + ((!g162) & (g167) & (g172) & (!g177) & (g42) & (!g43)) + ((!g162) & (g167) & (g172) & (g177) & (!g42) & (g43)) + ((!g162) & (g167) & (g172) & (g177) & (g42) & (!g43)) + ((!g162) & (g167) & (g172) & (g177) & (g42) & (g43)) + ((g162) & (!g167) & (!g172) & (!g177) & (!g42) & (!g43)) + ((g162) & (!g167) & (!g172) & (g177) & (!g42) & (!g43)) + ((g162) & (!g167) & (!g172) & (g177) & (g42) & (g43)) + ((g162) & (!g167) & (g172) & (!g177) & (!g42) & (!g43)) + ((g162) & (!g167) & (g172) & (!g177) & (!g42) & (g43)) + ((g162) & (!g167) & (g172) & (g177) & (!g42) & (!g43)) + ((g162) & (!g167) & (g172) & (g177) & (!g42) & (g43)) + ((g162) & (!g167) & (g172) & (g177) & (g42) & (g43)) + ((g162) & (g167) & (!g172) & (!g177) & (!g42) & (!g43)) + ((g162) & (g167) & (!g172) & (!g177) & (g42) & (!g43)) + ((g162) & (g167) & (!g172) & (g177) & (!g42) & (!g43)) + ((g162) & (g167) & (!g172) & (g177) & (g42) & (!g43)) + ((g162) & (g167) & (!g172) & (g177) & (g42) & (g43)) + ((g162) & (g167) & (g172) & (!g177) & (!g42) & (!g43)) + ((g162) & (g167) & (g172) & (!g177) & (!g42) & (g43)) + ((g162) & (g167) & (g172) & (!g177) & (g42) & (!g43)) + ((g162) & (g167) & (g172) & (g177) & (!g42) & (!g43)) + ((g162) & (g167) & (g172) & (g177) & (!g42) & (g43)) + ((g162) & (g167) & (g172) & (g177) & (g42) & (!g43)) + ((g162) & (g167) & (g172) & (g177) & (g42) & (g43)));
	assign g7239 = (((!g832) & (g999) & (!g179)) + ((!g832) & (g999) & (g179)) + ((g832) & (!g999) & (g179)) + ((g832) & (g999) & (g179)));
	assign g180 = (((!g34) & (!reset) & (!g178) & (g179)) + ((!g34) & (!reset) & (g178) & (g179)) + ((g34) & (!reset) & (g178) & (!g179)) + ((g34) & (!reset) & (g178) & (g179)));
	assign g185 = (((!g181) & (!g182) & (!g183) & (g184) & (g42) & (g43)) + ((!g181) & (!g182) & (g183) & (!g184) & (!g42) & (g43)) + ((!g181) & (!g182) & (g183) & (g184) & (!g42) & (g43)) + ((!g181) & (!g182) & (g183) & (g184) & (g42) & (g43)) + ((!g181) & (g182) & (!g183) & (!g184) & (g42) & (!g43)) + ((!g181) & (g182) & (!g183) & (g184) & (g42) & (!g43)) + ((!g181) & (g182) & (!g183) & (g184) & (g42) & (g43)) + ((!g181) & (g182) & (g183) & (!g184) & (!g42) & (g43)) + ((!g181) & (g182) & (g183) & (!g184) & (g42) & (!g43)) + ((!g181) & (g182) & (g183) & (g184) & (!g42) & (g43)) + ((!g181) & (g182) & (g183) & (g184) & (g42) & (!g43)) + ((!g181) & (g182) & (g183) & (g184) & (g42) & (g43)) + ((g181) & (!g182) & (!g183) & (!g184) & (!g42) & (!g43)) + ((g181) & (!g182) & (!g183) & (g184) & (!g42) & (!g43)) + ((g181) & (!g182) & (!g183) & (g184) & (g42) & (g43)) + ((g181) & (!g182) & (g183) & (!g184) & (!g42) & (!g43)) + ((g181) & (!g182) & (g183) & (!g184) & (!g42) & (g43)) + ((g181) & (!g182) & (g183) & (g184) & (!g42) & (!g43)) + ((g181) & (!g182) & (g183) & (g184) & (!g42) & (g43)) + ((g181) & (!g182) & (g183) & (g184) & (g42) & (g43)) + ((g181) & (g182) & (!g183) & (!g184) & (!g42) & (!g43)) + ((g181) & (g182) & (!g183) & (!g184) & (g42) & (!g43)) + ((g181) & (g182) & (!g183) & (g184) & (!g42) & (!g43)) + ((g181) & (g182) & (!g183) & (g184) & (g42) & (!g43)) + ((g181) & (g182) & (!g183) & (g184) & (g42) & (g43)) + ((g181) & (g182) & (g183) & (!g184) & (!g42) & (!g43)) + ((g181) & (g182) & (g183) & (!g184) & (!g42) & (g43)) + ((g181) & (g182) & (g183) & (!g184) & (g42) & (!g43)) + ((g181) & (g182) & (g183) & (g184) & (!g42) & (!g43)) + ((g181) & (g182) & (g183) & (g184) & (!g42) & (g43)) + ((g181) & (g182) & (g183) & (g184) & (g42) & (!g43)) + ((g181) & (g182) & (g183) & (g184) & (g42) & (g43)));
	assign g190 = (((!g186) & (!g187) & (!g188) & (g189) & (g42) & (g43)) + ((!g186) & (!g187) & (g188) & (!g189) & (!g42) & (g43)) + ((!g186) & (!g187) & (g188) & (g189) & (!g42) & (g43)) + ((!g186) & (!g187) & (g188) & (g189) & (g42) & (g43)) + ((!g186) & (g187) & (!g188) & (!g189) & (g42) & (!g43)) + ((!g186) & (g187) & (!g188) & (g189) & (g42) & (!g43)) + ((!g186) & (g187) & (!g188) & (g189) & (g42) & (g43)) + ((!g186) & (g187) & (g188) & (!g189) & (!g42) & (g43)) + ((!g186) & (g187) & (g188) & (!g189) & (g42) & (!g43)) + ((!g186) & (g187) & (g188) & (g189) & (!g42) & (g43)) + ((!g186) & (g187) & (g188) & (g189) & (g42) & (!g43)) + ((!g186) & (g187) & (g188) & (g189) & (g42) & (g43)) + ((g186) & (!g187) & (!g188) & (!g189) & (!g42) & (!g43)) + ((g186) & (!g187) & (!g188) & (g189) & (!g42) & (!g43)) + ((g186) & (!g187) & (!g188) & (g189) & (g42) & (g43)) + ((g186) & (!g187) & (g188) & (!g189) & (!g42) & (!g43)) + ((g186) & (!g187) & (g188) & (!g189) & (!g42) & (g43)) + ((g186) & (!g187) & (g188) & (g189) & (!g42) & (!g43)) + ((g186) & (!g187) & (g188) & (g189) & (!g42) & (g43)) + ((g186) & (!g187) & (g188) & (g189) & (g42) & (g43)) + ((g186) & (g187) & (!g188) & (!g189) & (!g42) & (!g43)) + ((g186) & (g187) & (!g188) & (!g189) & (g42) & (!g43)) + ((g186) & (g187) & (!g188) & (g189) & (!g42) & (!g43)) + ((g186) & (g187) & (!g188) & (g189) & (g42) & (!g43)) + ((g186) & (g187) & (!g188) & (g189) & (g42) & (g43)) + ((g186) & (g187) & (g188) & (!g189) & (!g42) & (!g43)) + ((g186) & (g187) & (g188) & (!g189) & (!g42) & (g43)) + ((g186) & (g187) & (g188) & (!g189) & (g42) & (!g43)) + ((g186) & (g187) & (g188) & (g189) & (!g42) & (!g43)) + ((g186) & (g187) & (g188) & (g189) & (!g42) & (g43)) + ((g186) & (g187) & (g188) & (g189) & (g42) & (!g43)) + ((g186) & (g187) & (g188) & (g189) & (g42) & (g43)));
	assign g195 = (((!g191) & (!g192) & (!g193) & (g194) & (g42) & (g43)) + ((!g191) & (!g192) & (g193) & (!g194) & (!g42) & (g43)) + ((!g191) & (!g192) & (g193) & (g194) & (!g42) & (g43)) + ((!g191) & (!g192) & (g193) & (g194) & (g42) & (g43)) + ((!g191) & (g192) & (!g193) & (!g194) & (g42) & (!g43)) + ((!g191) & (g192) & (!g193) & (g194) & (g42) & (!g43)) + ((!g191) & (g192) & (!g193) & (g194) & (g42) & (g43)) + ((!g191) & (g192) & (g193) & (!g194) & (!g42) & (g43)) + ((!g191) & (g192) & (g193) & (!g194) & (g42) & (!g43)) + ((!g191) & (g192) & (g193) & (g194) & (!g42) & (g43)) + ((!g191) & (g192) & (g193) & (g194) & (g42) & (!g43)) + ((!g191) & (g192) & (g193) & (g194) & (g42) & (g43)) + ((g191) & (!g192) & (!g193) & (!g194) & (!g42) & (!g43)) + ((g191) & (!g192) & (!g193) & (g194) & (!g42) & (!g43)) + ((g191) & (!g192) & (!g193) & (g194) & (g42) & (g43)) + ((g191) & (!g192) & (g193) & (!g194) & (!g42) & (!g43)) + ((g191) & (!g192) & (g193) & (!g194) & (!g42) & (g43)) + ((g191) & (!g192) & (g193) & (g194) & (!g42) & (!g43)) + ((g191) & (!g192) & (g193) & (g194) & (!g42) & (g43)) + ((g191) & (!g192) & (g193) & (g194) & (g42) & (g43)) + ((g191) & (g192) & (!g193) & (!g194) & (!g42) & (!g43)) + ((g191) & (g192) & (!g193) & (!g194) & (g42) & (!g43)) + ((g191) & (g192) & (!g193) & (g194) & (!g42) & (!g43)) + ((g191) & (g192) & (!g193) & (g194) & (g42) & (!g43)) + ((g191) & (g192) & (!g193) & (g194) & (g42) & (g43)) + ((g191) & (g192) & (g193) & (!g194) & (!g42) & (!g43)) + ((g191) & (g192) & (g193) & (!g194) & (!g42) & (g43)) + ((g191) & (g192) & (g193) & (!g194) & (g42) & (!g43)) + ((g191) & (g192) & (g193) & (g194) & (!g42) & (!g43)) + ((g191) & (g192) & (g193) & (g194) & (!g42) & (g43)) + ((g191) & (g192) & (g193) & (g194) & (g42) & (!g43)) + ((g191) & (g192) & (g193) & (g194) & (g42) & (g43)));
	assign g200 = (((!g196) & (!g197) & (!g198) & (g199) & (g42) & (g43)) + ((!g196) & (!g197) & (g198) & (!g199) & (!g42) & (g43)) + ((!g196) & (!g197) & (g198) & (g199) & (!g42) & (g43)) + ((!g196) & (!g197) & (g198) & (g199) & (g42) & (g43)) + ((!g196) & (g197) & (!g198) & (!g199) & (g42) & (!g43)) + ((!g196) & (g197) & (!g198) & (g199) & (g42) & (!g43)) + ((!g196) & (g197) & (!g198) & (g199) & (g42) & (g43)) + ((!g196) & (g197) & (g198) & (!g199) & (!g42) & (g43)) + ((!g196) & (g197) & (g198) & (!g199) & (g42) & (!g43)) + ((!g196) & (g197) & (g198) & (g199) & (!g42) & (g43)) + ((!g196) & (g197) & (g198) & (g199) & (g42) & (!g43)) + ((!g196) & (g197) & (g198) & (g199) & (g42) & (g43)) + ((g196) & (!g197) & (!g198) & (!g199) & (!g42) & (!g43)) + ((g196) & (!g197) & (!g198) & (g199) & (!g42) & (!g43)) + ((g196) & (!g197) & (!g198) & (g199) & (g42) & (g43)) + ((g196) & (!g197) & (g198) & (!g199) & (!g42) & (!g43)) + ((g196) & (!g197) & (g198) & (!g199) & (!g42) & (g43)) + ((g196) & (!g197) & (g198) & (g199) & (!g42) & (!g43)) + ((g196) & (!g197) & (g198) & (g199) & (!g42) & (g43)) + ((g196) & (!g197) & (g198) & (g199) & (g42) & (g43)) + ((g196) & (g197) & (!g198) & (!g199) & (!g42) & (!g43)) + ((g196) & (g197) & (!g198) & (!g199) & (g42) & (!g43)) + ((g196) & (g197) & (!g198) & (g199) & (!g42) & (!g43)) + ((g196) & (g197) & (!g198) & (g199) & (g42) & (!g43)) + ((g196) & (g197) & (!g198) & (g199) & (g42) & (g43)) + ((g196) & (g197) & (g198) & (!g199) & (!g42) & (!g43)) + ((g196) & (g197) & (g198) & (!g199) & (!g42) & (g43)) + ((g196) & (g197) & (g198) & (!g199) & (g42) & (!g43)) + ((g196) & (g197) & (g198) & (g199) & (!g42) & (!g43)) + ((g196) & (g197) & (g198) & (g199) & (!g42) & (g43)) + ((g196) & (g197) & (g198) & (g199) & (g42) & (!g43)) + ((g196) & (g197) & (g198) & (g199) & (g42) & (g43)));
	assign g201 = (((!g185) & (!g190) & (!g195) & (g200) & (g60) & (g61)) + ((!g185) & (!g190) & (g195) & (!g200) & (!g60) & (g61)) + ((!g185) & (!g190) & (g195) & (g200) & (!g60) & (g61)) + ((!g185) & (!g190) & (g195) & (g200) & (g60) & (g61)) + ((!g185) & (g190) & (!g195) & (!g200) & (g60) & (!g61)) + ((!g185) & (g190) & (!g195) & (g200) & (g60) & (!g61)) + ((!g185) & (g190) & (!g195) & (g200) & (g60) & (g61)) + ((!g185) & (g190) & (g195) & (!g200) & (!g60) & (g61)) + ((!g185) & (g190) & (g195) & (!g200) & (g60) & (!g61)) + ((!g185) & (g190) & (g195) & (g200) & (!g60) & (g61)) + ((!g185) & (g190) & (g195) & (g200) & (g60) & (!g61)) + ((!g185) & (g190) & (g195) & (g200) & (g60) & (g61)) + ((g185) & (!g190) & (!g195) & (!g200) & (!g60) & (!g61)) + ((g185) & (!g190) & (!g195) & (g200) & (!g60) & (!g61)) + ((g185) & (!g190) & (!g195) & (g200) & (g60) & (g61)) + ((g185) & (!g190) & (g195) & (!g200) & (!g60) & (!g61)) + ((g185) & (!g190) & (g195) & (!g200) & (!g60) & (g61)) + ((g185) & (!g190) & (g195) & (g200) & (!g60) & (!g61)) + ((g185) & (!g190) & (g195) & (g200) & (!g60) & (g61)) + ((g185) & (!g190) & (g195) & (g200) & (g60) & (g61)) + ((g185) & (g190) & (!g195) & (!g200) & (!g60) & (!g61)) + ((g185) & (g190) & (!g195) & (!g200) & (g60) & (!g61)) + ((g185) & (g190) & (!g195) & (g200) & (!g60) & (!g61)) + ((g185) & (g190) & (!g195) & (g200) & (g60) & (!g61)) + ((g185) & (g190) & (!g195) & (g200) & (g60) & (g61)) + ((g185) & (g190) & (g195) & (!g200) & (!g60) & (!g61)) + ((g185) & (g190) & (g195) & (!g200) & (!g60) & (g61)) + ((g185) & (g190) & (g195) & (!g200) & (g60) & (!g61)) + ((g185) & (g190) & (g195) & (g200) & (!g60) & (!g61)) + ((g185) & (g190) & (g195) & (g200) & (!g60) & (g61)) + ((g185) & (g190) & (g195) & (g200) & (g60) & (!g61)) + ((g185) & (g190) & (g195) & (g200) & (g60) & (g61)));
	assign g7240 = (((!g832) & (g1033) & (!g202)) + ((!g832) & (g1033) & (g202)) + ((g832) & (!g1033) & (g202)) + ((g832) & (g1033) & (g202)));
	assign g203 = (((!g34) & (!reset) & (!g201) & (g202)) + ((!g34) & (!reset) & (g201) & (g202)) + ((g34) & (!reset) & (g201) & (!g202)) + ((g34) & (!reset) & (g201) & (g202)));
	assign g208 = (((!g204) & (!g205) & (!g206) & (g207) & (g60) & (g61)) + ((!g204) & (!g205) & (g206) & (!g207) & (!g60) & (g61)) + ((!g204) & (!g205) & (g206) & (g207) & (!g60) & (g61)) + ((!g204) & (!g205) & (g206) & (g207) & (g60) & (g61)) + ((!g204) & (g205) & (!g206) & (!g207) & (g60) & (!g61)) + ((!g204) & (g205) & (!g206) & (g207) & (g60) & (!g61)) + ((!g204) & (g205) & (!g206) & (g207) & (g60) & (g61)) + ((!g204) & (g205) & (g206) & (!g207) & (!g60) & (g61)) + ((!g204) & (g205) & (g206) & (!g207) & (g60) & (!g61)) + ((!g204) & (g205) & (g206) & (g207) & (!g60) & (g61)) + ((!g204) & (g205) & (g206) & (g207) & (g60) & (!g61)) + ((!g204) & (g205) & (g206) & (g207) & (g60) & (g61)) + ((g204) & (!g205) & (!g206) & (!g207) & (!g60) & (!g61)) + ((g204) & (!g205) & (!g206) & (g207) & (!g60) & (!g61)) + ((g204) & (!g205) & (!g206) & (g207) & (g60) & (g61)) + ((g204) & (!g205) & (g206) & (!g207) & (!g60) & (!g61)) + ((g204) & (!g205) & (g206) & (!g207) & (!g60) & (g61)) + ((g204) & (!g205) & (g206) & (g207) & (!g60) & (!g61)) + ((g204) & (!g205) & (g206) & (g207) & (!g60) & (g61)) + ((g204) & (!g205) & (g206) & (g207) & (g60) & (g61)) + ((g204) & (g205) & (!g206) & (!g207) & (!g60) & (!g61)) + ((g204) & (g205) & (!g206) & (!g207) & (g60) & (!g61)) + ((g204) & (g205) & (!g206) & (g207) & (!g60) & (!g61)) + ((g204) & (g205) & (!g206) & (g207) & (g60) & (!g61)) + ((g204) & (g205) & (!g206) & (g207) & (g60) & (g61)) + ((g204) & (g205) & (g206) & (!g207) & (!g60) & (!g61)) + ((g204) & (g205) & (g206) & (!g207) & (!g60) & (g61)) + ((g204) & (g205) & (g206) & (!g207) & (g60) & (!g61)) + ((g204) & (g205) & (g206) & (g207) & (!g60) & (!g61)) + ((g204) & (g205) & (g206) & (g207) & (!g60) & (g61)) + ((g204) & (g205) & (g206) & (g207) & (g60) & (!g61)) + ((g204) & (g205) & (g206) & (g207) & (g60) & (g61)));
	assign g213 = (((!g209) & (!g210) & (!g211) & (g212) & (g60) & (g61)) + ((!g209) & (!g210) & (g211) & (!g212) & (!g60) & (g61)) + ((!g209) & (!g210) & (g211) & (g212) & (!g60) & (g61)) + ((!g209) & (!g210) & (g211) & (g212) & (g60) & (g61)) + ((!g209) & (g210) & (!g211) & (!g212) & (g60) & (!g61)) + ((!g209) & (g210) & (!g211) & (g212) & (g60) & (!g61)) + ((!g209) & (g210) & (!g211) & (g212) & (g60) & (g61)) + ((!g209) & (g210) & (g211) & (!g212) & (!g60) & (g61)) + ((!g209) & (g210) & (g211) & (!g212) & (g60) & (!g61)) + ((!g209) & (g210) & (g211) & (g212) & (!g60) & (g61)) + ((!g209) & (g210) & (g211) & (g212) & (g60) & (!g61)) + ((!g209) & (g210) & (g211) & (g212) & (g60) & (g61)) + ((g209) & (!g210) & (!g211) & (!g212) & (!g60) & (!g61)) + ((g209) & (!g210) & (!g211) & (g212) & (!g60) & (!g61)) + ((g209) & (!g210) & (!g211) & (g212) & (g60) & (g61)) + ((g209) & (!g210) & (g211) & (!g212) & (!g60) & (!g61)) + ((g209) & (!g210) & (g211) & (!g212) & (!g60) & (g61)) + ((g209) & (!g210) & (g211) & (g212) & (!g60) & (!g61)) + ((g209) & (!g210) & (g211) & (g212) & (!g60) & (g61)) + ((g209) & (!g210) & (g211) & (g212) & (g60) & (g61)) + ((g209) & (g210) & (!g211) & (!g212) & (!g60) & (!g61)) + ((g209) & (g210) & (!g211) & (!g212) & (g60) & (!g61)) + ((g209) & (g210) & (!g211) & (g212) & (!g60) & (!g61)) + ((g209) & (g210) & (!g211) & (g212) & (g60) & (!g61)) + ((g209) & (g210) & (!g211) & (g212) & (g60) & (g61)) + ((g209) & (g210) & (g211) & (!g212) & (!g60) & (!g61)) + ((g209) & (g210) & (g211) & (!g212) & (!g60) & (g61)) + ((g209) & (g210) & (g211) & (!g212) & (g60) & (!g61)) + ((g209) & (g210) & (g211) & (g212) & (!g60) & (!g61)) + ((g209) & (g210) & (g211) & (g212) & (!g60) & (g61)) + ((g209) & (g210) & (g211) & (g212) & (g60) & (!g61)) + ((g209) & (g210) & (g211) & (g212) & (g60) & (g61)));
	assign g218 = (((!g214) & (!g215) & (!g216) & (g217) & (g60) & (g61)) + ((!g214) & (!g215) & (g216) & (!g217) & (!g60) & (g61)) + ((!g214) & (!g215) & (g216) & (g217) & (!g60) & (g61)) + ((!g214) & (!g215) & (g216) & (g217) & (g60) & (g61)) + ((!g214) & (g215) & (!g216) & (!g217) & (g60) & (!g61)) + ((!g214) & (g215) & (!g216) & (g217) & (g60) & (!g61)) + ((!g214) & (g215) & (!g216) & (g217) & (g60) & (g61)) + ((!g214) & (g215) & (g216) & (!g217) & (!g60) & (g61)) + ((!g214) & (g215) & (g216) & (!g217) & (g60) & (!g61)) + ((!g214) & (g215) & (g216) & (g217) & (!g60) & (g61)) + ((!g214) & (g215) & (g216) & (g217) & (g60) & (!g61)) + ((!g214) & (g215) & (g216) & (g217) & (g60) & (g61)) + ((g214) & (!g215) & (!g216) & (!g217) & (!g60) & (!g61)) + ((g214) & (!g215) & (!g216) & (g217) & (!g60) & (!g61)) + ((g214) & (!g215) & (!g216) & (g217) & (g60) & (g61)) + ((g214) & (!g215) & (g216) & (!g217) & (!g60) & (!g61)) + ((g214) & (!g215) & (g216) & (!g217) & (!g60) & (g61)) + ((g214) & (!g215) & (g216) & (g217) & (!g60) & (!g61)) + ((g214) & (!g215) & (g216) & (g217) & (!g60) & (g61)) + ((g214) & (!g215) & (g216) & (g217) & (g60) & (g61)) + ((g214) & (g215) & (!g216) & (!g217) & (!g60) & (!g61)) + ((g214) & (g215) & (!g216) & (!g217) & (g60) & (!g61)) + ((g214) & (g215) & (!g216) & (g217) & (!g60) & (!g61)) + ((g214) & (g215) & (!g216) & (g217) & (g60) & (!g61)) + ((g214) & (g215) & (!g216) & (g217) & (g60) & (g61)) + ((g214) & (g215) & (g216) & (!g217) & (!g60) & (!g61)) + ((g214) & (g215) & (g216) & (!g217) & (!g60) & (g61)) + ((g214) & (g215) & (g216) & (!g217) & (g60) & (!g61)) + ((g214) & (g215) & (g216) & (g217) & (!g60) & (!g61)) + ((g214) & (g215) & (g216) & (g217) & (!g60) & (g61)) + ((g214) & (g215) & (g216) & (g217) & (g60) & (!g61)) + ((g214) & (g215) & (g216) & (g217) & (g60) & (g61)));
	assign g223 = (((!g219) & (!g220) & (!g221) & (g222) & (g60) & (g61)) + ((!g219) & (!g220) & (g221) & (!g222) & (!g60) & (g61)) + ((!g219) & (!g220) & (g221) & (g222) & (!g60) & (g61)) + ((!g219) & (!g220) & (g221) & (g222) & (g60) & (g61)) + ((!g219) & (g220) & (!g221) & (!g222) & (g60) & (!g61)) + ((!g219) & (g220) & (!g221) & (g222) & (g60) & (!g61)) + ((!g219) & (g220) & (!g221) & (g222) & (g60) & (g61)) + ((!g219) & (g220) & (g221) & (!g222) & (!g60) & (g61)) + ((!g219) & (g220) & (g221) & (!g222) & (g60) & (!g61)) + ((!g219) & (g220) & (g221) & (g222) & (!g60) & (g61)) + ((!g219) & (g220) & (g221) & (g222) & (g60) & (!g61)) + ((!g219) & (g220) & (g221) & (g222) & (g60) & (g61)) + ((g219) & (!g220) & (!g221) & (!g222) & (!g60) & (!g61)) + ((g219) & (!g220) & (!g221) & (g222) & (!g60) & (!g61)) + ((g219) & (!g220) & (!g221) & (g222) & (g60) & (g61)) + ((g219) & (!g220) & (g221) & (!g222) & (!g60) & (!g61)) + ((g219) & (!g220) & (g221) & (!g222) & (!g60) & (g61)) + ((g219) & (!g220) & (g221) & (g222) & (!g60) & (!g61)) + ((g219) & (!g220) & (g221) & (g222) & (!g60) & (g61)) + ((g219) & (!g220) & (g221) & (g222) & (g60) & (g61)) + ((g219) & (g220) & (!g221) & (!g222) & (!g60) & (!g61)) + ((g219) & (g220) & (!g221) & (!g222) & (g60) & (!g61)) + ((g219) & (g220) & (!g221) & (g222) & (!g60) & (!g61)) + ((g219) & (g220) & (!g221) & (g222) & (g60) & (!g61)) + ((g219) & (g220) & (!g221) & (g222) & (g60) & (g61)) + ((g219) & (g220) & (g221) & (!g222) & (!g60) & (!g61)) + ((g219) & (g220) & (g221) & (!g222) & (!g60) & (g61)) + ((g219) & (g220) & (g221) & (!g222) & (g60) & (!g61)) + ((g219) & (g220) & (g221) & (g222) & (!g60) & (!g61)) + ((g219) & (g220) & (g221) & (g222) & (!g60) & (g61)) + ((g219) & (g220) & (g221) & (g222) & (g60) & (!g61)) + ((g219) & (g220) & (g221) & (g222) & (g60) & (g61)));
	assign g224 = (((!g208) & (!g213) & (!g218) & (g223) & (g42) & (g43)) + ((!g208) & (!g213) & (g218) & (!g223) & (!g42) & (g43)) + ((!g208) & (!g213) & (g218) & (g223) & (!g42) & (g43)) + ((!g208) & (!g213) & (g218) & (g223) & (g42) & (g43)) + ((!g208) & (g213) & (!g218) & (!g223) & (g42) & (!g43)) + ((!g208) & (g213) & (!g218) & (g223) & (g42) & (!g43)) + ((!g208) & (g213) & (!g218) & (g223) & (g42) & (g43)) + ((!g208) & (g213) & (g218) & (!g223) & (!g42) & (g43)) + ((!g208) & (g213) & (g218) & (!g223) & (g42) & (!g43)) + ((!g208) & (g213) & (g218) & (g223) & (!g42) & (g43)) + ((!g208) & (g213) & (g218) & (g223) & (g42) & (!g43)) + ((!g208) & (g213) & (g218) & (g223) & (g42) & (g43)) + ((g208) & (!g213) & (!g218) & (!g223) & (!g42) & (!g43)) + ((g208) & (!g213) & (!g218) & (g223) & (!g42) & (!g43)) + ((g208) & (!g213) & (!g218) & (g223) & (g42) & (g43)) + ((g208) & (!g213) & (g218) & (!g223) & (!g42) & (!g43)) + ((g208) & (!g213) & (g218) & (!g223) & (!g42) & (g43)) + ((g208) & (!g213) & (g218) & (g223) & (!g42) & (!g43)) + ((g208) & (!g213) & (g218) & (g223) & (!g42) & (g43)) + ((g208) & (!g213) & (g218) & (g223) & (g42) & (g43)) + ((g208) & (g213) & (!g218) & (!g223) & (!g42) & (!g43)) + ((g208) & (g213) & (!g218) & (!g223) & (g42) & (!g43)) + ((g208) & (g213) & (!g218) & (g223) & (!g42) & (!g43)) + ((g208) & (g213) & (!g218) & (g223) & (g42) & (!g43)) + ((g208) & (g213) & (!g218) & (g223) & (g42) & (g43)) + ((g208) & (g213) & (g218) & (!g223) & (!g42) & (!g43)) + ((g208) & (g213) & (g218) & (!g223) & (!g42) & (g43)) + ((g208) & (g213) & (g218) & (!g223) & (g42) & (!g43)) + ((g208) & (g213) & (g218) & (g223) & (!g42) & (!g43)) + ((g208) & (g213) & (g218) & (g223) & (!g42) & (g43)) + ((g208) & (g213) & (g218) & (g223) & (g42) & (!g43)) + ((g208) & (g213) & (g218) & (g223) & (g42) & (g43)));
	assign g7241 = (((!g832) & (g1066) & (!g225)) + ((!g832) & (g1066) & (g225)) + ((g832) & (!g1066) & (g225)) + ((g832) & (g1066) & (g225)));
	assign g226 = (((!g34) & (!reset) & (!g224) & (g225)) + ((!g34) & (!reset) & (g224) & (g225)) + ((g34) & (!reset) & (g224) & (!g225)) + ((g34) & (!reset) & (g224) & (g225)));
	assign g231 = (((!g227) & (!g228) & (!g229) & (g230) & (g42) & (g43)) + ((!g227) & (!g228) & (g229) & (!g230) & (!g42) & (g43)) + ((!g227) & (!g228) & (g229) & (g230) & (!g42) & (g43)) + ((!g227) & (!g228) & (g229) & (g230) & (g42) & (g43)) + ((!g227) & (g228) & (!g229) & (!g230) & (g42) & (!g43)) + ((!g227) & (g228) & (!g229) & (g230) & (g42) & (!g43)) + ((!g227) & (g228) & (!g229) & (g230) & (g42) & (g43)) + ((!g227) & (g228) & (g229) & (!g230) & (!g42) & (g43)) + ((!g227) & (g228) & (g229) & (!g230) & (g42) & (!g43)) + ((!g227) & (g228) & (g229) & (g230) & (!g42) & (g43)) + ((!g227) & (g228) & (g229) & (g230) & (g42) & (!g43)) + ((!g227) & (g228) & (g229) & (g230) & (g42) & (g43)) + ((g227) & (!g228) & (!g229) & (!g230) & (!g42) & (!g43)) + ((g227) & (!g228) & (!g229) & (g230) & (!g42) & (!g43)) + ((g227) & (!g228) & (!g229) & (g230) & (g42) & (g43)) + ((g227) & (!g228) & (g229) & (!g230) & (!g42) & (!g43)) + ((g227) & (!g228) & (g229) & (!g230) & (!g42) & (g43)) + ((g227) & (!g228) & (g229) & (g230) & (!g42) & (!g43)) + ((g227) & (!g228) & (g229) & (g230) & (!g42) & (g43)) + ((g227) & (!g228) & (g229) & (g230) & (g42) & (g43)) + ((g227) & (g228) & (!g229) & (!g230) & (!g42) & (!g43)) + ((g227) & (g228) & (!g229) & (!g230) & (g42) & (!g43)) + ((g227) & (g228) & (!g229) & (g230) & (!g42) & (!g43)) + ((g227) & (g228) & (!g229) & (g230) & (g42) & (!g43)) + ((g227) & (g228) & (!g229) & (g230) & (g42) & (g43)) + ((g227) & (g228) & (g229) & (!g230) & (!g42) & (!g43)) + ((g227) & (g228) & (g229) & (!g230) & (!g42) & (g43)) + ((g227) & (g228) & (g229) & (!g230) & (g42) & (!g43)) + ((g227) & (g228) & (g229) & (g230) & (!g42) & (!g43)) + ((g227) & (g228) & (g229) & (g230) & (!g42) & (g43)) + ((g227) & (g228) & (g229) & (g230) & (g42) & (!g43)) + ((g227) & (g228) & (g229) & (g230) & (g42) & (g43)));
	assign g236 = (((!g232) & (!g233) & (!g234) & (g235) & (g42) & (g43)) + ((!g232) & (!g233) & (g234) & (!g235) & (!g42) & (g43)) + ((!g232) & (!g233) & (g234) & (g235) & (!g42) & (g43)) + ((!g232) & (!g233) & (g234) & (g235) & (g42) & (g43)) + ((!g232) & (g233) & (!g234) & (!g235) & (g42) & (!g43)) + ((!g232) & (g233) & (!g234) & (g235) & (g42) & (!g43)) + ((!g232) & (g233) & (!g234) & (g235) & (g42) & (g43)) + ((!g232) & (g233) & (g234) & (!g235) & (!g42) & (g43)) + ((!g232) & (g233) & (g234) & (!g235) & (g42) & (!g43)) + ((!g232) & (g233) & (g234) & (g235) & (!g42) & (g43)) + ((!g232) & (g233) & (g234) & (g235) & (g42) & (!g43)) + ((!g232) & (g233) & (g234) & (g235) & (g42) & (g43)) + ((g232) & (!g233) & (!g234) & (!g235) & (!g42) & (!g43)) + ((g232) & (!g233) & (!g234) & (g235) & (!g42) & (!g43)) + ((g232) & (!g233) & (!g234) & (g235) & (g42) & (g43)) + ((g232) & (!g233) & (g234) & (!g235) & (!g42) & (!g43)) + ((g232) & (!g233) & (g234) & (!g235) & (!g42) & (g43)) + ((g232) & (!g233) & (g234) & (g235) & (!g42) & (!g43)) + ((g232) & (!g233) & (g234) & (g235) & (!g42) & (g43)) + ((g232) & (!g233) & (g234) & (g235) & (g42) & (g43)) + ((g232) & (g233) & (!g234) & (!g235) & (!g42) & (!g43)) + ((g232) & (g233) & (!g234) & (!g235) & (g42) & (!g43)) + ((g232) & (g233) & (!g234) & (g235) & (!g42) & (!g43)) + ((g232) & (g233) & (!g234) & (g235) & (g42) & (!g43)) + ((g232) & (g233) & (!g234) & (g235) & (g42) & (g43)) + ((g232) & (g233) & (g234) & (!g235) & (!g42) & (!g43)) + ((g232) & (g233) & (g234) & (!g235) & (!g42) & (g43)) + ((g232) & (g233) & (g234) & (!g235) & (g42) & (!g43)) + ((g232) & (g233) & (g234) & (g235) & (!g42) & (!g43)) + ((g232) & (g233) & (g234) & (g235) & (!g42) & (g43)) + ((g232) & (g233) & (g234) & (g235) & (g42) & (!g43)) + ((g232) & (g233) & (g234) & (g235) & (g42) & (g43)));
	assign g241 = (((!g237) & (!g238) & (!g239) & (g240) & (g42) & (g43)) + ((!g237) & (!g238) & (g239) & (!g240) & (!g42) & (g43)) + ((!g237) & (!g238) & (g239) & (g240) & (!g42) & (g43)) + ((!g237) & (!g238) & (g239) & (g240) & (g42) & (g43)) + ((!g237) & (g238) & (!g239) & (!g240) & (g42) & (!g43)) + ((!g237) & (g238) & (!g239) & (g240) & (g42) & (!g43)) + ((!g237) & (g238) & (!g239) & (g240) & (g42) & (g43)) + ((!g237) & (g238) & (g239) & (!g240) & (!g42) & (g43)) + ((!g237) & (g238) & (g239) & (!g240) & (g42) & (!g43)) + ((!g237) & (g238) & (g239) & (g240) & (!g42) & (g43)) + ((!g237) & (g238) & (g239) & (g240) & (g42) & (!g43)) + ((!g237) & (g238) & (g239) & (g240) & (g42) & (g43)) + ((g237) & (!g238) & (!g239) & (!g240) & (!g42) & (!g43)) + ((g237) & (!g238) & (!g239) & (g240) & (!g42) & (!g43)) + ((g237) & (!g238) & (!g239) & (g240) & (g42) & (g43)) + ((g237) & (!g238) & (g239) & (!g240) & (!g42) & (!g43)) + ((g237) & (!g238) & (g239) & (!g240) & (!g42) & (g43)) + ((g237) & (!g238) & (g239) & (g240) & (!g42) & (!g43)) + ((g237) & (!g238) & (g239) & (g240) & (!g42) & (g43)) + ((g237) & (!g238) & (g239) & (g240) & (g42) & (g43)) + ((g237) & (g238) & (!g239) & (!g240) & (!g42) & (!g43)) + ((g237) & (g238) & (!g239) & (!g240) & (g42) & (!g43)) + ((g237) & (g238) & (!g239) & (g240) & (!g42) & (!g43)) + ((g237) & (g238) & (!g239) & (g240) & (g42) & (!g43)) + ((g237) & (g238) & (!g239) & (g240) & (g42) & (g43)) + ((g237) & (g238) & (g239) & (!g240) & (!g42) & (!g43)) + ((g237) & (g238) & (g239) & (!g240) & (!g42) & (g43)) + ((g237) & (g238) & (g239) & (!g240) & (g42) & (!g43)) + ((g237) & (g238) & (g239) & (g240) & (!g42) & (!g43)) + ((g237) & (g238) & (g239) & (g240) & (!g42) & (g43)) + ((g237) & (g238) & (g239) & (g240) & (g42) & (!g43)) + ((g237) & (g238) & (g239) & (g240) & (g42) & (g43)));
	assign g246 = (((!g242) & (!g243) & (!g244) & (g245) & (g42) & (g43)) + ((!g242) & (!g243) & (g244) & (!g245) & (!g42) & (g43)) + ((!g242) & (!g243) & (g244) & (g245) & (!g42) & (g43)) + ((!g242) & (!g243) & (g244) & (g245) & (g42) & (g43)) + ((!g242) & (g243) & (!g244) & (!g245) & (g42) & (!g43)) + ((!g242) & (g243) & (!g244) & (g245) & (g42) & (!g43)) + ((!g242) & (g243) & (!g244) & (g245) & (g42) & (g43)) + ((!g242) & (g243) & (g244) & (!g245) & (!g42) & (g43)) + ((!g242) & (g243) & (g244) & (!g245) & (g42) & (!g43)) + ((!g242) & (g243) & (g244) & (g245) & (!g42) & (g43)) + ((!g242) & (g243) & (g244) & (g245) & (g42) & (!g43)) + ((!g242) & (g243) & (g244) & (g245) & (g42) & (g43)) + ((g242) & (!g243) & (!g244) & (!g245) & (!g42) & (!g43)) + ((g242) & (!g243) & (!g244) & (g245) & (!g42) & (!g43)) + ((g242) & (!g243) & (!g244) & (g245) & (g42) & (g43)) + ((g242) & (!g243) & (g244) & (!g245) & (!g42) & (!g43)) + ((g242) & (!g243) & (g244) & (!g245) & (!g42) & (g43)) + ((g242) & (!g243) & (g244) & (g245) & (!g42) & (!g43)) + ((g242) & (!g243) & (g244) & (g245) & (!g42) & (g43)) + ((g242) & (!g243) & (g244) & (g245) & (g42) & (g43)) + ((g242) & (g243) & (!g244) & (!g245) & (!g42) & (!g43)) + ((g242) & (g243) & (!g244) & (!g245) & (g42) & (!g43)) + ((g242) & (g243) & (!g244) & (g245) & (!g42) & (!g43)) + ((g242) & (g243) & (!g244) & (g245) & (g42) & (!g43)) + ((g242) & (g243) & (!g244) & (g245) & (g42) & (g43)) + ((g242) & (g243) & (g244) & (!g245) & (!g42) & (!g43)) + ((g242) & (g243) & (g244) & (!g245) & (!g42) & (g43)) + ((g242) & (g243) & (g244) & (!g245) & (g42) & (!g43)) + ((g242) & (g243) & (g244) & (g245) & (!g42) & (!g43)) + ((g242) & (g243) & (g244) & (g245) & (!g42) & (g43)) + ((g242) & (g243) & (g244) & (g245) & (g42) & (!g43)) + ((g242) & (g243) & (g244) & (g245) & (g42) & (g43)));
	assign g247 = (((!g231) & (!g236) & (!g241) & (g246) & (g60) & (g61)) + ((!g231) & (!g236) & (g241) & (!g246) & (!g60) & (g61)) + ((!g231) & (!g236) & (g241) & (g246) & (!g60) & (g61)) + ((!g231) & (!g236) & (g241) & (g246) & (g60) & (g61)) + ((!g231) & (g236) & (!g241) & (!g246) & (g60) & (!g61)) + ((!g231) & (g236) & (!g241) & (g246) & (g60) & (!g61)) + ((!g231) & (g236) & (!g241) & (g246) & (g60) & (g61)) + ((!g231) & (g236) & (g241) & (!g246) & (!g60) & (g61)) + ((!g231) & (g236) & (g241) & (!g246) & (g60) & (!g61)) + ((!g231) & (g236) & (g241) & (g246) & (!g60) & (g61)) + ((!g231) & (g236) & (g241) & (g246) & (g60) & (!g61)) + ((!g231) & (g236) & (g241) & (g246) & (g60) & (g61)) + ((g231) & (!g236) & (!g241) & (!g246) & (!g60) & (!g61)) + ((g231) & (!g236) & (!g241) & (g246) & (!g60) & (!g61)) + ((g231) & (!g236) & (!g241) & (g246) & (g60) & (g61)) + ((g231) & (!g236) & (g241) & (!g246) & (!g60) & (!g61)) + ((g231) & (!g236) & (g241) & (!g246) & (!g60) & (g61)) + ((g231) & (!g236) & (g241) & (g246) & (!g60) & (!g61)) + ((g231) & (!g236) & (g241) & (g246) & (!g60) & (g61)) + ((g231) & (!g236) & (g241) & (g246) & (g60) & (g61)) + ((g231) & (g236) & (!g241) & (!g246) & (!g60) & (!g61)) + ((g231) & (g236) & (!g241) & (!g246) & (g60) & (!g61)) + ((g231) & (g236) & (!g241) & (g246) & (!g60) & (!g61)) + ((g231) & (g236) & (!g241) & (g246) & (g60) & (!g61)) + ((g231) & (g236) & (!g241) & (g246) & (g60) & (g61)) + ((g231) & (g236) & (g241) & (!g246) & (!g60) & (!g61)) + ((g231) & (g236) & (g241) & (!g246) & (!g60) & (g61)) + ((g231) & (g236) & (g241) & (!g246) & (g60) & (!g61)) + ((g231) & (g236) & (g241) & (g246) & (!g60) & (!g61)) + ((g231) & (g236) & (g241) & (g246) & (!g60) & (g61)) + ((g231) & (g236) & (g241) & (g246) & (g60) & (!g61)) + ((g231) & (g236) & (g241) & (g246) & (g60) & (g61)));
	assign g7242 = (((!g832) & (g1100) & (!g248)) + ((!g832) & (g1100) & (g248)) + ((g832) & (!g1100) & (g248)) + ((g832) & (g1100) & (g248)));
	assign g249 = (((!g34) & (!reset) & (!g247) & (g248)) + ((!g34) & (!reset) & (g247) & (g248)) + ((g34) & (!reset) & (g247) & (!g248)) + ((g34) & (!reset) & (g247) & (g248)));
	assign g254 = (((!g250) & (!g251) & (!g252) & (g253) & (g60) & (g61)) + ((!g250) & (!g251) & (g252) & (!g253) & (!g60) & (g61)) + ((!g250) & (!g251) & (g252) & (g253) & (!g60) & (g61)) + ((!g250) & (!g251) & (g252) & (g253) & (g60) & (g61)) + ((!g250) & (g251) & (!g252) & (!g253) & (g60) & (!g61)) + ((!g250) & (g251) & (!g252) & (g253) & (g60) & (!g61)) + ((!g250) & (g251) & (!g252) & (g253) & (g60) & (g61)) + ((!g250) & (g251) & (g252) & (!g253) & (!g60) & (g61)) + ((!g250) & (g251) & (g252) & (!g253) & (g60) & (!g61)) + ((!g250) & (g251) & (g252) & (g253) & (!g60) & (g61)) + ((!g250) & (g251) & (g252) & (g253) & (g60) & (!g61)) + ((!g250) & (g251) & (g252) & (g253) & (g60) & (g61)) + ((g250) & (!g251) & (!g252) & (!g253) & (!g60) & (!g61)) + ((g250) & (!g251) & (!g252) & (g253) & (!g60) & (!g61)) + ((g250) & (!g251) & (!g252) & (g253) & (g60) & (g61)) + ((g250) & (!g251) & (g252) & (!g253) & (!g60) & (!g61)) + ((g250) & (!g251) & (g252) & (!g253) & (!g60) & (g61)) + ((g250) & (!g251) & (g252) & (g253) & (!g60) & (!g61)) + ((g250) & (!g251) & (g252) & (g253) & (!g60) & (g61)) + ((g250) & (!g251) & (g252) & (g253) & (g60) & (g61)) + ((g250) & (g251) & (!g252) & (!g253) & (!g60) & (!g61)) + ((g250) & (g251) & (!g252) & (!g253) & (g60) & (!g61)) + ((g250) & (g251) & (!g252) & (g253) & (!g60) & (!g61)) + ((g250) & (g251) & (!g252) & (g253) & (g60) & (!g61)) + ((g250) & (g251) & (!g252) & (g253) & (g60) & (g61)) + ((g250) & (g251) & (g252) & (!g253) & (!g60) & (!g61)) + ((g250) & (g251) & (g252) & (!g253) & (!g60) & (g61)) + ((g250) & (g251) & (g252) & (!g253) & (g60) & (!g61)) + ((g250) & (g251) & (g252) & (g253) & (!g60) & (!g61)) + ((g250) & (g251) & (g252) & (g253) & (!g60) & (g61)) + ((g250) & (g251) & (g252) & (g253) & (g60) & (!g61)) + ((g250) & (g251) & (g252) & (g253) & (g60) & (g61)));
	assign g259 = (((!g255) & (!g256) & (!g257) & (g258) & (g60) & (g61)) + ((!g255) & (!g256) & (g257) & (!g258) & (!g60) & (g61)) + ((!g255) & (!g256) & (g257) & (g258) & (!g60) & (g61)) + ((!g255) & (!g256) & (g257) & (g258) & (g60) & (g61)) + ((!g255) & (g256) & (!g257) & (!g258) & (g60) & (!g61)) + ((!g255) & (g256) & (!g257) & (g258) & (g60) & (!g61)) + ((!g255) & (g256) & (!g257) & (g258) & (g60) & (g61)) + ((!g255) & (g256) & (g257) & (!g258) & (!g60) & (g61)) + ((!g255) & (g256) & (g257) & (!g258) & (g60) & (!g61)) + ((!g255) & (g256) & (g257) & (g258) & (!g60) & (g61)) + ((!g255) & (g256) & (g257) & (g258) & (g60) & (!g61)) + ((!g255) & (g256) & (g257) & (g258) & (g60) & (g61)) + ((g255) & (!g256) & (!g257) & (!g258) & (!g60) & (!g61)) + ((g255) & (!g256) & (!g257) & (g258) & (!g60) & (!g61)) + ((g255) & (!g256) & (!g257) & (g258) & (g60) & (g61)) + ((g255) & (!g256) & (g257) & (!g258) & (!g60) & (!g61)) + ((g255) & (!g256) & (g257) & (!g258) & (!g60) & (g61)) + ((g255) & (!g256) & (g257) & (g258) & (!g60) & (!g61)) + ((g255) & (!g256) & (g257) & (g258) & (!g60) & (g61)) + ((g255) & (!g256) & (g257) & (g258) & (g60) & (g61)) + ((g255) & (g256) & (!g257) & (!g258) & (!g60) & (!g61)) + ((g255) & (g256) & (!g257) & (!g258) & (g60) & (!g61)) + ((g255) & (g256) & (!g257) & (g258) & (!g60) & (!g61)) + ((g255) & (g256) & (!g257) & (g258) & (g60) & (!g61)) + ((g255) & (g256) & (!g257) & (g258) & (g60) & (g61)) + ((g255) & (g256) & (g257) & (!g258) & (!g60) & (!g61)) + ((g255) & (g256) & (g257) & (!g258) & (!g60) & (g61)) + ((g255) & (g256) & (g257) & (!g258) & (g60) & (!g61)) + ((g255) & (g256) & (g257) & (g258) & (!g60) & (!g61)) + ((g255) & (g256) & (g257) & (g258) & (!g60) & (g61)) + ((g255) & (g256) & (g257) & (g258) & (g60) & (!g61)) + ((g255) & (g256) & (g257) & (g258) & (g60) & (g61)));
	assign g264 = (((!g260) & (!g261) & (!g262) & (g263) & (g60) & (g61)) + ((!g260) & (!g261) & (g262) & (!g263) & (!g60) & (g61)) + ((!g260) & (!g261) & (g262) & (g263) & (!g60) & (g61)) + ((!g260) & (!g261) & (g262) & (g263) & (g60) & (g61)) + ((!g260) & (g261) & (!g262) & (!g263) & (g60) & (!g61)) + ((!g260) & (g261) & (!g262) & (g263) & (g60) & (!g61)) + ((!g260) & (g261) & (!g262) & (g263) & (g60) & (g61)) + ((!g260) & (g261) & (g262) & (!g263) & (!g60) & (g61)) + ((!g260) & (g261) & (g262) & (!g263) & (g60) & (!g61)) + ((!g260) & (g261) & (g262) & (g263) & (!g60) & (g61)) + ((!g260) & (g261) & (g262) & (g263) & (g60) & (!g61)) + ((!g260) & (g261) & (g262) & (g263) & (g60) & (g61)) + ((g260) & (!g261) & (!g262) & (!g263) & (!g60) & (!g61)) + ((g260) & (!g261) & (!g262) & (g263) & (!g60) & (!g61)) + ((g260) & (!g261) & (!g262) & (g263) & (g60) & (g61)) + ((g260) & (!g261) & (g262) & (!g263) & (!g60) & (!g61)) + ((g260) & (!g261) & (g262) & (!g263) & (!g60) & (g61)) + ((g260) & (!g261) & (g262) & (g263) & (!g60) & (!g61)) + ((g260) & (!g261) & (g262) & (g263) & (!g60) & (g61)) + ((g260) & (!g261) & (g262) & (g263) & (g60) & (g61)) + ((g260) & (g261) & (!g262) & (!g263) & (!g60) & (!g61)) + ((g260) & (g261) & (!g262) & (!g263) & (g60) & (!g61)) + ((g260) & (g261) & (!g262) & (g263) & (!g60) & (!g61)) + ((g260) & (g261) & (!g262) & (g263) & (g60) & (!g61)) + ((g260) & (g261) & (!g262) & (g263) & (g60) & (g61)) + ((g260) & (g261) & (g262) & (!g263) & (!g60) & (!g61)) + ((g260) & (g261) & (g262) & (!g263) & (!g60) & (g61)) + ((g260) & (g261) & (g262) & (!g263) & (g60) & (!g61)) + ((g260) & (g261) & (g262) & (g263) & (!g60) & (!g61)) + ((g260) & (g261) & (g262) & (g263) & (!g60) & (g61)) + ((g260) & (g261) & (g262) & (g263) & (g60) & (!g61)) + ((g260) & (g261) & (g262) & (g263) & (g60) & (g61)));
	assign g269 = (((!g265) & (!g266) & (!g267) & (g268) & (g60) & (g61)) + ((!g265) & (!g266) & (g267) & (!g268) & (!g60) & (g61)) + ((!g265) & (!g266) & (g267) & (g268) & (!g60) & (g61)) + ((!g265) & (!g266) & (g267) & (g268) & (g60) & (g61)) + ((!g265) & (g266) & (!g267) & (!g268) & (g60) & (!g61)) + ((!g265) & (g266) & (!g267) & (g268) & (g60) & (!g61)) + ((!g265) & (g266) & (!g267) & (g268) & (g60) & (g61)) + ((!g265) & (g266) & (g267) & (!g268) & (!g60) & (g61)) + ((!g265) & (g266) & (g267) & (!g268) & (g60) & (!g61)) + ((!g265) & (g266) & (g267) & (g268) & (!g60) & (g61)) + ((!g265) & (g266) & (g267) & (g268) & (g60) & (!g61)) + ((!g265) & (g266) & (g267) & (g268) & (g60) & (g61)) + ((g265) & (!g266) & (!g267) & (!g268) & (!g60) & (!g61)) + ((g265) & (!g266) & (!g267) & (g268) & (!g60) & (!g61)) + ((g265) & (!g266) & (!g267) & (g268) & (g60) & (g61)) + ((g265) & (!g266) & (g267) & (!g268) & (!g60) & (!g61)) + ((g265) & (!g266) & (g267) & (!g268) & (!g60) & (g61)) + ((g265) & (!g266) & (g267) & (g268) & (!g60) & (!g61)) + ((g265) & (!g266) & (g267) & (g268) & (!g60) & (g61)) + ((g265) & (!g266) & (g267) & (g268) & (g60) & (g61)) + ((g265) & (g266) & (!g267) & (!g268) & (!g60) & (!g61)) + ((g265) & (g266) & (!g267) & (!g268) & (g60) & (!g61)) + ((g265) & (g266) & (!g267) & (g268) & (!g60) & (!g61)) + ((g265) & (g266) & (!g267) & (g268) & (g60) & (!g61)) + ((g265) & (g266) & (!g267) & (g268) & (g60) & (g61)) + ((g265) & (g266) & (g267) & (!g268) & (!g60) & (!g61)) + ((g265) & (g266) & (g267) & (!g268) & (!g60) & (g61)) + ((g265) & (g266) & (g267) & (!g268) & (g60) & (!g61)) + ((g265) & (g266) & (g267) & (g268) & (!g60) & (!g61)) + ((g265) & (g266) & (g267) & (g268) & (!g60) & (g61)) + ((g265) & (g266) & (g267) & (g268) & (g60) & (!g61)) + ((g265) & (g266) & (g267) & (g268) & (g60) & (g61)));
	assign g270 = (((!g254) & (!g259) & (!g264) & (g269) & (g42) & (g43)) + ((!g254) & (!g259) & (g264) & (!g269) & (!g42) & (g43)) + ((!g254) & (!g259) & (g264) & (g269) & (!g42) & (g43)) + ((!g254) & (!g259) & (g264) & (g269) & (g42) & (g43)) + ((!g254) & (g259) & (!g264) & (!g269) & (g42) & (!g43)) + ((!g254) & (g259) & (!g264) & (g269) & (g42) & (!g43)) + ((!g254) & (g259) & (!g264) & (g269) & (g42) & (g43)) + ((!g254) & (g259) & (g264) & (!g269) & (!g42) & (g43)) + ((!g254) & (g259) & (g264) & (!g269) & (g42) & (!g43)) + ((!g254) & (g259) & (g264) & (g269) & (!g42) & (g43)) + ((!g254) & (g259) & (g264) & (g269) & (g42) & (!g43)) + ((!g254) & (g259) & (g264) & (g269) & (g42) & (g43)) + ((g254) & (!g259) & (!g264) & (!g269) & (!g42) & (!g43)) + ((g254) & (!g259) & (!g264) & (g269) & (!g42) & (!g43)) + ((g254) & (!g259) & (!g264) & (g269) & (g42) & (g43)) + ((g254) & (!g259) & (g264) & (!g269) & (!g42) & (!g43)) + ((g254) & (!g259) & (g264) & (!g269) & (!g42) & (g43)) + ((g254) & (!g259) & (g264) & (g269) & (!g42) & (!g43)) + ((g254) & (!g259) & (g264) & (g269) & (!g42) & (g43)) + ((g254) & (!g259) & (g264) & (g269) & (g42) & (g43)) + ((g254) & (g259) & (!g264) & (!g269) & (!g42) & (!g43)) + ((g254) & (g259) & (!g264) & (!g269) & (g42) & (!g43)) + ((g254) & (g259) & (!g264) & (g269) & (!g42) & (!g43)) + ((g254) & (g259) & (!g264) & (g269) & (g42) & (!g43)) + ((g254) & (g259) & (!g264) & (g269) & (g42) & (g43)) + ((g254) & (g259) & (g264) & (!g269) & (!g42) & (!g43)) + ((g254) & (g259) & (g264) & (!g269) & (!g42) & (g43)) + ((g254) & (g259) & (g264) & (!g269) & (g42) & (!g43)) + ((g254) & (g259) & (g264) & (g269) & (!g42) & (!g43)) + ((g254) & (g259) & (g264) & (g269) & (!g42) & (g43)) + ((g254) & (g259) & (g264) & (g269) & (g42) & (!g43)) + ((g254) & (g259) & (g264) & (g269) & (g42) & (g43)));
	assign g7243 = (((!g832) & (g1133) & (!g271)) + ((!g832) & (g1133) & (g271)) + ((g832) & (!g1133) & (g271)) + ((g832) & (g1133) & (g271)));
	assign g272 = (((!g34) & (!reset) & (!g270) & (g271)) + ((!g34) & (!reset) & (g270) & (g271)) + ((g34) & (!reset) & (g270) & (!g271)) + ((g34) & (!reset) & (g270) & (g271)));
	assign g277 = (((!g273) & (!g274) & (!g275) & (g276) & (g42) & (g43)) + ((!g273) & (!g274) & (g275) & (!g276) & (!g42) & (g43)) + ((!g273) & (!g274) & (g275) & (g276) & (!g42) & (g43)) + ((!g273) & (!g274) & (g275) & (g276) & (g42) & (g43)) + ((!g273) & (g274) & (!g275) & (!g276) & (g42) & (!g43)) + ((!g273) & (g274) & (!g275) & (g276) & (g42) & (!g43)) + ((!g273) & (g274) & (!g275) & (g276) & (g42) & (g43)) + ((!g273) & (g274) & (g275) & (!g276) & (!g42) & (g43)) + ((!g273) & (g274) & (g275) & (!g276) & (g42) & (!g43)) + ((!g273) & (g274) & (g275) & (g276) & (!g42) & (g43)) + ((!g273) & (g274) & (g275) & (g276) & (g42) & (!g43)) + ((!g273) & (g274) & (g275) & (g276) & (g42) & (g43)) + ((g273) & (!g274) & (!g275) & (!g276) & (!g42) & (!g43)) + ((g273) & (!g274) & (!g275) & (g276) & (!g42) & (!g43)) + ((g273) & (!g274) & (!g275) & (g276) & (g42) & (g43)) + ((g273) & (!g274) & (g275) & (!g276) & (!g42) & (!g43)) + ((g273) & (!g274) & (g275) & (!g276) & (!g42) & (g43)) + ((g273) & (!g274) & (g275) & (g276) & (!g42) & (!g43)) + ((g273) & (!g274) & (g275) & (g276) & (!g42) & (g43)) + ((g273) & (!g274) & (g275) & (g276) & (g42) & (g43)) + ((g273) & (g274) & (!g275) & (!g276) & (!g42) & (!g43)) + ((g273) & (g274) & (!g275) & (!g276) & (g42) & (!g43)) + ((g273) & (g274) & (!g275) & (g276) & (!g42) & (!g43)) + ((g273) & (g274) & (!g275) & (g276) & (g42) & (!g43)) + ((g273) & (g274) & (!g275) & (g276) & (g42) & (g43)) + ((g273) & (g274) & (g275) & (!g276) & (!g42) & (!g43)) + ((g273) & (g274) & (g275) & (!g276) & (!g42) & (g43)) + ((g273) & (g274) & (g275) & (!g276) & (g42) & (!g43)) + ((g273) & (g274) & (g275) & (g276) & (!g42) & (!g43)) + ((g273) & (g274) & (g275) & (g276) & (!g42) & (g43)) + ((g273) & (g274) & (g275) & (g276) & (g42) & (!g43)) + ((g273) & (g274) & (g275) & (g276) & (g42) & (g43)));
	assign g282 = (((!g278) & (!g279) & (!g280) & (g281) & (g42) & (g43)) + ((!g278) & (!g279) & (g280) & (!g281) & (!g42) & (g43)) + ((!g278) & (!g279) & (g280) & (g281) & (!g42) & (g43)) + ((!g278) & (!g279) & (g280) & (g281) & (g42) & (g43)) + ((!g278) & (g279) & (!g280) & (!g281) & (g42) & (!g43)) + ((!g278) & (g279) & (!g280) & (g281) & (g42) & (!g43)) + ((!g278) & (g279) & (!g280) & (g281) & (g42) & (g43)) + ((!g278) & (g279) & (g280) & (!g281) & (!g42) & (g43)) + ((!g278) & (g279) & (g280) & (!g281) & (g42) & (!g43)) + ((!g278) & (g279) & (g280) & (g281) & (!g42) & (g43)) + ((!g278) & (g279) & (g280) & (g281) & (g42) & (!g43)) + ((!g278) & (g279) & (g280) & (g281) & (g42) & (g43)) + ((g278) & (!g279) & (!g280) & (!g281) & (!g42) & (!g43)) + ((g278) & (!g279) & (!g280) & (g281) & (!g42) & (!g43)) + ((g278) & (!g279) & (!g280) & (g281) & (g42) & (g43)) + ((g278) & (!g279) & (g280) & (!g281) & (!g42) & (!g43)) + ((g278) & (!g279) & (g280) & (!g281) & (!g42) & (g43)) + ((g278) & (!g279) & (g280) & (g281) & (!g42) & (!g43)) + ((g278) & (!g279) & (g280) & (g281) & (!g42) & (g43)) + ((g278) & (!g279) & (g280) & (g281) & (g42) & (g43)) + ((g278) & (g279) & (!g280) & (!g281) & (!g42) & (!g43)) + ((g278) & (g279) & (!g280) & (!g281) & (g42) & (!g43)) + ((g278) & (g279) & (!g280) & (g281) & (!g42) & (!g43)) + ((g278) & (g279) & (!g280) & (g281) & (g42) & (!g43)) + ((g278) & (g279) & (!g280) & (g281) & (g42) & (g43)) + ((g278) & (g279) & (g280) & (!g281) & (!g42) & (!g43)) + ((g278) & (g279) & (g280) & (!g281) & (!g42) & (g43)) + ((g278) & (g279) & (g280) & (!g281) & (g42) & (!g43)) + ((g278) & (g279) & (g280) & (g281) & (!g42) & (!g43)) + ((g278) & (g279) & (g280) & (g281) & (!g42) & (g43)) + ((g278) & (g279) & (g280) & (g281) & (g42) & (!g43)) + ((g278) & (g279) & (g280) & (g281) & (g42) & (g43)));
	assign g287 = (((!g283) & (!g284) & (!g285) & (g286) & (g42) & (g43)) + ((!g283) & (!g284) & (g285) & (!g286) & (!g42) & (g43)) + ((!g283) & (!g284) & (g285) & (g286) & (!g42) & (g43)) + ((!g283) & (!g284) & (g285) & (g286) & (g42) & (g43)) + ((!g283) & (g284) & (!g285) & (!g286) & (g42) & (!g43)) + ((!g283) & (g284) & (!g285) & (g286) & (g42) & (!g43)) + ((!g283) & (g284) & (!g285) & (g286) & (g42) & (g43)) + ((!g283) & (g284) & (g285) & (!g286) & (!g42) & (g43)) + ((!g283) & (g284) & (g285) & (!g286) & (g42) & (!g43)) + ((!g283) & (g284) & (g285) & (g286) & (!g42) & (g43)) + ((!g283) & (g284) & (g285) & (g286) & (g42) & (!g43)) + ((!g283) & (g284) & (g285) & (g286) & (g42) & (g43)) + ((g283) & (!g284) & (!g285) & (!g286) & (!g42) & (!g43)) + ((g283) & (!g284) & (!g285) & (g286) & (!g42) & (!g43)) + ((g283) & (!g284) & (!g285) & (g286) & (g42) & (g43)) + ((g283) & (!g284) & (g285) & (!g286) & (!g42) & (!g43)) + ((g283) & (!g284) & (g285) & (!g286) & (!g42) & (g43)) + ((g283) & (!g284) & (g285) & (g286) & (!g42) & (!g43)) + ((g283) & (!g284) & (g285) & (g286) & (!g42) & (g43)) + ((g283) & (!g284) & (g285) & (g286) & (g42) & (g43)) + ((g283) & (g284) & (!g285) & (!g286) & (!g42) & (!g43)) + ((g283) & (g284) & (!g285) & (!g286) & (g42) & (!g43)) + ((g283) & (g284) & (!g285) & (g286) & (!g42) & (!g43)) + ((g283) & (g284) & (!g285) & (g286) & (g42) & (!g43)) + ((g283) & (g284) & (!g285) & (g286) & (g42) & (g43)) + ((g283) & (g284) & (g285) & (!g286) & (!g42) & (!g43)) + ((g283) & (g284) & (g285) & (!g286) & (!g42) & (g43)) + ((g283) & (g284) & (g285) & (!g286) & (g42) & (!g43)) + ((g283) & (g284) & (g285) & (g286) & (!g42) & (!g43)) + ((g283) & (g284) & (g285) & (g286) & (!g42) & (g43)) + ((g283) & (g284) & (g285) & (g286) & (g42) & (!g43)) + ((g283) & (g284) & (g285) & (g286) & (g42) & (g43)));
	assign g292 = (((!g288) & (!g289) & (!g290) & (g291) & (g42) & (g43)) + ((!g288) & (!g289) & (g290) & (!g291) & (!g42) & (g43)) + ((!g288) & (!g289) & (g290) & (g291) & (!g42) & (g43)) + ((!g288) & (!g289) & (g290) & (g291) & (g42) & (g43)) + ((!g288) & (g289) & (!g290) & (!g291) & (g42) & (!g43)) + ((!g288) & (g289) & (!g290) & (g291) & (g42) & (!g43)) + ((!g288) & (g289) & (!g290) & (g291) & (g42) & (g43)) + ((!g288) & (g289) & (g290) & (!g291) & (!g42) & (g43)) + ((!g288) & (g289) & (g290) & (!g291) & (g42) & (!g43)) + ((!g288) & (g289) & (g290) & (g291) & (!g42) & (g43)) + ((!g288) & (g289) & (g290) & (g291) & (g42) & (!g43)) + ((!g288) & (g289) & (g290) & (g291) & (g42) & (g43)) + ((g288) & (!g289) & (!g290) & (!g291) & (!g42) & (!g43)) + ((g288) & (!g289) & (!g290) & (g291) & (!g42) & (!g43)) + ((g288) & (!g289) & (!g290) & (g291) & (g42) & (g43)) + ((g288) & (!g289) & (g290) & (!g291) & (!g42) & (!g43)) + ((g288) & (!g289) & (g290) & (!g291) & (!g42) & (g43)) + ((g288) & (!g289) & (g290) & (g291) & (!g42) & (!g43)) + ((g288) & (!g289) & (g290) & (g291) & (!g42) & (g43)) + ((g288) & (!g289) & (g290) & (g291) & (g42) & (g43)) + ((g288) & (g289) & (!g290) & (!g291) & (!g42) & (!g43)) + ((g288) & (g289) & (!g290) & (!g291) & (g42) & (!g43)) + ((g288) & (g289) & (!g290) & (g291) & (!g42) & (!g43)) + ((g288) & (g289) & (!g290) & (g291) & (g42) & (!g43)) + ((g288) & (g289) & (!g290) & (g291) & (g42) & (g43)) + ((g288) & (g289) & (g290) & (!g291) & (!g42) & (!g43)) + ((g288) & (g289) & (g290) & (!g291) & (!g42) & (g43)) + ((g288) & (g289) & (g290) & (!g291) & (g42) & (!g43)) + ((g288) & (g289) & (g290) & (g291) & (!g42) & (!g43)) + ((g288) & (g289) & (g290) & (g291) & (!g42) & (g43)) + ((g288) & (g289) & (g290) & (g291) & (g42) & (!g43)) + ((g288) & (g289) & (g290) & (g291) & (g42) & (g43)));
	assign g293 = (((!g277) & (!g282) & (!g287) & (g292) & (g60) & (g61)) + ((!g277) & (!g282) & (g287) & (!g292) & (!g60) & (g61)) + ((!g277) & (!g282) & (g287) & (g292) & (!g60) & (g61)) + ((!g277) & (!g282) & (g287) & (g292) & (g60) & (g61)) + ((!g277) & (g282) & (!g287) & (!g292) & (g60) & (!g61)) + ((!g277) & (g282) & (!g287) & (g292) & (g60) & (!g61)) + ((!g277) & (g282) & (!g287) & (g292) & (g60) & (g61)) + ((!g277) & (g282) & (g287) & (!g292) & (!g60) & (g61)) + ((!g277) & (g282) & (g287) & (!g292) & (g60) & (!g61)) + ((!g277) & (g282) & (g287) & (g292) & (!g60) & (g61)) + ((!g277) & (g282) & (g287) & (g292) & (g60) & (!g61)) + ((!g277) & (g282) & (g287) & (g292) & (g60) & (g61)) + ((g277) & (!g282) & (!g287) & (!g292) & (!g60) & (!g61)) + ((g277) & (!g282) & (!g287) & (g292) & (!g60) & (!g61)) + ((g277) & (!g282) & (!g287) & (g292) & (g60) & (g61)) + ((g277) & (!g282) & (g287) & (!g292) & (!g60) & (!g61)) + ((g277) & (!g282) & (g287) & (!g292) & (!g60) & (g61)) + ((g277) & (!g282) & (g287) & (g292) & (!g60) & (!g61)) + ((g277) & (!g282) & (g287) & (g292) & (!g60) & (g61)) + ((g277) & (!g282) & (g287) & (g292) & (g60) & (g61)) + ((g277) & (g282) & (!g287) & (!g292) & (!g60) & (!g61)) + ((g277) & (g282) & (!g287) & (!g292) & (g60) & (!g61)) + ((g277) & (g282) & (!g287) & (g292) & (!g60) & (!g61)) + ((g277) & (g282) & (!g287) & (g292) & (g60) & (!g61)) + ((g277) & (g282) & (!g287) & (g292) & (g60) & (g61)) + ((g277) & (g282) & (g287) & (!g292) & (!g60) & (!g61)) + ((g277) & (g282) & (g287) & (!g292) & (!g60) & (g61)) + ((g277) & (g282) & (g287) & (!g292) & (g60) & (!g61)) + ((g277) & (g282) & (g287) & (g292) & (!g60) & (!g61)) + ((g277) & (g282) & (g287) & (g292) & (!g60) & (g61)) + ((g277) & (g282) & (g287) & (g292) & (g60) & (!g61)) + ((g277) & (g282) & (g287) & (g292) & (g60) & (g61)));
	assign g7244 = (((!g832) & (g1167) & (!g294)) + ((!g832) & (g1167) & (g294)) + ((g832) & (!g1167) & (g294)) + ((g832) & (g1167) & (g294)));
	assign g295 = (((!g34) & (!reset) & (!g293) & (g294)) + ((!g34) & (!reset) & (g293) & (g294)) + ((g34) & (!reset) & (g293) & (!g294)) + ((g34) & (!reset) & (g293) & (g294)));
	assign g300 = (((!g296) & (!g297) & (!g298) & (g299) & (g60) & (g61)) + ((!g296) & (!g297) & (g298) & (!g299) & (!g60) & (g61)) + ((!g296) & (!g297) & (g298) & (g299) & (!g60) & (g61)) + ((!g296) & (!g297) & (g298) & (g299) & (g60) & (g61)) + ((!g296) & (g297) & (!g298) & (!g299) & (g60) & (!g61)) + ((!g296) & (g297) & (!g298) & (g299) & (g60) & (!g61)) + ((!g296) & (g297) & (!g298) & (g299) & (g60) & (g61)) + ((!g296) & (g297) & (g298) & (!g299) & (!g60) & (g61)) + ((!g296) & (g297) & (g298) & (!g299) & (g60) & (!g61)) + ((!g296) & (g297) & (g298) & (g299) & (!g60) & (g61)) + ((!g296) & (g297) & (g298) & (g299) & (g60) & (!g61)) + ((!g296) & (g297) & (g298) & (g299) & (g60) & (g61)) + ((g296) & (!g297) & (!g298) & (!g299) & (!g60) & (!g61)) + ((g296) & (!g297) & (!g298) & (g299) & (!g60) & (!g61)) + ((g296) & (!g297) & (!g298) & (g299) & (g60) & (g61)) + ((g296) & (!g297) & (g298) & (!g299) & (!g60) & (!g61)) + ((g296) & (!g297) & (g298) & (!g299) & (!g60) & (g61)) + ((g296) & (!g297) & (g298) & (g299) & (!g60) & (!g61)) + ((g296) & (!g297) & (g298) & (g299) & (!g60) & (g61)) + ((g296) & (!g297) & (g298) & (g299) & (g60) & (g61)) + ((g296) & (g297) & (!g298) & (!g299) & (!g60) & (!g61)) + ((g296) & (g297) & (!g298) & (!g299) & (g60) & (!g61)) + ((g296) & (g297) & (!g298) & (g299) & (!g60) & (!g61)) + ((g296) & (g297) & (!g298) & (g299) & (g60) & (!g61)) + ((g296) & (g297) & (!g298) & (g299) & (g60) & (g61)) + ((g296) & (g297) & (g298) & (!g299) & (!g60) & (!g61)) + ((g296) & (g297) & (g298) & (!g299) & (!g60) & (g61)) + ((g296) & (g297) & (g298) & (!g299) & (g60) & (!g61)) + ((g296) & (g297) & (g298) & (g299) & (!g60) & (!g61)) + ((g296) & (g297) & (g298) & (g299) & (!g60) & (g61)) + ((g296) & (g297) & (g298) & (g299) & (g60) & (!g61)) + ((g296) & (g297) & (g298) & (g299) & (g60) & (g61)));
	assign g305 = (((!g301) & (!g302) & (!g303) & (g304) & (g60) & (g61)) + ((!g301) & (!g302) & (g303) & (!g304) & (!g60) & (g61)) + ((!g301) & (!g302) & (g303) & (g304) & (!g60) & (g61)) + ((!g301) & (!g302) & (g303) & (g304) & (g60) & (g61)) + ((!g301) & (g302) & (!g303) & (!g304) & (g60) & (!g61)) + ((!g301) & (g302) & (!g303) & (g304) & (g60) & (!g61)) + ((!g301) & (g302) & (!g303) & (g304) & (g60) & (g61)) + ((!g301) & (g302) & (g303) & (!g304) & (!g60) & (g61)) + ((!g301) & (g302) & (g303) & (!g304) & (g60) & (!g61)) + ((!g301) & (g302) & (g303) & (g304) & (!g60) & (g61)) + ((!g301) & (g302) & (g303) & (g304) & (g60) & (!g61)) + ((!g301) & (g302) & (g303) & (g304) & (g60) & (g61)) + ((g301) & (!g302) & (!g303) & (!g304) & (!g60) & (!g61)) + ((g301) & (!g302) & (!g303) & (g304) & (!g60) & (!g61)) + ((g301) & (!g302) & (!g303) & (g304) & (g60) & (g61)) + ((g301) & (!g302) & (g303) & (!g304) & (!g60) & (!g61)) + ((g301) & (!g302) & (g303) & (!g304) & (!g60) & (g61)) + ((g301) & (!g302) & (g303) & (g304) & (!g60) & (!g61)) + ((g301) & (!g302) & (g303) & (g304) & (!g60) & (g61)) + ((g301) & (!g302) & (g303) & (g304) & (g60) & (g61)) + ((g301) & (g302) & (!g303) & (!g304) & (!g60) & (!g61)) + ((g301) & (g302) & (!g303) & (!g304) & (g60) & (!g61)) + ((g301) & (g302) & (!g303) & (g304) & (!g60) & (!g61)) + ((g301) & (g302) & (!g303) & (g304) & (g60) & (!g61)) + ((g301) & (g302) & (!g303) & (g304) & (g60) & (g61)) + ((g301) & (g302) & (g303) & (!g304) & (!g60) & (!g61)) + ((g301) & (g302) & (g303) & (!g304) & (!g60) & (g61)) + ((g301) & (g302) & (g303) & (!g304) & (g60) & (!g61)) + ((g301) & (g302) & (g303) & (g304) & (!g60) & (!g61)) + ((g301) & (g302) & (g303) & (g304) & (!g60) & (g61)) + ((g301) & (g302) & (g303) & (g304) & (g60) & (!g61)) + ((g301) & (g302) & (g303) & (g304) & (g60) & (g61)));
	assign g310 = (((!g306) & (!g307) & (!g308) & (g309) & (g60) & (g61)) + ((!g306) & (!g307) & (g308) & (!g309) & (!g60) & (g61)) + ((!g306) & (!g307) & (g308) & (g309) & (!g60) & (g61)) + ((!g306) & (!g307) & (g308) & (g309) & (g60) & (g61)) + ((!g306) & (g307) & (!g308) & (!g309) & (g60) & (!g61)) + ((!g306) & (g307) & (!g308) & (g309) & (g60) & (!g61)) + ((!g306) & (g307) & (!g308) & (g309) & (g60) & (g61)) + ((!g306) & (g307) & (g308) & (!g309) & (!g60) & (g61)) + ((!g306) & (g307) & (g308) & (!g309) & (g60) & (!g61)) + ((!g306) & (g307) & (g308) & (g309) & (!g60) & (g61)) + ((!g306) & (g307) & (g308) & (g309) & (g60) & (!g61)) + ((!g306) & (g307) & (g308) & (g309) & (g60) & (g61)) + ((g306) & (!g307) & (!g308) & (!g309) & (!g60) & (!g61)) + ((g306) & (!g307) & (!g308) & (g309) & (!g60) & (!g61)) + ((g306) & (!g307) & (!g308) & (g309) & (g60) & (g61)) + ((g306) & (!g307) & (g308) & (!g309) & (!g60) & (!g61)) + ((g306) & (!g307) & (g308) & (!g309) & (!g60) & (g61)) + ((g306) & (!g307) & (g308) & (g309) & (!g60) & (!g61)) + ((g306) & (!g307) & (g308) & (g309) & (!g60) & (g61)) + ((g306) & (!g307) & (g308) & (g309) & (g60) & (g61)) + ((g306) & (g307) & (!g308) & (!g309) & (!g60) & (!g61)) + ((g306) & (g307) & (!g308) & (!g309) & (g60) & (!g61)) + ((g306) & (g307) & (!g308) & (g309) & (!g60) & (!g61)) + ((g306) & (g307) & (!g308) & (g309) & (g60) & (!g61)) + ((g306) & (g307) & (!g308) & (g309) & (g60) & (g61)) + ((g306) & (g307) & (g308) & (!g309) & (!g60) & (!g61)) + ((g306) & (g307) & (g308) & (!g309) & (!g60) & (g61)) + ((g306) & (g307) & (g308) & (!g309) & (g60) & (!g61)) + ((g306) & (g307) & (g308) & (g309) & (!g60) & (!g61)) + ((g306) & (g307) & (g308) & (g309) & (!g60) & (g61)) + ((g306) & (g307) & (g308) & (g309) & (g60) & (!g61)) + ((g306) & (g307) & (g308) & (g309) & (g60) & (g61)));
	assign g315 = (((!g311) & (!g312) & (!g313) & (g314) & (g60) & (g61)) + ((!g311) & (!g312) & (g313) & (!g314) & (!g60) & (g61)) + ((!g311) & (!g312) & (g313) & (g314) & (!g60) & (g61)) + ((!g311) & (!g312) & (g313) & (g314) & (g60) & (g61)) + ((!g311) & (g312) & (!g313) & (!g314) & (g60) & (!g61)) + ((!g311) & (g312) & (!g313) & (g314) & (g60) & (!g61)) + ((!g311) & (g312) & (!g313) & (g314) & (g60) & (g61)) + ((!g311) & (g312) & (g313) & (!g314) & (!g60) & (g61)) + ((!g311) & (g312) & (g313) & (!g314) & (g60) & (!g61)) + ((!g311) & (g312) & (g313) & (g314) & (!g60) & (g61)) + ((!g311) & (g312) & (g313) & (g314) & (g60) & (!g61)) + ((!g311) & (g312) & (g313) & (g314) & (g60) & (g61)) + ((g311) & (!g312) & (!g313) & (!g314) & (!g60) & (!g61)) + ((g311) & (!g312) & (!g313) & (g314) & (!g60) & (!g61)) + ((g311) & (!g312) & (!g313) & (g314) & (g60) & (g61)) + ((g311) & (!g312) & (g313) & (!g314) & (!g60) & (!g61)) + ((g311) & (!g312) & (g313) & (!g314) & (!g60) & (g61)) + ((g311) & (!g312) & (g313) & (g314) & (!g60) & (!g61)) + ((g311) & (!g312) & (g313) & (g314) & (!g60) & (g61)) + ((g311) & (!g312) & (g313) & (g314) & (g60) & (g61)) + ((g311) & (g312) & (!g313) & (!g314) & (!g60) & (!g61)) + ((g311) & (g312) & (!g313) & (!g314) & (g60) & (!g61)) + ((g311) & (g312) & (!g313) & (g314) & (!g60) & (!g61)) + ((g311) & (g312) & (!g313) & (g314) & (g60) & (!g61)) + ((g311) & (g312) & (!g313) & (g314) & (g60) & (g61)) + ((g311) & (g312) & (g313) & (!g314) & (!g60) & (!g61)) + ((g311) & (g312) & (g313) & (!g314) & (!g60) & (g61)) + ((g311) & (g312) & (g313) & (!g314) & (g60) & (!g61)) + ((g311) & (g312) & (g313) & (g314) & (!g60) & (!g61)) + ((g311) & (g312) & (g313) & (g314) & (!g60) & (g61)) + ((g311) & (g312) & (g313) & (g314) & (g60) & (!g61)) + ((g311) & (g312) & (g313) & (g314) & (g60) & (g61)));
	assign g316 = (((!g300) & (!g305) & (!g310) & (g315) & (g42) & (g43)) + ((!g300) & (!g305) & (g310) & (!g315) & (!g42) & (g43)) + ((!g300) & (!g305) & (g310) & (g315) & (!g42) & (g43)) + ((!g300) & (!g305) & (g310) & (g315) & (g42) & (g43)) + ((!g300) & (g305) & (!g310) & (!g315) & (g42) & (!g43)) + ((!g300) & (g305) & (!g310) & (g315) & (g42) & (!g43)) + ((!g300) & (g305) & (!g310) & (g315) & (g42) & (g43)) + ((!g300) & (g305) & (g310) & (!g315) & (!g42) & (g43)) + ((!g300) & (g305) & (g310) & (!g315) & (g42) & (!g43)) + ((!g300) & (g305) & (g310) & (g315) & (!g42) & (g43)) + ((!g300) & (g305) & (g310) & (g315) & (g42) & (!g43)) + ((!g300) & (g305) & (g310) & (g315) & (g42) & (g43)) + ((g300) & (!g305) & (!g310) & (!g315) & (!g42) & (!g43)) + ((g300) & (!g305) & (!g310) & (g315) & (!g42) & (!g43)) + ((g300) & (!g305) & (!g310) & (g315) & (g42) & (g43)) + ((g300) & (!g305) & (g310) & (!g315) & (!g42) & (!g43)) + ((g300) & (!g305) & (g310) & (!g315) & (!g42) & (g43)) + ((g300) & (!g305) & (g310) & (g315) & (!g42) & (!g43)) + ((g300) & (!g305) & (g310) & (g315) & (!g42) & (g43)) + ((g300) & (!g305) & (g310) & (g315) & (g42) & (g43)) + ((g300) & (g305) & (!g310) & (!g315) & (!g42) & (!g43)) + ((g300) & (g305) & (!g310) & (!g315) & (g42) & (!g43)) + ((g300) & (g305) & (!g310) & (g315) & (!g42) & (!g43)) + ((g300) & (g305) & (!g310) & (g315) & (g42) & (!g43)) + ((g300) & (g305) & (!g310) & (g315) & (g42) & (g43)) + ((g300) & (g305) & (g310) & (!g315) & (!g42) & (!g43)) + ((g300) & (g305) & (g310) & (!g315) & (!g42) & (g43)) + ((g300) & (g305) & (g310) & (!g315) & (g42) & (!g43)) + ((g300) & (g305) & (g310) & (g315) & (!g42) & (!g43)) + ((g300) & (g305) & (g310) & (g315) & (!g42) & (g43)) + ((g300) & (g305) & (g310) & (g315) & (g42) & (!g43)) + ((g300) & (g305) & (g310) & (g315) & (g42) & (g43)));
	assign g7245 = (((!g832) & (g1204) & (!g317)) + ((!g832) & (g1204) & (g317)) + ((g832) & (!g1204) & (g317)) + ((g832) & (g1204) & (g317)));
	assign g318 = (((!g34) & (!reset) & (!g316) & (g317)) + ((!g34) & (!reset) & (g316) & (g317)) + ((g34) & (!reset) & (g316) & (!g317)) + ((g34) & (!reset) & (g316) & (g317)));
	assign g323 = (((!g319) & (!g320) & (!g321) & (g322) & (g42) & (g43)) + ((!g319) & (!g320) & (g321) & (!g322) & (!g42) & (g43)) + ((!g319) & (!g320) & (g321) & (g322) & (!g42) & (g43)) + ((!g319) & (!g320) & (g321) & (g322) & (g42) & (g43)) + ((!g319) & (g320) & (!g321) & (!g322) & (g42) & (!g43)) + ((!g319) & (g320) & (!g321) & (g322) & (g42) & (!g43)) + ((!g319) & (g320) & (!g321) & (g322) & (g42) & (g43)) + ((!g319) & (g320) & (g321) & (!g322) & (!g42) & (g43)) + ((!g319) & (g320) & (g321) & (!g322) & (g42) & (!g43)) + ((!g319) & (g320) & (g321) & (g322) & (!g42) & (g43)) + ((!g319) & (g320) & (g321) & (g322) & (g42) & (!g43)) + ((!g319) & (g320) & (g321) & (g322) & (g42) & (g43)) + ((g319) & (!g320) & (!g321) & (!g322) & (!g42) & (!g43)) + ((g319) & (!g320) & (!g321) & (g322) & (!g42) & (!g43)) + ((g319) & (!g320) & (!g321) & (g322) & (g42) & (g43)) + ((g319) & (!g320) & (g321) & (!g322) & (!g42) & (!g43)) + ((g319) & (!g320) & (g321) & (!g322) & (!g42) & (g43)) + ((g319) & (!g320) & (g321) & (g322) & (!g42) & (!g43)) + ((g319) & (!g320) & (g321) & (g322) & (!g42) & (g43)) + ((g319) & (!g320) & (g321) & (g322) & (g42) & (g43)) + ((g319) & (g320) & (!g321) & (!g322) & (!g42) & (!g43)) + ((g319) & (g320) & (!g321) & (!g322) & (g42) & (!g43)) + ((g319) & (g320) & (!g321) & (g322) & (!g42) & (!g43)) + ((g319) & (g320) & (!g321) & (g322) & (g42) & (!g43)) + ((g319) & (g320) & (!g321) & (g322) & (g42) & (g43)) + ((g319) & (g320) & (g321) & (!g322) & (!g42) & (!g43)) + ((g319) & (g320) & (g321) & (!g322) & (!g42) & (g43)) + ((g319) & (g320) & (g321) & (!g322) & (g42) & (!g43)) + ((g319) & (g320) & (g321) & (g322) & (!g42) & (!g43)) + ((g319) & (g320) & (g321) & (g322) & (!g42) & (g43)) + ((g319) & (g320) & (g321) & (g322) & (g42) & (!g43)) + ((g319) & (g320) & (g321) & (g322) & (g42) & (g43)));
	assign g328 = (((!g324) & (!g325) & (!g326) & (g327) & (g42) & (g43)) + ((!g324) & (!g325) & (g326) & (!g327) & (!g42) & (g43)) + ((!g324) & (!g325) & (g326) & (g327) & (!g42) & (g43)) + ((!g324) & (!g325) & (g326) & (g327) & (g42) & (g43)) + ((!g324) & (g325) & (!g326) & (!g327) & (g42) & (!g43)) + ((!g324) & (g325) & (!g326) & (g327) & (g42) & (!g43)) + ((!g324) & (g325) & (!g326) & (g327) & (g42) & (g43)) + ((!g324) & (g325) & (g326) & (!g327) & (!g42) & (g43)) + ((!g324) & (g325) & (g326) & (!g327) & (g42) & (!g43)) + ((!g324) & (g325) & (g326) & (g327) & (!g42) & (g43)) + ((!g324) & (g325) & (g326) & (g327) & (g42) & (!g43)) + ((!g324) & (g325) & (g326) & (g327) & (g42) & (g43)) + ((g324) & (!g325) & (!g326) & (!g327) & (!g42) & (!g43)) + ((g324) & (!g325) & (!g326) & (g327) & (!g42) & (!g43)) + ((g324) & (!g325) & (!g326) & (g327) & (g42) & (g43)) + ((g324) & (!g325) & (g326) & (!g327) & (!g42) & (!g43)) + ((g324) & (!g325) & (g326) & (!g327) & (!g42) & (g43)) + ((g324) & (!g325) & (g326) & (g327) & (!g42) & (!g43)) + ((g324) & (!g325) & (g326) & (g327) & (!g42) & (g43)) + ((g324) & (!g325) & (g326) & (g327) & (g42) & (g43)) + ((g324) & (g325) & (!g326) & (!g327) & (!g42) & (!g43)) + ((g324) & (g325) & (!g326) & (!g327) & (g42) & (!g43)) + ((g324) & (g325) & (!g326) & (g327) & (!g42) & (!g43)) + ((g324) & (g325) & (!g326) & (g327) & (g42) & (!g43)) + ((g324) & (g325) & (!g326) & (g327) & (g42) & (g43)) + ((g324) & (g325) & (g326) & (!g327) & (!g42) & (!g43)) + ((g324) & (g325) & (g326) & (!g327) & (!g42) & (g43)) + ((g324) & (g325) & (g326) & (!g327) & (g42) & (!g43)) + ((g324) & (g325) & (g326) & (g327) & (!g42) & (!g43)) + ((g324) & (g325) & (g326) & (g327) & (!g42) & (g43)) + ((g324) & (g325) & (g326) & (g327) & (g42) & (!g43)) + ((g324) & (g325) & (g326) & (g327) & (g42) & (g43)));
	assign g333 = (((!g329) & (!g330) & (!g331) & (g332) & (g42) & (g43)) + ((!g329) & (!g330) & (g331) & (!g332) & (!g42) & (g43)) + ((!g329) & (!g330) & (g331) & (g332) & (!g42) & (g43)) + ((!g329) & (!g330) & (g331) & (g332) & (g42) & (g43)) + ((!g329) & (g330) & (!g331) & (!g332) & (g42) & (!g43)) + ((!g329) & (g330) & (!g331) & (g332) & (g42) & (!g43)) + ((!g329) & (g330) & (!g331) & (g332) & (g42) & (g43)) + ((!g329) & (g330) & (g331) & (!g332) & (!g42) & (g43)) + ((!g329) & (g330) & (g331) & (!g332) & (g42) & (!g43)) + ((!g329) & (g330) & (g331) & (g332) & (!g42) & (g43)) + ((!g329) & (g330) & (g331) & (g332) & (g42) & (!g43)) + ((!g329) & (g330) & (g331) & (g332) & (g42) & (g43)) + ((g329) & (!g330) & (!g331) & (!g332) & (!g42) & (!g43)) + ((g329) & (!g330) & (!g331) & (g332) & (!g42) & (!g43)) + ((g329) & (!g330) & (!g331) & (g332) & (g42) & (g43)) + ((g329) & (!g330) & (g331) & (!g332) & (!g42) & (!g43)) + ((g329) & (!g330) & (g331) & (!g332) & (!g42) & (g43)) + ((g329) & (!g330) & (g331) & (g332) & (!g42) & (!g43)) + ((g329) & (!g330) & (g331) & (g332) & (!g42) & (g43)) + ((g329) & (!g330) & (g331) & (g332) & (g42) & (g43)) + ((g329) & (g330) & (!g331) & (!g332) & (!g42) & (!g43)) + ((g329) & (g330) & (!g331) & (!g332) & (g42) & (!g43)) + ((g329) & (g330) & (!g331) & (g332) & (!g42) & (!g43)) + ((g329) & (g330) & (!g331) & (g332) & (g42) & (!g43)) + ((g329) & (g330) & (!g331) & (g332) & (g42) & (g43)) + ((g329) & (g330) & (g331) & (!g332) & (!g42) & (!g43)) + ((g329) & (g330) & (g331) & (!g332) & (!g42) & (g43)) + ((g329) & (g330) & (g331) & (!g332) & (g42) & (!g43)) + ((g329) & (g330) & (g331) & (g332) & (!g42) & (!g43)) + ((g329) & (g330) & (g331) & (g332) & (!g42) & (g43)) + ((g329) & (g330) & (g331) & (g332) & (g42) & (!g43)) + ((g329) & (g330) & (g331) & (g332) & (g42) & (g43)));
	assign g338 = (((!g334) & (!g335) & (!g336) & (g337) & (g42) & (g43)) + ((!g334) & (!g335) & (g336) & (!g337) & (!g42) & (g43)) + ((!g334) & (!g335) & (g336) & (g337) & (!g42) & (g43)) + ((!g334) & (!g335) & (g336) & (g337) & (g42) & (g43)) + ((!g334) & (g335) & (!g336) & (!g337) & (g42) & (!g43)) + ((!g334) & (g335) & (!g336) & (g337) & (g42) & (!g43)) + ((!g334) & (g335) & (!g336) & (g337) & (g42) & (g43)) + ((!g334) & (g335) & (g336) & (!g337) & (!g42) & (g43)) + ((!g334) & (g335) & (g336) & (!g337) & (g42) & (!g43)) + ((!g334) & (g335) & (g336) & (g337) & (!g42) & (g43)) + ((!g334) & (g335) & (g336) & (g337) & (g42) & (!g43)) + ((!g334) & (g335) & (g336) & (g337) & (g42) & (g43)) + ((g334) & (!g335) & (!g336) & (!g337) & (!g42) & (!g43)) + ((g334) & (!g335) & (!g336) & (g337) & (!g42) & (!g43)) + ((g334) & (!g335) & (!g336) & (g337) & (g42) & (g43)) + ((g334) & (!g335) & (g336) & (!g337) & (!g42) & (!g43)) + ((g334) & (!g335) & (g336) & (!g337) & (!g42) & (g43)) + ((g334) & (!g335) & (g336) & (g337) & (!g42) & (!g43)) + ((g334) & (!g335) & (g336) & (g337) & (!g42) & (g43)) + ((g334) & (!g335) & (g336) & (g337) & (g42) & (g43)) + ((g334) & (g335) & (!g336) & (!g337) & (!g42) & (!g43)) + ((g334) & (g335) & (!g336) & (!g337) & (g42) & (!g43)) + ((g334) & (g335) & (!g336) & (g337) & (!g42) & (!g43)) + ((g334) & (g335) & (!g336) & (g337) & (g42) & (!g43)) + ((g334) & (g335) & (!g336) & (g337) & (g42) & (g43)) + ((g334) & (g335) & (g336) & (!g337) & (!g42) & (!g43)) + ((g334) & (g335) & (g336) & (!g337) & (!g42) & (g43)) + ((g334) & (g335) & (g336) & (!g337) & (g42) & (!g43)) + ((g334) & (g335) & (g336) & (g337) & (!g42) & (!g43)) + ((g334) & (g335) & (g336) & (g337) & (!g42) & (g43)) + ((g334) & (g335) & (g336) & (g337) & (g42) & (!g43)) + ((g334) & (g335) & (g336) & (g337) & (g42) & (g43)));
	assign g339 = (((!g323) & (!g328) & (!g333) & (g338) & (g60) & (g61)) + ((!g323) & (!g328) & (g333) & (!g338) & (!g60) & (g61)) + ((!g323) & (!g328) & (g333) & (g338) & (!g60) & (g61)) + ((!g323) & (!g328) & (g333) & (g338) & (g60) & (g61)) + ((!g323) & (g328) & (!g333) & (!g338) & (g60) & (!g61)) + ((!g323) & (g328) & (!g333) & (g338) & (g60) & (!g61)) + ((!g323) & (g328) & (!g333) & (g338) & (g60) & (g61)) + ((!g323) & (g328) & (g333) & (!g338) & (!g60) & (g61)) + ((!g323) & (g328) & (g333) & (!g338) & (g60) & (!g61)) + ((!g323) & (g328) & (g333) & (g338) & (!g60) & (g61)) + ((!g323) & (g328) & (g333) & (g338) & (g60) & (!g61)) + ((!g323) & (g328) & (g333) & (g338) & (g60) & (g61)) + ((g323) & (!g328) & (!g333) & (!g338) & (!g60) & (!g61)) + ((g323) & (!g328) & (!g333) & (g338) & (!g60) & (!g61)) + ((g323) & (!g328) & (!g333) & (g338) & (g60) & (g61)) + ((g323) & (!g328) & (g333) & (!g338) & (!g60) & (!g61)) + ((g323) & (!g328) & (g333) & (!g338) & (!g60) & (g61)) + ((g323) & (!g328) & (g333) & (g338) & (!g60) & (!g61)) + ((g323) & (!g328) & (g333) & (g338) & (!g60) & (g61)) + ((g323) & (!g328) & (g333) & (g338) & (g60) & (g61)) + ((g323) & (g328) & (!g333) & (!g338) & (!g60) & (!g61)) + ((g323) & (g328) & (!g333) & (!g338) & (g60) & (!g61)) + ((g323) & (g328) & (!g333) & (g338) & (!g60) & (!g61)) + ((g323) & (g328) & (!g333) & (g338) & (g60) & (!g61)) + ((g323) & (g328) & (!g333) & (g338) & (g60) & (g61)) + ((g323) & (g328) & (g333) & (!g338) & (!g60) & (!g61)) + ((g323) & (g328) & (g333) & (!g338) & (!g60) & (g61)) + ((g323) & (g328) & (g333) & (!g338) & (g60) & (!g61)) + ((g323) & (g328) & (g333) & (g338) & (!g60) & (!g61)) + ((g323) & (g328) & (g333) & (g338) & (!g60) & (g61)) + ((g323) & (g328) & (g333) & (g338) & (g60) & (!g61)) + ((g323) & (g328) & (g333) & (g338) & (g60) & (g61)));
	assign g7246 = (((!g832) & (g1237) & (!g340)) + ((!g832) & (g1237) & (g340)) + ((g832) & (!g1237) & (g340)) + ((g832) & (g1237) & (g340)));
	assign g341 = (((!g34) & (!reset) & (!g339) & (g340)) + ((!g34) & (!reset) & (g339) & (g340)) + ((g34) & (!reset) & (g339) & (!g340)) + ((g34) & (!reset) & (g339) & (g340)));
	assign g346 = (((!g342) & (!g343) & (!g344) & (g345) & (g60) & (g61)) + ((!g342) & (!g343) & (g344) & (!g345) & (!g60) & (g61)) + ((!g342) & (!g343) & (g344) & (g345) & (!g60) & (g61)) + ((!g342) & (!g343) & (g344) & (g345) & (g60) & (g61)) + ((!g342) & (g343) & (!g344) & (!g345) & (g60) & (!g61)) + ((!g342) & (g343) & (!g344) & (g345) & (g60) & (!g61)) + ((!g342) & (g343) & (!g344) & (g345) & (g60) & (g61)) + ((!g342) & (g343) & (g344) & (!g345) & (!g60) & (g61)) + ((!g342) & (g343) & (g344) & (!g345) & (g60) & (!g61)) + ((!g342) & (g343) & (g344) & (g345) & (!g60) & (g61)) + ((!g342) & (g343) & (g344) & (g345) & (g60) & (!g61)) + ((!g342) & (g343) & (g344) & (g345) & (g60) & (g61)) + ((g342) & (!g343) & (!g344) & (!g345) & (!g60) & (!g61)) + ((g342) & (!g343) & (!g344) & (g345) & (!g60) & (!g61)) + ((g342) & (!g343) & (!g344) & (g345) & (g60) & (g61)) + ((g342) & (!g343) & (g344) & (!g345) & (!g60) & (!g61)) + ((g342) & (!g343) & (g344) & (!g345) & (!g60) & (g61)) + ((g342) & (!g343) & (g344) & (g345) & (!g60) & (!g61)) + ((g342) & (!g343) & (g344) & (g345) & (!g60) & (g61)) + ((g342) & (!g343) & (g344) & (g345) & (g60) & (g61)) + ((g342) & (g343) & (!g344) & (!g345) & (!g60) & (!g61)) + ((g342) & (g343) & (!g344) & (!g345) & (g60) & (!g61)) + ((g342) & (g343) & (!g344) & (g345) & (!g60) & (!g61)) + ((g342) & (g343) & (!g344) & (g345) & (g60) & (!g61)) + ((g342) & (g343) & (!g344) & (g345) & (g60) & (g61)) + ((g342) & (g343) & (g344) & (!g345) & (!g60) & (!g61)) + ((g342) & (g343) & (g344) & (!g345) & (!g60) & (g61)) + ((g342) & (g343) & (g344) & (!g345) & (g60) & (!g61)) + ((g342) & (g343) & (g344) & (g345) & (!g60) & (!g61)) + ((g342) & (g343) & (g344) & (g345) & (!g60) & (g61)) + ((g342) & (g343) & (g344) & (g345) & (g60) & (!g61)) + ((g342) & (g343) & (g344) & (g345) & (g60) & (g61)));
	assign g351 = (((!g347) & (!g348) & (!g349) & (g350) & (g60) & (g61)) + ((!g347) & (!g348) & (g349) & (!g350) & (!g60) & (g61)) + ((!g347) & (!g348) & (g349) & (g350) & (!g60) & (g61)) + ((!g347) & (!g348) & (g349) & (g350) & (g60) & (g61)) + ((!g347) & (g348) & (!g349) & (!g350) & (g60) & (!g61)) + ((!g347) & (g348) & (!g349) & (g350) & (g60) & (!g61)) + ((!g347) & (g348) & (!g349) & (g350) & (g60) & (g61)) + ((!g347) & (g348) & (g349) & (!g350) & (!g60) & (g61)) + ((!g347) & (g348) & (g349) & (!g350) & (g60) & (!g61)) + ((!g347) & (g348) & (g349) & (g350) & (!g60) & (g61)) + ((!g347) & (g348) & (g349) & (g350) & (g60) & (!g61)) + ((!g347) & (g348) & (g349) & (g350) & (g60) & (g61)) + ((g347) & (!g348) & (!g349) & (!g350) & (!g60) & (!g61)) + ((g347) & (!g348) & (!g349) & (g350) & (!g60) & (!g61)) + ((g347) & (!g348) & (!g349) & (g350) & (g60) & (g61)) + ((g347) & (!g348) & (g349) & (!g350) & (!g60) & (!g61)) + ((g347) & (!g348) & (g349) & (!g350) & (!g60) & (g61)) + ((g347) & (!g348) & (g349) & (g350) & (!g60) & (!g61)) + ((g347) & (!g348) & (g349) & (g350) & (!g60) & (g61)) + ((g347) & (!g348) & (g349) & (g350) & (g60) & (g61)) + ((g347) & (g348) & (!g349) & (!g350) & (!g60) & (!g61)) + ((g347) & (g348) & (!g349) & (!g350) & (g60) & (!g61)) + ((g347) & (g348) & (!g349) & (g350) & (!g60) & (!g61)) + ((g347) & (g348) & (!g349) & (g350) & (g60) & (!g61)) + ((g347) & (g348) & (!g349) & (g350) & (g60) & (g61)) + ((g347) & (g348) & (g349) & (!g350) & (!g60) & (!g61)) + ((g347) & (g348) & (g349) & (!g350) & (!g60) & (g61)) + ((g347) & (g348) & (g349) & (!g350) & (g60) & (!g61)) + ((g347) & (g348) & (g349) & (g350) & (!g60) & (!g61)) + ((g347) & (g348) & (g349) & (g350) & (!g60) & (g61)) + ((g347) & (g348) & (g349) & (g350) & (g60) & (!g61)) + ((g347) & (g348) & (g349) & (g350) & (g60) & (g61)));
	assign g356 = (((!g352) & (!g353) & (!g354) & (g355) & (g60) & (g61)) + ((!g352) & (!g353) & (g354) & (!g355) & (!g60) & (g61)) + ((!g352) & (!g353) & (g354) & (g355) & (!g60) & (g61)) + ((!g352) & (!g353) & (g354) & (g355) & (g60) & (g61)) + ((!g352) & (g353) & (!g354) & (!g355) & (g60) & (!g61)) + ((!g352) & (g353) & (!g354) & (g355) & (g60) & (!g61)) + ((!g352) & (g353) & (!g354) & (g355) & (g60) & (g61)) + ((!g352) & (g353) & (g354) & (!g355) & (!g60) & (g61)) + ((!g352) & (g353) & (g354) & (!g355) & (g60) & (!g61)) + ((!g352) & (g353) & (g354) & (g355) & (!g60) & (g61)) + ((!g352) & (g353) & (g354) & (g355) & (g60) & (!g61)) + ((!g352) & (g353) & (g354) & (g355) & (g60) & (g61)) + ((g352) & (!g353) & (!g354) & (!g355) & (!g60) & (!g61)) + ((g352) & (!g353) & (!g354) & (g355) & (!g60) & (!g61)) + ((g352) & (!g353) & (!g354) & (g355) & (g60) & (g61)) + ((g352) & (!g353) & (g354) & (!g355) & (!g60) & (!g61)) + ((g352) & (!g353) & (g354) & (!g355) & (!g60) & (g61)) + ((g352) & (!g353) & (g354) & (g355) & (!g60) & (!g61)) + ((g352) & (!g353) & (g354) & (g355) & (!g60) & (g61)) + ((g352) & (!g353) & (g354) & (g355) & (g60) & (g61)) + ((g352) & (g353) & (!g354) & (!g355) & (!g60) & (!g61)) + ((g352) & (g353) & (!g354) & (!g355) & (g60) & (!g61)) + ((g352) & (g353) & (!g354) & (g355) & (!g60) & (!g61)) + ((g352) & (g353) & (!g354) & (g355) & (g60) & (!g61)) + ((g352) & (g353) & (!g354) & (g355) & (g60) & (g61)) + ((g352) & (g353) & (g354) & (!g355) & (!g60) & (!g61)) + ((g352) & (g353) & (g354) & (!g355) & (!g60) & (g61)) + ((g352) & (g353) & (g354) & (!g355) & (g60) & (!g61)) + ((g352) & (g353) & (g354) & (g355) & (!g60) & (!g61)) + ((g352) & (g353) & (g354) & (g355) & (!g60) & (g61)) + ((g352) & (g353) & (g354) & (g355) & (g60) & (!g61)) + ((g352) & (g353) & (g354) & (g355) & (g60) & (g61)));
	assign g361 = (((!g357) & (!g358) & (!g359) & (g360) & (g60) & (g61)) + ((!g357) & (!g358) & (g359) & (!g360) & (!g60) & (g61)) + ((!g357) & (!g358) & (g359) & (g360) & (!g60) & (g61)) + ((!g357) & (!g358) & (g359) & (g360) & (g60) & (g61)) + ((!g357) & (g358) & (!g359) & (!g360) & (g60) & (!g61)) + ((!g357) & (g358) & (!g359) & (g360) & (g60) & (!g61)) + ((!g357) & (g358) & (!g359) & (g360) & (g60) & (g61)) + ((!g357) & (g358) & (g359) & (!g360) & (!g60) & (g61)) + ((!g357) & (g358) & (g359) & (!g360) & (g60) & (!g61)) + ((!g357) & (g358) & (g359) & (g360) & (!g60) & (g61)) + ((!g357) & (g358) & (g359) & (g360) & (g60) & (!g61)) + ((!g357) & (g358) & (g359) & (g360) & (g60) & (g61)) + ((g357) & (!g358) & (!g359) & (!g360) & (!g60) & (!g61)) + ((g357) & (!g358) & (!g359) & (g360) & (!g60) & (!g61)) + ((g357) & (!g358) & (!g359) & (g360) & (g60) & (g61)) + ((g357) & (!g358) & (g359) & (!g360) & (!g60) & (!g61)) + ((g357) & (!g358) & (g359) & (!g360) & (!g60) & (g61)) + ((g357) & (!g358) & (g359) & (g360) & (!g60) & (!g61)) + ((g357) & (!g358) & (g359) & (g360) & (!g60) & (g61)) + ((g357) & (!g358) & (g359) & (g360) & (g60) & (g61)) + ((g357) & (g358) & (!g359) & (!g360) & (!g60) & (!g61)) + ((g357) & (g358) & (!g359) & (!g360) & (g60) & (!g61)) + ((g357) & (g358) & (!g359) & (g360) & (!g60) & (!g61)) + ((g357) & (g358) & (!g359) & (g360) & (g60) & (!g61)) + ((g357) & (g358) & (!g359) & (g360) & (g60) & (g61)) + ((g357) & (g358) & (g359) & (!g360) & (!g60) & (!g61)) + ((g357) & (g358) & (g359) & (!g360) & (!g60) & (g61)) + ((g357) & (g358) & (g359) & (!g360) & (g60) & (!g61)) + ((g357) & (g358) & (g359) & (g360) & (!g60) & (!g61)) + ((g357) & (g358) & (g359) & (g360) & (!g60) & (g61)) + ((g357) & (g358) & (g359) & (g360) & (g60) & (!g61)) + ((g357) & (g358) & (g359) & (g360) & (g60) & (g61)));
	assign g362 = (((!g346) & (!g351) & (!g356) & (g361) & (g42) & (g43)) + ((!g346) & (!g351) & (g356) & (!g361) & (!g42) & (g43)) + ((!g346) & (!g351) & (g356) & (g361) & (!g42) & (g43)) + ((!g346) & (!g351) & (g356) & (g361) & (g42) & (g43)) + ((!g346) & (g351) & (!g356) & (!g361) & (g42) & (!g43)) + ((!g346) & (g351) & (!g356) & (g361) & (g42) & (!g43)) + ((!g346) & (g351) & (!g356) & (g361) & (g42) & (g43)) + ((!g346) & (g351) & (g356) & (!g361) & (!g42) & (g43)) + ((!g346) & (g351) & (g356) & (!g361) & (g42) & (!g43)) + ((!g346) & (g351) & (g356) & (g361) & (!g42) & (g43)) + ((!g346) & (g351) & (g356) & (g361) & (g42) & (!g43)) + ((!g346) & (g351) & (g356) & (g361) & (g42) & (g43)) + ((g346) & (!g351) & (!g356) & (!g361) & (!g42) & (!g43)) + ((g346) & (!g351) & (!g356) & (g361) & (!g42) & (!g43)) + ((g346) & (!g351) & (!g356) & (g361) & (g42) & (g43)) + ((g346) & (!g351) & (g356) & (!g361) & (!g42) & (!g43)) + ((g346) & (!g351) & (g356) & (!g361) & (!g42) & (g43)) + ((g346) & (!g351) & (g356) & (g361) & (!g42) & (!g43)) + ((g346) & (!g351) & (g356) & (g361) & (!g42) & (g43)) + ((g346) & (!g351) & (g356) & (g361) & (g42) & (g43)) + ((g346) & (g351) & (!g356) & (!g361) & (!g42) & (!g43)) + ((g346) & (g351) & (!g356) & (!g361) & (g42) & (!g43)) + ((g346) & (g351) & (!g356) & (g361) & (!g42) & (!g43)) + ((g346) & (g351) & (!g356) & (g361) & (g42) & (!g43)) + ((g346) & (g351) & (!g356) & (g361) & (g42) & (g43)) + ((g346) & (g351) & (g356) & (!g361) & (!g42) & (!g43)) + ((g346) & (g351) & (g356) & (!g361) & (!g42) & (g43)) + ((g346) & (g351) & (g356) & (!g361) & (g42) & (!g43)) + ((g346) & (g351) & (g356) & (g361) & (!g42) & (!g43)) + ((g346) & (g351) & (g356) & (g361) & (!g42) & (g43)) + ((g346) & (g351) & (g356) & (g361) & (g42) & (!g43)) + ((g346) & (g351) & (g356) & (g361) & (g42) & (g43)));
	assign g7247 = (((!g832) & (g1271) & (!g363)) + ((!g832) & (g1271) & (g363)) + ((g832) & (!g1271) & (g363)) + ((g832) & (g1271) & (g363)));
	assign g364 = (((!g34) & (!reset) & (!g362) & (g363)) + ((!g34) & (!reset) & (g362) & (g363)) + ((g34) & (!reset) & (g362) & (!g363)) + ((g34) & (!reset) & (g362) & (g363)));
	assign g369 = (((!g365) & (!g366) & (!g367) & (g368) & (g42) & (g43)) + ((!g365) & (!g366) & (g367) & (!g368) & (!g42) & (g43)) + ((!g365) & (!g366) & (g367) & (g368) & (!g42) & (g43)) + ((!g365) & (!g366) & (g367) & (g368) & (g42) & (g43)) + ((!g365) & (g366) & (!g367) & (!g368) & (g42) & (!g43)) + ((!g365) & (g366) & (!g367) & (g368) & (g42) & (!g43)) + ((!g365) & (g366) & (!g367) & (g368) & (g42) & (g43)) + ((!g365) & (g366) & (g367) & (!g368) & (!g42) & (g43)) + ((!g365) & (g366) & (g367) & (!g368) & (g42) & (!g43)) + ((!g365) & (g366) & (g367) & (g368) & (!g42) & (g43)) + ((!g365) & (g366) & (g367) & (g368) & (g42) & (!g43)) + ((!g365) & (g366) & (g367) & (g368) & (g42) & (g43)) + ((g365) & (!g366) & (!g367) & (!g368) & (!g42) & (!g43)) + ((g365) & (!g366) & (!g367) & (g368) & (!g42) & (!g43)) + ((g365) & (!g366) & (!g367) & (g368) & (g42) & (g43)) + ((g365) & (!g366) & (g367) & (!g368) & (!g42) & (!g43)) + ((g365) & (!g366) & (g367) & (!g368) & (!g42) & (g43)) + ((g365) & (!g366) & (g367) & (g368) & (!g42) & (!g43)) + ((g365) & (!g366) & (g367) & (g368) & (!g42) & (g43)) + ((g365) & (!g366) & (g367) & (g368) & (g42) & (g43)) + ((g365) & (g366) & (!g367) & (!g368) & (!g42) & (!g43)) + ((g365) & (g366) & (!g367) & (!g368) & (g42) & (!g43)) + ((g365) & (g366) & (!g367) & (g368) & (!g42) & (!g43)) + ((g365) & (g366) & (!g367) & (g368) & (g42) & (!g43)) + ((g365) & (g366) & (!g367) & (g368) & (g42) & (g43)) + ((g365) & (g366) & (g367) & (!g368) & (!g42) & (!g43)) + ((g365) & (g366) & (g367) & (!g368) & (!g42) & (g43)) + ((g365) & (g366) & (g367) & (!g368) & (g42) & (!g43)) + ((g365) & (g366) & (g367) & (g368) & (!g42) & (!g43)) + ((g365) & (g366) & (g367) & (g368) & (!g42) & (g43)) + ((g365) & (g366) & (g367) & (g368) & (g42) & (!g43)) + ((g365) & (g366) & (g367) & (g368) & (g42) & (g43)));
	assign g374 = (((!g370) & (!g371) & (!g372) & (g373) & (g42) & (g43)) + ((!g370) & (!g371) & (g372) & (!g373) & (!g42) & (g43)) + ((!g370) & (!g371) & (g372) & (g373) & (!g42) & (g43)) + ((!g370) & (!g371) & (g372) & (g373) & (g42) & (g43)) + ((!g370) & (g371) & (!g372) & (!g373) & (g42) & (!g43)) + ((!g370) & (g371) & (!g372) & (g373) & (g42) & (!g43)) + ((!g370) & (g371) & (!g372) & (g373) & (g42) & (g43)) + ((!g370) & (g371) & (g372) & (!g373) & (!g42) & (g43)) + ((!g370) & (g371) & (g372) & (!g373) & (g42) & (!g43)) + ((!g370) & (g371) & (g372) & (g373) & (!g42) & (g43)) + ((!g370) & (g371) & (g372) & (g373) & (g42) & (!g43)) + ((!g370) & (g371) & (g372) & (g373) & (g42) & (g43)) + ((g370) & (!g371) & (!g372) & (!g373) & (!g42) & (!g43)) + ((g370) & (!g371) & (!g372) & (g373) & (!g42) & (!g43)) + ((g370) & (!g371) & (!g372) & (g373) & (g42) & (g43)) + ((g370) & (!g371) & (g372) & (!g373) & (!g42) & (!g43)) + ((g370) & (!g371) & (g372) & (!g373) & (!g42) & (g43)) + ((g370) & (!g371) & (g372) & (g373) & (!g42) & (!g43)) + ((g370) & (!g371) & (g372) & (g373) & (!g42) & (g43)) + ((g370) & (!g371) & (g372) & (g373) & (g42) & (g43)) + ((g370) & (g371) & (!g372) & (!g373) & (!g42) & (!g43)) + ((g370) & (g371) & (!g372) & (!g373) & (g42) & (!g43)) + ((g370) & (g371) & (!g372) & (g373) & (!g42) & (!g43)) + ((g370) & (g371) & (!g372) & (g373) & (g42) & (!g43)) + ((g370) & (g371) & (!g372) & (g373) & (g42) & (g43)) + ((g370) & (g371) & (g372) & (!g373) & (!g42) & (!g43)) + ((g370) & (g371) & (g372) & (!g373) & (!g42) & (g43)) + ((g370) & (g371) & (g372) & (!g373) & (g42) & (!g43)) + ((g370) & (g371) & (g372) & (g373) & (!g42) & (!g43)) + ((g370) & (g371) & (g372) & (g373) & (!g42) & (g43)) + ((g370) & (g371) & (g372) & (g373) & (g42) & (!g43)) + ((g370) & (g371) & (g372) & (g373) & (g42) & (g43)));
	assign g379 = (((!g375) & (!g376) & (!g377) & (g378) & (g42) & (g43)) + ((!g375) & (!g376) & (g377) & (!g378) & (!g42) & (g43)) + ((!g375) & (!g376) & (g377) & (g378) & (!g42) & (g43)) + ((!g375) & (!g376) & (g377) & (g378) & (g42) & (g43)) + ((!g375) & (g376) & (!g377) & (!g378) & (g42) & (!g43)) + ((!g375) & (g376) & (!g377) & (g378) & (g42) & (!g43)) + ((!g375) & (g376) & (!g377) & (g378) & (g42) & (g43)) + ((!g375) & (g376) & (g377) & (!g378) & (!g42) & (g43)) + ((!g375) & (g376) & (g377) & (!g378) & (g42) & (!g43)) + ((!g375) & (g376) & (g377) & (g378) & (!g42) & (g43)) + ((!g375) & (g376) & (g377) & (g378) & (g42) & (!g43)) + ((!g375) & (g376) & (g377) & (g378) & (g42) & (g43)) + ((g375) & (!g376) & (!g377) & (!g378) & (!g42) & (!g43)) + ((g375) & (!g376) & (!g377) & (g378) & (!g42) & (!g43)) + ((g375) & (!g376) & (!g377) & (g378) & (g42) & (g43)) + ((g375) & (!g376) & (g377) & (!g378) & (!g42) & (!g43)) + ((g375) & (!g376) & (g377) & (!g378) & (!g42) & (g43)) + ((g375) & (!g376) & (g377) & (g378) & (!g42) & (!g43)) + ((g375) & (!g376) & (g377) & (g378) & (!g42) & (g43)) + ((g375) & (!g376) & (g377) & (g378) & (g42) & (g43)) + ((g375) & (g376) & (!g377) & (!g378) & (!g42) & (!g43)) + ((g375) & (g376) & (!g377) & (!g378) & (g42) & (!g43)) + ((g375) & (g376) & (!g377) & (g378) & (!g42) & (!g43)) + ((g375) & (g376) & (!g377) & (g378) & (g42) & (!g43)) + ((g375) & (g376) & (!g377) & (g378) & (g42) & (g43)) + ((g375) & (g376) & (g377) & (!g378) & (!g42) & (!g43)) + ((g375) & (g376) & (g377) & (!g378) & (!g42) & (g43)) + ((g375) & (g376) & (g377) & (!g378) & (g42) & (!g43)) + ((g375) & (g376) & (g377) & (g378) & (!g42) & (!g43)) + ((g375) & (g376) & (g377) & (g378) & (!g42) & (g43)) + ((g375) & (g376) & (g377) & (g378) & (g42) & (!g43)) + ((g375) & (g376) & (g377) & (g378) & (g42) & (g43)));
	assign g384 = (((!g380) & (!g381) & (!g382) & (g383) & (g42) & (g43)) + ((!g380) & (!g381) & (g382) & (!g383) & (!g42) & (g43)) + ((!g380) & (!g381) & (g382) & (g383) & (!g42) & (g43)) + ((!g380) & (!g381) & (g382) & (g383) & (g42) & (g43)) + ((!g380) & (g381) & (!g382) & (!g383) & (g42) & (!g43)) + ((!g380) & (g381) & (!g382) & (g383) & (g42) & (!g43)) + ((!g380) & (g381) & (!g382) & (g383) & (g42) & (g43)) + ((!g380) & (g381) & (g382) & (!g383) & (!g42) & (g43)) + ((!g380) & (g381) & (g382) & (!g383) & (g42) & (!g43)) + ((!g380) & (g381) & (g382) & (g383) & (!g42) & (g43)) + ((!g380) & (g381) & (g382) & (g383) & (g42) & (!g43)) + ((!g380) & (g381) & (g382) & (g383) & (g42) & (g43)) + ((g380) & (!g381) & (!g382) & (!g383) & (!g42) & (!g43)) + ((g380) & (!g381) & (!g382) & (g383) & (!g42) & (!g43)) + ((g380) & (!g381) & (!g382) & (g383) & (g42) & (g43)) + ((g380) & (!g381) & (g382) & (!g383) & (!g42) & (!g43)) + ((g380) & (!g381) & (g382) & (!g383) & (!g42) & (g43)) + ((g380) & (!g381) & (g382) & (g383) & (!g42) & (!g43)) + ((g380) & (!g381) & (g382) & (g383) & (!g42) & (g43)) + ((g380) & (!g381) & (g382) & (g383) & (g42) & (g43)) + ((g380) & (g381) & (!g382) & (!g383) & (!g42) & (!g43)) + ((g380) & (g381) & (!g382) & (!g383) & (g42) & (!g43)) + ((g380) & (g381) & (!g382) & (g383) & (!g42) & (!g43)) + ((g380) & (g381) & (!g382) & (g383) & (g42) & (!g43)) + ((g380) & (g381) & (!g382) & (g383) & (g42) & (g43)) + ((g380) & (g381) & (g382) & (!g383) & (!g42) & (!g43)) + ((g380) & (g381) & (g382) & (!g383) & (!g42) & (g43)) + ((g380) & (g381) & (g382) & (!g383) & (g42) & (!g43)) + ((g380) & (g381) & (g382) & (g383) & (!g42) & (!g43)) + ((g380) & (g381) & (g382) & (g383) & (!g42) & (g43)) + ((g380) & (g381) & (g382) & (g383) & (g42) & (!g43)) + ((g380) & (g381) & (g382) & (g383) & (g42) & (g43)));
	assign g385 = (((!g369) & (!g374) & (!g379) & (g384) & (g60) & (g61)) + ((!g369) & (!g374) & (g379) & (!g384) & (!g60) & (g61)) + ((!g369) & (!g374) & (g379) & (g384) & (!g60) & (g61)) + ((!g369) & (!g374) & (g379) & (g384) & (g60) & (g61)) + ((!g369) & (g374) & (!g379) & (!g384) & (g60) & (!g61)) + ((!g369) & (g374) & (!g379) & (g384) & (g60) & (!g61)) + ((!g369) & (g374) & (!g379) & (g384) & (g60) & (g61)) + ((!g369) & (g374) & (g379) & (!g384) & (!g60) & (g61)) + ((!g369) & (g374) & (g379) & (!g384) & (g60) & (!g61)) + ((!g369) & (g374) & (g379) & (g384) & (!g60) & (g61)) + ((!g369) & (g374) & (g379) & (g384) & (g60) & (!g61)) + ((!g369) & (g374) & (g379) & (g384) & (g60) & (g61)) + ((g369) & (!g374) & (!g379) & (!g384) & (!g60) & (!g61)) + ((g369) & (!g374) & (!g379) & (g384) & (!g60) & (!g61)) + ((g369) & (!g374) & (!g379) & (g384) & (g60) & (g61)) + ((g369) & (!g374) & (g379) & (!g384) & (!g60) & (!g61)) + ((g369) & (!g374) & (g379) & (!g384) & (!g60) & (g61)) + ((g369) & (!g374) & (g379) & (g384) & (!g60) & (!g61)) + ((g369) & (!g374) & (g379) & (g384) & (!g60) & (g61)) + ((g369) & (!g374) & (g379) & (g384) & (g60) & (g61)) + ((g369) & (g374) & (!g379) & (!g384) & (!g60) & (!g61)) + ((g369) & (g374) & (!g379) & (!g384) & (g60) & (!g61)) + ((g369) & (g374) & (!g379) & (g384) & (!g60) & (!g61)) + ((g369) & (g374) & (!g379) & (g384) & (g60) & (!g61)) + ((g369) & (g374) & (!g379) & (g384) & (g60) & (g61)) + ((g369) & (g374) & (g379) & (!g384) & (!g60) & (!g61)) + ((g369) & (g374) & (g379) & (!g384) & (!g60) & (g61)) + ((g369) & (g374) & (g379) & (!g384) & (g60) & (!g61)) + ((g369) & (g374) & (g379) & (g384) & (!g60) & (!g61)) + ((g369) & (g374) & (g379) & (g384) & (!g60) & (g61)) + ((g369) & (g374) & (g379) & (g384) & (g60) & (!g61)) + ((g369) & (g374) & (g379) & (g384) & (g60) & (g61)));
	assign g7248 = (((!g832) & (g1305) & (!g386)) + ((!g832) & (g1305) & (g386)) + ((g832) & (!g1305) & (g386)) + ((g832) & (g1305) & (g386)));
	assign g387 = (((!g34) & (!reset) & (!g385) & (g386)) + ((!g34) & (!reset) & (g385) & (g386)) + ((g34) & (!reset) & (g385) & (!g386)) + ((g34) & (!reset) & (g385) & (g386)));
	assign g392 = (((!g388) & (!g389) & (!g390) & (g391) & (g60) & (g61)) + ((!g388) & (!g389) & (g390) & (!g391) & (!g60) & (g61)) + ((!g388) & (!g389) & (g390) & (g391) & (!g60) & (g61)) + ((!g388) & (!g389) & (g390) & (g391) & (g60) & (g61)) + ((!g388) & (g389) & (!g390) & (!g391) & (g60) & (!g61)) + ((!g388) & (g389) & (!g390) & (g391) & (g60) & (!g61)) + ((!g388) & (g389) & (!g390) & (g391) & (g60) & (g61)) + ((!g388) & (g389) & (g390) & (!g391) & (!g60) & (g61)) + ((!g388) & (g389) & (g390) & (!g391) & (g60) & (!g61)) + ((!g388) & (g389) & (g390) & (g391) & (!g60) & (g61)) + ((!g388) & (g389) & (g390) & (g391) & (g60) & (!g61)) + ((!g388) & (g389) & (g390) & (g391) & (g60) & (g61)) + ((g388) & (!g389) & (!g390) & (!g391) & (!g60) & (!g61)) + ((g388) & (!g389) & (!g390) & (g391) & (!g60) & (!g61)) + ((g388) & (!g389) & (!g390) & (g391) & (g60) & (g61)) + ((g388) & (!g389) & (g390) & (!g391) & (!g60) & (!g61)) + ((g388) & (!g389) & (g390) & (!g391) & (!g60) & (g61)) + ((g388) & (!g389) & (g390) & (g391) & (!g60) & (!g61)) + ((g388) & (!g389) & (g390) & (g391) & (!g60) & (g61)) + ((g388) & (!g389) & (g390) & (g391) & (g60) & (g61)) + ((g388) & (g389) & (!g390) & (!g391) & (!g60) & (!g61)) + ((g388) & (g389) & (!g390) & (!g391) & (g60) & (!g61)) + ((g388) & (g389) & (!g390) & (g391) & (!g60) & (!g61)) + ((g388) & (g389) & (!g390) & (g391) & (g60) & (!g61)) + ((g388) & (g389) & (!g390) & (g391) & (g60) & (g61)) + ((g388) & (g389) & (g390) & (!g391) & (!g60) & (!g61)) + ((g388) & (g389) & (g390) & (!g391) & (!g60) & (g61)) + ((g388) & (g389) & (g390) & (!g391) & (g60) & (!g61)) + ((g388) & (g389) & (g390) & (g391) & (!g60) & (!g61)) + ((g388) & (g389) & (g390) & (g391) & (!g60) & (g61)) + ((g388) & (g389) & (g390) & (g391) & (g60) & (!g61)) + ((g388) & (g389) & (g390) & (g391) & (g60) & (g61)));
	assign g397 = (((!g393) & (!g394) & (!g395) & (g396) & (g60) & (g61)) + ((!g393) & (!g394) & (g395) & (!g396) & (!g60) & (g61)) + ((!g393) & (!g394) & (g395) & (g396) & (!g60) & (g61)) + ((!g393) & (!g394) & (g395) & (g396) & (g60) & (g61)) + ((!g393) & (g394) & (!g395) & (!g396) & (g60) & (!g61)) + ((!g393) & (g394) & (!g395) & (g396) & (g60) & (!g61)) + ((!g393) & (g394) & (!g395) & (g396) & (g60) & (g61)) + ((!g393) & (g394) & (g395) & (!g396) & (!g60) & (g61)) + ((!g393) & (g394) & (g395) & (!g396) & (g60) & (!g61)) + ((!g393) & (g394) & (g395) & (g396) & (!g60) & (g61)) + ((!g393) & (g394) & (g395) & (g396) & (g60) & (!g61)) + ((!g393) & (g394) & (g395) & (g396) & (g60) & (g61)) + ((g393) & (!g394) & (!g395) & (!g396) & (!g60) & (!g61)) + ((g393) & (!g394) & (!g395) & (g396) & (!g60) & (!g61)) + ((g393) & (!g394) & (!g395) & (g396) & (g60) & (g61)) + ((g393) & (!g394) & (g395) & (!g396) & (!g60) & (!g61)) + ((g393) & (!g394) & (g395) & (!g396) & (!g60) & (g61)) + ((g393) & (!g394) & (g395) & (g396) & (!g60) & (!g61)) + ((g393) & (!g394) & (g395) & (g396) & (!g60) & (g61)) + ((g393) & (!g394) & (g395) & (g396) & (g60) & (g61)) + ((g393) & (g394) & (!g395) & (!g396) & (!g60) & (!g61)) + ((g393) & (g394) & (!g395) & (!g396) & (g60) & (!g61)) + ((g393) & (g394) & (!g395) & (g396) & (!g60) & (!g61)) + ((g393) & (g394) & (!g395) & (g396) & (g60) & (!g61)) + ((g393) & (g394) & (!g395) & (g396) & (g60) & (g61)) + ((g393) & (g394) & (g395) & (!g396) & (!g60) & (!g61)) + ((g393) & (g394) & (g395) & (!g396) & (!g60) & (g61)) + ((g393) & (g394) & (g395) & (!g396) & (g60) & (!g61)) + ((g393) & (g394) & (g395) & (g396) & (!g60) & (!g61)) + ((g393) & (g394) & (g395) & (g396) & (!g60) & (g61)) + ((g393) & (g394) & (g395) & (g396) & (g60) & (!g61)) + ((g393) & (g394) & (g395) & (g396) & (g60) & (g61)));
	assign g402 = (((!g398) & (!g399) & (!g400) & (g401) & (g60) & (g61)) + ((!g398) & (!g399) & (g400) & (!g401) & (!g60) & (g61)) + ((!g398) & (!g399) & (g400) & (g401) & (!g60) & (g61)) + ((!g398) & (!g399) & (g400) & (g401) & (g60) & (g61)) + ((!g398) & (g399) & (!g400) & (!g401) & (g60) & (!g61)) + ((!g398) & (g399) & (!g400) & (g401) & (g60) & (!g61)) + ((!g398) & (g399) & (!g400) & (g401) & (g60) & (g61)) + ((!g398) & (g399) & (g400) & (!g401) & (!g60) & (g61)) + ((!g398) & (g399) & (g400) & (!g401) & (g60) & (!g61)) + ((!g398) & (g399) & (g400) & (g401) & (!g60) & (g61)) + ((!g398) & (g399) & (g400) & (g401) & (g60) & (!g61)) + ((!g398) & (g399) & (g400) & (g401) & (g60) & (g61)) + ((g398) & (!g399) & (!g400) & (!g401) & (!g60) & (!g61)) + ((g398) & (!g399) & (!g400) & (g401) & (!g60) & (!g61)) + ((g398) & (!g399) & (!g400) & (g401) & (g60) & (g61)) + ((g398) & (!g399) & (g400) & (!g401) & (!g60) & (!g61)) + ((g398) & (!g399) & (g400) & (!g401) & (!g60) & (g61)) + ((g398) & (!g399) & (g400) & (g401) & (!g60) & (!g61)) + ((g398) & (!g399) & (g400) & (g401) & (!g60) & (g61)) + ((g398) & (!g399) & (g400) & (g401) & (g60) & (g61)) + ((g398) & (g399) & (!g400) & (!g401) & (!g60) & (!g61)) + ((g398) & (g399) & (!g400) & (!g401) & (g60) & (!g61)) + ((g398) & (g399) & (!g400) & (g401) & (!g60) & (!g61)) + ((g398) & (g399) & (!g400) & (g401) & (g60) & (!g61)) + ((g398) & (g399) & (!g400) & (g401) & (g60) & (g61)) + ((g398) & (g399) & (g400) & (!g401) & (!g60) & (!g61)) + ((g398) & (g399) & (g400) & (!g401) & (!g60) & (g61)) + ((g398) & (g399) & (g400) & (!g401) & (g60) & (!g61)) + ((g398) & (g399) & (g400) & (g401) & (!g60) & (!g61)) + ((g398) & (g399) & (g400) & (g401) & (!g60) & (g61)) + ((g398) & (g399) & (g400) & (g401) & (g60) & (!g61)) + ((g398) & (g399) & (g400) & (g401) & (g60) & (g61)));
	assign g407 = (((!g403) & (!g404) & (!g405) & (g406) & (g60) & (g61)) + ((!g403) & (!g404) & (g405) & (!g406) & (!g60) & (g61)) + ((!g403) & (!g404) & (g405) & (g406) & (!g60) & (g61)) + ((!g403) & (!g404) & (g405) & (g406) & (g60) & (g61)) + ((!g403) & (g404) & (!g405) & (!g406) & (g60) & (!g61)) + ((!g403) & (g404) & (!g405) & (g406) & (g60) & (!g61)) + ((!g403) & (g404) & (!g405) & (g406) & (g60) & (g61)) + ((!g403) & (g404) & (g405) & (!g406) & (!g60) & (g61)) + ((!g403) & (g404) & (g405) & (!g406) & (g60) & (!g61)) + ((!g403) & (g404) & (g405) & (g406) & (!g60) & (g61)) + ((!g403) & (g404) & (g405) & (g406) & (g60) & (!g61)) + ((!g403) & (g404) & (g405) & (g406) & (g60) & (g61)) + ((g403) & (!g404) & (!g405) & (!g406) & (!g60) & (!g61)) + ((g403) & (!g404) & (!g405) & (g406) & (!g60) & (!g61)) + ((g403) & (!g404) & (!g405) & (g406) & (g60) & (g61)) + ((g403) & (!g404) & (g405) & (!g406) & (!g60) & (!g61)) + ((g403) & (!g404) & (g405) & (!g406) & (!g60) & (g61)) + ((g403) & (!g404) & (g405) & (g406) & (!g60) & (!g61)) + ((g403) & (!g404) & (g405) & (g406) & (!g60) & (g61)) + ((g403) & (!g404) & (g405) & (g406) & (g60) & (g61)) + ((g403) & (g404) & (!g405) & (!g406) & (!g60) & (!g61)) + ((g403) & (g404) & (!g405) & (!g406) & (g60) & (!g61)) + ((g403) & (g404) & (!g405) & (g406) & (!g60) & (!g61)) + ((g403) & (g404) & (!g405) & (g406) & (g60) & (!g61)) + ((g403) & (g404) & (!g405) & (g406) & (g60) & (g61)) + ((g403) & (g404) & (g405) & (!g406) & (!g60) & (!g61)) + ((g403) & (g404) & (g405) & (!g406) & (!g60) & (g61)) + ((g403) & (g404) & (g405) & (!g406) & (g60) & (!g61)) + ((g403) & (g404) & (g405) & (g406) & (!g60) & (!g61)) + ((g403) & (g404) & (g405) & (g406) & (!g60) & (g61)) + ((g403) & (g404) & (g405) & (g406) & (g60) & (!g61)) + ((g403) & (g404) & (g405) & (g406) & (g60) & (g61)));
	assign g408 = (((!g392) & (!g397) & (!g402) & (g407) & (g42) & (g43)) + ((!g392) & (!g397) & (g402) & (!g407) & (!g42) & (g43)) + ((!g392) & (!g397) & (g402) & (g407) & (!g42) & (g43)) + ((!g392) & (!g397) & (g402) & (g407) & (g42) & (g43)) + ((!g392) & (g397) & (!g402) & (!g407) & (g42) & (!g43)) + ((!g392) & (g397) & (!g402) & (g407) & (g42) & (!g43)) + ((!g392) & (g397) & (!g402) & (g407) & (g42) & (g43)) + ((!g392) & (g397) & (g402) & (!g407) & (!g42) & (g43)) + ((!g392) & (g397) & (g402) & (!g407) & (g42) & (!g43)) + ((!g392) & (g397) & (g402) & (g407) & (!g42) & (g43)) + ((!g392) & (g397) & (g402) & (g407) & (g42) & (!g43)) + ((!g392) & (g397) & (g402) & (g407) & (g42) & (g43)) + ((g392) & (!g397) & (!g402) & (!g407) & (!g42) & (!g43)) + ((g392) & (!g397) & (!g402) & (g407) & (!g42) & (!g43)) + ((g392) & (!g397) & (!g402) & (g407) & (g42) & (g43)) + ((g392) & (!g397) & (g402) & (!g407) & (!g42) & (!g43)) + ((g392) & (!g397) & (g402) & (!g407) & (!g42) & (g43)) + ((g392) & (!g397) & (g402) & (g407) & (!g42) & (!g43)) + ((g392) & (!g397) & (g402) & (g407) & (!g42) & (g43)) + ((g392) & (!g397) & (g402) & (g407) & (g42) & (g43)) + ((g392) & (g397) & (!g402) & (!g407) & (!g42) & (!g43)) + ((g392) & (g397) & (!g402) & (!g407) & (g42) & (!g43)) + ((g392) & (g397) & (!g402) & (g407) & (!g42) & (!g43)) + ((g392) & (g397) & (!g402) & (g407) & (g42) & (!g43)) + ((g392) & (g397) & (!g402) & (g407) & (g42) & (g43)) + ((g392) & (g397) & (g402) & (!g407) & (!g42) & (!g43)) + ((g392) & (g397) & (g402) & (!g407) & (!g42) & (g43)) + ((g392) & (g397) & (g402) & (!g407) & (g42) & (!g43)) + ((g392) & (g397) & (g402) & (g407) & (!g42) & (!g43)) + ((g392) & (g397) & (g402) & (g407) & (!g42) & (g43)) + ((g392) & (g397) & (g402) & (g407) & (g42) & (!g43)) + ((g392) & (g397) & (g402) & (g407) & (g42) & (g43)));
	assign g7249 = (((!g832) & (g1338) & (!g409)) + ((!g832) & (g1338) & (g409)) + ((g832) & (!g1338) & (g409)) + ((g832) & (g1338) & (g409)));
	assign g410 = (((!g34) & (!reset) & (!g408) & (g409)) + ((!g34) & (!reset) & (g408) & (g409)) + ((g34) & (!reset) & (g408) & (!g409)) + ((g34) & (!reset) & (g408) & (g409)));
	assign g415 = (((!g411) & (!g412) & (!g413) & (g414) & (g42) & (g43)) + ((!g411) & (!g412) & (g413) & (!g414) & (!g42) & (g43)) + ((!g411) & (!g412) & (g413) & (g414) & (!g42) & (g43)) + ((!g411) & (!g412) & (g413) & (g414) & (g42) & (g43)) + ((!g411) & (g412) & (!g413) & (!g414) & (g42) & (!g43)) + ((!g411) & (g412) & (!g413) & (g414) & (g42) & (!g43)) + ((!g411) & (g412) & (!g413) & (g414) & (g42) & (g43)) + ((!g411) & (g412) & (g413) & (!g414) & (!g42) & (g43)) + ((!g411) & (g412) & (g413) & (!g414) & (g42) & (!g43)) + ((!g411) & (g412) & (g413) & (g414) & (!g42) & (g43)) + ((!g411) & (g412) & (g413) & (g414) & (g42) & (!g43)) + ((!g411) & (g412) & (g413) & (g414) & (g42) & (g43)) + ((g411) & (!g412) & (!g413) & (!g414) & (!g42) & (!g43)) + ((g411) & (!g412) & (!g413) & (g414) & (!g42) & (!g43)) + ((g411) & (!g412) & (!g413) & (g414) & (g42) & (g43)) + ((g411) & (!g412) & (g413) & (!g414) & (!g42) & (!g43)) + ((g411) & (!g412) & (g413) & (!g414) & (!g42) & (g43)) + ((g411) & (!g412) & (g413) & (g414) & (!g42) & (!g43)) + ((g411) & (!g412) & (g413) & (g414) & (!g42) & (g43)) + ((g411) & (!g412) & (g413) & (g414) & (g42) & (g43)) + ((g411) & (g412) & (!g413) & (!g414) & (!g42) & (!g43)) + ((g411) & (g412) & (!g413) & (!g414) & (g42) & (!g43)) + ((g411) & (g412) & (!g413) & (g414) & (!g42) & (!g43)) + ((g411) & (g412) & (!g413) & (g414) & (g42) & (!g43)) + ((g411) & (g412) & (!g413) & (g414) & (g42) & (g43)) + ((g411) & (g412) & (g413) & (!g414) & (!g42) & (!g43)) + ((g411) & (g412) & (g413) & (!g414) & (!g42) & (g43)) + ((g411) & (g412) & (g413) & (!g414) & (g42) & (!g43)) + ((g411) & (g412) & (g413) & (g414) & (!g42) & (!g43)) + ((g411) & (g412) & (g413) & (g414) & (!g42) & (g43)) + ((g411) & (g412) & (g413) & (g414) & (g42) & (!g43)) + ((g411) & (g412) & (g413) & (g414) & (g42) & (g43)));
	assign g420 = (((!g416) & (!g417) & (!g418) & (g419) & (g42) & (g43)) + ((!g416) & (!g417) & (g418) & (!g419) & (!g42) & (g43)) + ((!g416) & (!g417) & (g418) & (g419) & (!g42) & (g43)) + ((!g416) & (!g417) & (g418) & (g419) & (g42) & (g43)) + ((!g416) & (g417) & (!g418) & (!g419) & (g42) & (!g43)) + ((!g416) & (g417) & (!g418) & (g419) & (g42) & (!g43)) + ((!g416) & (g417) & (!g418) & (g419) & (g42) & (g43)) + ((!g416) & (g417) & (g418) & (!g419) & (!g42) & (g43)) + ((!g416) & (g417) & (g418) & (!g419) & (g42) & (!g43)) + ((!g416) & (g417) & (g418) & (g419) & (!g42) & (g43)) + ((!g416) & (g417) & (g418) & (g419) & (g42) & (!g43)) + ((!g416) & (g417) & (g418) & (g419) & (g42) & (g43)) + ((g416) & (!g417) & (!g418) & (!g419) & (!g42) & (!g43)) + ((g416) & (!g417) & (!g418) & (g419) & (!g42) & (!g43)) + ((g416) & (!g417) & (!g418) & (g419) & (g42) & (g43)) + ((g416) & (!g417) & (g418) & (!g419) & (!g42) & (!g43)) + ((g416) & (!g417) & (g418) & (!g419) & (!g42) & (g43)) + ((g416) & (!g417) & (g418) & (g419) & (!g42) & (!g43)) + ((g416) & (!g417) & (g418) & (g419) & (!g42) & (g43)) + ((g416) & (!g417) & (g418) & (g419) & (g42) & (g43)) + ((g416) & (g417) & (!g418) & (!g419) & (!g42) & (!g43)) + ((g416) & (g417) & (!g418) & (!g419) & (g42) & (!g43)) + ((g416) & (g417) & (!g418) & (g419) & (!g42) & (!g43)) + ((g416) & (g417) & (!g418) & (g419) & (g42) & (!g43)) + ((g416) & (g417) & (!g418) & (g419) & (g42) & (g43)) + ((g416) & (g417) & (g418) & (!g419) & (!g42) & (!g43)) + ((g416) & (g417) & (g418) & (!g419) & (!g42) & (g43)) + ((g416) & (g417) & (g418) & (!g419) & (g42) & (!g43)) + ((g416) & (g417) & (g418) & (g419) & (!g42) & (!g43)) + ((g416) & (g417) & (g418) & (g419) & (!g42) & (g43)) + ((g416) & (g417) & (g418) & (g419) & (g42) & (!g43)) + ((g416) & (g417) & (g418) & (g419) & (g42) & (g43)));
	assign g425 = (((!g421) & (!g422) & (!g423) & (g424) & (g42) & (g43)) + ((!g421) & (!g422) & (g423) & (!g424) & (!g42) & (g43)) + ((!g421) & (!g422) & (g423) & (g424) & (!g42) & (g43)) + ((!g421) & (!g422) & (g423) & (g424) & (g42) & (g43)) + ((!g421) & (g422) & (!g423) & (!g424) & (g42) & (!g43)) + ((!g421) & (g422) & (!g423) & (g424) & (g42) & (!g43)) + ((!g421) & (g422) & (!g423) & (g424) & (g42) & (g43)) + ((!g421) & (g422) & (g423) & (!g424) & (!g42) & (g43)) + ((!g421) & (g422) & (g423) & (!g424) & (g42) & (!g43)) + ((!g421) & (g422) & (g423) & (g424) & (!g42) & (g43)) + ((!g421) & (g422) & (g423) & (g424) & (g42) & (!g43)) + ((!g421) & (g422) & (g423) & (g424) & (g42) & (g43)) + ((g421) & (!g422) & (!g423) & (!g424) & (!g42) & (!g43)) + ((g421) & (!g422) & (!g423) & (g424) & (!g42) & (!g43)) + ((g421) & (!g422) & (!g423) & (g424) & (g42) & (g43)) + ((g421) & (!g422) & (g423) & (!g424) & (!g42) & (!g43)) + ((g421) & (!g422) & (g423) & (!g424) & (!g42) & (g43)) + ((g421) & (!g422) & (g423) & (g424) & (!g42) & (!g43)) + ((g421) & (!g422) & (g423) & (g424) & (!g42) & (g43)) + ((g421) & (!g422) & (g423) & (g424) & (g42) & (g43)) + ((g421) & (g422) & (!g423) & (!g424) & (!g42) & (!g43)) + ((g421) & (g422) & (!g423) & (!g424) & (g42) & (!g43)) + ((g421) & (g422) & (!g423) & (g424) & (!g42) & (!g43)) + ((g421) & (g422) & (!g423) & (g424) & (g42) & (!g43)) + ((g421) & (g422) & (!g423) & (g424) & (g42) & (g43)) + ((g421) & (g422) & (g423) & (!g424) & (!g42) & (!g43)) + ((g421) & (g422) & (g423) & (!g424) & (!g42) & (g43)) + ((g421) & (g422) & (g423) & (!g424) & (g42) & (!g43)) + ((g421) & (g422) & (g423) & (g424) & (!g42) & (!g43)) + ((g421) & (g422) & (g423) & (g424) & (!g42) & (g43)) + ((g421) & (g422) & (g423) & (g424) & (g42) & (!g43)) + ((g421) & (g422) & (g423) & (g424) & (g42) & (g43)));
	assign g430 = (((!g426) & (!g427) & (!g428) & (g429) & (g42) & (g43)) + ((!g426) & (!g427) & (g428) & (!g429) & (!g42) & (g43)) + ((!g426) & (!g427) & (g428) & (g429) & (!g42) & (g43)) + ((!g426) & (!g427) & (g428) & (g429) & (g42) & (g43)) + ((!g426) & (g427) & (!g428) & (!g429) & (g42) & (!g43)) + ((!g426) & (g427) & (!g428) & (g429) & (g42) & (!g43)) + ((!g426) & (g427) & (!g428) & (g429) & (g42) & (g43)) + ((!g426) & (g427) & (g428) & (!g429) & (!g42) & (g43)) + ((!g426) & (g427) & (g428) & (!g429) & (g42) & (!g43)) + ((!g426) & (g427) & (g428) & (g429) & (!g42) & (g43)) + ((!g426) & (g427) & (g428) & (g429) & (g42) & (!g43)) + ((!g426) & (g427) & (g428) & (g429) & (g42) & (g43)) + ((g426) & (!g427) & (!g428) & (!g429) & (!g42) & (!g43)) + ((g426) & (!g427) & (!g428) & (g429) & (!g42) & (!g43)) + ((g426) & (!g427) & (!g428) & (g429) & (g42) & (g43)) + ((g426) & (!g427) & (g428) & (!g429) & (!g42) & (!g43)) + ((g426) & (!g427) & (g428) & (!g429) & (!g42) & (g43)) + ((g426) & (!g427) & (g428) & (g429) & (!g42) & (!g43)) + ((g426) & (!g427) & (g428) & (g429) & (!g42) & (g43)) + ((g426) & (!g427) & (g428) & (g429) & (g42) & (g43)) + ((g426) & (g427) & (!g428) & (!g429) & (!g42) & (!g43)) + ((g426) & (g427) & (!g428) & (!g429) & (g42) & (!g43)) + ((g426) & (g427) & (!g428) & (g429) & (!g42) & (!g43)) + ((g426) & (g427) & (!g428) & (g429) & (g42) & (!g43)) + ((g426) & (g427) & (!g428) & (g429) & (g42) & (g43)) + ((g426) & (g427) & (g428) & (!g429) & (!g42) & (!g43)) + ((g426) & (g427) & (g428) & (!g429) & (!g42) & (g43)) + ((g426) & (g427) & (g428) & (!g429) & (g42) & (!g43)) + ((g426) & (g427) & (g428) & (g429) & (!g42) & (!g43)) + ((g426) & (g427) & (g428) & (g429) & (!g42) & (g43)) + ((g426) & (g427) & (g428) & (g429) & (g42) & (!g43)) + ((g426) & (g427) & (g428) & (g429) & (g42) & (g43)));
	assign g431 = (((!g415) & (!g420) & (!g425) & (g430) & (g60) & (g61)) + ((!g415) & (!g420) & (g425) & (!g430) & (!g60) & (g61)) + ((!g415) & (!g420) & (g425) & (g430) & (!g60) & (g61)) + ((!g415) & (!g420) & (g425) & (g430) & (g60) & (g61)) + ((!g415) & (g420) & (!g425) & (!g430) & (g60) & (!g61)) + ((!g415) & (g420) & (!g425) & (g430) & (g60) & (!g61)) + ((!g415) & (g420) & (!g425) & (g430) & (g60) & (g61)) + ((!g415) & (g420) & (g425) & (!g430) & (!g60) & (g61)) + ((!g415) & (g420) & (g425) & (!g430) & (g60) & (!g61)) + ((!g415) & (g420) & (g425) & (g430) & (!g60) & (g61)) + ((!g415) & (g420) & (g425) & (g430) & (g60) & (!g61)) + ((!g415) & (g420) & (g425) & (g430) & (g60) & (g61)) + ((g415) & (!g420) & (!g425) & (!g430) & (!g60) & (!g61)) + ((g415) & (!g420) & (!g425) & (g430) & (!g60) & (!g61)) + ((g415) & (!g420) & (!g425) & (g430) & (g60) & (g61)) + ((g415) & (!g420) & (g425) & (!g430) & (!g60) & (!g61)) + ((g415) & (!g420) & (g425) & (!g430) & (!g60) & (g61)) + ((g415) & (!g420) & (g425) & (g430) & (!g60) & (!g61)) + ((g415) & (!g420) & (g425) & (g430) & (!g60) & (g61)) + ((g415) & (!g420) & (g425) & (g430) & (g60) & (g61)) + ((g415) & (g420) & (!g425) & (!g430) & (!g60) & (!g61)) + ((g415) & (g420) & (!g425) & (!g430) & (g60) & (!g61)) + ((g415) & (g420) & (!g425) & (g430) & (!g60) & (!g61)) + ((g415) & (g420) & (!g425) & (g430) & (g60) & (!g61)) + ((g415) & (g420) & (!g425) & (g430) & (g60) & (g61)) + ((g415) & (g420) & (g425) & (!g430) & (!g60) & (!g61)) + ((g415) & (g420) & (g425) & (!g430) & (!g60) & (g61)) + ((g415) & (g420) & (g425) & (!g430) & (g60) & (!g61)) + ((g415) & (g420) & (g425) & (g430) & (!g60) & (!g61)) + ((g415) & (g420) & (g425) & (g430) & (!g60) & (g61)) + ((g415) & (g420) & (g425) & (g430) & (g60) & (!g61)) + ((g415) & (g420) & (g425) & (g430) & (g60) & (g61)));
	assign g7250 = (((!g832) & (g1374) & (!g432)) + ((!g832) & (g1374) & (g432)) + ((g832) & (!g1374) & (g432)) + ((g832) & (g1374) & (g432)));
	assign g433 = (((!g34) & (!reset) & (!g431) & (g432)) + ((!g34) & (!reset) & (g431) & (g432)) + ((g34) & (!reset) & (g431) & (!g432)) + ((g34) & (!reset) & (g431) & (g432)));
	assign g438 = (((!g434) & (!g435) & (!g436) & (g437) & (g60) & (g61)) + ((!g434) & (!g435) & (g436) & (!g437) & (!g60) & (g61)) + ((!g434) & (!g435) & (g436) & (g437) & (!g60) & (g61)) + ((!g434) & (!g435) & (g436) & (g437) & (g60) & (g61)) + ((!g434) & (g435) & (!g436) & (!g437) & (g60) & (!g61)) + ((!g434) & (g435) & (!g436) & (g437) & (g60) & (!g61)) + ((!g434) & (g435) & (!g436) & (g437) & (g60) & (g61)) + ((!g434) & (g435) & (g436) & (!g437) & (!g60) & (g61)) + ((!g434) & (g435) & (g436) & (!g437) & (g60) & (!g61)) + ((!g434) & (g435) & (g436) & (g437) & (!g60) & (g61)) + ((!g434) & (g435) & (g436) & (g437) & (g60) & (!g61)) + ((!g434) & (g435) & (g436) & (g437) & (g60) & (g61)) + ((g434) & (!g435) & (!g436) & (!g437) & (!g60) & (!g61)) + ((g434) & (!g435) & (!g436) & (g437) & (!g60) & (!g61)) + ((g434) & (!g435) & (!g436) & (g437) & (g60) & (g61)) + ((g434) & (!g435) & (g436) & (!g437) & (!g60) & (!g61)) + ((g434) & (!g435) & (g436) & (!g437) & (!g60) & (g61)) + ((g434) & (!g435) & (g436) & (g437) & (!g60) & (!g61)) + ((g434) & (!g435) & (g436) & (g437) & (!g60) & (g61)) + ((g434) & (!g435) & (g436) & (g437) & (g60) & (g61)) + ((g434) & (g435) & (!g436) & (!g437) & (!g60) & (!g61)) + ((g434) & (g435) & (!g436) & (!g437) & (g60) & (!g61)) + ((g434) & (g435) & (!g436) & (g437) & (!g60) & (!g61)) + ((g434) & (g435) & (!g436) & (g437) & (g60) & (!g61)) + ((g434) & (g435) & (!g436) & (g437) & (g60) & (g61)) + ((g434) & (g435) & (g436) & (!g437) & (!g60) & (!g61)) + ((g434) & (g435) & (g436) & (!g437) & (!g60) & (g61)) + ((g434) & (g435) & (g436) & (!g437) & (g60) & (!g61)) + ((g434) & (g435) & (g436) & (g437) & (!g60) & (!g61)) + ((g434) & (g435) & (g436) & (g437) & (!g60) & (g61)) + ((g434) & (g435) & (g436) & (g437) & (g60) & (!g61)) + ((g434) & (g435) & (g436) & (g437) & (g60) & (g61)));
	assign g443 = (((!g439) & (!g440) & (!g441) & (g442) & (g60) & (g61)) + ((!g439) & (!g440) & (g441) & (!g442) & (!g60) & (g61)) + ((!g439) & (!g440) & (g441) & (g442) & (!g60) & (g61)) + ((!g439) & (!g440) & (g441) & (g442) & (g60) & (g61)) + ((!g439) & (g440) & (!g441) & (!g442) & (g60) & (!g61)) + ((!g439) & (g440) & (!g441) & (g442) & (g60) & (!g61)) + ((!g439) & (g440) & (!g441) & (g442) & (g60) & (g61)) + ((!g439) & (g440) & (g441) & (!g442) & (!g60) & (g61)) + ((!g439) & (g440) & (g441) & (!g442) & (g60) & (!g61)) + ((!g439) & (g440) & (g441) & (g442) & (!g60) & (g61)) + ((!g439) & (g440) & (g441) & (g442) & (g60) & (!g61)) + ((!g439) & (g440) & (g441) & (g442) & (g60) & (g61)) + ((g439) & (!g440) & (!g441) & (!g442) & (!g60) & (!g61)) + ((g439) & (!g440) & (!g441) & (g442) & (!g60) & (!g61)) + ((g439) & (!g440) & (!g441) & (g442) & (g60) & (g61)) + ((g439) & (!g440) & (g441) & (!g442) & (!g60) & (!g61)) + ((g439) & (!g440) & (g441) & (!g442) & (!g60) & (g61)) + ((g439) & (!g440) & (g441) & (g442) & (!g60) & (!g61)) + ((g439) & (!g440) & (g441) & (g442) & (!g60) & (g61)) + ((g439) & (!g440) & (g441) & (g442) & (g60) & (g61)) + ((g439) & (g440) & (!g441) & (!g442) & (!g60) & (!g61)) + ((g439) & (g440) & (!g441) & (!g442) & (g60) & (!g61)) + ((g439) & (g440) & (!g441) & (g442) & (!g60) & (!g61)) + ((g439) & (g440) & (!g441) & (g442) & (g60) & (!g61)) + ((g439) & (g440) & (!g441) & (g442) & (g60) & (g61)) + ((g439) & (g440) & (g441) & (!g442) & (!g60) & (!g61)) + ((g439) & (g440) & (g441) & (!g442) & (!g60) & (g61)) + ((g439) & (g440) & (g441) & (!g442) & (g60) & (!g61)) + ((g439) & (g440) & (g441) & (g442) & (!g60) & (!g61)) + ((g439) & (g440) & (g441) & (g442) & (!g60) & (g61)) + ((g439) & (g440) & (g441) & (g442) & (g60) & (!g61)) + ((g439) & (g440) & (g441) & (g442) & (g60) & (g61)));
	assign g448 = (((!g444) & (!g445) & (!g446) & (g447) & (g60) & (g61)) + ((!g444) & (!g445) & (g446) & (!g447) & (!g60) & (g61)) + ((!g444) & (!g445) & (g446) & (g447) & (!g60) & (g61)) + ((!g444) & (!g445) & (g446) & (g447) & (g60) & (g61)) + ((!g444) & (g445) & (!g446) & (!g447) & (g60) & (!g61)) + ((!g444) & (g445) & (!g446) & (g447) & (g60) & (!g61)) + ((!g444) & (g445) & (!g446) & (g447) & (g60) & (g61)) + ((!g444) & (g445) & (g446) & (!g447) & (!g60) & (g61)) + ((!g444) & (g445) & (g446) & (!g447) & (g60) & (!g61)) + ((!g444) & (g445) & (g446) & (g447) & (!g60) & (g61)) + ((!g444) & (g445) & (g446) & (g447) & (g60) & (!g61)) + ((!g444) & (g445) & (g446) & (g447) & (g60) & (g61)) + ((g444) & (!g445) & (!g446) & (!g447) & (!g60) & (!g61)) + ((g444) & (!g445) & (!g446) & (g447) & (!g60) & (!g61)) + ((g444) & (!g445) & (!g446) & (g447) & (g60) & (g61)) + ((g444) & (!g445) & (g446) & (!g447) & (!g60) & (!g61)) + ((g444) & (!g445) & (g446) & (!g447) & (!g60) & (g61)) + ((g444) & (!g445) & (g446) & (g447) & (!g60) & (!g61)) + ((g444) & (!g445) & (g446) & (g447) & (!g60) & (g61)) + ((g444) & (!g445) & (g446) & (g447) & (g60) & (g61)) + ((g444) & (g445) & (!g446) & (!g447) & (!g60) & (!g61)) + ((g444) & (g445) & (!g446) & (!g447) & (g60) & (!g61)) + ((g444) & (g445) & (!g446) & (g447) & (!g60) & (!g61)) + ((g444) & (g445) & (!g446) & (g447) & (g60) & (!g61)) + ((g444) & (g445) & (!g446) & (g447) & (g60) & (g61)) + ((g444) & (g445) & (g446) & (!g447) & (!g60) & (!g61)) + ((g444) & (g445) & (g446) & (!g447) & (!g60) & (g61)) + ((g444) & (g445) & (g446) & (!g447) & (g60) & (!g61)) + ((g444) & (g445) & (g446) & (g447) & (!g60) & (!g61)) + ((g444) & (g445) & (g446) & (g447) & (!g60) & (g61)) + ((g444) & (g445) & (g446) & (g447) & (g60) & (!g61)) + ((g444) & (g445) & (g446) & (g447) & (g60) & (g61)));
	assign g453 = (((!g449) & (!g450) & (!g451) & (g452) & (g60) & (g61)) + ((!g449) & (!g450) & (g451) & (!g452) & (!g60) & (g61)) + ((!g449) & (!g450) & (g451) & (g452) & (!g60) & (g61)) + ((!g449) & (!g450) & (g451) & (g452) & (g60) & (g61)) + ((!g449) & (g450) & (!g451) & (!g452) & (g60) & (!g61)) + ((!g449) & (g450) & (!g451) & (g452) & (g60) & (!g61)) + ((!g449) & (g450) & (!g451) & (g452) & (g60) & (g61)) + ((!g449) & (g450) & (g451) & (!g452) & (!g60) & (g61)) + ((!g449) & (g450) & (g451) & (!g452) & (g60) & (!g61)) + ((!g449) & (g450) & (g451) & (g452) & (!g60) & (g61)) + ((!g449) & (g450) & (g451) & (g452) & (g60) & (!g61)) + ((!g449) & (g450) & (g451) & (g452) & (g60) & (g61)) + ((g449) & (!g450) & (!g451) & (!g452) & (!g60) & (!g61)) + ((g449) & (!g450) & (!g451) & (g452) & (!g60) & (!g61)) + ((g449) & (!g450) & (!g451) & (g452) & (g60) & (g61)) + ((g449) & (!g450) & (g451) & (!g452) & (!g60) & (!g61)) + ((g449) & (!g450) & (g451) & (!g452) & (!g60) & (g61)) + ((g449) & (!g450) & (g451) & (g452) & (!g60) & (!g61)) + ((g449) & (!g450) & (g451) & (g452) & (!g60) & (g61)) + ((g449) & (!g450) & (g451) & (g452) & (g60) & (g61)) + ((g449) & (g450) & (!g451) & (!g452) & (!g60) & (!g61)) + ((g449) & (g450) & (!g451) & (!g452) & (g60) & (!g61)) + ((g449) & (g450) & (!g451) & (g452) & (!g60) & (!g61)) + ((g449) & (g450) & (!g451) & (g452) & (g60) & (!g61)) + ((g449) & (g450) & (!g451) & (g452) & (g60) & (g61)) + ((g449) & (g450) & (g451) & (!g452) & (!g60) & (!g61)) + ((g449) & (g450) & (g451) & (!g452) & (!g60) & (g61)) + ((g449) & (g450) & (g451) & (!g452) & (g60) & (!g61)) + ((g449) & (g450) & (g451) & (g452) & (!g60) & (!g61)) + ((g449) & (g450) & (g451) & (g452) & (!g60) & (g61)) + ((g449) & (g450) & (g451) & (g452) & (g60) & (!g61)) + ((g449) & (g450) & (g451) & (g452) & (g60) & (g61)));
	assign g454 = (((!g438) & (!g443) & (!g448) & (g453) & (g42) & (g43)) + ((!g438) & (!g443) & (g448) & (!g453) & (!g42) & (g43)) + ((!g438) & (!g443) & (g448) & (g453) & (!g42) & (g43)) + ((!g438) & (!g443) & (g448) & (g453) & (g42) & (g43)) + ((!g438) & (g443) & (!g448) & (!g453) & (g42) & (!g43)) + ((!g438) & (g443) & (!g448) & (g453) & (g42) & (!g43)) + ((!g438) & (g443) & (!g448) & (g453) & (g42) & (g43)) + ((!g438) & (g443) & (g448) & (!g453) & (!g42) & (g43)) + ((!g438) & (g443) & (g448) & (!g453) & (g42) & (!g43)) + ((!g438) & (g443) & (g448) & (g453) & (!g42) & (g43)) + ((!g438) & (g443) & (g448) & (g453) & (g42) & (!g43)) + ((!g438) & (g443) & (g448) & (g453) & (g42) & (g43)) + ((g438) & (!g443) & (!g448) & (!g453) & (!g42) & (!g43)) + ((g438) & (!g443) & (!g448) & (g453) & (!g42) & (!g43)) + ((g438) & (!g443) & (!g448) & (g453) & (g42) & (g43)) + ((g438) & (!g443) & (g448) & (!g453) & (!g42) & (!g43)) + ((g438) & (!g443) & (g448) & (!g453) & (!g42) & (g43)) + ((g438) & (!g443) & (g448) & (g453) & (!g42) & (!g43)) + ((g438) & (!g443) & (g448) & (g453) & (!g42) & (g43)) + ((g438) & (!g443) & (g448) & (g453) & (g42) & (g43)) + ((g438) & (g443) & (!g448) & (!g453) & (!g42) & (!g43)) + ((g438) & (g443) & (!g448) & (!g453) & (g42) & (!g43)) + ((g438) & (g443) & (!g448) & (g453) & (!g42) & (!g43)) + ((g438) & (g443) & (!g448) & (g453) & (g42) & (!g43)) + ((g438) & (g443) & (!g448) & (g453) & (g42) & (g43)) + ((g438) & (g443) & (g448) & (!g453) & (!g42) & (!g43)) + ((g438) & (g443) & (g448) & (!g453) & (!g42) & (g43)) + ((g438) & (g443) & (g448) & (!g453) & (g42) & (!g43)) + ((g438) & (g443) & (g448) & (g453) & (!g42) & (!g43)) + ((g438) & (g443) & (g448) & (g453) & (!g42) & (g43)) + ((g438) & (g443) & (g448) & (g453) & (g42) & (!g43)) + ((g438) & (g443) & (g448) & (g453) & (g42) & (g43)));
	assign g7251 = (((!g832) & (g1407) & (!g455)) + ((!g832) & (g1407) & (g455)) + ((g832) & (!g1407) & (g455)) + ((g832) & (g1407) & (g455)));
	assign g456 = (((!g34) & (!reset) & (!g454) & (g455)) + ((!g34) & (!reset) & (g454) & (g455)) + ((g34) & (!reset) & (g454) & (!g455)) + ((g34) & (!reset) & (g454) & (g455)));
	assign g461 = (((!g457) & (!g458) & (!g459) & (g460) & (g42) & (g43)) + ((!g457) & (!g458) & (g459) & (!g460) & (!g42) & (g43)) + ((!g457) & (!g458) & (g459) & (g460) & (!g42) & (g43)) + ((!g457) & (!g458) & (g459) & (g460) & (g42) & (g43)) + ((!g457) & (g458) & (!g459) & (!g460) & (g42) & (!g43)) + ((!g457) & (g458) & (!g459) & (g460) & (g42) & (!g43)) + ((!g457) & (g458) & (!g459) & (g460) & (g42) & (g43)) + ((!g457) & (g458) & (g459) & (!g460) & (!g42) & (g43)) + ((!g457) & (g458) & (g459) & (!g460) & (g42) & (!g43)) + ((!g457) & (g458) & (g459) & (g460) & (!g42) & (g43)) + ((!g457) & (g458) & (g459) & (g460) & (g42) & (!g43)) + ((!g457) & (g458) & (g459) & (g460) & (g42) & (g43)) + ((g457) & (!g458) & (!g459) & (!g460) & (!g42) & (!g43)) + ((g457) & (!g458) & (!g459) & (g460) & (!g42) & (!g43)) + ((g457) & (!g458) & (!g459) & (g460) & (g42) & (g43)) + ((g457) & (!g458) & (g459) & (!g460) & (!g42) & (!g43)) + ((g457) & (!g458) & (g459) & (!g460) & (!g42) & (g43)) + ((g457) & (!g458) & (g459) & (g460) & (!g42) & (!g43)) + ((g457) & (!g458) & (g459) & (g460) & (!g42) & (g43)) + ((g457) & (!g458) & (g459) & (g460) & (g42) & (g43)) + ((g457) & (g458) & (!g459) & (!g460) & (!g42) & (!g43)) + ((g457) & (g458) & (!g459) & (!g460) & (g42) & (!g43)) + ((g457) & (g458) & (!g459) & (g460) & (!g42) & (!g43)) + ((g457) & (g458) & (!g459) & (g460) & (g42) & (!g43)) + ((g457) & (g458) & (!g459) & (g460) & (g42) & (g43)) + ((g457) & (g458) & (g459) & (!g460) & (!g42) & (!g43)) + ((g457) & (g458) & (g459) & (!g460) & (!g42) & (g43)) + ((g457) & (g458) & (g459) & (!g460) & (g42) & (!g43)) + ((g457) & (g458) & (g459) & (g460) & (!g42) & (!g43)) + ((g457) & (g458) & (g459) & (g460) & (!g42) & (g43)) + ((g457) & (g458) & (g459) & (g460) & (g42) & (!g43)) + ((g457) & (g458) & (g459) & (g460) & (g42) & (g43)));
	assign g466 = (((!g462) & (!g463) & (!g464) & (g465) & (g42) & (g43)) + ((!g462) & (!g463) & (g464) & (!g465) & (!g42) & (g43)) + ((!g462) & (!g463) & (g464) & (g465) & (!g42) & (g43)) + ((!g462) & (!g463) & (g464) & (g465) & (g42) & (g43)) + ((!g462) & (g463) & (!g464) & (!g465) & (g42) & (!g43)) + ((!g462) & (g463) & (!g464) & (g465) & (g42) & (!g43)) + ((!g462) & (g463) & (!g464) & (g465) & (g42) & (g43)) + ((!g462) & (g463) & (g464) & (!g465) & (!g42) & (g43)) + ((!g462) & (g463) & (g464) & (!g465) & (g42) & (!g43)) + ((!g462) & (g463) & (g464) & (g465) & (!g42) & (g43)) + ((!g462) & (g463) & (g464) & (g465) & (g42) & (!g43)) + ((!g462) & (g463) & (g464) & (g465) & (g42) & (g43)) + ((g462) & (!g463) & (!g464) & (!g465) & (!g42) & (!g43)) + ((g462) & (!g463) & (!g464) & (g465) & (!g42) & (!g43)) + ((g462) & (!g463) & (!g464) & (g465) & (g42) & (g43)) + ((g462) & (!g463) & (g464) & (!g465) & (!g42) & (!g43)) + ((g462) & (!g463) & (g464) & (!g465) & (!g42) & (g43)) + ((g462) & (!g463) & (g464) & (g465) & (!g42) & (!g43)) + ((g462) & (!g463) & (g464) & (g465) & (!g42) & (g43)) + ((g462) & (!g463) & (g464) & (g465) & (g42) & (g43)) + ((g462) & (g463) & (!g464) & (!g465) & (!g42) & (!g43)) + ((g462) & (g463) & (!g464) & (!g465) & (g42) & (!g43)) + ((g462) & (g463) & (!g464) & (g465) & (!g42) & (!g43)) + ((g462) & (g463) & (!g464) & (g465) & (g42) & (!g43)) + ((g462) & (g463) & (!g464) & (g465) & (g42) & (g43)) + ((g462) & (g463) & (g464) & (!g465) & (!g42) & (!g43)) + ((g462) & (g463) & (g464) & (!g465) & (!g42) & (g43)) + ((g462) & (g463) & (g464) & (!g465) & (g42) & (!g43)) + ((g462) & (g463) & (g464) & (g465) & (!g42) & (!g43)) + ((g462) & (g463) & (g464) & (g465) & (!g42) & (g43)) + ((g462) & (g463) & (g464) & (g465) & (g42) & (!g43)) + ((g462) & (g463) & (g464) & (g465) & (g42) & (g43)));
	assign g471 = (((!g467) & (!g468) & (!g469) & (g470) & (g42) & (g43)) + ((!g467) & (!g468) & (g469) & (!g470) & (!g42) & (g43)) + ((!g467) & (!g468) & (g469) & (g470) & (!g42) & (g43)) + ((!g467) & (!g468) & (g469) & (g470) & (g42) & (g43)) + ((!g467) & (g468) & (!g469) & (!g470) & (g42) & (!g43)) + ((!g467) & (g468) & (!g469) & (g470) & (g42) & (!g43)) + ((!g467) & (g468) & (!g469) & (g470) & (g42) & (g43)) + ((!g467) & (g468) & (g469) & (!g470) & (!g42) & (g43)) + ((!g467) & (g468) & (g469) & (!g470) & (g42) & (!g43)) + ((!g467) & (g468) & (g469) & (g470) & (!g42) & (g43)) + ((!g467) & (g468) & (g469) & (g470) & (g42) & (!g43)) + ((!g467) & (g468) & (g469) & (g470) & (g42) & (g43)) + ((g467) & (!g468) & (!g469) & (!g470) & (!g42) & (!g43)) + ((g467) & (!g468) & (!g469) & (g470) & (!g42) & (!g43)) + ((g467) & (!g468) & (!g469) & (g470) & (g42) & (g43)) + ((g467) & (!g468) & (g469) & (!g470) & (!g42) & (!g43)) + ((g467) & (!g468) & (g469) & (!g470) & (!g42) & (g43)) + ((g467) & (!g468) & (g469) & (g470) & (!g42) & (!g43)) + ((g467) & (!g468) & (g469) & (g470) & (!g42) & (g43)) + ((g467) & (!g468) & (g469) & (g470) & (g42) & (g43)) + ((g467) & (g468) & (!g469) & (!g470) & (!g42) & (!g43)) + ((g467) & (g468) & (!g469) & (!g470) & (g42) & (!g43)) + ((g467) & (g468) & (!g469) & (g470) & (!g42) & (!g43)) + ((g467) & (g468) & (!g469) & (g470) & (g42) & (!g43)) + ((g467) & (g468) & (!g469) & (g470) & (g42) & (g43)) + ((g467) & (g468) & (g469) & (!g470) & (!g42) & (!g43)) + ((g467) & (g468) & (g469) & (!g470) & (!g42) & (g43)) + ((g467) & (g468) & (g469) & (!g470) & (g42) & (!g43)) + ((g467) & (g468) & (g469) & (g470) & (!g42) & (!g43)) + ((g467) & (g468) & (g469) & (g470) & (!g42) & (g43)) + ((g467) & (g468) & (g469) & (g470) & (g42) & (!g43)) + ((g467) & (g468) & (g469) & (g470) & (g42) & (g43)));
	assign g476 = (((!g472) & (!g473) & (!g474) & (g475) & (g42) & (g43)) + ((!g472) & (!g473) & (g474) & (!g475) & (!g42) & (g43)) + ((!g472) & (!g473) & (g474) & (g475) & (!g42) & (g43)) + ((!g472) & (!g473) & (g474) & (g475) & (g42) & (g43)) + ((!g472) & (g473) & (!g474) & (!g475) & (g42) & (!g43)) + ((!g472) & (g473) & (!g474) & (g475) & (g42) & (!g43)) + ((!g472) & (g473) & (!g474) & (g475) & (g42) & (g43)) + ((!g472) & (g473) & (g474) & (!g475) & (!g42) & (g43)) + ((!g472) & (g473) & (g474) & (!g475) & (g42) & (!g43)) + ((!g472) & (g473) & (g474) & (g475) & (!g42) & (g43)) + ((!g472) & (g473) & (g474) & (g475) & (g42) & (!g43)) + ((!g472) & (g473) & (g474) & (g475) & (g42) & (g43)) + ((g472) & (!g473) & (!g474) & (!g475) & (!g42) & (!g43)) + ((g472) & (!g473) & (!g474) & (g475) & (!g42) & (!g43)) + ((g472) & (!g473) & (!g474) & (g475) & (g42) & (g43)) + ((g472) & (!g473) & (g474) & (!g475) & (!g42) & (!g43)) + ((g472) & (!g473) & (g474) & (!g475) & (!g42) & (g43)) + ((g472) & (!g473) & (g474) & (g475) & (!g42) & (!g43)) + ((g472) & (!g473) & (g474) & (g475) & (!g42) & (g43)) + ((g472) & (!g473) & (g474) & (g475) & (g42) & (g43)) + ((g472) & (g473) & (!g474) & (!g475) & (!g42) & (!g43)) + ((g472) & (g473) & (!g474) & (!g475) & (g42) & (!g43)) + ((g472) & (g473) & (!g474) & (g475) & (!g42) & (!g43)) + ((g472) & (g473) & (!g474) & (g475) & (g42) & (!g43)) + ((g472) & (g473) & (!g474) & (g475) & (g42) & (g43)) + ((g472) & (g473) & (g474) & (!g475) & (!g42) & (!g43)) + ((g472) & (g473) & (g474) & (!g475) & (!g42) & (g43)) + ((g472) & (g473) & (g474) & (!g475) & (g42) & (!g43)) + ((g472) & (g473) & (g474) & (g475) & (!g42) & (!g43)) + ((g472) & (g473) & (g474) & (g475) & (!g42) & (g43)) + ((g472) & (g473) & (g474) & (g475) & (g42) & (!g43)) + ((g472) & (g473) & (g474) & (g475) & (g42) & (g43)));
	assign g477 = (((!g461) & (!g466) & (!g471) & (g476) & (g60) & (g61)) + ((!g461) & (!g466) & (g471) & (!g476) & (!g60) & (g61)) + ((!g461) & (!g466) & (g471) & (g476) & (!g60) & (g61)) + ((!g461) & (!g466) & (g471) & (g476) & (g60) & (g61)) + ((!g461) & (g466) & (!g471) & (!g476) & (g60) & (!g61)) + ((!g461) & (g466) & (!g471) & (g476) & (g60) & (!g61)) + ((!g461) & (g466) & (!g471) & (g476) & (g60) & (g61)) + ((!g461) & (g466) & (g471) & (!g476) & (!g60) & (g61)) + ((!g461) & (g466) & (g471) & (!g476) & (g60) & (!g61)) + ((!g461) & (g466) & (g471) & (g476) & (!g60) & (g61)) + ((!g461) & (g466) & (g471) & (g476) & (g60) & (!g61)) + ((!g461) & (g466) & (g471) & (g476) & (g60) & (g61)) + ((g461) & (!g466) & (!g471) & (!g476) & (!g60) & (!g61)) + ((g461) & (!g466) & (!g471) & (g476) & (!g60) & (!g61)) + ((g461) & (!g466) & (!g471) & (g476) & (g60) & (g61)) + ((g461) & (!g466) & (g471) & (!g476) & (!g60) & (!g61)) + ((g461) & (!g466) & (g471) & (!g476) & (!g60) & (g61)) + ((g461) & (!g466) & (g471) & (g476) & (!g60) & (!g61)) + ((g461) & (!g466) & (g471) & (g476) & (!g60) & (g61)) + ((g461) & (!g466) & (g471) & (g476) & (g60) & (g61)) + ((g461) & (g466) & (!g471) & (!g476) & (!g60) & (!g61)) + ((g461) & (g466) & (!g471) & (!g476) & (g60) & (!g61)) + ((g461) & (g466) & (!g471) & (g476) & (!g60) & (!g61)) + ((g461) & (g466) & (!g471) & (g476) & (g60) & (!g61)) + ((g461) & (g466) & (!g471) & (g476) & (g60) & (g61)) + ((g461) & (g466) & (g471) & (!g476) & (!g60) & (!g61)) + ((g461) & (g466) & (g471) & (!g476) & (!g60) & (g61)) + ((g461) & (g466) & (g471) & (!g476) & (g60) & (!g61)) + ((g461) & (g466) & (g471) & (g476) & (!g60) & (!g61)) + ((g461) & (g466) & (g471) & (g476) & (!g60) & (g61)) + ((g461) & (g466) & (g471) & (g476) & (g60) & (!g61)) + ((g461) & (g466) & (g471) & (g476) & (g60) & (g61)));
	assign g7252 = (((!g832) & (g1441) & (!g478)) + ((!g832) & (g1441) & (g478)) + ((g832) & (!g1441) & (g478)) + ((g832) & (g1441) & (g478)));
	assign g479 = (((!g34) & (!reset) & (!g477) & (g478)) + ((!g34) & (!reset) & (g477) & (g478)) + ((g34) & (!reset) & (g477) & (!g478)) + ((g34) & (!reset) & (g477) & (g478)));
	assign g484 = (((!g480) & (!g481) & (!g482) & (g483) & (g60) & (g61)) + ((!g480) & (!g481) & (g482) & (!g483) & (!g60) & (g61)) + ((!g480) & (!g481) & (g482) & (g483) & (!g60) & (g61)) + ((!g480) & (!g481) & (g482) & (g483) & (g60) & (g61)) + ((!g480) & (g481) & (!g482) & (!g483) & (g60) & (!g61)) + ((!g480) & (g481) & (!g482) & (g483) & (g60) & (!g61)) + ((!g480) & (g481) & (!g482) & (g483) & (g60) & (g61)) + ((!g480) & (g481) & (g482) & (!g483) & (!g60) & (g61)) + ((!g480) & (g481) & (g482) & (!g483) & (g60) & (!g61)) + ((!g480) & (g481) & (g482) & (g483) & (!g60) & (g61)) + ((!g480) & (g481) & (g482) & (g483) & (g60) & (!g61)) + ((!g480) & (g481) & (g482) & (g483) & (g60) & (g61)) + ((g480) & (!g481) & (!g482) & (!g483) & (!g60) & (!g61)) + ((g480) & (!g481) & (!g482) & (g483) & (!g60) & (!g61)) + ((g480) & (!g481) & (!g482) & (g483) & (g60) & (g61)) + ((g480) & (!g481) & (g482) & (!g483) & (!g60) & (!g61)) + ((g480) & (!g481) & (g482) & (!g483) & (!g60) & (g61)) + ((g480) & (!g481) & (g482) & (g483) & (!g60) & (!g61)) + ((g480) & (!g481) & (g482) & (g483) & (!g60) & (g61)) + ((g480) & (!g481) & (g482) & (g483) & (g60) & (g61)) + ((g480) & (g481) & (!g482) & (!g483) & (!g60) & (!g61)) + ((g480) & (g481) & (!g482) & (!g483) & (g60) & (!g61)) + ((g480) & (g481) & (!g482) & (g483) & (!g60) & (!g61)) + ((g480) & (g481) & (!g482) & (g483) & (g60) & (!g61)) + ((g480) & (g481) & (!g482) & (g483) & (g60) & (g61)) + ((g480) & (g481) & (g482) & (!g483) & (!g60) & (!g61)) + ((g480) & (g481) & (g482) & (!g483) & (!g60) & (g61)) + ((g480) & (g481) & (g482) & (!g483) & (g60) & (!g61)) + ((g480) & (g481) & (g482) & (g483) & (!g60) & (!g61)) + ((g480) & (g481) & (g482) & (g483) & (!g60) & (g61)) + ((g480) & (g481) & (g482) & (g483) & (g60) & (!g61)) + ((g480) & (g481) & (g482) & (g483) & (g60) & (g61)));
	assign g489 = (((!g485) & (!g486) & (!g487) & (g488) & (g60) & (g61)) + ((!g485) & (!g486) & (g487) & (!g488) & (!g60) & (g61)) + ((!g485) & (!g486) & (g487) & (g488) & (!g60) & (g61)) + ((!g485) & (!g486) & (g487) & (g488) & (g60) & (g61)) + ((!g485) & (g486) & (!g487) & (!g488) & (g60) & (!g61)) + ((!g485) & (g486) & (!g487) & (g488) & (g60) & (!g61)) + ((!g485) & (g486) & (!g487) & (g488) & (g60) & (g61)) + ((!g485) & (g486) & (g487) & (!g488) & (!g60) & (g61)) + ((!g485) & (g486) & (g487) & (!g488) & (g60) & (!g61)) + ((!g485) & (g486) & (g487) & (g488) & (!g60) & (g61)) + ((!g485) & (g486) & (g487) & (g488) & (g60) & (!g61)) + ((!g485) & (g486) & (g487) & (g488) & (g60) & (g61)) + ((g485) & (!g486) & (!g487) & (!g488) & (!g60) & (!g61)) + ((g485) & (!g486) & (!g487) & (g488) & (!g60) & (!g61)) + ((g485) & (!g486) & (!g487) & (g488) & (g60) & (g61)) + ((g485) & (!g486) & (g487) & (!g488) & (!g60) & (!g61)) + ((g485) & (!g486) & (g487) & (!g488) & (!g60) & (g61)) + ((g485) & (!g486) & (g487) & (g488) & (!g60) & (!g61)) + ((g485) & (!g486) & (g487) & (g488) & (!g60) & (g61)) + ((g485) & (!g486) & (g487) & (g488) & (g60) & (g61)) + ((g485) & (g486) & (!g487) & (!g488) & (!g60) & (!g61)) + ((g485) & (g486) & (!g487) & (!g488) & (g60) & (!g61)) + ((g485) & (g486) & (!g487) & (g488) & (!g60) & (!g61)) + ((g485) & (g486) & (!g487) & (g488) & (g60) & (!g61)) + ((g485) & (g486) & (!g487) & (g488) & (g60) & (g61)) + ((g485) & (g486) & (g487) & (!g488) & (!g60) & (!g61)) + ((g485) & (g486) & (g487) & (!g488) & (!g60) & (g61)) + ((g485) & (g486) & (g487) & (!g488) & (g60) & (!g61)) + ((g485) & (g486) & (g487) & (g488) & (!g60) & (!g61)) + ((g485) & (g486) & (g487) & (g488) & (!g60) & (g61)) + ((g485) & (g486) & (g487) & (g488) & (g60) & (!g61)) + ((g485) & (g486) & (g487) & (g488) & (g60) & (g61)));
	assign g494 = (((!g490) & (!g491) & (!g492) & (g493) & (g60) & (g61)) + ((!g490) & (!g491) & (g492) & (!g493) & (!g60) & (g61)) + ((!g490) & (!g491) & (g492) & (g493) & (!g60) & (g61)) + ((!g490) & (!g491) & (g492) & (g493) & (g60) & (g61)) + ((!g490) & (g491) & (!g492) & (!g493) & (g60) & (!g61)) + ((!g490) & (g491) & (!g492) & (g493) & (g60) & (!g61)) + ((!g490) & (g491) & (!g492) & (g493) & (g60) & (g61)) + ((!g490) & (g491) & (g492) & (!g493) & (!g60) & (g61)) + ((!g490) & (g491) & (g492) & (!g493) & (g60) & (!g61)) + ((!g490) & (g491) & (g492) & (g493) & (!g60) & (g61)) + ((!g490) & (g491) & (g492) & (g493) & (g60) & (!g61)) + ((!g490) & (g491) & (g492) & (g493) & (g60) & (g61)) + ((g490) & (!g491) & (!g492) & (!g493) & (!g60) & (!g61)) + ((g490) & (!g491) & (!g492) & (g493) & (!g60) & (!g61)) + ((g490) & (!g491) & (!g492) & (g493) & (g60) & (g61)) + ((g490) & (!g491) & (g492) & (!g493) & (!g60) & (!g61)) + ((g490) & (!g491) & (g492) & (!g493) & (!g60) & (g61)) + ((g490) & (!g491) & (g492) & (g493) & (!g60) & (!g61)) + ((g490) & (!g491) & (g492) & (g493) & (!g60) & (g61)) + ((g490) & (!g491) & (g492) & (g493) & (g60) & (g61)) + ((g490) & (g491) & (!g492) & (!g493) & (!g60) & (!g61)) + ((g490) & (g491) & (!g492) & (!g493) & (g60) & (!g61)) + ((g490) & (g491) & (!g492) & (g493) & (!g60) & (!g61)) + ((g490) & (g491) & (!g492) & (g493) & (g60) & (!g61)) + ((g490) & (g491) & (!g492) & (g493) & (g60) & (g61)) + ((g490) & (g491) & (g492) & (!g493) & (!g60) & (!g61)) + ((g490) & (g491) & (g492) & (!g493) & (!g60) & (g61)) + ((g490) & (g491) & (g492) & (!g493) & (g60) & (!g61)) + ((g490) & (g491) & (g492) & (g493) & (!g60) & (!g61)) + ((g490) & (g491) & (g492) & (g493) & (!g60) & (g61)) + ((g490) & (g491) & (g492) & (g493) & (g60) & (!g61)) + ((g490) & (g491) & (g492) & (g493) & (g60) & (g61)));
	assign g499 = (((!g495) & (!g496) & (!g497) & (g498) & (g60) & (g61)) + ((!g495) & (!g496) & (g497) & (!g498) & (!g60) & (g61)) + ((!g495) & (!g496) & (g497) & (g498) & (!g60) & (g61)) + ((!g495) & (!g496) & (g497) & (g498) & (g60) & (g61)) + ((!g495) & (g496) & (!g497) & (!g498) & (g60) & (!g61)) + ((!g495) & (g496) & (!g497) & (g498) & (g60) & (!g61)) + ((!g495) & (g496) & (!g497) & (g498) & (g60) & (g61)) + ((!g495) & (g496) & (g497) & (!g498) & (!g60) & (g61)) + ((!g495) & (g496) & (g497) & (!g498) & (g60) & (!g61)) + ((!g495) & (g496) & (g497) & (g498) & (!g60) & (g61)) + ((!g495) & (g496) & (g497) & (g498) & (g60) & (!g61)) + ((!g495) & (g496) & (g497) & (g498) & (g60) & (g61)) + ((g495) & (!g496) & (!g497) & (!g498) & (!g60) & (!g61)) + ((g495) & (!g496) & (!g497) & (g498) & (!g60) & (!g61)) + ((g495) & (!g496) & (!g497) & (g498) & (g60) & (g61)) + ((g495) & (!g496) & (g497) & (!g498) & (!g60) & (!g61)) + ((g495) & (!g496) & (g497) & (!g498) & (!g60) & (g61)) + ((g495) & (!g496) & (g497) & (g498) & (!g60) & (!g61)) + ((g495) & (!g496) & (g497) & (g498) & (!g60) & (g61)) + ((g495) & (!g496) & (g497) & (g498) & (g60) & (g61)) + ((g495) & (g496) & (!g497) & (!g498) & (!g60) & (!g61)) + ((g495) & (g496) & (!g497) & (!g498) & (g60) & (!g61)) + ((g495) & (g496) & (!g497) & (g498) & (!g60) & (!g61)) + ((g495) & (g496) & (!g497) & (g498) & (g60) & (!g61)) + ((g495) & (g496) & (!g497) & (g498) & (g60) & (g61)) + ((g495) & (g496) & (g497) & (!g498) & (!g60) & (!g61)) + ((g495) & (g496) & (g497) & (!g498) & (!g60) & (g61)) + ((g495) & (g496) & (g497) & (!g498) & (g60) & (!g61)) + ((g495) & (g496) & (g497) & (g498) & (!g60) & (!g61)) + ((g495) & (g496) & (g497) & (g498) & (!g60) & (g61)) + ((g495) & (g496) & (g497) & (g498) & (g60) & (!g61)) + ((g495) & (g496) & (g497) & (g498) & (g60) & (g61)));
	assign g500 = (((!g484) & (!g489) & (!g494) & (g499) & (g42) & (g43)) + ((!g484) & (!g489) & (g494) & (!g499) & (!g42) & (g43)) + ((!g484) & (!g489) & (g494) & (g499) & (!g42) & (g43)) + ((!g484) & (!g489) & (g494) & (g499) & (g42) & (g43)) + ((!g484) & (g489) & (!g494) & (!g499) & (g42) & (!g43)) + ((!g484) & (g489) & (!g494) & (g499) & (g42) & (!g43)) + ((!g484) & (g489) & (!g494) & (g499) & (g42) & (g43)) + ((!g484) & (g489) & (g494) & (!g499) & (!g42) & (g43)) + ((!g484) & (g489) & (g494) & (!g499) & (g42) & (!g43)) + ((!g484) & (g489) & (g494) & (g499) & (!g42) & (g43)) + ((!g484) & (g489) & (g494) & (g499) & (g42) & (!g43)) + ((!g484) & (g489) & (g494) & (g499) & (g42) & (g43)) + ((g484) & (!g489) & (!g494) & (!g499) & (!g42) & (!g43)) + ((g484) & (!g489) & (!g494) & (g499) & (!g42) & (!g43)) + ((g484) & (!g489) & (!g494) & (g499) & (g42) & (g43)) + ((g484) & (!g489) & (g494) & (!g499) & (!g42) & (!g43)) + ((g484) & (!g489) & (g494) & (!g499) & (!g42) & (g43)) + ((g484) & (!g489) & (g494) & (g499) & (!g42) & (!g43)) + ((g484) & (!g489) & (g494) & (g499) & (!g42) & (g43)) + ((g484) & (!g489) & (g494) & (g499) & (g42) & (g43)) + ((g484) & (g489) & (!g494) & (!g499) & (!g42) & (!g43)) + ((g484) & (g489) & (!g494) & (!g499) & (g42) & (!g43)) + ((g484) & (g489) & (!g494) & (g499) & (!g42) & (!g43)) + ((g484) & (g489) & (!g494) & (g499) & (g42) & (!g43)) + ((g484) & (g489) & (!g494) & (g499) & (g42) & (g43)) + ((g484) & (g489) & (g494) & (!g499) & (!g42) & (!g43)) + ((g484) & (g489) & (g494) & (!g499) & (!g42) & (g43)) + ((g484) & (g489) & (g494) & (!g499) & (g42) & (!g43)) + ((g484) & (g489) & (g494) & (g499) & (!g42) & (!g43)) + ((g484) & (g489) & (g494) & (g499) & (!g42) & (g43)) + ((g484) & (g489) & (g494) & (g499) & (g42) & (!g43)) + ((g484) & (g489) & (g494) & (g499) & (g42) & (g43)));
	assign g7253 = (((!g832) & (g1475) & (!g501)) + ((!g832) & (g1475) & (g501)) + ((g832) & (!g1475) & (g501)) + ((g832) & (g1475) & (g501)));
	assign g502 = (((!g34) & (!reset) & (!g500) & (g501)) + ((!g34) & (!reset) & (g500) & (g501)) + ((g34) & (!reset) & (g500) & (!g501)) + ((g34) & (!reset) & (g500) & (g501)));
	assign g507 = (((!g503) & (!g504) & (!g505) & (g506) & (g42) & (g43)) + ((!g503) & (!g504) & (g505) & (!g506) & (!g42) & (g43)) + ((!g503) & (!g504) & (g505) & (g506) & (!g42) & (g43)) + ((!g503) & (!g504) & (g505) & (g506) & (g42) & (g43)) + ((!g503) & (g504) & (!g505) & (!g506) & (g42) & (!g43)) + ((!g503) & (g504) & (!g505) & (g506) & (g42) & (!g43)) + ((!g503) & (g504) & (!g505) & (g506) & (g42) & (g43)) + ((!g503) & (g504) & (g505) & (!g506) & (!g42) & (g43)) + ((!g503) & (g504) & (g505) & (!g506) & (g42) & (!g43)) + ((!g503) & (g504) & (g505) & (g506) & (!g42) & (g43)) + ((!g503) & (g504) & (g505) & (g506) & (g42) & (!g43)) + ((!g503) & (g504) & (g505) & (g506) & (g42) & (g43)) + ((g503) & (!g504) & (!g505) & (!g506) & (!g42) & (!g43)) + ((g503) & (!g504) & (!g505) & (g506) & (!g42) & (!g43)) + ((g503) & (!g504) & (!g505) & (g506) & (g42) & (g43)) + ((g503) & (!g504) & (g505) & (!g506) & (!g42) & (!g43)) + ((g503) & (!g504) & (g505) & (!g506) & (!g42) & (g43)) + ((g503) & (!g504) & (g505) & (g506) & (!g42) & (!g43)) + ((g503) & (!g504) & (g505) & (g506) & (!g42) & (g43)) + ((g503) & (!g504) & (g505) & (g506) & (g42) & (g43)) + ((g503) & (g504) & (!g505) & (!g506) & (!g42) & (!g43)) + ((g503) & (g504) & (!g505) & (!g506) & (g42) & (!g43)) + ((g503) & (g504) & (!g505) & (g506) & (!g42) & (!g43)) + ((g503) & (g504) & (!g505) & (g506) & (g42) & (!g43)) + ((g503) & (g504) & (!g505) & (g506) & (g42) & (g43)) + ((g503) & (g504) & (g505) & (!g506) & (!g42) & (!g43)) + ((g503) & (g504) & (g505) & (!g506) & (!g42) & (g43)) + ((g503) & (g504) & (g505) & (!g506) & (g42) & (!g43)) + ((g503) & (g504) & (g505) & (g506) & (!g42) & (!g43)) + ((g503) & (g504) & (g505) & (g506) & (!g42) & (g43)) + ((g503) & (g504) & (g505) & (g506) & (g42) & (!g43)) + ((g503) & (g504) & (g505) & (g506) & (g42) & (g43)));
	assign g512 = (((!g508) & (!g509) & (!g510) & (g511) & (g42) & (g43)) + ((!g508) & (!g509) & (g510) & (!g511) & (!g42) & (g43)) + ((!g508) & (!g509) & (g510) & (g511) & (!g42) & (g43)) + ((!g508) & (!g509) & (g510) & (g511) & (g42) & (g43)) + ((!g508) & (g509) & (!g510) & (!g511) & (g42) & (!g43)) + ((!g508) & (g509) & (!g510) & (g511) & (g42) & (!g43)) + ((!g508) & (g509) & (!g510) & (g511) & (g42) & (g43)) + ((!g508) & (g509) & (g510) & (!g511) & (!g42) & (g43)) + ((!g508) & (g509) & (g510) & (!g511) & (g42) & (!g43)) + ((!g508) & (g509) & (g510) & (g511) & (!g42) & (g43)) + ((!g508) & (g509) & (g510) & (g511) & (g42) & (!g43)) + ((!g508) & (g509) & (g510) & (g511) & (g42) & (g43)) + ((g508) & (!g509) & (!g510) & (!g511) & (!g42) & (!g43)) + ((g508) & (!g509) & (!g510) & (g511) & (!g42) & (!g43)) + ((g508) & (!g509) & (!g510) & (g511) & (g42) & (g43)) + ((g508) & (!g509) & (g510) & (!g511) & (!g42) & (!g43)) + ((g508) & (!g509) & (g510) & (!g511) & (!g42) & (g43)) + ((g508) & (!g509) & (g510) & (g511) & (!g42) & (!g43)) + ((g508) & (!g509) & (g510) & (g511) & (!g42) & (g43)) + ((g508) & (!g509) & (g510) & (g511) & (g42) & (g43)) + ((g508) & (g509) & (!g510) & (!g511) & (!g42) & (!g43)) + ((g508) & (g509) & (!g510) & (!g511) & (g42) & (!g43)) + ((g508) & (g509) & (!g510) & (g511) & (!g42) & (!g43)) + ((g508) & (g509) & (!g510) & (g511) & (g42) & (!g43)) + ((g508) & (g509) & (!g510) & (g511) & (g42) & (g43)) + ((g508) & (g509) & (g510) & (!g511) & (!g42) & (!g43)) + ((g508) & (g509) & (g510) & (!g511) & (!g42) & (g43)) + ((g508) & (g509) & (g510) & (!g511) & (g42) & (!g43)) + ((g508) & (g509) & (g510) & (g511) & (!g42) & (!g43)) + ((g508) & (g509) & (g510) & (g511) & (!g42) & (g43)) + ((g508) & (g509) & (g510) & (g511) & (g42) & (!g43)) + ((g508) & (g509) & (g510) & (g511) & (g42) & (g43)));
	assign g517 = (((!g513) & (!g514) & (!g515) & (g516) & (g42) & (g43)) + ((!g513) & (!g514) & (g515) & (!g516) & (!g42) & (g43)) + ((!g513) & (!g514) & (g515) & (g516) & (!g42) & (g43)) + ((!g513) & (!g514) & (g515) & (g516) & (g42) & (g43)) + ((!g513) & (g514) & (!g515) & (!g516) & (g42) & (!g43)) + ((!g513) & (g514) & (!g515) & (g516) & (g42) & (!g43)) + ((!g513) & (g514) & (!g515) & (g516) & (g42) & (g43)) + ((!g513) & (g514) & (g515) & (!g516) & (!g42) & (g43)) + ((!g513) & (g514) & (g515) & (!g516) & (g42) & (!g43)) + ((!g513) & (g514) & (g515) & (g516) & (!g42) & (g43)) + ((!g513) & (g514) & (g515) & (g516) & (g42) & (!g43)) + ((!g513) & (g514) & (g515) & (g516) & (g42) & (g43)) + ((g513) & (!g514) & (!g515) & (!g516) & (!g42) & (!g43)) + ((g513) & (!g514) & (!g515) & (g516) & (!g42) & (!g43)) + ((g513) & (!g514) & (!g515) & (g516) & (g42) & (g43)) + ((g513) & (!g514) & (g515) & (!g516) & (!g42) & (!g43)) + ((g513) & (!g514) & (g515) & (!g516) & (!g42) & (g43)) + ((g513) & (!g514) & (g515) & (g516) & (!g42) & (!g43)) + ((g513) & (!g514) & (g515) & (g516) & (!g42) & (g43)) + ((g513) & (!g514) & (g515) & (g516) & (g42) & (g43)) + ((g513) & (g514) & (!g515) & (!g516) & (!g42) & (!g43)) + ((g513) & (g514) & (!g515) & (!g516) & (g42) & (!g43)) + ((g513) & (g514) & (!g515) & (g516) & (!g42) & (!g43)) + ((g513) & (g514) & (!g515) & (g516) & (g42) & (!g43)) + ((g513) & (g514) & (!g515) & (g516) & (g42) & (g43)) + ((g513) & (g514) & (g515) & (!g516) & (!g42) & (!g43)) + ((g513) & (g514) & (g515) & (!g516) & (!g42) & (g43)) + ((g513) & (g514) & (g515) & (!g516) & (g42) & (!g43)) + ((g513) & (g514) & (g515) & (g516) & (!g42) & (!g43)) + ((g513) & (g514) & (g515) & (g516) & (!g42) & (g43)) + ((g513) & (g514) & (g515) & (g516) & (g42) & (!g43)) + ((g513) & (g514) & (g515) & (g516) & (g42) & (g43)));
	assign g522 = (((!g518) & (!g519) & (!g520) & (g521) & (g42) & (g43)) + ((!g518) & (!g519) & (g520) & (!g521) & (!g42) & (g43)) + ((!g518) & (!g519) & (g520) & (g521) & (!g42) & (g43)) + ((!g518) & (!g519) & (g520) & (g521) & (g42) & (g43)) + ((!g518) & (g519) & (!g520) & (!g521) & (g42) & (!g43)) + ((!g518) & (g519) & (!g520) & (g521) & (g42) & (!g43)) + ((!g518) & (g519) & (!g520) & (g521) & (g42) & (g43)) + ((!g518) & (g519) & (g520) & (!g521) & (!g42) & (g43)) + ((!g518) & (g519) & (g520) & (!g521) & (g42) & (!g43)) + ((!g518) & (g519) & (g520) & (g521) & (!g42) & (g43)) + ((!g518) & (g519) & (g520) & (g521) & (g42) & (!g43)) + ((!g518) & (g519) & (g520) & (g521) & (g42) & (g43)) + ((g518) & (!g519) & (!g520) & (!g521) & (!g42) & (!g43)) + ((g518) & (!g519) & (!g520) & (g521) & (!g42) & (!g43)) + ((g518) & (!g519) & (!g520) & (g521) & (g42) & (g43)) + ((g518) & (!g519) & (g520) & (!g521) & (!g42) & (!g43)) + ((g518) & (!g519) & (g520) & (!g521) & (!g42) & (g43)) + ((g518) & (!g519) & (g520) & (g521) & (!g42) & (!g43)) + ((g518) & (!g519) & (g520) & (g521) & (!g42) & (g43)) + ((g518) & (!g519) & (g520) & (g521) & (g42) & (g43)) + ((g518) & (g519) & (!g520) & (!g521) & (!g42) & (!g43)) + ((g518) & (g519) & (!g520) & (!g521) & (g42) & (!g43)) + ((g518) & (g519) & (!g520) & (g521) & (!g42) & (!g43)) + ((g518) & (g519) & (!g520) & (g521) & (g42) & (!g43)) + ((g518) & (g519) & (!g520) & (g521) & (g42) & (g43)) + ((g518) & (g519) & (g520) & (!g521) & (!g42) & (!g43)) + ((g518) & (g519) & (g520) & (!g521) & (!g42) & (g43)) + ((g518) & (g519) & (g520) & (!g521) & (g42) & (!g43)) + ((g518) & (g519) & (g520) & (g521) & (!g42) & (!g43)) + ((g518) & (g519) & (g520) & (g521) & (!g42) & (g43)) + ((g518) & (g519) & (g520) & (g521) & (g42) & (!g43)) + ((g518) & (g519) & (g520) & (g521) & (g42) & (g43)));
	assign g523 = (((!g507) & (!g512) & (!g517) & (g522) & (g60) & (g61)) + ((!g507) & (!g512) & (g517) & (!g522) & (!g60) & (g61)) + ((!g507) & (!g512) & (g517) & (g522) & (!g60) & (g61)) + ((!g507) & (!g512) & (g517) & (g522) & (g60) & (g61)) + ((!g507) & (g512) & (!g517) & (!g522) & (g60) & (!g61)) + ((!g507) & (g512) & (!g517) & (g522) & (g60) & (!g61)) + ((!g507) & (g512) & (!g517) & (g522) & (g60) & (g61)) + ((!g507) & (g512) & (g517) & (!g522) & (!g60) & (g61)) + ((!g507) & (g512) & (g517) & (!g522) & (g60) & (!g61)) + ((!g507) & (g512) & (g517) & (g522) & (!g60) & (g61)) + ((!g507) & (g512) & (g517) & (g522) & (g60) & (!g61)) + ((!g507) & (g512) & (g517) & (g522) & (g60) & (g61)) + ((g507) & (!g512) & (!g517) & (!g522) & (!g60) & (!g61)) + ((g507) & (!g512) & (!g517) & (g522) & (!g60) & (!g61)) + ((g507) & (!g512) & (!g517) & (g522) & (g60) & (g61)) + ((g507) & (!g512) & (g517) & (!g522) & (!g60) & (!g61)) + ((g507) & (!g512) & (g517) & (!g522) & (!g60) & (g61)) + ((g507) & (!g512) & (g517) & (g522) & (!g60) & (!g61)) + ((g507) & (!g512) & (g517) & (g522) & (!g60) & (g61)) + ((g507) & (!g512) & (g517) & (g522) & (g60) & (g61)) + ((g507) & (g512) & (!g517) & (!g522) & (!g60) & (!g61)) + ((g507) & (g512) & (!g517) & (!g522) & (g60) & (!g61)) + ((g507) & (g512) & (!g517) & (g522) & (!g60) & (!g61)) + ((g507) & (g512) & (!g517) & (g522) & (g60) & (!g61)) + ((g507) & (g512) & (!g517) & (g522) & (g60) & (g61)) + ((g507) & (g512) & (g517) & (!g522) & (!g60) & (!g61)) + ((g507) & (g512) & (g517) & (!g522) & (!g60) & (g61)) + ((g507) & (g512) & (g517) & (!g522) & (g60) & (!g61)) + ((g507) & (g512) & (g517) & (g522) & (!g60) & (!g61)) + ((g507) & (g512) & (g517) & (g522) & (!g60) & (g61)) + ((g507) & (g512) & (g517) & (g522) & (g60) & (!g61)) + ((g507) & (g512) & (g517) & (g522) & (g60) & (g61)));
	assign g7254 = (((!g832) & (g1508) & (!g524)) + ((!g832) & (g1508) & (g524)) + ((g832) & (!g1508) & (g524)) + ((g832) & (g1508) & (g524)));
	assign g525 = (((!g34) & (!reset) & (!g523) & (g524)) + ((!g34) & (!reset) & (g523) & (g524)) + ((g34) & (!reset) & (g523) & (!g524)) + ((g34) & (!reset) & (g523) & (g524)));
	assign g530 = (((!g526) & (!g527) & (!g528) & (g529) & (g60) & (g61)) + ((!g526) & (!g527) & (g528) & (!g529) & (!g60) & (g61)) + ((!g526) & (!g527) & (g528) & (g529) & (!g60) & (g61)) + ((!g526) & (!g527) & (g528) & (g529) & (g60) & (g61)) + ((!g526) & (g527) & (!g528) & (!g529) & (g60) & (!g61)) + ((!g526) & (g527) & (!g528) & (g529) & (g60) & (!g61)) + ((!g526) & (g527) & (!g528) & (g529) & (g60) & (g61)) + ((!g526) & (g527) & (g528) & (!g529) & (!g60) & (g61)) + ((!g526) & (g527) & (g528) & (!g529) & (g60) & (!g61)) + ((!g526) & (g527) & (g528) & (g529) & (!g60) & (g61)) + ((!g526) & (g527) & (g528) & (g529) & (g60) & (!g61)) + ((!g526) & (g527) & (g528) & (g529) & (g60) & (g61)) + ((g526) & (!g527) & (!g528) & (!g529) & (!g60) & (!g61)) + ((g526) & (!g527) & (!g528) & (g529) & (!g60) & (!g61)) + ((g526) & (!g527) & (!g528) & (g529) & (g60) & (g61)) + ((g526) & (!g527) & (g528) & (!g529) & (!g60) & (!g61)) + ((g526) & (!g527) & (g528) & (!g529) & (!g60) & (g61)) + ((g526) & (!g527) & (g528) & (g529) & (!g60) & (!g61)) + ((g526) & (!g527) & (g528) & (g529) & (!g60) & (g61)) + ((g526) & (!g527) & (g528) & (g529) & (g60) & (g61)) + ((g526) & (g527) & (!g528) & (!g529) & (!g60) & (!g61)) + ((g526) & (g527) & (!g528) & (!g529) & (g60) & (!g61)) + ((g526) & (g527) & (!g528) & (g529) & (!g60) & (!g61)) + ((g526) & (g527) & (!g528) & (g529) & (g60) & (!g61)) + ((g526) & (g527) & (!g528) & (g529) & (g60) & (g61)) + ((g526) & (g527) & (g528) & (!g529) & (!g60) & (!g61)) + ((g526) & (g527) & (g528) & (!g529) & (!g60) & (g61)) + ((g526) & (g527) & (g528) & (!g529) & (g60) & (!g61)) + ((g526) & (g527) & (g528) & (g529) & (!g60) & (!g61)) + ((g526) & (g527) & (g528) & (g529) & (!g60) & (g61)) + ((g526) & (g527) & (g528) & (g529) & (g60) & (!g61)) + ((g526) & (g527) & (g528) & (g529) & (g60) & (g61)));
	assign g535 = (((!g531) & (!g532) & (!g533) & (g534) & (g60) & (g61)) + ((!g531) & (!g532) & (g533) & (!g534) & (!g60) & (g61)) + ((!g531) & (!g532) & (g533) & (g534) & (!g60) & (g61)) + ((!g531) & (!g532) & (g533) & (g534) & (g60) & (g61)) + ((!g531) & (g532) & (!g533) & (!g534) & (g60) & (!g61)) + ((!g531) & (g532) & (!g533) & (g534) & (g60) & (!g61)) + ((!g531) & (g532) & (!g533) & (g534) & (g60) & (g61)) + ((!g531) & (g532) & (g533) & (!g534) & (!g60) & (g61)) + ((!g531) & (g532) & (g533) & (!g534) & (g60) & (!g61)) + ((!g531) & (g532) & (g533) & (g534) & (!g60) & (g61)) + ((!g531) & (g532) & (g533) & (g534) & (g60) & (!g61)) + ((!g531) & (g532) & (g533) & (g534) & (g60) & (g61)) + ((g531) & (!g532) & (!g533) & (!g534) & (!g60) & (!g61)) + ((g531) & (!g532) & (!g533) & (g534) & (!g60) & (!g61)) + ((g531) & (!g532) & (!g533) & (g534) & (g60) & (g61)) + ((g531) & (!g532) & (g533) & (!g534) & (!g60) & (!g61)) + ((g531) & (!g532) & (g533) & (!g534) & (!g60) & (g61)) + ((g531) & (!g532) & (g533) & (g534) & (!g60) & (!g61)) + ((g531) & (!g532) & (g533) & (g534) & (!g60) & (g61)) + ((g531) & (!g532) & (g533) & (g534) & (g60) & (g61)) + ((g531) & (g532) & (!g533) & (!g534) & (!g60) & (!g61)) + ((g531) & (g532) & (!g533) & (!g534) & (g60) & (!g61)) + ((g531) & (g532) & (!g533) & (g534) & (!g60) & (!g61)) + ((g531) & (g532) & (!g533) & (g534) & (g60) & (!g61)) + ((g531) & (g532) & (!g533) & (g534) & (g60) & (g61)) + ((g531) & (g532) & (g533) & (!g534) & (!g60) & (!g61)) + ((g531) & (g532) & (g533) & (!g534) & (!g60) & (g61)) + ((g531) & (g532) & (g533) & (!g534) & (g60) & (!g61)) + ((g531) & (g532) & (g533) & (g534) & (!g60) & (!g61)) + ((g531) & (g532) & (g533) & (g534) & (!g60) & (g61)) + ((g531) & (g532) & (g533) & (g534) & (g60) & (!g61)) + ((g531) & (g532) & (g533) & (g534) & (g60) & (g61)));
	assign g540 = (((!g536) & (!g537) & (!g538) & (g539) & (g60) & (g61)) + ((!g536) & (!g537) & (g538) & (!g539) & (!g60) & (g61)) + ((!g536) & (!g537) & (g538) & (g539) & (!g60) & (g61)) + ((!g536) & (!g537) & (g538) & (g539) & (g60) & (g61)) + ((!g536) & (g537) & (!g538) & (!g539) & (g60) & (!g61)) + ((!g536) & (g537) & (!g538) & (g539) & (g60) & (!g61)) + ((!g536) & (g537) & (!g538) & (g539) & (g60) & (g61)) + ((!g536) & (g537) & (g538) & (!g539) & (!g60) & (g61)) + ((!g536) & (g537) & (g538) & (!g539) & (g60) & (!g61)) + ((!g536) & (g537) & (g538) & (g539) & (!g60) & (g61)) + ((!g536) & (g537) & (g538) & (g539) & (g60) & (!g61)) + ((!g536) & (g537) & (g538) & (g539) & (g60) & (g61)) + ((g536) & (!g537) & (!g538) & (!g539) & (!g60) & (!g61)) + ((g536) & (!g537) & (!g538) & (g539) & (!g60) & (!g61)) + ((g536) & (!g537) & (!g538) & (g539) & (g60) & (g61)) + ((g536) & (!g537) & (g538) & (!g539) & (!g60) & (!g61)) + ((g536) & (!g537) & (g538) & (!g539) & (!g60) & (g61)) + ((g536) & (!g537) & (g538) & (g539) & (!g60) & (!g61)) + ((g536) & (!g537) & (g538) & (g539) & (!g60) & (g61)) + ((g536) & (!g537) & (g538) & (g539) & (g60) & (g61)) + ((g536) & (g537) & (!g538) & (!g539) & (!g60) & (!g61)) + ((g536) & (g537) & (!g538) & (!g539) & (g60) & (!g61)) + ((g536) & (g537) & (!g538) & (g539) & (!g60) & (!g61)) + ((g536) & (g537) & (!g538) & (g539) & (g60) & (!g61)) + ((g536) & (g537) & (!g538) & (g539) & (g60) & (g61)) + ((g536) & (g537) & (g538) & (!g539) & (!g60) & (!g61)) + ((g536) & (g537) & (g538) & (!g539) & (!g60) & (g61)) + ((g536) & (g537) & (g538) & (!g539) & (g60) & (!g61)) + ((g536) & (g537) & (g538) & (g539) & (!g60) & (!g61)) + ((g536) & (g537) & (g538) & (g539) & (!g60) & (g61)) + ((g536) & (g537) & (g538) & (g539) & (g60) & (!g61)) + ((g536) & (g537) & (g538) & (g539) & (g60) & (g61)));
	assign g545 = (((!g541) & (!g542) & (!g543) & (g544) & (g60) & (g61)) + ((!g541) & (!g542) & (g543) & (!g544) & (!g60) & (g61)) + ((!g541) & (!g542) & (g543) & (g544) & (!g60) & (g61)) + ((!g541) & (!g542) & (g543) & (g544) & (g60) & (g61)) + ((!g541) & (g542) & (!g543) & (!g544) & (g60) & (!g61)) + ((!g541) & (g542) & (!g543) & (g544) & (g60) & (!g61)) + ((!g541) & (g542) & (!g543) & (g544) & (g60) & (g61)) + ((!g541) & (g542) & (g543) & (!g544) & (!g60) & (g61)) + ((!g541) & (g542) & (g543) & (!g544) & (g60) & (!g61)) + ((!g541) & (g542) & (g543) & (g544) & (!g60) & (g61)) + ((!g541) & (g542) & (g543) & (g544) & (g60) & (!g61)) + ((!g541) & (g542) & (g543) & (g544) & (g60) & (g61)) + ((g541) & (!g542) & (!g543) & (!g544) & (!g60) & (!g61)) + ((g541) & (!g542) & (!g543) & (g544) & (!g60) & (!g61)) + ((g541) & (!g542) & (!g543) & (g544) & (g60) & (g61)) + ((g541) & (!g542) & (g543) & (!g544) & (!g60) & (!g61)) + ((g541) & (!g542) & (g543) & (!g544) & (!g60) & (g61)) + ((g541) & (!g542) & (g543) & (g544) & (!g60) & (!g61)) + ((g541) & (!g542) & (g543) & (g544) & (!g60) & (g61)) + ((g541) & (!g542) & (g543) & (g544) & (g60) & (g61)) + ((g541) & (g542) & (!g543) & (!g544) & (!g60) & (!g61)) + ((g541) & (g542) & (!g543) & (!g544) & (g60) & (!g61)) + ((g541) & (g542) & (!g543) & (g544) & (!g60) & (!g61)) + ((g541) & (g542) & (!g543) & (g544) & (g60) & (!g61)) + ((g541) & (g542) & (!g543) & (g544) & (g60) & (g61)) + ((g541) & (g542) & (g543) & (!g544) & (!g60) & (!g61)) + ((g541) & (g542) & (g543) & (!g544) & (!g60) & (g61)) + ((g541) & (g542) & (g543) & (!g544) & (g60) & (!g61)) + ((g541) & (g542) & (g543) & (g544) & (!g60) & (!g61)) + ((g541) & (g542) & (g543) & (g544) & (!g60) & (g61)) + ((g541) & (g542) & (g543) & (g544) & (g60) & (!g61)) + ((g541) & (g542) & (g543) & (g544) & (g60) & (g61)));
	assign g546 = (((!g530) & (!g535) & (!g540) & (g545) & (g42) & (g43)) + ((!g530) & (!g535) & (g540) & (!g545) & (!g42) & (g43)) + ((!g530) & (!g535) & (g540) & (g545) & (!g42) & (g43)) + ((!g530) & (!g535) & (g540) & (g545) & (g42) & (g43)) + ((!g530) & (g535) & (!g540) & (!g545) & (g42) & (!g43)) + ((!g530) & (g535) & (!g540) & (g545) & (g42) & (!g43)) + ((!g530) & (g535) & (!g540) & (g545) & (g42) & (g43)) + ((!g530) & (g535) & (g540) & (!g545) & (!g42) & (g43)) + ((!g530) & (g535) & (g540) & (!g545) & (g42) & (!g43)) + ((!g530) & (g535) & (g540) & (g545) & (!g42) & (g43)) + ((!g530) & (g535) & (g540) & (g545) & (g42) & (!g43)) + ((!g530) & (g535) & (g540) & (g545) & (g42) & (g43)) + ((g530) & (!g535) & (!g540) & (!g545) & (!g42) & (!g43)) + ((g530) & (!g535) & (!g540) & (g545) & (!g42) & (!g43)) + ((g530) & (!g535) & (!g540) & (g545) & (g42) & (g43)) + ((g530) & (!g535) & (g540) & (!g545) & (!g42) & (!g43)) + ((g530) & (!g535) & (g540) & (!g545) & (!g42) & (g43)) + ((g530) & (!g535) & (g540) & (g545) & (!g42) & (!g43)) + ((g530) & (!g535) & (g540) & (g545) & (!g42) & (g43)) + ((g530) & (!g535) & (g540) & (g545) & (g42) & (g43)) + ((g530) & (g535) & (!g540) & (!g545) & (!g42) & (!g43)) + ((g530) & (g535) & (!g540) & (!g545) & (g42) & (!g43)) + ((g530) & (g535) & (!g540) & (g545) & (!g42) & (!g43)) + ((g530) & (g535) & (!g540) & (g545) & (g42) & (!g43)) + ((g530) & (g535) & (!g540) & (g545) & (g42) & (g43)) + ((g530) & (g535) & (g540) & (!g545) & (!g42) & (!g43)) + ((g530) & (g535) & (g540) & (!g545) & (!g42) & (g43)) + ((g530) & (g535) & (g540) & (!g545) & (g42) & (!g43)) + ((g530) & (g535) & (g540) & (g545) & (!g42) & (!g43)) + ((g530) & (g535) & (g540) & (g545) & (!g42) & (g43)) + ((g530) & (g535) & (g540) & (g545) & (g42) & (!g43)) + ((g530) & (g535) & (g540) & (g545) & (g42) & (g43)));
	assign g7255 = (((!g832) & (g1545) & (!g547)) + ((!g832) & (g1545) & (g547)) + ((g832) & (!g1545) & (g547)) + ((g832) & (g1545) & (g547)));
	assign g548 = (((!g34) & (!reset) & (!g546) & (g547)) + ((!g34) & (!reset) & (g546) & (g547)) + ((g34) & (!reset) & (g546) & (!g547)) + ((g34) & (!reset) & (g546) & (g547)));
	assign g553 = (((!g549) & (!g550) & (!g551) & (g552) & (g42) & (g43)) + ((!g549) & (!g550) & (g551) & (!g552) & (!g42) & (g43)) + ((!g549) & (!g550) & (g551) & (g552) & (!g42) & (g43)) + ((!g549) & (!g550) & (g551) & (g552) & (g42) & (g43)) + ((!g549) & (g550) & (!g551) & (!g552) & (g42) & (!g43)) + ((!g549) & (g550) & (!g551) & (g552) & (g42) & (!g43)) + ((!g549) & (g550) & (!g551) & (g552) & (g42) & (g43)) + ((!g549) & (g550) & (g551) & (!g552) & (!g42) & (g43)) + ((!g549) & (g550) & (g551) & (!g552) & (g42) & (!g43)) + ((!g549) & (g550) & (g551) & (g552) & (!g42) & (g43)) + ((!g549) & (g550) & (g551) & (g552) & (g42) & (!g43)) + ((!g549) & (g550) & (g551) & (g552) & (g42) & (g43)) + ((g549) & (!g550) & (!g551) & (!g552) & (!g42) & (!g43)) + ((g549) & (!g550) & (!g551) & (g552) & (!g42) & (!g43)) + ((g549) & (!g550) & (!g551) & (g552) & (g42) & (g43)) + ((g549) & (!g550) & (g551) & (!g552) & (!g42) & (!g43)) + ((g549) & (!g550) & (g551) & (!g552) & (!g42) & (g43)) + ((g549) & (!g550) & (g551) & (g552) & (!g42) & (!g43)) + ((g549) & (!g550) & (g551) & (g552) & (!g42) & (g43)) + ((g549) & (!g550) & (g551) & (g552) & (g42) & (g43)) + ((g549) & (g550) & (!g551) & (!g552) & (!g42) & (!g43)) + ((g549) & (g550) & (!g551) & (!g552) & (g42) & (!g43)) + ((g549) & (g550) & (!g551) & (g552) & (!g42) & (!g43)) + ((g549) & (g550) & (!g551) & (g552) & (g42) & (!g43)) + ((g549) & (g550) & (!g551) & (g552) & (g42) & (g43)) + ((g549) & (g550) & (g551) & (!g552) & (!g42) & (!g43)) + ((g549) & (g550) & (g551) & (!g552) & (!g42) & (g43)) + ((g549) & (g550) & (g551) & (!g552) & (g42) & (!g43)) + ((g549) & (g550) & (g551) & (g552) & (!g42) & (!g43)) + ((g549) & (g550) & (g551) & (g552) & (!g42) & (g43)) + ((g549) & (g550) & (g551) & (g552) & (g42) & (!g43)) + ((g549) & (g550) & (g551) & (g552) & (g42) & (g43)));
	assign g558 = (((!g554) & (!g555) & (!g556) & (g557) & (g42) & (g43)) + ((!g554) & (!g555) & (g556) & (!g557) & (!g42) & (g43)) + ((!g554) & (!g555) & (g556) & (g557) & (!g42) & (g43)) + ((!g554) & (!g555) & (g556) & (g557) & (g42) & (g43)) + ((!g554) & (g555) & (!g556) & (!g557) & (g42) & (!g43)) + ((!g554) & (g555) & (!g556) & (g557) & (g42) & (!g43)) + ((!g554) & (g555) & (!g556) & (g557) & (g42) & (g43)) + ((!g554) & (g555) & (g556) & (!g557) & (!g42) & (g43)) + ((!g554) & (g555) & (g556) & (!g557) & (g42) & (!g43)) + ((!g554) & (g555) & (g556) & (g557) & (!g42) & (g43)) + ((!g554) & (g555) & (g556) & (g557) & (g42) & (!g43)) + ((!g554) & (g555) & (g556) & (g557) & (g42) & (g43)) + ((g554) & (!g555) & (!g556) & (!g557) & (!g42) & (!g43)) + ((g554) & (!g555) & (!g556) & (g557) & (!g42) & (!g43)) + ((g554) & (!g555) & (!g556) & (g557) & (g42) & (g43)) + ((g554) & (!g555) & (g556) & (!g557) & (!g42) & (!g43)) + ((g554) & (!g555) & (g556) & (!g557) & (!g42) & (g43)) + ((g554) & (!g555) & (g556) & (g557) & (!g42) & (!g43)) + ((g554) & (!g555) & (g556) & (g557) & (!g42) & (g43)) + ((g554) & (!g555) & (g556) & (g557) & (g42) & (g43)) + ((g554) & (g555) & (!g556) & (!g557) & (!g42) & (!g43)) + ((g554) & (g555) & (!g556) & (!g557) & (g42) & (!g43)) + ((g554) & (g555) & (!g556) & (g557) & (!g42) & (!g43)) + ((g554) & (g555) & (!g556) & (g557) & (g42) & (!g43)) + ((g554) & (g555) & (!g556) & (g557) & (g42) & (g43)) + ((g554) & (g555) & (g556) & (!g557) & (!g42) & (!g43)) + ((g554) & (g555) & (g556) & (!g557) & (!g42) & (g43)) + ((g554) & (g555) & (g556) & (!g557) & (g42) & (!g43)) + ((g554) & (g555) & (g556) & (g557) & (!g42) & (!g43)) + ((g554) & (g555) & (g556) & (g557) & (!g42) & (g43)) + ((g554) & (g555) & (g556) & (g557) & (g42) & (!g43)) + ((g554) & (g555) & (g556) & (g557) & (g42) & (g43)));
	assign g563 = (((!g559) & (!g560) & (!g561) & (g562) & (g42) & (g43)) + ((!g559) & (!g560) & (g561) & (!g562) & (!g42) & (g43)) + ((!g559) & (!g560) & (g561) & (g562) & (!g42) & (g43)) + ((!g559) & (!g560) & (g561) & (g562) & (g42) & (g43)) + ((!g559) & (g560) & (!g561) & (!g562) & (g42) & (!g43)) + ((!g559) & (g560) & (!g561) & (g562) & (g42) & (!g43)) + ((!g559) & (g560) & (!g561) & (g562) & (g42) & (g43)) + ((!g559) & (g560) & (g561) & (!g562) & (!g42) & (g43)) + ((!g559) & (g560) & (g561) & (!g562) & (g42) & (!g43)) + ((!g559) & (g560) & (g561) & (g562) & (!g42) & (g43)) + ((!g559) & (g560) & (g561) & (g562) & (g42) & (!g43)) + ((!g559) & (g560) & (g561) & (g562) & (g42) & (g43)) + ((g559) & (!g560) & (!g561) & (!g562) & (!g42) & (!g43)) + ((g559) & (!g560) & (!g561) & (g562) & (!g42) & (!g43)) + ((g559) & (!g560) & (!g561) & (g562) & (g42) & (g43)) + ((g559) & (!g560) & (g561) & (!g562) & (!g42) & (!g43)) + ((g559) & (!g560) & (g561) & (!g562) & (!g42) & (g43)) + ((g559) & (!g560) & (g561) & (g562) & (!g42) & (!g43)) + ((g559) & (!g560) & (g561) & (g562) & (!g42) & (g43)) + ((g559) & (!g560) & (g561) & (g562) & (g42) & (g43)) + ((g559) & (g560) & (!g561) & (!g562) & (!g42) & (!g43)) + ((g559) & (g560) & (!g561) & (!g562) & (g42) & (!g43)) + ((g559) & (g560) & (!g561) & (g562) & (!g42) & (!g43)) + ((g559) & (g560) & (!g561) & (g562) & (g42) & (!g43)) + ((g559) & (g560) & (!g561) & (g562) & (g42) & (g43)) + ((g559) & (g560) & (g561) & (!g562) & (!g42) & (!g43)) + ((g559) & (g560) & (g561) & (!g562) & (!g42) & (g43)) + ((g559) & (g560) & (g561) & (!g562) & (g42) & (!g43)) + ((g559) & (g560) & (g561) & (g562) & (!g42) & (!g43)) + ((g559) & (g560) & (g561) & (g562) & (!g42) & (g43)) + ((g559) & (g560) & (g561) & (g562) & (g42) & (!g43)) + ((g559) & (g560) & (g561) & (g562) & (g42) & (g43)));
	assign g568 = (((!g564) & (!g565) & (!g566) & (g567) & (g42) & (g43)) + ((!g564) & (!g565) & (g566) & (!g567) & (!g42) & (g43)) + ((!g564) & (!g565) & (g566) & (g567) & (!g42) & (g43)) + ((!g564) & (!g565) & (g566) & (g567) & (g42) & (g43)) + ((!g564) & (g565) & (!g566) & (!g567) & (g42) & (!g43)) + ((!g564) & (g565) & (!g566) & (g567) & (g42) & (!g43)) + ((!g564) & (g565) & (!g566) & (g567) & (g42) & (g43)) + ((!g564) & (g565) & (g566) & (!g567) & (!g42) & (g43)) + ((!g564) & (g565) & (g566) & (!g567) & (g42) & (!g43)) + ((!g564) & (g565) & (g566) & (g567) & (!g42) & (g43)) + ((!g564) & (g565) & (g566) & (g567) & (g42) & (!g43)) + ((!g564) & (g565) & (g566) & (g567) & (g42) & (g43)) + ((g564) & (!g565) & (!g566) & (!g567) & (!g42) & (!g43)) + ((g564) & (!g565) & (!g566) & (g567) & (!g42) & (!g43)) + ((g564) & (!g565) & (!g566) & (g567) & (g42) & (g43)) + ((g564) & (!g565) & (g566) & (!g567) & (!g42) & (!g43)) + ((g564) & (!g565) & (g566) & (!g567) & (!g42) & (g43)) + ((g564) & (!g565) & (g566) & (g567) & (!g42) & (!g43)) + ((g564) & (!g565) & (g566) & (g567) & (!g42) & (g43)) + ((g564) & (!g565) & (g566) & (g567) & (g42) & (g43)) + ((g564) & (g565) & (!g566) & (!g567) & (!g42) & (!g43)) + ((g564) & (g565) & (!g566) & (!g567) & (g42) & (!g43)) + ((g564) & (g565) & (!g566) & (g567) & (!g42) & (!g43)) + ((g564) & (g565) & (!g566) & (g567) & (g42) & (!g43)) + ((g564) & (g565) & (!g566) & (g567) & (g42) & (g43)) + ((g564) & (g565) & (g566) & (!g567) & (!g42) & (!g43)) + ((g564) & (g565) & (g566) & (!g567) & (!g42) & (g43)) + ((g564) & (g565) & (g566) & (!g567) & (g42) & (!g43)) + ((g564) & (g565) & (g566) & (g567) & (!g42) & (!g43)) + ((g564) & (g565) & (g566) & (g567) & (!g42) & (g43)) + ((g564) & (g565) & (g566) & (g567) & (g42) & (!g43)) + ((g564) & (g565) & (g566) & (g567) & (g42) & (g43)));
	assign g569 = (((!g553) & (!g558) & (!g563) & (g568) & (g60) & (g61)) + ((!g553) & (!g558) & (g563) & (!g568) & (!g60) & (g61)) + ((!g553) & (!g558) & (g563) & (g568) & (!g60) & (g61)) + ((!g553) & (!g558) & (g563) & (g568) & (g60) & (g61)) + ((!g553) & (g558) & (!g563) & (!g568) & (g60) & (!g61)) + ((!g553) & (g558) & (!g563) & (g568) & (g60) & (!g61)) + ((!g553) & (g558) & (!g563) & (g568) & (g60) & (g61)) + ((!g553) & (g558) & (g563) & (!g568) & (!g60) & (g61)) + ((!g553) & (g558) & (g563) & (!g568) & (g60) & (!g61)) + ((!g553) & (g558) & (g563) & (g568) & (!g60) & (g61)) + ((!g553) & (g558) & (g563) & (g568) & (g60) & (!g61)) + ((!g553) & (g558) & (g563) & (g568) & (g60) & (g61)) + ((g553) & (!g558) & (!g563) & (!g568) & (!g60) & (!g61)) + ((g553) & (!g558) & (!g563) & (g568) & (!g60) & (!g61)) + ((g553) & (!g558) & (!g563) & (g568) & (g60) & (g61)) + ((g553) & (!g558) & (g563) & (!g568) & (!g60) & (!g61)) + ((g553) & (!g558) & (g563) & (!g568) & (!g60) & (g61)) + ((g553) & (!g558) & (g563) & (g568) & (!g60) & (!g61)) + ((g553) & (!g558) & (g563) & (g568) & (!g60) & (g61)) + ((g553) & (!g558) & (g563) & (g568) & (g60) & (g61)) + ((g553) & (g558) & (!g563) & (!g568) & (!g60) & (!g61)) + ((g553) & (g558) & (!g563) & (!g568) & (g60) & (!g61)) + ((g553) & (g558) & (!g563) & (g568) & (!g60) & (!g61)) + ((g553) & (g558) & (!g563) & (g568) & (g60) & (!g61)) + ((g553) & (g558) & (!g563) & (g568) & (g60) & (g61)) + ((g553) & (g558) & (g563) & (!g568) & (!g60) & (!g61)) + ((g553) & (g558) & (g563) & (!g568) & (!g60) & (g61)) + ((g553) & (g558) & (g563) & (!g568) & (g60) & (!g61)) + ((g553) & (g558) & (g563) & (g568) & (!g60) & (!g61)) + ((g553) & (g558) & (g563) & (g568) & (!g60) & (g61)) + ((g553) & (g558) & (g563) & (g568) & (g60) & (!g61)) + ((g553) & (g558) & (g563) & (g568) & (g60) & (g61)));
	assign g7256 = (((!g832) & (g1578) & (!g570)) + ((!g832) & (g1578) & (g570)) + ((g832) & (!g1578) & (g570)) + ((g832) & (g1578) & (g570)));
	assign g571 = (((!g34) & (!reset) & (!g569) & (g570)) + ((!g34) & (!reset) & (g569) & (g570)) + ((g34) & (!reset) & (g569) & (!g570)) + ((g34) & (!reset) & (g569) & (g570)));
	assign g576 = (((!g572) & (!g573) & (!g574) & (g575) & (g60) & (g61)) + ((!g572) & (!g573) & (g574) & (!g575) & (!g60) & (g61)) + ((!g572) & (!g573) & (g574) & (g575) & (!g60) & (g61)) + ((!g572) & (!g573) & (g574) & (g575) & (g60) & (g61)) + ((!g572) & (g573) & (!g574) & (!g575) & (g60) & (!g61)) + ((!g572) & (g573) & (!g574) & (g575) & (g60) & (!g61)) + ((!g572) & (g573) & (!g574) & (g575) & (g60) & (g61)) + ((!g572) & (g573) & (g574) & (!g575) & (!g60) & (g61)) + ((!g572) & (g573) & (g574) & (!g575) & (g60) & (!g61)) + ((!g572) & (g573) & (g574) & (g575) & (!g60) & (g61)) + ((!g572) & (g573) & (g574) & (g575) & (g60) & (!g61)) + ((!g572) & (g573) & (g574) & (g575) & (g60) & (g61)) + ((g572) & (!g573) & (!g574) & (!g575) & (!g60) & (!g61)) + ((g572) & (!g573) & (!g574) & (g575) & (!g60) & (!g61)) + ((g572) & (!g573) & (!g574) & (g575) & (g60) & (g61)) + ((g572) & (!g573) & (g574) & (!g575) & (!g60) & (!g61)) + ((g572) & (!g573) & (g574) & (!g575) & (!g60) & (g61)) + ((g572) & (!g573) & (g574) & (g575) & (!g60) & (!g61)) + ((g572) & (!g573) & (g574) & (g575) & (!g60) & (g61)) + ((g572) & (!g573) & (g574) & (g575) & (g60) & (g61)) + ((g572) & (g573) & (!g574) & (!g575) & (!g60) & (!g61)) + ((g572) & (g573) & (!g574) & (!g575) & (g60) & (!g61)) + ((g572) & (g573) & (!g574) & (g575) & (!g60) & (!g61)) + ((g572) & (g573) & (!g574) & (g575) & (g60) & (!g61)) + ((g572) & (g573) & (!g574) & (g575) & (g60) & (g61)) + ((g572) & (g573) & (g574) & (!g575) & (!g60) & (!g61)) + ((g572) & (g573) & (g574) & (!g575) & (!g60) & (g61)) + ((g572) & (g573) & (g574) & (!g575) & (g60) & (!g61)) + ((g572) & (g573) & (g574) & (g575) & (!g60) & (!g61)) + ((g572) & (g573) & (g574) & (g575) & (!g60) & (g61)) + ((g572) & (g573) & (g574) & (g575) & (g60) & (!g61)) + ((g572) & (g573) & (g574) & (g575) & (g60) & (g61)));
	assign g581 = (((!g577) & (!g578) & (!g579) & (g580) & (g60) & (g61)) + ((!g577) & (!g578) & (g579) & (!g580) & (!g60) & (g61)) + ((!g577) & (!g578) & (g579) & (g580) & (!g60) & (g61)) + ((!g577) & (!g578) & (g579) & (g580) & (g60) & (g61)) + ((!g577) & (g578) & (!g579) & (!g580) & (g60) & (!g61)) + ((!g577) & (g578) & (!g579) & (g580) & (g60) & (!g61)) + ((!g577) & (g578) & (!g579) & (g580) & (g60) & (g61)) + ((!g577) & (g578) & (g579) & (!g580) & (!g60) & (g61)) + ((!g577) & (g578) & (g579) & (!g580) & (g60) & (!g61)) + ((!g577) & (g578) & (g579) & (g580) & (!g60) & (g61)) + ((!g577) & (g578) & (g579) & (g580) & (g60) & (!g61)) + ((!g577) & (g578) & (g579) & (g580) & (g60) & (g61)) + ((g577) & (!g578) & (!g579) & (!g580) & (!g60) & (!g61)) + ((g577) & (!g578) & (!g579) & (g580) & (!g60) & (!g61)) + ((g577) & (!g578) & (!g579) & (g580) & (g60) & (g61)) + ((g577) & (!g578) & (g579) & (!g580) & (!g60) & (!g61)) + ((g577) & (!g578) & (g579) & (!g580) & (!g60) & (g61)) + ((g577) & (!g578) & (g579) & (g580) & (!g60) & (!g61)) + ((g577) & (!g578) & (g579) & (g580) & (!g60) & (g61)) + ((g577) & (!g578) & (g579) & (g580) & (g60) & (g61)) + ((g577) & (g578) & (!g579) & (!g580) & (!g60) & (!g61)) + ((g577) & (g578) & (!g579) & (!g580) & (g60) & (!g61)) + ((g577) & (g578) & (!g579) & (g580) & (!g60) & (!g61)) + ((g577) & (g578) & (!g579) & (g580) & (g60) & (!g61)) + ((g577) & (g578) & (!g579) & (g580) & (g60) & (g61)) + ((g577) & (g578) & (g579) & (!g580) & (!g60) & (!g61)) + ((g577) & (g578) & (g579) & (!g580) & (!g60) & (g61)) + ((g577) & (g578) & (g579) & (!g580) & (g60) & (!g61)) + ((g577) & (g578) & (g579) & (g580) & (!g60) & (!g61)) + ((g577) & (g578) & (g579) & (g580) & (!g60) & (g61)) + ((g577) & (g578) & (g579) & (g580) & (g60) & (!g61)) + ((g577) & (g578) & (g579) & (g580) & (g60) & (g61)));
	assign g586 = (((!g582) & (!g583) & (!g584) & (g585) & (g60) & (g61)) + ((!g582) & (!g583) & (g584) & (!g585) & (!g60) & (g61)) + ((!g582) & (!g583) & (g584) & (g585) & (!g60) & (g61)) + ((!g582) & (!g583) & (g584) & (g585) & (g60) & (g61)) + ((!g582) & (g583) & (!g584) & (!g585) & (g60) & (!g61)) + ((!g582) & (g583) & (!g584) & (g585) & (g60) & (!g61)) + ((!g582) & (g583) & (!g584) & (g585) & (g60) & (g61)) + ((!g582) & (g583) & (g584) & (!g585) & (!g60) & (g61)) + ((!g582) & (g583) & (g584) & (!g585) & (g60) & (!g61)) + ((!g582) & (g583) & (g584) & (g585) & (!g60) & (g61)) + ((!g582) & (g583) & (g584) & (g585) & (g60) & (!g61)) + ((!g582) & (g583) & (g584) & (g585) & (g60) & (g61)) + ((g582) & (!g583) & (!g584) & (!g585) & (!g60) & (!g61)) + ((g582) & (!g583) & (!g584) & (g585) & (!g60) & (!g61)) + ((g582) & (!g583) & (!g584) & (g585) & (g60) & (g61)) + ((g582) & (!g583) & (g584) & (!g585) & (!g60) & (!g61)) + ((g582) & (!g583) & (g584) & (!g585) & (!g60) & (g61)) + ((g582) & (!g583) & (g584) & (g585) & (!g60) & (!g61)) + ((g582) & (!g583) & (g584) & (g585) & (!g60) & (g61)) + ((g582) & (!g583) & (g584) & (g585) & (g60) & (g61)) + ((g582) & (g583) & (!g584) & (!g585) & (!g60) & (!g61)) + ((g582) & (g583) & (!g584) & (!g585) & (g60) & (!g61)) + ((g582) & (g583) & (!g584) & (g585) & (!g60) & (!g61)) + ((g582) & (g583) & (!g584) & (g585) & (g60) & (!g61)) + ((g582) & (g583) & (!g584) & (g585) & (g60) & (g61)) + ((g582) & (g583) & (g584) & (!g585) & (!g60) & (!g61)) + ((g582) & (g583) & (g584) & (!g585) & (!g60) & (g61)) + ((g582) & (g583) & (g584) & (!g585) & (g60) & (!g61)) + ((g582) & (g583) & (g584) & (g585) & (!g60) & (!g61)) + ((g582) & (g583) & (g584) & (g585) & (!g60) & (g61)) + ((g582) & (g583) & (g584) & (g585) & (g60) & (!g61)) + ((g582) & (g583) & (g584) & (g585) & (g60) & (g61)));
	assign g591 = (((!g587) & (!g588) & (!g589) & (g590) & (g60) & (g61)) + ((!g587) & (!g588) & (g589) & (!g590) & (!g60) & (g61)) + ((!g587) & (!g588) & (g589) & (g590) & (!g60) & (g61)) + ((!g587) & (!g588) & (g589) & (g590) & (g60) & (g61)) + ((!g587) & (g588) & (!g589) & (!g590) & (g60) & (!g61)) + ((!g587) & (g588) & (!g589) & (g590) & (g60) & (!g61)) + ((!g587) & (g588) & (!g589) & (g590) & (g60) & (g61)) + ((!g587) & (g588) & (g589) & (!g590) & (!g60) & (g61)) + ((!g587) & (g588) & (g589) & (!g590) & (g60) & (!g61)) + ((!g587) & (g588) & (g589) & (g590) & (!g60) & (g61)) + ((!g587) & (g588) & (g589) & (g590) & (g60) & (!g61)) + ((!g587) & (g588) & (g589) & (g590) & (g60) & (g61)) + ((g587) & (!g588) & (!g589) & (!g590) & (!g60) & (!g61)) + ((g587) & (!g588) & (!g589) & (g590) & (!g60) & (!g61)) + ((g587) & (!g588) & (!g589) & (g590) & (g60) & (g61)) + ((g587) & (!g588) & (g589) & (!g590) & (!g60) & (!g61)) + ((g587) & (!g588) & (g589) & (!g590) & (!g60) & (g61)) + ((g587) & (!g588) & (g589) & (g590) & (!g60) & (!g61)) + ((g587) & (!g588) & (g589) & (g590) & (!g60) & (g61)) + ((g587) & (!g588) & (g589) & (g590) & (g60) & (g61)) + ((g587) & (g588) & (!g589) & (!g590) & (!g60) & (!g61)) + ((g587) & (g588) & (!g589) & (!g590) & (g60) & (!g61)) + ((g587) & (g588) & (!g589) & (g590) & (!g60) & (!g61)) + ((g587) & (g588) & (!g589) & (g590) & (g60) & (!g61)) + ((g587) & (g588) & (!g589) & (g590) & (g60) & (g61)) + ((g587) & (g588) & (g589) & (!g590) & (!g60) & (!g61)) + ((g587) & (g588) & (g589) & (!g590) & (!g60) & (g61)) + ((g587) & (g588) & (g589) & (!g590) & (g60) & (!g61)) + ((g587) & (g588) & (g589) & (g590) & (!g60) & (!g61)) + ((g587) & (g588) & (g589) & (g590) & (!g60) & (g61)) + ((g587) & (g588) & (g589) & (g590) & (g60) & (!g61)) + ((g587) & (g588) & (g589) & (g590) & (g60) & (g61)));
	assign g592 = (((!g576) & (!g581) & (!g586) & (g591) & (g42) & (g43)) + ((!g576) & (!g581) & (g586) & (!g591) & (!g42) & (g43)) + ((!g576) & (!g581) & (g586) & (g591) & (!g42) & (g43)) + ((!g576) & (!g581) & (g586) & (g591) & (g42) & (g43)) + ((!g576) & (g581) & (!g586) & (!g591) & (g42) & (!g43)) + ((!g576) & (g581) & (!g586) & (g591) & (g42) & (!g43)) + ((!g576) & (g581) & (!g586) & (g591) & (g42) & (g43)) + ((!g576) & (g581) & (g586) & (!g591) & (!g42) & (g43)) + ((!g576) & (g581) & (g586) & (!g591) & (g42) & (!g43)) + ((!g576) & (g581) & (g586) & (g591) & (!g42) & (g43)) + ((!g576) & (g581) & (g586) & (g591) & (g42) & (!g43)) + ((!g576) & (g581) & (g586) & (g591) & (g42) & (g43)) + ((g576) & (!g581) & (!g586) & (!g591) & (!g42) & (!g43)) + ((g576) & (!g581) & (!g586) & (g591) & (!g42) & (!g43)) + ((g576) & (!g581) & (!g586) & (g591) & (g42) & (g43)) + ((g576) & (!g581) & (g586) & (!g591) & (!g42) & (!g43)) + ((g576) & (!g581) & (g586) & (!g591) & (!g42) & (g43)) + ((g576) & (!g581) & (g586) & (g591) & (!g42) & (!g43)) + ((g576) & (!g581) & (g586) & (g591) & (!g42) & (g43)) + ((g576) & (!g581) & (g586) & (g591) & (g42) & (g43)) + ((g576) & (g581) & (!g586) & (!g591) & (!g42) & (!g43)) + ((g576) & (g581) & (!g586) & (!g591) & (g42) & (!g43)) + ((g576) & (g581) & (!g586) & (g591) & (!g42) & (!g43)) + ((g576) & (g581) & (!g586) & (g591) & (g42) & (!g43)) + ((g576) & (g581) & (!g586) & (g591) & (g42) & (g43)) + ((g576) & (g581) & (g586) & (!g591) & (!g42) & (!g43)) + ((g576) & (g581) & (g586) & (!g591) & (!g42) & (g43)) + ((g576) & (g581) & (g586) & (!g591) & (g42) & (!g43)) + ((g576) & (g581) & (g586) & (g591) & (!g42) & (!g43)) + ((g576) & (g581) & (g586) & (g591) & (!g42) & (g43)) + ((g576) & (g581) & (g586) & (g591) & (g42) & (!g43)) + ((g576) & (g581) & (g586) & (g591) & (g42) & (g43)));
	assign g7257 = (((!g832) & (g1612) & (!g593)) + ((!g832) & (g1612) & (g593)) + ((g832) & (!g1612) & (g593)) + ((g832) & (g1612) & (g593)));
	assign g594 = (((!g34) & (!reset) & (!g592) & (g593)) + ((!g34) & (!reset) & (g592) & (g593)) + ((g34) & (!reset) & (g592) & (!g593)) + ((g34) & (!reset) & (g592) & (g593)));
	assign g599 = (((!g595) & (!g596) & (!g597) & (g598) & (g42) & (g43)) + ((!g595) & (!g596) & (g597) & (!g598) & (!g42) & (g43)) + ((!g595) & (!g596) & (g597) & (g598) & (!g42) & (g43)) + ((!g595) & (!g596) & (g597) & (g598) & (g42) & (g43)) + ((!g595) & (g596) & (!g597) & (!g598) & (g42) & (!g43)) + ((!g595) & (g596) & (!g597) & (g598) & (g42) & (!g43)) + ((!g595) & (g596) & (!g597) & (g598) & (g42) & (g43)) + ((!g595) & (g596) & (g597) & (!g598) & (!g42) & (g43)) + ((!g595) & (g596) & (g597) & (!g598) & (g42) & (!g43)) + ((!g595) & (g596) & (g597) & (g598) & (!g42) & (g43)) + ((!g595) & (g596) & (g597) & (g598) & (g42) & (!g43)) + ((!g595) & (g596) & (g597) & (g598) & (g42) & (g43)) + ((g595) & (!g596) & (!g597) & (!g598) & (!g42) & (!g43)) + ((g595) & (!g596) & (!g597) & (g598) & (!g42) & (!g43)) + ((g595) & (!g596) & (!g597) & (g598) & (g42) & (g43)) + ((g595) & (!g596) & (g597) & (!g598) & (!g42) & (!g43)) + ((g595) & (!g596) & (g597) & (!g598) & (!g42) & (g43)) + ((g595) & (!g596) & (g597) & (g598) & (!g42) & (!g43)) + ((g595) & (!g596) & (g597) & (g598) & (!g42) & (g43)) + ((g595) & (!g596) & (g597) & (g598) & (g42) & (g43)) + ((g595) & (g596) & (!g597) & (!g598) & (!g42) & (!g43)) + ((g595) & (g596) & (!g597) & (!g598) & (g42) & (!g43)) + ((g595) & (g596) & (!g597) & (g598) & (!g42) & (!g43)) + ((g595) & (g596) & (!g597) & (g598) & (g42) & (!g43)) + ((g595) & (g596) & (!g597) & (g598) & (g42) & (g43)) + ((g595) & (g596) & (g597) & (!g598) & (!g42) & (!g43)) + ((g595) & (g596) & (g597) & (!g598) & (!g42) & (g43)) + ((g595) & (g596) & (g597) & (!g598) & (g42) & (!g43)) + ((g595) & (g596) & (g597) & (g598) & (!g42) & (!g43)) + ((g595) & (g596) & (g597) & (g598) & (!g42) & (g43)) + ((g595) & (g596) & (g597) & (g598) & (g42) & (!g43)) + ((g595) & (g596) & (g597) & (g598) & (g42) & (g43)));
	assign g604 = (((!g600) & (!g601) & (!g602) & (g603) & (g42) & (g43)) + ((!g600) & (!g601) & (g602) & (!g603) & (!g42) & (g43)) + ((!g600) & (!g601) & (g602) & (g603) & (!g42) & (g43)) + ((!g600) & (!g601) & (g602) & (g603) & (g42) & (g43)) + ((!g600) & (g601) & (!g602) & (!g603) & (g42) & (!g43)) + ((!g600) & (g601) & (!g602) & (g603) & (g42) & (!g43)) + ((!g600) & (g601) & (!g602) & (g603) & (g42) & (g43)) + ((!g600) & (g601) & (g602) & (!g603) & (!g42) & (g43)) + ((!g600) & (g601) & (g602) & (!g603) & (g42) & (!g43)) + ((!g600) & (g601) & (g602) & (g603) & (!g42) & (g43)) + ((!g600) & (g601) & (g602) & (g603) & (g42) & (!g43)) + ((!g600) & (g601) & (g602) & (g603) & (g42) & (g43)) + ((g600) & (!g601) & (!g602) & (!g603) & (!g42) & (!g43)) + ((g600) & (!g601) & (!g602) & (g603) & (!g42) & (!g43)) + ((g600) & (!g601) & (!g602) & (g603) & (g42) & (g43)) + ((g600) & (!g601) & (g602) & (!g603) & (!g42) & (!g43)) + ((g600) & (!g601) & (g602) & (!g603) & (!g42) & (g43)) + ((g600) & (!g601) & (g602) & (g603) & (!g42) & (!g43)) + ((g600) & (!g601) & (g602) & (g603) & (!g42) & (g43)) + ((g600) & (!g601) & (g602) & (g603) & (g42) & (g43)) + ((g600) & (g601) & (!g602) & (!g603) & (!g42) & (!g43)) + ((g600) & (g601) & (!g602) & (!g603) & (g42) & (!g43)) + ((g600) & (g601) & (!g602) & (g603) & (!g42) & (!g43)) + ((g600) & (g601) & (!g602) & (g603) & (g42) & (!g43)) + ((g600) & (g601) & (!g602) & (g603) & (g42) & (g43)) + ((g600) & (g601) & (g602) & (!g603) & (!g42) & (!g43)) + ((g600) & (g601) & (g602) & (!g603) & (!g42) & (g43)) + ((g600) & (g601) & (g602) & (!g603) & (g42) & (!g43)) + ((g600) & (g601) & (g602) & (g603) & (!g42) & (!g43)) + ((g600) & (g601) & (g602) & (g603) & (!g42) & (g43)) + ((g600) & (g601) & (g602) & (g603) & (g42) & (!g43)) + ((g600) & (g601) & (g602) & (g603) & (g42) & (g43)));
	assign g609 = (((!g605) & (!g606) & (!g607) & (g608) & (g42) & (g43)) + ((!g605) & (!g606) & (g607) & (!g608) & (!g42) & (g43)) + ((!g605) & (!g606) & (g607) & (g608) & (!g42) & (g43)) + ((!g605) & (!g606) & (g607) & (g608) & (g42) & (g43)) + ((!g605) & (g606) & (!g607) & (!g608) & (g42) & (!g43)) + ((!g605) & (g606) & (!g607) & (g608) & (g42) & (!g43)) + ((!g605) & (g606) & (!g607) & (g608) & (g42) & (g43)) + ((!g605) & (g606) & (g607) & (!g608) & (!g42) & (g43)) + ((!g605) & (g606) & (g607) & (!g608) & (g42) & (!g43)) + ((!g605) & (g606) & (g607) & (g608) & (!g42) & (g43)) + ((!g605) & (g606) & (g607) & (g608) & (g42) & (!g43)) + ((!g605) & (g606) & (g607) & (g608) & (g42) & (g43)) + ((g605) & (!g606) & (!g607) & (!g608) & (!g42) & (!g43)) + ((g605) & (!g606) & (!g607) & (g608) & (!g42) & (!g43)) + ((g605) & (!g606) & (!g607) & (g608) & (g42) & (g43)) + ((g605) & (!g606) & (g607) & (!g608) & (!g42) & (!g43)) + ((g605) & (!g606) & (g607) & (!g608) & (!g42) & (g43)) + ((g605) & (!g606) & (g607) & (g608) & (!g42) & (!g43)) + ((g605) & (!g606) & (g607) & (g608) & (!g42) & (g43)) + ((g605) & (!g606) & (g607) & (g608) & (g42) & (g43)) + ((g605) & (g606) & (!g607) & (!g608) & (!g42) & (!g43)) + ((g605) & (g606) & (!g607) & (!g608) & (g42) & (!g43)) + ((g605) & (g606) & (!g607) & (g608) & (!g42) & (!g43)) + ((g605) & (g606) & (!g607) & (g608) & (g42) & (!g43)) + ((g605) & (g606) & (!g607) & (g608) & (g42) & (g43)) + ((g605) & (g606) & (g607) & (!g608) & (!g42) & (!g43)) + ((g605) & (g606) & (g607) & (!g608) & (!g42) & (g43)) + ((g605) & (g606) & (g607) & (!g608) & (g42) & (!g43)) + ((g605) & (g606) & (g607) & (g608) & (!g42) & (!g43)) + ((g605) & (g606) & (g607) & (g608) & (!g42) & (g43)) + ((g605) & (g606) & (g607) & (g608) & (g42) & (!g43)) + ((g605) & (g606) & (g607) & (g608) & (g42) & (g43)));
	assign g614 = (((!g610) & (!g611) & (!g612) & (g613) & (g42) & (g43)) + ((!g610) & (!g611) & (g612) & (!g613) & (!g42) & (g43)) + ((!g610) & (!g611) & (g612) & (g613) & (!g42) & (g43)) + ((!g610) & (!g611) & (g612) & (g613) & (g42) & (g43)) + ((!g610) & (g611) & (!g612) & (!g613) & (g42) & (!g43)) + ((!g610) & (g611) & (!g612) & (g613) & (g42) & (!g43)) + ((!g610) & (g611) & (!g612) & (g613) & (g42) & (g43)) + ((!g610) & (g611) & (g612) & (!g613) & (!g42) & (g43)) + ((!g610) & (g611) & (g612) & (!g613) & (g42) & (!g43)) + ((!g610) & (g611) & (g612) & (g613) & (!g42) & (g43)) + ((!g610) & (g611) & (g612) & (g613) & (g42) & (!g43)) + ((!g610) & (g611) & (g612) & (g613) & (g42) & (g43)) + ((g610) & (!g611) & (!g612) & (!g613) & (!g42) & (!g43)) + ((g610) & (!g611) & (!g612) & (g613) & (!g42) & (!g43)) + ((g610) & (!g611) & (!g612) & (g613) & (g42) & (g43)) + ((g610) & (!g611) & (g612) & (!g613) & (!g42) & (!g43)) + ((g610) & (!g611) & (g612) & (!g613) & (!g42) & (g43)) + ((g610) & (!g611) & (g612) & (g613) & (!g42) & (!g43)) + ((g610) & (!g611) & (g612) & (g613) & (!g42) & (g43)) + ((g610) & (!g611) & (g612) & (g613) & (g42) & (g43)) + ((g610) & (g611) & (!g612) & (!g613) & (!g42) & (!g43)) + ((g610) & (g611) & (!g612) & (!g613) & (g42) & (!g43)) + ((g610) & (g611) & (!g612) & (g613) & (!g42) & (!g43)) + ((g610) & (g611) & (!g612) & (g613) & (g42) & (!g43)) + ((g610) & (g611) & (!g612) & (g613) & (g42) & (g43)) + ((g610) & (g611) & (g612) & (!g613) & (!g42) & (!g43)) + ((g610) & (g611) & (g612) & (!g613) & (!g42) & (g43)) + ((g610) & (g611) & (g612) & (!g613) & (g42) & (!g43)) + ((g610) & (g611) & (g612) & (g613) & (!g42) & (!g43)) + ((g610) & (g611) & (g612) & (g613) & (!g42) & (g43)) + ((g610) & (g611) & (g612) & (g613) & (g42) & (!g43)) + ((g610) & (g611) & (g612) & (g613) & (g42) & (g43)));
	assign g615 = (((!g599) & (!g604) & (!g609) & (g614) & (g60) & (g61)) + ((!g599) & (!g604) & (g609) & (!g614) & (!g60) & (g61)) + ((!g599) & (!g604) & (g609) & (g614) & (!g60) & (g61)) + ((!g599) & (!g604) & (g609) & (g614) & (g60) & (g61)) + ((!g599) & (g604) & (!g609) & (!g614) & (g60) & (!g61)) + ((!g599) & (g604) & (!g609) & (g614) & (g60) & (!g61)) + ((!g599) & (g604) & (!g609) & (g614) & (g60) & (g61)) + ((!g599) & (g604) & (g609) & (!g614) & (!g60) & (g61)) + ((!g599) & (g604) & (g609) & (!g614) & (g60) & (!g61)) + ((!g599) & (g604) & (g609) & (g614) & (!g60) & (g61)) + ((!g599) & (g604) & (g609) & (g614) & (g60) & (!g61)) + ((!g599) & (g604) & (g609) & (g614) & (g60) & (g61)) + ((g599) & (!g604) & (!g609) & (!g614) & (!g60) & (!g61)) + ((g599) & (!g604) & (!g609) & (g614) & (!g60) & (!g61)) + ((g599) & (!g604) & (!g609) & (g614) & (g60) & (g61)) + ((g599) & (!g604) & (g609) & (!g614) & (!g60) & (!g61)) + ((g599) & (!g604) & (g609) & (!g614) & (!g60) & (g61)) + ((g599) & (!g604) & (g609) & (g614) & (!g60) & (!g61)) + ((g599) & (!g604) & (g609) & (g614) & (!g60) & (g61)) + ((g599) & (!g604) & (g609) & (g614) & (g60) & (g61)) + ((g599) & (g604) & (!g609) & (!g614) & (!g60) & (!g61)) + ((g599) & (g604) & (!g609) & (!g614) & (g60) & (!g61)) + ((g599) & (g604) & (!g609) & (g614) & (!g60) & (!g61)) + ((g599) & (g604) & (!g609) & (g614) & (g60) & (!g61)) + ((g599) & (g604) & (!g609) & (g614) & (g60) & (g61)) + ((g599) & (g604) & (g609) & (!g614) & (!g60) & (!g61)) + ((g599) & (g604) & (g609) & (!g614) & (!g60) & (g61)) + ((g599) & (g604) & (g609) & (!g614) & (g60) & (!g61)) + ((g599) & (g604) & (g609) & (g614) & (!g60) & (!g61)) + ((g599) & (g604) & (g609) & (g614) & (!g60) & (g61)) + ((g599) & (g604) & (g609) & (g614) & (g60) & (!g61)) + ((g599) & (g604) & (g609) & (g614) & (g60) & (g61)));
	assign g7258 = (((!g832) & (g1645) & (!g616)) + ((!g832) & (g1645) & (g616)) + ((g832) & (!g1645) & (g616)) + ((g832) & (g1645) & (g616)));
	assign g617 = (((!g34) & (!reset) & (!g615) & (g616)) + ((!g34) & (!reset) & (g615) & (g616)) + ((g34) & (!reset) & (g615) & (!g616)) + ((g34) & (!reset) & (g615) & (g616)));
	assign g622 = (((!g618) & (!g619) & (!g620) & (g621) & (g60) & (g61)) + ((!g618) & (!g619) & (g620) & (!g621) & (!g60) & (g61)) + ((!g618) & (!g619) & (g620) & (g621) & (!g60) & (g61)) + ((!g618) & (!g619) & (g620) & (g621) & (g60) & (g61)) + ((!g618) & (g619) & (!g620) & (!g621) & (g60) & (!g61)) + ((!g618) & (g619) & (!g620) & (g621) & (g60) & (!g61)) + ((!g618) & (g619) & (!g620) & (g621) & (g60) & (g61)) + ((!g618) & (g619) & (g620) & (!g621) & (!g60) & (g61)) + ((!g618) & (g619) & (g620) & (!g621) & (g60) & (!g61)) + ((!g618) & (g619) & (g620) & (g621) & (!g60) & (g61)) + ((!g618) & (g619) & (g620) & (g621) & (g60) & (!g61)) + ((!g618) & (g619) & (g620) & (g621) & (g60) & (g61)) + ((g618) & (!g619) & (!g620) & (!g621) & (!g60) & (!g61)) + ((g618) & (!g619) & (!g620) & (g621) & (!g60) & (!g61)) + ((g618) & (!g619) & (!g620) & (g621) & (g60) & (g61)) + ((g618) & (!g619) & (g620) & (!g621) & (!g60) & (!g61)) + ((g618) & (!g619) & (g620) & (!g621) & (!g60) & (g61)) + ((g618) & (!g619) & (g620) & (g621) & (!g60) & (!g61)) + ((g618) & (!g619) & (g620) & (g621) & (!g60) & (g61)) + ((g618) & (!g619) & (g620) & (g621) & (g60) & (g61)) + ((g618) & (g619) & (!g620) & (!g621) & (!g60) & (!g61)) + ((g618) & (g619) & (!g620) & (!g621) & (g60) & (!g61)) + ((g618) & (g619) & (!g620) & (g621) & (!g60) & (!g61)) + ((g618) & (g619) & (!g620) & (g621) & (g60) & (!g61)) + ((g618) & (g619) & (!g620) & (g621) & (g60) & (g61)) + ((g618) & (g619) & (g620) & (!g621) & (!g60) & (!g61)) + ((g618) & (g619) & (g620) & (!g621) & (!g60) & (g61)) + ((g618) & (g619) & (g620) & (!g621) & (g60) & (!g61)) + ((g618) & (g619) & (g620) & (g621) & (!g60) & (!g61)) + ((g618) & (g619) & (g620) & (g621) & (!g60) & (g61)) + ((g618) & (g619) & (g620) & (g621) & (g60) & (!g61)) + ((g618) & (g619) & (g620) & (g621) & (g60) & (g61)));
	assign g627 = (((!g623) & (!g624) & (!g625) & (g626) & (g60) & (g61)) + ((!g623) & (!g624) & (g625) & (!g626) & (!g60) & (g61)) + ((!g623) & (!g624) & (g625) & (g626) & (!g60) & (g61)) + ((!g623) & (!g624) & (g625) & (g626) & (g60) & (g61)) + ((!g623) & (g624) & (!g625) & (!g626) & (g60) & (!g61)) + ((!g623) & (g624) & (!g625) & (g626) & (g60) & (!g61)) + ((!g623) & (g624) & (!g625) & (g626) & (g60) & (g61)) + ((!g623) & (g624) & (g625) & (!g626) & (!g60) & (g61)) + ((!g623) & (g624) & (g625) & (!g626) & (g60) & (!g61)) + ((!g623) & (g624) & (g625) & (g626) & (!g60) & (g61)) + ((!g623) & (g624) & (g625) & (g626) & (g60) & (!g61)) + ((!g623) & (g624) & (g625) & (g626) & (g60) & (g61)) + ((g623) & (!g624) & (!g625) & (!g626) & (!g60) & (!g61)) + ((g623) & (!g624) & (!g625) & (g626) & (!g60) & (!g61)) + ((g623) & (!g624) & (!g625) & (g626) & (g60) & (g61)) + ((g623) & (!g624) & (g625) & (!g626) & (!g60) & (!g61)) + ((g623) & (!g624) & (g625) & (!g626) & (!g60) & (g61)) + ((g623) & (!g624) & (g625) & (g626) & (!g60) & (!g61)) + ((g623) & (!g624) & (g625) & (g626) & (!g60) & (g61)) + ((g623) & (!g624) & (g625) & (g626) & (g60) & (g61)) + ((g623) & (g624) & (!g625) & (!g626) & (!g60) & (!g61)) + ((g623) & (g624) & (!g625) & (!g626) & (g60) & (!g61)) + ((g623) & (g624) & (!g625) & (g626) & (!g60) & (!g61)) + ((g623) & (g624) & (!g625) & (g626) & (g60) & (!g61)) + ((g623) & (g624) & (!g625) & (g626) & (g60) & (g61)) + ((g623) & (g624) & (g625) & (!g626) & (!g60) & (!g61)) + ((g623) & (g624) & (g625) & (!g626) & (!g60) & (g61)) + ((g623) & (g624) & (g625) & (!g626) & (g60) & (!g61)) + ((g623) & (g624) & (g625) & (g626) & (!g60) & (!g61)) + ((g623) & (g624) & (g625) & (g626) & (!g60) & (g61)) + ((g623) & (g624) & (g625) & (g626) & (g60) & (!g61)) + ((g623) & (g624) & (g625) & (g626) & (g60) & (g61)));
	assign g632 = (((!g628) & (!g629) & (!g630) & (g631) & (g60) & (g61)) + ((!g628) & (!g629) & (g630) & (!g631) & (!g60) & (g61)) + ((!g628) & (!g629) & (g630) & (g631) & (!g60) & (g61)) + ((!g628) & (!g629) & (g630) & (g631) & (g60) & (g61)) + ((!g628) & (g629) & (!g630) & (!g631) & (g60) & (!g61)) + ((!g628) & (g629) & (!g630) & (g631) & (g60) & (!g61)) + ((!g628) & (g629) & (!g630) & (g631) & (g60) & (g61)) + ((!g628) & (g629) & (g630) & (!g631) & (!g60) & (g61)) + ((!g628) & (g629) & (g630) & (!g631) & (g60) & (!g61)) + ((!g628) & (g629) & (g630) & (g631) & (!g60) & (g61)) + ((!g628) & (g629) & (g630) & (g631) & (g60) & (!g61)) + ((!g628) & (g629) & (g630) & (g631) & (g60) & (g61)) + ((g628) & (!g629) & (!g630) & (!g631) & (!g60) & (!g61)) + ((g628) & (!g629) & (!g630) & (g631) & (!g60) & (!g61)) + ((g628) & (!g629) & (!g630) & (g631) & (g60) & (g61)) + ((g628) & (!g629) & (g630) & (!g631) & (!g60) & (!g61)) + ((g628) & (!g629) & (g630) & (!g631) & (!g60) & (g61)) + ((g628) & (!g629) & (g630) & (g631) & (!g60) & (!g61)) + ((g628) & (!g629) & (g630) & (g631) & (!g60) & (g61)) + ((g628) & (!g629) & (g630) & (g631) & (g60) & (g61)) + ((g628) & (g629) & (!g630) & (!g631) & (!g60) & (!g61)) + ((g628) & (g629) & (!g630) & (!g631) & (g60) & (!g61)) + ((g628) & (g629) & (!g630) & (g631) & (!g60) & (!g61)) + ((g628) & (g629) & (!g630) & (g631) & (g60) & (!g61)) + ((g628) & (g629) & (!g630) & (g631) & (g60) & (g61)) + ((g628) & (g629) & (g630) & (!g631) & (!g60) & (!g61)) + ((g628) & (g629) & (g630) & (!g631) & (!g60) & (g61)) + ((g628) & (g629) & (g630) & (!g631) & (g60) & (!g61)) + ((g628) & (g629) & (g630) & (g631) & (!g60) & (!g61)) + ((g628) & (g629) & (g630) & (g631) & (!g60) & (g61)) + ((g628) & (g629) & (g630) & (g631) & (g60) & (!g61)) + ((g628) & (g629) & (g630) & (g631) & (g60) & (g61)));
	assign g637 = (((!g633) & (!g634) & (!g635) & (g636) & (g60) & (g61)) + ((!g633) & (!g634) & (g635) & (!g636) & (!g60) & (g61)) + ((!g633) & (!g634) & (g635) & (g636) & (!g60) & (g61)) + ((!g633) & (!g634) & (g635) & (g636) & (g60) & (g61)) + ((!g633) & (g634) & (!g635) & (!g636) & (g60) & (!g61)) + ((!g633) & (g634) & (!g635) & (g636) & (g60) & (!g61)) + ((!g633) & (g634) & (!g635) & (g636) & (g60) & (g61)) + ((!g633) & (g634) & (g635) & (!g636) & (!g60) & (g61)) + ((!g633) & (g634) & (g635) & (!g636) & (g60) & (!g61)) + ((!g633) & (g634) & (g635) & (g636) & (!g60) & (g61)) + ((!g633) & (g634) & (g635) & (g636) & (g60) & (!g61)) + ((!g633) & (g634) & (g635) & (g636) & (g60) & (g61)) + ((g633) & (!g634) & (!g635) & (!g636) & (!g60) & (!g61)) + ((g633) & (!g634) & (!g635) & (g636) & (!g60) & (!g61)) + ((g633) & (!g634) & (!g635) & (g636) & (g60) & (g61)) + ((g633) & (!g634) & (g635) & (!g636) & (!g60) & (!g61)) + ((g633) & (!g634) & (g635) & (!g636) & (!g60) & (g61)) + ((g633) & (!g634) & (g635) & (g636) & (!g60) & (!g61)) + ((g633) & (!g634) & (g635) & (g636) & (!g60) & (g61)) + ((g633) & (!g634) & (g635) & (g636) & (g60) & (g61)) + ((g633) & (g634) & (!g635) & (!g636) & (!g60) & (!g61)) + ((g633) & (g634) & (!g635) & (!g636) & (g60) & (!g61)) + ((g633) & (g634) & (!g635) & (g636) & (!g60) & (!g61)) + ((g633) & (g634) & (!g635) & (g636) & (g60) & (!g61)) + ((g633) & (g634) & (!g635) & (g636) & (g60) & (g61)) + ((g633) & (g634) & (g635) & (!g636) & (!g60) & (!g61)) + ((g633) & (g634) & (g635) & (!g636) & (!g60) & (g61)) + ((g633) & (g634) & (g635) & (!g636) & (g60) & (!g61)) + ((g633) & (g634) & (g635) & (g636) & (!g60) & (!g61)) + ((g633) & (g634) & (g635) & (g636) & (!g60) & (g61)) + ((g633) & (g634) & (g635) & (g636) & (g60) & (!g61)) + ((g633) & (g634) & (g635) & (g636) & (g60) & (g61)));
	assign g638 = (((!g622) & (!g627) & (!g632) & (g637) & (g42) & (g43)) + ((!g622) & (!g627) & (g632) & (!g637) & (!g42) & (g43)) + ((!g622) & (!g627) & (g632) & (g637) & (!g42) & (g43)) + ((!g622) & (!g627) & (g632) & (g637) & (g42) & (g43)) + ((!g622) & (g627) & (!g632) & (!g637) & (g42) & (!g43)) + ((!g622) & (g627) & (!g632) & (g637) & (g42) & (!g43)) + ((!g622) & (g627) & (!g632) & (g637) & (g42) & (g43)) + ((!g622) & (g627) & (g632) & (!g637) & (!g42) & (g43)) + ((!g622) & (g627) & (g632) & (!g637) & (g42) & (!g43)) + ((!g622) & (g627) & (g632) & (g637) & (!g42) & (g43)) + ((!g622) & (g627) & (g632) & (g637) & (g42) & (!g43)) + ((!g622) & (g627) & (g632) & (g637) & (g42) & (g43)) + ((g622) & (!g627) & (!g632) & (!g637) & (!g42) & (!g43)) + ((g622) & (!g627) & (!g632) & (g637) & (!g42) & (!g43)) + ((g622) & (!g627) & (!g632) & (g637) & (g42) & (g43)) + ((g622) & (!g627) & (g632) & (!g637) & (!g42) & (!g43)) + ((g622) & (!g627) & (g632) & (!g637) & (!g42) & (g43)) + ((g622) & (!g627) & (g632) & (g637) & (!g42) & (!g43)) + ((g622) & (!g627) & (g632) & (g637) & (!g42) & (g43)) + ((g622) & (!g627) & (g632) & (g637) & (g42) & (g43)) + ((g622) & (g627) & (!g632) & (!g637) & (!g42) & (!g43)) + ((g622) & (g627) & (!g632) & (!g637) & (g42) & (!g43)) + ((g622) & (g627) & (!g632) & (g637) & (!g42) & (!g43)) + ((g622) & (g627) & (!g632) & (g637) & (g42) & (!g43)) + ((g622) & (g627) & (!g632) & (g637) & (g42) & (g43)) + ((g622) & (g627) & (g632) & (!g637) & (!g42) & (!g43)) + ((g622) & (g627) & (g632) & (!g637) & (!g42) & (g43)) + ((g622) & (g627) & (g632) & (!g637) & (g42) & (!g43)) + ((g622) & (g627) & (g632) & (g637) & (!g42) & (!g43)) + ((g622) & (g627) & (g632) & (g637) & (!g42) & (g43)) + ((g622) & (g627) & (g632) & (g637) & (g42) & (!g43)) + ((g622) & (g627) & (g632) & (g637) & (g42) & (g43)));
	assign g7259 = (((!g832) & (g1679) & (!g639)) + ((!g832) & (g1679) & (g639)) + ((g832) & (!g1679) & (g639)) + ((g832) & (g1679) & (g639)));
	assign g640 = (((!g34) & (!reset) & (!g638) & (g639)) + ((!g34) & (!reset) & (g638) & (g639)) + ((g34) & (!reset) & (g638) & (!g639)) + ((g34) & (!reset) & (g638) & (g639)));
	assign g645 = (((!g641) & (!g642) & (!g643) & (g644) & (g42) & (g43)) + ((!g641) & (!g642) & (g643) & (!g644) & (!g42) & (g43)) + ((!g641) & (!g642) & (g643) & (g644) & (!g42) & (g43)) + ((!g641) & (!g642) & (g643) & (g644) & (g42) & (g43)) + ((!g641) & (g642) & (!g643) & (!g644) & (g42) & (!g43)) + ((!g641) & (g642) & (!g643) & (g644) & (g42) & (!g43)) + ((!g641) & (g642) & (!g643) & (g644) & (g42) & (g43)) + ((!g641) & (g642) & (g643) & (!g644) & (!g42) & (g43)) + ((!g641) & (g642) & (g643) & (!g644) & (g42) & (!g43)) + ((!g641) & (g642) & (g643) & (g644) & (!g42) & (g43)) + ((!g641) & (g642) & (g643) & (g644) & (g42) & (!g43)) + ((!g641) & (g642) & (g643) & (g644) & (g42) & (g43)) + ((g641) & (!g642) & (!g643) & (!g644) & (!g42) & (!g43)) + ((g641) & (!g642) & (!g643) & (g644) & (!g42) & (!g43)) + ((g641) & (!g642) & (!g643) & (g644) & (g42) & (g43)) + ((g641) & (!g642) & (g643) & (!g644) & (!g42) & (!g43)) + ((g641) & (!g642) & (g643) & (!g644) & (!g42) & (g43)) + ((g641) & (!g642) & (g643) & (g644) & (!g42) & (!g43)) + ((g641) & (!g642) & (g643) & (g644) & (!g42) & (g43)) + ((g641) & (!g642) & (g643) & (g644) & (g42) & (g43)) + ((g641) & (g642) & (!g643) & (!g644) & (!g42) & (!g43)) + ((g641) & (g642) & (!g643) & (!g644) & (g42) & (!g43)) + ((g641) & (g642) & (!g643) & (g644) & (!g42) & (!g43)) + ((g641) & (g642) & (!g643) & (g644) & (g42) & (!g43)) + ((g641) & (g642) & (!g643) & (g644) & (g42) & (g43)) + ((g641) & (g642) & (g643) & (!g644) & (!g42) & (!g43)) + ((g641) & (g642) & (g643) & (!g644) & (!g42) & (g43)) + ((g641) & (g642) & (g643) & (!g644) & (g42) & (!g43)) + ((g641) & (g642) & (g643) & (g644) & (!g42) & (!g43)) + ((g641) & (g642) & (g643) & (g644) & (!g42) & (g43)) + ((g641) & (g642) & (g643) & (g644) & (g42) & (!g43)) + ((g641) & (g642) & (g643) & (g644) & (g42) & (g43)));
	assign g650 = (((!g646) & (!g647) & (!g648) & (g649) & (g42) & (g43)) + ((!g646) & (!g647) & (g648) & (!g649) & (!g42) & (g43)) + ((!g646) & (!g647) & (g648) & (g649) & (!g42) & (g43)) + ((!g646) & (!g647) & (g648) & (g649) & (g42) & (g43)) + ((!g646) & (g647) & (!g648) & (!g649) & (g42) & (!g43)) + ((!g646) & (g647) & (!g648) & (g649) & (g42) & (!g43)) + ((!g646) & (g647) & (!g648) & (g649) & (g42) & (g43)) + ((!g646) & (g647) & (g648) & (!g649) & (!g42) & (g43)) + ((!g646) & (g647) & (g648) & (!g649) & (g42) & (!g43)) + ((!g646) & (g647) & (g648) & (g649) & (!g42) & (g43)) + ((!g646) & (g647) & (g648) & (g649) & (g42) & (!g43)) + ((!g646) & (g647) & (g648) & (g649) & (g42) & (g43)) + ((g646) & (!g647) & (!g648) & (!g649) & (!g42) & (!g43)) + ((g646) & (!g647) & (!g648) & (g649) & (!g42) & (!g43)) + ((g646) & (!g647) & (!g648) & (g649) & (g42) & (g43)) + ((g646) & (!g647) & (g648) & (!g649) & (!g42) & (!g43)) + ((g646) & (!g647) & (g648) & (!g649) & (!g42) & (g43)) + ((g646) & (!g647) & (g648) & (g649) & (!g42) & (!g43)) + ((g646) & (!g647) & (g648) & (g649) & (!g42) & (g43)) + ((g646) & (!g647) & (g648) & (g649) & (g42) & (g43)) + ((g646) & (g647) & (!g648) & (!g649) & (!g42) & (!g43)) + ((g646) & (g647) & (!g648) & (!g649) & (g42) & (!g43)) + ((g646) & (g647) & (!g648) & (g649) & (!g42) & (!g43)) + ((g646) & (g647) & (!g648) & (g649) & (g42) & (!g43)) + ((g646) & (g647) & (!g648) & (g649) & (g42) & (g43)) + ((g646) & (g647) & (g648) & (!g649) & (!g42) & (!g43)) + ((g646) & (g647) & (g648) & (!g649) & (!g42) & (g43)) + ((g646) & (g647) & (g648) & (!g649) & (g42) & (!g43)) + ((g646) & (g647) & (g648) & (g649) & (!g42) & (!g43)) + ((g646) & (g647) & (g648) & (g649) & (!g42) & (g43)) + ((g646) & (g647) & (g648) & (g649) & (g42) & (!g43)) + ((g646) & (g647) & (g648) & (g649) & (g42) & (g43)));
	assign g655 = (((!g651) & (!g652) & (!g653) & (g654) & (g42) & (g43)) + ((!g651) & (!g652) & (g653) & (!g654) & (!g42) & (g43)) + ((!g651) & (!g652) & (g653) & (g654) & (!g42) & (g43)) + ((!g651) & (!g652) & (g653) & (g654) & (g42) & (g43)) + ((!g651) & (g652) & (!g653) & (!g654) & (g42) & (!g43)) + ((!g651) & (g652) & (!g653) & (g654) & (g42) & (!g43)) + ((!g651) & (g652) & (!g653) & (g654) & (g42) & (g43)) + ((!g651) & (g652) & (g653) & (!g654) & (!g42) & (g43)) + ((!g651) & (g652) & (g653) & (!g654) & (g42) & (!g43)) + ((!g651) & (g652) & (g653) & (g654) & (!g42) & (g43)) + ((!g651) & (g652) & (g653) & (g654) & (g42) & (!g43)) + ((!g651) & (g652) & (g653) & (g654) & (g42) & (g43)) + ((g651) & (!g652) & (!g653) & (!g654) & (!g42) & (!g43)) + ((g651) & (!g652) & (!g653) & (g654) & (!g42) & (!g43)) + ((g651) & (!g652) & (!g653) & (g654) & (g42) & (g43)) + ((g651) & (!g652) & (g653) & (!g654) & (!g42) & (!g43)) + ((g651) & (!g652) & (g653) & (!g654) & (!g42) & (g43)) + ((g651) & (!g652) & (g653) & (g654) & (!g42) & (!g43)) + ((g651) & (!g652) & (g653) & (g654) & (!g42) & (g43)) + ((g651) & (!g652) & (g653) & (g654) & (g42) & (g43)) + ((g651) & (g652) & (!g653) & (!g654) & (!g42) & (!g43)) + ((g651) & (g652) & (!g653) & (!g654) & (g42) & (!g43)) + ((g651) & (g652) & (!g653) & (g654) & (!g42) & (!g43)) + ((g651) & (g652) & (!g653) & (g654) & (g42) & (!g43)) + ((g651) & (g652) & (!g653) & (g654) & (g42) & (g43)) + ((g651) & (g652) & (g653) & (!g654) & (!g42) & (!g43)) + ((g651) & (g652) & (g653) & (!g654) & (!g42) & (g43)) + ((g651) & (g652) & (g653) & (!g654) & (g42) & (!g43)) + ((g651) & (g652) & (g653) & (g654) & (!g42) & (!g43)) + ((g651) & (g652) & (g653) & (g654) & (!g42) & (g43)) + ((g651) & (g652) & (g653) & (g654) & (g42) & (!g43)) + ((g651) & (g652) & (g653) & (g654) & (g42) & (g43)));
	assign g660 = (((!g656) & (!g657) & (!g658) & (g659) & (g42) & (g43)) + ((!g656) & (!g657) & (g658) & (!g659) & (!g42) & (g43)) + ((!g656) & (!g657) & (g658) & (g659) & (!g42) & (g43)) + ((!g656) & (!g657) & (g658) & (g659) & (g42) & (g43)) + ((!g656) & (g657) & (!g658) & (!g659) & (g42) & (!g43)) + ((!g656) & (g657) & (!g658) & (g659) & (g42) & (!g43)) + ((!g656) & (g657) & (!g658) & (g659) & (g42) & (g43)) + ((!g656) & (g657) & (g658) & (!g659) & (!g42) & (g43)) + ((!g656) & (g657) & (g658) & (!g659) & (g42) & (!g43)) + ((!g656) & (g657) & (g658) & (g659) & (!g42) & (g43)) + ((!g656) & (g657) & (g658) & (g659) & (g42) & (!g43)) + ((!g656) & (g657) & (g658) & (g659) & (g42) & (g43)) + ((g656) & (!g657) & (!g658) & (!g659) & (!g42) & (!g43)) + ((g656) & (!g657) & (!g658) & (g659) & (!g42) & (!g43)) + ((g656) & (!g657) & (!g658) & (g659) & (g42) & (g43)) + ((g656) & (!g657) & (g658) & (!g659) & (!g42) & (!g43)) + ((g656) & (!g657) & (g658) & (!g659) & (!g42) & (g43)) + ((g656) & (!g657) & (g658) & (g659) & (!g42) & (!g43)) + ((g656) & (!g657) & (g658) & (g659) & (!g42) & (g43)) + ((g656) & (!g657) & (g658) & (g659) & (g42) & (g43)) + ((g656) & (g657) & (!g658) & (!g659) & (!g42) & (!g43)) + ((g656) & (g657) & (!g658) & (!g659) & (g42) & (!g43)) + ((g656) & (g657) & (!g658) & (g659) & (!g42) & (!g43)) + ((g656) & (g657) & (!g658) & (g659) & (g42) & (!g43)) + ((g656) & (g657) & (!g658) & (g659) & (g42) & (g43)) + ((g656) & (g657) & (g658) & (!g659) & (!g42) & (!g43)) + ((g656) & (g657) & (g658) & (!g659) & (!g42) & (g43)) + ((g656) & (g657) & (g658) & (!g659) & (g42) & (!g43)) + ((g656) & (g657) & (g658) & (g659) & (!g42) & (!g43)) + ((g656) & (g657) & (g658) & (g659) & (!g42) & (g43)) + ((g656) & (g657) & (g658) & (g659) & (g42) & (!g43)) + ((g656) & (g657) & (g658) & (g659) & (g42) & (g43)));
	assign g661 = (((!g645) & (!g650) & (!g655) & (g660) & (g60) & (g61)) + ((!g645) & (!g650) & (g655) & (!g660) & (!g60) & (g61)) + ((!g645) & (!g650) & (g655) & (g660) & (!g60) & (g61)) + ((!g645) & (!g650) & (g655) & (g660) & (g60) & (g61)) + ((!g645) & (g650) & (!g655) & (!g660) & (g60) & (!g61)) + ((!g645) & (g650) & (!g655) & (g660) & (g60) & (!g61)) + ((!g645) & (g650) & (!g655) & (g660) & (g60) & (g61)) + ((!g645) & (g650) & (g655) & (!g660) & (!g60) & (g61)) + ((!g645) & (g650) & (g655) & (!g660) & (g60) & (!g61)) + ((!g645) & (g650) & (g655) & (g660) & (!g60) & (g61)) + ((!g645) & (g650) & (g655) & (g660) & (g60) & (!g61)) + ((!g645) & (g650) & (g655) & (g660) & (g60) & (g61)) + ((g645) & (!g650) & (!g655) & (!g660) & (!g60) & (!g61)) + ((g645) & (!g650) & (!g655) & (g660) & (!g60) & (!g61)) + ((g645) & (!g650) & (!g655) & (g660) & (g60) & (g61)) + ((g645) & (!g650) & (g655) & (!g660) & (!g60) & (!g61)) + ((g645) & (!g650) & (g655) & (!g660) & (!g60) & (g61)) + ((g645) & (!g650) & (g655) & (g660) & (!g60) & (!g61)) + ((g645) & (!g650) & (g655) & (g660) & (!g60) & (g61)) + ((g645) & (!g650) & (g655) & (g660) & (g60) & (g61)) + ((g645) & (g650) & (!g655) & (!g660) & (!g60) & (!g61)) + ((g645) & (g650) & (!g655) & (!g660) & (g60) & (!g61)) + ((g645) & (g650) & (!g655) & (g660) & (!g60) & (!g61)) + ((g645) & (g650) & (!g655) & (g660) & (g60) & (!g61)) + ((g645) & (g650) & (!g655) & (g660) & (g60) & (g61)) + ((g645) & (g650) & (g655) & (!g660) & (!g60) & (!g61)) + ((g645) & (g650) & (g655) & (!g660) & (!g60) & (g61)) + ((g645) & (g650) & (g655) & (!g660) & (g60) & (!g61)) + ((g645) & (g650) & (g655) & (g660) & (!g60) & (!g61)) + ((g645) & (g650) & (g655) & (g660) & (!g60) & (g61)) + ((g645) & (g650) & (g655) & (g660) & (g60) & (!g61)) + ((g645) & (g650) & (g655) & (g660) & (g60) & (g61)));
	assign g7260 = (((!g832) & (g1712) & (!g662)) + ((!g832) & (g1712) & (g662)) + ((g832) & (!g1712) & (g662)) + ((g832) & (g1712) & (g662)));
	assign g663 = (((!g34) & (!reset) & (!g661) & (g662)) + ((!g34) & (!reset) & (g661) & (g662)) + ((g34) & (!reset) & (g661) & (!g662)) + ((g34) & (!reset) & (g661) & (g662)));
	assign g668 = (((!g664) & (!g665) & (!g666) & (g667) & (g60) & (g61)) + ((!g664) & (!g665) & (g666) & (!g667) & (!g60) & (g61)) + ((!g664) & (!g665) & (g666) & (g667) & (!g60) & (g61)) + ((!g664) & (!g665) & (g666) & (g667) & (g60) & (g61)) + ((!g664) & (g665) & (!g666) & (!g667) & (g60) & (!g61)) + ((!g664) & (g665) & (!g666) & (g667) & (g60) & (!g61)) + ((!g664) & (g665) & (!g666) & (g667) & (g60) & (g61)) + ((!g664) & (g665) & (g666) & (!g667) & (!g60) & (g61)) + ((!g664) & (g665) & (g666) & (!g667) & (g60) & (!g61)) + ((!g664) & (g665) & (g666) & (g667) & (!g60) & (g61)) + ((!g664) & (g665) & (g666) & (g667) & (g60) & (!g61)) + ((!g664) & (g665) & (g666) & (g667) & (g60) & (g61)) + ((g664) & (!g665) & (!g666) & (!g667) & (!g60) & (!g61)) + ((g664) & (!g665) & (!g666) & (g667) & (!g60) & (!g61)) + ((g664) & (!g665) & (!g666) & (g667) & (g60) & (g61)) + ((g664) & (!g665) & (g666) & (!g667) & (!g60) & (!g61)) + ((g664) & (!g665) & (g666) & (!g667) & (!g60) & (g61)) + ((g664) & (!g665) & (g666) & (g667) & (!g60) & (!g61)) + ((g664) & (!g665) & (g666) & (g667) & (!g60) & (g61)) + ((g664) & (!g665) & (g666) & (g667) & (g60) & (g61)) + ((g664) & (g665) & (!g666) & (!g667) & (!g60) & (!g61)) + ((g664) & (g665) & (!g666) & (!g667) & (g60) & (!g61)) + ((g664) & (g665) & (!g666) & (g667) & (!g60) & (!g61)) + ((g664) & (g665) & (!g666) & (g667) & (g60) & (!g61)) + ((g664) & (g665) & (!g666) & (g667) & (g60) & (g61)) + ((g664) & (g665) & (g666) & (!g667) & (!g60) & (!g61)) + ((g664) & (g665) & (g666) & (!g667) & (!g60) & (g61)) + ((g664) & (g665) & (g666) & (!g667) & (g60) & (!g61)) + ((g664) & (g665) & (g666) & (g667) & (!g60) & (!g61)) + ((g664) & (g665) & (g666) & (g667) & (!g60) & (g61)) + ((g664) & (g665) & (g666) & (g667) & (g60) & (!g61)) + ((g664) & (g665) & (g666) & (g667) & (g60) & (g61)));
	assign g673 = (((!g669) & (!g670) & (!g671) & (g672) & (g60) & (g61)) + ((!g669) & (!g670) & (g671) & (!g672) & (!g60) & (g61)) + ((!g669) & (!g670) & (g671) & (g672) & (!g60) & (g61)) + ((!g669) & (!g670) & (g671) & (g672) & (g60) & (g61)) + ((!g669) & (g670) & (!g671) & (!g672) & (g60) & (!g61)) + ((!g669) & (g670) & (!g671) & (g672) & (g60) & (!g61)) + ((!g669) & (g670) & (!g671) & (g672) & (g60) & (g61)) + ((!g669) & (g670) & (g671) & (!g672) & (!g60) & (g61)) + ((!g669) & (g670) & (g671) & (!g672) & (g60) & (!g61)) + ((!g669) & (g670) & (g671) & (g672) & (!g60) & (g61)) + ((!g669) & (g670) & (g671) & (g672) & (g60) & (!g61)) + ((!g669) & (g670) & (g671) & (g672) & (g60) & (g61)) + ((g669) & (!g670) & (!g671) & (!g672) & (!g60) & (!g61)) + ((g669) & (!g670) & (!g671) & (g672) & (!g60) & (!g61)) + ((g669) & (!g670) & (!g671) & (g672) & (g60) & (g61)) + ((g669) & (!g670) & (g671) & (!g672) & (!g60) & (!g61)) + ((g669) & (!g670) & (g671) & (!g672) & (!g60) & (g61)) + ((g669) & (!g670) & (g671) & (g672) & (!g60) & (!g61)) + ((g669) & (!g670) & (g671) & (g672) & (!g60) & (g61)) + ((g669) & (!g670) & (g671) & (g672) & (g60) & (g61)) + ((g669) & (g670) & (!g671) & (!g672) & (!g60) & (!g61)) + ((g669) & (g670) & (!g671) & (!g672) & (g60) & (!g61)) + ((g669) & (g670) & (!g671) & (g672) & (!g60) & (!g61)) + ((g669) & (g670) & (!g671) & (g672) & (g60) & (!g61)) + ((g669) & (g670) & (!g671) & (g672) & (g60) & (g61)) + ((g669) & (g670) & (g671) & (!g672) & (!g60) & (!g61)) + ((g669) & (g670) & (g671) & (!g672) & (!g60) & (g61)) + ((g669) & (g670) & (g671) & (!g672) & (g60) & (!g61)) + ((g669) & (g670) & (g671) & (g672) & (!g60) & (!g61)) + ((g669) & (g670) & (g671) & (g672) & (!g60) & (g61)) + ((g669) & (g670) & (g671) & (g672) & (g60) & (!g61)) + ((g669) & (g670) & (g671) & (g672) & (g60) & (g61)));
	assign g678 = (((!g674) & (!g675) & (!g676) & (g677) & (g60) & (g61)) + ((!g674) & (!g675) & (g676) & (!g677) & (!g60) & (g61)) + ((!g674) & (!g675) & (g676) & (g677) & (!g60) & (g61)) + ((!g674) & (!g675) & (g676) & (g677) & (g60) & (g61)) + ((!g674) & (g675) & (!g676) & (!g677) & (g60) & (!g61)) + ((!g674) & (g675) & (!g676) & (g677) & (g60) & (!g61)) + ((!g674) & (g675) & (!g676) & (g677) & (g60) & (g61)) + ((!g674) & (g675) & (g676) & (!g677) & (!g60) & (g61)) + ((!g674) & (g675) & (g676) & (!g677) & (g60) & (!g61)) + ((!g674) & (g675) & (g676) & (g677) & (!g60) & (g61)) + ((!g674) & (g675) & (g676) & (g677) & (g60) & (!g61)) + ((!g674) & (g675) & (g676) & (g677) & (g60) & (g61)) + ((g674) & (!g675) & (!g676) & (!g677) & (!g60) & (!g61)) + ((g674) & (!g675) & (!g676) & (g677) & (!g60) & (!g61)) + ((g674) & (!g675) & (!g676) & (g677) & (g60) & (g61)) + ((g674) & (!g675) & (g676) & (!g677) & (!g60) & (!g61)) + ((g674) & (!g675) & (g676) & (!g677) & (!g60) & (g61)) + ((g674) & (!g675) & (g676) & (g677) & (!g60) & (!g61)) + ((g674) & (!g675) & (g676) & (g677) & (!g60) & (g61)) + ((g674) & (!g675) & (g676) & (g677) & (g60) & (g61)) + ((g674) & (g675) & (!g676) & (!g677) & (!g60) & (!g61)) + ((g674) & (g675) & (!g676) & (!g677) & (g60) & (!g61)) + ((g674) & (g675) & (!g676) & (g677) & (!g60) & (!g61)) + ((g674) & (g675) & (!g676) & (g677) & (g60) & (!g61)) + ((g674) & (g675) & (!g676) & (g677) & (g60) & (g61)) + ((g674) & (g675) & (g676) & (!g677) & (!g60) & (!g61)) + ((g674) & (g675) & (g676) & (!g677) & (!g60) & (g61)) + ((g674) & (g675) & (g676) & (!g677) & (g60) & (!g61)) + ((g674) & (g675) & (g676) & (g677) & (!g60) & (!g61)) + ((g674) & (g675) & (g676) & (g677) & (!g60) & (g61)) + ((g674) & (g675) & (g676) & (g677) & (g60) & (!g61)) + ((g674) & (g675) & (g676) & (g677) & (g60) & (g61)));
	assign g683 = (((!g679) & (!g680) & (!g681) & (g682) & (g60) & (g61)) + ((!g679) & (!g680) & (g681) & (!g682) & (!g60) & (g61)) + ((!g679) & (!g680) & (g681) & (g682) & (!g60) & (g61)) + ((!g679) & (!g680) & (g681) & (g682) & (g60) & (g61)) + ((!g679) & (g680) & (!g681) & (!g682) & (g60) & (!g61)) + ((!g679) & (g680) & (!g681) & (g682) & (g60) & (!g61)) + ((!g679) & (g680) & (!g681) & (g682) & (g60) & (g61)) + ((!g679) & (g680) & (g681) & (!g682) & (!g60) & (g61)) + ((!g679) & (g680) & (g681) & (!g682) & (g60) & (!g61)) + ((!g679) & (g680) & (g681) & (g682) & (!g60) & (g61)) + ((!g679) & (g680) & (g681) & (g682) & (g60) & (!g61)) + ((!g679) & (g680) & (g681) & (g682) & (g60) & (g61)) + ((g679) & (!g680) & (!g681) & (!g682) & (!g60) & (!g61)) + ((g679) & (!g680) & (!g681) & (g682) & (!g60) & (!g61)) + ((g679) & (!g680) & (!g681) & (g682) & (g60) & (g61)) + ((g679) & (!g680) & (g681) & (!g682) & (!g60) & (!g61)) + ((g679) & (!g680) & (g681) & (!g682) & (!g60) & (g61)) + ((g679) & (!g680) & (g681) & (g682) & (!g60) & (!g61)) + ((g679) & (!g680) & (g681) & (g682) & (!g60) & (g61)) + ((g679) & (!g680) & (g681) & (g682) & (g60) & (g61)) + ((g679) & (g680) & (!g681) & (!g682) & (!g60) & (!g61)) + ((g679) & (g680) & (!g681) & (!g682) & (g60) & (!g61)) + ((g679) & (g680) & (!g681) & (g682) & (!g60) & (!g61)) + ((g679) & (g680) & (!g681) & (g682) & (g60) & (!g61)) + ((g679) & (g680) & (!g681) & (g682) & (g60) & (g61)) + ((g679) & (g680) & (g681) & (!g682) & (!g60) & (!g61)) + ((g679) & (g680) & (g681) & (!g682) & (!g60) & (g61)) + ((g679) & (g680) & (g681) & (!g682) & (g60) & (!g61)) + ((g679) & (g680) & (g681) & (g682) & (!g60) & (!g61)) + ((g679) & (g680) & (g681) & (g682) & (!g60) & (g61)) + ((g679) & (g680) & (g681) & (g682) & (g60) & (!g61)) + ((g679) & (g680) & (g681) & (g682) & (g60) & (g61)));
	assign g684 = (((!g668) & (!g673) & (!g678) & (g683) & (g42) & (g43)) + ((!g668) & (!g673) & (g678) & (!g683) & (!g42) & (g43)) + ((!g668) & (!g673) & (g678) & (g683) & (!g42) & (g43)) + ((!g668) & (!g673) & (g678) & (g683) & (g42) & (g43)) + ((!g668) & (g673) & (!g678) & (!g683) & (g42) & (!g43)) + ((!g668) & (g673) & (!g678) & (g683) & (g42) & (!g43)) + ((!g668) & (g673) & (!g678) & (g683) & (g42) & (g43)) + ((!g668) & (g673) & (g678) & (!g683) & (!g42) & (g43)) + ((!g668) & (g673) & (g678) & (!g683) & (g42) & (!g43)) + ((!g668) & (g673) & (g678) & (g683) & (!g42) & (g43)) + ((!g668) & (g673) & (g678) & (g683) & (g42) & (!g43)) + ((!g668) & (g673) & (g678) & (g683) & (g42) & (g43)) + ((g668) & (!g673) & (!g678) & (!g683) & (!g42) & (!g43)) + ((g668) & (!g673) & (!g678) & (g683) & (!g42) & (!g43)) + ((g668) & (!g673) & (!g678) & (g683) & (g42) & (g43)) + ((g668) & (!g673) & (g678) & (!g683) & (!g42) & (!g43)) + ((g668) & (!g673) & (g678) & (!g683) & (!g42) & (g43)) + ((g668) & (!g673) & (g678) & (g683) & (!g42) & (!g43)) + ((g668) & (!g673) & (g678) & (g683) & (!g42) & (g43)) + ((g668) & (!g673) & (g678) & (g683) & (g42) & (g43)) + ((g668) & (g673) & (!g678) & (!g683) & (!g42) & (!g43)) + ((g668) & (g673) & (!g678) & (!g683) & (g42) & (!g43)) + ((g668) & (g673) & (!g678) & (g683) & (!g42) & (!g43)) + ((g668) & (g673) & (!g678) & (g683) & (g42) & (!g43)) + ((g668) & (g673) & (!g678) & (g683) & (g42) & (g43)) + ((g668) & (g673) & (g678) & (!g683) & (!g42) & (!g43)) + ((g668) & (g673) & (g678) & (!g683) & (!g42) & (g43)) + ((g668) & (g673) & (g678) & (!g683) & (g42) & (!g43)) + ((g668) & (g673) & (g678) & (g683) & (!g42) & (!g43)) + ((g668) & (g673) & (g678) & (g683) & (!g42) & (g43)) + ((g668) & (g673) & (g678) & (g683) & (g42) & (!g43)) + ((g668) & (g673) & (g678) & (g683) & (g42) & (g43)));
	assign g7261 = (((!g832) & (g1746) & (!g685)) + ((!g832) & (g1746) & (g685)) + ((g832) & (!g1746) & (g685)) + ((g832) & (g1746) & (g685)));
	assign g686 = (((!g34) & (!reset) & (!g684) & (g685)) + ((!g34) & (!reset) & (g684) & (g685)) + ((g34) & (!reset) & (g684) & (!g685)) + ((g34) & (!reset) & (g684) & (g685)));
	assign g691 = (((!g687) & (!g688) & (!g689) & (g690) & (g42) & (g43)) + ((!g687) & (!g688) & (g689) & (!g690) & (!g42) & (g43)) + ((!g687) & (!g688) & (g689) & (g690) & (!g42) & (g43)) + ((!g687) & (!g688) & (g689) & (g690) & (g42) & (g43)) + ((!g687) & (g688) & (!g689) & (!g690) & (g42) & (!g43)) + ((!g687) & (g688) & (!g689) & (g690) & (g42) & (!g43)) + ((!g687) & (g688) & (!g689) & (g690) & (g42) & (g43)) + ((!g687) & (g688) & (g689) & (!g690) & (!g42) & (g43)) + ((!g687) & (g688) & (g689) & (!g690) & (g42) & (!g43)) + ((!g687) & (g688) & (g689) & (g690) & (!g42) & (g43)) + ((!g687) & (g688) & (g689) & (g690) & (g42) & (!g43)) + ((!g687) & (g688) & (g689) & (g690) & (g42) & (g43)) + ((g687) & (!g688) & (!g689) & (!g690) & (!g42) & (!g43)) + ((g687) & (!g688) & (!g689) & (g690) & (!g42) & (!g43)) + ((g687) & (!g688) & (!g689) & (g690) & (g42) & (g43)) + ((g687) & (!g688) & (g689) & (!g690) & (!g42) & (!g43)) + ((g687) & (!g688) & (g689) & (!g690) & (!g42) & (g43)) + ((g687) & (!g688) & (g689) & (g690) & (!g42) & (!g43)) + ((g687) & (!g688) & (g689) & (g690) & (!g42) & (g43)) + ((g687) & (!g688) & (g689) & (g690) & (g42) & (g43)) + ((g687) & (g688) & (!g689) & (!g690) & (!g42) & (!g43)) + ((g687) & (g688) & (!g689) & (!g690) & (g42) & (!g43)) + ((g687) & (g688) & (!g689) & (g690) & (!g42) & (!g43)) + ((g687) & (g688) & (!g689) & (g690) & (g42) & (!g43)) + ((g687) & (g688) & (!g689) & (g690) & (g42) & (g43)) + ((g687) & (g688) & (g689) & (!g690) & (!g42) & (!g43)) + ((g687) & (g688) & (g689) & (!g690) & (!g42) & (g43)) + ((g687) & (g688) & (g689) & (!g690) & (g42) & (!g43)) + ((g687) & (g688) & (g689) & (g690) & (!g42) & (!g43)) + ((g687) & (g688) & (g689) & (g690) & (!g42) & (g43)) + ((g687) & (g688) & (g689) & (g690) & (g42) & (!g43)) + ((g687) & (g688) & (g689) & (g690) & (g42) & (g43)));
	assign g696 = (((!g692) & (!g693) & (!g694) & (g695) & (g42) & (g43)) + ((!g692) & (!g693) & (g694) & (!g695) & (!g42) & (g43)) + ((!g692) & (!g693) & (g694) & (g695) & (!g42) & (g43)) + ((!g692) & (!g693) & (g694) & (g695) & (g42) & (g43)) + ((!g692) & (g693) & (!g694) & (!g695) & (g42) & (!g43)) + ((!g692) & (g693) & (!g694) & (g695) & (g42) & (!g43)) + ((!g692) & (g693) & (!g694) & (g695) & (g42) & (g43)) + ((!g692) & (g693) & (g694) & (!g695) & (!g42) & (g43)) + ((!g692) & (g693) & (g694) & (!g695) & (g42) & (!g43)) + ((!g692) & (g693) & (g694) & (g695) & (!g42) & (g43)) + ((!g692) & (g693) & (g694) & (g695) & (g42) & (!g43)) + ((!g692) & (g693) & (g694) & (g695) & (g42) & (g43)) + ((g692) & (!g693) & (!g694) & (!g695) & (!g42) & (!g43)) + ((g692) & (!g693) & (!g694) & (g695) & (!g42) & (!g43)) + ((g692) & (!g693) & (!g694) & (g695) & (g42) & (g43)) + ((g692) & (!g693) & (g694) & (!g695) & (!g42) & (!g43)) + ((g692) & (!g693) & (g694) & (!g695) & (!g42) & (g43)) + ((g692) & (!g693) & (g694) & (g695) & (!g42) & (!g43)) + ((g692) & (!g693) & (g694) & (g695) & (!g42) & (g43)) + ((g692) & (!g693) & (g694) & (g695) & (g42) & (g43)) + ((g692) & (g693) & (!g694) & (!g695) & (!g42) & (!g43)) + ((g692) & (g693) & (!g694) & (!g695) & (g42) & (!g43)) + ((g692) & (g693) & (!g694) & (g695) & (!g42) & (!g43)) + ((g692) & (g693) & (!g694) & (g695) & (g42) & (!g43)) + ((g692) & (g693) & (!g694) & (g695) & (g42) & (g43)) + ((g692) & (g693) & (g694) & (!g695) & (!g42) & (!g43)) + ((g692) & (g693) & (g694) & (!g695) & (!g42) & (g43)) + ((g692) & (g693) & (g694) & (!g695) & (g42) & (!g43)) + ((g692) & (g693) & (g694) & (g695) & (!g42) & (!g43)) + ((g692) & (g693) & (g694) & (g695) & (!g42) & (g43)) + ((g692) & (g693) & (g694) & (g695) & (g42) & (!g43)) + ((g692) & (g693) & (g694) & (g695) & (g42) & (g43)));
	assign g701 = (((!g697) & (!g698) & (!g699) & (g700) & (g42) & (g43)) + ((!g697) & (!g698) & (g699) & (!g700) & (!g42) & (g43)) + ((!g697) & (!g698) & (g699) & (g700) & (!g42) & (g43)) + ((!g697) & (!g698) & (g699) & (g700) & (g42) & (g43)) + ((!g697) & (g698) & (!g699) & (!g700) & (g42) & (!g43)) + ((!g697) & (g698) & (!g699) & (g700) & (g42) & (!g43)) + ((!g697) & (g698) & (!g699) & (g700) & (g42) & (g43)) + ((!g697) & (g698) & (g699) & (!g700) & (!g42) & (g43)) + ((!g697) & (g698) & (g699) & (!g700) & (g42) & (!g43)) + ((!g697) & (g698) & (g699) & (g700) & (!g42) & (g43)) + ((!g697) & (g698) & (g699) & (g700) & (g42) & (!g43)) + ((!g697) & (g698) & (g699) & (g700) & (g42) & (g43)) + ((g697) & (!g698) & (!g699) & (!g700) & (!g42) & (!g43)) + ((g697) & (!g698) & (!g699) & (g700) & (!g42) & (!g43)) + ((g697) & (!g698) & (!g699) & (g700) & (g42) & (g43)) + ((g697) & (!g698) & (g699) & (!g700) & (!g42) & (!g43)) + ((g697) & (!g698) & (g699) & (!g700) & (!g42) & (g43)) + ((g697) & (!g698) & (g699) & (g700) & (!g42) & (!g43)) + ((g697) & (!g698) & (g699) & (g700) & (!g42) & (g43)) + ((g697) & (!g698) & (g699) & (g700) & (g42) & (g43)) + ((g697) & (g698) & (!g699) & (!g700) & (!g42) & (!g43)) + ((g697) & (g698) & (!g699) & (!g700) & (g42) & (!g43)) + ((g697) & (g698) & (!g699) & (g700) & (!g42) & (!g43)) + ((g697) & (g698) & (!g699) & (g700) & (g42) & (!g43)) + ((g697) & (g698) & (!g699) & (g700) & (g42) & (g43)) + ((g697) & (g698) & (g699) & (!g700) & (!g42) & (!g43)) + ((g697) & (g698) & (g699) & (!g700) & (!g42) & (g43)) + ((g697) & (g698) & (g699) & (!g700) & (g42) & (!g43)) + ((g697) & (g698) & (g699) & (g700) & (!g42) & (!g43)) + ((g697) & (g698) & (g699) & (g700) & (!g42) & (g43)) + ((g697) & (g698) & (g699) & (g700) & (g42) & (!g43)) + ((g697) & (g698) & (g699) & (g700) & (g42) & (g43)));
	assign g706 = (((!g702) & (!g703) & (!g704) & (g705) & (g42) & (g43)) + ((!g702) & (!g703) & (g704) & (!g705) & (!g42) & (g43)) + ((!g702) & (!g703) & (g704) & (g705) & (!g42) & (g43)) + ((!g702) & (!g703) & (g704) & (g705) & (g42) & (g43)) + ((!g702) & (g703) & (!g704) & (!g705) & (g42) & (!g43)) + ((!g702) & (g703) & (!g704) & (g705) & (g42) & (!g43)) + ((!g702) & (g703) & (!g704) & (g705) & (g42) & (g43)) + ((!g702) & (g703) & (g704) & (!g705) & (!g42) & (g43)) + ((!g702) & (g703) & (g704) & (!g705) & (g42) & (!g43)) + ((!g702) & (g703) & (g704) & (g705) & (!g42) & (g43)) + ((!g702) & (g703) & (g704) & (g705) & (g42) & (!g43)) + ((!g702) & (g703) & (g704) & (g705) & (g42) & (g43)) + ((g702) & (!g703) & (!g704) & (!g705) & (!g42) & (!g43)) + ((g702) & (!g703) & (!g704) & (g705) & (!g42) & (!g43)) + ((g702) & (!g703) & (!g704) & (g705) & (g42) & (g43)) + ((g702) & (!g703) & (g704) & (!g705) & (!g42) & (!g43)) + ((g702) & (!g703) & (g704) & (!g705) & (!g42) & (g43)) + ((g702) & (!g703) & (g704) & (g705) & (!g42) & (!g43)) + ((g702) & (!g703) & (g704) & (g705) & (!g42) & (g43)) + ((g702) & (!g703) & (g704) & (g705) & (g42) & (g43)) + ((g702) & (g703) & (!g704) & (!g705) & (!g42) & (!g43)) + ((g702) & (g703) & (!g704) & (!g705) & (g42) & (!g43)) + ((g702) & (g703) & (!g704) & (g705) & (!g42) & (!g43)) + ((g702) & (g703) & (!g704) & (g705) & (g42) & (!g43)) + ((g702) & (g703) & (!g704) & (g705) & (g42) & (g43)) + ((g702) & (g703) & (g704) & (!g705) & (!g42) & (!g43)) + ((g702) & (g703) & (g704) & (!g705) & (!g42) & (g43)) + ((g702) & (g703) & (g704) & (!g705) & (g42) & (!g43)) + ((g702) & (g703) & (g704) & (g705) & (!g42) & (!g43)) + ((g702) & (g703) & (g704) & (g705) & (!g42) & (g43)) + ((g702) & (g703) & (g704) & (g705) & (g42) & (!g43)) + ((g702) & (g703) & (g704) & (g705) & (g42) & (g43)));
	assign g707 = (((!g691) & (!g696) & (!g701) & (g706) & (g60) & (g61)) + ((!g691) & (!g696) & (g701) & (!g706) & (!g60) & (g61)) + ((!g691) & (!g696) & (g701) & (g706) & (!g60) & (g61)) + ((!g691) & (!g696) & (g701) & (g706) & (g60) & (g61)) + ((!g691) & (g696) & (!g701) & (!g706) & (g60) & (!g61)) + ((!g691) & (g696) & (!g701) & (g706) & (g60) & (!g61)) + ((!g691) & (g696) & (!g701) & (g706) & (g60) & (g61)) + ((!g691) & (g696) & (g701) & (!g706) & (!g60) & (g61)) + ((!g691) & (g696) & (g701) & (!g706) & (g60) & (!g61)) + ((!g691) & (g696) & (g701) & (g706) & (!g60) & (g61)) + ((!g691) & (g696) & (g701) & (g706) & (g60) & (!g61)) + ((!g691) & (g696) & (g701) & (g706) & (g60) & (g61)) + ((g691) & (!g696) & (!g701) & (!g706) & (!g60) & (!g61)) + ((g691) & (!g696) & (!g701) & (g706) & (!g60) & (!g61)) + ((g691) & (!g696) & (!g701) & (g706) & (g60) & (g61)) + ((g691) & (!g696) & (g701) & (!g706) & (!g60) & (!g61)) + ((g691) & (!g696) & (g701) & (!g706) & (!g60) & (g61)) + ((g691) & (!g696) & (g701) & (g706) & (!g60) & (!g61)) + ((g691) & (!g696) & (g701) & (g706) & (!g60) & (g61)) + ((g691) & (!g696) & (g701) & (g706) & (g60) & (g61)) + ((g691) & (g696) & (!g701) & (!g706) & (!g60) & (!g61)) + ((g691) & (g696) & (!g701) & (!g706) & (g60) & (!g61)) + ((g691) & (g696) & (!g701) & (g706) & (!g60) & (!g61)) + ((g691) & (g696) & (!g701) & (g706) & (g60) & (!g61)) + ((g691) & (g696) & (!g701) & (g706) & (g60) & (g61)) + ((g691) & (g696) & (g701) & (!g706) & (!g60) & (!g61)) + ((g691) & (g696) & (g701) & (!g706) & (!g60) & (g61)) + ((g691) & (g696) & (g701) & (!g706) & (g60) & (!g61)) + ((g691) & (g696) & (g701) & (g706) & (!g60) & (!g61)) + ((g691) & (g696) & (g701) & (g706) & (!g60) & (g61)) + ((g691) & (g696) & (g701) & (g706) & (g60) & (!g61)) + ((g691) & (g696) & (g701) & (g706) & (g60) & (g61)));
	assign g7262 = (((!g832) & (g1782) & (!g708)) + ((!g832) & (g1782) & (g708)) + ((g832) & (!g1782) & (g708)) + ((g832) & (g1782) & (g708)));
	assign g709 = (((!g34) & (!reset) & (!g707) & (g708)) + ((!g34) & (!reset) & (g707) & (g708)) + ((g34) & (!reset) & (g707) & (!g708)) + ((g34) & (!reset) & (g707) & (g708)));
	assign g714 = (((!g710) & (!g711) & (!g712) & (g713) & (g60) & (g61)) + ((!g710) & (!g711) & (g712) & (!g713) & (!g60) & (g61)) + ((!g710) & (!g711) & (g712) & (g713) & (!g60) & (g61)) + ((!g710) & (!g711) & (g712) & (g713) & (g60) & (g61)) + ((!g710) & (g711) & (!g712) & (!g713) & (g60) & (!g61)) + ((!g710) & (g711) & (!g712) & (g713) & (g60) & (!g61)) + ((!g710) & (g711) & (!g712) & (g713) & (g60) & (g61)) + ((!g710) & (g711) & (g712) & (!g713) & (!g60) & (g61)) + ((!g710) & (g711) & (g712) & (!g713) & (g60) & (!g61)) + ((!g710) & (g711) & (g712) & (g713) & (!g60) & (g61)) + ((!g710) & (g711) & (g712) & (g713) & (g60) & (!g61)) + ((!g710) & (g711) & (g712) & (g713) & (g60) & (g61)) + ((g710) & (!g711) & (!g712) & (!g713) & (!g60) & (!g61)) + ((g710) & (!g711) & (!g712) & (g713) & (!g60) & (!g61)) + ((g710) & (!g711) & (!g712) & (g713) & (g60) & (g61)) + ((g710) & (!g711) & (g712) & (!g713) & (!g60) & (!g61)) + ((g710) & (!g711) & (g712) & (!g713) & (!g60) & (g61)) + ((g710) & (!g711) & (g712) & (g713) & (!g60) & (!g61)) + ((g710) & (!g711) & (g712) & (g713) & (!g60) & (g61)) + ((g710) & (!g711) & (g712) & (g713) & (g60) & (g61)) + ((g710) & (g711) & (!g712) & (!g713) & (!g60) & (!g61)) + ((g710) & (g711) & (!g712) & (!g713) & (g60) & (!g61)) + ((g710) & (g711) & (!g712) & (g713) & (!g60) & (!g61)) + ((g710) & (g711) & (!g712) & (g713) & (g60) & (!g61)) + ((g710) & (g711) & (!g712) & (g713) & (g60) & (g61)) + ((g710) & (g711) & (g712) & (!g713) & (!g60) & (!g61)) + ((g710) & (g711) & (g712) & (!g713) & (!g60) & (g61)) + ((g710) & (g711) & (g712) & (!g713) & (g60) & (!g61)) + ((g710) & (g711) & (g712) & (g713) & (!g60) & (!g61)) + ((g710) & (g711) & (g712) & (g713) & (!g60) & (g61)) + ((g710) & (g711) & (g712) & (g713) & (g60) & (!g61)) + ((g710) & (g711) & (g712) & (g713) & (g60) & (g61)));
	assign g719 = (((!g715) & (!g716) & (!g717) & (g718) & (g60) & (g61)) + ((!g715) & (!g716) & (g717) & (!g718) & (!g60) & (g61)) + ((!g715) & (!g716) & (g717) & (g718) & (!g60) & (g61)) + ((!g715) & (!g716) & (g717) & (g718) & (g60) & (g61)) + ((!g715) & (g716) & (!g717) & (!g718) & (g60) & (!g61)) + ((!g715) & (g716) & (!g717) & (g718) & (g60) & (!g61)) + ((!g715) & (g716) & (!g717) & (g718) & (g60) & (g61)) + ((!g715) & (g716) & (g717) & (!g718) & (!g60) & (g61)) + ((!g715) & (g716) & (g717) & (!g718) & (g60) & (!g61)) + ((!g715) & (g716) & (g717) & (g718) & (!g60) & (g61)) + ((!g715) & (g716) & (g717) & (g718) & (g60) & (!g61)) + ((!g715) & (g716) & (g717) & (g718) & (g60) & (g61)) + ((g715) & (!g716) & (!g717) & (!g718) & (!g60) & (!g61)) + ((g715) & (!g716) & (!g717) & (g718) & (!g60) & (!g61)) + ((g715) & (!g716) & (!g717) & (g718) & (g60) & (g61)) + ((g715) & (!g716) & (g717) & (!g718) & (!g60) & (!g61)) + ((g715) & (!g716) & (g717) & (!g718) & (!g60) & (g61)) + ((g715) & (!g716) & (g717) & (g718) & (!g60) & (!g61)) + ((g715) & (!g716) & (g717) & (g718) & (!g60) & (g61)) + ((g715) & (!g716) & (g717) & (g718) & (g60) & (g61)) + ((g715) & (g716) & (!g717) & (!g718) & (!g60) & (!g61)) + ((g715) & (g716) & (!g717) & (!g718) & (g60) & (!g61)) + ((g715) & (g716) & (!g717) & (g718) & (!g60) & (!g61)) + ((g715) & (g716) & (!g717) & (g718) & (g60) & (!g61)) + ((g715) & (g716) & (!g717) & (g718) & (g60) & (g61)) + ((g715) & (g716) & (g717) & (!g718) & (!g60) & (!g61)) + ((g715) & (g716) & (g717) & (!g718) & (!g60) & (g61)) + ((g715) & (g716) & (g717) & (!g718) & (g60) & (!g61)) + ((g715) & (g716) & (g717) & (g718) & (!g60) & (!g61)) + ((g715) & (g716) & (g717) & (g718) & (!g60) & (g61)) + ((g715) & (g716) & (g717) & (g718) & (g60) & (!g61)) + ((g715) & (g716) & (g717) & (g718) & (g60) & (g61)));
	assign g724 = (((!g720) & (!g721) & (!g722) & (g723) & (g60) & (g61)) + ((!g720) & (!g721) & (g722) & (!g723) & (!g60) & (g61)) + ((!g720) & (!g721) & (g722) & (g723) & (!g60) & (g61)) + ((!g720) & (!g721) & (g722) & (g723) & (g60) & (g61)) + ((!g720) & (g721) & (!g722) & (!g723) & (g60) & (!g61)) + ((!g720) & (g721) & (!g722) & (g723) & (g60) & (!g61)) + ((!g720) & (g721) & (!g722) & (g723) & (g60) & (g61)) + ((!g720) & (g721) & (g722) & (!g723) & (!g60) & (g61)) + ((!g720) & (g721) & (g722) & (!g723) & (g60) & (!g61)) + ((!g720) & (g721) & (g722) & (g723) & (!g60) & (g61)) + ((!g720) & (g721) & (g722) & (g723) & (g60) & (!g61)) + ((!g720) & (g721) & (g722) & (g723) & (g60) & (g61)) + ((g720) & (!g721) & (!g722) & (!g723) & (!g60) & (!g61)) + ((g720) & (!g721) & (!g722) & (g723) & (!g60) & (!g61)) + ((g720) & (!g721) & (!g722) & (g723) & (g60) & (g61)) + ((g720) & (!g721) & (g722) & (!g723) & (!g60) & (!g61)) + ((g720) & (!g721) & (g722) & (!g723) & (!g60) & (g61)) + ((g720) & (!g721) & (g722) & (g723) & (!g60) & (!g61)) + ((g720) & (!g721) & (g722) & (g723) & (!g60) & (g61)) + ((g720) & (!g721) & (g722) & (g723) & (g60) & (g61)) + ((g720) & (g721) & (!g722) & (!g723) & (!g60) & (!g61)) + ((g720) & (g721) & (!g722) & (!g723) & (g60) & (!g61)) + ((g720) & (g721) & (!g722) & (g723) & (!g60) & (!g61)) + ((g720) & (g721) & (!g722) & (g723) & (g60) & (!g61)) + ((g720) & (g721) & (!g722) & (g723) & (g60) & (g61)) + ((g720) & (g721) & (g722) & (!g723) & (!g60) & (!g61)) + ((g720) & (g721) & (g722) & (!g723) & (!g60) & (g61)) + ((g720) & (g721) & (g722) & (!g723) & (g60) & (!g61)) + ((g720) & (g721) & (g722) & (g723) & (!g60) & (!g61)) + ((g720) & (g721) & (g722) & (g723) & (!g60) & (g61)) + ((g720) & (g721) & (g722) & (g723) & (g60) & (!g61)) + ((g720) & (g721) & (g722) & (g723) & (g60) & (g61)));
	assign g729 = (((!g725) & (!g726) & (!g727) & (g728) & (g60) & (g61)) + ((!g725) & (!g726) & (g727) & (!g728) & (!g60) & (g61)) + ((!g725) & (!g726) & (g727) & (g728) & (!g60) & (g61)) + ((!g725) & (!g726) & (g727) & (g728) & (g60) & (g61)) + ((!g725) & (g726) & (!g727) & (!g728) & (g60) & (!g61)) + ((!g725) & (g726) & (!g727) & (g728) & (g60) & (!g61)) + ((!g725) & (g726) & (!g727) & (g728) & (g60) & (g61)) + ((!g725) & (g726) & (g727) & (!g728) & (!g60) & (g61)) + ((!g725) & (g726) & (g727) & (!g728) & (g60) & (!g61)) + ((!g725) & (g726) & (g727) & (g728) & (!g60) & (g61)) + ((!g725) & (g726) & (g727) & (g728) & (g60) & (!g61)) + ((!g725) & (g726) & (g727) & (g728) & (g60) & (g61)) + ((g725) & (!g726) & (!g727) & (!g728) & (!g60) & (!g61)) + ((g725) & (!g726) & (!g727) & (g728) & (!g60) & (!g61)) + ((g725) & (!g726) & (!g727) & (g728) & (g60) & (g61)) + ((g725) & (!g726) & (g727) & (!g728) & (!g60) & (!g61)) + ((g725) & (!g726) & (g727) & (!g728) & (!g60) & (g61)) + ((g725) & (!g726) & (g727) & (g728) & (!g60) & (!g61)) + ((g725) & (!g726) & (g727) & (g728) & (!g60) & (g61)) + ((g725) & (!g726) & (g727) & (g728) & (g60) & (g61)) + ((g725) & (g726) & (!g727) & (!g728) & (!g60) & (!g61)) + ((g725) & (g726) & (!g727) & (!g728) & (g60) & (!g61)) + ((g725) & (g726) & (!g727) & (g728) & (!g60) & (!g61)) + ((g725) & (g726) & (!g727) & (g728) & (g60) & (!g61)) + ((g725) & (g726) & (!g727) & (g728) & (g60) & (g61)) + ((g725) & (g726) & (g727) & (!g728) & (!g60) & (!g61)) + ((g725) & (g726) & (g727) & (!g728) & (!g60) & (g61)) + ((g725) & (g726) & (g727) & (!g728) & (g60) & (!g61)) + ((g725) & (g726) & (g727) & (g728) & (!g60) & (!g61)) + ((g725) & (g726) & (g727) & (g728) & (!g60) & (g61)) + ((g725) & (g726) & (g727) & (g728) & (g60) & (!g61)) + ((g725) & (g726) & (g727) & (g728) & (g60) & (g61)));
	assign g730 = (((!g714) & (!g719) & (!g724) & (g729) & (g42) & (g43)) + ((!g714) & (!g719) & (g724) & (!g729) & (!g42) & (g43)) + ((!g714) & (!g719) & (g724) & (g729) & (!g42) & (g43)) + ((!g714) & (!g719) & (g724) & (g729) & (g42) & (g43)) + ((!g714) & (g719) & (!g724) & (!g729) & (g42) & (!g43)) + ((!g714) & (g719) & (!g724) & (g729) & (g42) & (!g43)) + ((!g714) & (g719) & (!g724) & (g729) & (g42) & (g43)) + ((!g714) & (g719) & (g724) & (!g729) & (!g42) & (g43)) + ((!g714) & (g719) & (g724) & (!g729) & (g42) & (!g43)) + ((!g714) & (g719) & (g724) & (g729) & (!g42) & (g43)) + ((!g714) & (g719) & (g724) & (g729) & (g42) & (!g43)) + ((!g714) & (g719) & (g724) & (g729) & (g42) & (g43)) + ((g714) & (!g719) & (!g724) & (!g729) & (!g42) & (!g43)) + ((g714) & (!g719) & (!g724) & (g729) & (!g42) & (!g43)) + ((g714) & (!g719) & (!g724) & (g729) & (g42) & (g43)) + ((g714) & (!g719) & (g724) & (!g729) & (!g42) & (!g43)) + ((g714) & (!g719) & (g724) & (!g729) & (!g42) & (g43)) + ((g714) & (!g719) & (g724) & (g729) & (!g42) & (!g43)) + ((g714) & (!g719) & (g724) & (g729) & (!g42) & (g43)) + ((g714) & (!g719) & (g724) & (g729) & (g42) & (g43)) + ((g714) & (g719) & (!g724) & (!g729) & (!g42) & (!g43)) + ((g714) & (g719) & (!g724) & (!g729) & (g42) & (!g43)) + ((g714) & (g719) & (!g724) & (g729) & (!g42) & (!g43)) + ((g714) & (g719) & (!g724) & (g729) & (g42) & (!g43)) + ((g714) & (g719) & (!g724) & (g729) & (g42) & (g43)) + ((g714) & (g719) & (g724) & (!g729) & (!g42) & (!g43)) + ((g714) & (g719) & (g724) & (!g729) & (!g42) & (g43)) + ((g714) & (g719) & (g724) & (!g729) & (g42) & (!g43)) + ((g714) & (g719) & (g724) & (g729) & (!g42) & (!g43)) + ((g714) & (g719) & (g724) & (g729) & (!g42) & (g43)) + ((g714) & (g719) & (g724) & (g729) & (g42) & (!g43)) + ((g714) & (g719) & (g724) & (g729) & (g42) & (g43)));
	assign g7263 = (((!g832) & (g1815) & (!g731)) + ((!g832) & (g1815) & (g731)) + ((g832) & (!g1815) & (g731)) + ((g832) & (g1815) & (g731)));
	assign g732 = (((!g34) & (!reset) & (!g730) & (g731)) + ((!g34) & (!reset) & (g730) & (g731)) + ((g34) & (!reset) & (g730) & (!g731)) + ((g34) & (!reset) & (g730) & (g731)));
	assign g737 = (((!g733) & (!g734) & (!g735) & (g736) & (g42) & (g43)) + ((!g733) & (!g734) & (g735) & (!g736) & (!g42) & (g43)) + ((!g733) & (!g734) & (g735) & (g736) & (!g42) & (g43)) + ((!g733) & (!g734) & (g735) & (g736) & (g42) & (g43)) + ((!g733) & (g734) & (!g735) & (!g736) & (g42) & (!g43)) + ((!g733) & (g734) & (!g735) & (g736) & (g42) & (!g43)) + ((!g733) & (g734) & (!g735) & (g736) & (g42) & (g43)) + ((!g733) & (g734) & (g735) & (!g736) & (!g42) & (g43)) + ((!g733) & (g734) & (g735) & (!g736) & (g42) & (!g43)) + ((!g733) & (g734) & (g735) & (g736) & (!g42) & (g43)) + ((!g733) & (g734) & (g735) & (g736) & (g42) & (!g43)) + ((!g733) & (g734) & (g735) & (g736) & (g42) & (g43)) + ((g733) & (!g734) & (!g735) & (!g736) & (!g42) & (!g43)) + ((g733) & (!g734) & (!g735) & (g736) & (!g42) & (!g43)) + ((g733) & (!g734) & (!g735) & (g736) & (g42) & (g43)) + ((g733) & (!g734) & (g735) & (!g736) & (!g42) & (!g43)) + ((g733) & (!g734) & (g735) & (!g736) & (!g42) & (g43)) + ((g733) & (!g734) & (g735) & (g736) & (!g42) & (!g43)) + ((g733) & (!g734) & (g735) & (g736) & (!g42) & (g43)) + ((g733) & (!g734) & (g735) & (g736) & (g42) & (g43)) + ((g733) & (g734) & (!g735) & (!g736) & (!g42) & (!g43)) + ((g733) & (g734) & (!g735) & (!g736) & (g42) & (!g43)) + ((g733) & (g734) & (!g735) & (g736) & (!g42) & (!g43)) + ((g733) & (g734) & (!g735) & (g736) & (g42) & (!g43)) + ((g733) & (g734) & (!g735) & (g736) & (g42) & (g43)) + ((g733) & (g734) & (g735) & (!g736) & (!g42) & (!g43)) + ((g733) & (g734) & (g735) & (!g736) & (!g42) & (g43)) + ((g733) & (g734) & (g735) & (!g736) & (g42) & (!g43)) + ((g733) & (g734) & (g735) & (g736) & (!g42) & (!g43)) + ((g733) & (g734) & (g735) & (g736) & (!g42) & (g43)) + ((g733) & (g734) & (g735) & (g736) & (g42) & (!g43)) + ((g733) & (g734) & (g735) & (g736) & (g42) & (g43)));
	assign g742 = (((!g738) & (!g739) & (!g740) & (g741) & (g42) & (g43)) + ((!g738) & (!g739) & (g740) & (!g741) & (!g42) & (g43)) + ((!g738) & (!g739) & (g740) & (g741) & (!g42) & (g43)) + ((!g738) & (!g739) & (g740) & (g741) & (g42) & (g43)) + ((!g738) & (g739) & (!g740) & (!g741) & (g42) & (!g43)) + ((!g738) & (g739) & (!g740) & (g741) & (g42) & (!g43)) + ((!g738) & (g739) & (!g740) & (g741) & (g42) & (g43)) + ((!g738) & (g739) & (g740) & (!g741) & (!g42) & (g43)) + ((!g738) & (g739) & (g740) & (!g741) & (g42) & (!g43)) + ((!g738) & (g739) & (g740) & (g741) & (!g42) & (g43)) + ((!g738) & (g739) & (g740) & (g741) & (g42) & (!g43)) + ((!g738) & (g739) & (g740) & (g741) & (g42) & (g43)) + ((g738) & (!g739) & (!g740) & (!g741) & (!g42) & (!g43)) + ((g738) & (!g739) & (!g740) & (g741) & (!g42) & (!g43)) + ((g738) & (!g739) & (!g740) & (g741) & (g42) & (g43)) + ((g738) & (!g739) & (g740) & (!g741) & (!g42) & (!g43)) + ((g738) & (!g739) & (g740) & (!g741) & (!g42) & (g43)) + ((g738) & (!g739) & (g740) & (g741) & (!g42) & (!g43)) + ((g738) & (!g739) & (g740) & (g741) & (!g42) & (g43)) + ((g738) & (!g739) & (g740) & (g741) & (g42) & (g43)) + ((g738) & (g739) & (!g740) & (!g741) & (!g42) & (!g43)) + ((g738) & (g739) & (!g740) & (!g741) & (g42) & (!g43)) + ((g738) & (g739) & (!g740) & (g741) & (!g42) & (!g43)) + ((g738) & (g739) & (!g740) & (g741) & (g42) & (!g43)) + ((g738) & (g739) & (!g740) & (g741) & (g42) & (g43)) + ((g738) & (g739) & (g740) & (!g741) & (!g42) & (!g43)) + ((g738) & (g739) & (g740) & (!g741) & (!g42) & (g43)) + ((g738) & (g739) & (g740) & (!g741) & (g42) & (!g43)) + ((g738) & (g739) & (g740) & (g741) & (!g42) & (!g43)) + ((g738) & (g739) & (g740) & (g741) & (!g42) & (g43)) + ((g738) & (g739) & (g740) & (g741) & (g42) & (!g43)) + ((g738) & (g739) & (g740) & (g741) & (g42) & (g43)));
	assign g747 = (((!g743) & (!g744) & (!g745) & (g746) & (g42) & (g43)) + ((!g743) & (!g744) & (g745) & (!g746) & (!g42) & (g43)) + ((!g743) & (!g744) & (g745) & (g746) & (!g42) & (g43)) + ((!g743) & (!g744) & (g745) & (g746) & (g42) & (g43)) + ((!g743) & (g744) & (!g745) & (!g746) & (g42) & (!g43)) + ((!g743) & (g744) & (!g745) & (g746) & (g42) & (!g43)) + ((!g743) & (g744) & (!g745) & (g746) & (g42) & (g43)) + ((!g743) & (g744) & (g745) & (!g746) & (!g42) & (g43)) + ((!g743) & (g744) & (g745) & (!g746) & (g42) & (!g43)) + ((!g743) & (g744) & (g745) & (g746) & (!g42) & (g43)) + ((!g743) & (g744) & (g745) & (g746) & (g42) & (!g43)) + ((!g743) & (g744) & (g745) & (g746) & (g42) & (g43)) + ((g743) & (!g744) & (!g745) & (!g746) & (!g42) & (!g43)) + ((g743) & (!g744) & (!g745) & (g746) & (!g42) & (!g43)) + ((g743) & (!g744) & (!g745) & (g746) & (g42) & (g43)) + ((g743) & (!g744) & (g745) & (!g746) & (!g42) & (!g43)) + ((g743) & (!g744) & (g745) & (!g746) & (!g42) & (g43)) + ((g743) & (!g744) & (g745) & (g746) & (!g42) & (!g43)) + ((g743) & (!g744) & (g745) & (g746) & (!g42) & (g43)) + ((g743) & (!g744) & (g745) & (g746) & (g42) & (g43)) + ((g743) & (g744) & (!g745) & (!g746) & (!g42) & (!g43)) + ((g743) & (g744) & (!g745) & (!g746) & (g42) & (!g43)) + ((g743) & (g744) & (!g745) & (g746) & (!g42) & (!g43)) + ((g743) & (g744) & (!g745) & (g746) & (g42) & (!g43)) + ((g743) & (g744) & (!g745) & (g746) & (g42) & (g43)) + ((g743) & (g744) & (g745) & (!g746) & (!g42) & (!g43)) + ((g743) & (g744) & (g745) & (!g746) & (!g42) & (g43)) + ((g743) & (g744) & (g745) & (!g746) & (g42) & (!g43)) + ((g743) & (g744) & (g745) & (g746) & (!g42) & (!g43)) + ((g743) & (g744) & (g745) & (g746) & (!g42) & (g43)) + ((g743) & (g744) & (g745) & (g746) & (g42) & (!g43)) + ((g743) & (g744) & (g745) & (g746) & (g42) & (g43)));
	assign g752 = (((!g748) & (!g749) & (!g750) & (g751) & (g42) & (g43)) + ((!g748) & (!g749) & (g750) & (!g751) & (!g42) & (g43)) + ((!g748) & (!g749) & (g750) & (g751) & (!g42) & (g43)) + ((!g748) & (!g749) & (g750) & (g751) & (g42) & (g43)) + ((!g748) & (g749) & (!g750) & (!g751) & (g42) & (!g43)) + ((!g748) & (g749) & (!g750) & (g751) & (g42) & (!g43)) + ((!g748) & (g749) & (!g750) & (g751) & (g42) & (g43)) + ((!g748) & (g749) & (g750) & (!g751) & (!g42) & (g43)) + ((!g748) & (g749) & (g750) & (!g751) & (g42) & (!g43)) + ((!g748) & (g749) & (g750) & (g751) & (!g42) & (g43)) + ((!g748) & (g749) & (g750) & (g751) & (g42) & (!g43)) + ((!g748) & (g749) & (g750) & (g751) & (g42) & (g43)) + ((g748) & (!g749) & (!g750) & (!g751) & (!g42) & (!g43)) + ((g748) & (!g749) & (!g750) & (g751) & (!g42) & (!g43)) + ((g748) & (!g749) & (!g750) & (g751) & (g42) & (g43)) + ((g748) & (!g749) & (g750) & (!g751) & (!g42) & (!g43)) + ((g748) & (!g749) & (g750) & (!g751) & (!g42) & (g43)) + ((g748) & (!g749) & (g750) & (g751) & (!g42) & (!g43)) + ((g748) & (!g749) & (g750) & (g751) & (!g42) & (g43)) + ((g748) & (!g749) & (g750) & (g751) & (g42) & (g43)) + ((g748) & (g749) & (!g750) & (!g751) & (!g42) & (!g43)) + ((g748) & (g749) & (!g750) & (!g751) & (g42) & (!g43)) + ((g748) & (g749) & (!g750) & (g751) & (!g42) & (!g43)) + ((g748) & (g749) & (!g750) & (g751) & (g42) & (!g43)) + ((g748) & (g749) & (!g750) & (g751) & (g42) & (g43)) + ((g748) & (g749) & (g750) & (!g751) & (!g42) & (!g43)) + ((g748) & (g749) & (g750) & (!g751) & (!g42) & (g43)) + ((g748) & (g749) & (g750) & (!g751) & (g42) & (!g43)) + ((g748) & (g749) & (g750) & (g751) & (!g42) & (!g43)) + ((g748) & (g749) & (g750) & (g751) & (!g42) & (g43)) + ((g748) & (g749) & (g750) & (g751) & (g42) & (!g43)) + ((g748) & (g749) & (g750) & (g751) & (g42) & (g43)));
	assign g753 = (((!g737) & (!g742) & (!g747) & (g752) & (g60) & (g61)) + ((!g737) & (!g742) & (g747) & (!g752) & (!g60) & (g61)) + ((!g737) & (!g742) & (g747) & (g752) & (!g60) & (g61)) + ((!g737) & (!g742) & (g747) & (g752) & (g60) & (g61)) + ((!g737) & (g742) & (!g747) & (!g752) & (g60) & (!g61)) + ((!g737) & (g742) & (!g747) & (g752) & (g60) & (!g61)) + ((!g737) & (g742) & (!g747) & (g752) & (g60) & (g61)) + ((!g737) & (g742) & (g747) & (!g752) & (!g60) & (g61)) + ((!g737) & (g742) & (g747) & (!g752) & (g60) & (!g61)) + ((!g737) & (g742) & (g747) & (g752) & (!g60) & (g61)) + ((!g737) & (g742) & (g747) & (g752) & (g60) & (!g61)) + ((!g737) & (g742) & (g747) & (g752) & (g60) & (g61)) + ((g737) & (!g742) & (!g747) & (!g752) & (!g60) & (!g61)) + ((g737) & (!g742) & (!g747) & (g752) & (!g60) & (!g61)) + ((g737) & (!g742) & (!g747) & (g752) & (g60) & (g61)) + ((g737) & (!g742) & (g747) & (!g752) & (!g60) & (!g61)) + ((g737) & (!g742) & (g747) & (!g752) & (!g60) & (g61)) + ((g737) & (!g742) & (g747) & (g752) & (!g60) & (!g61)) + ((g737) & (!g742) & (g747) & (g752) & (!g60) & (g61)) + ((g737) & (!g742) & (g747) & (g752) & (g60) & (g61)) + ((g737) & (g742) & (!g747) & (!g752) & (!g60) & (!g61)) + ((g737) & (g742) & (!g747) & (!g752) & (g60) & (!g61)) + ((g737) & (g742) & (!g747) & (g752) & (!g60) & (!g61)) + ((g737) & (g742) & (!g747) & (g752) & (g60) & (!g61)) + ((g737) & (g742) & (!g747) & (g752) & (g60) & (g61)) + ((g737) & (g742) & (g747) & (!g752) & (!g60) & (!g61)) + ((g737) & (g742) & (g747) & (!g752) & (!g60) & (g61)) + ((g737) & (g742) & (g747) & (!g752) & (g60) & (!g61)) + ((g737) & (g742) & (g747) & (g752) & (!g60) & (!g61)) + ((g737) & (g742) & (g747) & (g752) & (!g60) & (g61)) + ((g737) & (g742) & (g747) & (g752) & (g60) & (!g61)) + ((g737) & (g742) & (g747) & (g752) & (g60) & (g61)));
	assign g7264 = (((!g832) & (g1849) & (!g754)) + ((!g832) & (g1849) & (g754)) + ((g832) & (!g1849) & (g754)) + ((g832) & (g1849) & (g754)));
	assign g755 = (((!g34) & (!reset) & (!g753) & (g754)) + ((!g34) & (!reset) & (g753) & (g754)) + ((g34) & (!reset) & (g753) & (!g754)) + ((g34) & (!reset) & (g753) & (g754)));
	assign g760 = (((!g756) & (!g757) & (!g758) & (g759) & (g60) & (g61)) + ((!g756) & (!g757) & (g758) & (!g759) & (!g60) & (g61)) + ((!g756) & (!g757) & (g758) & (g759) & (!g60) & (g61)) + ((!g756) & (!g757) & (g758) & (g759) & (g60) & (g61)) + ((!g756) & (g757) & (!g758) & (!g759) & (g60) & (!g61)) + ((!g756) & (g757) & (!g758) & (g759) & (g60) & (!g61)) + ((!g756) & (g757) & (!g758) & (g759) & (g60) & (g61)) + ((!g756) & (g757) & (g758) & (!g759) & (!g60) & (g61)) + ((!g756) & (g757) & (g758) & (!g759) & (g60) & (!g61)) + ((!g756) & (g757) & (g758) & (g759) & (!g60) & (g61)) + ((!g756) & (g757) & (g758) & (g759) & (g60) & (!g61)) + ((!g756) & (g757) & (g758) & (g759) & (g60) & (g61)) + ((g756) & (!g757) & (!g758) & (!g759) & (!g60) & (!g61)) + ((g756) & (!g757) & (!g758) & (g759) & (!g60) & (!g61)) + ((g756) & (!g757) & (!g758) & (g759) & (g60) & (g61)) + ((g756) & (!g757) & (g758) & (!g759) & (!g60) & (!g61)) + ((g756) & (!g757) & (g758) & (!g759) & (!g60) & (g61)) + ((g756) & (!g757) & (g758) & (g759) & (!g60) & (!g61)) + ((g756) & (!g757) & (g758) & (g759) & (!g60) & (g61)) + ((g756) & (!g757) & (g758) & (g759) & (g60) & (g61)) + ((g756) & (g757) & (!g758) & (!g759) & (!g60) & (!g61)) + ((g756) & (g757) & (!g758) & (!g759) & (g60) & (!g61)) + ((g756) & (g757) & (!g758) & (g759) & (!g60) & (!g61)) + ((g756) & (g757) & (!g758) & (g759) & (g60) & (!g61)) + ((g756) & (g757) & (!g758) & (g759) & (g60) & (g61)) + ((g756) & (g757) & (g758) & (!g759) & (!g60) & (!g61)) + ((g756) & (g757) & (g758) & (!g759) & (!g60) & (g61)) + ((g756) & (g757) & (g758) & (!g759) & (g60) & (!g61)) + ((g756) & (g757) & (g758) & (g759) & (!g60) & (!g61)) + ((g756) & (g757) & (g758) & (g759) & (!g60) & (g61)) + ((g756) & (g757) & (g758) & (g759) & (g60) & (!g61)) + ((g756) & (g757) & (g758) & (g759) & (g60) & (g61)));
	assign g765 = (((!g761) & (!g762) & (!g763) & (g764) & (g60) & (g61)) + ((!g761) & (!g762) & (g763) & (!g764) & (!g60) & (g61)) + ((!g761) & (!g762) & (g763) & (g764) & (!g60) & (g61)) + ((!g761) & (!g762) & (g763) & (g764) & (g60) & (g61)) + ((!g761) & (g762) & (!g763) & (!g764) & (g60) & (!g61)) + ((!g761) & (g762) & (!g763) & (g764) & (g60) & (!g61)) + ((!g761) & (g762) & (!g763) & (g764) & (g60) & (g61)) + ((!g761) & (g762) & (g763) & (!g764) & (!g60) & (g61)) + ((!g761) & (g762) & (g763) & (!g764) & (g60) & (!g61)) + ((!g761) & (g762) & (g763) & (g764) & (!g60) & (g61)) + ((!g761) & (g762) & (g763) & (g764) & (g60) & (!g61)) + ((!g761) & (g762) & (g763) & (g764) & (g60) & (g61)) + ((g761) & (!g762) & (!g763) & (!g764) & (!g60) & (!g61)) + ((g761) & (!g762) & (!g763) & (g764) & (!g60) & (!g61)) + ((g761) & (!g762) & (!g763) & (g764) & (g60) & (g61)) + ((g761) & (!g762) & (g763) & (!g764) & (!g60) & (!g61)) + ((g761) & (!g762) & (g763) & (!g764) & (!g60) & (g61)) + ((g761) & (!g762) & (g763) & (g764) & (!g60) & (!g61)) + ((g761) & (!g762) & (g763) & (g764) & (!g60) & (g61)) + ((g761) & (!g762) & (g763) & (g764) & (g60) & (g61)) + ((g761) & (g762) & (!g763) & (!g764) & (!g60) & (!g61)) + ((g761) & (g762) & (!g763) & (!g764) & (g60) & (!g61)) + ((g761) & (g762) & (!g763) & (g764) & (!g60) & (!g61)) + ((g761) & (g762) & (!g763) & (g764) & (g60) & (!g61)) + ((g761) & (g762) & (!g763) & (g764) & (g60) & (g61)) + ((g761) & (g762) & (g763) & (!g764) & (!g60) & (!g61)) + ((g761) & (g762) & (g763) & (!g764) & (!g60) & (g61)) + ((g761) & (g762) & (g763) & (!g764) & (g60) & (!g61)) + ((g761) & (g762) & (g763) & (g764) & (!g60) & (!g61)) + ((g761) & (g762) & (g763) & (g764) & (!g60) & (g61)) + ((g761) & (g762) & (g763) & (g764) & (g60) & (!g61)) + ((g761) & (g762) & (g763) & (g764) & (g60) & (g61)));
	assign g770 = (((!g766) & (!g767) & (!g768) & (g769) & (g60) & (g61)) + ((!g766) & (!g767) & (g768) & (!g769) & (!g60) & (g61)) + ((!g766) & (!g767) & (g768) & (g769) & (!g60) & (g61)) + ((!g766) & (!g767) & (g768) & (g769) & (g60) & (g61)) + ((!g766) & (g767) & (!g768) & (!g769) & (g60) & (!g61)) + ((!g766) & (g767) & (!g768) & (g769) & (g60) & (!g61)) + ((!g766) & (g767) & (!g768) & (g769) & (g60) & (g61)) + ((!g766) & (g767) & (g768) & (!g769) & (!g60) & (g61)) + ((!g766) & (g767) & (g768) & (!g769) & (g60) & (!g61)) + ((!g766) & (g767) & (g768) & (g769) & (!g60) & (g61)) + ((!g766) & (g767) & (g768) & (g769) & (g60) & (!g61)) + ((!g766) & (g767) & (g768) & (g769) & (g60) & (g61)) + ((g766) & (!g767) & (!g768) & (!g769) & (!g60) & (!g61)) + ((g766) & (!g767) & (!g768) & (g769) & (!g60) & (!g61)) + ((g766) & (!g767) & (!g768) & (g769) & (g60) & (g61)) + ((g766) & (!g767) & (g768) & (!g769) & (!g60) & (!g61)) + ((g766) & (!g767) & (g768) & (!g769) & (!g60) & (g61)) + ((g766) & (!g767) & (g768) & (g769) & (!g60) & (!g61)) + ((g766) & (!g767) & (g768) & (g769) & (!g60) & (g61)) + ((g766) & (!g767) & (g768) & (g769) & (g60) & (g61)) + ((g766) & (g767) & (!g768) & (!g769) & (!g60) & (!g61)) + ((g766) & (g767) & (!g768) & (!g769) & (g60) & (!g61)) + ((g766) & (g767) & (!g768) & (g769) & (!g60) & (!g61)) + ((g766) & (g767) & (!g768) & (g769) & (g60) & (!g61)) + ((g766) & (g767) & (!g768) & (g769) & (g60) & (g61)) + ((g766) & (g767) & (g768) & (!g769) & (!g60) & (!g61)) + ((g766) & (g767) & (g768) & (!g769) & (!g60) & (g61)) + ((g766) & (g767) & (g768) & (!g769) & (g60) & (!g61)) + ((g766) & (g767) & (g768) & (g769) & (!g60) & (!g61)) + ((g766) & (g767) & (g768) & (g769) & (!g60) & (g61)) + ((g766) & (g767) & (g768) & (g769) & (g60) & (!g61)) + ((g766) & (g767) & (g768) & (g769) & (g60) & (g61)));
	assign g775 = (((!g771) & (!g772) & (!g773) & (g774) & (g60) & (g61)) + ((!g771) & (!g772) & (g773) & (!g774) & (!g60) & (g61)) + ((!g771) & (!g772) & (g773) & (g774) & (!g60) & (g61)) + ((!g771) & (!g772) & (g773) & (g774) & (g60) & (g61)) + ((!g771) & (g772) & (!g773) & (!g774) & (g60) & (!g61)) + ((!g771) & (g772) & (!g773) & (g774) & (g60) & (!g61)) + ((!g771) & (g772) & (!g773) & (g774) & (g60) & (g61)) + ((!g771) & (g772) & (g773) & (!g774) & (!g60) & (g61)) + ((!g771) & (g772) & (g773) & (!g774) & (g60) & (!g61)) + ((!g771) & (g772) & (g773) & (g774) & (!g60) & (g61)) + ((!g771) & (g772) & (g773) & (g774) & (g60) & (!g61)) + ((!g771) & (g772) & (g773) & (g774) & (g60) & (g61)) + ((g771) & (!g772) & (!g773) & (!g774) & (!g60) & (!g61)) + ((g771) & (!g772) & (!g773) & (g774) & (!g60) & (!g61)) + ((g771) & (!g772) & (!g773) & (g774) & (g60) & (g61)) + ((g771) & (!g772) & (g773) & (!g774) & (!g60) & (!g61)) + ((g771) & (!g772) & (g773) & (!g774) & (!g60) & (g61)) + ((g771) & (!g772) & (g773) & (g774) & (!g60) & (!g61)) + ((g771) & (!g772) & (g773) & (g774) & (!g60) & (g61)) + ((g771) & (!g772) & (g773) & (g774) & (g60) & (g61)) + ((g771) & (g772) & (!g773) & (!g774) & (!g60) & (!g61)) + ((g771) & (g772) & (!g773) & (!g774) & (g60) & (!g61)) + ((g771) & (g772) & (!g773) & (g774) & (!g60) & (!g61)) + ((g771) & (g772) & (!g773) & (g774) & (g60) & (!g61)) + ((g771) & (g772) & (!g773) & (g774) & (g60) & (g61)) + ((g771) & (g772) & (g773) & (!g774) & (!g60) & (!g61)) + ((g771) & (g772) & (g773) & (!g774) & (!g60) & (g61)) + ((g771) & (g772) & (g773) & (!g774) & (g60) & (!g61)) + ((g771) & (g772) & (g773) & (g774) & (!g60) & (!g61)) + ((g771) & (g772) & (g773) & (g774) & (!g60) & (g61)) + ((g771) & (g772) & (g773) & (g774) & (g60) & (!g61)) + ((g771) & (g772) & (g773) & (g774) & (g60) & (g61)));
	assign g776 = (((!g760) & (!g765) & (!g770) & (g775) & (g42) & (g43)) + ((!g760) & (!g765) & (g770) & (!g775) & (!g42) & (g43)) + ((!g760) & (!g765) & (g770) & (g775) & (!g42) & (g43)) + ((!g760) & (!g765) & (g770) & (g775) & (g42) & (g43)) + ((!g760) & (g765) & (!g770) & (!g775) & (g42) & (!g43)) + ((!g760) & (g765) & (!g770) & (g775) & (g42) & (!g43)) + ((!g760) & (g765) & (!g770) & (g775) & (g42) & (g43)) + ((!g760) & (g765) & (g770) & (!g775) & (!g42) & (g43)) + ((!g760) & (g765) & (g770) & (!g775) & (g42) & (!g43)) + ((!g760) & (g765) & (g770) & (g775) & (!g42) & (g43)) + ((!g760) & (g765) & (g770) & (g775) & (g42) & (!g43)) + ((!g760) & (g765) & (g770) & (g775) & (g42) & (g43)) + ((g760) & (!g765) & (!g770) & (!g775) & (!g42) & (!g43)) + ((g760) & (!g765) & (!g770) & (g775) & (!g42) & (!g43)) + ((g760) & (!g765) & (!g770) & (g775) & (g42) & (g43)) + ((g760) & (!g765) & (g770) & (!g775) & (!g42) & (!g43)) + ((g760) & (!g765) & (g770) & (!g775) & (!g42) & (g43)) + ((g760) & (!g765) & (g770) & (g775) & (!g42) & (!g43)) + ((g760) & (!g765) & (g770) & (g775) & (!g42) & (g43)) + ((g760) & (!g765) & (g770) & (g775) & (g42) & (g43)) + ((g760) & (g765) & (!g770) & (!g775) & (!g42) & (!g43)) + ((g760) & (g765) & (!g770) & (!g775) & (g42) & (!g43)) + ((g760) & (g765) & (!g770) & (g775) & (!g42) & (!g43)) + ((g760) & (g765) & (!g770) & (g775) & (g42) & (!g43)) + ((g760) & (g765) & (!g770) & (g775) & (g42) & (g43)) + ((g760) & (g765) & (g770) & (!g775) & (!g42) & (!g43)) + ((g760) & (g765) & (g770) & (!g775) & (!g42) & (g43)) + ((g760) & (g765) & (g770) & (!g775) & (g42) & (!g43)) + ((g760) & (g765) & (g770) & (g775) & (!g42) & (!g43)) + ((g760) & (g765) & (g770) & (g775) & (!g42) & (g43)) + ((g760) & (g765) & (g770) & (g775) & (g42) & (!g43)) + ((g760) & (g765) & (g770) & (g775) & (g42) & (g43)));
	assign g7265 = (((!g832) & (g1882) & (!g777)) + ((!g832) & (g1882) & (g777)) + ((g832) & (!g1882) & (g777)) + ((g832) & (g1882) & (g777)));
	assign g778 = (((!g34) & (!reset) & (!g776) & (g777)) + ((!g34) & (!reset) & (g776) & (g777)) + ((g34) & (!reset) & (g776) & (!g777)) + ((g34) & (!reset) & (g776) & (g777)));
	assign g780 = (((g43) & (g60) & (g61)));
	assign g781 = (((g42) & (g780)));
	assign g782 = (((!g34) & (g36) & (!g781)) + ((!g34) & (g36) & (g781)) + ((g34) & (g36) & (!g781)));
	assign g783 = (((!g34) & (!g35) & (!reset) & (!g779) & (!data_req) & (g782)) + ((!g34) & (!g35) & (!reset) & (!g779) & (data_req) & (g782)) + ((!g34) & (!g35) & (!reset) & (g779) & (!data_req) & (g782)) + ((!g34) & (!g35) & (!reset) & (g779) & (data_req) & (g782)) + ((!g34) & (g35) & (!reset) & (!g779) & (!data_req) & (g782)) + ((!g34) & (g35) & (!reset) & (!g779) & (data_req) & (g782)) + ((!g34) & (g35) & (!reset) & (g779) & (!data_req) & (g782)) + ((!g34) & (g35) & (!reset) & (g779) & (data_req) & (g782)) + ((g34) & (!g35) & (!reset) & (!g779) & (!data_req) & (g782)) + ((g34) & (!g35) & (!reset) & (!g779) & (data_req) & (g782)) + ((g34) & (!g35) & (!reset) & (g779) & (!data_req) & (!g782)) + ((g34) & (!g35) & (!reset) & (g779) & (!data_req) & (g782)) + ((g34) & (!g35) & (!reset) & (g779) & (data_req) & (g782)) + ((g34) & (g35) & (!reset) & (!g779) & (!data_req) & (!g782)) + ((g34) & (g35) & (!reset) & (!g779) & (!data_req) & (g782)) + ((g34) & (g35) & (!reset) & (!g779) & (data_req) & (!g782)) + ((g34) & (g35) & (!reset) & (!g779) & (data_req) & (g782)) + ((g34) & (g35) & (!reset) & (g779) & (!data_req) & (!g782)) + ((g34) & (g35) & (!reset) & (g779) & (!data_req) & (g782)) + ((g34) & (g35) & (!reset) & (g779) & (data_req) & (!g782)) + ((g34) & (g35) & (!reset) & (g779) & (data_req) & (g782)));
	assign g784 = (((!g34) & (!g35) & (!g36) & (!reset) & (!g781) & (data_req)) + ((!g34) & (!g35) & (!g36) & (!reset) & (g781) & (data_req)) + ((!g34) & (!g35) & (g36) & (!reset) & (!g781) & (!data_req)) + ((!g34) & (!g35) & (g36) & (!reset) & (g781) & (!data_req)) + ((!g34) & (g35) & (!g36) & (!reset) & (!g781) & (!data_req)) + ((!g34) & (g35) & (!g36) & (!reset) & (!g781) & (data_req)) + ((!g34) & (g35) & (!g36) & (!reset) & (g781) & (!data_req)) + ((!g34) & (g35) & (!g36) & (!reset) & (g781) & (data_req)) + ((!g34) & (g35) & (g36) & (!reset) & (!g781) & (!data_req)) + ((!g34) & (g35) & (g36) & (!reset) & (g781) & (!data_req)) + ((g34) & (!g35) & (!g36) & (!reset) & (!g781) & (data_req)) + ((g34) & (!g35) & (!g36) & (!reset) & (g781) & (data_req)) + ((g34) & (!g35) & (g36) & (!reset) & (!g781) & (!data_req)) + ((g34) & (!g35) & (g36) & (!reset) & (g781) & (data_req)) + ((g34) & (g35) & (!g36) & (!reset) & (!g781) & (!data_req)) + ((g34) & (g35) & (!g36) & (!reset) & (g781) & (!data_req)) + ((g34) & (g35) & (g36) & (!reset) & (!g781) & (!data_req)) + ((g34) & (g35) & (g36) & (!reset) & (!g781) & (data_req)) + ((g34) & (g35) & (g36) & (!reset) & (g781) & (!data_req)) + ((g34) & (g35) & (g36) & (!reset) & (g781) & (data_req)));
	assign g785 = (((!g34) & (!g35) & (g36)) + ((!g34) & (g35) & (g36)) + ((g34) & (g35) & (!g36)));
	assign g786 = (((g35) & (g36)));
	assign g787 = (((g36) & (!g781)));
	assign g788 = (((!reset) & (!g785) & (!g786) & (!g787) & (!g779) & (!data_req)) + ((!reset) & (!g785) & (!g786) & (!g787) & (!g779) & (data_req)) + ((!reset) & (!g785) & (!g786) & (g787) & (!g779) & (data_req)) + ((!reset) & (!g785) & (!g786) & (g787) & (g779) & (data_req)) + ((!reset) & (!g785) & (g786) & (!g787) & (!g779) & (!data_req)) + ((!reset) & (!g785) & (g786) & (!g787) & (!g779) & (data_req)) + ((!reset) & (!g785) & (g786) & (!g787) & (g779) & (!data_req)) + ((!reset) & (!g785) & (g786) & (!g787) & (g779) & (data_req)) + ((!reset) & (!g785) & (g786) & (g787) & (!g779) & (!data_req)) + ((!reset) & (!g785) & (g786) & (g787) & (!g779) & (data_req)) + ((!reset) & (!g785) & (g786) & (g787) & (g779) & (!data_req)) + ((!reset) & (!g785) & (g786) & (g787) & (g779) & (data_req)) + ((!reset) & (g785) & (!g786) & (!g787) & (!g779) & (data_req)) + ((!reset) & (g785) & (!g786) & (!g787) & (g779) & (data_req)) + ((!reset) & (g785) & (!g786) & (g787) & (!g779) & (data_req)) + ((!reset) & (g785) & (!g786) & (g787) & (g779) & (data_req)) + ((!reset) & (g785) & (g786) & (!g787) & (!g779) & (data_req)) + ((!reset) & (g785) & (g786) & (!g787) & (g779) & (data_req)) + ((!reset) & (g785) & (g786) & (g787) & (!g779) & (data_req)) + ((!reset) & (g785) & (g786) & (g787) & (g779) & (data_req)));
	assign g789 = (((!g34) & (!g36) & (!reset) & (g38) & (!g63)) + ((!g34) & (!g36) & (!reset) & (g38) & (g63)) + ((!g34) & (g36) & (!reset) & (!g38) & (g63)) + ((!g34) & (g36) & (!reset) & (g38) & (g63)) + ((g34) & (!g36) & (!reset) & (g38) & (!g63)) + ((g34) & (!g36) & (!reset) & (g38) & (g63)) + ((g34) & (g36) & (!reset) & (g38) & (!g63)) + ((g34) & (g36) & (!reset) & (g38) & (g63)));
	assign g7266 = (((!g832) & (g1885) & (!g790)) + ((!g832) & (g1885) & (g790)) + ((g832) & (!g1885) & (g790)) + ((g832) & (g1885) & (g790)));
	assign g791 = (((!g34) & (!g36) & (!reset) & (g39) & (!g790)) + ((!g34) & (!g36) & (!reset) & (g39) & (g790)) + ((!g34) & (g36) & (!reset) & (!g39) & (g790)) + ((!g34) & (g36) & (!reset) & (g39) & (g790)) + ((g34) & (!g36) & (!reset) & (g39) & (!g790)) + ((g34) & (!g36) & (!reset) & (g39) & (g790)) + ((g34) & (g36) & (!reset) & (g39) & (!g790)) + ((g34) & (g36) & (!reset) & (g39) & (g790)));
	assign g7267 = (((!g832) & (g1887) & (!g792)) + ((!g832) & (g1887) & (g792)) + ((g832) & (!g1887) & (g792)) + ((g832) & (g1887) & (g792)));
	assign g793 = (((!g34) & (!g36) & (!reset) & (g40) & (!g792)) + ((!g34) & (!g36) & (!reset) & (g40) & (g792)) + ((!g34) & (g36) & (!reset) & (!g40) & (g792)) + ((!g34) & (g36) & (!reset) & (g40) & (g792)) + ((g34) & (!g36) & (!reset) & (g40) & (!g792)) + ((g34) & (!g36) & (!reset) & (g40) & (g792)) + ((g34) & (g36) & (!reset) & (g40) & (!g792)) + ((g34) & (g36) & (!reset) & (g40) & (g792)));
	assign g7268 = (((!g832) & (g1889) & (!g794)) + ((!g832) & (g1889) & (g794)) + ((g832) & (!g1889) & (g794)) + ((g832) & (g1889) & (g794)));
	assign g795 = (((!g34) & (!g36) & (!reset) & (g41) & (!g794)) + ((!g34) & (!g36) & (!reset) & (g41) & (g794)) + ((!g34) & (g36) & (!reset) & (!g41) & (g794)) + ((!g34) & (g36) & (!reset) & (g41) & (g794)) + ((g34) & (!g36) & (!reset) & (g41) & (!g794)) + ((g34) & (!g36) & (!reset) & (g41) & (g794)) + ((g34) & (g36) & (!reset) & (g41) & (!g794)) + ((g34) & (g36) & (!reset) & (g41) & (g794)));
	assign g796 = (((!g34) & (g35) & (g36) & (!reset) & (!g42) & (g780)) + ((!g34) & (g35) & (g36) & (!reset) & (g42) & (!g780)) + ((g34) & (!g35) & (g36) & (!reset) & (!g42) & (g780)) + ((g34) & (!g35) & (g36) & (!reset) & (g42) & (!g780)) + ((g34) & (g35) & (g36) & (!reset) & (!g42) & (g780)) + ((g34) & (g35) & (g36) & (!reset) & (g42) & (!g780)));
	assign g797 = (((g34) & (g35) & (!reset)));
	assign g798 = (((!g43) & (g60) & (g61)) + ((g43) & (!g60) & (!g61)) + ((g43) & (!g60) & (g61)) + ((g43) & (g60) & (!g61)));
	assign g799 = (((!g34) & (g35) & (g36) & (!reset) & (!g781) & (g798)) + ((!g34) & (g35) & (g36) & (!reset) & (g781) & (g798)) + ((g34) & (!g35) & (g36) & (!reset) & (!g781) & (g798)) + ((g34) & (g35) & (g36) & (!reset) & (!g781) & (g798)));
	assign g7269 = (((!g832) & (g1891) & (!g800)) + ((!g832) & (g1891) & (g800)) + ((g832) & (!g1891) & (g800)) + ((g832) & (g1891) & (g800)));
	assign g801 = (((!g34) & (!g36) & (!reset) & (g45) & (!g800)) + ((!g34) & (!g36) & (!reset) & (g45) & (g800)) + ((!g34) & (g36) & (!reset) & (!g45) & (g800)) + ((!g34) & (g36) & (!reset) & (g45) & (g800)) + ((g34) & (!g36) & (!reset) & (g45) & (!g800)) + ((g34) & (!g36) & (!reset) & (g45) & (g800)) + ((g34) & (g36) & (!reset) & (g45) & (!g800)) + ((g34) & (g36) & (!reset) & (g45) & (g800)));
	assign g7270 = (((!g832) & (g1893) & (!g802)) + ((!g832) & (g1893) & (g802)) + ((g832) & (!g1893) & (g802)) + ((g832) & (g1893) & (g802)));
	assign g803 = (((!g34) & (!g36) & (!reset) & (g46) & (!g802)) + ((!g34) & (!g36) & (!reset) & (g46) & (g802)) + ((!g34) & (g36) & (!reset) & (!g46) & (g802)) + ((!g34) & (g36) & (!reset) & (g46) & (g802)) + ((g34) & (!g36) & (!reset) & (g46) & (!g802)) + ((g34) & (!g36) & (!reset) & (g46) & (g802)) + ((g34) & (g36) & (!reset) & (g46) & (!g802)) + ((g34) & (g36) & (!reset) & (g46) & (g802)));
	assign g7271 = (((!g832) & (g1895) & (!g804)) + ((!g832) & (g1895) & (g804)) + ((g832) & (!g1895) & (g804)) + ((g832) & (g1895) & (g804)));
	assign g805 = (((!g34) & (!g36) & (!reset) & (g47) & (!g804)) + ((!g34) & (!g36) & (!reset) & (g47) & (g804)) + ((!g34) & (g36) & (!reset) & (!g47) & (g804)) + ((!g34) & (g36) & (!reset) & (g47) & (g804)) + ((g34) & (!g36) & (!reset) & (g47) & (!g804)) + ((g34) & (!g36) & (!reset) & (g47) & (g804)) + ((g34) & (g36) & (!reset) & (g47) & (!g804)) + ((g34) & (g36) & (!reset) & (g47) & (g804)));
	assign g7272 = (((!g832) & (g1897) & (!g806)) + ((!g832) & (g1897) & (g806)) + ((g832) & (!g1897) & (g806)) + ((g832) & (g1897) & (g806)));
	assign g807 = (((!g34) & (!g36) & (!reset) & (g48) & (!g806)) + ((!g34) & (!g36) & (!reset) & (g48) & (g806)) + ((!g34) & (g36) & (!reset) & (!g48) & (g806)) + ((!g34) & (g36) & (!reset) & (g48) & (g806)) + ((g34) & (!g36) & (!reset) & (g48) & (!g806)) + ((g34) & (!g36) & (!reset) & (g48) & (g806)) + ((g34) & (g36) & (!reset) & (g48) & (!g806)) + ((g34) & (g36) & (!reset) & (g48) & (g806)));
	assign g7273 = (((!g832) & (g1899) & (!g808)) + ((!g832) & (g1899) & (g808)) + ((g832) & (!g1899) & (g808)) + ((g832) & (g1899) & (g808)));
	assign g809 = (((!g34) & (!g36) & (!reset) & (g50) & (!g808)) + ((!g34) & (!g36) & (!reset) & (g50) & (g808)) + ((!g34) & (g36) & (!reset) & (!g50) & (g808)) + ((!g34) & (g36) & (!reset) & (g50) & (g808)) + ((g34) & (!g36) & (!reset) & (g50) & (!g808)) + ((g34) & (!g36) & (!reset) & (g50) & (g808)) + ((g34) & (g36) & (!reset) & (g50) & (!g808)) + ((g34) & (g36) & (!reset) & (g50) & (g808)));
	assign g7274 = (((!g832) & (g1901) & (!g810)) + ((!g832) & (g1901) & (g810)) + ((g832) & (!g1901) & (g810)) + ((g832) & (g1901) & (g810)));
	assign g811 = (((!g34) & (!g36) & (!reset) & (g51) & (!g810)) + ((!g34) & (!g36) & (!reset) & (g51) & (g810)) + ((!g34) & (g36) & (!reset) & (!g51) & (g810)) + ((!g34) & (g36) & (!reset) & (g51) & (g810)) + ((g34) & (!g36) & (!reset) & (g51) & (!g810)) + ((g34) & (!g36) & (!reset) & (g51) & (g810)) + ((g34) & (g36) & (!reset) & (g51) & (!g810)) + ((g34) & (g36) & (!reset) & (g51) & (g810)));
	assign g7275 = (((!g832) & (g1903) & (!g812)) + ((!g832) & (g1903) & (g812)) + ((g832) & (!g1903) & (g812)) + ((g832) & (g1903) & (g812)));
	assign g813 = (((!g34) & (!g36) & (!reset) & (g52) & (!g812)) + ((!g34) & (!g36) & (!reset) & (g52) & (g812)) + ((!g34) & (g36) & (!reset) & (!g52) & (g812)) + ((!g34) & (g36) & (!reset) & (g52) & (g812)) + ((g34) & (!g36) & (!reset) & (g52) & (!g812)) + ((g34) & (!g36) & (!reset) & (g52) & (g812)) + ((g34) & (g36) & (!reset) & (g52) & (!g812)) + ((g34) & (g36) & (!reset) & (g52) & (g812)));
	assign g7276 = (((!g832) & (g1905) & (!g814)) + ((!g832) & (g1905) & (g814)) + ((g832) & (!g1905) & (g814)) + ((g832) & (g1905) & (g814)));
	assign g815 = (((!g34) & (!g36) & (!reset) & (g53) & (!g814)) + ((!g34) & (!g36) & (!reset) & (g53) & (g814)) + ((!g34) & (g36) & (!reset) & (!g53) & (g814)) + ((!g34) & (g36) & (!reset) & (g53) & (g814)) + ((g34) & (!g36) & (!reset) & (g53) & (!g814)) + ((g34) & (!g36) & (!reset) & (g53) & (g814)) + ((g34) & (g36) & (!reset) & (g53) & (!g814)) + ((g34) & (g36) & (!reset) & (g53) & (g814)));
	assign g7277 = (((!g832) & (g1907) & (!g816)) + ((!g832) & (g1907) & (g816)) + ((g832) & (!g1907) & (g816)) + ((g832) & (g1907) & (g816)));
	assign g817 = (((!g34) & (!g36) & (!reset) & (g55) & (!g816)) + ((!g34) & (!g36) & (!reset) & (g55) & (g816)) + ((!g34) & (g36) & (!reset) & (!g55) & (g816)) + ((!g34) & (g36) & (!reset) & (g55) & (g816)) + ((g34) & (!g36) & (!reset) & (g55) & (!g816)) + ((g34) & (!g36) & (!reset) & (g55) & (g816)) + ((g34) & (g36) & (!reset) & (g55) & (!g816)) + ((g34) & (g36) & (!reset) & (g55) & (g816)));
	assign g7278 = (((!g832) & (g1909) & (!g818)) + ((!g832) & (g1909) & (g818)) + ((g832) & (!g1909) & (g818)) + ((g832) & (g1909) & (g818)));
	assign g819 = (((!g34) & (!g36) & (!reset) & (g56) & (!g818)) + ((!g34) & (!g36) & (!reset) & (g56) & (g818)) + ((!g34) & (g36) & (!reset) & (!g56) & (g818)) + ((!g34) & (g36) & (!reset) & (g56) & (g818)) + ((g34) & (!g36) & (!reset) & (g56) & (!g818)) + ((g34) & (!g36) & (!reset) & (g56) & (g818)) + ((g34) & (g36) & (!reset) & (g56) & (!g818)) + ((g34) & (g36) & (!reset) & (g56) & (g818)));
	assign g7279 = (((!g832) & (g1911) & (!g820)) + ((!g832) & (g1911) & (g820)) + ((g832) & (!g1911) & (g820)) + ((g832) & (g1911) & (g820)));
	assign g821 = (((!g34) & (!g36) & (!reset) & (g57) & (!g820)) + ((!g34) & (!g36) & (!reset) & (g57) & (g820)) + ((!g34) & (g36) & (!reset) & (!g57) & (g820)) + ((!g34) & (g36) & (!reset) & (g57) & (g820)) + ((g34) & (!g36) & (!reset) & (g57) & (!g820)) + ((g34) & (!g36) & (!reset) & (g57) & (g820)) + ((g34) & (g36) & (!reset) & (g57) & (!g820)) + ((g34) & (g36) & (!reset) & (g57) & (g820)));
	assign g7280 = (((!g832) & (g1913) & (!g822)) + ((!g832) & (g1913) & (g822)) + ((g832) & (!g1913) & (g822)) + ((g832) & (g1913) & (g822)));
	assign g823 = (((!g34) & (!g36) & (!reset) & (g58) & (!g822)) + ((!g34) & (!g36) & (!reset) & (g58) & (g822)) + ((!g34) & (g36) & (!reset) & (!g58) & (g822)) + ((!g34) & (g36) & (!reset) & (g58) & (g822)) + ((g34) & (!g36) & (!reset) & (g58) & (!g822)) + ((g34) & (!g36) & (!reset) & (g58) & (g822)) + ((g34) & (g36) & (!reset) & (g58) & (!g822)) + ((g34) & (g36) & (!reset) & (g58) & (g822)));
	assign g824 = (((!g60) & (g61)) + ((g60) & (!g61)));
	assign g825 = (((!g34) & (g35) & (g36) & (!reset) & (!g781) & (g824)) + ((!g34) & (g35) & (g36) & (!reset) & (g781) & (g824)) + ((g34) & (!g35) & (g36) & (!reset) & (!g781) & (g824)) + ((g34) & (g35) & (g36) & (!reset) & (!g781) & (g824)));
	assign g826 = (((!g34) & (!g35) & (!g36) & (!reset) & (!g61) & (!g781)) + ((!g34) & (!g35) & (!g36) & (!reset) & (!g61) & (g781)) + ((!g34) & (!g35) & (!g36) & (!reset) & (g61) & (!g781)) + ((!g34) & (!g35) & (!g36) & (!reset) & (g61) & (g781)) + ((!g34) & (!g35) & (!g36) & (reset) & (!g61) & (!g781)) + ((!g34) & (!g35) & (!g36) & (reset) & (!g61) & (g781)) + ((!g34) & (!g35) & (!g36) & (reset) & (g61) & (!g781)) + ((!g34) & (!g35) & (!g36) & (reset) & (g61) & (g781)) + ((!g34) & (!g35) & (g36) & (!reset) & (!g61) & (!g781)) + ((!g34) & (!g35) & (g36) & (!reset) & (!g61) & (g781)) + ((!g34) & (!g35) & (g36) & (!reset) & (g61) & (!g781)) + ((!g34) & (!g35) & (g36) & (!reset) & (g61) & (g781)) + ((!g34) & (!g35) & (g36) & (reset) & (!g61) & (!g781)) + ((!g34) & (!g35) & (g36) & (reset) & (!g61) & (g781)) + ((!g34) & (!g35) & (g36) & (reset) & (g61) & (!g781)) + ((!g34) & (!g35) & (g36) & (reset) & (g61) & (g781)) + ((!g34) & (g35) & (!g36) & (!reset) & (!g61) & (!g781)) + ((!g34) & (g35) & (!g36) & (!reset) & (!g61) & (g781)) + ((!g34) & (g35) & (!g36) & (!reset) & (g61) & (!g781)) + ((!g34) & (g35) & (!g36) & (!reset) & (g61) & (g781)) + ((!g34) & (g35) & (!g36) & (reset) & (!g61) & (!g781)) + ((!g34) & (g35) & (!g36) & (reset) & (!g61) & (g781)) + ((!g34) & (g35) & (!g36) & (reset) & (g61) & (!g781)) + ((!g34) & (g35) & (!g36) & (reset) & (g61) & (g781)) + ((!g34) & (g35) & (g36) & (!reset) & (g61) & (!g781)) + ((!g34) & (g35) & (g36) & (!reset) & (g61) & (g781)) + ((!g34) & (g35) & (g36) & (reset) & (!g61) & (!g781)) + ((!g34) & (g35) & (g36) & (reset) & (!g61) & (g781)) + ((!g34) & (g35) & (g36) & (reset) & (g61) & (!g781)) + ((!g34) & (g35) & (g36) & (reset) & (g61) & (g781)) + ((g34) & (!g35) & (!g36) & (!reset) & (!g61) & (!g781)) + ((g34) & (!g35) & (!g36) & (!reset) & (!g61) & (g781)) + ((g34) & (!g35) & (!g36) & (!reset) & (g61) & (!g781)) + ((g34) & (!g35) & (!g36) & (!reset) & (g61) & (g781)) + ((g34) & (!g35) & (!g36) & (reset) & (!g61) & (!g781)) + ((g34) & (!g35) & (!g36) & (reset) & (!g61) & (g781)) + ((g34) & (!g35) & (!g36) & (reset) & (g61) & (!g781)) + ((g34) & (!g35) & (!g36) & (reset) & (g61) & (g781)) + ((g34) & (!g35) & (g36) & (!reset) & (!g61) & (g781)) + ((g34) & (!g35) & (g36) & (!reset) & (g61) & (!g781)) + ((g34) & (!g35) & (g36) & (!reset) & (g61) & (g781)) + ((g34) & (!g35) & (g36) & (reset) & (!g61) & (!g781)) + ((g34) & (!g35) & (g36) & (reset) & (!g61) & (g781)) + ((g34) & (!g35) & (g36) & (reset) & (g61) & (!g781)) + ((g34) & (!g35) & (g36) & (reset) & (g61) & (g781)) + ((g34) & (g35) & (!g36) & (!reset) & (!g61) & (!g781)) + ((g34) & (g35) & (!g36) & (!reset) & (!g61) & (g781)) + ((g34) & (g35) & (!g36) & (!reset) & (g61) & (!g781)) + ((g34) & (g35) & (!g36) & (!reset) & (g61) & (g781)) + ((g34) & (g35) & (!g36) & (reset) & (!g61) & (!g781)) + ((g34) & (g35) & (!g36) & (reset) & (!g61) & (g781)) + ((g34) & (g35) & (!g36) & (reset) & (g61) & (!g781)) + ((g34) & (g35) & (!g36) & (reset) & (g61) & (g781)) + ((g34) & (g35) & (g36) & (!reset) & (!g61) & (g781)) + ((g34) & (g35) & (g36) & (!reset) & (g61) & (!g781)) + ((g34) & (g35) & (g36) & (!reset) & (g61) & (g781)) + ((g34) & (g35) & (g36) & (reset) & (!g61) & (!g781)) + ((g34) & (g35) & (g36) & (reset) & (!g61) & (g781)) + ((g34) & (g35) & (g36) & (reset) & (g61) & (!g781)) + ((g34) & (g35) & (g36) & (reset) & (g61) & (g781)));
	assign g7281 = (((!g1938) & (g1937) & (!g827)) + ((!g1938) & (g1937) & (g827)) + ((g1938) & (!g1937) & (g827)) + ((g1938) & (g1937) & (g827)));
	assign g7282 = (((!g2017) & (g7190) & (!g828)) + ((!g2017) & (g7190) & (g828)) + ((g2017) & (!g7190) & (g828)) + ((g2017) & (g7190) & (g828)));
	assign g829 = (((!g63) & (!g827) & (g828)) + ((!g63) & (g827) & (g828)) + ((g63) & (!g827) & (g828)) + ((g63) & (g827) & (!g828)));
	assign g832 = (((!reset) & (!g827) & (!g830) & (!g831)) + ((!reset) & (!g827) & (!g830) & (g831)) + ((!reset) & (!g827) & (g830) & (g831)) + ((!reset) & (g827) & (!g830) & (g831)) + ((!reset) & (g827) & (g830) & (!g831)) + ((!reset) & (g827) & (g830) & (g831)) + ((reset) & (!g827) & (!g830) & (!g831)) + ((reset) & (!g827) & (!g830) & (g831)) + ((reset) & (!g827) & (g830) & (!g831)) + ((reset) & (!g827) & (g830) & (g831)) + ((reset) & (g827) & (!g830) & (!g831)) + ((reset) & (g827) & (!g830) & (g831)) + ((reset) & (g827) & (g830) & (!g831)) + ((reset) & (g827) & (g830) & (g831)));
	assign g833 = (((!g34) & (!g36) & (!reset) & (g66) & (!g87)) + ((!g34) & (!g36) & (!reset) & (g66) & (g87)) + ((!g34) & (g36) & (!reset) & (!g66) & (g87)) + ((!g34) & (g36) & (!reset) & (g66) & (g87)) + ((g34) & (!g36) & (!reset) & (g66) & (!g87)) + ((g34) & (!g36) & (!reset) & (g66) & (g87)) + ((g34) & (g36) & (!reset) & (g66) & (!g87)) + ((g34) & (g36) & (!reset) & (g66) & (g87)));
	assign g7283 = (((!g832) & (g2021) & (!g834)) + ((!g832) & (g2021) & (g834)) + ((g832) & (!g2021) & (g834)) + ((g832) & (g2021) & (g834)));
	assign g835 = (((!g34) & (!g36) & (!reset) & (g67) & (!g834)) + ((!g34) & (!g36) & (!reset) & (g67) & (g834)) + ((!g34) & (g36) & (!reset) & (!g67) & (g834)) + ((!g34) & (g36) & (!reset) & (g67) & (g834)) + ((g34) & (!g36) & (!reset) & (g67) & (!g834)) + ((g34) & (!g36) & (!reset) & (g67) & (g834)) + ((g34) & (g36) & (!reset) & (g67) & (!g834)) + ((g34) & (g36) & (!reset) & (g67) & (g834)));
	assign g7284 = (((!g832) & (g2023) & (!g836)) + ((!g832) & (g2023) & (g836)) + ((g832) & (!g2023) & (g836)) + ((g832) & (g2023) & (g836)));
	assign g837 = (((!g34) & (!g36) & (!reset) & (g68) & (!g836)) + ((!g34) & (!g36) & (!reset) & (g68) & (g836)) + ((!g34) & (g36) & (!reset) & (!g68) & (g836)) + ((!g34) & (g36) & (!reset) & (g68) & (g836)) + ((g34) & (!g36) & (!reset) & (g68) & (!g836)) + ((g34) & (!g36) & (!reset) & (g68) & (g836)) + ((g34) & (g36) & (!reset) & (g68) & (!g836)) + ((g34) & (g36) & (!reset) & (g68) & (g836)));
	assign g7285 = (((!g832) & (g2024) & (!g838)) + ((!g832) & (g2024) & (g838)) + ((g832) & (!g2024) & (g838)) + ((g832) & (g2024) & (g838)));
	assign g839 = (((!g34) & (!g36) & (!reset) & (g69) & (!g838)) + ((!g34) & (!g36) & (!reset) & (g69) & (g838)) + ((!g34) & (g36) & (!reset) & (!g69) & (g838)) + ((!g34) & (g36) & (!reset) & (g69) & (g838)) + ((g34) & (!g36) & (!reset) & (g69) & (!g838)) + ((g34) & (!g36) & (!reset) & (g69) & (g838)) + ((g34) & (g36) & (!reset) & (g69) & (!g838)) + ((g34) & (g36) & (!reset) & (g69) & (g838)));
	assign g7286 = (((!g832) & (g2025) & (!g840)) + ((!g832) & (g2025) & (g840)) + ((g832) & (!g2025) & (g840)) + ((g832) & (g2025) & (g840)));
	assign g841 = (((!g34) & (!g36) & (!reset) & (g71) & (!g840)) + ((!g34) & (!g36) & (!reset) & (g71) & (g840)) + ((!g34) & (g36) & (!reset) & (!g71) & (g840)) + ((!g34) & (g36) & (!reset) & (g71) & (g840)) + ((g34) & (!g36) & (!reset) & (g71) & (!g840)) + ((g34) & (!g36) & (!reset) & (g71) & (g840)) + ((g34) & (g36) & (!reset) & (g71) & (!g840)) + ((g34) & (g36) & (!reset) & (g71) & (g840)));
	assign g7287 = (((!g832) & (g2027) & (!g842)) + ((!g832) & (g2027) & (g842)) + ((g832) & (!g2027) & (g842)) + ((g832) & (g2027) & (g842)));
	assign g843 = (((!g34) & (!g36) & (!reset) & (g72) & (!g842)) + ((!g34) & (!g36) & (!reset) & (g72) & (g842)) + ((!g34) & (g36) & (!reset) & (!g72) & (g842)) + ((!g34) & (g36) & (!reset) & (g72) & (g842)) + ((g34) & (!g36) & (!reset) & (g72) & (!g842)) + ((g34) & (!g36) & (!reset) & (g72) & (g842)) + ((g34) & (g36) & (!reset) & (g72) & (!g842)) + ((g34) & (g36) & (!reset) & (g72) & (g842)));
	assign g7288 = (((!g832) & (g2029) & (!g844)) + ((!g832) & (g2029) & (g844)) + ((g832) & (!g2029) & (g844)) + ((g832) & (g2029) & (g844)));
	assign g845 = (((!g34) & (!g36) & (!reset) & (g73) & (!g844)) + ((!g34) & (!g36) & (!reset) & (g73) & (g844)) + ((!g34) & (g36) & (!reset) & (!g73) & (g844)) + ((!g34) & (g36) & (!reset) & (g73) & (g844)) + ((g34) & (!g36) & (!reset) & (g73) & (!g844)) + ((g34) & (!g36) & (!reset) & (g73) & (g844)) + ((g34) & (g36) & (!reset) & (g73) & (!g844)) + ((g34) & (g36) & (!reset) & (g73) & (g844)));
	assign g7289 = (((!g832) & (g2031) & (!g846)) + ((!g832) & (g2031) & (g846)) + ((g832) & (!g2031) & (g846)) + ((g832) & (g2031) & (g846)));
	assign g847 = (((!g34) & (!g36) & (!reset) & (g74) & (!g846)) + ((!g34) & (!g36) & (!reset) & (g74) & (g846)) + ((!g34) & (g36) & (!reset) & (!g74) & (g846)) + ((!g34) & (g36) & (!reset) & (g74) & (g846)) + ((g34) & (!g36) & (!reset) & (g74) & (!g846)) + ((g34) & (!g36) & (!reset) & (g74) & (g846)) + ((g34) & (g36) & (!reset) & (g74) & (!g846)) + ((g34) & (g36) & (!reset) & (g74) & (g846)));
	assign g7290 = (((!g832) & (g2033) & (!g848)) + ((!g832) & (g2033) & (g848)) + ((g832) & (!g2033) & (g848)) + ((g832) & (g2033) & (g848)));
	assign g849 = (((!g34) & (!g36) & (!reset) & (g76) & (!g848)) + ((!g34) & (!g36) & (!reset) & (g76) & (g848)) + ((!g34) & (g36) & (!reset) & (!g76) & (g848)) + ((!g34) & (g36) & (!reset) & (g76) & (g848)) + ((g34) & (!g36) & (!reset) & (g76) & (!g848)) + ((g34) & (!g36) & (!reset) & (g76) & (g848)) + ((g34) & (g36) & (!reset) & (g76) & (!g848)) + ((g34) & (g36) & (!reset) & (g76) & (g848)));
	assign g7291 = (((!g832) & (g2035) & (!g850)) + ((!g832) & (g2035) & (g850)) + ((g832) & (!g2035) & (g850)) + ((g832) & (g2035) & (g850)));
	assign g851 = (((!g34) & (!g36) & (!reset) & (g77) & (!g850)) + ((!g34) & (!g36) & (!reset) & (g77) & (g850)) + ((!g34) & (g36) & (!reset) & (!g77) & (g850)) + ((!g34) & (g36) & (!reset) & (g77) & (g850)) + ((g34) & (!g36) & (!reset) & (g77) & (!g850)) + ((g34) & (!g36) & (!reset) & (g77) & (g850)) + ((g34) & (g36) & (!reset) & (g77) & (!g850)) + ((g34) & (g36) & (!reset) & (g77) & (g850)));
	assign g7292 = (((!g832) & (g2037) & (!g852)) + ((!g832) & (g2037) & (g852)) + ((g832) & (!g2037) & (g852)) + ((g832) & (g2037) & (g852)));
	assign g853 = (((!g34) & (!g36) & (!reset) & (g78) & (!g852)) + ((!g34) & (!g36) & (!reset) & (g78) & (g852)) + ((!g34) & (g36) & (!reset) & (!g78) & (g852)) + ((!g34) & (g36) & (!reset) & (g78) & (g852)) + ((g34) & (!g36) & (!reset) & (g78) & (!g852)) + ((g34) & (!g36) & (!reset) & (g78) & (g852)) + ((g34) & (g36) & (!reset) & (g78) & (!g852)) + ((g34) & (g36) & (!reset) & (g78) & (g852)));
	assign g7293 = (((!g832) & (g2039) & (!g854)) + ((!g832) & (g2039) & (g854)) + ((g832) & (!g2039) & (g854)) + ((g832) & (g2039) & (g854)));
	assign g855 = (((!g34) & (!g36) & (!reset) & (g79) & (!g854)) + ((!g34) & (!g36) & (!reset) & (g79) & (g854)) + ((!g34) & (g36) & (!reset) & (!g79) & (g854)) + ((!g34) & (g36) & (!reset) & (g79) & (g854)) + ((g34) & (!g36) & (!reset) & (g79) & (!g854)) + ((g34) & (!g36) & (!reset) & (g79) & (g854)) + ((g34) & (g36) & (!reset) & (g79) & (!g854)) + ((g34) & (g36) & (!reset) & (g79) & (g854)));
	assign g7294 = (((!g832) & (g2040) & (!g856)) + ((!g832) & (g2040) & (g856)) + ((g832) & (!g2040) & (g856)) + ((g832) & (g2040) & (g856)));
	assign g857 = (((!g34) & (!g36) & (!reset) & (g81) & (!g856)) + ((!g34) & (!g36) & (!reset) & (g81) & (g856)) + ((!g34) & (g36) & (!reset) & (!g81) & (g856)) + ((!g34) & (g36) & (!reset) & (g81) & (g856)) + ((g34) & (!g36) & (!reset) & (g81) & (!g856)) + ((g34) & (!g36) & (!reset) & (g81) & (g856)) + ((g34) & (g36) & (!reset) & (g81) & (!g856)) + ((g34) & (g36) & (!reset) & (g81) & (g856)));
	assign g7295 = (((!g832) & (g2042) & (!g858)) + ((!g832) & (g2042) & (g858)) + ((g832) & (!g2042) & (g858)) + ((g832) & (g2042) & (g858)));
	assign g859 = (((!g34) & (!g36) & (!reset) & (g82) & (!g858)) + ((!g34) & (!g36) & (!reset) & (g82) & (g858)) + ((!g34) & (g36) & (!reset) & (!g82) & (g858)) + ((!g34) & (g36) & (!reset) & (g82) & (g858)) + ((g34) & (!g36) & (!reset) & (g82) & (!g858)) + ((g34) & (!g36) & (!reset) & (g82) & (g858)) + ((g34) & (g36) & (!reset) & (g82) & (!g858)) + ((g34) & (g36) & (!reset) & (g82) & (g858)));
	assign g7296 = (((!g832) & (g2044) & (!g860)) + ((!g832) & (g2044) & (g860)) + ((g832) & (!g2044) & (g860)) + ((g832) & (g2044) & (g860)));
	assign g861 = (((!g34) & (!g36) & (!reset) & (g83) & (!g860)) + ((!g34) & (!g36) & (!reset) & (g83) & (g860)) + ((!g34) & (g36) & (!reset) & (!g83) & (g860)) + ((!g34) & (g36) & (!reset) & (g83) & (g860)) + ((g34) & (!g36) & (!reset) & (g83) & (!g860)) + ((g34) & (!g36) & (!reset) & (g83) & (g860)) + ((g34) & (g36) & (!reset) & (g83) & (!g860)) + ((g34) & (g36) & (!reset) & (g83) & (g860)));
	assign g7297 = (((!g832) & (g2046) & (!g862)) + ((!g832) & (g2046) & (g862)) + ((g832) & (!g2046) & (g862)) + ((g832) & (g2046) & (g862)));
	assign g863 = (((!g34) & (!g36) & (!reset) & (g84) & (!g862)) + ((!g34) & (!g36) & (!reset) & (g84) & (g862)) + ((!g34) & (g36) & (!reset) & (!g84) & (g862)) + ((!g34) & (g36) & (!reset) & (g84) & (g862)) + ((g34) & (!g36) & (!reset) & (g84) & (!g862)) + ((g34) & (!g36) & (!reset) & (g84) & (g862)) + ((g34) & (g36) & (!reset) & (g84) & (!g862)) + ((g34) & (g36) & (!reset) & (g84) & (g862)));
	assign g7298 = (((!g2017) & (g7184) & (!g864)) + ((!g2017) & (g7184) & (g864)) + ((g2017) & (!g7184) & (g864)) + ((g2017) & (g7184) & (g864)));
	assign g865 = (((!g63) & (!g827) & (!g87) & (!g828) & (g864)) + ((!g63) & (!g827) & (!g87) & (g828) & (g864)) + ((!g63) & (!g827) & (g87) & (!g828) & (g864)) + ((!g63) & (!g827) & (g87) & (g828) & (g864)) + ((!g63) & (g827) & (!g87) & (!g828) & (g864)) + ((!g63) & (g827) & (!g87) & (g828) & (g864)) + ((!g63) & (g827) & (g87) & (!g828) & (!g864)) + ((!g63) & (g827) & (g87) & (g828) & (!g864)) + ((g63) & (!g827) & (!g87) & (!g828) & (g864)) + ((g63) & (!g827) & (!g87) & (g828) & (g864)) + ((g63) & (!g827) & (g87) & (!g828) & (g864)) + ((g63) & (!g827) & (g87) & (g828) & (g864)) + ((g63) & (g827) & (!g87) & (!g828) & (g864)) + ((g63) & (g827) & (!g87) & (g828) & (!g864)) + ((g63) & (g827) & (g87) & (!g828) & (!g864)) + ((g63) & (g827) & (g87) & (g828) & (g864)));
	assign g866 = (((!g34) & (!g36) & (!reset) & (g89) & (!g110)) + ((!g34) & (!g36) & (!reset) & (g89) & (g110)) + ((!g34) & (g36) & (!reset) & (!g89) & (g110)) + ((!g34) & (g36) & (!reset) & (g89) & (g110)) + ((g34) & (!g36) & (!reset) & (g89) & (!g110)) + ((g34) & (!g36) & (!reset) & (g89) & (g110)) + ((g34) & (g36) & (!reset) & (g89) & (!g110)) + ((g34) & (g36) & (!reset) & (g89) & (g110)));
	assign g7299 = (((!g832) & (g2054) & (!g867)) + ((!g832) & (g2054) & (g867)) + ((g832) & (!g2054) & (g867)) + ((g832) & (g2054) & (g867)));
	assign g868 = (((!g34) & (!g36) & (!reset) & (g90) & (!g867)) + ((!g34) & (!g36) & (!reset) & (g90) & (g867)) + ((!g34) & (g36) & (!reset) & (!g90) & (g867)) + ((!g34) & (g36) & (!reset) & (g90) & (g867)) + ((g34) & (!g36) & (!reset) & (g90) & (!g867)) + ((g34) & (!g36) & (!reset) & (g90) & (g867)) + ((g34) & (g36) & (!reset) & (g90) & (!g867)) + ((g34) & (g36) & (!reset) & (g90) & (g867)));
	assign g7300 = (((!g832) & (g2057) & (!g869)) + ((!g832) & (g2057) & (g869)) + ((g832) & (!g2057) & (g869)) + ((g832) & (g2057) & (g869)));
	assign g870 = (((!g34) & (!g36) & (!reset) & (g91) & (!g869)) + ((!g34) & (!g36) & (!reset) & (g91) & (g869)) + ((!g34) & (g36) & (!reset) & (!g91) & (g869)) + ((!g34) & (g36) & (!reset) & (g91) & (g869)) + ((g34) & (!g36) & (!reset) & (g91) & (!g869)) + ((g34) & (!g36) & (!reset) & (g91) & (g869)) + ((g34) & (g36) & (!reset) & (g91) & (!g869)) + ((g34) & (g36) & (!reset) & (g91) & (g869)));
	assign g7301 = (((!g832) & (g2059) & (!g871)) + ((!g832) & (g2059) & (g871)) + ((g832) & (!g2059) & (g871)) + ((g832) & (g2059) & (g871)));
	assign g872 = (((!g34) & (!g36) & (!reset) & (g92) & (!g871)) + ((!g34) & (!g36) & (!reset) & (g92) & (g871)) + ((!g34) & (g36) & (!reset) & (!g92) & (g871)) + ((!g34) & (g36) & (!reset) & (g92) & (g871)) + ((g34) & (!g36) & (!reset) & (g92) & (!g871)) + ((g34) & (!g36) & (!reset) & (g92) & (g871)) + ((g34) & (g36) & (!reset) & (g92) & (!g871)) + ((g34) & (g36) & (!reset) & (g92) & (g871)));
	assign g7302 = (((!g832) & (g2061) & (!g873)) + ((!g832) & (g2061) & (g873)) + ((g832) & (!g2061) & (g873)) + ((g832) & (g2061) & (g873)));
	assign g874 = (((!g34) & (!g36) & (!reset) & (g94) & (!g873)) + ((!g34) & (!g36) & (!reset) & (g94) & (g873)) + ((!g34) & (g36) & (!reset) & (!g94) & (g873)) + ((!g34) & (g36) & (!reset) & (g94) & (g873)) + ((g34) & (!g36) & (!reset) & (g94) & (!g873)) + ((g34) & (!g36) & (!reset) & (g94) & (g873)) + ((g34) & (g36) & (!reset) & (g94) & (!g873)) + ((g34) & (g36) & (!reset) & (g94) & (g873)));
	assign g7303 = (((!g832) & (g2064) & (!g875)) + ((!g832) & (g2064) & (g875)) + ((g832) & (!g2064) & (g875)) + ((g832) & (g2064) & (g875)));
	assign g876 = (((!g34) & (!g36) & (!reset) & (g95) & (!g875)) + ((!g34) & (!g36) & (!reset) & (g95) & (g875)) + ((!g34) & (g36) & (!reset) & (!g95) & (g875)) + ((!g34) & (g36) & (!reset) & (g95) & (g875)) + ((g34) & (!g36) & (!reset) & (g95) & (!g875)) + ((g34) & (!g36) & (!reset) & (g95) & (g875)) + ((g34) & (g36) & (!reset) & (g95) & (!g875)) + ((g34) & (g36) & (!reset) & (g95) & (g875)));
	assign g7304 = (((!g832) & (g2067) & (!g877)) + ((!g832) & (g2067) & (g877)) + ((g832) & (!g2067) & (g877)) + ((g832) & (g2067) & (g877)));
	assign g878 = (((!g34) & (!g36) & (!reset) & (g96) & (!g877)) + ((!g34) & (!g36) & (!reset) & (g96) & (g877)) + ((!g34) & (g36) & (!reset) & (!g96) & (g877)) + ((!g34) & (g36) & (!reset) & (g96) & (g877)) + ((g34) & (!g36) & (!reset) & (g96) & (!g877)) + ((g34) & (!g36) & (!reset) & (g96) & (g877)) + ((g34) & (g36) & (!reset) & (g96) & (!g877)) + ((g34) & (g36) & (!reset) & (g96) & (g877)));
	assign g7305 = (((!g832) & (g2070) & (!g879)) + ((!g832) & (g2070) & (g879)) + ((g832) & (!g2070) & (g879)) + ((g832) & (g2070) & (g879)));
	assign g880 = (((!g34) & (!g36) & (!reset) & (g97) & (!g879)) + ((!g34) & (!g36) & (!reset) & (g97) & (g879)) + ((!g34) & (g36) & (!reset) & (!g97) & (g879)) + ((!g34) & (g36) & (!reset) & (g97) & (g879)) + ((g34) & (!g36) & (!reset) & (g97) & (!g879)) + ((g34) & (!g36) & (!reset) & (g97) & (g879)) + ((g34) & (g36) & (!reset) & (g97) & (!g879)) + ((g34) & (g36) & (!reset) & (g97) & (g879)));
	assign g7306 = (((!g832) & (g2073) & (!g881)) + ((!g832) & (g2073) & (g881)) + ((g832) & (!g2073) & (g881)) + ((g832) & (g2073) & (g881)));
	assign g882 = (((!g34) & (!g36) & (!reset) & (g99) & (!g881)) + ((!g34) & (!g36) & (!reset) & (g99) & (g881)) + ((!g34) & (g36) & (!reset) & (!g99) & (g881)) + ((!g34) & (g36) & (!reset) & (g99) & (g881)) + ((g34) & (!g36) & (!reset) & (g99) & (!g881)) + ((g34) & (!g36) & (!reset) & (g99) & (g881)) + ((g34) & (g36) & (!reset) & (g99) & (!g881)) + ((g34) & (g36) & (!reset) & (g99) & (g881)));
	assign g7307 = (((!g832) & (g2076) & (!g883)) + ((!g832) & (g2076) & (g883)) + ((g832) & (!g2076) & (g883)) + ((g832) & (g2076) & (g883)));
	assign g884 = (((!g34) & (!g36) & (!reset) & (g100) & (!g883)) + ((!g34) & (!g36) & (!reset) & (g100) & (g883)) + ((!g34) & (g36) & (!reset) & (!g100) & (g883)) + ((!g34) & (g36) & (!reset) & (g100) & (g883)) + ((g34) & (!g36) & (!reset) & (g100) & (!g883)) + ((g34) & (!g36) & (!reset) & (g100) & (g883)) + ((g34) & (g36) & (!reset) & (g100) & (!g883)) + ((g34) & (g36) & (!reset) & (g100) & (g883)));
	assign g7308 = (((!g832) & (g2079) & (!g885)) + ((!g832) & (g2079) & (g885)) + ((g832) & (!g2079) & (g885)) + ((g832) & (g2079) & (g885)));
	assign g886 = (((!g34) & (!g36) & (!reset) & (g101) & (!g885)) + ((!g34) & (!g36) & (!reset) & (g101) & (g885)) + ((!g34) & (g36) & (!reset) & (!g101) & (g885)) + ((!g34) & (g36) & (!reset) & (g101) & (g885)) + ((g34) & (!g36) & (!reset) & (g101) & (!g885)) + ((g34) & (!g36) & (!reset) & (g101) & (g885)) + ((g34) & (g36) & (!reset) & (g101) & (!g885)) + ((g34) & (g36) & (!reset) & (g101) & (g885)));
	assign g7309 = (((!g832) & (g2082) & (!g887)) + ((!g832) & (g2082) & (g887)) + ((g832) & (!g2082) & (g887)) + ((g832) & (g2082) & (g887)));
	assign g888 = (((!g34) & (!g36) & (!reset) & (g102) & (!g887)) + ((!g34) & (!g36) & (!reset) & (g102) & (g887)) + ((!g34) & (g36) & (!reset) & (!g102) & (g887)) + ((!g34) & (g36) & (!reset) & (g102) & (g887)) + ((g34) & (!g36) & (!reset) & (g102) & (!g887)) + ((g34) & (!g36) & (!reset) & (g102) & (g887)) + ((g34) & (g36) & (!reset) & (g102) & (!g887)) + ((g34) & (g36) & (!reset) & (g102) & (g887)));
	assign g7310 = (((!g832) & (g2084) & (!g889)) + ((!g832) & (g2084) & (g889)) + ((g832) & (!g2084) & (g889)) + ((g832) & (g2084) & (g889)));
	assign g890 = (((!g34) & (!g36) & (!reset) & (g104) & (!g889)) + ((!g34) & (!g36) & (!reset) & (g104) & (g889)) + ((!g34) & (g36) & (!reset) & (!g104) & (g889)) + ((!g34) & (g36) & (!reset) & (g104) & (g889)) + ((g34) & (!g36) & (!reset) & (g104) & (!g889)) + ((g34) & (!g36) & (!reset) & (g104) & (g889)) + ((g34) & (g36) & (!reset) & (g104) & (!g889)) + ((g34) & (g36) & (!reset) & (g104) & (g889)));
	assign g7311 = (((!g832) & (g2087) & (!g891)) + ((!g832) & (g2087) & (g891)) + ((g832) & (!g2087) & (g891)) + ((g832) & (g2087) & (g891)));
	assign g892 = (((!g34) & (!g36) & (!reset) & (g105) & (!g891)) + ((!g34) & (!g36) & (!reset) & (g105) & (g891)) + ((!g34) & (g36) & (!reset) & (!g105) & (g891)) + ((!g34) & (g36) & (!reset) & (g105) & (g891)) + ((g34) & (!g36) & (!reset) & (g105) & (!g891)) + ((g34) & (!g36) & (!reset) & (g105) & (g891)) + ((g34) & (g36) & (!reset) & (g105) & (!g891)) + ((g34) & (g36) & (!reset) & (g105) & (g891)));
	assign g7312 = (((!g832) & (g2090) & (!g893)) + ((!g832) & (g2090) & (g893)) + ((g832) & (!g2090) & (g893)) + ((g832) & (g2090) & (g893)));
	assign g894 = (((!g34) & (!g36) & (!reset) & (g106) & (!g893)) + ((!g34) & (!g36) & (!reset) & (g106) & (g893)) + ((!g34) & (g36) & (!reset) & (!g106) & (g893)) + ((!g34) & (g36) & (!reset) & (g106) & (g893)) + ((g34) & (!g36) & (!reset) & (g106) & (!g893)) + ((g34) & (!g36) & (!reset) & (g106) & (g893)) + ((g34) & (g36) & (!reset) & (g106) & (!g893)) + ((g34) & (g36) & (!reset) & (g106) & (g893)));
	assign g7313 = (((!g832) & (g2093) & (!g895)) + ((!g832) & (g2093) & (g895)) + ((g832) & (!g2093) & (g895)) + ((g832) & (g2093) & (g895)));
	assign g896 = (((!g34) & (!g36) & (!reset) & (g107) & (!g895)) + ((!g34) & (!g36) & (!reset) & (g107) & (g895)) + ((!g34) & (g36) & (!reset) & (!g107) & (g895)) + ((!g34) & (g36) & (!reset) & (g107) & (g895)) + ((g34) & (!g36) & (!reset) & (g107) & (!g895)) + ((g34) & (!g36) & (!reset) & (g107) & (g895)) + ((g34) & (g36) & (!reset) & (g107) & (!g895)) + ((g34) & (g36) & (!reset) & (g107) & (g895)));
	assign g7314 = (((!g2017) & (g7177) & (!g897)) + ((!g2017) & (g7177) & (g897)) + ((g2017) & (!g7177) & (g897)) + ((g2017) & (g7177) & (g897)));
	assign g898 = (((!g63) & (g87) & (!g828) & (g864)) + ((!g63) & (g87) & (g828) & (g864)) + ((g63) & (!g87) & (g828) & (g864)) + ((g63) & (g87) & (!g828) & (g864)) + ((g63) & (g87) & (g828) & (!g864)) + ((g63) & (g87) & (g828) & (g864)));
	assign g899 = (((!g827) & (!g110) & (g897) & (!g898)) + ((!g827) & (!g110) & (g897) & (g898)) + ((!g827) & (g110) & (g897) & (!g898)) + ((!g827) & (g110) & (g897) & (g898)) + ((g827) & (!g110) & (!g897) & (g898)) + ((g827) & (!g110) & (g897) & (!g898)) + ((g827) & (g110) & (!g897) & (!g898)) + ((g827) & (g110) & (g897) & (g898)));
	assign g900 = (((!g34) & (!g36) & (!reset) & (g112) & (!g133)) + ((!g34) & (!g36) & (!reset) & (g112) & (g133)) + ((!g34) & (g36) & (!reset) & (!g112) & (g133)) + ((!g34) & (g36) & (!reset) & (g112) & (g133)) + ((g34) & (!g36) & (!reset) & (g112) & (!g133)) + ((g34) & (!g36) & (!reset) & (g112) & (g133)) + ((g34) & (g36) & (!reset) & (g112) & (!g133)) + ((g34) & (g36) & (!reset) & (g112) & (g133)));
	assign g7315 = (((!g832) & (g2103) & (!g901)) + ((!g832) & (g2103) & (g901)) + ((g832) & (!g2103) & (g901)) + ((g832) & (g2103) & (g901)));
	assign g902 = (((!g34) & (!g36) & (!reset) & (g113) & (!g901)) + ((!g34) & (!g36) & (!reset) & (g113) & (g901)) + ((!g34) & (g36) & (!reset) & (!g113) & (g901)) + ((!g34) & (g36) & (!reset) & (g113) & (g901)) + ((g34) & (!g36) & (!reset) & (g113) & (!g901)) + ((g34) & (!g36) & (!reset) & (g113) & (g901)) + ((g34) & (g36) & (!reset) & (g113) & (!g901)) + ((g34) & (g36) & (!reset) & (g113) & (g901)));
	assign g7316 = (((!g832) & (g2105) & (!g903)) + ((!g832) & (g2105) & (g903)) + ((g832) & (!g2105) & (g903)) + ((g832) & (g2105) & (g903)));
	assign g904 = (((!g34) & (!g36) & (!reset) & (g114) & (!g903)) + ((!g34) & (!g36) & (!reset) & (g114) & (g903)) + ((!g34) & (g36) & (!reset) & (!g114) & (g903)) + ((!g34) & (g36) & (!reset) & (g114) & (g903)) + ((g34) & (!g36) & (!reset) & (g114) & (!g903)) + ((g34) & (!g36) & (!reset) & (g114) & (g903)) + ((g34) & (g36) & (!reset) & (g114) & (!g903)) + ((g34) & (g36) & (!reset) & (g114) & (g903)));
	assign g7317 = (((!g832) & (g2106) & (!g905)) + ((!g832) & (g2106) & (g905)) + ((g832) & (!g2106) & (g905)) + ((g832) & (g2106) & (g905)));
	assign g906 = (((!g34) & (!g36) & (!reset) & (g115) & (!g905)) + ((!g34) & (!g36) & (!reset) & (g115) & (g905)) + ((!g34) & (g36) & (!reset) & (!g115) & (g905)) + ((!g34) & (g36) & (!reset) & (g115) & (g905)) + ((g34) & (!g36) & (!reset) & (g115) & (!g905)) + ((g34) & (!g36) & (!reset) & (g115) & (g905)) + ((g34) & (g36) & (!reset) & (g115) & (!g905)) + ((g34) & (g36) & (!reset) & (g115) & (g905)));
	assign g7318 = (((!g832) & (g2107) & (!g907)) + ((!g832) & (g2107) & (g907)) + ((g832) & (!g2107) & (g907)) + ((g832) & (g2107) & (g907)));
	assign g908 = (((!g34) & (!g36) & (!reset) & (g117) & (!g907)) + ((!g34) & (!g36) & (!reset) & (g117) & (g907)) + ((!g34) & (g36) & (!reset) & (!g117) & (g907)) + ((!g34) & (g36) & (!reset) & (g117) & (g907)) + ((g34) & (!g36) & (!reset) & (g117) & (!g907)) + ((g34) & (!g36) & (!reset) & (g117) & (g907)) + ((g34) & (g36) & (!reset) & (g117) & (!g907)) + ((g34) & (g36) & (!reset) & (g117) & (g907)));
	assign g7319 = (((!g832) & (g2109) & (!g909)) + ((!g832) & (g2109) & (g909)) + ((g832) & (!g2109) & (g909)) + ((g832) & (g2109) & (g909)));
	assign g910 = (((!g34) & (!g36) & (!reset) & (g118) & (!g909)) + ((!g34) & (!g36) & (!reset) & (g118) & (g909)) + ((!g34) & (g36) & (!reset) & (!g118) & (g909)) + ((!g34) & (g36) & (!reset) & (g118) & (g909)) + ((g34) & (!g36) & (!reset) & (g118) & (!g909)) + ((g34) & (!g36) & (!reset) & (g118) & (g909)) + ((g34) & (g36) & (!reset) & (g118) & (!g909)) + ((g34) & (g36) & (!reset) & (g118) & (g909)));
	assign g7320 = (((!g832) & (g2111) & (!g911)) + ((!g832) & (g2111) & (g911)) + ((g832) & (!g2111) & (g911)) + ((g832) & (g2111) & (g911)));
	assign g912 = (((!g34) & (!g36) & (!reset) & (g119) & (!g911)) + ((!g34) & (!g36) & (!reset) & (g119) & (g911)) + ((!g34) & (g36) & (!reset) & (!g119) & (g911)) + ((!g34) & (g36) & (!reset) & (g119) & (g911)) + ((g34) & (!g36) & (!reset) & (g119) & (!g911)) + ((g34) & (!g36) & (!reset) & (g119) & (g911)) + ((g34) & (g36) & (!reset) & (g119) & (!g911)) + ((g34) & (g36) & (!reset) & (g119) & (g911)));
	assign g7321 = (((!g832) & (g2113) & (!g913)) + ((!g832) & (g2113) & (g913)) + ((g832) & (!g2113) & (g913)) + ((g832) & (g2113) & (g913)));
	assign g914 = (((!g34) & (!g36) & (!reset) & (g120) & (!g913)) + ((!g34) & (!g36) & (!reset) & (g120) & (g913)) + ((!g34) & (g36) & (!reset) & (!g120) & (g913)) + ((!g34) & (g36) & (!reset) & (g120) & (g913)) + ((g34) & (!g36) & (!reset) & (g120) & (!g913)) + ((g34) & (!g36) & (!reset) & (g120) & (g913)) + ((g34) & (g36) & (!reset) & (g120) & (!g913)) + ((g34) & (g36) & (!reset) & (g120) & (g913)));
	assign g7322 = (((!g832) & (g2115) & (!g915)) + ((!g832) & (g2115) & (g915)) + ((g832) & (!g2115) & (g915)) + ((g832) & (g2115) & (g915)));
	assign g916 = (((!g34) & (!g36) & (!reset) & (g122) & (!g915)) + ((!g34) & (!g36) & (!reset) & (g122) & (g915)) + ((!g34) & (g36) & (!reset) & (!g122) & (g915)) + ((!g34) & (g36) & (!reset) & (g122) & (g915)) + ((g34) & (!g36) & (!reset) & (g122) & (!g915)) + ((g34) & (!g36) & (!reset) & (g122) & (g915)) + ((g34) & (g36) & (!reset) & (g122) & (!g915)) + ((g34) & (g36) & (!reset) & (g122) & (g915)));
	assign g7323 = (((!g832) & (g2117) & (!g917)) + ((!g832) & (g2117) & (g917)) + ((g832) & (!g2117) & (g917)) + ((g832) & (g2117) & (g917)));
	assign g918 = (((!g34) & (!g36) & (!reset) & (g123) & (!g917)) + ((!g34) & (!g36) & (!reset) & (g123) & (g917)) + ((!g34) & (g36) & (!reset) & (!g123) & (g917)) + ((!g34) & (g36) & (!reset) & (g123) & (g917)) + ((g34) & (!g36) & (!reset) & (g123) & (!g917)) + ((g34) & (!g36) & (!reset) & (g123) & (g917)) + ((g34) & (g36) & (!reset) & (g123) & (!g917)) + ((g34) & (g36) & (!reset) & (g123) & (g917)));
	assign g7324 = (((!g832) & (g2119) & (!g919)) + ((!g832) & (g2119) & (g919)) + ((g832) & (!g2119) & (g919)) + ((g832) & (g2119) & (g919)));
	assign g920 = (((!g34) & (!g36) & (!reset) & (g124) & (!g919)) + ((!g34) & (!g36) & (!reset) & (g124) & (g919)) + ((!g34) & (g36) & (!reset) & (!g124) & (g919)) + ((!g34) & (g36) & (!reset) & (g124) & (g919)) + ((g34) & (!g36) & (!reset) & (g124) & (!g919)) + ((g34) & (!g36) & (!reset) & (g124) & (g919)) + ((g34) & (g36) & (!reset) & (g124) & (!g919)) + ((g34) & (g36) & (!reset) & (g124) & (g919)));
	assign g7325 = (((!g832) & (g2121) & (!g921)) + ((!g832) & (g2121) & (g921)) + ((g832) & (!g2121) & (g921)) + ((g832) & (g2121) & (g921)));
	assign g922 = (((!g34) & (!g36) & (!reset) & (g125) & (!g921)) + ((!g34) & (!g36) & (!reset) & (g125) & (g921)) + ((!g34) & (g36) & (!reset) & (!g125) & (g921)) + ((!g34) & (g36) & (!reset) & (g125) & (g921)) + ((g34) & (!g36) & (!reset) & (g125) & (!g921)) + ((g34) & (!g36) & (!reset) & (g125) & (g921)) + ((g34) & (g36) & (!reset) & (g125) & (!g921)) + ((g34) & (g36) & (!reset) & (g125) & (g921)));
	assign g7326 = (((!g832) & (g2122) & (!g923)) + ((!g832) & (g2122) & (g923)) + ((g832) & (!g2122) & (g923)) + ((g832) & (g2122) & (g923)));
	assign g924 = (((!g34) & (!g36) & (!reset) & (g127) & (!g923)) + ((!g34) & (!g36) & (!reset) & (g127) & (g923)) + ((!g34) & (g36) & (!reset) & (!g127) & (g923)) + ((!g34) & (g36) & (!reset) & (g127) & (g923)) + ((g34) & (!g36) & (!reset) & (g127) & (!g923)) + ((g34) & (!g36) & (!reset) & (g127) & (g923)) + ((g34) & (g36) & (!reset) & (g127) & (!g923)) + ((g34) & (g36) & (!reset) & (g127) & (g923)));
	assign g7327 = (((!g832) & (g2124) & (!g925)) + ((!g832) & (g2124) & (g925)) + ((g832) & (!g2124) & (g925)) + ((g832) & (g2124) & (g925)));
	assign g926 = (((!g34) & (!g36) & (!reset) & (g128) & (!g925)) + ((!g34) & (!g36) & (!reset) & (g128) & (g925)) + ((!g34) & (g36) & (!reset) & (!g128) & (g925)) + ((!g34) & (g36) & (!reset) & (g128) & (g925)) + ((g34) & (!g36) & (!reset) & (g128) & (!g925)) + ((g34) & (!g36) & (!reset) & (g128) & (g925)) + ((g34) & (g36) & (!reset) & (g128) & (!g925)) + ((g34) & (g36) & (!reset) & (g128) & (g925)));
	assign g7328 = (((!g832) & (g2126) & (!g927)) + ((!g832) & (g2126) & (g927)) + ((g832) & (!g2126) & (g927)) + ((g832) & (g2126) & (g927)));
	assign g928 = (((!g34) & (!g36) & (!reset) & (g129) & (!g927)) + ((!g34) & (!g36) & (!reset) & (g129) & (g927)) + ((!g34) & (g36) & (!reset) & (!g129) & (g927)) + ((!g34) & (g36) & (!reset) & (g129) & (g927)) + ((g34) & (!g36) & (!reset) & (g129) & (!g927)) + ((g34) & (!g36) & (!reset) & (g129) & (g927)) + ((g34) & (g36) & (!reset) & (g129) & (!g927)) + ((g34) & (g36) & (!reset) & (g129) & (g927)));
	assign g7329 = (((!g832) & (g2128) & (!g929)) + ((!g832) & (g2128) & (g929)) + ((g832) & (!g2128) & (g929)) + ((g832) & (g2128) & (g929)));
	assign g930 = (((!g34) & (!g36) & (!reset) & (g130) & (!g929)) + ((!g34) & (!g36) & (!reset) & (g130) & (g929)) + ((!g34) & (g36) & (!reset) & (!g130) & (g929)) + ((!g34) & (g36) & (!reset) & (g130) & (g929)) + ((g34) & (!g36) & (!reset) & (g130) & (!g929)) + ((g34) & (!g36) & (!reset) & (g130) & (g929)) + ((g34) & (g36) & (!reset) & (g130) & (!g929)) + ((g34) & (g36) & (!reset) & (g130) & (g929)));
	assign g7330 = (((!g2017) & (g7171) & (!g931)) + ((!g2017) & (g7171) & (g931)) + ((g2017) & (!g7171) & (g931)) + ((g2017) & (g7171) & (g931)));
	assign g932 = (((!g827) & (!g110) & (!g133) & (!g897) & (g931) & (!g898)) + ((!g827) & (!g110) & (!g133) & (!g897) & (g931) & (g898)) + ((!g827) & (!g110) & (!g133) & (g897) & (g931) & (!g898)) + ((!g827) & (!g110) & (!g133) & (g897) & (g931) & (g898)) + ((!g827) & (!g110) & (g133) & (!g897) & (g931) & (!g898)) + ((!g827) & (!g110) & (g133) & (!g897) & (g931) & (g898)) + ((!g827) & (!g110) & (g133) & (g897) & (g931) & (!g898)) + ((!g827) & (!g110) & (g133) & (g897) & (g931) & (g898)) + ((!g827) & (g110) & (!g133) & (!g897) & (g931) & (!g898)) + ((!g827) & (g110) & (!g133) & (!g897) & (g931) & (g898)) + ((!g827) & (g110) & (!g133) & (g897) & (g931) & (!g898)) + ((!g827) & (g110) & (!g133) & (g897) & (g931) & (g898)) + ((!g827) & (g110) & (g133) & (!g897) & (g931) & (!g898)) + ((!g827) & (g110) & (g133) & (!g897) & (g931) & (g898)) + ((!g827) & (g110) & (g133) & (g897) & (g931) & (!g898)) + ((!g827) & (g110) & (g133) & (g897) & (g931) & (g898)) + ((g827) & (!g110) & (!g133) & (!g897) & (g931) & (!g898)) + ((g827) & (!g110) & (!g133) & (!g897) & (g931) & (g898)) + ((g827) & (!g110) & (!g133) & (g897) & (!g931) & (g898)) + ((g827) & (!g110) & (!g133) & (g897) & (g931) & (!g898)) + ((g827) & (!g110) & (g133) & (!g897) & (!g931) & (!g898)) + ((g827) & (!g110) & (g133) & (!g897) & (!g931) & (g898)) + ((g827) & (!g110) & (g133) & (g897) & (!g931) & (!g898)) + ((g827) & (!g110) & (g133) & (g897) & (g931) & (g898)) + ((g827) & (g110) & (!g133) & (!g897) & (!g931) & (g898)) + ((g827) & (g110) & (!g133) & (!g897) & (g931) & (!g898)) + ((g827) & (g110) & (!g133) & (g897) & (!g931) & (!g898)) + ((g827) & (g110) & (!g133) & (g897) & (!g931) & (g898)) + ((g827) & (g110) & (g133) & (!g897) & (!g931) & (!g898)) + ((g827) & (g110) & (g133) & (!g897) & (g931) & (g898)) + ((g827) & (g110) & (g133) & (g897) & (g931) & (!g898)) + ((g827) & (g110) & (g133) & (g897) & (g931) & (g898)));
	assign g933 = (((!g34) & (!g36) & (!reset) & (g135) & (!g156)) + ((!g34) & (!g36) & (!reset) & (g135) & (g156)) + ((!g34) & (g36) & (!reset) & (!g135) & (g156)) + ((!g34) & (g36) & (!reset) & (g135) & (g156)) + ((g34) & (!g36) & (!reset) & (g135) & (!g156)) + ((g34) & (!g36) & (!reset) & (g135) & (g156)) + ((g34) & (g36) & (!reset) & (g135) & (!g156)) + ((g34) & (g36) & (!reset) & (g135) & (g156)));
	assign g7331 = (((!g832) & (g2136) & (!g934)) + ((!g832) & (g2136) & (g934)) + ((g832) & (!g2136) & (g934)) + ((g832) & (g2136) & (g934)));
	assign g935 = (((!g34) & (!g36) & (!reset) & (g136) & (!g934)) + ((!g34) & (!g36) & (!reset) & (g136) & (g934)) + ((!g34) & (g36) & (!reset) & (!g136) & (g934)) + ((!g34) & (g36) & (!reset) & (g136) & (g934)) + ((g34) & (!g36) & (!reset) & (g136) & (!g934)) + ((g34) & (!g36) & (!reset) & (g136) & (g934)) + ((g34) & (g36) & (!reset) & (g136) & (!g934)) + ((g34) & (g36) & (!reset) & (g136) & (g934)));
	assign g7332 = (((!g832) & (g2139) & (!g936)) + ((!g832) & (g2139) & (g936)) + ((g832) & (!g2139) & (g936)) + ((g832) & (g2139) & (g936)));
	assign g937 = (((!g34) & (!g36) & (!reset) & (g137) & (!g936)) + ((!g34) & (!g36) & (!reset) & (g137) & (g936)) + ((!g34) & (g36) & (!reset) & (!g137) & (g936)) + ((!g34) & (g36) & (!reset) & (g137) & (g936)) + ((g34) & (!g36) & (!reset) & (g137) & (!g936)) + ((g34) & (!g36) & (!reset) & (g137) & (g936)) + ((g34) & (g36) & (!reset) & (g137) & (!g936)) + ((g34) & (g36) & (!reset) & (g137) & (g936)));
	assign g7333 = (((!g832) & (g2141) & (!g938)) + ((!g832) & (g2141) & (g938)) + ((g832) & (!g2141) & (g938)) + ((g832) & (g2141) & (g938)));
	assign g939 = (((!g34) & (!g36) & (!reset) & (g138) & (!g938)) + ((!g34) & (!g36) & (!reset) & (g138) & (g938)) + ((!g34) & (g36) & (!reset) & (!g138) & (g938)) + ((!g34) & (g36) & (!reset) & (g138) & (g938)) + ((g34) & (!g36) & (!reset) & (g138) & (!g938)) + ((g34) & (!g36) & (!reset) & (g138) & (g938)) + ((g34) & (g36) & (!reset) & (g138) & (!g938)) + ((g34) & (g36) & (!reset) & (g138) & (g938)));
	assign g7334 = (((!g832) & (g2143) & (!g940)) + ((!g832) & (g2143) & (g940)) + ((g832) & (!g2143) & (g940)) + ((g832) & (g2143) & (g940)));
	assign g941 = (((!g34) & (!g36) & (!reset) & (g140) & (!g940)) + ((!g34) & (!g36) & (!reset) & (g140) & (g940)) + ((!g34) & (g36) & (!reset) & (!g140) & (g940)) + ((!g34) & (g36) & (!reset) & (g140) & (g940)) + ((g34) & (!g36) & (!reset) & (g140) & (!g940)) + ((g34) & (!g36) & (!reset) & (g140) & (g940)) + ((g34) & (g36) & (!reset) & (g140) & (!g940)) + ((g34) & (g36) & (!reset) & (g140) & (g940)));
	assign g7335 = (((!g832) & (g2146) & (!g942)) + ((!g832) & (g2146) & (g942)) + ((g832) & (!g2146) & (g942)) + ((g832) & (g2146) & (g942)));
	assign g943 = (((!g34) & (!g36) & (!reset) & (g141) & (!g942)) + ((!g34) & (!g36) & (!reset) & (g141) & (g942)) + ((!g34) & (g36) & (!reset) & (!g141) & (g942)) + ((!g34) & (g36) & (!reset) & (g141) & (g942)) + ((g34) & (!g36) & (!reset) & (g141) & (!g942)) + ((g34) & (!g36) & (!reset) & (g141) & (g942)) + ((g34) & (g36) & (!reset) & (g141) & (!g942)) + ((g34) & (g36) & (!reset) & (g141) & (g942)));
	assign g7336 = (((!g832) & (g2149) & (!g944)) + ((!g832) & (g2149) & (g944)) + ((g832) & (!g2149) & (g944)) + ((g832) & (g2149) & (g944)));
	assign g945 = (((!g34) & (!g36) & (!reset) & (g142) & (!g944)) + ((!g34) & (!g36) & (!reset) & (g142) & (g944)) + ((!g34) & (g36) & (!reset) & (!g142) & (g944)) + ((!g34) & (g36) & (!reset) & (g142) & (g944)) + ((g34) & (!g36) & (!reset) & (g142) & (!g944)) + ((g34) & (!g36) & (!reset) & (g142) & (g944)) + ((g34) & (g36) & (!reset) & (g142) & (!g944)) + ((g34) & (g36) & (!reset) & (g142) & (g944)));
	assign g7337 = (((!g832) & (g2152) & (!g946)) + ((!g832) & (g2152) & (g946)) + ((g832) & (!g2152) & (g946)) + ((g832) & (g2152) & (g946)));
	assign g947 = (((!g34) & (!g36) & (!reset) & (g143) & (!g946)) + ((!g34) & (!g36) & (!reset) & (g143) & (g946)) + ((!g34) & (g36) & (!reset) & (!g143) & (g946)) + ((!g34) & (g36) & (!reset) & (g143) & (g946)) + ((g34) & (!g36) & (!reset) & (g143) & (!g946)) + ((g34) & (!g36) & (!reset) & (g143) & (g946)) + ((g34) & (g36) & (!reset) & (g143) & (!g946)) + ((g34) & (g36) & (!reset) & (g143) & (g946)));
	assign g7338 = (((!g832) & (g2155) & (!g948)) + ((!g832) & (g2155) & (g948)) + ((g832) & (!g2155) & (g948)) + ((g832) & (g2155) & (g948)));
	assign g949 = (((!g34) & (!g36) & (!reset) & (g145) & (!g948)) + ((!g34) & (!g36) & (!reset) & (g145) & (g948)) + ((!g34) & (g36) & (!reset) & (!g145) & (g948)) + ((!g34) & (g36) & (!reset) & (g145) & (g948)) + ((g34) & (!g36) & (!reset) & (g145) & (!g948)) + ((g34) & (!g36) & (!reset) & (g145) & (g948)) + ((g34) & (g36) & (!reset) & (g145) & (!g948)) + ((g34) & (g36) & (!reset) & (g145) & (g948)));
	assign g7339 = (((!g832) & (g2158) & (!g950)) + ((!g832) & (g2158) & (g950)) + ((g832) & (!g2158) & (g950)) + ((g832) & (g2158) & (g950)));
	assign g951 = (((!g34) & (!g36) & (!reset) & (g146) & (!g950)) + ((!g34) & (!g36) & (!reset) & (g146) & (g950)) + ((!g34) & (g36) & (!reset) & (!g146) & (g950)) + ((!g34) & (g36) & (!reset) & (g146) & (g950)) + ((g34) & (!g36) & (!reset) & (g146) & (!g950)) + ((g34) & (!g36) & (!reset) & (g146) & (g950)) + ((g34) & (g36) & (!reset) & (g146) & (!g950)) + ((g34) & (g36) & (!reset) & (g146) & (g950)));
	assign g7340 = (((!g832) & (g2161) & (!g952)) + ((!g832) & (g2161) & (g952)) + ((g832) & (!g2161) & (g952)) + ((g832) & (g2161) & (g952)));
	assign g953 = (((!g34) & (!g36) & (!reset) & (g147) & (!g952)) + ((!g34) & (!g36) & (!reset) & (g147) & (g952)) + ((!g34) & (g36) & (!reset) & (!g147) & (g952)) + ((!g34) & (g36) & (!reset) & (g147) & (g952)) + ((g34) & (!g36) & (!reset) & (g147) & (!g952)) + ((g34) & (!g36) & (!reset) & (g147) & (g952)) + ((g34) & (g36) & (!reset) & (g147) & (!g952)) + ((g34) & (g36) & (!reset) & (g147) & (g952)));
	assign g7341 = (((!g832) & (g2164) & (!g954)) + ((!g832) & (g2164) & (g954)) + ((g832) & (!g2164) & (g954)) + ((g832) & (g2164) & (g954)));
	assign g955 = (((!g34) & (!g36) & (!reset) & (g148) & (!g954)) + ((!g34) & (!g36) & (!reset) & (g148) & (g954)) + ((!g34) & (g36) & (!reset) & (!g148) & (g954)) + ((!g34) & (g36) & (!reset) & (g148) & (g954)) + ((g34) & (!g36) & (!reset) & (g148) & (!g954)) + ((g34) & (!g36) & (!reset) & (g148) & (g954)) + ((g34) & (g36) & (!reset) & (g148) & (!g954)) + ((g34) & (g36) & (!reset) & (g148) & (g954)));
	assign g7342 = (((!g832) & (g2166) & (!g956)) + ((!g832) & (g2166) & (g956)) + ((g832) & (!g2166) & (g956)) + ((g832) & (g2166) & (g956)));
	assign g957 = (((!g34) & (!g36) & (!reset) & (g150) & (!g956)) + ((!g34) & (!g36) & (!reset) & (g150) & (g956)) + ((!g34) & (g36) & (!reset) & (!g150) & (g956)) + ((!g34) & (g36) & (!reset) & (g150) & (g956)) + ((g34) & (!g36) & (!reset) & (g150) & (!g956)) + ((g34) & (!g36) & (!reset) & (g150) & (g956)) + ((g34) & (g36) & (!reset) & (g150) & (!g956)) + ((g34) & (g36) & (!reset) & (g150) & (g956)));
	assign g7343 = (((!g832) & (g2169) & (!g958)) + ((!g832) & (g2169) & (g958)) + ((g832) & (!g2169) & (g958)) + ((g832) & (g2169) & (g958)));
	assign g959 = (((!g34) & (!g36) & (!reset) & (g151) & (!g958)) + ((!g34) & (!g36) & (!reset) & (g151) & (g958)) + ((!g34) & (g36) & (!reset) & (!g151) & (g958)) + ((!g34) & (g36) & (!reset) & (g151) & (g958)) + ((g34) & (!g36) & (!reset) & (g151) & (!g958)) + ((g34) & (!g36) & (!reset) & (g151) & (g958)) + ((g34) & (g36) & (!reset) & (g151) & (!g958)) + ((g34) & (g36) & (!reset) & (g151) & (g958)));
	assign g7344 = (((!g832) & (g2172) & (!g960)) + ((!g832) & (g2172) & (g960)) + ((g832) & (!g2172) & (g960)) + ((g832) & (g2172) & (g960)));
	assign g961 = (((!g34) & (!g36) & (!reset) & (g152) & (!g960)) + ((!g34) & (!g36) & (!reset) & (g152) & (g960)) + ((!g34) & (g36) & (!reset) & (!g152) & (g960)) + ((!g34) & (g36) & (!reset) & (g152) & (g960)) + ((g34) & (!g36) & (!reset) & (g152) & (!g960)) + ((g34) & (!g36) & (!reset) & (g152) & (g960)) + ((g34) & (g36) & (!reset) & (g152) & (!g960)) + ((g34) & (g36) & (!reset) & (g152) & (g960)));
	assign g7345 = (((!g832) & (g2175) & (!g962)) + ((!g832) & (g2175) & (g962)) + ((g832) & (!g2175) & (g962)) + ((g832) & (g2175) & (g962)));
	assign g963 = (((!g34) & (!g36) & (!reset) & (g153) & (!g962)) + ((!g34) & (!g36) & (!reset) & (g153) & (g962)) + ((!g34) & (g36) & (!reset) & (!g153) & (g962)) + ((!g34) & (g36) & (!reset) & (g153) & (g962)) + ((g34) & (!g36) & (!reset) & (g153) & (!g962)) + ((g34) & (!g36) & (!reset) & (g153) & (g962)) + ((g34) & (g36) & (!reset) & (g153) & (!g962)) + ((g34) & (g36) & (!reset) & (g153) & (g962)));
	assign g7346 = (((!g2017) & (g7165) & (!g964)) + ((!g2017) & (g7165) & (g964)) + ((g2017) & (!g7165) & (g964)) + ((g2017) & (g7165) & (g964)));
	assign g965 = (((!g110) & (!g133) & (g897) & (g931) & (g898)) + ((!g110) & (g133) & (!g897) & (g931) & (!g898)) + ((!g110) & (g133) & (!g897) & (g931) & (g898)) + ((!g110) & (g133) & (g897) & (!g931) & (g898)) + ((!g110) & (g133) & (g897) & (g931) & (!g898)) + ((!g110) & (g133) & (g897) & (g931) & (g898)) + ((g110) & (!g133) & (!g897) & (g931) & (g898)) + ((g110) & (!g133) & (g897) & (g931) & (!g898)) + ((g110) & (!g133) & (g897) & (g931) & (g898)) + ((g110) & (g133) & (!g897) & (!g931) & (g898)) + ((g110) & (g133) & (!g897) & (g931) & (!g898)) + ((g110) & (g133) & (!g897) & (g931) & (g898)) + ((g110) & (g133) & (g897) & (!g931) & (!g898)) + ((g110) & (g133) & (g897) & (!g931) & (g898)) + ((g110) & (g133) & (g897) & (g931) & (!g898)) + ((g110) & (g133) & (g897) & (g931) & (g898)));
	assign g966 = (((!g827) & (!g156) & (g964) & (!g965)) + ((!g827) & (!g156) & (g964) & (g965)) + ((!g827) & (g156) & (g964) & (!g965)) + ((!g827) & (g156) & (g964) & (g965)) + ((g827) & (!g156) & (!g964) & (g965)) + ((g827) & (!g156) & (g964) & (!g965)) + ((g827) & (g156) & (!g964) & (!g965)) + ((g827) & (g156) & (g964) & (g965)));
	assign g967 = (((!g34) & (!g36) & (!reset) & (g158) & (!g179)) + ((!g34) & (!g36) & (!reset) & (g158) & (g179)) + ((!g34) & (g36) & (!reset) & (!g158) & (g179)) + ((!g34) & (g36) & (!reset) & (g158) & (g179)) + ((g34) & (!g36) & (!reset) & (g158) & (!g179)) + ((g34) & (!g36) & (!reset) & (g158) & (g179)) + ((g34) & (g36) & (!reset) & (g158) & (!g179)) + ((g34) & (g36) & (!reset) & (g158) & (g179)));
	assign g7347 = (((!g832) & (g2183) & (!g968)) + ((!g832) & (g2183) & (g968)) + ((g832) & (!g2183) & (g968)) + ((g832) & (g2183) & (g968)));
	assign g969 = (((!g34) & (!g36) & (!reset) & (g159) & (!g968)) + ((!g34) & (!g36) & (!reset) & (g159) & (g968)) + ((!g34) & (g36) & (!reset) & (!g159) & (g968)) + ((!g34) & (g36) & (!reset) & (g159) & (g968)) + ((g34) & (!g36) & (!reset) & (g159) & (!g968)) + ((g34) & (!g36) & (!reset) & (g159) & (g968)) + ((g34) & (g36) & (!reset) & (g159) & (!g968)) + ((g34) & (g36) & (!reset) & (g159) & (g968)));
	assign g7348 = (((!g832) & (g2185) & (!g970)) + ((!g832) & (g2185) & (g970)) + ((g832) & (!g2185) & (g970)) + ((g832) & (g2185) & (g970)));
	assign g971 = (((!g34) & (!g36) & (!reset) & (g160) & (!g970)) + ((!g34) & (!g36) & (!reset) & (g160) & (g970)) + ((!g34) & (g36) & (!reset) & (!g160) & (g970)) + ((!g34) & (g36) & (!reset) & (g160) & (g970)) + ((g34) & (!g36) & (!reset) & (g160) & (!g970)) + ((g34) & (!g36) & (!reset) & (g160) & (g970)) + ((g34) & (g36) & (!reset) & (g160) & (!g970)) + ((g34) & (g36) & (!reset) & (g160) & (g970)));
	assign g7349 = (((!g832) & (g2186) & (!g972)) + ((!g832) & (g2186) & (g972)) + ((g832) & (!g2186) & (g972)) + ((g832) & (g2186) & (g972)));
	assign g973 = (((!g34) & (!g36) & (!reset) & (g161) & (!g972)) + ((!g34) & (!g36) & (!reset) & (g161) & (g972)) + ((!g34) & (g36) & (!reset) & (!g161) & (g972)) + ((!g34) & (g36) & (!reset) & (g161) & (g972)) + ((g34) & (!g36) & (!reset) & (g161) & (!g972)) + ((g34) & (!g36) & (!reset) & (g161) & (g972)) + ((g34) & (g36) & (!reset) & (g161) & (!g972)) + ((g34) & (g36) & (!reset) & (g161) & (g972)));
	assign g7350 = (((!g832) & (g2187) & (!g974)) + ((!g832) & (g2187) & (g974)) + ((g832) & (!g2187) & (g974)) + ((g832) & (g2187) & (g974)));
	assign g975 = (((!g34) & (!g36) & (!reset) & (g163) & (!g974)) + ((!g34) & (!g36) & (!reset) & (g163) & (g974)) + ((!g34) & (g36) & (!reset) & (!g163) & (g974)) + ((!g34) & (g36) & (!reset) & (g163) & (g974)) + ((g34) & (!g36) & (!reset) & (g163) & (!g974)) + ((g34) & (!g36) & (!reset) & (g163) & (g974)) + ((g34) & (g36) & (!reset) & (g163) & (!g974)) + ((g34) & (g36) & (!reset) & (g163) & (g974)));
	assign g7351 = (((!g832) & (g2189) & (!g976)) + ((!g832) & (g2189) & (g976)) + ((g832) & (!g2189) & (g976)) + ((g832) & (g2189) & (g976)));
	assign g977 = (((!g34) & (!g36) & (!reset) & (g164) & (!g976)) + ((!g34) & (!g36) & (!reset) & (g164) & (g976)) + ((!g34) & (g36) & (!reset) & (!g164) & (g976)) + ((!g34) & (g36) & (!reset) & (g164) & (g976)) + ((g34) & (!g36) & (!reset) & (g164) & (!g976)) + ((g34) & (!g36) & (!reset) & (g164) & (g976)) + ((g34) & (g36) & (!reset) & (g164) & (!g976)) + ((g34) & (g36) & (!reset) & (g164) & (g976)));
	assign g7352 = (((!g832) & (g2191) & (!g978)) + ((!g832) & (g2191) & (g978)) + ((g832) & (!g2191) & (g978)) + ((g832) & (g2191) & (g978)));
	assign g979 = (((!g34) & (!g36) & (!reset) & (g165) & (!g978)) + ((!g34) & (!g36) & (!reset) & (g165) & (g978)) + ((!g34) & (g36) & (!reset) & (!g165) & (g978)) + ((!g34) & (g36) & (!reset) & (g165) & (g978)) + ((g34) & (!g36) & (!reset) & (g165) & (!g978)) + ((g34) & (!g36) & (!reset) & (g165) & (g978)) + ((g34) & (g36) & (!reset) & (g165) & (!g978)) + ((g34) & (g36) & (!reset) & (g165) & (g978)));
	assign g7353 = (((!g832) & (g2193) & (!g980)) + ((!g832) & (g2193) & (g980)) + ((g832) & (!g2193) & (g980)) + ((g832) & (g2193) & (g980)));
	assign g981 = (((!g34) & (!g36) & (!reset) & (g166) & (!g980)) + ((!g34) & (!g36) & (!reset) & (g166) & (g980)) + ((!g34) & (g36) & (!reset) & (!g166) & (g980)) + ((!g34) & (g36) & (!reset) & (g166) & (g980)) + ((g34) & (!g36) & (!reset) & (g166) & (!g980)) + ((g34) & (!g36) & (!reset) & (g166) & (g980)) + ((g34) & (g36) & (!reset) & (g166) & (!g980)) + ((g34) & (g36) & (!reset) & (g166) & (g980)));
	assign g7354 = (((!g832) & (g2195) & (!g982)) + ((!g832) & (g2195) & (g982)) + ((g832) & (!g2195) & (g982)) + ((g832) & (g2195) & (g982)));
	assign g983 = (((!g34) & (!g36) & (!reset) & (g168) & (!g982)) + ((!g34) & (!g36) & (!reset) & (g168) & (g982)) + ((!g34) & (g36) & (!reset) & (!g168) & (g982)) + ((!g34) & (g36) & (!reset) & (g168) & (g982)) + ((g34) & (!g36) & (!reset) & (g168) & (!g982)) + ((g34) & (!g36) & (!reset) & (g168) & (g982)) + ((g34) & (g36) & (!reset) & (g168) & (!g982)) + ((g34) & (g36) & (!reset) & (g168) & (g982)));
	assign g7355 = (((!g832) & (g2197) & (!g984)) + ((!g832) & (g2197) & (g984)) + ((g832) & (!g2197) & (g984)) + ((g832) & (g2197) & (g984)));
	assign g985 = (((!g34) & (!g36) & (!reset) & (g169) & (!g984)) + ((!g34) & (!g36) & (!reset) & (g169) & (g984)) + ((!g34) & (g36) & (!reset) & (!g169) & (g984)) + ((!g34) & (g36) & (!reset) & (g169) & (g984)) + ((g34) & (!g36) & (!reset) & (g169) & (!g984)) + ((g34) & (!g36) & (!reset) & (g169) & (g984)) + ((g34) & (g36) & (!reset) & (g169) & (!g984)) + ((g34) & (g36) & (!reset) & (g169) & (g984)));
	assign g7356 = (((!g832) & (g2199) & (!g986)) + ((!g832) & (g2199) & (g986)) + ((g832) & (!g2199) & (g986)) + ((g832) & (g2199) & (g986)));
	assign g987 = (((!g34) & (!g36) & (!reset) & (g170) & (!g986)) + ((!g34) & (!g36) & (!reset) & (g170) & (g986)) + ((!g34) & (g36) & (!reset) & (!g170) & (g986)) + ((!g34) & (g36) & (!reset) & (g170) & (g986)) + ((g34) & (!g36) & (!reset) & (g170) & (!g986)) + ((g34) & (!g36) & (!reset) & (g170) & (g986)) + ((g34) & (g36) & (!reset) & (g170) & (!g986)) + ((g34) & (g36) & (!reset) & (g170) & (g986)));
	assign g7357 = (((!g832) & (g2201) & (!g988)) + ((!g832) & (g2201) & (g988)) + ((g832) & (!g2201) & (g988)) + ((g832) & (g2201) & (g988)));
	assign g989 = (((!g34) & (!g36) & (!reset) & (g171) & (!g988)) + ((!g34) & (!g36) & (!reset) & (g171) & (g988)) + ((!g34) & (g36) & (!reset) & (!g171) & (g988)) + ((!g34) & (g36) & (!reset) & (g171) & (g988)) + ((g34) & (!g36) & (!reset) & (g171) & (!g988)) + ((g34) & (!g36) & (!reset) & (g171) & (g988)) + ((g34) & (g36) & (!reset) & (g171) & (!g988)) + ((g34) & (g36) & (!reset) & (g171) & (g988)));
	assign g7358 = (((!g832) & (g2202) & (!g990)) + ((!g832) & (g2202) & (g990)) + ((g832) & (!g2202) & (g990)) + ((g832) & (g2202) & (g990)));
	assign g991 = (((!g34) & (!g36) & (!reset) & (g173) & (!g990)) + ((!g34) & (!g36) & (!reset) & (g173) & (g990)) + ((!g34) & (g36) & (!reset) & (!g173) & (g990)) + ((!g34) & (g36) & (!reset) & (g173) & (g990)) + ((g34) & (!g36) & (!reset) & (g173) & (!g990)) + ((g34) & (!g36) & (!reset) & (g173) & (g990)) + ((g34) & (g36) & (!reset) & (g173) & (!g990)) + ((g34) & (g36) & (!reset) & (g173) & (g990)));
	assign g7359 = (((!g832) & (g2204) & (!g992)) + ((!g832) & (g2204) & (g992)) + ((g832) & (!g2204) & (g992)) + ((g832) & (g2204) & (g992)));
	assign g993 = (((!g34) & (!g36) & (!reset) & (g174) & (!g992)) + ((!g34) & (!g36) & (!reset) & (g174) & (g992)) + ((!g34) & (g36) & (!reset) & (!g174) & (g992)) + ((!g34) & (g36) & (!reset) & (g174) & (g992)) + ((g34) & (!g36) & (!reset) & (g174) & (!g992)) + ((g34) & (!g36) & (!reset) & (g174) & (g992)) + ((g34) & (g36) & (!reset) & (g174) & (!g992)) + ((g34) & (g36) & (!reset) & (g174) & (g992)));
	assign g7360 = (((!g832) & (g2206) & (!g994)) + ((!g832) & (g2206) & (g994)) + ((g832) & (!g2206) & (g994)) + ((g832) & (g2206) & (g994)));
	assign g995 = (((!g34) & (!g36) & (!reset) & (g175) & (!g994)) + ((!g34) & (!g36) & (!reset) & (g175) & (g994)) + ((!g34) & (g36) & (!reset) & (!g175) & (g994)) + ((!g34) & (g36) & (!reset) & (g175) & (g994)) + ((g34) & (!g36) & (!reset) & (g175) & (!g994)) + ((g34) & (!g36) & (!reset) & (g175) & (g994)) + ((g34) & (g36) & (!reset) & (g175) & (!g994)) + ((g34) & (g36) & (!reset) & (g175) & (g994)));
	assign g7361 = (((!g832) & (g2208) & (!g996)) + ((!g832) & (g2208) & (g996)) + ((g832) & (!g2208) & (g996)) + ((g832) & (g2208) & (g996)));
	assign g997 = (((!g34) & (!g36) & (!reset) & (g176) & (!g996)) + ((!g34) & (!g36) & (!reset) & (g176) & (g996)) + ((!g34) & (g36) & (!reset) & (!g176) & (g996)) + ((!g34) & (g36) & (!reset) & (g176) & (g996)) + ((g34) & (!g36) & (!reset) & (g176) & (!g996)) + ((g34) & (!g36) & (!reset) & (g176) & (g996)) + ((g34) & (g36) & (!reset) & (g176) & (!g996)) + ((g34) & (g36) & (!reset) & (g176) & (g996)));
	assign g7362 = (((!g2017) & (g7158) & (!g998)) + ((!g2017) & (g7158) & (g998)) + ((g2017) & (!g7158) & (g998)) + ((g2017) & (g7158) & (g998)));
	assign g999 = (((!g827) & (!g156) & (!g179) & (!g964) & (g998) & (!g965)) + ((!g827) & (!g156) & (!g179) & (!g964) & (g998) & (g965)) + ((!g827) & (!g156) & (!g179) & (g964) & (g998) & (!g965)) + ((!g827) & (!g156) & (!g179) & (g964) & (g998) & (g965)) + ((!g827) & (!g156) & (g179) & (!g964) & (g998) & (!g965)) + ((!g827) & (!g156) & (g179) & (!g964) & (g998) & (g965)) + ((!g827) & (!g156) & (g179) & (g964) & (g998) & (!g965)) + ((!g827) & (!g156) & (g179) & (g964) & (g998) & (g965)) + ((!g827) & (g156) & (!g179) & (!g964) & (g998) & (!g965)) + ((!g827) & (g156) & (!g179) & (!g964) & (g998) & (g965)) + ((!g827) & (g156) & (!g179) & (g964) & (g998) & (!g965)) + ((!g827) & (g156) & (!g179) & (g964) & (g998) & (g965)) + ((!g827) & (g156) & (g179) & (!g964) & (g998) & (!g965)) + ((!g827) & (g156) & (g179) & (!g964) & (g998) & (g965)) + ((!g827) & (g156) & (g179) & (g964) & (g998) & (!g965)) + ((!g827) & (g156) & (g179) & (g964) & (g998) & (g965)) + ((g827) & (!g156) & (!g179) & (!g964) & (g998) & (!g965)) + ((g827) & (!g156) & (!g179) & (!g964) & (g998) & (g965)) + ((g827) & (!g156) & (!g179) & (g964) & (!g998) & (g965)) + ((g827) & (!g156) & (!g179) & (g964) & (g998) & (!g965)) + ((g827) & (!g156) & (g179) & (!g964) & (!g998) & (!g965)) + ((g827) & (!g156) & (g179) & (!g964) & (!g998) & (g965)) + ((g827) & (!g156) & (g179) & (g964) & (!g998) & (!g965)) + ((g827) & (!g156) & (g179) & (g964) & (g998) & (g965)) + ((g827) & (g156) & (!g179) & (!g964) & (!g998) & (g965)) + ((g827) & (g156) & (!g179) & (!g964) & (g998) & (!g965)) + ((g827) & (g156) & (!g179) & (g964) & (!g998) & (!g965)) + ((g827) & (g156) & (!g179) & (g964) & (!g998) & (g965)) + ((g827) & (g156) & (g179) & (!g964) & (!g998) & (!g965)) + ((g827) & (g156) & (g179) & (!g964) & (g998) & (g965)) + ((g827) & (g156) & (g179) & (g964) & (g998) & (!g965)) + ((g827) & (g156) & (g179) & (g964) & (g998) & (g965)));
	assign g1000 = (((!g34) & (!g36) & (!reset) & (g181) & (!g202)) + ((!g34) & (!g36) & (!reset) & (g181) & (g202)) + ((!g34) & (g36) & (!reset) & (!g181) & (g202)) + ((!g34) & (g36) & (!reset) & (g181) & (g202)) + ((g34) & (!g36) & (!reset) & (g181) & (!g202)) + ((g34) & (!g36) & (!reset) & (g181) & (g202)) + ((g34) & (g36) & (!reset) & (g181) & (!g202)) + ((g34) & (g36) & (!reset) & (g181) & (g202)));
	assign g7363 = (((!g832) & (g2216) & (!g1001)) + ((!g832) & (g2216) & (g1001)) + ((g832) & (!g2216) & (g1001)) + ((g832) & (g2216) & (g1001)));
	assign g1002 = (((!g34) & (!g36) & (!reset) & (g182) & (!g1001)) + ((!g34) & (!g36) & (!reset) & (g182) & (g1001)) + ((!g34) & (g36) & (!reset) & (!g182) & (g1001)) + ((!g34) & (g36) & (!reset) & (g182) & (g1001)) + ((g34) & (!g36) & (!reset) & (g182) & (!g1001)) + ((g34) & (!g36) & (!reset) & (g182) & (g1001)) + ((g34) & (g36) & (!reset) & (g182) & (!g1001)) + ((g34) & (g36) & (!reset) & (g182) & (g1001)));
	assign g7364 = (((!g832) & (g2219) & (!g1003)) + ((!g832) & (g2219) & (g1003)) + ((g832) & (!g2219) & (g1003)) + ((g832) & (g2219) & (g1003)));
	assign g1004 = (((!g34) & (!g36) & (!reset) & (g183) & (!g1003)) + ((!g34) & (!g36) & (!reset) & (g183) & (g1003)) + ((!g34) & (g36) & (!reset) & (!g183) & (g1003)) + ((!g34) & (g36) & (!reset) & (g183) & (g1003)) + ((g34) & (!g36) & (!reset) & (g183) & (!g1003)) + ((g34) & (!g36) & (!reset) & (g183) & (g1003)) + ((g34) & (g36) & (!reset) & (g183) & (!g1003)) + ((g34) & (g36) & (!reset) & (g183) & (g1003)));
	assign g7365 = (((!g832) & (g2221) & (!g1005)) + ((!g832) & (g2221) & (g1005)) + ((g832) & (!g2221) & (g1005)) + ((g832) & (g2221) & (g1005)));
	assign g1006 = (((!g34) & (!g36) & (!reset) & (g184) & (!g1005)) + ((!g34) & (!g36) & (!reset) & (g184) & (g1005)) + ((!g34) & (g36) & (!reset) & (!g184) & (g1005)) + ((!g34) & (g36) & (!reset) & (g184) & (g1005)) + ((g34) & (!g36) & (!reset) & (g184) & (!g1005)) + ((g34) & (!g36) & (!reset) & (g184) & (g1005)) + ((g34) & (g36) & (!reset) & (g184) & (!g1005)) + ((g34) & (g36) & (!reset) & (g184) & (g1005)));
	assign g7366 = (((!g832) & (g2223) & (!g1007)) + ((!g832) & (g2223) & (g1007)) + ((g832) & (!g2223) & (g1007)) + ((g832) & (g2223) & (g1007)));
	assign g1008 = (((!g34) & (!g36) & (!reset) & (g186) & (!g1007)) + ((!g34) & (!g36) & (!reset) & (g186) & (g1007)) + ((!g34) & (g36) & (!reset) & (!g186) & (g1007)) + ((!g34) & (g36) & (!reset) & (g186) & (g1007)) + ((g34) & (!g36) & (!reset) & (g186) & (!g1007)) + ((g34) & (!g36) & (!reset) & (g186) & (g1007)) + ((g34) & (g36) & (!reset) & (g186) & (!g1007)) + ((g34) & (g36) & (!reset) & (g186) & (g1007)));
	assign g7367 = (((!g832) & (g2226) & (!g1009)) + ((!g832) & (g2226) & (g1009)) + ((g832) & (!g2226) & (g1009)) + ((g832) & (g2226) & (g1009)));
	assign g1010 = (((!g34) & (!g36) & (!reset) & (g187) & (!g1009)) + ((!g34) & (!g36) & (!reset) & (g187) & (g1009)) + ((!g34) & (g36) & (!reset) & (!g187) & (g1009)) + ((!g34) & (g36) & (!reset) & (g187) & (g1009)) + ((g34) & (!g36) & (!reset) & (g187) & (!g1009)) + ((g34) & (!g36) & (!reset) & (g187) & (g1009)) + ((g34) & (g36) & (!reset) & (g187) & (!g1009)) + ((g34) & (g36) & (!reset) & (g187) & (g1009)));
	assign g7368 = (((!g832) & (g2229) & (!g1011)) + ((!g832) & (g2229) & (g1011)) + ((g832) & (!g2229) & (g1011)) + ((g832) & (g2229) & (g1011)));
	assign g1012 = (((!g34) & (!g36) & (!reset) & (g188) & (!g1011)) + ((!g34) & (!g36) & (!reset) & (g188) & (g1011)) + ((!g34) & (g36) & (!reset) & (!g188) & (g1011)) + ((!g34) & (g36) & (!reset) & (g188) & (g1011)) + ((g34) & (!g36) & (!reset) & (g188) & (!g1011)) + ((g34) & (!g36) & (!reset) & (g188) & (g1011)) + ((g34) & (g36) & (!reset) & (g188) & (!g1011)) + ((g34) & (g36) & (!reset) & (g188) & (g1011)));
	assign g7369 = (((!g832) & (g2232) & (!g1013)) + ((!g832) & (g2232) & (g1013)) + ((g832) & (!g2232) & (g1013)) + ((g832) & (g2232) & (g1013)));
	assign g1014 = (((!g34) & (!g36) & (!reset) & (g189) & (!g1013)) + ((!g34) & (!g36) & (!reset) & (g189) & (g1013)) + ((!g34) & (g36) & (!reset) & (!g189) & (g1013)) + ((!g34) & (g36) & (!reset) & (g189) & (g1013)) + ((g34) & (!g36) & (!reset) & (g189) & (!g1013)) + ((g34) & (!g36) & (!reset) & (g189) & (g1013)) + ((g34) & (g36) & (!reset) & (g189) & (!g1013)) + ((g34) & (g36) & (!reset) & (g189) & (g1013)));
	assign g7370 = (((!g832) & (g2235) & (!g1015)) + ((!g832) & (g2235) & (g1015)) + ((g832) & (!g2235) & (g1015)) + ((g832) & (g2235) & (g1015)));
	assign g1016 = (((!g34) & (!g36) & (!reset) & (g191) & (!g1015)) + ((!g34) & (!g36) & (!reset) & (g191) & (g1015)) + ((!g34) & (g36) & (!reset) & (!g191) & (g1015)) + ((!g34) & (g36) & (!reset) & (g191) & (g1015)) + ((g34) & (!g36) & (!reset) & (g191) & (!g1015)) + ((g34) & (!g36) & (!reset) & (g191) & (g1015)) + ((g34) & (g36) & (!reset) & (g191) & (!g1015)) + ((g34) & (g36) & (!reset) & (g191) & (g1015)));
	assign g7371 = (((!g832) & (g2238) & (!g1017)) + ((!g832) & (g2238) & (g1017)) + ((g832) & (!g2238) & (g1017)) + ((g832) & (g2238) & (g1017)));
	assign g1018 = (((!g34) & (!g36) & (!reset) & (g192) & (!g1017)) + ((!g34) & (!g36) & (!reset) & (g192) & (g1017)) + ((!g34) & (g36) & (!reset) & (!g192) & (g1017)) + ((!g34) & (g36) & (!reset) & (g192) & (g1017)) + ((g34) & (!g36) & (!reset) & (g192) & (!g1017)) + ((g34) & (!g36) & (!reset) & (g192) & (g1017)) + ((g34) & (g36) & (!reset) & (g192) & (!g1017)) + ((g34) & (g36) & (!reset) & (g192) & (g1017)));
	assign g7372 = (((!g832) & (g2241) & (!g1019)) + ((!g832) & (g2241) & (g1019)) + ((g832) & (!g2241) & (g1019)) + ((g832) & (g2241) & (g1019)));
	assign g1020 = (((!g34) & (!g36) & (!reset) & (g193) & (!g1019)) + ((!g34) & (!g36) & (!reset) & (g193) & (g1019)) + ((!g34) & (g36) & (!reset) & (!g193) & (g1019)) + ((!g34) & (g36) & (!reset) & (g193) & (g1019)) + ((g34) & (!g36) & (!reset) & (g193) & (!g1019)) + ((g34) & (!g36) & (!reset) & (g193) & (g1019)) + ((g34) & (g36) & (!reset) & (g193) & (!g1019)) + ((g34) & (g36) & (!reset) & (g193) & (g1019)));
	assign g7373 = (((!g832) & (g2244) & (!g1021)) + ((!g832) & (g2244) & (g1021)) + ((g832) & (!g2244) & (g1021)) + ((g832) & (g2244) & (g1021)));
	assign g1022 = (((!g34) & (!g36) & (!reset) & (g194) & (!g1021)) + ((!g34) & (!g36) & (!reset) & (g194) & (g1021)) + ((!g34) & (g36) & (!reset) & (!g194) & (g1021)) + ((!g34) & (g36) & (!reset) & (g194) & (g1021)) + ((g34) & (!g36) & (!reset) & (g194) & (!g1021)) + ((g34) & (!g36) & (!reset) & (g194) & (g1021)) + ((g34) & (g36) & (!reset) & (g194) & (!g1021)) + ((g34) & (g36) & (!reset) & (g194) & (g1021)));
	assign g7374 = (((!g832) & (g2246) & (!g1023)) + ((!g832) & (g2246) & (g1023)) + ((g832) & (!g2246) & (g1023)) + ((g832) & (g2246) & (g1023)));
	assign g1024 = (((!g34) & (!g36) & (!reset) & (g196) & (!g1023)) + ((!g34) & (!g36) & (!reset) & (g196) & (g1023)) + ((!g34) & (g36) & (!reset) & (!g196) & (g1023)) + ((!g34) & (g36) & (!reset) & (g196) & (g1023)) + ((g34) & (!g36) & (!reset) & (g196) & (!g1023)) + ((g34) & (!g36) & (!reset) & (g196) & (g1023)) + ((g34) & (g36) & (!reset) & (g196) & (!g1023)) + ((g34) & (g36) & (!reset) & (g196) & (g1023)));
	assign g7375 = (((!g832) & (g2249) & (!g1025)) + ((!g832) & (g2249) & (g1025)) + ((g832) & (!g2249) & (g1025)) + ((g832) & (g2249) & (g1025)));
	assign g1026 = (((!g34) & (!g36) & (!reset) & (g197) & (!g1025)) + ((!g34) & (!g36) & (!reset) & (g197) & (g1025)) + ((!g34) & (g36) & (!reset) & (!g197) & (g1025)) + ((!g34) & (g36) & (!reset) & (g197) & (g1025)) + ((g34) & (!g36) & (!reset) & (g197) & (!g1025)) + ((g34) & (!g36) & (!reset) & (g197) & (g1025)) + ((g34) & (g36) & (!reset) & (g197) & (!g1025)) + ((g34) & (g36) & (!reset) & (g197) & (g1025)));
	assign g7376 = (((!g832) & (g2252) & (!g1027)) + ((!g832) & (g2252) & (g1027)) + ((g832) & (!g2252) & (g1027)) + ((g832) & (g2252) & (g1027)));
	assign g1028 = (((!g34) & (!g36) & (!reset) & (g198) & (!g1027)) + ((!g34) & (!g36) & (!reset) & (g198) & (g1027)) + ((!g34) & (g36) & (!reset) & (!g198) & (g1027)) + ((!g34) & (g36) & (!reset) & (g198) & (g1027)) + ((g34) & (!g36) & (!reset) & (g198) & (!g1027)) + ((g34) & (!g36) & (!reset) & (g198) & (g1027)) + ((g34) & (g36) & (!reset) & (g198) & (!g1027)) + ((g34) & (g36) & (!reset) & (g198) & (g1027)));
	assign g7377 = (((!g832) & (g2255) & (!g1029)) + ((!g832) & (g2255) & (g1029)) + ((g832) & (!g2255) & (g1029)) + ((g832) & (g2255) & (g1029)));
	assign g1030 = (((!g34) & (!g36) & (!reset) & (g199) & (!g1029)) + ((!g34) & (!g36) & (!reset) & (g199) & (g1029)) + ((!g34) & (g36) & (!reset) & (!g199) & (g1029)) + ((!g34) & (g36) & (!reset) & (g199) & (g1029)) + ((g34) & (!g36) & (!reset) & (g199) & (!g1029)) + ((g34) & (!g36) & (!reset) & (g199) & (g1029)) + ((g34) & (g36) & (!reset) & (g199) & (!g1029)) + ((g34) & (g36) & (!reset) & (g199) & (g1029)));
	assign g7378 = (((!g2017) & (g2265) & (!g1031)) + ((!g2017) & (g2265) & (g1031)) + ((g2017) & (!g2265) & (g1031)) + ((g2017) & (g2265) & (g1031)));
	assign g1032 = (((!g156) & (!g179) & (g964) & (g998) & (g965)) + ((!g156) & (g179) & (!g964) & (g998) & (!g965)) + ((!g156) & (g179) & (!g964) & (g998) & (g965)) + ((!g156) & (g179) & (g964) & (!g998) & (g965)) + ((!g156) & (g179) & (g964) & (g998) & (!g965)) + ((!g156) & (g179) & (g964) & (g998) & (g965)) + ((g156) & (!g179) & (!g964) & (g998) & (g965)) + ((g156) & (!g179) & (g964) & (g998) & (!g965)) + ((g156) & (!g179) & (g964) & (g998) & (g965)) + ((g156) & (g179) & (!g964) & (!g998) & (g965)) + ((g156) & (g179) & (!g964) & (g998) & (!g965)) + ((g156) & (g179) & (!g964) & (g998) & (g965)) + ((g156) & (g179) & (g964) & (!g998) & (!g965)) + ((g156) & (g179) & (g964) & (!g998) & (g965)) + ((g156) & (g179) & (g964) & (g998) & (!g965)) + ((g156) & (g179) & (g964) & (g998) & (g965)));
	assign g1033 = (((!g827) & (!g202) & (g1031) & (!g1032)) + ((!g827) & (!g202) & (g1031) & (g1032)) + ((!g827) & (g202) & (g1031) & (!g1032)) + ((!g827) & (g202) & (g1031) & (g1032)) + ((g827) & (!g202) & (!g1031) & (g1032)) + ((g827) & (!g202) & (g1031) & (!g1032)) + ((g827) & (g202) & (!g1031) & (!g1032)) + ((g827) & (g202) & (g1031) & (g1032)));
	assign g1034 = (((!g34) & (!g36) & (!reset) & (g204) & (!g225)) + ((!g34) & (!g36) & (!reset) & (g204) & (g225)) + ((!g34) & (g36) & (!reset) & (!g204) & (g225)) + ((!g34) & (g36) & (!reset) & (g204) & (g225)) + ((g34) & (!g36) & (!reset) & (g204) & (!g225)) + ((g34) & (!g36) & (!reset) & (g204) & (g225)) + ((g34) & (g36) & (!reset) & (g204) & (!g225)) + ((g34) & (g36) & (!reset) & (g204) & (g225)));
	assign g7379 = (((!g832) & (g2266) & (!g1035)) + ((!g832) & (g2266) & (g1035)) + ((g832) & (!g2266) & (g1035)) + ((g832) & (g2266) & (g1035)));
	assign g1036 = (((!g34) & (!g36) & (!reset) & (g205) & (!g1035)) + ((!g34) & (!g36) & (!reset) & (g205) & (g1035)) + ((!g34) & (g36) & (!reset) & (!g205) & (g1035)) + ((!g34) & (g36) & (!reset) & (g205) & (g1035)) + ((g34) & (!g36) & (!reset) & (g205) & (!g1035)) + ((g34) & (!g36) & (!reset) & (g205) & (g1035)) + ((g34) & (g36) & (!reset) & (g205) & (!g1035)) + ((g34) & (g36) & (!reset) & (g205) & (g1035)));
	assign g7380 = (((!g832) & (g2268) & (!g1037)) + ((!g832) & (g2268) & (g1037)) + ((g832) & (!g2268) & (g1037)) + ((g832) & (g2268) & (g1037)));
	assign g1038 = (((!g34) & (!g36) & (!reset) & (g206) & (!g1037)) + ((!g34) & (!g36) & (!reset) & (g206) & (g1037)) + ((!g34) & (g36) & (!reset) & (!g206) & (g1037)) + ((!g34) & (g36) & (!reset) & (g206) & (g1037)) + ((g34) & (!g36) & (!reset) & (g206) & (!g1037)) + ((g34) & (!g36) & (!reset) & (g206) & (g1037)) + ((g34) & (g36) & (!reset) & (g206) & (!g1037)) + ((g34) & (g36) & (!reset) & (g206) & (g1037)));
	assign g7381 = (((!g832) & (g2269) & (!g1039)) + ((!g832) & (g2269) & (g1039)) + ((g832) & (!g2269) & (g1039)) + ((g832) & (g2269) & (g1039)));
	assign g1040 = (((!g34) & (!g36) & (!reset) & (g207) & (!g1039)) + ((!g34) & (!g36) & (!reset) & (g207) & (g1039)) + ((!g34) & (g36) & (!reset) & (!g207) & (g1039)) + ((!g34) & (g36) & (!reset) & (g207) & (g1039)) + ((g34) & (!g36) & (!reset) & (g207) & (!g1039)) + ((g34) & (!g36) & (!reset) & (g207) & (g1039)) + ((g34) & (g36) & (!reset) & (g207) & (!g1039)) + ((g34) & (g36) & (!reset) & (g207) & (g1039)));
	assign g7382 = (((!g832) & (g2270) & (!g1041)) + ((!g832) & (g2270) & (g1041)) + ((g832) & (!g2270) & (g1041)) + ((g832) & (g2270) & (g1041)));
	assign g1042 = (((!g34) & (!g36) & (!reset) & (g209) & (!g1041)) + ((!g34) & (!g36) & (!reset) & (g209) & (g1041)) + ((!g34) & (g36) & (!reset) & (!g209) & (g1041)) + ((!g34) & (g36) & (!reset) & (g209) & (g1041)) + ((g34) & (!g36) & (!reset) & (g209) & (!g1041)) + ((g34) & (!g36) & (!reset) & (g209) & (g1041)) + ((g34) & (g36) & (!reset) & (g209) & (!g1041)) + ((g34) & (g36) & (!reset) & (g209) & (g1041)));
	assign g7383 = (((!g832) & (g2272) & (!g1043)) + ((!g832) & (g2272) & (g1043)) + ((g832) & (!g2272) & (g1043)) + ((g832) & (g2272) & (g1043)));
	assign g1044 = (((!g34) & (!g36) & (!reset) & (g210) & (!g1043)) + ((!g34) & (!g36) & (!reset) & (g210) & (g1043)) + ((!g34) & (g36) & (!reset) & (!g210) & (g1043)) + ((!g34) & (g36) & (!reset) & (g210) & (g1043)) + ((g34) & (!g36) & (!reset) & (g210) & (!g1043)) + ((g34) & (!g36) & (!reset) & (g210) & (g1043)) + ((g34) & (g36) & (!reset) & (g210) & (!g1043)) + ((g34) & (g36) & (!reset) & (g210) & (g1043)));
	assign g7384 = (((!g832) & (g2274) & (!g1045)) + ((!g832) & (g2274) & (g1045)) + ((g832) & (!g2274) & (g1045)) + ((g832) & (g2274) & (g1045)));
	assign g1046 = (((!g34) & (!g36) & (!reset) & (g211) & (!g1045)) + ((!g34) & (!g36) & (!reset) & (g211) & (g1045)) + ((!g34) & (g36) & (!reset) & (!g211) & (g1045)) + ((!g34) & (g36) & (!reset) & (g211) & (g1045)) + ((g34) & (!g36) & (!reset) & (g211) & (!g1045)) + ((g34) & (!g36) & (!reset) & (g211) & (g1045)) + ((g34) & (g36) & (!reset) & (g211) & (!g1045)) + ((g34) & (g36) & (!reset) & (g211) & (g1045)));
	assign g7385 = (((!g832) & (g2276) & (!g1047)) + ((!g832) & (g2276) & (g1047)) + ((g832) & (!g2276) & (g1047)) + ((g832) & (g2276) & (g1047)));
	assign g1048 = (((!g34) & (!g36) & (!reset) & (g212) & (!g1047)) + ((!g34) & (!g36) & (!reset) & (g212) & (g1047)) + ((!g34) & (g36) & (!reset) & (!g212) & (g1047)) + ((!g34) & (g36) & (!reset) & (g212) & (g1047)) + ((g34) & (!g36) & (!reset) & (g212) & (!g1047)) + ((g34) & (!g36) & (!reset) & (g212) & (g1047)) + ((g34) & (g36) & (!reset) & (g212) & (!g1047)) + ((g34) & (g36) & (!reset) & (g212) & (g1047)));
	assign g7386 = (((!g832) & (g2278) & (!g1049)) + ((!g832) & (g2278) & (g1049)) + ((g832) & (!g2278) & (g1049)) + ((g832) & (g2278) & (g1049)));
	assign g1050 = (((!g34) & (!g36) & (!reset) & (g214) & (!g1049)) + ((!g34) & (!g36) & (!reset) & (g214) & (g1049)) + ((!g34) & (g36) & (!reset) & (!g214) & (g1049)) + ((!g34) & (g36) & (!reset) & (g214) & (g1049)) + ((g34) & (!g36) & (!reset) & (g214) & (!g1049)) + ((g34) & (!g36) & (!reset) & (g214) & (g1049)) + ((g34) & (g36) & (!reset) & (g214) & (!g1049)) + ((g34) & (g36) & (!reset) & (g214) & (g1049)));
	assign g7387 = (((!g832) & (g2280) & (!g1051)) + ((!g832) & (g2280) & (g1051)) + ((g832) & (!g2280) & (g1051)) + ((g832) & (g2280) & (g1051)));
	assign g1052 = (((!g34) & (!g36) & (!reset) & (g215) & (!g1051)) + ((!g34) & (!g36) & (!reset) & (g215) & (g1051)) + ((!g34) & (g36) & (!reset) & (!g215) & (g1051)) + ((!g34) & (g36) & (!reset) & (g215) & (g1051)) + ((g34) & (!g36) & (!reset) & (g215) & (!g1051)) + ((g34) & (!g36) & (!reset) & (g215) & (g1051)) + ((g34) & (g36) & (!reset) & (g215) & (!g1051)) + ((g34) & (g36) & (!reset) & (g215) & (g1051)));
	assign g7388 = (((!g832) & (g2282) & (!g1053)) + ((!g832) & (g2282) & (g1053)) + ((g832) & (!g2282) & (g1053)) + ((g832) & (g2282) & (g1053)));
	assign g1054 = (((!g34) & (!g36) & (!reset) & (g216) & (!g1053)) + ((!g34) & (!g36) & (!reset) & (g216) & (g1053)) + ((!g34) & (g36) & (!reset) & (!g216) & (g1053)) + ((!g34) & (g36) & (!reset) & (g216) & (g1053)) + ((g34) & (!g36) & (!reset) & (g216) & (!g1053)) + ((g34) & (!g36) & (!reset) & (g216) & (g1053)) + ((g34) & (g36) & (!reset) & (g216) & (!g1053)) + ((g34) & (g36) & (!reset) & (g216) & (g1053)));
	assign g7389 = (((!g832) & (g2284) & (!g1055)) + ((!g832) & (g2284) & (g1055)) + ((g832) & (!g2284) & (g1055)) + ((g832) & (g2284) & (g1055)));
	assign g1056 = (((!g34) & (!g36) & (!reset) & (g217) & (!g1055)) + ((!g34) & (!g36) & (!reset) & (g217) & (g1055)) + ((!g34) & (g36) & (!reset) & (!g217) & (g1055)) + ((!g34) & (g36) & (!reset) & (g217) & (g1055)) + ((g34) & (!g36) & (!reset) & (g217) & (!g1055)) + ((g34) & (!g36) & (!reset) & (g217) & (g1055)) + ((g34) & (g36) & (!reset) & (g217) & (!g1055)) + ((g34) & (g36) & (!reset) & (g217) & (g1055)));
	assign g7390 = (((!g832) & (g2285) & (!g1057)) + ((!g832) & (g2285) & (g1057)) + ((g832) & (!g2285) & (g1057)) + ((g832) & (g2285) & (g1057)));
	assign g1058 = (((!g34) & (!g36) & (!reset) & (g219) & (!g1057)) + ((!g34) & (!g36) & (!reset) & (g219) & (g1057)) + ((!g34) & (g36) & (!reset) & (!g219) & (g1057)) + ((!g34) & (g36) & (!reset) & (g219) & (g1057)) + ((g34) & (!g36) & (!reset) & (g219) & (!g1057)) + ((g34) & (!g36) & (!reset) & (g219) & (g1057)) + ((g34) & (g36) & (!reset) & (g219) & (!g1057)) + ((g34) & (g36) & (!reset) & (g219) & (g1057)));
	assign g7391 = (((!g832) & (g2287) & (!g1059)) + ((!g832) & (g2287) & (g1059)) + ((g832) & (!g2287) & (g1059)) + ((g832) & (g2287) & (g1059)));
	assign g1060 = (((!g34) & (!g36) & (!reset) & (g220) & (!g1059)) + ((!g34) & (!g36) & (!reset) & (g220) & (g1059)) + ((!g34) & (g36) & (!reset) & (!g220) & (g1059)) + ((!g34) & (g36) & (!reset) & (g220) & (g1059)) + ((g34) & (!g36) & (!reset) & (g220) & (!g1059)) + ((g34) & (!g36) & (!reset) & (g220) & (g1059)) + ((g34) & (g36) & (!reset) & (g220) & (!g1059)) + ((g34) & (g36) & (!reset) & (g220) & (g1059)));
	assign g7392 = (((!g832) & (g2289) & (!g1061)) + ((!g832) & (g2289) & (g1061)) + ((g832) & (!g2289) & (g1061)) + ((g832) & (g2289) & (g1061)));
	assign g1062 = (((!g34) & (!g36) & (!reset) & (g221) & (!g1061)) + ((!g34) & (!g36) & (!reset) & (g221) & (g1061)) + ((!g34) & (g36) & (!reset) & (!g221) & (g1061)) + ((!g34) & (g36) & (!reset) & (g221) & (g1061)) + ((g34) & (!g36) & (!reset) & (g221) & (!g1061)) + ((g34) & (!g36) & (!reset) & (g221) & (g1061)) + ((g34) & (g36) & (!reset) & (g221) & (!g1061)) + ((g34) & (g36) & (!reset) & (g221) & (g1061)));
	assign g7393 = (((!g832) & (g2291) & (!g1063)) + ((!g832) & (g2291) & (g1063)) + ((g832) & (!g2291) & (g1063)) + ((g832) & (g2291) & (g1063)));
	assign g1064 = (((!g34) & (!g36) & (!reset) & (g222) & (!g1063)) + ((!g34) & (!g36) & (!reset) & (g222) & (g1063)) + ((!g34) & (g36) & (!reset) & (!g222) & (g1063)) + ((!g34) & (g36) & (!reset) & (g222) & (g1063)) + ((g34) & (!g36) & (!reset) & (g222) & (!g1063)) + ((g34) & (!g36) & (!reset) & (g222) & (g1063)) + ((g34) & (g36) & (!reset) & (g222) & (!g1063)) + ((g34) & (g36) & (!reset) & (g222) & (g1063)));
	assign g7394 = (((!g2017) & (g2301) & (!g1065)) + ((!g2017) & (g2301) & (g1065)) + ((g2017) & (!g2301) & (g1065)) + ((g2017) & (g2301) & (g1065)));
	assign g1066 = (((!g827) & (!g202) & (!g225) & (!g1031) & (g1065) & (!g1032)) + ((!g827) & (!g202) & (!g225) & (!g1031) & (g1065) & (g1032)) + ((!g827) & (!g202) & (!g225) & (g1031) & (g1065) & (!g1032)) + ((!g827) & (!g202) & (!g225) & (g1031) & (g1065) & (g1032)) + ((!g827) & (!g202) & (g225) & (!g1031) & (g1065) & (!g1032)) + ((!g827) & (!g202) & (g225) & (!g1031) & (g1065) & (g1032)) + ((!g827) & (!g202) & (g225) & (g1031) & (g1065) & (!g1032)) + ((!g827) & (!g202) & (g225) & (g1031) & (g1065) & (g1032)) + ((!g827) & (g202) & (!g225) & (!g1031) & (g1065) & (!g1032)) + ((!g827) & (g202) & (!g225) & (!g1031) & (g1065) & (g1032)) + ((!g827) & (g202) & (!g225) & (g1031) & (g1065) & (!g1032)) + ((!g827) & (g202) & (!g225) & (g1031) & (g1065) & (g1032)) + ((!g827) & (g202) & (g225) & (!g1031) & (g1065) & (!g1032)) + ((!g827) & (g202) & (g225) & (!g1031) & (g1065) & (g1032)) + ((!g827) & (g202) & (g225) & (g1031) & (g1065) & (!g1032)) + ((!g827) & (g202) & (g225) & (g1031) & (g1065) & (g1032)) + ((g827) & (!g202) & (!g225) & (!g1031) & (g1065) & (!g1032)) + ((g827) & (!g202) & (!g225) & (!g1031) & (g1065) & (g1032)) + ((g827) & (!g202) & (!g225) & (g1031) & (!g1065) & (g1032)) + ((g827) & (!g202) & (!g225) & (g1031) & (g1065) & (!g1032)) + ((g827) & (!g202) & (g225) & (!g1031) & (!g1065) & (!g1032)) + ((g827) & (!g202) & (g225) & (!g1031) & (!g1065) & (g1032)) + ((g827) & (!g202) & (g225) & (g1031) & (!g1065) & (!g1032)) + ((g827) & (!g202) & (g225) & (g1031) & (g1065) & (g1032)) + ((g827) & (g202) & (!g225) & (!g1031) & (!g1065) & (g1032)) + ((g827) & (g202) & (!g225) & (!g1031) & (g1065) & (!g1032)) + ((g827) & (g202) & (!g225) & (g1031) & (!g1065) & (!g1032)) + ((g827) & (g202) & (!g225) & (g1031) & (!g1065) & (g1032)) + ((g827) & (g202) & (g225) & (!g1031) & (!g1065) & (!g1032)) + ((g827) & (g202) & (g225) & (!g1031) & (g1065) & (g1032)) + ((g827) & (g202) & (g225) & (g1031) & (g1065) & (!g1032)) + ((g827) & (g202) & (g225) & (g1031) & (g1065) & (g1032)));
	assign g1067 = (((!g34) & (!g36) & (!reset) & (g227) & (!g248)) + ((!g34) & (!g36) & (!reset) & (g227) & (g248)) + ((!g34) & (g36) & (!reset) & (!g227) & (g248)) + ((!g34) & (g36) & (!reset) & (g227) & (g248)) + ((g34) & (!g36) & (!reset) & (g227) & (!g248)) + ((g34) & (!g36) & (!reset) & (g227) & (g248)) + ((g34) & (g36) & (!reset) & (g227) & (!g248)) + ((g34) & (g36) & (!reset) & (g227) & (g248)));
	assign g7395 = (((!g832) & (g2303) & (!g1068)) + ((!g832) & (g2303) & (g1068)) + ((g832) & (!g2303) & (g1068)) + ((g832) & (g2303) & (g1068)));
	assign g1069 = (((!g34) & (!g36) & (!reset) & (g228) & (!g1068)) + ((!g34) & (!g36) & (!reset) & (g228) & (g1068)) + ((!g34) & (g36) & (!reset) & (!g228) & (g1068)) + ((!g34) & (g36) & (!reset) & (g228) & (g1068)) + ((g34) & (!g36) & (!reset) & (g228) & (!g1068)) + ((g34) & (!g36) & (!reset) & (g228) & (g1068)) + ((g34) & (g36) & (!reset) & (g228) & (!g1068)) + ((g34) & (g36) & (!reset) & (g228) & (g1068)));
	assign g7396 = (((!g832) & (g2306) & (!g1070)) + ((!g832) & (g2306) & (g1070)) + ((g832) & (!g2306) & (g1070)) + ((g832) & (g2306) & (g1070)));
	assign g1071 = (((!g34) & (!g36) & (!reset) & (g229) & (!g1070)) + ((!g34) & (!g36) & (!reset) & (g229) & (g1070)) + ((!g34) & (g36) & (!reset) & (!g229) & (g1070)) + ((!g34) & (g36) & (!reset) & (g229) & (g1070)) + ((g34) & (!g36) & (!reset) & (g229) & (!g1070)) + ((g34) & (!g36) & (!reset) & (g229) & (g1070)) + ((g34) & (g36) & (!reset) & (g229) & (!g1070)) + ((g34) & (g36) & (!reset) & (g229) & (g1070)));
	assign g7397 = (((!g832) & (g2308) & (!g1072)) + ((!g832) & (g2308) & (g1072)) + ((g832) & (!g2308) & (g1072)) + ((g832) & (g2308) & (g1072)));
	assign g1073 = (((!g34) & (!g36) & (!reset) & (g230) & (!g1072)) + ((!g34) & (!g36) & (!reset) & (g230) & (g1072)) + ((!g34) & (g36) & (!reset) & (!g230) & (g1072)) + ((!g34) & (g36) & (!reset) & (g230) & (g1072)) + ((g34) & (!g36) & (!reset) & (g230) & (!g1072)) + ((g34) & (!g36) & (!reset) & (g230) & (g1072)) + ((g34) & (g36) & (!reset) & (g230) & (!g1072)) + ((g34) & (g36) & (!reset) & (g230) & (g1072)));
	assign g7398 = (((!g832) & (g2310) & (!g1074)) + ((!g832) & (g2310) & (g1074)) + ((g832) & (!g2310) & (g1074)) + ((g832) & (g2310) & (g1074)));
	assign g1075 = (((!g34) & (!g36) & (!reset) & (g232) & (!g1074)) + ((!g34) & (!g36) & (!reset) & (g232) & (g1074)) + ((!g34) & (g36) & (!reset) & (!g232) & (g1074)) + ((!g34) & (g36) & (!reset) & (g232) & (g1074)) + ((g34) & (!g36) & (!reset) & (g232) & (!g1074)) + ((g34) & (!g36) & (!reset) & (g232) & (g1074)) + ((g34) & (g36) & (!reset) & (g232) & (!g1074)) + ((g34) & (g36) & (!reset) & (g232) & (g1074)));
	assign g7399 = (((!g832) & (g2313) & (!g1076)) + ((!g832) & (g2313) & (g1076)) + ((g832) & (!g2313) & (g1076)) + ((g832) & (g2313) & (g1076)));
	assign g1077 = (((!g34) & (!g36) & (!reset) & (g233) & (!g1076)) + ((!g34) & (!g36) & (!reset) & (g233) & (g1076)) + ((!g34) & (g36) & (!reset) & (!g233) & (g1076)) + ((!g34) & (g36) & (!reset) & (g233) & (g1076)) + ((g34) & (!g36) & (!reset) & (g233) & (!g1076)) + ((g34) & (!g36) & (!reset) & (g233) & (g1076)) + ((g34) & (g36) & (!reset) & (g233) & (!g1076)) + ((g34) & (g36) & (!reset) & (g233) & (g1076)));
	assign g7400 = (((!g832) & (g2316) & (!g1078)) + ((!g832) & (g2316) & (g1078)) + ((g832) & (!g2316) & (g1078)) + ((g832) & (g2316) & (g1078)));
	assign g1079 = (((!g34) & (!g36) & (!reset) & (g234) & (!g1078)) + ((!g34) & (!g36) & (!reset) & (g234) & (g1078)) + ((!g34) & (g36) & (!reset) & (!g234) & (g1078)) + ((!g34) & (g36) & (!reset) & (g234) & (g1078)) + ((g34) & (!g36) & (!reset) & (g234) & (!g1078)) + ((g34) & (!g36) & (!reset) & (g234) & (g1078)) + ((g34) & (g36) & (!reset) & (g234) & (!g1078)) + ((g34) & (g36) & (!reset) & (g234) & (g1078)));
	assign g7401 = (((!g832) & (g2319) & (!g1080)) + ((!g832) & (g2319) & (g1080)) + ((g832) & (!g2319) & (g1080)) + ((g832) & (g2319) & (g1080)));
	assign g1081 = (((!g34) & (!g36) & (!reset) & (g235) & (!g1080)) + ((!g34) & (!g36) & (!reset) & (g235) & (g1080)) + ((!g34) & (g36) & (!reset) & (!g235) & (g1080)) + ((!g34) & (g36) & (!reset) & (g235) & (g1080)) + ((g34) & (!g36) & (!reset) & (g235) & (!g1080)) + ((g34) & (!g36) & (!reset) & (g235) & (g1080)) + ((g34) & (g36) & (!reset) & (g235) & (!g1080)) + ((g34) & (g36) & (!reset) & (g235) & (g1080)));
	assign g7402 = (((!g832) & (g2322) & (!g1082)) + ((!g832) & (g2322) & (g1082)) + ((g832) & (!g2322) & (g1082)) + ((g832) & (g2322) & (g1082)));
	assign g1083 = (((!g34) & (!g36) & (!reset) & (g237) & (!g1082)) + ((!g34) & (!g36) & (!reset) & (g237) & (g1082)) + ((!g34) & (g36) & (!reset) & (!g237) & (g1082)) + ((!g34) & (g36) & (!reset) & (g237) & (g1082)) + ((g34) & (!g36) & (!reset) & (g237) & (!g1082)) + ((g34) & (!g36) & (!reset) & (g237) & (g1082)) + ((g34) & (g36) & (!reset) & (g237) & (!g1082)) + ((g34) & (g36) & (!reset) & (g237) & (g1082)));
	assign g7403 = (((!g832) & (g2325) & (!g1084)) + ((!g832) & (g2325) & (g1084)) + ((g832) & (!g2325) & (g1084)) + ((g832) & (g2325) & (g1084)));
	assign g1085 = (((!g34) & (!g36) & (!reset) & (g238) & (!g1084)) + ((!g34) & (!g36) & (!reset) & (g238) & (g1084)) + ((!g34) & (g36) & (!reset) & (!g238) & (g1084)) + ((!g34) & (g36) & (!reset) & (g238) & (g1084)) + ((g34) & (!g36) & (!reset) & (g238) & (!g1084)) + ((g34) & (!g36) & (!reset) & (g238) & (g1084)) + ((g34) & (g36) & (!reset) & (g238) & (!g1084)) + ((g34) & (g36) & (!reset) & (g238) & (g1084)));
	assign g7404 = (((!g832) & (g2328) & (!g1086)) + ((!g832) & (g2328) & (g1086)) + ((g832) & (!g2328) & (g1086)) + ((g832) & (g2328) & (g1086)));
	assign g1087 = (((!g34) & (!g36) & (!reset) & (g239) & (!g1086)) + ((!g34) & (!g36) & (!reset) & (g239) & (g1086)) + ((!g34) & (g36) & (!reset) & (!g239) & (g1086)) + ((!g34) & (g36) & (!reset) & (g239) & (g1086)) + ((g34) & (!g36) & (!reset) & (g239) & (!g1086)) + ((g34) & (!g36) & (!reset) & (g239) & (g1086)) + ((g34) & (g36) & (!reset) & (g239) & (!g1086)) + ((g34) & (g36) & (!reset) & (g239) & (g1086)));
	assign g7405 = (((!g832) & (g2331) & (!g1088)) + ((!g832) & (g2331) & (g1088)) + ((g832) & (!g2331) & (g1088)) + ((g832) & (g2331) & (g1088)));
	assign g1089 = (((!g34) & (!g36) & (!reset) & (g240) & (!g1088)) + ((!g34) & (!g36) & (!reset) & (g240) & (g1088)) + ((!g34) & (g36) & (!reset) & (!g240) & (g1088)) + ((!g34) & (g36) & (!reset) & (g240) & (g1088)) + ((g34) & (!g36) & (!reset) & (g240) & (!g1088)) + ((g34) & (!g36) & (!reset) & (g240) & (g1088)) + ((g34) & (g36) & (!reset) & (g240) & (!g1088)) + ((g34) & (g36) & (!reset) & (g240) & (g1088)));
	assign g7406 = (((!g832) & (g2333) & (!g1090)) + ((!g832) & (g2333) & (g1090)) + ((g832) & (!g2333) & (g1090)) + ((g832) & (g2333) & (g1090)));
	assign g1091 = (((!g34) & (!g36) & (!reset) & (g242) & (!g1090)) + ((!g34) & (!g36) & (!reset) & (g242) & (g1090)) + ((!g34) & (g36) & (!reset) & (!g242) & (g1090)) + ((!g34) & (g36) & (!reset) & (g242) & (g1090)) + ((g34) & (!g36) & (!reset) & (g242) & (!g1090)) + ((g34) & (!g36) & (!reset) & (g242) & (g1090)) + ((g34) & (g36) & (!reset) & (g242) & (!g1090)) + ((g34) & (g36) & (!reset) & (g242) & (g1090)));
	assign g7407 = (((!g832) & (g2336) & (!g1092)) + ((!g832) & (g2336) & (g1092)) + ((g832) & (!g2336) & (g1092)) + ((g832) & (g2336) & (g1092)));
	assign g1093 = (((!g34) & (!g36) & (!reset) & (g243) & (!g1092)) + ((!g34) & (!g36) & (!reset) & (g243) & (g1092)) + ((!g34) & (g36) & (!reset) & (!g243) & (g1092)) + ((!g34) & (g36) & (!reset) & (g243) & (g1092)) + ((g34) & (!g36) & (!reset) & (g243) & (!g1092)) + ((g34) & (!g36) & (!reset) & (g243) & (g1092)) + ((g34) & (g36) & (!reset) & (g243) & (!g1092)) + ((g34) & (g36) & (!reset) & (g243) & (g1092)));
	assign g7408 = (((!g832) & (g2339) & (!g1094)) + ((!g832) & (g2339) & (g1094)) + ((g832) & (!g2339) & (g1094)) + ((g832) & (g2339) & (g1094)));
	assign g1095 = (((!g34) & (!g36) & (!reset) & (g244) & (!g1094)) + ((!g34) & (!g36) & (!reset) & (g244) & (g1094)) + ((!g34) & (g36) & (!reset) & (!g244) & (g1094)) + ((!g34) & (g36) & (!reset) & (g244) & (g1094)) + ((g34) & (!g36) & (!reset) & (g244) & (!g1094)) + ((g34) & (!g36) & (!reset) & (g244) & (g1094)) + ((g34) & (g36) & (!reset) & (g244) & (!g1094)) + ((g34) & (g36) & (!reset) & (g244) & (g1094)));
	assign g7409 = (((!g832) & (g2342) & (!g1096)) + ((!g832) & (g2342) & (g1096)) + ((g832) & (!g2342) & (g1096)) + ((g832) & (g2342) & (g1096)));
	assign g1097 = (((!g34) & (!g36) & (!reset) & (g245) & (!g1096)) + ((!g34) & (!g36) & (!reset) & (g245) & (g1096)) + ((!g34) & (g36) & (!reset) & (!g245) & (g1096)) + ((!g34) & (g36) & (!reset) & (g245) & (g1096)) + ((g34) & (!g36) & (!reset) & (g245) & (!g1096)) + ((g34) & (!g36) & (!reset) & (g245) & (g1096)) + ((g34) & (g36) & (!reset) & (g245) & (!g1096)) + ((g34) & (g36) & (!reset) & (g245) & (g1096)));
	assign g7410 = (((!g2017) & (g7152) & (!g1098)) + ((!g2017) & (g7152) & (g1098)) + ((g2017) & (!g7152) & (g1098)) + ((g2017) & (g7152) & (g1098)));
	assign g1099 = (((!g202) & (!g225) & (g1031) & (g1065) & (g1032)) + ((!g202) & (g225) & (!g1031) & (g1065) & (!g1032)) + ((!g202) & (g225) & (!g1031) & (g1065) & (g1032)) + ((!g202) & (g225) & (g1031) & (!g1065) & (g1032)) + ((!g202) & (g225) & (g1031) & (g1065) & (!g1032)) + ((!g202) & (g225) & (g1031) & (g1065) & (g1032)) + ((g202) & (!g225) & (!g1031) & (g1065) & (g1032)) + ((g202) & (!g225) & (g1031) & (g1065) & (!g1032)) + ((g202) & (!g225) & (g1031) & (g1065) & (g1032)) + ((g202) & (g225) & (!g1031) & (!g1065) & (g1032)) + ((g202) & (g225) & (!g1031) & (g1065) & (!g1032)) + ((g202) & (g225) & (!g1031) & (g1065) & (g1032)) + ((g202) & (g225) & (g1031) & (!g1065) & (!g1032)) + ((g202) & (g225) & (g1031) & (!g1065) & (g1032)) + ((g202) & (g225) & (g1031) & (g1065) & (!g1032)) + ((g202) & (g225) & (g1031) & (g1065) & (g1032)));
	assign g1100 = (((!g827) & (!g248) & (g1098) & (!g1099)) + ((!g827) & (!g248) & (g1098) & (g1099)) + ((!g827) & (g248) & (g1098) & (!g1099)) + ((!g827) & (g248) & (g1098) & (g1099)) + ((g827) & (!g248) & (!g1098) & (g1099)) + ((g827) & (!g248) & (g1098) & (!g1099)) + ((g827) & (g248) & (!g1098) & (!g1099)) + ((g827) & (g248) & (g1098) & (g1099)));
	assign g1101 = (((!g34) & (!g36) & (!reset) & (g250) & (!g271)) + ((!g34) & (!g36) & (!reset) & (g250) & (g271)) + ((!g34) & (g36) & (!reset) & (!g250) & (g271)) + ((!g34) & (g36) & (!reset) & (g250) & (g271)) + ((g34) & (!g36) & (!reset) & (g250) & (!g271)) + ((g34) & (!g36) & (!reset) & (g250) & (g271)) + ((g34) & (g36) & (!reset) & (g250) & (!g271)) + ((g34) & (g36) & (!reset) & (g250) & (g271)));
	assign g7411 = (((!g832) & (g2349) & (!g1102)) + ((!g832) & (g2349) & (g1102)) + ((g832) & (!g2349) & (g1102)) + ((g832) & (g2349) & (g1102)));
	assign g1103 = (((!g34) & (!g36) & (!reset) & (g251) & (!g1102)) + ((!g34) & (!g36) & (!reset) & (g251) & (g1102)) + ((!g34) & (g36) & (!reset) & (!g251) & (g1102)) + ((!g34) & (g36) & (!reset) & (g251) & (g1102)) + ((g34) & (!g36) & (!reset) & (g251) & (!g1102)) + ((g34) & (!g36) & (!reset) & (g251) & (g1102)) + ((g34) & (g36) & (!reset) & (g251) & (!g1102)) + ((g34) & (g36) & (!reset) & (g251) & (g1102)));
	assign g7412 = (((!g832) & (g2351) & (!g1104)) + ((!g832) & (g2351) & (g1104)) + ((g832) & (!g2351) & (g1104)) + ((g832) & (g2351) & (g1104)));
	assign g1105 = (((!g34) & (!g36) & (!reset) & (g252) & (!g1104)) + ((!g34) & (!g36) & (!reset) & (g252) & (g1104)) + ((!g34) & (g36) & (!reset) & (!g252) & (g1104)) + ((!g34) & (g36) & (!reset) & (g252) & (g1104)) + ((g34) & (!g36) & (!reset) & (g252) & (!g1104)) + ((g34) & (!g36) & (!reset) & (g252) & (g1104)) + ((g34) & (g36) & (!reset) & (g252) & (!g1104)) + ((g34) & (g36) & (!reset) & (g252) & (g1104)));
	assign g7413 = (((!g832) & (g2352) & (!g1106)) + ((!g832) & (g2352) & (g1106)) + ((g832) & (!g2352) & (g1106)) + ((g832) & (g2352) & (g1106)));
	assign g1107 = (((!g34) & (!g36) & (!reset) & (g253) & (!g1106)) + ((!g34) & (!g36) & (!reset) & (g253) & (g1106)) + ((!g34) & (g36) & (!reset) & (!g253) & (g1106)) + ((!g34) & (g36) & (!reset) & (g253) & (g1106)) + ((g34) & (!g36) & (!reset) & (g253) & (!g1106)) + ((g34) & (!g36) & (!reset) & (g253) & (g1106)) + ((g34) & (g36) & (!reset) & (g253) & (!g1106)) + ((g34) & (g36) & (!reset) & (g253) & (g1106)));
	assign g7414 = (((!g832) & (g2353) & (!g1108)) + ((!g832) & (g2353) & (g1108)) + ((g832) & (!g2353) & (g1108)) + ((g832) & (g2353) & (g1108)));
	assign g1109 = (((!g34) & (!g36) & (!reset) & (g255) & (!g1108)) + ((!g34) & (!g36) & (!reset) & (g255) & (g1108)) + ((!g34) & (g36) & (!reset) & (!g255) & (g1108)) + ((!g34) & (g36) & (!reset) & (g255) & (g1108)) + ((g34) & (!g36) & (!reset) & (g255) & (!g1108)) + ((g34) & (!g36) & (!reset) & (g255) & (g1108)) + ((g34) & (g36) & (!reset) & (g255) & (!g1108)) + ((g34) & (g36) & (!reset) & (g255) & (g1108)));
	assign g7415 = (((!g832) & (g2355) & (!g1110)) + ((!g832) & (g2355) & (g1110)) + ((g832) & (!g2355) & (g1110)) + ((g832) & (g2355) & (g1110)));
	assign g1111 = (((!g34) & (!g36) & (!reset) & (g256) & (!g1110)) + ((!g34) & (!g36) & (!reset) & (g256) & (g1110)) + ((!g34) & (g36) & (!reset) & (!g256) & (g1110)) + ((!g34) & (g36) & (!reset) & (g256) & (g1110)) + ((g34) & (!g36) & (!reset) & (g256) & (!g1110)) + ((g34) & (!g36) & (!reset) & (g256) & (g1110)) + ((g34) & (g36) & (!reset) & (g256) & (!g1110)) + ((g34) & (g36) & (!reset) & (g256) & (g1110)));
	assign g7416 = (((!g832) & (g2357) & (!g1112)) + ((!g832) & (g2357) & (g1112)) + ((g832) & (!g2357) & (g1112)) + ((g832) & (g2357) & (g1112)));
	assign g1113 = (((!g34) & (!g36) & (!reset) & (g257) & (!g1112)) + ((!g34) & (!g36) & (!reset) & (g257) & (g1112)) + ((!g34) & (g36) & (!reset) & (!g257) & (g1112)) + ((!g34) & (g36) & (!reset) & (g257) & (g1112)) + ((g34) & (!g36) & (!reset) & (g257) & (!g1112)) + ((g34) & (!g36) & (!reset) & (g257) & (g1112)) + ((g34) & (g36) & (!reset) & (g257) & (!g1112)) + ((g34) & (g36) & (!reset) & (g257) & (g1112)));
	assign g7417 = (((!g832) & (g2359) & (!g1114)) + ((!g832) & (g2359) & (g1114)) + ((g832) & (!g2359) & (g1114)) + ((g832) & (g2359) & (g1114)));
	assign g1115 = (((!g34) & (!g36) & (!reset) & (g258) & (!g1114)) + ((!g34) & (!g36) & (!reset) & (g258) & (g1114)) + ((!g34) & (g36) & (!reset) & (!g258) & (g1114)) + ((!g34) & (g36) & (!reset) & (g258) & (g1114)) + ((g34) & (!g36) & (!reset) & (g258) & (!g1114)) + ((g34) & (!g36) & (!reset) & (g258) & (g1114)) + ((g34) & (g36) & (!reset) & (g258) & (!g1114)) + ((g34) & (g36) & (!reset) & (g258) & (g1114)));
	assign g7418 = (((!g832) & (g2361) & (!g1116)) + ((!g832) & (g2361) & (g1116)) + ((g832) & (!g2361) & (g1116)) + ((g832) & (g2361) & (g1116)));
	assign g1117 = (((!g34) & (!g36) & (!reset) & (g260) & (!g1116)) + ((!g34) & (!g36) & (!reset) & (g260) & (g1116)) + ((!g34) & (g36) & (!reset) & (!g260) & (g1116)) + ((!g34) & (g36) & (!reset) & (g260) & (g1116)) + ((g34) & (!g36) & (!reset) & (g260) & (!g1116)) + ((g34) & (!g36) & (!reset) & (g260) & (g1116)) + ((g34) & (g36) & (!reset) & (g260) & (!g1116)) + ((g34) & (g36) & (!reset) & (g260) & (g1116)));
	assign g7419 = (((!g832) & (g2363) & (!g1118)) + ((!g832) & (g2363) & (g1118)) + ((g832) & (!g2363) & (g1118)) + ((g832) & (g2363) & (g1118)));
	assign g1119 = (((!g34) & (!g36) & (!reset) & (g261) & (!g1118)) + ((!g34) & (!g36) & (!reset) & (g261) & (g1118)) + ((!g34) & (g36) & (!reset) & (!g261) & (g1118)) + ((!g34) & (g36) & (!reset) & (g261) & (g1118)) + ((g34) & (!g36) & (!reset) & (g261) & (!g1118)) + ((g34) & (!g36) & (!reset) & (g261) & (g1118)) + ((g34) & (g36) & (!reset) & (g261) & (!g1118)) + ((g34) & (g36) & (!reset) & (g261) & (g1118)));
	assign g7420 = (((!g832) & (g2365) & (!g1120)) + ((!g832) & (g2365) & (g1120)) + ((g832) & (!g2365) & (g1120)) + ((g832) & (g2365) & (g1120)));
	assign g1121 = (((!g34) & (!g36) & (!reset) & (g262) & (!g1120)) + ((!g34) & (!g36) & (!reset) & (g262) & (g1120)) + ((!g34) & (g36) & (!reset) & (!g262) & (g1120)) + ((!g34) & (g36) & (!reset) & (g262) & (g1120)) + ((g34) & (!g36) & (!reset) & (g262) & (!g1120)) + ((g34) & (!g36) & (!reset) & (g262) & (g1120)) + ((g34) & (g36) & (!reset) & (g262) & (!g1120)) + ((g34) & (g36) & (!reset) & (g262) & (g1120)));
	assign g7421 = (((!g832) & (g2367) & (!g1122)) + ((!g832) & (g2367) & (g1122)) + ((g832) & (!g2367) & (g1122)) + ((g832) & (g2367) & (g1122)));
	assign g1123 = (((!g34) & (!g36) & (!reset) & (g263) & (!g1122)) + ((!g34) & (!g36) & (!reset) & (g263) & (g1122)) + ((!g34) & (g36) & (!reset) & (!g263) & (g1122)) + ((!g34) & (g36) & (!reset) & (g263) & (g1122)) + ((g34) & (!g36) & (!reset) & (g263) & (!g1122)) + ((g34) & (!g36) & (!reset) & (g263) & (g1122)) + ((g34) & (g36) & (!reset) & (g263) & (!g1122)) + ((g34) & (g36) & (!reset) & (g263) & (g1122)));
	assign g7422 = (((!g832) & (g2368) & (!g1124)) + ((!g832) & (g2368) & (g1124)) + ((g832) & (!g2368) & (g1124)) + ((g832) & (g2368) & (g1124)));
	assign g1125 = (((!g34) & (!g36) & (!reset) & (g265) & (!g1124)) + ((!g34) & (!g36) & (!reset) & (g265) & (g1124)) + ((!g34) & (g36) & (!reset) & (!g265) & (g1124)) + ((!g34) & (g36) & (!reset) & (g265) & (g1124)) + ((g34) & (!g36) & (!reset) & (g265) & (!g1124)) + ((g34) & (!g36) & (!reset) & (g265) & (g1124)) + ((g34) & (g36) & (!reset) & (g265) & (!g1124)) + ((g34) & (g36) & (!reset) & (g265) & (g1124)));
	assign g7423 = (((!g832) & (g2370) & (!g1126)) + ((!g832) & (g2370) & (g1126)) + ((g832) & (!g2370) & (g1126)) + ((g832) & (g2370) & (g1126)));
	assign g1127 = (((!g34) & (!g36) & (!reset) & (g266) & (!g1126)) + ((!g34) & (!g36) & (!reset) & (g266) & (g1126)) + ((!g34) & (g36) & (!reset) & (!g266) & (g1126)) + ((!g34) & (g36) & (!reset) & (g266) & (g1126)) + ((g34) & (!g36) & (!reset) & (g266) & (!g1126)) + ((g34) & (!g36) & (!reset) & (g266) & (g1126)) + ((g34) & (g36) & (!reset) & (g266) & (!g1126)) + ((g34) & (g36) & (!reset) & (g266) & (g1126)));
	assign g7424 = (((!g832) & (g2372) & (!g1128)) + ((!g832) & (g2372) & (g1128)) + ((g832) & (!g2372) & (g1128)) + ((g832) & (g2372) & (g1128)));
	assign g1129 = (((!g34) & (!g36) & (!reset) & (g267) & (!g1128)) + ((!g34) & (!g36) & (!reset) & (g267) & (g1128)) + ((!g34) & (g36) & (!reset) & (!g267) & (g1128)) + ((!g34) & (g36) & (!reset) & (g267) & (g1128)) + ((g34) & (!g36) & (!reset) & (g267) & (!g1128)) + ((g34) & (!g36) & (!reset) & (g267) & (g1128)) + ((g34) & (g36) & (!reset) & (g267) & (!g1128)) + ((g34) & (g36) & (!reset) & (g267) & (g1128)));
	assign g7425 = (((!g832) & (g2374) & (!g1130)) + ((!g832) & (g2374) & (g1130)) + ((g832) & (!g2374) & (g1130)) + ((g832) & (g2374) & (g1130)));
	assign g1131 = (((!g34) & (!g36) & (!reset) & (g268) & (!g1130)) + ((!g34) & (!g36) & (!reset) & (g268) & (g1130)) + ((!g34) & (g36) & (!reset) & (!g268) & (g1130)) + ((!g34) & (g36) & (!reset) & (g268) & (g1130)) + ((g34) & (!g36) & (!reset) & (g268) & (!g1130)) + ((g34) & (!g36) & (!reset) & (g268) & (g1130)) + ((g34) & (g36) & (!reset) & (g268) & (!g1130)) + ((g34) & (g36) & (!reset) & (g268) & (g1130)));
	assign g7426 = (((!g2017) & (g7146) & (!g1132)) + ((!g2017) & (g7146) & (g1132)) + ((g2017) & (!g7146) & (g1132)) + ((g2017) & (g7146) & (g1132)));
	assign g1133 = (((!g827) & (!g248) & (!g271) & (!g1098) & (g1132) & (!g1099)) + ((!g827) & (!g248) & (!g271) & (!g1098) & (g1132) & (g1099)) + ((!g827) & (!g248) & (!g271) & (g1098) & (g1132) & (!g1099)) + ((!g827) & (!g248) & (!g271) & (g1098) & (g1132) & (g1099)) + ((!g827) & (!g248) & (g271) & (!g1098) & (g1132) & (!g1099)) + ((!g827) & (!g248) & (g271) & (!g1098) & (g1132) & (g1099)) + ((!g827) & (!g248) & (g271) & (g1098) & (g1132) & (!g1099)) + ((!g827) & (!g248) & (g271) & (g1098) & (g1132) & (g1099)) + ((!g827) & (g248) & (!g271) & (!g1098) & (g1132) & (!g1099)) + ((!g827) & (g248) & (!g271) & (!g1098) & (g1132) & (g1099)) + ((!g827) & (g248) & (!g271) & (g1098) & (g1132) & (!g1099)) + ((!g827) & (g248) & (!g271) & (g1098) & (g1132) & (g1099)) + ((!g827) & (g248) & (g271) & (!g1098) & (g1132) & (!g1099)) + ((!g827) & (g248) & (g271) & (!g1098) & (g1132) & (g1099)) + ((!g827) & (g248) & (g271) & (g1098) & (g1132) & (!g1099)) + ((!g827) & (g248) & (g271) & (g1098) & (g1132) & (g1099)) + ((g827) & (!g248) & (!g271) & (!g1098) & (g1132) & (!g1099)) + ((g827) & (!g248) & (!g271) & (!g1098) & (g1132) & (g1099)) + ((g827) & (!g248) & (!g271) & (g1098) & (!g1132) & (g1099)) + ((g827) & (!g248) & (!g271) & (g1098) & (g1132) & (!g1099)) + ((g827) & (!g248) & (g271) & (!g1098) & (!g1132) & (!g1099)) + ((g827) & (!g248) & (g271) & (!g1098) & (!g1132) & (g1099)) + ((g827) & (!g248) & (g271) & (g1098) & (!g1132) & (!g1099)) + ((g827) & (!g248) & (g271) & (g1098) & (g1132) & (g1099)) + ((g827) & (g248) & (!g271) & (!g1098) & (!g1132) & (g1099)) + ((g827) & (g248) & (!g271) & (!g1098) & (g1132) & (!g1099)) + ((g827) & (g248) & (!g271) & (g1098) & (!g1132) & (!g1099)) + ((g827) & (g248) & (!g271) & (g1098) & (!g1132) & (g1099)) + ((g827) & (g248) & (g271) & (!g1098) & (!g1132) & (!g1099)) + ((g827) & (g248) & (g271) & (!g1098) & (g1132) & (g1099)) + ((g827) & (g248) & (g271) & (g1098) & (g1132) & (!g1099)) + ((g827) & (g248) & (g271) & (g1098) & (g1132) & (g1099)));
	assign g1134 = (((!g34) & (!g36) & (!reset) & (g273) & (!g294)) + ((!g34) & (!g36) & (!reset) & (g273) & (g294)) + ((!g34) & (g36) & (!reset) & (!g273) & (g294)) + ((!g34) & (g36) & (!reset) & (g273) & (g294)) + ((g34) & (!g36) & (!reset) & (g273) & (!g294)) + ((g34) & (!g36) & (!reset) & (g273) & (g294)) + ((g34) & (g36) & (!reset) & (g273) & (!g294)) + ((g34) & (g36) & (!reset) & (g273) & (g294)));
	assign g7427 = (((!g832) & (g2382) & (!g1135)) + ((!g832) & (g2382) & (g1135)) + ((g832) & (!g2382) & (g1135)) + ((g832) & (g2382) & (g1135)));
	assign g1136 = (((!g34) & (!g36) & (!reset) & (g274) & (!g1135)) + ((!g34) & (!g36) & (!reset) & (g274) & (g1135)) + ((!g34) & (g36) & (!reset) & (!g274) & (g1135)) + ((!g34) & (g36) & (!reset) & (g274) & (g1135)) + ((g34) & (!g36) & (!reset) & (g274) & (!g1135)) + ((g34) & (!g36) & (!reset) & (g274) & (g1135)) + ((g34) & (g36) & (!reset) & (g274) & (!g1135)) + ((g34) & (g36) & (!reset) & (g274) & (g1135)));
	assign g7428 = (((!g832) & (g2385) & (!g1137)) + ((!g832) & (g2385) & (g1137)) + ((g832) & (!g2385) & (g1137)) + ((g832) & (g2385) & (g1137)));
	assign g1138 = (((!g34) & (!g36) & (!reset) & (g275) & (!g1137)) + ((!g34) & (!g36) & (!reset) & (g275) & (g1137)) + ((!g34) & (g36) & (!reset) & (!g275) & (g1137)) + ((!g34) & (g36) & (!reset) & (g275) & (g1137)) + ((g34) & (!g36) & (!reset) & (g275) & (!g1137)) + ((g34) & (!g36) & (!reset) & (g275) & (g1137)) + ((g34) & (g36) & (!reset) & (g275) & (!g1137)) + ((g34) & (g36) & (!reset) & (g275) & (g1137)));
	assign g7429 = (((!g832) & (g2387) & (!g1139)) + ((!g832) & (g2387) & (g1139)) + ((g832) & (!g2387) & (g1139)) + ((g832) & (g2387) & (g1139)));
	assign g1140 = (((!g34) & (!g36) & (!reset) & (g276) & (!g1139)) + ((!g34) & (!g36) & (!reset) & (g276) & (g1139)) + ((!g34) & (g36) & (!reset) & (!g276) & (g1139)) + ((!g34) & (g36) & (!reset) & (g276) & (g1139)) + ((g34) & (!g36) & (!reset) & (g276) & (!g1139)) + ((g34) & (!g36) & (!reset) & (g276) & (g1139)) + ((g34) & (g36) & (!reset) & (g276) & (!g1139)) + ((g34) & (g36) & (!reset) & (g276) & (g1139)));
	assign g7430 = (((!g832) & (g2389) & (!g1141)) + ((!g832) & (g2389) & (g1141)) + ((g832) & (!g2389) & (g1141)) + ((g832) & (g2389) & (g1141)));
	assign g1142 = (((!g34) & (!g36) & (!reset) & (g278) & (!g1141)) + ((!g34) & (!g36) & (!reset) & (g278) & (g1141)) + ((!g34) & (g36) & (!reset) & (!g278) & (g1141)) + ((!g34) & (g36) & (!reset) & (g278) & (g1141)) + ((g34) & (!g36) & (!reset) & (g278) & (!g1141)) + ((g34) & (!g36) & (!reset) & (g278) & (g1141)) + ((g34) & (g36) & (!reset) & (g278) & (!g1141)) + ((g34) & (g36) & (!reset) & (g278) & (g1141)));
	assign g7431 = (((!g832) & (g2392) & (!g1143)) + ((!g832) & (g2392) & (g1143)) + ((g832) & (!g2392) & (g1143)) + ((g832) & (g2392) & (g1143)));
	assign g1144 = (((!g34) & (!g36) & (!reset) & (g279) & (!g1143)) + ((!g34) & (!g36) & (!reset) & (g279) & (g1143)) + ((!g34) & (g36) & (!reset) & (!g279) & (g1143)) + ((!g34) & (g36) & (!reset) & (g279) & (g1143)) + ((g34) & (!g36) & (!reset) & (g279) & (!g1143)) + ((g34) & (!g36) & (!reset) & (g279) & (g1143)) + ((g34) & (g36) & (!reset) & (g279) & (!g1143)) + ((g34) & (g36) & (!reset) & (g279) & (g1143)));
	assign g7432 = (((!g832) & (g2395) & (!g1145)) + ((!g832) & (g2395) & (g1145)) + ((g832) & (!g2395) & (g1145)) + ((g832) & (g2395) & (g1145)));
	assign g1146 = (((!g34) & (!g36) & (!reset) & (g280) & (!g1145)) + ((!g34) & (!g36) & (!reset) & (g280) & (g1145)) + ((!g34) & (g36) & (!reset) & (!g280) & (g1145)) + ((!g34) & (g36) & (!reset) & (g280) & (g1145)) + ((g34) & (!g36) & (!reset) & (g280) & (!g1145)) + ((g34) & (!g36) & (!reset) & (g280) & (g1145)) + ((g34) & (g36) & (!reset) & (g280) & (!g1145)) + ((g34) & (g36) & (!reset) & (g280) & (g1145)));
	assign g7433 = (((!g832) & (g2398) & (!g1147)) + ((!g832) & (g2398) & (g1147)) + ((g832) & (!g2398) & (g1147)) + ((g832) & (g2398) & (g1147)));
	assign g1148 = (((!g34) & (!g36) & (!reset) & (g281) & (!g1147)) + ((!g34) & (!g36) & (!reset) & (g281) & (g1147)) + ((!g34) & (g36) & (!reset) & (!g281) & (g1147)) + ((!g34) & (g36) & (!reset) & (g281) & (g1147)) + ((g34) & (!g36) & (!reset) & (g281) & (!g1147)) + ((g34) & (!g36) & (!reset) & (g281) & (g1147)) + ((g34) & (g36) & (!reset) & (g281) & (!g1147)) + ((g34) & (g36) & (!reset) & (g281) & (g1147)));
	assign g7434 = (((!g832) & (g2401) & (!g1149)) + ((!g832) & (g2401) & (g1149)) + ((g832) & (!g2401) & (g1149)) + ((g832) & (g2401) & (g1149)));
	assign g1150 = (((!g34) & (!g36) & (!reset) & (g283) & (!g1149)) + ((!g34) & (!g36) & (!reset) & (g283) & (g1149)) + ((!g34) & (g36) & (!reset) & (!g283) & (g1149)) + ((!g34) & (g36) & (!reset) & (g283) & (g1149)) + ((g34) & (!g36) & (!reset) & (g283) & (!g1149)) + ((g34) & (!g36) & (!reset) & (g283) & (g1149)) + ((g34) & (g36) & (!reset) & (g283) & (!g1149)) + ((g34) & (g36) & (!reset) & (g283) & (g1149)));
	assign g7435 = (((!g832) & (g2404) & (!g1151)) + ((!g832) & (g2404) & (g1151)) + ((g832) & (!g2404) & (g1151)) + ((g832) & (g2404) & (g1151)));
	assign g1152 = (((!g34) & (!g36) & (!reset) & (g284) & (!g1151)) + ((!g34) & (!g36) & (!reset) & (g284) & (g1151)) + ((!g34) & (g36) & (!reset) & (!g284) & (g1151)) + ((!g34) & (g36) & (!reset) & (g284) & (g1151)) + ((g34) & (!g36) & (!reset) & (g284) & (!g1151)) + ((g34) & (!g36) & (!reset) & (g284) & (g1151)) + ((g34) & (g36) & (!reset) & (g284) & (!g1151)) + ((g34) & (g36) & (!reset) & (g284) & (g1151)));
	assign g7436 = (((!g832) & (g2407) & (!g1153)) + ((!g832) & (g2407) & (g1153)) + ((g832) & (!g2407) & (g1153)) + ((g832) & (g2407) & (g1153)));
	assign g1154 = (((!g34) & (!g36) & (!reset) & (g285) & (!g1153)) + ((!g34) & (!g36) & (!reset) & (g285) & (g1153)) + ((!g34) & (g36) & (!reset) & (!g285) & (g1153)) + ((!g34) & (g36) & (!reset) & (g285) & (g1153)) + ((g34) & (!g36) & (!reset) & (g285) & (!g1153)) + ((g34) & (!g36) & (!reset) & (g285) & (g1153)) + ((g34) & (g36) & (!reset) & (g285) & (!g1153)) + ((g34) & (g36) & (!reset) & (g285) & (g1153)));
	assign g7437 = (((!g832) & (g2410) & (!g1155)) + ((!g832) & (g2410) & (g1155)) + ((g832) & (!g2410) & (g1155)) + ((g832) & (g2410) & (g1155)));
	assign g1156 = (((!g34) & (!g36) & (!reset) & (g286) & (!g1155)) + ((!g34) & (!g36) & (!reset) & (g286) & (g1155)) + ((!g34) & (g36) & (!reset) & (!g286) & (g1155)) + ((!g34) & (g36) & (!reset) & (g286) & (g1155)) + ((g34) & (!g36) & (!reset) & (g286) & (!g1155)) + ((g34) & (!g36) & (!reset) & (g286) & (g1155)) + ((g34) & (g36) & (!reset) & (g286) & (!g1155)) + ((g34) & (g36) & (!reset) & (g286) & (g1155)));
	assign g7438 = (((!g832) & (g2412) & (!g1157)) + ((!g832) & (g2412) & (g1157)) + ((g832) & (!g2412) & (g1157)) + ((g832) & (g2412) & (g1157)));
	assign g1158 = (((!g34) & (!g36) & (!reset) & (g288) & (!g1157)) + ((!g34) & (!g36) & (!reset) & (g288) & (g1157)) + ((!g34) & (g36) & (!reset) & (!g288) & (g1157)) + ((!g34) & (g36) & (!reset) & (g288) & (g1157)) + ((g34) & (!g36) & (!reset) & (g288) & (!g1157)) + ((g34) & (!g36) & (!reset) & (g288) & (g1157)) + ((g34) & (g36) & (!reset) & (g288) & (!g1157)) + ((g34) & (g36) & (!reset) & (g288) & (g1157)));
	assign g7439 = (((!g832) & (g2415) & (!g1159)) + ((!g832) & (g2415) & (g1159)) + ((g832) & (!g2415) & (g1159)) + ((g832) & (g2415) & (g1159)));
	assign g1160 = (((!g34) & (!g36) & (!reset) & (g289) & (!g1159)) + ((!g34) & (!g36) & (!reset) & (g289) & (g1159)) + ((!g34) & (g36) & (!reset) & (!g289) & (g1159)) + ((!g34) & (g36) & (!reset) & (g289) & (g1159)) + ((g34) & (!g36) & (!reset) & (g289) & (!g1159)) + ((g34) & (!g36) & (!reset) & (g289) & (g1159)) + ((g34) & (g36) & (!reset) & (g289) & (!g1159)) + ((g34) & (g36) & (!reset) & (g289) & (g1159)));
	assign g7440 = (((!g832) & (g2418) & (!g1161)) + ((!g832) & (g2418) & (g1161)) + ((g832) & (!g2418) & (g1161)) + ((g832) & (g2418) & (g1161)));
	assign g1162 = (((!g34) & (!g36) & (!reset) & (g290) & (!g1161)) + ((!g34) & (!g36) & (!reset) & (g290) & (g1161)) + ((!g34) & (g36) & (!reset) & (!g290) & (g1161)) + ((!g34) & (g36) & (!reset) & (g290) & (g1161)) + ((g34) & (!g36) & (!reset) & (g290) & (!g1161)) + ((g34) & (!g36) & (!reset) & (g290) & (g1161)) + ((g34) & (g36) & (!reset) & (g290) & (!g1161)) + ((g34) & (g36) & (!reset) & (g290) & (g1161)));
	assign g7441 = (((!g832) & (g2421) & (!g1163)) + ((!g832) & (g2421) & (g1163)) + ((g832) & (!g2421) & (g1163)) + ((g832) & (g2421) & (g1163)));
	assign g1164 = (((!g34) & (!g36) & (!reset) & (g291) & (!g1163)) + ((!g34) & (!g36) & (!reset) & (g291) & (g1163)) + ((!g34) & (g36) & (!reset) & (!g291) & (g1163)) + ((!g34) & (g36) & (!reset) & (g291) & (g1163)) + ((g34) & (!g36) & (!reset) & (g291) & (!g1163)) + ((g34) & (!g36) & (!reset) & (g291) & (g1163)) + ((g34) & (g36) & (!reset) & (g291) & (!g1163)) + ((g34) & (g36) & (!reset) & (g291) & (g1163)));
	assign g7442 = (((!g2017) & (g7140) & (!g1165)) + ((!g2017) & (g7140) & (g1165)) + ((g2017) & (!g7140) & (g1165)) + ((g2017) & (g7140) & (g1165)));
	assign g1166 = (((!g248) & (!g271) & (g1098) & (g1132) & (g1099)) + ((!g248) & (g271) & (!g1098) & (g1132) & (!g1099)) + ((!g248) & (g271) & (!g1098) & (g1132) & (g1099)) + ((!g248) & (g271) & (g1098) & (!g1132) & (g1099)) + ((!g248) & (g271) & (g1098) & (g1132) & (!g1099)) + ((!g248) & (g271) & (g1098) & (g1132) & (g1099)) + ((g248) & (!g271) & (!g1098) & (g1132) & (g1099)) + ((g248) & (!g271) & (g1098) & (g1132) & (!g1099)) + ((g248) & (!g271) & (g1098) & (g1132) & (g1099)) + ((g248) & (g271) & (!g1098) & (!g1132) & (g1099)) + ((g248) & (g271) & (!g1098) & (g1132) & (!g1099)) + ((g248) & (g271) & (!g1098) & (g1132) & (g1099)) + ((g248) & (g271) & (g1098) & (!g1132) & (!g1099)) + ((g248) & (g271) & (g1098) & (!g1132) & (g1099)) + ((g248) & (g271) & (g1098) & (g1132) & (!g1099)) + ((g248) & (g271) & (g1098) & (g1132) & (g1099)));
	assign g1167 = (((!g827) & (!g294) & (g1165) & (!g1166)) + ((!g827) & (!g294) & (g1165) & (g1166)) + ((!g827) & (g294) & (g1165) & (!g1166)) + ((!g827) & (g294) & (g1165) & (g1166)) + ((g827) & (!g294) & (!g1165) & (g1166)) + ((g827) & (!g294) & (g1165) & (!g1166)) + ((g827) & (g294) & (!g1165) & (!g1166)) + ((g827) & (g294) & (g1165) & (g1166)));
	assign g1168 = (((!g34) & (!g36) & (!reset) & (g296) & (!g317)) + ((!g34) & (!g36) & (!reset) & (g296) & (g317)) + ((!g34) & (g36) & (!reset) & (!g296) & (g317)) + ((!g34) & (g36) & (!reset) & (g296) & (g317)) + ((g34) & (!g36) & (!reset) & (g296) & (!g317)) + ((g34) & (!g36) & (!reset) & (g296) & (g317)) + ((g34) & (g36) & (!reset) & (g296) & (!g317)) + ((g34) & (g36) & (!reset) & (g296) & (g317)));
	assign g7443 = (((!g832) & (g2433) & (!g1169)) + ((!g832) & (g2433) & (g1169)) + ((g832) & (!g2433) & (g1169)) + ((g832) & (g2433) & (g1169)));
	assign g1170 = (((!g34) & (!g36) & (!reset) & (g297) & (!g1169)) + ((!g34) & (!g36) & (!reset) & (g297) & (g1169)) + ((!g34) & (g36) & (!reset) & (!g297) & (g1169)) + ((!g34) & (g36) & (!reset) & (g297) & (g1169)) + ((g34) & (!g36) & (!reset) & (g297) & (!g1169)) + ((g34) & (!g36) & (!reset) & (g297) & (g1169)) + ((g34) & (g36) & (!reset) & (g297) & (!g1169)) + ((g34) & (g36) & (!reset) & (g297) & (g1169)));
	assign g7444 = (((!g832) & (g2439) & (!g1171)) + ((!g832) & (g2439) & (g1171)) + ((g832) & (!g2439) & (g1171)) + ((g832) & (g2439) & (g1171)));
	assign g1172 = (((!g34) & (!g36) & (!reset) & (g298) & (!g1171)) + ((!g34) & (!g36) & (!reset) & (g298) & (g1171)) + ((!g34) & (g36) & (!reset) & (!g298) & (g1171)) + ((!g34) & (g36) & (!reset) & (g298) & (g1171)) + ((g34) & (!g36) & (!reset) & (g298) & (!g1171)) + ((g34) & (!g36) & (!reset) & (g298) & (g1171)) + ((g34) & (g36) & (!reset) & (g298) & (!g1171)) + ((g34) & (g36) & (!reset) & (g298) & (g1171)));
	assign g7445 = (((!g832) & (g2444) & (!g1173)) + ((!g832) & (g2444) & (g1173)) + ((g832) & (!g2444) & (g1173)) + ((g832) & (g2444) & (g1173)));
	assign g1174 = (((!g34) & (!g36) & (!reset) & (g299) & (!g1173)) + ((!g34) & (!g36) & (!reset) & (g299) & (g1173)) + ((!g34) & (g36) & (!reset) & (!g299) & (g1173)) + ((!g34) & (g36) & (!reset) & (g299) & (g1173)) + ((g34) & (!g36) & (!reset) & (g299) & (!g1173)) + ((g34) & (!g36) & (!reset) & (g299) & (g1173)) + ((g34) & (g36) & (!reset) & (g299) & (!g1173)) + ((g34) & (g36) & (!reset) & (g299) & (g1173)));
	assign g7446 = (((!g832) & (g2449) & (!g1175)) + ((!g832) & (g2449) & (g1175)) + ((g832) & (!g2449) & (g1175)) + ((g832) & (g2449) & (g1175)));
	assign g1176 = (((!g34) & (!g36) & (!reset) & (g301) & (!g1175)) + ((!g34) & (!g36) & (!reset) & (g301) & (g1175)) + ((!g34) & (g36) & (!reset) & (!g301) & (g1175)) + ((!g34) & (g36) & (!reset) & (g301) & (g1175)) + ((g34) & (!g36) & (!reset) & (g301) & (!g1175)) + ((g34) & (!g36) & (!reset) & (g301) & (g1175)) + ((g34) & (g36) & (!reset) & (g301) & (!g1175)) + ((g34) & (g36) & (!reset) & (g301) & (g1175)));
	assign g7447 = (((!g832) & (g2455) & (!g1177)) + ((!g832) & (g2455) & (g1177)) + ((g832) & (!g2455) & (g1177)) + ((g832) & (g2455) & (g1177)));
	assign g1178 = (((!g34) & (!g36) & (!reset) & (g302) & (!g1177)) + ((!g34) & (!g36) & (!reset) & (g302) & (g1177)) + ((!g34) & (g36) & (!reset) & (!g302) & (g1177)) + ((!g34) & (g36) & (!reset) & (g302) & (g1177)) + ((g34) & (!g36) & (!reset) & (g302) & (!g1177)) + ((g34) & (!g36) & (!reset) & (g302) & (g1177)) + ((g34) & (g36) & (!reset) & (g302) & (!g1177)) + ((g34) & (g36) & (!reset) & (g302) & (g1177)));
	assign g7448 = (((!g832) & (g2461) & (!g1179)) + ((!g832) & (g2461) & (g1179)) + ((g832) & (!g2461) & (g1179)) + ((g832) & (g2461) & (g1179)));
	assign g1180 = (((!g34) & (!g36) & (!reset) & (g303) & (!g1179)) + ((!g34) & (!g36) & (!reset) & (g303) & (g1179)) + ((!g34) & (g36) & (!reset) & (!g303) & (g1179)) + ((!g34) & (g36) & (!reset) & (g303) & (g1179)) + ((g34) & (!g36) & (!reset) & (g303) & (!g1179)) + ((g34) & (!g36) & (!reset) & (g303) & (g1179)) + ((g34) & (g36) & (!reset) & (g303) & (!g1179)) + ((g34) & (g36) & (!reset) & (g303) & (g1179)));
	assign g7449 = (((!g832) & (g2467) & (!g1181)) + ((!g832) & (g2467) & (g1181)) + ((g832) & (!g2467) & (g1181)) + ((g832) & (g2467) & (g1181)));
	assign g1182 = (((!g34) & (!g36) & (!reset) & (g304) & (!g1181)) + ((!g34) & (!g36) & (!reset) & (g304) & (g1181)) + ((!g34) & (g36) & (!reset) & (!g304) & (g1181)) + ((!g34) & (g36) & (!reset) & (g304) & (g1181)) + ((g34) & (!g36) & (!reset) & (g304) & (!g1181)) + ((g34) & (!g36) & (!reset) & (g304) & (g1181)) + ((g34) & (g36) & (!reset) & (g304) & (!g1181)) + ((g34) & (g36) & (!reset) & (g304) & (g1181)));
	assign g7450 = (((!g832) & (g2473) & (!g1183)) + ((!g832) & (g2473) & (g1183)) + ((g832) & (!g2473) & (g1183)) + ((g832) & (g2473) & (g1183)));
	assign g1184 = (((!g34) & (!g36) & (!reset) & (g306) & (!g1183)) + ((!g34) & (!g36) & (!reset) & (g306) & (g1183)) + ((!g34) & (g36) & (!reset) & (!g306) & (g1183)) + ((!g34) & (g36) & (!reset) & (g306) & (g1183)) + ((g34) & (!g36) & (!reset) & (g306) & (!g1183)) + ((g34) & (!g36) & (!reset) & (g306) & (g1183)) + ((g34) & (g36) & (!reset) & (g306) & (!g1183)) + ((g34) & (g36) & (!reset) & (g306) & (g1183)));
	assign g7451 = (((!g832) & (g2479) & (!g1185)) + ((!g832) & (g2479) & (g1185)) + ((g832) & (!g2479) & (g1185)) + ((g832) & (g2479) & (g1185)));
	assign g1186 = (((!g34) & (!g36) & (!reset) & (g307) & (!g1185)) + ((!g34) & (!g36) & (!reset) & (g307) & (g1185)) + ((!g34) & (g36) & (!reset) & (!g307) & (g1185)) + ((!g34) & (g36) & (!reset) & (g307) & (g1185)) + ((g34) & (!g36) & (!reset) & (g307) & (!g1185)) + ((g34) & (!g36) & (!reset) & (g307) & (g1185)) + ((g34) & (g36) & (!reset) & (g307) & (!g1185)) + ((g34) & (g36) & (!reset) & (g307) & (g1185)));
	assign g7452 = (((!g832) & (g2485) & (!g1187)) + ((!g832) & (g2485) & (g1187)) + ((g832) & (!g2485) & (g1187)) + ((g832) & (g2485) & (g1187)));
	assign g1188 = (((!g34) & (!g36) & (!reset) & (g308) & (!g1187)) + ((!g34) & (!g36) & (!reset) & (g308) & (g1187)) + ((!g34) & (g36) & (!reset) & (!g308) & (g1187)) + ((!g34) & (g36) & (!reset) & (g308) & (g1187)) + ((g34) & (!g36) & (!reset) & (g308) & (!g1187)) + ((g34) & (!g36) & (!reset) & (g308) & (g1187)) + ((g34) & (g36) & (!reset) & (g308) & (!g1187)) + ((g34) & (g36) & (!reset) & (g308) & (g1187)));
	assign g7453 = (((!g832) & (g2491) & (!g1189)) + ((!g832) & (g2491) & (g1189)) + ((g832) & (!g2491) & (g1189)) + ((g832) & (g2491) & (g1189)));
	assign g1190 = (((!g34) & (!g36) & (!reset) & (g309) & (!g1189)) + ((!g34) & (!g36) & (!reset) & (g309) & (g1189)) + ((!g34) & (g36) & (!reset) & (!g309) & (g1189)) + ((!g34) & (g36) & (!reset) & (g309) & (g1189)) + ((g34) & (!g36) & (!reset) & (g309) & (!g1189)) + ((g34) & (!g36) & (!reset) & (g309) & (g1189)) + ((g34) & (g36) & (!reset) & (g309) & (!g1189)) + ((g34) & (g36) & (!reset) & (g309) & (g1189)));
	assign g7454 = (((!g832) & (g2496) & (!g1191)) + ((!g832) & (g2496) & (g1191)) + ((g832) & (!g2496) & (g1191)) + ((g832) & (g2496) & (g1191)));
	assign g1192 = (((!g34) & (!g36) & (!reset) & (g311) & (!g1191)) + ((!g34) & (!g36) & (!reset) & (g311) & (g1191)) + ((!g34) & (g36) & (!reset) & (!g311) & (g1191)) + ((!g34) & (g36) & (!reset) & (g311) & (g1191)) + ((g34) & (!g36) & (!reset) & (g311) & (!g1191)) + ((g34) & (!g36) & (!reset) & (g311) & (g1191)) + ((g34) & (g36) & (!reset) & (g311) & (!g1191)) + ((g34) & (g36) & (!reset) & (g311) & (g1191)));
	assign g7455 = (((!g832) & (g2502) & (!g1193)) + ((!g832) & (g2502) & (g1193)) + ((g832) & (!g2502) & (g1193)) + ((g832) & (g2502) & (g1193)));
	assign g1194 = (((!g34) & (!g36) & (!reset) & (g312) & (!g1193)) + ((!g34) & (!g36) & (!reset) & (g312) & (g1193)) + ((!g34) & (g36) & (!reset) & (!g312) & (g1193)) + ((!g34) & (g36) & (!reset) & (g312) & (g1193)) + ((g34) & (!g36) & (!reset) & (g312) & (!g1193)) + ((g34) & (!g36) & (!reset) & (g312) & (g1193)) + ((g34) & (g36) & (!reset) & (g312) & (!g1193)) + ((g34) & (g36) & (!reset) & (g312) & (g1193)));
	assign g7456 = (((!g832) & (g2508) & (!g1195)) + ((!g832) & (g2508) & (g1195)) + ((g832) & (!g2508) & (g1195)) + ((g832) & (g2508) & (g1195)));
	assign g1196 = (((!g34) & (!g36) & (!reset) & (g313) & (!g1195)) + ((!g34) & (!g36) & (!reset) & (g313) & (g1195)) + ((!g34) & (g36) & (!reset) & (!g313) & (g1195)) + ((!g34) & (g36) & (!reset) & (g313) & (g1195)) + ((g34) & (!g36) & (!reset) & (g313) & (!g1195)) + ((g34) & (!g36) & (!reset) & (g313) & (g1195)) + ((g34) & (g36) & (!reset) & (g313) & (!g1195)) + ((g34) & (g36) & (!reset) & (g313) & (g1195)));
	assign g7457 = (((!g832) & (g2514) & (!g1197)) + ((!g832) & (g2514) & (g1197)) + ((g832) & (!g2514) & (g1197)) + ((g832) & (g2514) & (g1197)));
	assign g1198 = (((!g34) & (!g36) & (!reset) & (g314) & (!g1197)) + ((!g34) & (!g36) & (!reset) & (g314) & (g1197)) + ((!g34) & (g36) & (!reset) & (!g314) & (g1197)) + ((!g34) & (g36) & (!reset) & (g314) & (g1197)) + ((g34) & (!g36) & (!reset) & (g314) & (!g1197)) + ((g34) & (!g36) & (!reset) & (g314) & (g1197)) + ((g34) & (g36) & (!reset) & (g314) & (!g1197)) + ((g34) & (g36) & (!reset) & (g314) & (g1197)));
	assign g7458 = (((!g2017) & (g2521) & (!g1199)) + ((!g2017) & (g2521) & (g1199)) + ((g2017) & (!g2521) & (g1199)) + ((g2017) & (g2521) & (g1199)));
	assign g1200 = (((!g294) & (g1165)) + ((g294) & (!g1165)));
	assign g1201 = (((!g248) & (!g271) & (g1098) & (g1132) & (g1099) & (g1200)) + ((!g248) & (g271) & (!g1098) & (g1132) & (!g1099) & (g1200)) + ((!g248) & (g271) & (!g1098) & (g1132) & (g1099) & (g1200)) + ((!g248) & (g271) & (g1098) & (!g1132) & (g1099) & (g1200)) + ((!g248) & (g271) & (g1098) & (g1132) & (!g1099) & (g1200)) + ((!g248) & (g271) & (g1098) & (g1132) & (g1099) & (g1200)) + ((g248) & (!g271) & (!g1098) & (g1132) & (g1099) & (g1200)) + ((g248) & (!g271) & (g1098) & (g1132) & (!g1099) & (g1200)) + ((g248) & (!g271) & (g1098) & (g1132) & (g1099) & (g1200)) + ((g248) & (g271) & (!g1098) & (!g1132) & (g1099) & (g1200)) + ((g248) & (g271) & (!g1098) & (g1132) & (!g1099) & (g1200)) + ((g248) & (g271) & (!g1098) & (g1132) & (g1099) & (g1200)) + ((g248) & (g271) & (g1098) & (!g1132) & (!g1099) & (g1200)) + ((g248) & (g271) & (g1098) & (!g1132) & (g1099) & (g1200)) + ((g248) & (g271) & (g1098) & (g1132) & (!g1099) & (g1200)) + ((g248) & (g271) & (g1098) & (g1132) & (g1099) & (g1200)));
	assign g1202 = (((g294) & (g1165)));
	assign g1203 = (((!g1201) & (!g1202)));
	assign g1204 = (((!g827) & (!g317) & (g1199) & (!g1203)) + ((!g827) & (!g317) & (g1199) & (g1203)) + ((!g827) & (g317) & (g1199) & (!g1203)) + ((!g827) & (g317) & (g1199) & (g1203)) + ((g827) & (!g317) & (!g1199) & (!g1203)) + ((g827) & (!g317) & (g1199) & (g1203)) + ((g827) & (g317) & (!g1199) & (g1203)) + ((g827) & (g317) & (g1199) & (!g1203)));
	assign g1205 = (((!g34) & (!g36) & (!reset) & (g319) & (!g340)) + ((!g34) & (!g36) & (!reset) & (g319) & (g340)) + ((!g34) & (g36) & (!reset) & (!g319) & (g340)) + ((!g34) & (g36) & (!reset) & (g319) & (g340)) + ((g34) & (!g36) & (!reset) & (g319) & (!g340)) + ((g34) & (!g36) & (!reset) & (g319) & (g340)) + ((g34) & (g36) & (!reset) & (g319) & (!g340)) + ((g34) & (g36) & (!reset) & (g319) & (g340)));
	assign g7459 = (((!g832) & (g2522) & (!g1206)) + ((!g832) & (g2522) & (g1206)) + ((g832) & (!g2522) & (g1206)) + ((g832) & (g2522) & (g1206)));
	assign g1207 = (((!g34) & (!g36) & (!reset) & (g320) & (!g1206)) + ((!g34) & (!g36) & (!reset) & (g320) & (g1206)) + ((!g34) & (g36) & (!reset) & (!g320) & (g1206)) + ((!g34) & (g36) & (!reset) & (g320) & (g1206)) + ((g34) & (!g36) & (!reset) & (g320) & (!g1206)) + ((g34) & (!g36) & (!reset) & (g320) & (g1206)) + ((g34) & (g36) & (!reset) & (g320) & (!g1206)) + ((g34) & (g36) & (!reset) & (g320) & (g1206)));
	assign g7460 = (((!g832) & (g2524) & (!g1208)) + ((!g832) & (g2524) & (g1208)) + ((g832) & (!g2524) & (g1208)) + ((g832) & (g2524) & (g1208)));
	assign g1209 = (((!g34) & (!g36) & (!reset) & (g321) & (!g1208)) + ((!g34) & (!g36) & (!reset) & (g321) & (g1208)) + ((!g34) & (g36) & (!reset) & (!g321) & (g1208)) + ((!g34) & (g36) & (!reset) & (g321) & (g1208)) + ((g34) & (!g36) & (!reset) & (g321) & (!g1208)) + ((g34) & (!g36) & (!reset) & (g321) & (g1208)) + ((g34) & (g36) & (!reset) & (g321) & (!g1208)) + ((g34) & (g36) & (!reset) & (g321) & (g1208)));
	assign g7461 = (((!g832) & (g2525) & (!g1210)) + ((!g832) & (g2525) & (g1210)) + ((g832) & (!g2525) & (g1210)) + ((g832) & (g2525) & (g1210)));
	assign g1211 = (((!g34) & (!g36) & (!reset) & (g322) & (!g1210)) + ((!g34) & (!g36) & (!reset) & (g322) & (g1210)) + ((!g34) & (g36) & (!reset) & (!g322) & (g1210)) + ((!g34) & (g36) & (!reset) & (g322) & (g1210)) + ((g34) & (!g36) & (!reset) & (g322) & (!g1210)) + ((g34) & (!g36) & (!reset) & (g322) & (g1210)) + ((g34) & (g36) & (!reset) & (g322) & (!g1210)) + ((g34) & (g36) & (!reset) & (g322) & (g1210)));
	assign g7462 = (((!g832) & (g2526) & (!g1212)) + ((!g832) & (g2526) & (g1212)) + ((g832) & (!g2526) & (g1212)) + ((g832) & (g2526) & (g1212)));
	assign g1213 = (((!g34) & (!g36) & (!reset) & (g324) & (!g1212)) + ((!g34) & (!g36) & (!reset) & (g324) & (g1212)) + ((!g34) & (g36) & (!reset) & (!g324) & (g1212)) + ((!g34) & (g36) & (!reset) & (g324) & (g1212)) + ((g34) & (!g36) & (!reset) & (g324) & (!g1212)) + ((g34) & (!g36) & (!reset) & (g324) & (g1212)) + ((g34) & (g36) & (!reset) & (g324) & (!g1212)) + ((g34) & (g36) & (!reset) & (g324) & (g1212)));
	assign g7463 = (((!g832) & (g2528) & (!g1214)) + ((!g832) & (g2528) & (g1214)) + ((g832) & (!g2528) & (g1214)) + ((g832) & (g2528) & (g1214)));
	assign g1215 = (((!g34) & (!g36) & (!reset) & (g325) & (!g1214)) + ((!g34) & (!g36) & (!reset) & (g325) & (g1214)) + ((!g34) & (g36) & (!reset) & (!g325) & (g1214)) + ((!g34) & (g36) & (!reset) & (g325) & (g1214)) + ((g34) & (!g36) & (!reset) & (g325) & (!g1214)) + ((g34) & (!g36) & (!reset) & (g325) & (g1214)) + ((g34) & (g36) & (!reset) & (g325) & (!g1214)) + ((g34) & (g36) & (!reset) & (g325) & (g1214)));
	assign g7464 = (((!g832) & (g2530) & (!g1216)) + ((!g832) & (g2530) & (g1216)) + ((g832) & (!g2530) & (g1216)) + ((g832) & (g2530) & (g1216)));
	assign g1217 = (((!g34) & (!g36) & (!reset) & (g326) & (!g1216)) + ((!g34) & (!g36) & (!reset) & (g326) & (g1216)) + ((!g34) & (g36) & (!reset) & (!g326) & (g1216)) + ((!g34) & (g36) & (!reset) & (g326) & (g1216)) + ((g34) & (!g36) & (!reset) & (g326) & (!g1216)) + ((g34) & (!g36) & (!reset) & (g326) & (g1216)) + ((g34) & (g36) & (!reset) & (g326) & (!g1216)) + ((g34) & (g36) & (!reset) & (g326) & (g1216)));
	assign g7465 = (((!g832) & (g2532) & (!g1218)) + ((!g832) & (g2532) & (g1218)) + ((g832) & (!g2532) & (g1218)) + ((g832) & (g2532) & (g1218)));
	assign g1219 = (((!g34) & (!g36) & (!reset) & (g327) & (!g1218)) + ((!g34) & (!g36) & (!reset) & (g327) & (g1218)) + ((!g34) & (g36) & (!reset) & (!g327) & (g1218)) + ((!g34) & (g36) & (!reset) & (g327) & (g1218)) + ((g34) & (!g36) & (!reset) & (g327) & (!g1218)) + ((g34) & (!g36) & (!reset) & (g327) & (g1218)) + ((g34) & (g36) & (!reset) & (g327) & (!g1218)) + ((g34) & (g36) & (!reset) & (g327) & (g1218)));
	assign g7466 = (((!g832) & (g2534) & (!g1220)) + ((!g832) & (g2534) & (g1220)) + ((g832) & (!g2534) & (g1220)) + ((g832) & (g2534) & (g1220)));
	assign g1221 = (((!g34) & (!g36) & (!reset) & (g329) & (!g1220)) + ((!g34) & (!g36) & (!reset) & (g329) & (g1220)) + ((!g34) & (g36) & (!reset) & (!g329) & (g1220)) + ((!g34) & (g36) & (!reset) & (g329) & (g1220)) + ((g34) & (!g36) & (!reset) & (g329) & (!g1220)) + ((g34) & (!g36) & (!reset) & (g329) & (g1220)) + ((g34) & (g36) & (!reset) & (g329) & (!g1220)) + ((g34) & (g36) & (!reset) & (g329) & (g1220)));
	assign g7467 = (((!g832) & (g2536) & (!g1222)) + ((!g832) & (g2536) & (g1222)) + ((g832) & (!g2536) & (g1222)) + ((g832) & (g2536) & (g1222)));
	assign g1223 = (((!g34) & (!g36) & (!reset) & (g330) & (!g1222)) + ((!g34) & (!g36) & (!reset) & (g330) & (g1222)) + ((!g34) & (g36) & (!reset) & (!g330) & (g1222)) + ((!g34) & (g36) & (!reset) & (g330) & (g1222)) + ((g34) & (!g36) & (!reset) & (g330) & (!g1222)) + ((g34) & (!g36) & (!reset) & (g330) & (g1222)) + ((g34) & (g36) & (!reset) & (g330) & (!g1222)) + ((g34) & (g36) & (!reset) & (g330) & (g1222)));
	assign g7468 = (((!g832) & (g2538) & (!g1224)) + ((!g832) & (g2538) & (g1224)) + ((g832) & (!g2538) & (g1224)) + ((g832) & (g2538) & (g1224)));
	assign g1225 = (((!g34) & (!g36) & (!reset) & (g331) & (!g1224)) + ((!g34) & (!g36) & (!reset) & (g331) & (g1224)) + ((!g34) & (g36) & (!reset) & (!g331) & (g1224)) + ((!g34) & (g36) & (!reset) & (g331) & (g1224)) + ((g34) & (!g36) & (!reset) & (g331) & (!g1224)) + ((g34) & (!g36) & (!reset) & (g331) & (g1224)) + ((g34) & (g36) & (!reset) & (g331) & (!g1224)) + ((g34) & (g36) & (!reset) & (g331) & (g1224)));
	assign g7469 = (((!g832) & (g2540) & (!g1226)) + ((!g832) & (g2540) & (g1226)) + ((g832) & (!g2540) & (g1226)) + ((g832) & (g2540) & (g1226)));
	assign g1227 = (((!g34) & (!g36) & (!reset) & (g332) & (!g1226)) + ((!g34) & (!g36) & (!reset) & (g332) & (g1226)) + ((!g34) & (g36) & (!reset) & (!g332) & (g1226)) + ((!g34) & (g36) & (!reset) & (g332) & (g1226)) + ((g34) & (!g36) & (!reset) & (g332) & (!g1226)) + ((g34) & (!g36) & (!reset) & (g332) & (g1226)) + ((g34) & (g36) & (!reset) & (g332) & (!g1226)) + ((g34) & (g36) & (!reset) & (g332) & (g1226)));
	assign g7470 = (((!g832) & (g2541) & (!g1228)) + ((!g832) & (g2541) & (g1228)) + ((g832) & (!g2541) & (g1228)) + ((g832) & (g2541) & (g1228)));
	assign g1229 = (((!g34) & (!g36) & (!reset) & (g334) & (!g1228)) + ((!g34) & (!g36) & (!reset) & (g334) & (g1228)) + ((!g34) & (g36) & (!reset) & (!g334) & (g1228)) + ((!g34) & (g36) & (!reset) & (g334) & (g1228)) + ((g34) & (!g36) & (!reset) & (g334) & (!g1228)) + ((g34) & (!g36) & (!reset) & (g334) & (g1228)) + ((g34) & (g36) & (!reset) & (g334) & (!g1228)) + ((g34) & (g36) & (!reset) & (g334) & (g1228)));
	assign g7471 = (((!g832) & (g2543) & (!g1230)) + ((!g832) & (g2543) & (g1230)) + ((g832) & (!g2543) & (g1230)) + ((g832) & (g2543) & (g1230)));
	assign g1231 = (((!g34) & (!g36) & (!reset) & (g335) & (!g1230)) + ((!g34) & (!g36) & (!reset) & (g335) & (g1230)) + ((!g34) & (g36) & (!reset) & (!g335) & (g1230)) + ((!g34) & (g36) & (!reset) & (g335) & (g1230)) + ((g34) & (!g36) & (!reset) & (g335) & (!g1230)) + ((g34) & (!g36) & (!reset) & (g335) & (g1230)) + ((g34) & (g36) & (!reset) & (g335) & (!g1230)) + ((g34) & (g36) & (!reset) & (g335) & (g1230)));
	assign g7472 = (((!g832) & (g2545) & (!g1232)) + ((!g832) & (g2545) & (g1232)) + ((g832) & (!g2545) & (g1232)) + ((g832) & (g2545) & (g1232)));
	assign g1233 = (((!g34) & (!g36) & (!reset) & (g336) & (!g1232)) + ((!g34) & (!g36) & (!reset) & (g336) & (g1232)) + ((!g34) & (g36) & (!reset) & (!g336) & (g1232)) + ((!g34) & (g36) & (!reset) & (g336) & (g1232)) + ((g34) & (!g36) & (!reset) & (g336) & (!g1232)) + ((g34) & (!g36) & (!reset) & (g336) & (g1232)) + ((g34) & (g36) & (!reset) & (g336) & (!g1232)) + ((g34) & (g36) & (!reset) & (g336) & (g1232)));
	assign g7473 = (((!g832) & (g2547) & (!g1234)) + ((!g832) & (g2547) & (g1234)) + ((g832) & (!g2547) & (g1234)) + ((g832) & (g2547) & (g1234)));
	assign g1235 = (((!g34) & (!g36) & (!reset) & (g337) & (!g1234)) + ((!g34) & (!g36) & (!reset) & (g337) & (g1234)) + ((!g34) & (g36) & (!reset) & (!g337) & (g1234)) + ((!g34) & (g36) & (!reset) & (g337) & (g1234)) + ((g34) & (!g36) & (!reset) & (g337) & (!g1234)) + ((g34) & (!g36) & (!reset) & (g337) & (g1234)) + ((g34) & (g36) & (!reset) & (g337) & (!g1234)) + ((g34) & (g36) & (!reset) & (g337) & (g1234)));
	assign g7474 = (((!g2017) & (g7133) & (!g1236)) + ((!g2017) & (g7133) & (g1236)) + ((g2017) & (!g7133) & (g1236)) + ((g2017) & (g7133) & (g1236)));
	assign g1237 = (((!g827) & (!g317) & (!g340) & (!g1199) & (g1236) & (!g1203)) + ((!g827) & (!g317) & (!g340) & (!g1199) & (g1236) & (g1203)) + ((!g827) & (!g317) & (!g340) & (g1199) & (g1236) & (!g1203)) + ((!g827) & (!g317) & (!g340) & (g1199) & (g1236) & (g1203)) + ((!g827) & (!g317) & (g340) & (!g1199) & (g1236) & (!g1203)) + ((!g827) & (!g317) & (g340) & (!g1199) & (g1236) & (g1203)) + ((!g827) & (!g317) & (g340) & (g1199) & (g1236) & (!g1203)) + ((!g827) & (!g317) & (g340) & (g1199) & (g1236) & (g1203)) + ((!g827) & (g317) & (!g340) & (!g1199) & (g1236) & (!g1203)) + ((!g827) & (g317) & (!g340) & (!g1199) & (g1236) & (g1203)) + ((!g827) & (g317) & (!g340) & (g1199) & (g1236) & (!g1203)) + ((!g827) & (g317) & (!g340) & (g1199) & (g1236) & (g1203)) + ((!g827) & (g317) & (g340) & (!g1199) & (g1236) & (!g1203)) + ((!g827) & (g317) & (g340) & (!g1199) & (g1236) & (g1203)) + ((!g827) & (g317) & (g340) & (g1199) & (g1236) & (!g1203)) + ((!g827) & (g317) & (g340) & (g1199) & (g1236) & (g1203)) + ((g827) & (!g317) & (!g340) & (!g1199) & (g1236) & (!g1203)) + ((g827) & (!g317) & (!g340) & (!g1199) & (g1236) & (g1203)) + ((g827) & (!g317) & (!g340) & (g1199) & (!g1236) & (!g1203)) + ((g827) & (!g317) & (!g340) & (g1199) & (g1236) & (g1203)) + ((g827) & (!g317) & (g340) & (!g1199) & (!g1236) & (!g1203)) + ((g827) & (!g317) & (g340) & (!g1199) & (!g1236) & (g1203)) + ((g827) & (!g317) & (g340) & (g1199) & (!g1236) & (g1203)) + ((g827) & (!g317) & (g340) & (g1199) & (g1236) & (!g1203)) + ((g827) & (g317) & (!g340) & (!g1199) & (!g1236) & (!g1203)) + ((g827) & (g317) & (!g340) & (!g1199) & (g1236) & (g1203)) + ((g827) & (g317) & (!g340) & (g1199) & (!g1236) & (!g1203)) + ((g827) & (g317) & (!g340) & (g1199) & (!g1236) & (g1203)) + ((g827) & (g317) & (g340) & (!g1199) & (!g1236) & (g1203)) + ((g827) & (g317) & (g340) & (!g1199) & (g1236) & (!g1203)) + ((g827) & (g317) & (g340) & (g1199) & (g1236) & (!g1203)) + ((g827) & (g317) & (g340) & (g1199) & (g1236) & (g1203)));
	assign g1238 = (((!g34) & (!g36) & (!reset) & (g342) & (!g363)) + ((!g34) & (!g36) & (!reset) & (g342) & (g363)) + ((!g34) & (g36) & (!reset) & (!g342) & (g363)) + ((!g34) & (g36) & (!reset) & (g342) & (g363)) + ((g34) & (!g36) & (!reset) & (g342) & (!g363)) + ((g34) & (!g36) & (!reset) & (g342) & (g363)) + ((g34) & (g36) & (!reset) & (g342) & (!g363)) + ((g34) & (g36) & (!reset) & (g342) & (g363)));
	assign g7475 = (((!g832) & (g2558) & (!g1239)) + ((!g832) & (g2558) & (g1239)) + ((g832) & (!g2558) & (g1239)) + ((g832) & (g2558) & (g1239)));
	assign g1240 = (((!g34) & (!g36) & (!reset) & (g343) & (!g1239)) + ((!g34) & (!g36) & (!reset) & (g343) & (g1239)) + ((!g34) & (g36) & (!reset) & (!g343) & (g1239)) + ((!g34) & (g36) & (!reset) & (g343) & (g1239)) + ((g34) & (!g36) & (!reset) & (g343) & (!g1239)) + ((g34) & (!g36) & (!reset) & (g343) & (g1239)) + ((g34) & (g36) & (!reset) & (g343) & (!g1239)) + ((g34) & (g36) & (!reset) & (g343) & (g1239)));
	assign g7476 = (((!g832) & (g2561) & (!g1241)) + ((!g832) & (g2561) & (g1241)) + ((g832) & (!g2561) & (g1241)) + ((g832) & (g2561) & (g1241)));
	assign g1242 = (((!g34) & (!g36) & (!reset) & (g344) & (!g1241)) + ((!g34) & (!g36) & (!reset) & (g344) & (g1241)) + ((!g34) & (g36) & (!reset) & (!g344) & (g1241)) + ((!g34) & (g36) & (!reset) & (g344) & (g1241)) + ((g34) & (!g36) & (!reset) & (g344) & (!g1241)) + ((g34) & (!g36) & (!reset) & (g344) & (g1241)) + ((g34) & (g36) & (!reset) & (g344) & (!g1241)) + ((g34) & (g36) & (!reset) & (g344) & (g1241)));
	assign g7477 = (((!g832) & (g2563) & (!g1243)) + ((!g832) & (g2563) & (g1243)) + ((g832) & (!g2563) & (g1243)) + ((g832) & (g2563) & (g1243)));
	assign g1244 = (((!g34) & (!g36) & (!reset) & (g345) & (!g1243)) + ((!g34) & (!g36) & (!reset) & (g345) & (g1243)) + ((!g34) & (g36) & (!reset) & (!g345) & (g1243)) + ((!g34) & (g36) & (!reset) & (g345) & (g1243)) + ((g34) & (!g36) & (!reset) & (g345) & (!g1243)) + ((g34) & (!g36) & (!reset) & (g345) & (g1243)) + ((g34) & (g36) & (!reset) & (g345) & (!g1243)) + ((g34) & (g36) & (!reset) & (g345) & (g1243)));
	assign g7478 = (((!g832) & (g2565) & (!g1245)) + ((!g832) & (g2565) & (g1245)) + ((g832) & (!g2565) & (g1245)) + ((g832) & (g2565) & (g1245)));
	assign g1246 = (((!g34) & (!g36) & (!reset) & (g347) & (!g1245)) + ((!g34) & (!g36) & (!reset) & (g347) & (g1245)) + ((!g34) & (g36) & (!reset) & (!g347) & (g1245)) + ((!g34) & (g36) & (!reset) & (g347) & (g1245)) + ((g34) & (!g36) & (!reset) & (g347) & (!g1245)) + ((g34) & (!g36) & (!reset) & (g347) & (g1245)) + ((g34) & (g36) & (!reset) & (g347) & (!g1245)) + ((g34) & (g36) & (!reset) & (g347) & (g1245)));
	assign g7479 = (((!g832) & (g2568) & (!g1247)) + ((!g832) & (g2568) & (g1247)) + ((g832) & (!g2568) & (g1247)) + ((g832) & (g2568) & (g1247)));
	assign g1248 = (((!g34) & (!g36) & (!reset) & (g348) & (!g1247)) + ((!g34) & (!g36) & (!reset) & (g348) & (g1247)) + ((!g34) & (g36) & (!reset) & (!g348) & (g1247)) + ((!g34) & (g36) & (!reset) & (g348) & (g1247)) + ((g34) & (!g36) & (!reset) & (g348) & (!g1247)) + ((g34) & (!g36) & (!reset) & (g348) & (g1247)) + ((g34) & (g36) & (!reset) & (g348) & (!g1247)) + ((g34) & (g36) & (!reset) & (g348) & (g1247)));
	assign g7480 = (((!g832) & (g2571) & (!g1249)) + ((!g832) & (g2571) & (g1249)) + ((g832) & (!g2571) & (g1249)) + ((g832) & (g2571) & (g1249)));
	assign g1250 = (((!g34) & (!g36) & (!reset) & (g349) & (!g1249)) + ((!g34) & (!g36) & (!reset) & (g349) & (g1249)) + ((!g34) & (g36) & (!reset) & (!g349) & (g1249)) + ((!g34) & (g36) & (!reset) & (g349) & (g1249)) + ((g34) & (!g36) & (!reset) & (g349) & (!g1249)) + ((g34) & (!g36) & (!reset) & (g349) & (g1249)) + ((g34) & (g36) & (!reset) & (g349) & (!g1249)) + ((g34) & (g36) & (!reset) & (g349) & (g1249)));
	assign g7481 = (((!g832) & (g2574) & (!g1251)) + ((!g832) & (g2574) & (g1251)) + ((g832) & (!g2574) & (g1251)) + ((g832) & (g2574) & (g1251)));
	assign g1252 = (((!g34) & (!g36) & (!reset) & (g350) & (!g1251)) + ((!g34) & (!g36) & (!reset) & (g350) & (g1251)) + ((!g34) & (g36) & (!reset) & (!g350) & (g1251)) + ((!g34) & (g36) & (!reset) & (g350) & (g1251)) + ((g34) & (!g36) & (!reset) & (g350) & (!g1251)) + ((g34) & (!g36) & (!reset) & (g350) & (g1251)) + ((g34) & (g36) & (!reset) & (g350) & (!g1251)) + ((g34) & (g36) & (!reset) & (g350) & (g1251)));
	assign g7482 = (((!g832) & (g2577) & (!g1253)) + ((!g832) & (g2577) & (g1253)) + ((g832) & (!g2577) & (g1253)) + ((g832) & (g2577) & (g1253)));
	assign g1254 = (((!g34) & (!g36) & (!reset) & (g352) & (!g1253)) + ((!g34) & (!g36) & (!reset) & (g352) & (g1253)) + ((!g34) & (g36) & (!reset) & (!g352) & (g1253)) + ((!g34) & (g36) & (!reset) & (g352) & (g1253)) + ((g34) & (!g36) & (!reset) & (g352) & (!g1253)) + ((g34) & (!g36) & (!reset) & (g352) & (g1253)) + ((g34) & (g36) & (!reset) & (g352) & (!g1253)) + ((g34) & (g36) & (!reset) & (g352) & (g1253)));
	assign g7483 = (((!g832) & (g2580) & (!g1255)) + ((!g832) & (g2580) & (g1255)) + ((g832) & (!g2580) & (g1255)) + ((g832) & (g2580) & (g1255)));
	assign g1256 = (((!g34) & (!g36) & (!reset) & (g353) & (!g1255)) + ((!g34) & (!g36) & (!reset) & (g353) & (g1255)) + ((!g34) & (g36) & (!reset) & (!g353) & (g1255)) + ((!g34) & (g36) & (!reset) & (g353) & (g1255)) + ((g34) & (!g36) & (!reset) & (g353) & (!g1255)) + ((g34) & (!g36) & (!reset) & (g353) & (g1255)) + ((g34) & (g36) & (!reset) & (g353) & (!g1255)) + ((g34) & (g36) & (!reset) & (g353) & (g1255)));
	assign g7484 = (((!g832) & (g2583) & (!g1257)) + ((!g832) & (g2583) & (g1257)) + ((g832) & (!g2583) & (g1257)) + ((g832) & (g2583) & (g1257)));
	assign g1258 = (((!g34) & (!g36) & (!reset) & (g354) & (!g1257)) + ((!g34) & (!g36) & (!reset) & (g354) & (g1257)) + ((!g34) & (g36) & (!reset) & (!g354) & (g1257)) + ((!g34) & (g36) & (!reset) & (g354) & (g1257)) + ((g34) & (!g36) & (!reset) & (g354) & (!g1257)) + ((g34) & (!g36) & (!reset) & (g354) & (g1257)) + ((g34) & (g36) & (!reset) & (g354) & (!g1257)) + ((g34) & (g36) & (!reset) & (g354) & (g1257)));
	assign g7485 = (((!g832) & (g2586) & (!g1259)) + ((!g832) & (g2586) & (g1259)) + ((g832) & (!g2586) & (g1259)) + ((g832) & (g2586) & (g1259)));
	assign g1260 = (((!g34) & (!g36) & (!reset) & (g355) & (!g1259)) + ((!g34) & (!g36) & (!reset) & (g355) & (g1259)) + ((!g34) & (g36) & (!reset) & (!g355) & (g1259)) + ((!g34) & (g36) & (!reset) & (g355) & (g1259)) + ((g34) & (!g36) & (!reset) & (g355) & (!g1259)) + ((g34) & (!g36) & (!reset) & (g355) & (g1259)) + ((g34) & (g36) & (!reset) & (g355) & (!g1259)) + ((g34) & (g36) & (!reset) & (g355) & (g1259)));
	assign g7486 = (((!g832) & (g2588) & (!g1261)) + ((!g832) & (g2588) & (g1261)) + ((g832) & (!g2588) & (g1261)) + ((g832) & (g2588) & (g1261)));
	assign g1262 = (((!g34) & (!g36) & (!reset) & (g357) & (!g1261)) + ((!g34) & (!g36) & (!reset) & (g357) & (g1261)) + ((!g34) & (g36) & (!reset) & (!g357) & (g1261)) + ((!g34) & (g36) & (!reset) & (g357) & (g1261)) + ((g34) & (!g36) & (!reset) & (g357) & (!g1261)) + ((g34) & (!g36) & (!reset) & (g357) & (g1261)) + ((g34) & (g36) & (!reset) & (g357) & (!g1261)) + ((g34) & (g36) & (!reset) & (g357) & (g1261)));
	assign g7487 = (((!g832) & (g2591) & (!g1263)) + ((!g832) & (g2591) & (g1263)) + ((g832) & (!g2591) & (g1263)) + ((g832) & (g2591) & (g1263)));
	assign g1264 = (((!g34) & (!g36) & (!reset) & (g358) & (!g1263)) + ((!g34) & (!g36) & (!reset) & (g358) & (g1263)) + ((!g34) & (g36) & (!reset) & (!g358) & (g1263)) + ((!g34) & (g36) & (!reset) & (g358) & (g1263)) + ((g34) & (!g36) & (!reset) & (g358) & (!g1263)) + ((g34) & (!g36) & (!reset) & (g358) & (g1263)) + ((g34) & (g36) & (!reset) & (g358) & (!g1263)) + ((g34) & (g36) & (!reset) & (g358) & (g1263)));
	assign g7488 = (((!g832) & (g2594) & (!g1265)) + ((!g832) & (g2594) & (g1265)) + ((g832) & (!g2594) & (g1265)) + ((g832) & (g2594) & (g1265)));
	assign g1266 = (((!g34) & (!g36) & (!reset) & (g359) & (!g1265)) + ((!g34) & (!g36) & (!reset) & (g359) & (g1265)) + ((!g34) & (g36) & (!reset) & (!g359) & (g1265)) + ((!g34) & (g36) & (!reset) & (g359) & (g1265)) + ((g34) & (!g36) & (!reset) & (g359) & (!g1265)) + ((g34) & (!g36) & (!reset) & (g359) & (g1265)) + ((g34) & (g36) & (!reset) & (g359) & (!g1265)) + ((g34) & (g36) & (!reset) & (g359) & (g1265)));
	assign g7489 = (((!g832) & (g2597) & (!g1267)) + ((!g832) & (g2597) & (g1267)) + ((g832) & (!g2597) & (g1267)) + ((g832) & (g2597) & (g1267)));
	assign g1268 = (((!g34) & (!g36) & (!reset) & (g360) & (!g1267)) + ((!g34) & (!g36) & (!reset) & (g360) & (g1267)) + ((!g34) & (g36) & (!reset) & (!g360) & (g1267)) + ((!g34) & (g36) & (!reset) & (g360) & (g1267)) + ((g34) & (!g36) & (!reset) & (g360) & (!g1267)) + ((g34) & (!g36) & (!reset) & (g360) & (g1267)) + ((g34) & (g36) & (!reset) & (g360) & (!g1267)) + ((g34) & (g36) & (!reset) & (g360) & (g1267)));
	assign g7490 = (((!g2017) & (g2604) & (!g1269)) + ((!g2017) & (g2604) & (g1269)) + ((g2017) & (!g2604) & (g1269)) + ((g2017) & (g2604) & (g1269)));
	assign g1270 = (((!g317) & (!g340) & (!g1199) & (!g1236) & (!g1201) & (!g1202)) + ((!g317) & (!g340) & (!g1199) & (!g1236) & (!g1201) & (g1202)) + ((!g317) & (!g340) & (!g1199) & (!g1236) & (g1201) & (!g1202)) + ((!g317) & (!g340) & (!g1199) & (!g1236) & (g1201) & (g1202)) + ((!g317) & (!g340) & (!g1199) & (g1236) & (!g1201) & (!g1202)) + ((!g317) & (!g340) & (!g1199) & (g1236) & (!g1201) & (g1202)) + ((!g317) & (!g340) & (!g1199) & (g1236) & (g1201) & (!g1202)) + ((!g317) & (!g340) & (!g1199) & (g1236) & (g1201) & (g1202)) + ((!g317) & (!g340) & (g1199) & (!g1236) & (!g1201) & (!g1202)) + ((!g317) & (!g340) & (g1199) & (!g1236) & (!g1201) & (g1202)) + ((!g317) & (!g340) & (g1199) & (!g1236) & (g1201) & (!g1202)) + ((!g317) & (!g340) & (g1199) & (!g1236) & (g1201) & (g1202)) + ((!g317) & (!g340) & (g1199) & (g1236) & (!g1201) & (!g1202)) + ((!g317) & (g340) & (!g1199) & (!g1236) & (!g1201) & (!g1202)) + ((!g317) & (g340) & (!g1199) & (!g1236) & (!g1201) & (g1202)) + ((!g317) & (g340) & (!g1199) & (!g1236) & (g1201) & (!g1202)) + ((!g317) & (g340) & (!g1199) & (!g1236) & (g1201) & (g1202)) + ((!g317) & (g340) & (g1199) & (!g1236) & (!g1201) & (!g1202)) + ((g317) & (!g340) & (!g1199) & (!g1236) & (!g1201) & (!g1202)) + ((g317) & (!g340) & (!g1199) & (!g1236) & (!g1201) & (g1202)) + ((g317) & (!g340) & (!g1199) & (!g1236) & (g1201) & (!g1202)) + ((g317) & (!g340) & (!g1199) & (!g1236) & (g1201) & (g1202)) + ((g317) & (!g340) & (!g1199) & (g1236) & (!g1201) & (!g1202)) + ((g317) & (!g340) & (g1199) & (!g1236) & (!g1201) & (!g1202)) + ((g317) & (!g340) & (g1199) & (!g1236) & (!g1201) & (g1202)) + ((g317) & (!g340) & (g1199) & (!g1236) & (g1201) & (!g1202)) + ((g317) & (!g340) & (g1199) & (!g1236) & (g1201) & (g1202)) + ((g317) & (g340) & (!g1199) & (!g1236) & (!g1201) & (!g1202)));
	assign g1271 = (((!g827) & (!g363) & (g1269) & (!g1270)) + ((!g827) & (!g363) & (g1269) & (g1270)) + ((!g827) & (g363) & (g1269) & (!g1270)) + ((!g827) & (g363) & (g1269) & (g1270)) + ((g827) & (!g363) & (!g1269) & (!g1270)) + ((g827) & (!g363) & (g1269) & (g1270)) + ((g827) & (g363) & (!g1269) & (g1270)) + ((g827) & (g363) & (g1269) & (!g1270)));
	assign g1272 = (((!g34) & (!g36) & (!reset) & (g365) & (!g386)) + ((!g34) & (!g36) & (!reset) & (g365) & (g386)) + ((!g34) & (g36) & (!reset) & (!g365) & (g386)) + ((!g34) & (g36) & (!reset) & (g365) & (g386)) + ((g34) & (!g36) & (!reset) & (g365) & (!g386)) + ((g34) & (!g36) & (!reset) & (g365) & (g386)) + ((g34) & (g36) & (!reset) & (g365) & (!g386)) + ((g34) & (g36) & (!reset) & (g365) & (g386)));
	assign g7491 = (((!g832) & (g2606) & (!g1273)) + ((!g832) & (g2606) & (g1273)) + ((g832) & (!g2606) & (g1273)) + ((g832) & (g2606) & (g1273)));
	assign g1274 = (((!g34) & (!g36) & (!reset) & (g366) & (!g1273)) + ((!g34) & (!g36) & (!reset) & (g366) & (g1273)) + ((!g34) & (g36) & (!reset) & (!g366) & (g1273)) + ((!g34) & (g36) & (!reset) & (g366) & (g1273)) + ((g34) & (!g36) & (!reset) & (g366) & (!g1273)) + ((g34) & (!g36) & (!reset) & (g366) & (g1273)) + ((g34) & (g36) & (!reset) & (g366) & (!g1273)) + ((g34) & (g36) & (!reset) & (g366) & (g1273)));
	assign g7492 = (((!g832) & (g2609) & (!g1275)) + ((!g832) & (g2609) & (g1275)) + ((g832) & (!g2609) & (g1275)) + ((g832) & (g2609) & (g1275)));
	assign g1276 = (((!g34) & (!g36) & (!reset) & (g367) & (!g1275)) + ((!g34) & (!g36) & (!reset) & (g367) & (g1275)) + ((!g34) & (g36) & (!reset) & (!g367) & (g1275)) + ((!g34) & (g36) & (!reset) & (g367) & (g1275)) + ((g34) & (!g36) & (!reset) & (g367) & (!g1275)) + ((g34) & (!g36) & (!reset) & (g367) & (g1275)) + ((g34) & (g36) & (!reset) & (g367) & (!g1275)) + ((g34) & (g36) & (!reset) & (g367) & (g1275)));
	assign g7493 = (((!g832) & (g2611) & (!g1277)) + ((!g832) & (g2611) & (g1277)) + ((g832) & (!g2611) & (g1277)) + ((g832) & (g2611) & (g1277)));
	assign g1278 = (((!g34) & (!g36) & (!reset) & (g368) & (!g1277)) + ((!g34) & (!g36) & (!reset) & (g368) & (g1277)) + ((!g34) & (g36) & (!reset) & (!g368) & (g1277)) + ((!g34) & (g36) & (!reset) & (g368) & (g1277)) + ((g34) & (!g36) & (!reset) & (g368) & (!g1277)) + ((g34) & (!g36) & (!reset) & (g368) & (g1277)) + ((g34) & (g36) & (!reset) & (g368) & (!g1277)) + ((g34) & (g36) & (!reset) & (g368) & (g1277)));
	assign g7494 = (((!g832) & (g2613) & (!g1279)) + ((!g832) & (g2613) & (g1279)) + ((g832) & (!g2613) & (g1279)) + ((g832) & (g2613) & (g1279)));
	assign g1280 = (((!g34) & (!g36) & (!reset) & (g370) & (!g1279)) + ((!g34) & (!g36) & (!reset) & (g370) & (g1279)) + ((!g34) & (g36) & (!reset) & (!g370) & (g1279)) + ((!g34) & (g36) & (!reset) & (g370) & (g1279)) + ((g34) & (!g36) & (!reset) & (g370) & (!g1279)) + ((g34) & (!g36) & (!reset) & (g370) & (g1279)) + ((g34) & (g36) & (!reset) & (g370) & (!g1279)) + ((g34) & (g36) & (!reset) & (g370) & (g1279)));
	assign g7495 = (((!g832) & (g2616) & (!g1281)) + ((!g832) & (g2616) & (g1281)) + ((g832) & (!g2616) & (g1281)) + ((g832) & (g2616) & (g1281)));
	assign g1282 = (((!g34) & (!g36) & (!reset) & (g371) & (!g1281)) + ((!g34) & (!g36) & (!reset) & (g371) & (g1281)) + ((!g34) & (g36) & (!reset) & (!g371) & (g1281)) + ((!g34) & (g36) & (!reset) & (g371) & (g1281)) + ((g34) & (!g36) & (!reset) & (g371) & (!g1281)) + ((g34) & (!g36) & (!reset) & (g371) & (g1281)) + ((g34) & (g36) & (!reset) & (g371) & (!g1281)) + ((g34) & (g36) & (!reset) & (g371) & (g1281)));
	assign g7496 = (((!g832) & (g2619) & (!g1283)) + ((!g832) & (g2619) & (g1283)) + ((g832) & (!g2619) & (g1283)) + ((g832) & (g2619) & (g1283)));
	assign g1284 = (((!g34) & (!g36) & (!reset) & (g372) & (!g1283)) + ((!g34) & (!g36) & (!reset) & (g372) & (g1283)) + ((!g34) & (g36) & (!reset) & (!g372) & (g1283)) + ((!g34) & (g36) & (!reset) & (g372) & (g1283)) + ((g34) & (!g36) & (!reset) & (g372) & (!g1283)) + ((g34) & (!g36) & (!reset) & (g372) & (g1283)) + ((g34) & (g36) & (!reset) & (g372) & (!g1283)) + ((g34) & (g36) & (!reset) & (g372) & (g1283)));
	assign g7497 = (((!g832) & (g2622) & (!g1285)) + ((!g832) & (g2622) & (g1285)) + ((g832) & (!g2622) & (g1285)) + ((g832) & (g2622) & (g1285)));
	assign g1286 = (((!g34) & (!g36) & (!reset) & (g373) & (!g1285)) + ((!g34) & (!g36) & (!reset) & (g373) & (g1285)) + ((!g34) & (g36) & (!reset) & (!g373) & (g1285)) + ((!g34) & (g36) & (!reset) & (g373) & (g1285)) + ((g34) & (!g36) & (!reset) & (g373) & (!g1285)) + ((g34) & (!g36) & (!reset) & (g373) & (g1285)) + ((g34) & (g36) & (!reset) & (g373) & (!g1285)) + ((g34) & (g36) & (!reset) & (g373) & (g1285)));
	assign g7498 = (((!g832) & (g2625) & (!g1287)) + ((!g832) & (g2625) & (g1287)) + ((g832) & (!g2625) & (g1287)) + ((g832) & (g2625) & (g1287)));
	assign g1288 = (((!g34) & (!g36) & (!reset) & (g375) & (!g1287)) + ((!g34) & (!g36) & (!reset) & (g375) & (g1287)) + ((!g34) & (g36) & (!reset) & (!g375) & (g1287)) + ((!g34) & (g36) & (!reset) & (g375) & (g1287)) + ((g34) & (!g36) & (!reset) & (g375) & (!g1287)) + ((g34) & (!g36) & (!reset) & (g375) & (g1287)) + ((g34) & (g36) & (!reset) & (g375) & (!g1287)) + ((g34) & (g36) & (!reset) & (g375) & (g1287)));
	assign g7499 = (((!g832) & (g2628) & (!g1289)) + ((!g832) & (g2628) & (g1289)) + ((g832) & (!g2628) & (g1289)) + ((g832) & (g2628) & (g1289)));
	assign g1290 = (((!g34) & (!g36) & (!reset) & (g376) & (!g1289)) + ((!g34) & (!g36) & (!reset) & (g376) & (g1289)) + ((!g34) & (g36) & (!reset) & (!g376) & (g1289)) + ((!g34) & (g36) & (!reset) & (g376) & (g1289)) + ((g34) & (!g36) & (!reset) & (g376) & (!g1289)) + ((g34) & (!g36) & (!reset) & (g376) & (g1289)) + ((g34) & (g36) & (!reset) & (g376) & (!g1289)) + ((g34) & (g36) & (!reset) & (g376) & (g1289)));
	assign g7500 = (((!g832) & (g2631) & (!g1291)) + ((!g832) & (g2631) & (g1291)) + ((g832) & (!g2631) & (g1291)) + ((g832) & (g2631) & (g1291)));
	assign g1292 = (((!g34) & (!g36) & (!reset) & (g377) & (!g1291)) + ((!g34) & (!g36) & (!reset) & (g377) & (g1291)) + ((!g34) & (g36) & (!reset) & (!g377) & (g1291)) + ((!g34) & (g36) & (!reset) & (g377) & (g1291)) + ((g34) & (!g36) & (!reset) & (g377) & (!g1291)) + ((g34) & (!g36) & (!reset) & (g377) & (g1291)) + ((g34) & (g36) & (!reset) & (g377) & (!g1291)) + ((g34) & (g36) & (!reset) & (g377) & (g1291)));
	assign g7501 = (((!g832) & (g2634) & (!g1293)) + ((!g832) & (g2634) & (g1293)) + ((g832) & (!g2634) & (g1293)) + ((g832) & (g2634) & (g1293)));
	assign g1294 = (((!g34) & (!g36) & (!reset) & (g378) & (!g1293)) + ((!g34) & (!g36) & (!reset) & (g378) & (g1293)) + ((!g34) & (g36) & (!reset) & (!g378) & (g1293)) + ((!g34) & (g36) & (!reset) & (g378) & (g1293)) + ((g34) & (!g36) & (!reset) & (g378) & (!g1293)) + ((g34) & (!g36) & (!reset) & (g378) & (g1293)) + ((g34) & (g36) & (!reset) & (g378) & (!g1293)) + ((g34) & (g36) & (!reset) & (g378) & (g1293)));
	assign g7502 = (((!g832) & (g2636) & (!g1295)) + ((!g832) & (g2636) & (g1295)) + ((g832) & (!g2636) & (g1295)) + ((g832) & (g2636) & (g1295)));
	assign g1296 = (((!g34) & (!g36) & (!reset) & (g380) & (!g1295)) + ((!g34) & (!g36) & (!reset) & (g380) & (g1295)) + ((!g34) & (g36) & (!reset) & (!g380) & (g1295)) + ((!g34) & (g36) & (!reset) & (g380) & (g1295)) + ((g34) & (!g36) & (!reset) & (g380) & (!g1295)) + ((g34) & (!g36) & (!reset) & (g380) & (g1295)) + ((g34) & (g36) & (!reset) & (g380) & (!g1295)) + ((g34) & (g36) & (!reset) & (g380) & (g1295)));
	assign g7503 = (((!g832) & (g2639) & (!g1297)) + ((!g832) & (g2639) & (g1297)) + ((g832) & (!g2639) & (g1297)) + ((g832) & (g2639) & (g1297)));
	assign g1298 = (((!g34) & (!g36) & (!reset) & (g381) & (!g1297)) + ((!g34) & (!g36) & (!reset) & (g381) & (g1297)) + ((!g34) & (g36) & (!reset) & (!g381) & (g1297)) + ((!g34) & (g36) & (!reset) & (g381) & (g1297)) + ((g34) & (!g36) & (!reset) & (g381) & (!g1297)) + ((g34) & (!g36) & (!reset) & (g381) & (g1297)) + ((g34) & (g36) & (!reset) & (g381) & (!g1297)) + ((g34) & (g36) & (!reset) & (g381) & (g1297)));
	assign g7504 = (((!g832) & (g2642) & (!g1299)) + ((!g832) & (g2642) & (g1299)) + ((g832) & (!g2642) & (g1299)) + ((g832) & (g2642) & (g1299)));
	assign g1300 = (((!g34) & (!g36) & (!reset) & (g382) & (!g1299)) + ((!g34) & (!g36) & (!reset) & (g382) & (g1299)) + ((!g34) & (g36) & (!reset) & (!g382) & (g1299)) + ((!g34) & (g36) & (!reset) & (g382) & (g1299)) + ((g34) & (!g36) & (!reset) & (g382) & (!g1299)) + ((g34) & (!g36) & (!reset) & (g382) & (g1299)) + ((g34) & (g36) & (!reset) & (g382) & (!g1299)) + ((g34) & (g36) & (!reset) & (g382) & (g1299)));
	assign g7505 = (((!g832) & (g2645) & (!g1301)) + ((!g832) & (g2645) & (g1301)) + ((g832) & (!g2645) & (g1301)) + ((g832) & (g2645) & (g1301)));
	assign g1302 = (((!g34) & (!g36) & (!reset) & (g383) & (!g1301)) + ((!g34) & (!g36) & (!reset) & (g383) & (g1301)) + ((!g34) & (g36) & (!reset) & (!g383) & (g1301)) + ((!g34) & (g36) & (!reset) & (g383) & (g1301)) + ((g34) & (!g36) & (!reset) & (g383) & (!g1301)) + ((g34) & (!g36) & (!reset) & (g383) & (g1301)) + ((g34) & (g36) & (!reset) & (g383) & (!g1301)) + ((g34) & (g36) & (!reset) & (g383) & (g1301)));
	assign g7506 = (((!g2017) & (g7126) & (!g1303)) + ((!g2017) & (g7126) & (g1303)) + ((g2017) & (!g7126) & (g1303)) + ((g2017) & (g7126) & (g1303)));
	assign g1304 = (((!g363) & (g1269) & (!g1270)) + ((g363) & (!g1269) & (!g1270)) + ((g363) & (g1269) & (!g1270)) + ((g363) & (g1269) & (g1270)));
	assign g1305 = (((!g827) & (!g386) & (g1303) & (!g1304)) + ((!g827) & (!g386) & (g1303) & (g1304)) + ((!g827) & (g386) & (g1303) & (!g1304)) + ((!g827) & (g386) & (g1303) & (g1304)) + ((g827) & (!g386) & (!g1303) & (g1304)) + ((g827) & (!g386) & (g1303) & (!g1304)) + ((g827) & (g386) & (!g1303) & (!g1304)) + ((g827) & (g386) & (g1303) & (g1304)));
	assign g1306 = (((!g34) & (!g36) & (!reset) & (g388) & (!g409)) + ((!g34) & (!g36) & (!reset) & (g388) & (g409)) + ((!g34) & (g36) & (!reset) & (!g388) & (g409)) + ((!g34) & (g36) & (!reset) & (g388) & (g409)) + ((g34) & (!g36) & (!reset) & (g388) & (!g409)) + ((g34) & (!g36) & (!reset) & (g388) & (g409)) + ((g34) & (g36) & (!reset) & (g388) & (!g409)) + ((g34) & (g36) & (!reset) & (g388) & (g409)));
	assign g7507 = (((!g832) & (g2652) & (!g1307)) + ((!g832) & (g2652) & (g1307)) + ((g832) & (!g2652) & (g1307)) + ((g832) & (g2652) & (g1307)));
	assign g1308 = (((!g34) & (!g36) & (!reset) & (g389) & (!g1307)) + ((!g34) & (!g36) & (!reset) & (g389) & (g1307)) + ((!g34) & (g36) & (!reset) & (!g389) & (g1307)) + ((!g34) & (g36) & (!reset) & (g389) & (g1307)) + ((g34) & (!g36) & (!reset) & (g389) & (!g1307)) + ((g34) & (!g36) & (!reset) & (g389) & (g1307)) + ((g34) & (g36) & (!reset) & (g389) & (!g1307)) + ((g34) & (g36) & (!reset) & (g389) & (g1307)));
	assign g7508 = (((!g832) & (g2654) & (!g1309)) + ((!g832) & (g2654) & (g1309)) + ((g832) & (!g2654) & (g1309)) + ((g832) & (g2654) & (g1309)));
	assign g1310 = (((!g34) & (!g36) & (!reset) & (g390) & (!g1309)) + ((!g34) & (!g36) & (!reset) & (g390) & (g1309)) + ((!g34) & (g36) & (!reset) & (!g390) & (g1309)) + ((!g34) & (g36) & (!reset) & (g390) & (g1309)) + ((g34) & (!g36) & (!reset) & (g390) & (!g1309)) + ((g34) & (!g36) & (!reset) & (g390) & (g1309)) + ((g34) & (g36) & (!reset) & (g390) & (!g1309)) + ((g34) & (g36) & (!reset) & (g390) & (g1309)));
	assign g7509 = (((!g832) & (g2655) & (!g1311)) + ((!g832) & (g2655) & (g1311)) + ((g832) & (!g2655) & (g1311)) + ((g832) & (g2655) & (g1311)));
	assign g1312 = (((!g34) & (!g36) & (!reset) & (g391) & (!g1311)) + ((!g34) & (!g36) & (!reset) & (g391) & (g1311)) + ((!g34) & (g36) & (!reset) & (!g391) & (g1311)) + ((!g34) & (g36) & (!reset) & (g391) & (g1311)) + ((g34) & (!g36) & (!reset) & (g391) & (!g1311)) + ((g34) & (!g36) & (!reset) & (g391) & (g1311)) + ((g34) & (g36) & (!reset) & (g391) & (!g1311)) + ((g34) & (g36) & (!reset) & (g391) & (g1311)));
	assign g7510 = (((!g832) & (g2656) & (!g1313)) + ((!g832) & (g2656) & (g1313)) + ((g832) & (!g2656) & (g1313)) + ((g832) & (g2656) & (g1313)));
	assign g1314 = (((!g34) & (!g36) & (!reset) & (g393) & (!g1313)) + ((!g34) & (!g36) & (!reset) & (g393) & (g1313)) + ((!g34) & (g36) & (!reset) & (!g393) & (g1313)) + ((!g34) & (g36) & (!reset) & (g393) & (g1313)) + ((g34) & (!g36) & (!reset) & (g393) & (!g1313)) + ((g34) & (!g36) & (!reset) & (g393) & (g1313)) + ((g34) & (g36) & (!reset) & (g393) & (!g1313)) + ((g34) & (g36) & (!reset) & (g393) & (g1313)));
	assign g7511 = (((!g832) & (g2658) & (!g1315)) + ((!g832) & (g2658) & (g1315)) + ((g832) & (!g2658) & (g1315)) + ((g832) & (g2658) & (g1315)));
	assign g1316 = (((!g34) & (!g36) & (!reset) & (g394) & (!g1315)) + ((!g34) & (!g36) & (!reset) & (g394) & (g1315)) + ((!g34) & (g36) & (!reset) & (!g394) & (g1315)) + ((!g34) & (g36) & (!reset) & (g394) & (g1315)) + ((g34) & (!g36) & (!reset) & (g394) & (!g1315)) + ((g34) & (!g36) & (!reset) & (g394) & (g1315)) + ((g34) & (g36) & (!reset) & (g394) & (!g1315)) + ((g34) & (g36) & (!reset) & (g394) & (g1315)));
	assign g7512 = (((!g832) & (g2660) & (!g1317)) + ((!g832) & (g2660) & (g1317)) + ((g832) & (!g2660) & (g1317)) + ((g832) & (g2660) & (g1317)));
	assign g1318 = (((!g34) & (!g36) & (!reset) & (g395) & (!g1317)) + ((!g34) & (!g36) & (!reset) & (g395) & (g1317)) + ((!g34) & (g36) & (!reset) & (!g395) & (g1317)) + ((!g34) & (g36) & (!reset) & (g395) & (g1317)) + ((g34) & (!g36) & (!reset) & (g395) & (!g1317)) + ((g34) & (!g36) & (!reset) & (g395) & (g1317)) + ((g34) & (g36) & (!reset) & (g395) & (!g1317)) + ((g34) & (g36) & (!reset) & (g395) & (g1317)));
	assign g7513 = (((!g832) & (g2662) & (!g1319)) + ((!g832) & (g2662) & (g1319)) + ((g832) & (!g2662) & (g1319)) + ((g832) & (g2662) & (g1319)));
	assign g1320 = (((!g34) & (!g36) & (!reset) & (g396) & (!g1319)) + ((!g34) & (!g36) & (!reset) & (g396) & (g1319)) + ((!g34) & (g36) & (!reset) & (!g396) & (g1319)) + ((!g34) & (g36) & (!reset) & (g396) & (g1319)) + ((g34) & (!g36) & (!reset) & (g396) & (!g1319)) + ((g34) & (!g36) & (!reset) & (g396) & (g1319)) + ((g34) & (g36) & (!reset) & (g396) & (!g1319)) + ((g34) & (g36) & (!reset) & (g396) & (g1319)));
	assign g7514 = (((!g832) & (g2664) & (!g1321)) + ((!g832) & (g2664) & (g1321)) + ((g832) & (!g2664) & (g1321)) + ((g832) & (g2664) & (g1321)));
	assign g1322 = (((!g34) & (!g36) & (!reset) & (g398) & (!g1321)) + ((!g34) & (!g36) & (!reset) & (g398) & (g1321)) + ((!g34) & (g36) & (!reset) & (!g398) & (g1321)) + ((!g34) & (g36) & (!reset) & (g398) & (g1321)) + ((g34) & (!g36) & (!reset) & (g398) & (!g1321)) + ((g34) & (!g36) & (!reset) & (g398) & (g1321)) + ((g34) & (g36) & (!reset) & (g398) & (!g1321)) + ((g34) & (g36) & (!reset) & (g398) & (g1321)));
	assign g7515 = (((!g832) & (g2666) & (!g1323)) + ((!g832) & (g2666) & (g1323)) + ((g832) & (!g2666) & (g1323)) + ((g832) & (g2666) & (g1323)));
	assign g1324 = (((!g34) & (!g36) & (!reset) & (g399) & (!g1323)) + ((!g34) & (!g36) & (!reset) & (g399) & (g1323)) + ((!g34) & (g36) & (!reset) & (!g399) & (g1323)) + ((!g34) & (g36) & (!reset) & (g399) & (g1323)) + ((g34) & (!g36) & (!reset) & (g399) & (!g1323)) + ((g34) & (!g36) & (!reset) & (g399) & (g1323)) + ((g34) & (g36) & (!reset) & (g399) & (!g1323)) + ((g34) & (g36) & (!reset) & (g399) & (g1323)));
	assign g7516 = (((!g832) & (g2668) & (!g1325)) + ((!g832) & (g2668) & (g1325)) + ((g832) & (!g2668) & (g1325)) + ((g832) & (g2668) & (g1325)));
	assign g1326 = (((!g34) & (!g36) & (!reset) & (g400) & (!g1325)) + ((!g34) & (!g36) & (!reset) & (g400) & (g1325)) + ((!g34) & (g36) & (!reset) & (!g400) & (g1325)) + ((!g34) & (g36) & (!reset) & (g400) & (g1325)) + ((g34) & (!g36) & (!reset) & (g400) & (!g1325)) + ((g34) & (!g36) & (!reset) & (g400) & (g1325)) + ((g34) & (g36) & (!reset) & (g400) & (!g1325)) + ((g34) & (g36) & (!reset) & (g400) & (g1325)));
	assign g7517 = (((!g832) & (g2670) & (!g1327)) + ((!g832) & (g2670) & (g1327)) + ((g832) & (!g2670) & (g1327)) + ((g832) & (g2670) & (g1327)));
	assign g1328 = (((!g34) & (!g36) & (!reset) & (g401) & (!g1327)) + ((!g34) & (!g36) & (!reset) & (g401) & (g1327)) + ((!g34) & (g36) & (!reset) & (!g401) & (g1327)) + ((!g34) & (g36) & (!reset) & (g401) & (g1327)) + ((g34) & (!g36) & (!reset) & (g401) & (!g1327)) + ((g34) & (!g36) & (!reset) & (g401) & (g1327)) + ((g34) & (g36) & (!reset) & (g401) & (!g1327)) + ((g34) & (g36) & (!reset) & (g401) & (g1327)));
	assign g7518 = (((!g832) & (g2671) & (!g1329)) + ((!g832) & (g2671) & (g1329)) + ((g832) & (!g2671) & (g1329)) + ((g832) & (g2671) & (g1329)));
	assign g1330 = (((!g34) & (!g36) & (!reset) & (g403) & (!g1329)) + ((!g34) & (!g36) & (!reset) & (g403) & (g1329)) + ((!g34) & (g36) & (!reset) & (!g403) & (g1329)) + ((!g34) & (g36) & (!reset) & (g403) & (g1329)) + ((g34) & (!g36) & (!reset) & (g403) & (!g1329)) + ((g34) & (!g36) & (!reset) & (g403) & (g1329)) + ((g34) & (g36) & (!reset) & (g403) & (!g1329)) + ((g34) & (g36) & (!reset) & (g403) & (g1329)));
	assign g7519 = (((!g832) & (g2673) & (!g1331)) + ((!g832) & (g2673) & (g1331)) + ((g832) & (!g2673) & (g1331)) + ((g832) & (g2673) & (g1331)));
	assign g1332 = (((!g34) & (!g36) & (!reset) & (g404) & (!g1331)) + ((!g34) & (!g36) & (!reset) & (g404) & (g1331)) + ((!g34) & (g36) & (!reset) & (!g404) & (g1331)) + ((!g34) & (g36) & (!reset) & (g404) & (g1331)) + ((g34) & (!g36) & (!reset) & (g404) & (!g1331)) + ((g34) & (!g36) & (!reset) & (g404) & (g1331)) + ((g34) & (g36) & (!reset) & (g404) & (!g1331)) + ((g34) & (g36) & (!reset) & (g404) & (g1331)));
	assign g7520 = (((!g832) & (g2675) & (!g1333)) + ((!g832) & (g2675) & (g1333)) + ((g832) & (!g2675) & (g1333)) + ((g832) & (g2675) & (g1333)));
	assign g1334 = (((!g34) & (!g36) & (!reset) & (g405) & (!g1333)) + ((!g34) & (!g36) & (!reset) & (g405) & (g1333)) + ((!g34) & (g36) & (!reset) & (!g405) & (g1333)) + ((!g34) & (g36) & (!reset) & (g405) & (g1333)) + ((g34) & (!g36) & (!reset) & (g405) & (!g1333)) + ((g34) & (!g36) & (!reset) & (g405) & (g1333)) + ((g34) & (g36) & (!reset) & (g405) & (!g1333)) + ((g34) & (g36) & (!reset) & (g405) & (g1333)));
	assign g7521 = (((!g832) & (g2677) & (!g1335)) + ((!g832) & (g2677) & (g1335)) + ((g832) & (!g2677) & (g1335)) + ((g832) & (g2677) & (g1335)));
	assign g1336 = (((!g34) & (!g36) & (!reset) & (g406) & (!g1335)) + ((!g34) & (!g36) & (!reset) & (g406) & (g1335)) + ((!g34) & (g36) & (!reset) & (!g406) & (g1335)) + ((!g34) & (g36) & (!reset) & (g406) & (g1335)) + ((g34) & (!g36) & (!reset) & (g406) & (!g1335)) + ((g34) & (!g36) & (!reset) & (g406) & (g1335)) + ((g34) & (g36) & (!reset) & (g406) & (!g1335)) + ((g34) & (g36) & (!reset) & (g406) & (g1335)));
	assign g7522 = (((!g2017) & (g2685) & (!g1337)) + ((!g2017) & (g2685) & (g1337)) + ((g2017) & (!g2685) & (g1337)) + ((g2017) & (g2685) & (g1337)));
	assign g1338 = (((!g827) & (!g386) & (!g409) & (!g1303) & (g1337) & (!g1304)) + ((!g827) & (!g386) & (!g409) & (!g1303) & (g1337) & (g1304)) + ((!g827) & (!g386) & (!g409) & (g1303) & (g1337) & (!g1304)) + ((!g827) & (!g386) & (!g409) & (g1303) & (g1337) & (g1304)) + ((!g827) & (!g386) & (g409) & (!g1303) & (g1337) & (!g1304)) + ((!g827) & (!g386) & (g409) & (!g1303) & (g1337) & (g1304)) + ((!g827) & (!g386) & (g409) & (g1303) & (g1337) & (!g1304)) + ((!g827) & (!g386) & (g409) & (g1303) & (g1337) & (g1304)) + ((!g827) & (g386) & (!g409) & (!g1303) & (g1337) & (!g1304)) + ((!g827) & (g386) & (!g409) & (!g1303) & (g1337) & (g1304)) + ((!g827) & (g386) & (!g409) & (g1303) & (g1337) & (!g1304)) + ((!g827) & (g386) & (!g409) & (g1303) & (g1337) & (g1304)) + ((!g827) & (g386) & (g409) & (!g1303) & (g1337) & (!g1304)) + ((!g827) & (g386) & (g409) & (!g1303) & (g1337) & (g1304)) + ((!g827) & (g386) & (g409) & (g1303) & (g1337) & (!g1304)) + ((!g827) & (g386) & (g409) & (g1303) & (g1337) & (g1304)) + ((g827) & (!g386) & (!g409) & (!g1303) & (g1337) & (!g1304)) + ((g827) & (!g386) & (!g409) & (!g1303) & (g1337) & (g1304)) + ((g827) & (!g386) & (!g409) & (g1303) & (!g1337) & (g1304)) + ((g827) & (!g386) & (!g409) & (g1303) & (g1337) & (!g1304)) + ((g827) & (!g386) & (g409) & (!g1303) & (!g1337) & (!g1304)) + ((g827) & (!g386) & (g409) & (!g1303) & (!g1337) & (g1304)) + ((g827) & (!g386) & (g409) & (g1303) & (!g1337) & (!g1304)) + ((g827) & (!g386) & (g409) & (g1303) & (g1337) & (g1304)) + ((g827) & (g386) & (!g409) & (!g1303) & (!g1337) & (g1304)) + ((g827) & (g386) & (!g409) & (!g1303) & (g1337) & (!g1304)) + ((g827) & (g386) & (!g409) & (g1303) & (!g1337) & (!g1304)) + ((g827) & (g386) & (!g409) & (g1303) & (!g1337) & (g1304)) + ((g827) & (g386) & (g409) & (!g1303) & (!g1337) & (!g1304)) + ((g827) & (g386) & (g409) & (!g1303) & (g1337) & (g1304)) + ((g827) & (g386) & (g409) & (g1303) & (g1337) & (!g1304)) + ((g827) & (g386) & (g409) & (g1303) & (g1337) & (g1304)));
	assign g1339 = (((!g34) & (!g36) & (!reset) & (g411) & (!g432)) + ((!g34) & (!g36) & (!reset) & (g411) & (g432)) + ((!g34) & (g36) & (!reset) & (!g411) & (g432)) + ((!g34) & (g36) & (!reset) & (g411) & (g432)) + ((g34) & (!g36) & (!reset) & (g411) & (!g432)) + ((g34) & (!g36) & (!reset) & (g411) & (g432)) + ((g34) & (g36) & (!reset) & (g411) & (!g432)) + ((g34) & (g36) & (!reset) & (g411) & (g432)));
	assign g7523 = (((!g832) & (g2689) & (!g1340)) + ((!g832) & (g2689) & (g1340)) + ((g832) & (!g2689) & (g1340)) + ((g832) & (g2689) & (g1340)));
	assign g1341 = (((!g34) & (!g36) & (!reset) & (g412) & (!g1340)) + ((!g34) & (!g36) & (!reset) & (g412) & (g1340)) + ((!g34) & (g36) & (!reset) & (!g412) & (g1340)) + ((!g34) & (g36) & (!reset) & (g412) & (g1340)) + ((g34) & (!g36) & (!reset) & (g412) & (!g1340)) + ((g34) & (!g36) & (!reset) & (g412) & (g1340)) + ((g34) & (g36) & (!reset) & (g412) & (!g1340)) + ((g34) & (g36) & (!reset) & (g412) & (g1340)));
	assign g7524 = (((!g832) & (g2694) & (!g1342)) + ((!g832) & (g2694) & (g1342)) + ((g832) & (!g2694) & (g1342)) + ((g832) & (g2694) & (g1342)));
	assign g1343 = (((!g34) & (!g36) & (!reset) & (g413) & (!g1342)) + ((!g34) & (!g36) & (!reset) & (g413) & (g1342)) + ((!g34) & (g36) & (!reset) & (!g413) & (g1342)) + ((!g34) & (g36) & (!reset) & (g413) & (g1342)) + ((g34) & (!g36) & (!reset) & (g413) & (!g1342)) + ((g34) & (!g36) & (!reset) & (g413) & (g1342)) + ((g34) & (g36) & (!reset) & (g413) & (!g1342)) + ((g34) & (g36) & (!reset) & (g413) & (g1342)));
	assign g7525 = (((!g832) & (g2698) & (!g1344)) + ((!g832) & (g2698) & (g1344)) + ((g832) & (!g2698) & (g1344)) + ((g832) & (g2698) & (g1344)));
	assign g1345 = (((!g34) & (!g36) & (!reset) & (g414) & (!g1344)) + ((!g34) & (!g36) & (!reset) & (g414) & (g1344)) + ((!g34) & (g36) & (!reset) & (!g414) & (g1344)) + ((!g34) & (g36) & (!reset) & (g414) & (g1344)) + ((g34) & (!g36) & (!reset) & (g414) & (!g1344)) + ((g34) & (!g36) & (!reset) & (g414) & (g1344)) + ((g34) & (g36) & (!reset) & (g414) & (!g1344)) + ((g34) & (g36) & (!reset) & (g414) & (g1344)));
	assign g7526 = (((!g832) & (g2702) & (!g1346)) + ((!g832) & (g2702) & (g1346)) + ((g832) & (!g2702) & (g1346)) + ((g832) & (g2702) & (g1346)));
	assign g1347 = (((!g34) & (!g36) & (!reset) & (g416) & (!g1346)) + ((!g34) & (!g36) & (!reset) & (g416) & (g1346)) + ((!g34) & (g36) & (!reset) & (!g416) & (g1346)) + ((!g34) & (g36) & (!reset) & (g416) & (g1346)) + ((g34) & (!g36) & (!reset) & (g416) & (!g1346)) + ((g34) & (!g36) & (!reset) & (g416) & (g1346)) + ((g34) & (g36) & (!reset) & (g416) & (!g1346)) + ((g34) & (g36) & (!reset) & (g416) & (g1346)));
	assign g7527 = (((!g832) & (g2707) & (!g1348)) + ((!g832) & (g2707) & (g1348)) + ((g832) & (!g2707) & (g1348)) + ((g832) & (g2707) & (g1348)));
	assign g1349 = (((!g34) & (!g36) & (!reset) & (g417) & (!g1348)) + ((!g34) & (!g36) & (!reset) & (g417) & (g1348)) + ((!g34) & (g36) & (!reset) & (!g417) & (g1348)) + ((!g34) & (g36) & (!reset) & (g417) & (g1348)) + ((g34) & (!g36) & (!reset) & (g417) & (!g1348)) + ((g34) & (!g36) & (!reset) & (g417) & (g1348)) + ((g34) & (g36) & (!reset) & (g417) & (!g1348)) + ((g34) & (g36) & (!reset) & (g417) & (g1348)));
	assign g7528 = (((!g832) & (g2712) & (!g1350)) + ((!g832) & (g2712) & (g1350)) + ((g832) & (!g2712) & (g1350)) + ((g832) & (g2712) & (g1350)));
	assign g1351 = (((!g34) & (!g36) & (!reset) & (g418) & (!g1350)) + ((!g34) & (!g36) & (!reset) & (g418) & (g1350)) + ((!g34) & (g36) & (!reset) & (!g418) & (g1350)) + ((!g34) & (g36) & (!reset) & (g418) & (g1350)) + ((g34) & (!g36) & (!reset) & (g418) & (!g1350)) + ((g34) & (!g36) & (!reset) & (g418) & (g1350)) + ((g34) & (g36) & (!reset) & (g418) & (!g1350)) + ((g34) & (g36) & (!reset) & (g418) & (g1350)));
	assign g7529 = (((!g832) & (g2717) & (!g1352)) + ((!g832) & (g2717) & (g1352)) + ((g832) & (!g2717) & (g1352)) + ((g832) & (g2717) & (g1352)));
	assign g1353 = (((!g34) & (!g36) & (!reset) & (g419) & (!g1352)) + ((!g34) & (!g36) & (!reset) & (g419) & (g1352)) + ((!g34) & (g36) & (!reset) & (!g419) & (g1352)) + ((!g34) & (g36) & (!reset) & (g419) & (g1352)) + ((g34) & (!g36) & (!reset) & (g419) & (!g1352)) + ((g34) & (!g36) & (!reset) & (g419) & (g1352)) + ((g34) & (g36) & (!reset) & (g419) & (!g1352)) + ((g34) & (g36) & (!reset) & (g419) & (g1352)));
	assign g7530 = (((!g832) & (g2722) & (!g1354)) + ((!g832) & (g2722) & (g1354)) + ((g832) & (!g2722) & (g1354)) + ((g832) & (g2722) & (g1354)));
	assign g1355 = (((!g34) & (!g36) & (!reset) & (g421) & (!g1354)) + ((!g34) & (!g36) & (!reset) & (g421) & (g1354)) + ((!g34) & (g36) & (!reset) & (!g421) & (g1354)) + ((!g34) & (g36) & (!reset) & (g421) & (g1354)) + ((g34) & (!g36) & (!reset) & (g421) & (!g1354)) + ((g34) & (!g36) & (!reset) & (g421) & (g1354)) + ((g34) & (g36) & (!reset) & (g421) & (!g1354)) + ((g34) & (g36) & (!reset) & (g421) & (g1354)));
	assign g7531 = (((!g832) & (g2727) & (!g1356)) + ((!g832) & (g2727) & (g1356)) + ((g832) & (!g2727) & (g1356)) + ((g832) & (g2727) & (g1356)));
	assign g1357 = (((!g34) & (!g36) & (!reset) & (g422) & (!g1356)) + ((!g34) & (!g36) & (!reset) & (g422) & (g1356)) + ((!g34) & (g36) & (!reset) & (!g422) & (g1356)) + ((!g34) & (g36) & (!reset) & (g422) & (g1356)) + ((g34) & (!g36) & (!reset) & (g422) & (!g1356)) + ((g34) & (!g36) & (!reset) & (g422) & (g1356)) + ((g34) & (g36) & (!reset) & (g422) & (!g1356)) + ((g34) & (g36) & (!reset) & (g422) & (g1356)));
	assign g7532 = (((!g832) & (g2732) & (!g1358)) + ((!g832) & (g2732) & (g1358)) + ((g832) & (!g2732) & (g1358)) + ((g832) & (g2732) & (g1358)));
	assign g1359 = (((!g34) & (!g36) & (!reset) & (g423) & (!g1358)) + ((!g34) & (!g36) & (!reset) & (g423) & (g1358)) + ((!g34) & (g36) & (!reset) & (!g423) & (g1358)) + ((!g34) & (g36) & (!reset) & (g423) & (g1358)) + ((g34) & (!g36) & (!reset) & (g423) & (!g1358)) + ((g34) & (!g36) & (!reset) & (g423) & (g1358)) + ((g34) & (g36) & (!reset) & (g423) & (!g1358)) + ((g34) & (g36) & (!reset) & (g423) & (g1358)));
	assign g7533 = (((!g832) & (g2737) & (!g1360)) + ((!g832) & (g2737) & (g1360)) + ((g832) & (!g2737) & (g1360)) + ((g832) & (g2737) & (g1360)));
	assign g1361 = (((!g34) & (!g36) & (!reset) & (g424) & (!g1360)) + ((!g34) & (!g36) & (!reset) & (g424) & (g1360)) + ((!g34) & (g36) & (!reset) & (!g424) & (g1360)) + ((!g34) & (g36) & (!reset) & (g424) & (g1360)) + ((g34) & (!g36) & (!reset) & (g424) & (!g1360)) + ((g34) & (!g36) & (!reset) & (g424) & (g1360)) + ((g34) & (g36) & (!reset) & (g424) & (!g1360)) + ((g34) & (g36) & (!reset) & (g424) & (g1360)));
	assign g7534 = (((!g832) & (g2741) & (!g1362)) + ((!g832) & (g2741) & (g1362)) + ((g832) & (!g2741) & (g1362)) + ((g832) & (g2741) & (g1362)));
	assign g1363 = (((!g34) & (!g36) & (!reset) & (g426) & (!g1362)) + ((!g34) & (!g36) & (!reset) & (g426) & (g1362)) + ((!g34) & (g36) & (!reset) & (!g426) & (g1362)) + ((!g34) & (g36) & (!reset) & (g426) & (g1362)) + ((g34) & (!g36) & (!reset) & (g426) & (!g1362)) + ((g34) & (!g36) & (!reset) & (g426) & (g1362)) + ((g34) & (g36) & (!reset) & (g426) & (!g1362)) + ((g34) & (g36) & (!reset) & (g426) & (g1362)));
	assign g7535 = (((!g832) & (g2746) & (!g1364)) + ((!g832) & (g2746) & (g1364)) + ((g832) & (!g2746) & (g1364)) + ((g832) & (g2746) & (g1364)));
	assign g1365 = (((!g34) & (!g36) & (!reset) & (g427) & (!g1364)) + ((!g34) & (!g36) & (!reset) & (g427) & (g1364)) + ((!g34) & (g36) & (!reset) & (!g427) & (g1364)) + ((!g34) & (g36) & (!reset) & (g427) & (g1364)) + ((g34) & (!g36) & (!reset) & (g427) & (!g1364)) + ((g34) & (!g36) & (!reset) & (g427) & (g1364)) + ((g34) & (g36) & (!reset) & (g427) & (!g1364)) + ((g34) & (g36) & (!reset) & (g427) & (g1364)));
	assign g7536 = (((!g832) & (g2751) & (!g1366)) + ((!g832) & (g2751) & (g1366)) + ((g832) & (!g2751) & (g1366)) + ((g832) & (g2751) & (g1366)));
	assign g1367 = (((!g34) & (!g36) & (!reset) & (g428) & (!g1366)) + ((!g34) & (!g36) & (!reset) & (g428) & (g1366)) + ((!g34) & (g36) & (!reset) & (!g428) & (g1366)) + ((!g34) & (g36) & (!reset) & (g428) & (g1366)) + ((g34) & (!g36) & (!reset) & (g428) & (!g1366)) + ((g34) & (!g36) & (!reset) & (g428) & (g1366)) + ((g34) & (g36) & (!reset) & (g428) & (!g1366)) + ((g34) & (g36) & (!reset) & (g428) & (g1366)));
	assign g7537 = (((!g832) & (g2756) & (!g1368)) + ((!g832) & (g2756) & (g1368)) + ((g832) & (!g2756) & (g1368)) + ((g832) & (g2756) & (g1368)));
	assign g1369 = (((!g34) & (!g36) & (!reset) & (g429) & (!g1368)) + ((!g34) & (!g36) & (!reset) & (g429) & (g1368)) + ((!g34) & (g36) & (!reset) & (!g429) & (g1368)) + ((!g34) & (g36) & (!reset) & (g429) & (g1368)) + ((g34) & (!g36) & (!reset) & (g429) & (!g1368)) + ((g34) & (!g36) & (!reset) & (g429) & (g1368)) + ((g34) & (g36) & (!reset) & (g429) & (!g1368)) + ((g34) & (g36) & (!reset) & (g429) & (g1368)));
	assign g7538 = (((!g2017) & (g2762) & (!g1370)) + ((!g2017) & (g2762) & (g1370)) + ((g2017) & (!g2762) & (g1370)) + ((g2017) & (g2762) & (g1370)));
	assign g1371 = (((!g317) & (!g1199) & (!g1201) & (!g1202) & (!g5721) & (g5722)) + ((!g317) & (!g1199) & (!g1201) & (g1202) & (!g5721) & (g5722)) + ((!g317) & (!g1199) & (g1201) & (!g1202) & (!g5721) & (g5722)) + ((!g317) & (!g1199) & (g1201) & (g1202) & (!g5721) & (g5722)) + ((!g317) & (g1199) & (!g1201) & (!g1202) & (!g5721) & (g5722)) + ((!g317) & (g1199) & (!g1201) & (g1202) & (!g5721) & (g5722)) + ((!g317) & (g1199) & (!g1201) & (g1202) & (g5721) & (g5722)) + ((!g317) & (g1199) & (g1201) & (!g1202) & (!g5721) & (g5722)) + ((!g317) & (g1199) & (g1201) & (!g1202) & (g5721) & (g5722)) + ((!g317) & (g1199) & (g1201) & (g1202) & (!g5721) & (g5722)) + ((!g317) & (g1199) & (g1201) & (g1202) & (g5721) & (g5722)) + ((g317) & (!g1199) & (!g1201) & (!g1202) & (!g5721) & (g5722)) + ((g317) & (!g1199) & (!g1201) & (g1202) & (!g5721) & (g5722)) + ((g317) & (!g1199) & (!g1201) & (g1202) & (g5721) & (g5722)) + ((g317) & (!g1199) & (g1201) & (!g1202) & (!g5721) & (g5722)) + ((g317) & (!g1199) & (g1201) & (!g1202) & (g5721) & (g5722)) + ((g317) & (!g1199) & (g1201) & (g1202) & (!g5721) & (g5722)) + ((g317) & (!g1199) & (g1201) & (g1202) & (g5721) & (g5722)) + ((g317) & (g1199) & (!g1201) & (!g1202) & (!g5721) & (g5722)) + ((g317) & (g1199) & (!g1201) & (!g1202) & (g5721) & (g5722)) + ((g317) & (g1199) & (!g1201) & (g1202) & (!g5721) & (g5722)) + ((g317) & (g1199) & (!g1201) & (g1202) & (g5721) & (g5722)) + ((g317) & (g1199) & (g1201) & (!g1202) & (!g5721) & (g5722)) + ((g317) & (g1199) & (g1201) & (!g1202) & (g5721) & (g5722)) + ((g317) & (g1199) & (g1201) & (g1202) & (!g5721) & (g5722)) + ((g317) & (g1199) & (g1201) & (g1202) & (g5721) & (g5722)));
	assign g1372 = (((g409) & (g1337)));
	assign g1373 = (((!g1371) & (!g1372)));
	assign g1374 = (((!g827) & (!g432) & (g1370) & (!g1373)) + ((!g827) & (!g432) & (g1370) & (g1373)) + ((!g827) & (g432) & (g1370) & (!g1373)) + ((!g827) & (g432) & (g1370) & (g1373)) + ((g827) & (!g432) & (!g1370) & (!g1373)) + ((g827) & (!g432) & (g1370) & (g1373)) + ((g827) & (g432) & (!g1370) & (g1373)) + ((g827) & (g432) & (g1370) & (!g1373)));
	assign g1375 = (((!g34) & (!g36) & (!reset) & (g434) & (!g455)) + ((!g34) & (!g36) & (!reset) & (g434) & (g455)) + ((!g34) & (g36) & (!reset) & (!g434) & (g455)) + ((!g34) & (g36) & (!reset) & (g434) & (g455)) + ((g34) & (!g36) & (!reset) & (g434) & (!g455)) + ((g34) & (!g36) & (!reset) & (g434) & (g455)) + ((g34) & (g36) & (!reset) & (g434) & (!g455)) + ((g34) & (g36) & (!reset) & (g434) & (g455)));
	assign g7539 = (((!g832) & (g2763) & (!g1376)) + ((!g832) & (g2763) & (g1376)) + ((g832) & (!g2763) & (g1376)) + ((g832) & (g2763) & (g1376)));
	assign g1377 = (((!g34) & (!g36) & (!reset) & (g435) & (!g1376)) + ((!g34) & (!g36) & (!reset) & (g435) & (g1376)) + ((!g34) & (g36) & (!reset) & (!g435) & (g1376)) + ((!g34) & (g36) & (!reset) & (g435) & (g1376)) + ((g34) & (!g36) & (!reset) & (g435) & (!g1376)) + ((g34) & (!g36) & (!reset) & (g435) & (g1376)) + ((g34) & (g36) & (!reset) & (g435) & (!g1376)) + ((g34) & (g36) & (!reset) & (g435) & (g1376)));
	assign g7540 = (((!g832) & (g2765) & (!g1378)) + ((!g832) & (g2765) & (g1378)) + ((g832) & (!g2765) & (g1378)) + ((g832) & (g2765) & (g1378)));
	assign g1379 = (((!g34) & (!g36) & (!reset) & (g436) & (!g1378)) + ((!g34) & (!g36) & (!reset) & (g436) & (g1378)) + ((!g34) & (g36) & (!reset) & (!g436) & (g1378)) + ((!g34) & (g36) & (!reset) & (g436) & (g1378)) + ((g34) & (!g36) & (!reset) & (g436) & (!g1378)) + ((g34) & (!g36) & (!reset) & (g436) & (g1378)) + ((g34) & (g36) & (!reset) & (g436) & (!g1378)) + ((g34) & (g36) & (!reset) & (g436) & (g1378)));
	assign g7541 = (((!g832) & (g2766) & (!g1380)) + ((!g832) & (g2766) & (g1380)) + ((g832) & (!g2766) & (g1380)) + ((g832) & (g2766) & (g1380)));
	assign g1381 = (((!g34) & (!g36) & (!reset) & (g437) & (!g1380)) + ((!g34) & (!g36) & (!reset) & (g437) & (g1380)) + ((!g34) & (g36) & (!reset) & (!g437) & (g1380)) + ((!g34) & (g36) & (!reset) & (g437) & (g1380)) + ((g34) & (!g36) & (!reset) & (g437) & (!g1380)) + ((g34) & (!g36) & (!reset) & (g437) & (g1380)) + ((g34) & (g36) & (!reset) & (g437) & (!g1380)) + ((g34) & (g36) & (!reset) & (g437) & (g1380)));
	assign g7542 = (((!g832) & (g2767) & (!g1382)) + ((!g832) & (g2767) & (g1382)) + ((g832) & (!g2767) & (g1382)) + ((g832) & (g2767) & (g1382)));
	assign g1383 = (((!g34) & (!g36) & (!reset) & (g439) & (!g1382)) + ((!g34) & (!g36) & (!reset) & (g439) & (g1382)) + ((!g34) & (g36) & (!reset) & (!g439) & (g1382)) + ((!g34) & (g36) & (!reset) & (g439) & (g1382)) + ((g34) & (!g36) & (!reset) & (g439) & (!g1382)) + ((g34) & (!g36) & (!reset) & (g439) & (g1382)) + ((g34) & (g36) & (!reset) & (g439) & (!g1382)) + ((g34) & (g36) & (!reset) & (g439) & (g1382)));
	assign g7543 = (((!g832) & (g2769) & (!g1384)) + ((!g832) & (g2769) & (g1384)) + ((g832) & (!g2769) & (g1384)) + ((g832) & (g2769) & (g1384)));
	assign g1385 = (((!g34) & (!g36) & (!reset) & (g440) & (!g1384)) + ((!g34) & (!g36) & (!reset) & (g440) & (g1384)) + ((!g34) & (g36) & (!reset) & (!g440) & (g1384)) + ((!g34) & (g36) & (!reset) & (g440) & (g1384)) + ((g34) & (!g36) & (!reset) & (g440) & (!g1384)) + ((g34) & (!g36) & (!reset) & (g440) & (g1384)) + ((g34) & (g36) & (!reset) & (g440) & (!g1384)) + ((g34) & (g36) & (!reset) & (g440) & (g1384)));
	assign g7544 = (((!g832) & (g2771) & (!g1386)) + ((!g832) & (g2771) & (g1386)) + ((g832) & (!g2771) & (g1386)) + ((g832) & (g2771) & (g1386)));
	assign g1387 = (((!g34) & (!g36) & (!reset) & (g441) & (!g1386)) + ((!g34) & (!g36) & (!reset) & (g441) & (g1386)) + ((!g34) & (g36) & (!reset) & (!g441) & (g1386)) + ((!g34) & (g36) & (!reset) & (g441) & (g1386)) + ((g34) & (!g36) & (!reset) & (g441) & (!g1386)) + ((g34) & (!g36) & (!reset) & (g441) & (g1386)) + ((g34) & (g36) & (!reset) & (g441) & (!g1386)) + ((g34) & (g36) & (!reset) & (g441) & (g1386)));
	assign g7545 = (((!g832) & (g2773) & (!g1388)) + ((!g832) & (g2773) & (g1388)) + ((g832) & (!g2773) & (g1388)) + ((g832) & (g2773) & (g1388)));
	assign g1389 = (((!g34) & (!g36) & (!reset) & (g442) & (!g1388)) + ((!g34) & (!g36) & (!reset) & (g442) & (g1388)) + ((!g34) & (g36) & (!reset) & (!g442) & (g1388)) + ((!g34) & (g36) & (!reset) & (g442) & (g1388)) + ((g34) & (!g36) & (!reset) & (g442) & (!g1388)) + ((g34) & (!g36) & (!reset) & (g442) & (g1388)) + ((g34) & (g36) & (!reset) & (g442) & (!g1388)) + ((g34) & (g36) & (!reset) & (g442) & (g1388)));
	assign g7546 = (((!g832) & (g2775) & (!g1390)) + ((!g832) & (g2775) & (g1390)) + ((g832) & (!g2775) & (g1390)) + ((g832) & (g2775) & (g1390)));
	assign g1391 = (((!g34) & (!g36) & (!reset) & (g444) & (!g1390)) + ((!g34) & (!g36) & (!reset) & (g444) & (g1390)) + ((!g34) & (g36) & (!reset) & (!g444) & (g1390)) + ((!g34) & (g36) & (!reset) & (g444) & (g1390)) + ((g34) & (!g36) & (!reset) & (g444) & (!g1390)) + ((g34) & (!g36) & (!reset) & (g444) & (g1390)) + ((g34) & (g36) & (!reset) & (g444) & (!g1390)) + ((g34) & (g36) & (!reset) & (g444) & (g1390)));
	assign g7547 = (((!g832) & (g2777) & (!g1392)) + ((!g832) & (g2777) & (g1392)) + ((g832) & (!g2777) & (g1392)) + ((g832) & (g2777) & (g1392)));
	assign g1393 = (((!g34) & (!g36) & (!reset) & (g445) & (!g1392)) + ((!g34) & (!g36) & (!reset) & (g445) & (g1392)) + ((!g34) & (g36) & (!reset) & (!g445) & (g1392)) + ((!g34) & (g36) & (!reset) & (g445) & (g1392)) + ((g34) & (!g36) & (!reset) & (g445) & (!g1392)) + ((g34) & (!g36) & (!reset) & (g445) & (g1392)) + ((g34) & (g36) & (!reset) & (g445) & (!g1392)) + ((g34) & (g36) & (!reset) & (g445) & (g1392)));
	assign g7548 = (((!g832) & (g2779) & (!g1394)) + ((!g832) & (g2779) & (g1394)) + ((g832) & (!g2779) & (g1394)) + ((g832) & (g2779) & (g1394)));
	assign g1395 = (((!g34) & (!g36) & (!reset) & (g446) & (!g1394)) + ((!g34) & (!g36) & (!reset) & (g446) & (g1394)) + ((!g34) & (g36) & (!reset) & (!g446) & (g1394)) + ((!g34) & (g36) & (!reset) & (g446) & (g1394)) + ((g34) & (!g36) & (!reset) & (g446) & (!g1394)) + ((g34) & (!g36) & (!reset) & (g446) & (g1394)) + ((g34) & (g36) & (!reset) & (g446) & (!g1394)) + ((g34) & (g36) & (!reset) & (g446) & (g1394)));
	assign g7549 = (((!g832) & (g2781) & (!g1396)) + ((!g832) & (g2781) & (g1396)) + ((g832) & (!g2781) & (g1396)) + ((g832) & (g2781) & (g1396)));
	assign g1397 = (((!g34) & (!g36) & (!reset) & (g447) & (!g1396)) + ((!g34) & (!g36) & (!reset) & (g447) & (g1396)) + ((!g34) & (g36) & (!reset) & (!g447) & (g1396)) + ((!g34) & (g36) & (!reset) & (g447) & (g1396)) + ((g34) & (!g36) & (!reset) & (g447) & (!g1396)) + ((g34) & (!g36) & (!reset) & (g447) & (g1396)) + ((g34) & (g36) & (!reset) & (g447) & (!g1396)) + ((g34) & (g36) & (!reset) & (g447) & (g1396)));
	assign g7550 = (((!g832) & (g2782) & (!g1398)) + ((!g832) & (g2782) & (g1398)) + ((g832) & (!g2782) & (g1398)) + ((g832) & (g2782) & (g1398)));
	assign g1399 = (((!g34) & (!g36) & (!reset) & (g449) & (!g1398)) + ((!g34) & (!g36) & (!reset) & (g449) & (g1398)) + ((!g34) & (g36) & (!reset) & (!g449) & (g1398)) + ((!g34) & (g36) & (!reset) & (g449) & (g1398)) + ((g34) & (!g36) & (!reset) & (g449) & (!g1398)) + ((g34) & (!g36) & (!reset) & (g449) & (g1398)) + ((g34) & (g36) & (!reset) & (g449) & (!g1398)) + ((g34) & (g36) & (!reset) & (g449) & (g1398)));
	assign g7551 = (((!g832) & (g2784) & (!g1400)) + ((!g832) & (g2784) & (g1400)) + ((g832) & (!g2784) & (g1400)) + ((g832) & (g2784) & (g1400)));
	assign g1401 = (((!g34) & (!g36) & (!reset) & (g450) & (!g1400)) + ((!g34) & (!g36) & (!reset) & (g450) & (g1400)) + ((!g34) & (g36) & (!reset) & (!g450) & (g1400)) + ((!g34) & (g36) & (!reset) & (g450) & (g1400)) + ((g34) & (!g36) & (!reset) & (g450) & (!g1400)) + ((g34) & (!g36) & (!reset) & (g450) & (g1400)) + ((g34) & (g36) & (!reset) & (g450) & (!g1400)) + ((g34) & (g36) & (!reset) & (g450) & (g1400)));
	assign g7552 = (((!g832) & (g2786) & (!g1402)) + ((!g832) & (g2786) & (g1402)) + ((g832) & (!g2786) & (g1402)) + ((g832) & (g2786) & (g1402)));
	assign g1403 = (((!g34) & (!g36) & (!reset) & (g451) & (!g1402)) + ((!g34) & (!g36) & (!reset) & (g451) & (g1402)) + ((!g34) & (g36) & (!reset) & (!g451) & (g1402)) + ((!g34) & (g36) & (!reset) & (g451) & (g1402)) + ((g34) & (!g36) & (!reset) & (g451) & (!g1402)) + ((g34) & (!g36) & (!reset) & (g451) & (g1402)) + ((g34) & (g36) & (!reset) & (g451) & (!g1402)) + ((g34) & (g36) & (!reset) & (g451) & (g1402)));
	assign g7553 = (((!g832) & (g2788) & (!g1404)) + ((!g832) & (g2788) & (g1404)) + ((g832) & (!g2788) & (g1404)) + ((g832) & (g2788) & (g1404)));
	assign g1405 = (((!g34) & (!g36) & (!reset) & (g452) & (!g1404)) + ((!g34) & (!g36) & (!reset) & (g452) & (g1404)) + ((!g34) & (g36) & (!reset) & (!g452) & (g1404)) + ((!g34) & (g36) & (!reset) & (g452) & (g1404)) + ((g34) & (!g36) & (!reset) & (g452) & (!g1404)) + ((g34) & (!g36) & (!reset) & (g452) & (g1404)) + ((g34) & (g36) & (!reset) & (g452) & (!g1404)) + ((g34) & (g36) & (!reset) & (g452) & (g1404)));
	assign g7554 = (((!g2017) & (g7120) & (!g1406)) + ((!g2017) & (g7120) & (g1406)) + ((g2017) & (!g7120) & (g1406)) + ((g2017) & (g7120) & (g1406)));
	assign g1407 = (((!g827) & (!g432) & (!g455) & (!g1370) & (g1406) & (!g1373)) + ((!g827) & (!g432) & (!g455) & (!g1370) & (g1406) & (g1373)) + ((!g827) & (!g432) & (!g455) & (g1370) & (g1406) & (!g1373)) + ((!g827) & (!g432) & (!g455) & (g1370) & (g1406) & (g1373)) + ((!g827) & (!g432) & (g455) & (!g1370) & (g1406) & (!g1373)) + ((!g827) & (!g432) & (g455) & (!g1370) & (g1406) & (g1373)) + ((!g827) & (!g432) & (g455) & (g1370) & (g1406) & (!g1373)) + ((!g827) & (!g432) & (g455) & (g1370) & (g1406) & (g1373)) + ((!g827) & (g432) & (!g455) & (!g1370) & (g1406) & (!g1373)) + ((!g827) & (g432) & (!g455) & (!g1370) & (g1406) & (g1373)) + ((!g827) & (g432) & (!g455) & (g1370) & (g1406) & (!g1373)) + ((!g827) & (g432) & (!g455) & (g1370) & (g1406) & (g1373)) + ((!g827) & (g432) & (g455) & (!g1370) & (g1406) & (!g1373)) + ((!g827) & (g432) & (g455) & (!g1370) & (g1406) & (g1373)) + ((!g827) & (g432) & (g455) & (g1370) & (g1406) & (!g1373)) + ((!g827) & (g432) & (g455) & (g1370) & (g1406) & (g1373)) + ((g827) & (!g432) & (!g455) & (!g1370) & (g1406) & (!g1373)) + ((g827) & (!g432) & (!g455) & (!g1370) & (g1406) & (g1373)) + ((g827) & (!g432) & (!g455) & (g1370) & (!g1406) & (!g1373)) + ((g827) & (!g432) & (!g455) & (g1370) & (g1406) & (g1373)) + ((g827) & (!g432) & (g455) & (!g1370) & (!g1406) & (!g1373)) + ((g827) & (!g432) & (g455) & (!g1370) & (!g1406) & (g1373)) + ((g827) & (!g432) & (g455) & (g1370) & (!g1406) & (g1373)) + ((g827) & (!g432) & (g455) & (g1370) & (g1406) & (!g1373)) + ((g827) & (g432) & (!g455) & (!g1370) & (!g1406) & (!g1373)) + ((g827) & (g432) & (!g455) & (!g1370) & (g1406) & (g1373)) + ((g827) & (g432) & (!g455) & (g1370) & (!g1406) & (!g1373)) + ((g827) & (g432) & (!g455) & (g1370) & (!g1406) & (g1373)) + ((g827) & (g432) & (g455) & (!g1370) & (!g1406) & (g1373)) + ((g827) & (g432) & (g455) & (!g1370) & (g1406) & (!g1373)) + ((g827) & (g432) & (g455) & (g1370) & (g1406) & (!g1373)) + ((g827) & (g432) & (g455) & (g1370) & (g1406) & (g1373)));
	assign g1408 = (((!g34) & (!g36) & (!reset) & (g457) & (!g478)) + ((!g34) & (!g36) & (!reset) & (g457) & (g478)) + ((!g34) & (g36) & (!reset) & (!g457) & (g478)) + ((!g34) & (g36) & (!reset) & (g457) & (g478)) + ((g34) & (!g36) & (!reset) & (g457) & (!g478)) + ((g34) & (!g36) & (!reset) & (g457) & (g478)) + ((g34) & (g36) & (!reset) & (g457) & (!g478)) + ((g34) & (g36) & (!reset) & (g457) & (g478)));
	assign g7555 = (((!g832) & (g2796) & (!g1409)) + ((!g832) & (g2796) & (g1409)) + ((g832) & (!g2796) & (g1409)) + ((g832) & (g2796) & (g1409)));
	assign g1410 = (((!g34) & (!g36) & (!reset) & (g458) & (!g1409)) + ((!g34) & (!g36) & (!reset) & (g458) & (g1409)) + ((!g34) & (g36) & (!reset) & (!g458) & (g1409)) + ((!g34) & (g36) & (!reset) & (g458) & (g1409)) + ((g34) & (!g36) & (!reset) & (g458) & (!g1409)) + ((g34) & (!g36) & (!reset) & (g458) & (g1409)) + ((g34) & (g36) & (!reset) & (g458) & (!g1409)) + ((g34) & (g36) & (!reset) & (g458) & (g1409)));
	assign g7556 = (((!g832) & (g2799) & (!g1411)) + ((!g832) & (g2799) & (g1411)) + ((g832) & (!g2799) & (g1411)) + ((g832) & (g2799) & (g1411)));
	assign g1412 = (((!g34) & (!g36) & (!reset) & (g459) & (!g1411)) + ((!g34) & (!g36) & (!reset) & (g459) & (g1411)) + ((!g34) & (g36) & (!reset) & (!g459) & (g1411)) + ((!g34) & (g36) & (!reset) & (g459) & (g1411)) + ((g34) & (!g36) & (!reset) & (g459) & (!g1411)) + ((g34) & (!g36) & (!reset) & (g459) & (g1411)) + ((g34) & (g36) & (!reset) & (g459) & (!g1411)) + ((g34) & (g36) & (!reset) & (g459) & (g1411)));
	assign g7557 = (((!g832) & (g2801) & (!g1413)) + ((!g832) & (g2801) & (g1413)) + ((g832) & (!g2801) & (g1413)) + ((g832) & (g2801) & (g1413)));
	assign g1414 = (((!g34) & (!g36) & (!reset) & (g460) & (!g1413)) + ((!g34) & (!g36) & (!reset) & (g460) & (g1413)) + ((!g34) & (g36) & (!reset) & (!g460) & (g1413)) + ((!g34) & (g36) & (!reset) & (g460) & (g1413)) + ((g34) & (!g36) & (!reset) & (g460) & (!g1413)) + ((g34) & (!g36) & (!reset) & (g460) & (g1413)) + ((g34) & (g36) & (!reset) & (g460) & (!g1413)) + ((g34) & (g36) & (!reset) & (g460) & (g1413)));
	assign g7558 = (((!g832) & (g2803) & (!g1415)) + ((!g832) & (g2803) & (g1415)) + ((g832) & (!g2803) & (g1415)) + ((g832) & (g2803) & (g1415)));
	assign g1416 = (((!g34) & (!g36) & (!reset) & (g462) & (!g1415)) + ((!g34) & (!g36) & (!reset) & (g462) & (g1415)) + ((!g34) & (g36) & (!reset) & (!g462) & (g1415)) + ((!g34) & (g36) & (!reset) & (g462) & (g1415)) + ((g34) & (!g36) & (!reset) & (g462) & (!g1415)) + ((g34) & (!g36) & (!reset) & (g462) & (g1415)) + ((g34) & (g36) & (!reset) & (g462) & (!g1415)) + ((g34) & (g36) & (!reset) & (g462) & (g1415)));
	assign g7559 = (((!g832) & (g2806) & (!g1417)) + ((!g832) & (g2806) & (g1417)) + ((g832) & (!g2806) & (g1417)) + ((g832) & (g2806) & (g1417)));
	assign g1418 = (((!g34) & (!g36) & (!reset) & (g463) & (!g1417)) + ((!g34) & (!g36) & (!reset) & (g463) & (g1417)) + ((!g34) & (g36) & (!reset) & (!g463) & (g1417)) + ((!g34) & (g36) & (!reset) & (g463) & (g1417)) + ((g34) & (!g36) & (!reset) & (g463) & (!g1417)) + ((g34) & (!g36) & (!reset) & (g463) & (g1417)) + ((g34) & (g36) & (!reset) & (g463) & (!g1417)) + ((g34) & (g36) & (!reset) & (g463) & (g1417)));
	assign g7560 = (((!g832) & (g2809) & (!g1419)) + ((!g832) & (g2809) & (g1419)) + ((g832) & (!g2809) & (g1419)) + ((g832) & (g2809) & (g1419)));
	assign g1420 = (((!g34) & (!g36) & (!reset) & (g464) & (!g1419)) + ((!g34) & (!g36) & (!reset) & (g464) & (g1419)) + ((!g34) & (g36) & (!reset) & (!g464) & (g1419)) + ((!g34) & (g36) & (!reset) & (g464) & (g1419)) + ((g34) & (!g36) & (!reset) & (g464) & (!g1419)) + ((g34) & (!g36) & (!reset) & (g464) & (g1419)) + ((g34) & (g36) & (!reset) & (g464) & (!g1419)) + ((g34) & (g36) & (!reset) & (g464) & (g1419)));
	assign g7561 = (((!g832) & (g2812) & (!g1421)) + ((!g832) & (g2812) & (g1421)) + ((g832) & (!g2812) & (g1421)) + ((g832) & (g2812) & (g1421)));
	assign g1422 = (((!g34) & (!g36) & (!reset) & (g465) & (!g1421)) + ((!g34) & (!g36) & (!reset) & (g465) & (g1421)) + ((!g34) & (g36) & (!reset) & (!g465) & (g1421)) + ((!g34) & (g36) & (!reset) & (g465) & (g1421)) + ((g34) & (!g36) & (!reset) & (g465) & (!g1421)) + ((g34) & (!g36) & (!reset) & (g465) & (g1421)) + ((g34) & (g36) & (!reset) & (g465) & (!g1421)) + ((g34) & (g36) & (!reset) & (g465) & (g1421)));
	assign g7562 = (((!g832) & (g2815) & (!g1423)) + ((!g832) & (g2815) & (g1423)) + ((g832) & (!g2815) & (g1423)) + ((g832) & (g2815) & (g1423)));
	assign g1424 = (((!g34) & (!g36) & (!reset) & (g467) & (!g1423)) + ((!g34) & (!g36) & (!reset) & (g467) & (g1423)) + ((!g34) & (g36) & (!reset) & (!g467) & (g1423)) + ((!g34) & (g36) & (!reset) & (g467) & (g1423)) + ((g34) & (!g36) & (!reset) & (g467) & (!g1423)) + ((g34) & (!g36) & (!reset) & (g467) & (g1423)) + ((g34) & (g36) & (!reset) & (g467) & (!g1423)) + ((g34) & (g36) & (!reset) & (g467) & (g1423)));
	assign g7563 = (((!g832) & (g2818) & (!g1425)) + ((!g832) & (g2818) & (g1425)) + ((g832) & (!g2818) & (g1425)) + ((g832) & (g2818) & (g1425)));
	assign g1426 = (((!g34) & (!g36) & (!reset) & (g468) & (!g1425)) + ((!g34) & (!g36) & (!reset) & (g468) & (g1425)) + ((!g34) & (g36) & (!reset) & (!g468) & (g1425)) + ((!g34) & (g36) & (!reset) & (g468) & (g1425)) + ((g34) & (!g36) & (!reset) & (g468) & (!g1425)) + ((g34) & (!g36) & (!reset) & (g468) & (g1425)) + ((g34) & (g36) & (!reset) & (g468) & (!g1425)) + ((g34) & (g36) & (!reset) & (g468) & (g1425)));
	assign g7564 = (((!g832) & (g2821) & (!g1427)) + ((!g832) & (g2821) & (g1427)) + ((g832) & (!g2821) & (g1427)) + ((g832) & (g2821) & (g1427)));
	assign g1428 = (((!g34) & (!g36) & (!reset) & (g469) & (!g1427)) + ((!g34) & (!g36) & (!reset) & (g469) & (g1427)) + ((!g34) & (g36) & (!reset) & (!g469) & (g1427)) + ((!g34) & (g36) & (!reset) & (g469) & (g1427)) + ((g34) & (!g36) & (!reset) & (g469) & (!g1427)) + ((g34) & (!g36) & (!reset) & (g469) & (g1427)) + ((g34) & (g36) & (!reset) & (g469) & (!g1427)) + ((g34) & (g36) & (!reset) & (g469) & (g1427)));
	assign g7565 = (((!g832) & (g2824) & (!g1429)) + ((!g832) & (g2824) & (g1429)) + ((g832) & (!g2824) & (g1429)) + ((g832) & (g2824) & (g1429)));
	assign g1430 = (((!g34) & (!g36) & (!reset) & (g470) & (!g1429)) + ((!g34) & (!g36) & (!reset) & (g470) & (g1429)) + ((!g34) & (g36) & (!reset) & (!g470) & (g1429)) + ((!g34) & (g36) & (!reset) & (g470) & (g1429)) + ((g34) & (!g36) & (!reset) & (g470) & (!g1429)) + ((g34) & (!g36) & (!reset) & (g470) & (g1429)) + ((g34) & (g36) & (!reset) & (g470) & (!g1429)) + ((g34) & (g36) & (!reset) & (g470) & (g1429)));
	assign g7566 = (((!g832) & (g2826) & (!g1431)) + ((!g832) & (g2826) & (g1431)) + ((g832) & (!g2826) & (g1431)) + ((g832) & (g2826) & (g1431)));
	assign g1432 = (((!g34) & (!g36) & (!reset) & (g472) & (!g1431)) + ((!g34) & (!g36) & (!reset) & (g472) & (g1431)) + ((!g34) & (g36) & (!reset) & (!g472) & (g1431)) + ((!g34) & (g36) & (!reset) & (g472) & (g1431)) + ((g34) & (!g36) & (!reset) & (g472) & (!g1431)) + ((g34) & (!g36) & (!reset) & (g472) & (g1431)) + ((g34) & (g36) & (!reset) & (g472) & (!g1431)) + ((g34) & (g36) & (!reset) & (g472) & (g1431)));
	assign g7567 = (((!g832) & (g2829) & (!g1433)) + ((!g832) & (g2829) & (g1433)) + ((g832) & (!g2829) & (g1433)) + ((g832) & (g2829) & (g1433)));
	assign g1434 = (((!g34) & (!g36) & (!reset) & (g473) & (!g1433)) + ((!g34) & (!g36) & (!reset) & (g473) & (g1433)) + ((!g34) & (g36) & (!reset) & (!g473) & (g1433)) + ((!g34) & (g36) & (!reset) & (g473) & (g1433)) + ((g34) & (!g36) & (!reset) & (g473) & (!g1433)) + ((g34) & (!g36) & (!reset) & (g473) & (g1433)) + ((g34) & (g36) & (!reset) & (g473) & (!g1433)) + ((g34) & (g36) & (!reset) & (g473) & (g1433)));
	assign g7568 = (((!g832) & (g2832) & (!g1435)) + ((!g832) & (g2832) & (g1435)) + ((g832) & (!g2832) & (g1435)) + ((g832) & (g2832) & (g1435)));
	assign g1436 = (((!g34) & (!g36) & (!reset) & (g474) & (!g1435)) + ((!g34) & (!g36) & (!reset) & (g474) & (g1435)) + ((!g34) & (g36) & (!reset) & (!g474) & (g1435)) + ((!g34) & (g36) & (!reset) & (g474) & (g1435)) + ((g34) & (!g36) & (!reset) & (g474) & (!g1435)) + ((g34) & (!g36) & (!reset) & (g474) & (g1435)) + ((g34) & (g36) & (!reset) & (g474) & (!g1435)) + ((g34) & (g36) & (!reset) & (g474) & (g1435)));
	assign g7569 = (((!g832) & (g2835) & (!g1437)) + ((!g832) & (g2835) & (g1437)) + ((g832) & (!g2835) & (g1437)) + ((g832) & (g2835) & (g1437)));
	assign g1438 = (((!g34) & (!g36) & (!reset) & (g475) & (!g1437)) + ((!g34) & (!g36) & (!reset) & (g475) & (g1437)) + ((!g34) & (g36) & (!reset) & (!g475) & (g1437)) + ((!g34) & (g36) & (!reset) & (g475) & (g1437)) + ((g34) & (!g36) & (!reset) & (g475) & (!g1437)) + ((g34) & (!g36) & (!reset) & (g475) & (g1437)) + ((g34) & (g36) & (!reset) & (g475) & (!g1437)) + ((g34) & (g36) & (!reset) & (g475) & (g1437)));
	assign g7570 = (((!g2017) & (g7114) & (!g1439)) + ((!g2017) & (g7114) & (g1439)) + ((g2017) & (!g7114) & (g1439)) + ((g2017) & (g7114) & (g1439)));
	assign g1440 = (((!g432) & (!g455) & (!g1370) & (!g1406) & (!g1371) & (!g1372)) + ((!g432) & (!g455) & (!g1370) & (!g1406) & (!g1371) & (g1372)) + ((!g432) & (!g455) & (!g1370) & (!g1406) & (g1371) & (!g1372)) + ((!g432) & (!g455) & (!g1370) & (!g1406) & (g1371) & (g1372)) + ((!g432) & (!g455) & (!g1370) & (g1406) & (!g1371) & (!g1372)) + ((!g432) & (!g455) & (!g1370) & (g1406) & (!g1371) & (g1372)) + ((!g432) & (!g455) & (!g1370) & (g1406) & (g1371) & (!g1372)) + ((!g432) & (!g455) & (!g1370) & (g1406) & (g1371) & (g1372)) + ((!g432) & (!g455) & (g1370) & (!g1406) & (!g1371) & (!g1372)) + ((!g432) & (!g455) & (g1370) & (!g1406) & (!g1371) & (g1372)) + ((!g432) & (!g455) & (g1370) & (!g1406) & (g1371) & (!g1372)) + ((!g432) & (!g455) & (g1370) & (!g1406) & (g1371) & (g1372)) + ((!g432) & (!g455) & (g1370) & (g1406) & (!g1371) & (!g1372)) + ((!g432) & (g455) & (!g1370) & (!g1406) & (!g1371) & (!g1372)) + ((!g432) & (g455) & (!g1370) & (!g1406) & (!g1371) & (g1372)) + ((!g432) & (g455) & (!g1370) & (!g1406) & (g1371) & (!g1372)) + ((!g432) & (g455) & (!g1370) & (!g1406) & (g1371) & (g1372)) + ((!g432) & (g455) & (g1370) & (!g1406) & (!g1371) & (!g1372)) + ((g432) & (!g455) & (!g1370) & (!g1406) & (!g1371) & (!g1372)) + ((g432) & (!g455) & (!g1370) & (!g1406) & (!g1371) & (g1372)) + ((g432) & (!g455) & (!g1370) & (!g1406) & (g1371) & (!g1372)) + ((g432) & (!g455) & (!g1370) & (!g1406) & (g1371) & (g1372)) + ((g432) & (!g455) & (!g1370) & (g1406) & (!g1371) & (!g1372)) + ((g432) & (!g455) & (g1370) & (!g1406) & (!g1371) & (!g1372)) + ((g432) & (!g455) & (g1370) & (!g1406) & (!g1371) & (g1372)) + ((g432) & (!g455) & (g1370) & (!g1406) & (g1371) & (!g1372)) + ((g432) & (!g455) & (g1370) & (!g1406) & (g1371) & (g1372)) + ((g432) & (g455) & (!g1370) & (!g1406) & (!g1371) & (!g1372)));
	assign g1441 = (((!g827) & (!g478) & (g1439) & (!g1440)) + ((!g827) & (!g478) & (g1439) & (g1440)) + ((!g827) & (g478) & (g1439) & (!g1440)) + ((!g827) & (g478) & (g1439) & (g1440)) + ((g827) & (!g478) & (!g1439) & (!g1440)) + ((g827) & (!g478) & (g1439) & (g1440)) + ((g827) & (g478) & (!g1439) & (g1440)) + ((g827) & (g478) & (g1439) & (!g1440)));
	assign g1442 = (((!g34) & (!g36) & (!reset) & (g480) & (!g501)) + ((!g34) & (!g36) & (!reset) & (g480) & (g501)) + ((!g34) & (g36) & (!reset) & (!g480) & (g501)) + ((!g34) & (g36) & (!reset) & (g480) & (g501)) + ((g34) & (!g36) & (!reset) & (g480) & (!g501)) + ((g34) & (!g36) & (!reset) & (g480) & (g501)) + ((g34) & (g36) & (!reset) & (g480) & (!g501)) + ((g34) & (g36) & (!reset) & (g480) & (g501)));
	assign g7571 = (((!g832) & (g2837) & (!g1443)) + ((!g832) & (g2837) & (g1443)) + ((g832) & (!g2837) & (g1443)) + ((g832) & (g2837) & (g1443)));
	assign g1444 = (((!g34) & (!g36) & (!reset) & (g481) & (!g1443)) + ((!g34) & (!g36) & (!reset) & (g481) & (g1443)) + ((!g34) & (g36) & (!reset) & (!g481) & (g1443)) + ((!g34) & (g36) & (!reset) & (g481) & (g1443)) + ((g34) & (!g36) & (!reset) & (g481) & (!g1443)) + ((g34) & (!g36) & (!reset) & (g481) & (g1443)) + ((g34) & (g36) & (!reset) & (g481) & (!g1443)) + ((g34) & (g36) & (!reset) & (g481) & (g1443)));
	assign g7572 = (((!g832) & (g2840) & (!g1445)) + ((!g832) & (g2840) & (g1445)) + ((g832) & (!g2840) & (g1445)) + ((g832) & (g2840) & (g1445)));
	assign g1446 = (((!g34) & (!g36) & (!reset) & (g482) & (!g1445)) + ((!g34) & (!g36) & (!reset) & (g482) & (g1445)) + ((!g34) & (g36) & (!reset) & (!g482) & (g1445)) + ((!g34) & (g36) & (!reset) & (g482) & (g1445)) + ((g34) & (!g36) & (!reset) & (g482) & (!g1445)) + ((g34) & (!g36) & (!reset) & (g482) & (g1445)) + ((g34) & (g36) & (!reset) & (g482) & (!g1445)) + ((g34) & (g36) & (!reset) & (g482) & (g1445)));
	assign g7573 = (((!g832) & (g2842) & (!g1447)) + ((!g832) & (g2842) & (g1447)) + ((g832) & (!g2842) & (g1447)) + ((g832) & (g2842) & (g1447)));
	assign g1448 = (((!g34) & (!g36) & (!reset) & (g483) & (!g1447)) + ((!g34) & (!g36) & (!reset) & (g483) & (g1447)) + ((!g34) & (g36) & (!reset) & (!g483) & (g1447)) + ((!g34) & (g36) & (!reset) & (g483) & (g1447)) + ((g34) & (!g36) & (!reset) & (g483) & (!g1447)) + ((g34) & (!g36) & (!reset) & (g483) & (g1447)) + ((g34) & (g36) & (!reset) & (g483) & (!g1447)) + ((g34) & (g36) & (!reset) & (g483) & (g1447)));
	assign g7574 = (((!g832) & (g2844) & (!g1449)) + ((!g832) & (g2844) & (g1449)) + ((g832) & (!g2844) & (g1449)) + ((g832) & (g2844) & (g1449)));
	assign g1450 = (((!g34) & (!g36) & (!reset) & (g485) & (!g1449)) + ((!g34) & (!g36) & (!reset) & (g485) & (g1449)) + ((!g34) & (g36) & (!reset) & (!g485) & (g1449)) + ((!g34) & (g36) & (!reset) & (g485) & (g1449)) + ((g34) & (!g36) & (!reset) & (g485) & (!g1449)) + ((g34) & (!g36) & (!reset) & (g485) & (g1449)) + ((g34) & (g36) & (!reset) & (g485) & (!g1449)) + ((g34) & (g36) & (!reset) & (g485) & (g1449)));
	assign g7575 = (((!g832) & (g2847) & (!g1451)) + ((!g832) & (g2847) & (g1451)) + ((g832) & (!g2847) & (g1451)) + ((g832) & (g2847) & (g1451)));
	assign g1452 = (((!g34) & (!g36) & (!reset) & (g486) & (!g1451)) + ((!g34) & (!g36) & (!reset) & (g486) & (g1451)) + ((!g34) & (g36) & (!reset) & (!g486) & (g1451)) + ((!g34) & (g36) & (!reset) & (g486) & (g1451)) + ((g34) & (!g36) & (!reset) & (g486) & (!g1451)) + ((g34) & (!g36) & (!reset) & (g486) & (g1451)) + ((g34) & (g36) & (!reset) & (g486) & (!g1451)) + ((g34) & (g36) & (!reset) & (g486) & (g1451)));
	assign g7576 = (((!g832) & (g2850) & (!g1453)) + ((!g832) & (g2850) & (g1453)) + ((g832) & (!g2850) & (g1453)) + ((g832) & (g2850) & (g1453)));
	assign g1454 = (((!g34) & (!g36) & (!reset) & (g487) & (!g1453)) + ((!g34) & (!g36) & (!reset) & (g487) & (g1453)) + ((!g34) & (g36) & (!reset) & (!g487) & (g1453)) + ((!g34) & (g36) & (!reset) & (g487) & (g1453)) + ((g34) & (!g36) & (!reset) & (g487) & (!g1453)) + ((g34) & (!g36) & (!reset) & (g487) & (g1453)) + ((g34) & (g36) & (!reset) & (g487) & (!g1453)) + ((g34) & (g36) & (!reset) & (g487) & (g1453)));
	assign g7577 = (((!g832) & (g2853) & (!g1455)) + ((!g832) & (g2853) & (g1455)) + ((g832) & (!g2853) & (g1455)) + ((g832) & (g2853) & (g1455)));
	assign g1456 = (((!g34) & (!g36) & (!reset) & (g488) & (!g1455)) + ((!g34) & (!g36) & (!reset) & (g488) & (g1455)) + ((!g34) & (g36) & (!reset) & (!g488) & (g1455)) + ((!g34) & (g36) & (!reset) & (g488) & (g1455)) + ((g34) & (!g36) & (!reset) & (g488) & (!g1455)) + ((g34) & (!g36) & (!reset) & (g488) & (g1455)) + ((g34) & (g36) & (!reset) & (g488) & (!g1455)) + ((g34) & (g36) & (!reset) & (g488) & (g1455)));
	assign g7578 = (((!g832) & (g2856) & (!g1457)) + ((!g832) & (g2856) & (g1457)) + ((g832) & (!g2856) & (g1457)) + ((g832) & (g2856) & (g1457)));
	assign g1458 = (((!g34) & (!g36) & (!reset) & (g490) & (!g1457)) + ((!g34) & (!g36) & (!reset) & (g490) & (g1457)) + ((!g34) & (g36) & (!reset) & (!g490) & (g1457)) + ((!g34) & (g36) & (!reset) & (g490) & (g1457)) + ((g34) & (!g36) & (!reset) & (g490) & (!g1457)) + ((g34) & (!g36) & (!reset) & (g490) & (g1457)) + ((g34) & (g36) & (!reset) & (g490) & (!g1457)) + ((g34) & (g36) & (!reset) & (g490) & (g1457)));
	assign g7579 = (((!g832) & (g2859) & (!g1459)) + ((!g832) & (g2859) & (g1459)) + ((g832) & (!g2859) & (g1459)) + ((g832) & (g2859) & (g1459)));
	assign g1460 = (((!g34) & (!g36) & (!reset) & (g491) & (!g1459)) + ((!g34) & (!g36) & (!reset) & (g491) & (g1459)) + ((!g34) & (g36) & (!reset) & (!g491) & (g1459)) + ((!g34) & (g36) & (!reset) & (g491) & (g1459)) + ((g34) & (!g36) & (!reset) & (g491) & (!g1459)) + ((g34) & (!g36) & (!reset) & (g491) & (g1459)) + ((g34) & (g36) & (!reset) & (g491) & (!g1459)) + ((g34) & (g36) & (!reset) & (g491) & (g1459)));
	assign g7580 = (((!g832) & (g2862) & (!g1461)) + ((!g832) & (g2862) & (g1461)) + ((g832) & (!g2862) & (g1461)) + ((g832) & (g2862) & (g1461)));
	assign g1462 = (((!g34) & (!g36) & (!reset) & (g492) & (!g1461)) + ((!g34) & (!g36) & (!reset) & (g492) & (g1461)) + ((!g34) & (g36) & (!reset) & (!g492) & (g1461)) + ((!g34) & (g36) & (!reset) & (g492) & (g1461)) + ((g34) & (!g36) & (!reset) & (g492) & (!g1461)) + ((g34) & (!g36) & (!reset) & (g492) & (g1461)) + ((g34) & (g36) & (!reset) & (g492) & (!g1461)) + ((g34) & (g36) & (!reset) & (g492) & (g1461)));
	assign g7581 = (((!g832) & (g2865) & (!g1463)) + ((!g832) & (g2865) & (g1463)) + ((g832) & (!g2865) & (g1463)) + ((g832) & (g2865) & (g1463)));
	assign g1464 = (((!g34) & (!g36) & (!reset) & (g493) & (!g1463)) + ((!g34) & (!g36) & (!reset) & (g493) & (g1463)) + ((!g34) & (g36) & (!reset) & (!g493) & (g1463)) + ((!g34) & (g36) & (!reset) & (g493) & (g1463)) + ((g34) & (!g36) & (!reset) & (g493) & (!g1463)) + ((g34) & (!g36) & (!reset) & (g493) & (g1463)) + ((g34) & (g36) & (!reset) & (g493) & (!g1463)) + ((g34) & (g36) & (!reset) & (g493) & (g1463)));
	assign g7582 = (((!g832) & (g2867) & (!g1465)) + ((!g832) & (g2867) & (g1465)) + ((g832) & (!g2867) & (g1465)) + ((g832) & (g2867) & (g1465)));
	assign g1466 = (((!g34) & (!g36) & (!reset) & (g495) & (!g1465)) + ((!g34) & (!g36) & (!reset) & (g495) & (g1465)) + ((!g34) & (g36) & (!reset) & (!g495) & (g1465)) + ((!g34) & (g36) & (!reset) & (g495) & (g1465)) + ((g34) & (!g36) & (!reset) & (g495) & (!g1465)) + ((g34) & (!g36) & (!reset) & (g495) & (g1465)) + ((g34) & (g36) & (!reset) & (g495) & (!g1465)) + ((g34) & (g36) & (!reset) & (g495) & (g1465)));
	assign g7583 = (((!g832) & (g2870) & (!g1467)) + ((!g832) & (g2870) & (g1467)) + ((g832) & (!g2870) & (g1467)) + ((g832) & (g2870) & (g1467)));
	assign g1468 = (((!g34) & (!g36) & (!reset) & (g496) & (!g1467)) + ((!g34) & (!g36) & (!reset) & (g496) & (g1467)) + ((!g34) & (g36) & (!reset) & (!g496) & (g1467)) + ((!g34) & (g36) & (!reset) & (g496) & (g1467)) + ((g34) & (!g36) & (!reset) & (g496) & (!g1467)) + ((g34) & (!g36) & (!reset) & (g496) & (g1467)) + ((g34) & (g36) & (!reset) & (g496) & (!g1467)) + ((g34) & (g36) & (!reset) & (g496) & (g1467)));
	assign g7584 = (((!g832) & (g2873) & (!g1469)) + ((!g832) & (g2873) & (g1469)) + ((g832) & (!g2873) & (g1469)) + ((g832) & (g2873) & (g1469)));
	assign g1470 = (((!g34) & (!g36) & (!reset) & (g497) & (!g1469)) + ((!g34) & (!g36) & (!reset) & (g497) & (g1469)) + ((!g34) & (g36) & (!reset) & (!g497) & (g1469)) + ((!g34) & (g36) & (!reset) & (g497) & (g1469)) + ((g34) & (!g36) & (!reset) & (g497) & (!g1469)) + ((g34) & (!g36) & (!reset) & (g497) & (g1469)) + ((g34) & (g36) & (!reset) & (g497) & (!g1469)) + ((g34) & (g36) & (!reset) & (g497) & (g1469)));
	assign g7585 = (((!g832) & (g2876) & (!g1471)) + ((!g832) & (g2876) & (g1471)) + ((g832) & (!g2876) & (g1471)) + ((g832) & (g2876) & (g1471)));
	assign g1472 = (((!g34) & (!g36) & (!reset) & (g498) & (!g1471)) + ((!g34) & (!g36) & (!reset) & (g498) & (g1471)) + ((!g34) & (g36) & (!reset) & (!g498) & (g1471)) + ((!g34) & (g36) & (!reset) & (g498) & (g1471)) + ((g34) & (!g36) & (!reset) & (g498) & (!g1471)) + ((g34) & (!g36) & (!reset) & (g498) & (g1471)) + ((g34) & (g36) & (!reset) & (g498) & (!g1471)) + ((g34) & (g36) & (!reset) & (g498) & (g1471)));
	assign g7586 = (((!g2017) & (g2879) & (!g1473)) + ((!g2017) & (g2879) & (g1473)) + ((g2017) & (!g2879) & (g1473)) + ((g2017) & (g2879) & (g1473)));
	assign g1474 = (((!g478) & (g1439) & (!g1440)) + ((g478) & (!g1439) & (!g1440)) + ((g478) & (g1439) & (!g1440)) + ((g478) & (g1439) & (g1440)));
	assign g1475 = (((!g827) & (!g501) & (g1473) & (!g1474)) + ((!g827) & (!g501) & (g1473) & (g1474)) + ((!g827) & (g501) & (g1473) & (!g1474)) + ((!g827) & (g501) & (g1473) & (g1474)) + ((g827) & (!g501) & (!g1473) & (g1474)) + ((g827) & (!g501) & (g1473) & (!g1474)) + ((g827) & (g501) & (!g1473) & (!g1474)) + ((g827) & (g501) & (g1473) & (g1474)));
	assign g1476 = (((!g34) & (!g36) & (!reset) & (g503) & (!g524)) + ((!g34) & (!g36) & (!reset) & (g503) & (g524)) + ((!g34) & (g36) & (!reset) & (!g503) & (g524)) + ((!g34) & (g36) & (!reset) & (g503) & (g524)) + ((g34) & (!g36) & (!reset) & (g503) & (!g524)) + ((g34) & (!g36) & (!reset) & (g503) & (g524)) + ((g34) & (g36) & (!reset) & (g503) & (!g524)) + ((g34) & (g36) & (!reset) & (g503) & (g524)));
	assign g7587 = (((!g832) & (g2880) & (!g1477)) + ((!g832) & (g2880) & (g1477)) + ((g832) & (!g2880) & (g1477)) + ((g832) & (g2880) & (g1477)));
	assign g1478 = (((!g34) & (!g36) & (!reset) & (g504) & (!g1477)) + ((!g34) & (!g36) & (!reset) & (g504) & (g1477)) + ((!g34) & (g36) & (!reset) & (!g504) & (g1477)) + ((!g34) & (g36) & (!reset) & (g504) & (g1477)) + ((g34) & (!g36) & (!reset) & (g504) & (!g1477)) + ((g34) & (!g36) & (!reset) & (g504) & (g1477)) + ((g34) & (g36) & (!reset) & (g504) & (!g1477)) + ((g34) & (g36) & (!reset) & (g504) & (g1477)));
	assign g7588 = (((!g832) & (g2882) & (!g1479)) + ((!g832) & (g2882) & (g1479)) + ((g832) & (!g2882) & (g1479)) + ((g832) & (g2882) & (g1479)));
	assign g1480 = (((!g34) & (!g36) & (!reset) & (g505) & (!g1479)) + ((!g34) & (!g36) & (!reset) & (g505) & (g1479)) + ((!g34) & (g36) & (!reset) & (!g505) & (g1479)) + ((!g34) & (g36) & (!reset) & (g505) & (g1479)) + ((g34) & (!g36) & (!reset) & (g505) & (!g1479)) + ((g34) & (!g36) & (!reset) & (g505) & (g1479)) + ((g34) & (g36) & (!reset) & (g505) & (!g1479)) + ((g34) & (g36) & (!reset) & (g505) & (g1479)));
	assign g7589 = (((!g832) & (g2883) & (!g1481)) + ((!g832) & (g2883) & (g1481)) + ((g832) & (!g2883) & (g1481)) + ((g832) & (g2883) & (g1481)));
	assign g1482 = (((!g34) & (!g36) & (!reset) & (g506) & (!g1481)) + ((!g34) & (!g36) & (!reset) & (g506) & (g1481)) + ((!g34) & (g36) & (!reset) & (!g506) & (g1481)) + ((!g34) & (g36) & (!reset) & (g506) & (g1481)) + ((g34) & (!g36) & (!reset) & (g506) & (!g1481)) + ((g34) & (!g36) & (!reset) & (g506) & (g1481)) + ((g34) & (g36) & (!reset) & (g506) & (!g1481)) + ((g34) & (g36) & (!reset) & (g506) & (g1481)));
	assign g7590 = (((!g832) & (g2884) & (!g1483)) + ((!g832) & (g2884) & (g1483)) + ((g832) & (!g2884) & (g1483)) + ((g832) & (g2884) & (g1483)));
	assign g1484 = (((!g34) & (!g36) & (!reset) & (g508) & (!g1483)) + ((!g34) & (!g36) & (!reset) & (g508) & (g1483)) + ((!g34) & (g36) & (!reset) & (!g508) & (g1483)) + ((!g34) & (g36) & (!reset) & (g508) & (g1483)) + ((g34) & (!g36) & (!reset) & (g508) & (!g1483)) + ((g34) & (!g36) & (!reset) & (g508) & (g1483)) + ((g34) & (g36) & (!reset) & (g508) & (!g1483)) + ((g34) & (g36) & (!reset) & (g508) & (g1483)));
	assign g7591 = (((!g832) & (g2886) & (!g1485)) + ((!g832) & (g2886) & (g1485)) + ((g832) & (!g2886) & (g1485)) + ((g832) & (g2886) & (g1485)));
	assign g1486 = (((!g34) & (!g36) & (!reset) & (g509) & (!g1485)) + ((!g34) & (!g36) & (!reset) & (g509) & (g1485)) + ((!g34) & (g36) & (!reset) & (!g509) & (g1485)) + ((!g34) & (g36) & (!reset) & (g509) & (g1485)) + ((g34) & (!g36) & (!reset) & (g509) & (!g1485)) + ((g34) & (!g36) & (!reset) & (g509) & (g1485)) + ((g34) & (g36) & (!reset) & (g509) & (!g1485)) + ((g34) & (g36) & (!reset) & (g509) & (g1485)));
	assign g7592 = (((!g832) & (g2888) & (!g1487)) + ((!g832) & (g2888) & (g1487)) + ((g832) & (!g2888) & (g1487)) + ((g832) & (g2888) & (g1487)));
	assign g1488 = (((!g34) & (!g36) & (!reset) & (g510) & (!g1487)) + ((!g34) & (!g36) & (!reset) & (g510) & (g1487)) + ((!g34) & (g36) & (!reset) & (!g510) & (g1487)) + ((!g34) & (g36) & (!reset) & (g510) & (g1487)) + ((g34) & (!g36) & (!reset) & (g510) & (!g1487)) + ((g34) & (!g36) & (!reset) & (g510) & (g1487)) + ((g34) & (g36) & (!reset) & (g510) & (!g1487)) + ((g34) & (g36) & (!reset) & (g510) & (g1487)));
	assign g7593 = (((!g832) & (g2890) & (!g1489)) + ((!g832) & (g2890) & (g1489)) + ((g832) & (!g2890) & (g1489)) + ((g832) & (g2890) & (g1489)));
	assign g1490 = (((!g34) & (!g36) & (!reset) & (g511) & (!g1489)) + ((!g34) & (!g36) & (!reset) & (g511) & (g1489)) + ((!g34) & (g36) & (!reset) & (!g511) & (g1489)) + ((!g34) & (g36) & (!reset) & (g511) & (g1489)) + ((g34) & (!g36) & (!reset) & (g511) & (!g1489)) + ((g34) & (!g36) & (!reset) & (g511) & (g1489)) + ((g34) & (g36) & (!reset) & (g511) & (!g1489)) + ((g34) & (g36) & (!reset) & (g511) & (g1489)));
	assign g7594 = (((!g832) & (g2892) & (!g1491)) + ((!g832) & (g2892) & (g1491)) + ((g832) & (!g2892) & (g1491)) + ((g832) & (g2892) & (g1491)));
	assign g1492 = (((!g34) & (!g36) & (!reset) & (g513) & (!g1491)) + ((!g34) & (!g36) & (!reset) & (g513) & (g1491)) + ((!g34) & (g36) & (!reset) & (!g513) & (g1491)) + ((!g34) & (g36) & (!reset) & (g513) & (g1491)) + ((g34) & (!g36) & (!reset) & (g513) & (!g1491)) + ((g34) & (!g36) & (!reset) & (g513) & (g1491)) + ((g34) & (g36) & (!reset) & (g513) & (!g1491)) + ((g34) & (g36) & (!reset) & (g513) & (g1491)));
	assign g7595 = (((!g832) & (g2894) & (!g1493)) + ((!g832) & (g2894) & (g1493)) + ((g832) & (!g2894) & (g1493)) + ((g832) & (g2894) & (g1493)));
	assign g1494 = (((!g34) & (!g36) & (!reset) & (g514) & (!g1493)) + ((!g34) & (!g36) & (!reset) & (g514) & (g1493)) + ((!g34) & (g36) & (!reset) & (!g514) & (g1493)) + ((!g34) & (g36) & (!reset) & (g514) & (g1493)) + ((g34) & (!g36) & (!reset) & (g514) & (!g1493)) + ((g34) & (!g36) & (!reset) & (g514) & (g1493)) + ((g34) & (g36) & (!reset) & (g514) & (!g1493)) + ((g34) & (g36) & (!reset) & (g514) & (g1493)));
	assign g7596 = (((!g832) & (g2896) & (!g1495)) + ((!g832) & (g2896) & (g1495)) + ((g832) & (!g2896) & (g1495)) + ((g832) & (g2896) & (g1495)));
	assign g1496 = (((!g34) & (!g36) & (!reset) & (g515) & (!g1495)) + ((!g34) & (!g36) & (!reset) & (g515) & (g1495)) + ((!g34) & (g36) & (!reset) & (!g515) & (g1495)) + ((!g34) & (g36) & (!reset) & (g515) & (g1495)) + ((g34) & (!g36) & (!reset) & (g515) & (!g1495)) + ((g34) & (!g36) & (!reset) & (g515) & (g1495)) + ((g34) & (g36) & (!reset) & (g515) & (!g1495)) + ((g34) & (g36) & (!reset) & (g515) & (g1495)));
	assign g7597 = (((!g832) & (g2898) & (!g1497)) + ((!g832) & (g2898) & (g1497)) + ((g832) & (!g2898) & (g1497)) + ((g832) & (g2898) & (g1497)));
	assign g1498 = (((!g34) & (!g36) & (!reset) & (g516) & (!g1497)) + ((!g34) & (!g36) & (!reset) & (g516) & (g1497)) + ((!g34) & (g36) & (!reset) & (!g516) & (g1497)) + ((!g34) & (g36) & (!reset) & (g516) & (g1497)) + ((g34) & (!g36) & (!reset) & (g516) & (!g1497)) + ((g34) & (!g36) & (!reset) & (g516) & (g1497)) + ((g34) & (g36) & (!reset) & (g516) & (!g1497)) + ((g34) & (g36) & (!reset) & (g516) & (g1497)));
	assign g7598 = (((!g832) & (g2899) & (!g1499)) + ((!g832) & (g2899) & (g1499)) + ((g832) & (!g2899) & (g1499)) + ((g832) & (g2899) & (g1499)));
	assign g1500 = (((!g34) & (!g36) & (!reset) & (g518) & (!g1499)) + ((!g34) & (!g36) & (!reset) & (g518) & (g1499)) + ((!g34) & (g36) & (!reset) & (!g518) & (g1499)) + ((!g34) & (g36) & (!reset) & (g518) & (g1499)) + ((g34) & (!g36) & (!reset) & (g518) & (!g1499)) + ((g34) & (!g36) & (!reset) & (g518) & (g1499)) + ((g34) & (g36) & (!reset) & (g518) & (!g1499)) + ((g34) & (g36) & (!reset) & (g518) & (g1499)));
	assign g7599 = (((!g832) & (g2901) & (!g1501)) + ((!g832) & (g2901) & (g1501)) + ((g832) & (!g2901) & (g1501)) + ((g832) & (g2901) & (g1501)));
	assign g1502 = (((!g34) & (!g36) & (!reset) & (g519) & (!g1501)) + ((!g34) & (!g36) & (!reset) & (g519) & (g1501)) + ((!g34) & (g36) & (!reset) & (!g519) & (g1501)) + ((!g34) & (g36) & (!reset) & (g519) & (g1501)) + ((g34) & (!g36) & (!reset) & (g519) & (!g1501)) + ((g34) & (!g36) & (!reset) & (g519) & (g1501)) + ((g34) & (g36) & (!reset) & (g519) & (!g1501)) + ((g34) & (g36) & (!reset) & (g519) & (g1501)));
	assign g7600 = (((!g832) & (g2903) & (!g1503)) + ((!g832) & (g2903) & (g1503)) + ((g832) & (!g2903) & (g1503)) + ((g832) & (g2903) & (g1503)));
	assign g1504 = (((!g34) & (!g36) & (!reset) & (g520) & (!g1503)) + ((!g34) & (!g36) & (!reset) & (g520) & (g1503)) + ((!g34) & (g36) & (!reset) & (!g520) & (g1503)) + ((!g34) & (g36) & (!reset) & (g520) & (g1503)) + ((g34) & (!g36) & (!reset) & (g520) & (!g1503)) + ((g34) & (!g36) & (!reset) & (g520) & (g1503)) + ((g34) & (g36) & (!reset) & (g520) & (!g1503)) + ((g34) & (g36) & (!reset) & (g520) & (g1503)));
	assign g7601 = (((!g832) & (g2905) & (!g1505)) + ((!g832) & (g2905) & (g1505)) + ((g832) & (!g2905) & (g1505)) + ((g832) & (g2905) & (g1505)));
	assign g1506 = (((!g34) & (!g36) & (!reset) & (g521) & (!g1505)) + ((!g34) & (!g36) & (!reset) & (g521) & (g1505)) + ((!g34) & (g36) & (!reset) & (!g521) & (g1505)) + ((!g34) & (g36) & (!reset) & (g521) & (g1505)) + ((g34) & (!g36) & (!reset) & (g521) & (!g1505)) + ((g34) & (!g36) & (!reset) & (g521) & (g1505)) + ((g34) & (g36) & (!reset) & (g521) & (!g1505)) + ((g34) & (g36) & (!reset) & (g521) & (g1505)));
	assign g7602 = (((!g2017) & (g2910) & (!g1507)) + ((!g2017) & (g2910) & (g1507)) + ((g2017) & (!g2910) & (g1507)) + ((g2017) & (g2910) & (g1507)));
	assign g1508 = (((!g827) & (!g501) & (!g524) & (!g1473) & (g1507) & (!g1474)) + ((!g827) & (!g501) & (!g524) & (!g1473) & (g1507) & (g1474)) + ((!g827) & (!g501) & (!g524) & (g1473) & (g1507) & (!g1474)) + ((!g827) & (!g501) & (!g524) & (g1473) & (g1507) & (g1474)) + ((!g827) & (!g501) & (g524) & (!g1473) & (g1507) & (!g1474)) + ((!g827) & (!g501) & (g524) & (!g1473) & (g1507) & (g1474)) + ((!g827) & (!g501) & (g524) & (g1473) & (g1507) & (!g1474)) + ((!g827) & (!g501) & (g524) & (g1473) & (g1507) & (g1474)) + ((!g827) & (g501) & (!g524) & (!g1473) & (g1507) & (!g1474)) + ((!g827) & (g501) & (!g524) & (!g1473) & (g1507) & (g1474)) + ((!g827) & (g501) & (!g524) & (g1473) & (g1507) & (!g1474)) + ((!g827) & (g501) & (!g524) & (g1473) & (g1507) & (g1474)) + ((!g827) & (g501) & (g524) & (!g1473) & (g1507) & (!g1474)) + ((!g827) & (g501) & (g524) & (!g1473) & (g1507) & (g1474)) + ((!g827) & (g501) & (g524) & (g1473) & (g1507) & (!g1474)) + ((!g827) & (g501) & (g524) & (g1473) & (g1507) & (g1474)) + ((g827) & (!g501) & (!g524) & (!g1473) & (g1507) & (!g1474)) + ((g827) & (!g501) & (!g524) & (!g1473) & (g1507) & (g1474)) + ((g827) & (!g501) & (!g524) & (g1473) & (!g1507) & (g1474)) + ((g827) & (!g501) & (!g524) & (g1473) & (g1507) & (!g1474)) + ((g827) & (!g501) & (g524) & (!g1473) & (!g1507) & (!g1474)) + ((g827) & (!g501) & (g524) & (!g1473) & (!g1507) & (g1474)) + ((g827) & (!g501) & (g524) & (g1473) & (!g1507) & (!g1474)) + ((g827) & (!g501) & (g524) & (g1473) & (g1507) & (g1474)) + ((g827) & (g501) & (!g524) & (!g1473) & (!g1507) & (g1474)) + ((g827) & (g501) & (!g524) & (!g1473) & (g1507) & (!g1474)) + ((g827) & (g501) & (!g524) & (g1473) & (!g1507) & (!g1474)) + ((g827) & (g501) & (!g524) & (g1473) & (!g1507) & (g1474)) + ((g827) & (g501) & (g524) & (!g1473) & (!g1507) & (!g1474)) + ((g827) & (g501) & (g524) & (!g1473) & (g1507) & (g1474)) + ((g827) & (g501) & (g524) & (g1473) & (g1507) & (!g1474)) + ((g827) & (g501) & (g524) & (g1473) & (g1507) & (g1474)));
	assign g1509 = (((!g34) & (!g36) & (!reset) & (g526) & (!g547)) + ((!g34) & (!g36) & (!reset) & (g526) & (g547)) + ((!g34) & (g36) & (!reset) & (!g526) & (g547)) + ((!g34) & (g36) & (!reset) & (g526) & (g547)) + ((g34) & (!g36) & (!reset) & (g526) & (!g547)) + ((g34) & (!g36) & (!reset) & (g526) & (g547)) + ((g34) & (g36) & (!reset) & (g526) & (!g547)) + ((g34) & (g36) & (!reset) & (g526) & (g547)));
	assign g7603 = (((!g832) & (g2915) & (!g1510)) + ((!g832) & (g2915) & (g1510)) + ((g832) & (!g2915) & (g1510)) + ((g832) & (g2915) & (g1510)));
	assign g1511 = (((!g34) & (!g36) & (!reset) & (g527) & (!g1510)) + ((!g34) & (!g36) & (!reset) & (g527) & (g1510)) + ((!g34) & (g36) & (!reset) & (!g527) & (g1510)) + ((!g34) & (g36) & (!reset) & (g527) & (g1510)) + ((g34) & (!g36) & (!reset) & (g527) & (!g1510)) + ((g34) & (!g36) & (!reset) & (g527) & (g1510)) + ((g34) & (g36) & (!reset) & (g527) & (!g1510)) + ((g34) & (g36) & (!reset) & (g527) & (g1510)));
	assign g7604 = (((!g832) & (g2921) & (!g1512)) + ((!g832) & (g2921) & (g1512)) + ((g832) & (!g2921) & (g1512)) + ((g832) & (g2921) & (g1512)));
	assign g1513 = (((!g34) & (!g36) & (!reset) & (g528) & (!g1512)) + ((!g34) & (!g36) & (!reset) & (g528) & (g1512)) + ((!g34) & (g36) & (!reset) & (!g528) & (g1512)) + ((!g34) & (g36) & (!reset) & (g528) & (g1512)) + ((g34) & (!g36) & (!reset) & (g528) & (!g1512)) + ((g34) & (!g36) & (!reset) & (g528) & (g1512)) + ((g34) & (g36) & (!reset) & (g528) & (!g1512)) + ((g34) & (g36) & (!reset) & (g528) & (g1512)));
	assign g7605 = (((!g832) & (g2926) & (!g1514)) + ((!g832) & (g2926) & (g1514)) + ((g832) & (!g2926) & (g1514)) + ((g832) & (g2926) & (g1514)));
	assign g1515 = (((!g34) & (!g36) & (!reset) & (g529) & (!g1514)) + ((!g34) & (!g36) & (!reset) & (g529) & (g1514)) + ((!g34) & (g36) & (!reset) & (!g529) & (g1514)) + ((!g34) & (g36) & (!reset) & (g529) & (g1514)) + ((g34) & (!g36) & (!reset) & (g529) & (!g1514)) + ((g34) & (!g36) & (!reset) & (g529) & (g1514)) + ((g34) & (g36) & (!reset) & (g529) & (!g1514)) + ((g34) & (g36) & (!reset) & (g529) & (g1514)));
	assign g7606 = (((!g832) & (g2931) & (!g1516)) + ((!g832) & (g2931) & (g1516)) + ((g832) & (!g2931) & (g1516)) + ((g832) & (g2931) & (g1516)));
	assign g1517 = (((!g34) & (!g36) & (!reset) & (g531) & (!g1516)) + ((!g34) & (!g36) & (!reset) & (g531) & (g1516)) + ((!g34) & (g36) & (!reset) & (!g531) & (g1516)) + ((!g34) & (g36) & (!reset) & (g531) & (g1516)) + ((g34) & (!g36) & (!reset) & (g531) & (!g1516)) + ((g34) & (!g36) & (!reset) & (g531) & (g1516)) + ((g34) & (g36) & (!reset) & (g531) & (!g1516)) + ((g34) & (g36) & (!reset) & (g531) & (g1516)));
	assign g7607 = (((!g832) & (g2937) & (!g1518)) + ((!g832) & (g2937) & (g1518)) + ((g832) & (!g2937) & (g1518)) + ((g832) & (g2937) & (g1518)));
	assign g1519 = (((!g34) & (!g36) & (!reset) & (g532) & (!g1518)) + ((!g34) & (!g36) & (!reset) & (g532) & (g1518)) + ((!g34) & (g36) & (!reset) & (!g532) & (g1518)) + ((!g34) & (g36) & (!reset) & (g532) & (g1518)) + ((g34) & (!g36) & (!reset) & (g532) & (!g1518)) + ((g34) & (!g36) & (!reset) & (g532) & (g1518)) + ((g34) & (g36) & (!reset) & (g532) & (!g1518)) + ((g34) & (g36) & (!reset) & (g532) & (g1518)));
	assign g7608 = (((!g832) & (g2943) & (!g1520)) + ((!g832) & (g2943) & (g1520)) + ((g832) & (!g2943) & (g1520)) + ((g832) & (g2943) & (g1520)));
	assign g1521 = (((!g34) & (!g36) & (!reset) & (g533) & (!g1520)) + ((!g34) & (!g36) & (!reset) & (g533) & (g1520)) + ((!g34) & (g36) & (!reset) & (!g533) & (g1520)) + ((!g34) & (g36) & (!reset) & (g533) & (g1520)) + ((g34) & (!g36) & (!reset) & (g533) & (!g1520)) + ((g34) & (!g36) & (!reset) & (g533) & (g1520)) + ((g34) & (g36) & (!reset) & (g533) & (!g1520)) + ((g34) & (g36) & (!reset) & (g533) & (g1520)));
	assign g7609 = (((!g832) & (g2949) & (!g1522)) + ((!g832) & (g2949) & (g1522)) + ((g832) & (!g2949) & (g1522)) + ((g832) & (g2949) & (g1522)));
	assign g1523 = (((!g34) & (!g36) & (!reset) & (g534) & (!g1522)) + ((!g34) & (!g36) & (!reset) & (g534) & (g1522)) + ((!g34) & (g36) & (!reset) & (!g534) & (g1522)) + ((!g34) & (g36) & (!reset) & (g534) & (g1522)) + ((g34) & (!g36) & (!reset) & (g534) & (!g1522)) + ((g34) & (!g36) & (!reset) & (g534) & (g1522)) + ((g34) & (g36) & (!reset) & (g534) & (!g1522)) + ((g34) & (g36) & (!reset) & (g534) & (g1522)));
	assign g7610 = (((!g832) & (g2955) & (!g1524)) + ((!g832) & (g2955) & (g1524)) + ((g832) & (!g2955) & (g1524)) + ((g832) & (g2955) & (g1524)));
	assign g1525 = (((!g34) & (!g36) & (!reset) & (g536) & (!g1524)) + ((!g34) & (!g36) & (!reset) & (g536) & (g1524)) + ((!g34) & (g36) & (!reset) & (!g536) & (g1524)) + ((!g34) & (g36) & (!reset) & (g536) & (g1524)) + ((g34) & (!g36) & (!reset) & (g536) & (!g1524)) + ((g34) & (!g36) & (!reset) & (g536) & (g1524)) + ((g34) & (g36) & (!reset) & (g536) & (!g1524)) + ((g34) & (g36) & (!reset) & (g536) & (g1524)));
	assign g7611 = (((!g832) & (g2961) & (!g1526)) + ((!g832) & (g2961) & (g1526)) + ((g832) & (!g2961) & (g1526)) + ((g832) & (g2961) & (g1526)));
	assign g1527 = (((!g34) & (!g36) & (!reset) & (g537) & (!g1526)) + ((!g34) & (!g36) & (!reset) & (g537) & (g1526)) + ((!g34) & (g36) & (!reset) & (!g537) & (g1526)) + ((!g34) & (g36) & (!reset) & (g537) & (g1526)) + ((g34) & (!g36) & (!reset) & (g537) & (!g1526)) + ((g34) & (!g36) & (!reset) & (g537) & (g1526)) + ((g34) & (g36) & (!reset) & (g537) & (!g1526)) + ((g34) & (g36) & (!reset) & (g537) & (g1526)));
	assign g7612 = (((!g832) & (g2967) & (!g1528)) + ((!g832) & (g2967) & (g1528)) + ((g832) & (!g2967) & (g1528)) + ((g832) & (g2967) & (g1528)));
	assign g1529 = (((!g34) & (!g36) & (!reset) & (g538) & (!g1528)) + ((!g34) & (!g36) & (!reset) & (g538) & (g1528)) + ((!g34) & (g36) & (!reset) & (!g538) & (g1528)) + ((!g34) & (g36) & (!reset) & (g538) & (g1528)) + ((g34) & (!g36) & (!reset) & (g538) & (!g1528)) + ((g34) & (!g36) & (!reset) & (g538) & (g1528)) + ((g34) & (g36) & (!reset) & (g538) & (!g1528)) + ((g34) & (g36) & (!reset) & (g538) & (g1528)));
	assign g7613 = (((!g832) & (g2973) & (!g1530)) + ((!g832) & (g2973) & (g1530)) + ((g832) & (!g2973) & (g1530)) + ((g832) & (g2973) & (g1530)));
	assign g1531 = (((!g34) & (!g36) & (!reset) & (g539) & (!g1530)) + ((!g34) & (!g36) & (!reset) & (g539) & (g1530)) + ((!g34) & (g36) & (!reset) & (!g539) & (g1530)) + ((!g34) & (g36) & (!reset) & (g539) & (g1530)) + ((g34) & (!g36) & (!reset) & (g539) & (!g1530)) + ((g34) & (!g36) & (!reset) & (g539) & (g1530)) + ((g34) & (g36) & (!reset) & (g539) & (!g1530)) + ((g34) & (g36) & (!reset) & (g539) & (g1530)));
	assign g7614 = (((!g832) & (g2978) & (!g1532)) + ((!g832) & (g2978) & (g1532)) + ((g832) & (!g2978) & (g1532)) + ((g832) & (g2978) & (g1532)));
	assign g1533 = (((!g34) & (!g36) & (!reset) & (g541) & (!g1532)) + ((!g34) & (!g36) & (!reset) & (g541) & (g1532)) + ((!g34) & (g36) & (!reset) & (!g541) & (g1532)) + ((!g34) & (g36) & (!reset) & (g541) & (g1532)) + ((g34) & (!g36) & (!reset) & (g541) & (!g1532)) + ((g34) & (!g36) & (!reset) & (g541) & (g1532)) + ((g34) & (g36) & (!reset) & (g541) & (!g1532)) + ((g34) & (g36) & (!reset) & (g541) & (g1532)));
	assign g7615 = (((!g832) & (g2984) & (!g1534)) + ((!g832) & (g2984) & (g1534)) + ((g832) & (!g2984) & (g1534)) + ((g832) & (g2984) & (g1534)));
	assign g1535 = (((!g34) & (!g36) & (!reset) & (g542) & (!g1534)) + ((!g34) & (!g36) & (!reset) & (g542) & (g1534)) + ((!g34) & (g36) & (!reset) & (!g542) & (g1534)) + ((!g34) & (g36) & (!reset) & (g542) & (g1534)) + ((g34) & (!g36) & (!reset) & (g542) & (!g1534)) + ((g34) & (!g36) & (!reset) & (g542) & (g1534)) + ((g34) & (g36) & (!reset) & (g542) & (!g1534)) + ((g34) & (g36) & (!reset) & (g542) & (g1534)));
	assign g7616 = (((!g832) & (g2990) & (!g1536)) + ((!g832) & (g2990) & (g1536)) + ((g832) & (!g2990) & (g1536)) + ((g832) & (g2990) & (g1536)));
	assign g1537 = (((!g34) & (!g36) & (!reset) & (g543) & (!g1536)) + ((!g34) & (!g36) & (!reset) & (g543) & (g1536)) + ((!g34) & (g36) & (!reset) & (!g543) & (g1536)) + ((!g34) & (g36) & (!reset) & (g543) & (g1536)) + ((g34) & (!g36) & (!reset) & (g543) & (!g1536)) + ((g34) & (!g36) & (!reset) & (g543) & (g1536)) + ((g34) & (g36) & (!reset) & (g543) & (!g1536)) + ((g34) & (g36) & (!reset) & (g543) & (g1536)));
	assign g7617 = (((!g832) & (g2996) & (!g1538)) + ((!g832) & (g2996) & (g1538)) + ((g832) & (!g2996) & (g1538)) + ((g832) & (g2996) & (g1538)));
	assign g1539 = (((!g34) & (!g36) & (!reset) & (g544) & (!g1538)) + ((!g34) & (!g36) & (!reset) & (g544) & (g1538)) + ((!g34) & (g36) & (!reset) & (!g544) & (g1538)) + ((!g34) & (g36) & (!reset) & (g544) & (g1538)) + ((g34) & (!g36) & (!reset) & (g544) & (!g1538)) + ((g34) & (!g36) & (!reset) & (g544) & (g1538)) + ((g34) & (g36) & (!reset) & (g544) & (!g1538)) + ((g34) & (g36) & (!reset) & (g544) & (g1538)));
	assign g7618 = (((!g2017) & (g7107) & (!g1540)) + ((!g2017) & (g7107) & (g1540)) + ((g2017) & (!g7107) & (g1540)) + ((g2017) & (g7107) & (g1540)));
	assign g1541 = (((!g524) & (g1507)) + ((g524) & (!g1507)));
	assign g1542 = (((!g478) & (!g501) & (g1439) & (g1473) & (!g1440) & (g1541)) + ((!g478) & (g501) & (!g1439) & (g1473) & (!g1440) & (g1541)) + ((!g478) & (g501) & (!g1439) & (g1473) & (g1440) & (g1541)) + ((!g478) & (g501) & (g1439) & (!g1473) & (!g1440) & (g1541)) + ((!g478) & (g501) & (g1439) & (g1473) & (!g1440) & (g1541)) + ((!g478) & (g501) & (g1439) & (g1473) & (g1440) & (g1541)) + ((g478) & (!g501) & (!g1439) & (g1473) & (!g1440) & (g1541)) + ((g478) & (!g501) & (g1439) & (g1473) & (!g1440) & (g1541)) + ((g478) & (!g501) & (g1439) & (g1473) & (g1440) & (g1541)) + ((g478) & (g501) & (!g1439) & (!g1473) & (!g1440) & (g1541)) + ((g478) & (g501) & (!g1439) & (g1473) & (!g1440) & (g1541)) + ((g478) & (g501) & (!g1439) & (g1473) & (g1440) & (g1541)) + ((g478) & (g501) & (g1439) & (!g1473) & (!g1440) & (g1541)) + ((g478) & (g501) & (g1439) & (!g1473) & (g1440) & (g1541)) + ((g478) & (g501) & (g1439) & (g1473) & (!g1440) & (g1541)) + ((g478) & (g501) & (g1439) & (g1473) & (g1440) & (g1541)));
	assign g1543 = (((g524) & (g1507)));
	assign g1544 = (((!g1542) & (!g1543)));
	assign g1545 = (((!g827) & (!g547) & (g1540) & (!g1544)) + ((!g827) & (!g547) & (g1540) & (g1544)) + ((!g827) & (g547) & (g1540) & (!g1544)) + ((!g827) & (g547) & (g1540) & (g1544)) + ((g827) & (!g547) & (!g1540) & (!g1544)) + ((g827) & (!g547) & (g1540) & (g1544)) + ((g827) & (g547) & (!g1540) & (g1544)) + ((g827) & (g547) & (g1540) & (!g1544)));
	assign g1546 = (((!g34) & (!g36) & (!reset) & (g549) & (!g570)) + ((!g34) & (!g36) & (!reset) & (g549) & (g570)) + ((!g34) & (g36) & (!reset) & (!g549) & (g570)) + ((!g34) & (g36) & (!reset) & (g549) & (g570)) + ((g34) & (!g36) & (!reset) & (g549) & (!g570)) + ((g34) & (!g36) & (!reset) & (g549) & (g570)) + ((g34) & (g36) & (!reset) & (g549) & (!g570)) + ((g34) & (g36) & (!reset) & (g549) & (g570)));
	assign g7619 = (((!g832) & (g2998) & (!g1547)) + ((!g832) & (g2998) & (g1547)) + ((g832) & (!g2998) & (g1547)) + ((g832) & (g2998) & (g1547)));
	assign g1548 = (((!g34) & (!g36) & (!reset) & (g550) & (!g1547)) + ((!g34) & (!g36) & (!reset) & (g550) & (g1547)) + ((!g34) & (g36) & (!reset) & (!g550) & (g1547)) + ((!g34) & (g36) & (!reset) & (g550) & (g1547)) + ((g34) & (!g36) & (!reset) & (g550) & (!g1547)) + ((g34) & (!g36) & (!reset) & (g550) & (g1547)) + ((g34) & (g36) & (!reset) & (g550) & (!g1547)) + ((g34) & (g36) & (!reset) & (g550) & (g1547)));
	assign g7620 = (((!g832) & (g3000) & (!g1549)) + ((!g832) & (g3000) & (g1549)) + ((g832) & (!g3000) & (g1549)) + ((g832) & (g3000) & (g1549)));
	assign g1550 = (((!g34) & (!g36) & (!reset) & (g551) & (!g1549)) + ((!g34) & (!g36) & (!reset) & (g551) & (g1549)) + ((!g34) & (g36) & (!reset) & (!g551) & (g1549)) + ((!g34) & (g36) & (!reset) & (g551) & (g1549)) + ((g34) & (!g36) & (!reset) & (g551) & (!g1549)) + ((g34) & (!g36) & (!reset) & (g551) & (g1549)) + ((g34) & (g36) & (!reset) & (g551) & (!g1549)) + ((g34) & (g36) & (!reset) & (g551) & (g1549)));
	assign g7621 = (((!g832) & (g3001) & (!g1551)) + ((!g832) & (g3001) & (g1551)) + ((g832) & (!g3001) & (g1551)) + ((g832) & (g3001) & (g1551)));
	assign g1552 = (((!g34) & (!g36) & (!reset) & (g552) & (!g1551)) + ((!g34) & (!g36) & (!reset) & (g552) & (g1551)) + ((!g34) & (g36) & (!reset) & (!g552) & (g1551)) + ((!g34) & (g36) & (!reset) & (g552) & (g1551)) + ((g34) & (!g36) & (!reset) & (g552) & (!g1551)) + ((g34) & (!g36) & (!reset) & (g552) & (g1551)) + ((g34) & (g36) & (!reset) & (g552) & (!g1551)) + ((g34) & (g36) & (!reset) & (g552) & (g1551)));
	assign g7622 = (((!g832) & (g3002) & (!g1553)) + ((!g832) & (g3002) & (g1553)) + ((g832) & (!g3002) & (g1553)) + ((g832) & (g3002) & (g1553)));
	assign g1554 = (((!g34) & (!g36) & (!reset) & (g554) & (!g1553)) + ((!g34) & (!g36) & (!reset) & (g554) & (g1553)) + ((!g34) & (g36) & (!reset) & (!g554) & (g1553)) + ((!g34) & (g36) & (!reset) & (g554) & (g1553)) + ((g34) & (!g36) & (!reset) & (g554) & (!g1553)) + ((g34) & (!g36) & (!reset) & (g554) & (g1553)) + ((g34) & (g36) & (!reset) & (g554) & (!g1553)) + ((g34) & (g36) & (!reset) & (g554) & (g1553)));
	assign g7623 = (((!g832) & (g3004) & (!g1555)) + ((!g832) & (g3004) & (g1555)) + ((g832) & (!g3004) & (g1555)) + ((g832) & (g3004) & (g1555)));
	assign g1556 = (((!g34) & (!g36) & (!reset) & (g555) & (!g1555)) + ((!g34) & (!g36) & (!reset) & (g555) & (g1555)) + ((!g34) & (g36) & (!reset) & (!g555) & (g1555)) + ((!g34) & (g36) & (!reset) & (g555) & (g1555)) + ((g34) & (!g36) & (!reset) & (g555) & (!g1555)) + ((g34) & (!g36) & (!reset) & (g555) & (g1555)) + ((g34) & (g36) & (!reset) & (g555) & (!g1555)) + ((g34) & (g36) & (!reset) & (g555) & (g1555)));
	assign g7624 = (((!g832) & (g3006) & (!g1557)) + ((!g832) & (g3006) & (g1557)) + ((g832) & (!g3006) & (g1557)) + ((g832) & (g3006) & (g1557)));
	assign g1558 = (((!g34) & (!g36) & (!reset) & (g556) & (!g1557)) + ((!g34) & (!g36) & (!reset) & (g556) & (g1557)) + ((!g34) & (g36) & (!reset) & (!g556) & (g1557)) + ((!g34) & (g36) & (!reset) & (g556) & (g1557)) + ((g34) & (!g36) & (!reset) & (g556) & (!g1557)) + ((g34) & (!g36) & (!reset) & (g556) & (g1557)) + ((g34) & (g36) & (!reset) & (g556) & (!g1557)) + ((g34) & (g36) & (!reset) & (g556) & (g1557)));
	assign g7625 = (((!g832) & (g3008) & (!g1559)) + ((!g832) & (g3008) & (g1559)) + ((g832) & (!g3008) & (g1559)) + ((g832) & (g3008) & (g1559)));
	assign g1560 = (((!g34) & (!g36) & (!reset) & (g557) & (!g1559)) + ((!g34) & (!g36) & (!reset) & (g557) & (g1559)) + ((!g34) & (g36) & (!reset) & (!g557) & (g1559)) + ((!g34) & (g36) & (!reset) & (g557) & (g1559)) + ((g34) & (!g36) & (!reset) & (g557) & (!g1559)) + ((g34) & (!g36) & (!reset) & (g557) & (g1559)) + ((g34) & (g36) & (!reset) & (g557) & (!g1559)) + ((g34) & (g36) & (!reset) & (g557) & (g1559)));
	assign g7626 = (((!g832) & (g3010) & (!g1561)) + ((!g832) & (g3010) & (g1561)) + ((g832) & (!g3010) & (g1561)) + ((g832) & (g3010) & (g1561)));
	assign g1562 = (((!g34) & (!g36) & (!reset) & (g559) & (!g1561)) + ((!g34) & (!g36) & (!reset) & (g559) & (g1561)) + ((!g34) & (g36) & (!reset) & (!g559) & (g1561)) + ((!g34) & (g36) & (!reset) & (g559) & (g1561)) + ((g34) & (!g36) & (!reset) & (g559) & (!g1561)) + ((g34) & (!g36) & (!reset) & (g559) & (g1561)) + ((g34) & (g36) & (!reset) & (g559) & (!g1561)) + ((g34) & (g36) & (!reset) & (g559) & (g1561)));
	assign g7627 = (((!g832) & (g3012) & (!g1563)) + ((!g832) & (g3012) & (g1563)) + ((g832) & (!g3012) & (g1563)) + ((g832) & (g3012) & (g1563)));
	assign g1564 = (((!g34) & (!g36) & (!reset) & (g560) & (!g1563)) + ((!g34) & (!g36) & (!reset) & (g560) & (g1563)) + ((!g34) & (g36) & (!reset) & (!g560) & (g1563)) + ((!g34) & (g36) & (!reset) & (g560) & (g1563)) + ((g34) & (!g36) & (!reset) & (g560) & (!g1563)) + ((g34) & (!g36) & (!reset) & (g560) & (g1563)) + ((g34) & (g36) & (!reset) & (g560) & (!g1563)) + ((g34) & (g36) & (!reset) & (g560) & (g1563)));
	assign g7628 = (((!g832) & (g3014) & (!g1565)) + ((!g832) & (g3014) & (g1565)) + ((g832) & (!g3014) & (g1565)) + ((g832) & (g3014) & (g1565)));
	assign g1566 = (((!g34) & (!g36) & (!reset) & (g561) & (!g1565)) + ((!g34) & (!g36) & (!reset) & (g561) & (g1565)) + ((!g34) & (g36) & (!reset) & (!g561) & (g1565)) + ((!g34) & (g36) & (!reset) & (g561) & (g1565)) + ((g34) & (!g36) & (!reset) & (g561) & (!g1565)) + ((g34) & (!g36) & (!reset) & (g561) & (g1565)) + ((g34) & (g36) & (!reset) & (g561) & (!g1565)) + ((g34) & (g36) & (!reset) & (g561) & (g1565)));
	assign g7629 = (((!g832) & (g3016) & (!g1567)) + ((!g832) & (g3016) & (g1567)) + ((g832) & (!g3016) & (g1567)) + ((g832) & (g3016) & (g1567)));
	assign g1568 = (((!g34) & (!g36) & (!reset) & (g562) & (!g1567)) + ((!g34) & (!g36) & (!reset) & (g562) & (g1567)) + ((!g34) & (g36) & (!reset) & (!g562) & (g1567)) + ((!g34) & (g36) & (!reset) & (g562) & (g1567)) + ((g34) & (!g36) & (!reset) & (g562) & (!g1567)) + ((g34) & (!g36) & (!reset) & (g562) & (g1567)) + ((g34) & (g36) & (!reset) & (g562) & (!g1567)) + ((g34) & (g36) & (!reset) & (g562) & (g1567)));
	assign g7630 = (((!g832) & (g3017) & (!g1569)) + ((!g832) & (g3017) & (g1569)) + ((g832) & (!g3017) & (g1569)) + ((g832) & (g3017) & (g1569)));
	assign g1570 = (((!g34) & (!g36) & (!reset) & (g564) & (!g1569)) + ((!g34) & (!g36) & (!reset) & (g564) & (g1569)) + ((!g34) & (g36) & (!reset) & (!g564) & (g1569)) + ((!g34) & (g36) & (!reset) & (g564) & (g1569)) + ((g34) & (!g36) & (!reset) & (g564) & (!g1569)) + ((g34) & (!g36) & (!reset) & (g564) & (g1569)) + ((g34) & (g36) & (!reset) & (g564) & (!g1569)) + ((g34) & (g36) & (!reset) & (g564) & (g1569)));
	assign g7631 = (((!g832) & (g3019) & (!g1571)) + ((!g832) & (g3019) & (g1571)) + ((g832) & (!g3019) & (g1571)) + ((g832) & (g3019) & (g1571)));
	assign g1572 = (((!g34) & (!g36) & (!reset) & (g565) & (!g1571)) + ((!g34) & (!g36) & (!reset) & (g565) & (g1571)) + ((!g34) & (g36) & (!reset) & (!g565) & (g1571)) + ((!g34) & (g36) & (!reset) & (g565) & (g1571)) + ((g34) & (!g36) & (!reset) & (g565) & (!g1571)) + ((g34) & (!g36) & (!reset) & (g565) & (g1571)) + ((g34) & (g36) & (!reset) & (g565) & (!g1571)) + ((g34) & (g36) & (!reset) & (g565) & (g1571)));
	assign g7632 = (((!g832) & (g3021) & (!g1573)) + ((!g832) & (g3021) & (g1573)) + ((g832) & (!g3021) & (g1573)) + ((g832) & (g3021) & (g1573)));
	assign g1574 = (((!g34) & (!g36) & (!reset) & (g566) & (!g1573)) + ((!g34) & (!g36) & (!reset) & (g566) & (g1573)) + ((!g34) & (g36) & (!reset) & (!g566) & (g1573)) + ((!g34) & (g36) & (!reset) & (g566) & (g1573)) + ((g34) & (!g36) & (!reset) & (g566) & (!g1573)) + ((g34) & (!g36) & (!reset) & (g566) & (g1573)) + ((g34) & (g36) & (!reset) & (g566) & (!g1573)) + ((g34) & (g36) & (!reset) & (g566) & (g1573)));
	assign g7633 = (((!g832) & (g3023) & (!g1575)) + ((!g832) & (g3023) & (g1575)) + ((g832) & (!g3023) & (g1575)) + ((g832) & (g3023) & (g1575)));
	assign g1576 = (((!g34) & (!g36) & (!reset) & (g567) & (!g1575)) + ((!g34) & (!g36) & (!reset) & (g567) & (g1575)) + ((!g34) & (g36) & (!reset) & (!g567) & (g1575)) + ((!g34) & (g36) & (!reset) & (g567) & (g1575)) + ((g34) & (!g36) & (!reset) & (g567) & (!g1575)) + ((g34) & (!g36) & (!reset) & (g567) & (g1575)) + ((g34) & (g36) & (!reset) & (g567) & (!g1575)) + ((g34) & (g36) & (!reset) & (g567) & (g1575)));
	assign g7634 = (((!g2017) & (g3028) & (!g1577)) + ((!g2017) & (g3028) & (g1577)) + ((g2017) & (!g3028) & (g1577)) + ((g2017) & (g3028) & (g1577)));
	assign g1578 = (((!g827) & (!g547) & (!g570) & (!g1540) & (g1577) & (!g1544)) + ((!g827) & (!g547) & (!g570) & (!g1540) & (g1577) & (g1544)) + ((!g827) & (!g547) & (!g570) & (g1540) & (g1577) & (!g1544)) + ((!g827) & (!g547) & (!g570) & (g1540) & (g1577) & (g1544)) + ((!g827) & (!g547) & (g570) & (!g1540) & (g1577) & (!g1544)) + ((!g827) & (!g547) & (g570) & (!g1540) & (g1577) & (g1544)) + ((!g827) & (!g547) & (g570) & (g1540) & (g1577) & (!g1544)) + ((!g827) & (!g547) & (g570) & (g1540) & (g1577) & (g1544)) + ((!g827) & (g547) & (!g570) & (!g1540) & (g1577) & (!g1544)) + ((!g827) & (g547) & (!g570) & (!g1540) & (g1577) & (g1544)) + ((!g827) & (g547) & (!g570) & (g1540) & (g1577) & (!g1544)) + ((!g827) & (g547) & (!g570) & (g1540) & (g1577) & (g1544)) + ((!g827) & (g547) & (g570) & (!g1540) & (g1577) & (!g1544)) + ((!g827) & (g547) & (g570) & (!g1540) & (g1577) & (g1544)) + ((!g827) & (g547) & (g570) & (g1540) & (g1577) & (!g1544)) + ((!g827) & (g547) & (g570) & (g1540) & (g1577) & (g1544)) + ((g827) & (!g547) & (!g570) & (!g1540) & (g1577) & (!g1544)) + ((g827) & (!g547) & (!g570) & (!g1540) & (g1577) & (g1544)) + ((g827) & (!g547) & (!g570) & (g1540) & (!g1577) & (!g1544)) + ((g827) & (!g547) & (!g570) & (g1540) & (g1577) & (g1544)) + ((g827) & (!g547) & (g570) & (!g1540) & (!g1577) & (!g1544)) + ((g827) & (!g547) & (g570) & (!g1540) & (!g1577) & (g1544)) + ((g827) & (!g547) & (g570) & (g1540) & (!g1577) & (g1544)) + ((g827) & (!g547) & (g570) & (g1540) & (g1577) & (!g1544)) + ((g827) & (g547) & (!g570) & (!g1540) & (!g1577) & (!g1544)) + ((g827) & (g547) & (!g570) & (!g1540) & (g1577) & (g1544)) + ((g827) & (g547) & (!g570) & (g1540) & (!g1577) & (!g1544)) + ((g827) & (g547) & (!g570) & (g1540) & (!g1577) & (g1544)) + ((g827) & (g547) & (g570) & (!g1540) & (!g1577) & (g1544)) + ((g827) & (g547) & (g570) & (!g1540) & (g1577) & (!g1544)) + ((g827) & (g547) & (g570) & (g1540) & (g1577) & (!g1544)) + ((g827) & (g547) & (g570) & (g1540) & (g1577) & (g1544)));
	assign g1579 = (((!g34) & (!g36) & (!reset) & (g572) & (!g593)) + ((!g34) & (!g36) & (!reset) & (g572) & (g593)) + ((!g34) & (g36) & (!reset) & (!g572) & (g593)) + ((!g34) & (g36) & (!reset) & (g572) & (g593)) + ((g34) & (!g36) & (!reset) & (g572) & (!g593)) + ((g34) & (!g36) & (!reset) & (g572) & (g593)) + ((g34) & (g36) & (!reset) & (g572) & (!g593)) + ((g34) & (g36) & (!reset) & (g572) & (g593)));
	assign g7635 = (((!g832) & (g3030) & (!g1580)) + ((!g832) & (g3030) & (g1580)) + ((g832) & (!g3030) & (g1580)) + ((g832) & (g3030) & (g1580)));
	assign g1581 = (((!g34) & (!g36) & (!reset) & (g573) & (!g1580)) + ((!g34) & (!g36) & (!reset) & (g573) & (g1580)) + ((!g34) & (g36) & (!reset) & (!g573) & (g1580)) + ((!g34) & (g36) & (!reset) & (g573) & (g1580)) + ((g34) & (!g36) & (!reset) & (g573) & (!g1580)) + ((g34) & (!g36) & (!reset) & (g573) & (g1580)) + ((g34) & (g36) & (!reset) & (g573) & (!g1580)) + ((g34) & (g36) & (!reset) & (g573) & (g1580)));
	assign g7636 = (((!g832) & (g3033) & (!g1582)) + ((!g832) & (g3033) & (g1582)) + ((g832) & (!g3033) & (g1582)) + ((g832) & (g3033) & (g1582)));
	assign g1583 = (((!g34) & (!g36) & (!reset) & (g574) & (!g1582)) + ((!g34) & (!g36) & (!reset) & (g574) & (g1582)) + ((!g34) & (g36) & (!reset) & (!g574) & (g1582)) + ((!g34) & (g36) & (!reset) & (g574) & (g1582)) + ((g34) & (!g36) & (!reset) & (g574) & (!g1582)) + ((g34) & (!g36) & (!reset) & (g574) & (g1582)) + ((g34) & (g36) & (!reset) & (g574) & (!g1582)) + ((g34) & (g36) & (!reset) & (g574) & (g1582)));
	assign g7637 = (((!g832) & (g3035) & (!g1584)) + ((!g832) & (g3035) & (g1584)) + ((g832) & (!g3035) & (g1584)) + ((g832) & (g3035) & (g1584)));
	assign g1585 = (((!g34) & (!g36) & (!reset) & (g575) & (!g1584)) + ((!g34) & (!g36) & (!reset) & (g575) & (g1584)) + ((!g34) & (g36) & (!reset) & (!g575) & (g1584)) + ((!g34) & (g36) & (!reset) & (g575) & (g1584)) + ((g34) & (!g36) & (!reset) & (g575) & (!g1584)) + ((g34) & (!g36) & (!reset) & (g575) & (g1584)) + ((g34) & (g36) & (!reset) & (g575) & (!g1584)) + ((g34) & (g36) & (!reset) & (g575) & (g1584)));
	assign g7638 = (((!g832) & (g3037) & (!g1586)) + ((!g832) & (g3037) & (g1586)) + ((g832) & (!g3037) & (g1586)) + ((g832) & (g3037) & (g1586)));
	assign g1587 = (((!g34) & (!g36) & (!reset) & (g577) & (!g1586)) + ((!g34) & (!g36) & (!reset) & (g577) & (g1586)) + ((!g34) & (g36) & (!reset) & (!g577) & (g1586)) + ((!g34) & (g36) & (!reset) & (g577) & (g1586)) + ((g34) & (!g36) & (!reset) & (g577) & (!g1586)) + ((g34) & (!g36) & (!reset) & (g577) & (g1586)) + ((g34) & (g36) & (!reset) & (g577) & (!g1586)) + ((g34) & (g36) & (!reset) & (g577) & (g1586)));
	assign g7639 = (((!g832) & (g3040) & (!g1588)) + ((!g832) & (g3040) & (g1588)) + ((g832) & (!g3040) & (g1588)) + ((g832) & (g3040) & (g1588)));
	assign g1589 = (((!g34) & (!g36) & (!reset) & (g578) & (!g1588)) + ((!g34) & (!g36) & (!reset) & (g578) & (g1588)) + ((!g34) & (g36) & (!reset) & (!g578) & (g1588)) + ((!g34) & (g36) & (!reset) & (g578) & (g1588)) + ((g34) & (!g36) & (!reset) & (g578) & (!g1588)) + ((g34) & (!g36) & (!reset) & (g578) & (g1588)) + ((g34) & (g36) & (!reset) & (g578) & (!g1588)) + ((g34) & (g36) & (!reset) & (g578) & (g1588)));
	assign g7640 = (((!g832) & (g3043) & (!g1590)) + ((!g832) & (g3043) & (g1590)) + ((g832) & (!g3043) & (g1590)) + ((g832) & (g3043) & (g1590)));
	assign g1591 = (((!g34) & (!g36) & (!reset) & (g579) & (!g1590)) + ((!g34) & (!g36) & (!reset) & (g579) & (g1590)) + ((!g34) & (g36) & (!reset) & (!g579) & (g1590)) + ((!g34) & (g36) & (!reset) & (g579) & (g1590)) + ((g34) & (!g36) & (!reset) & (g579) & (!g1590)) + ((g34) & (!g36) & (!reset) & (g579) & (g1590)) + ((g34) & (g36) & (!reset) & (g579) & (!g1590)) + ((g34) & (g36) & (!reset) & (g579) & (g1590)));
	assign g7641 = (((!g832) & (g3046) & (!g1592)) + ((!g832) & (g3046) & (g1592)) + ((g832) & (!g3046) & (g1592)) + ((g832) & (g3046) & (g1592)));
	assign g1593 = (((!g34) & (!g36) & (!reset) & (g580) & (!g1592)) + ((!g34) & (!g36) & (!reset) & (g580) & (g1592)) + ((!g34) & (g36) & (!reset) & (!g580) & (g1592)) + ((!g34) & (g36) & (!reset) & (g580) & (g1592)) + ((g34) & (!g36) & (!reset) & (g580) & (!g1592)) + ((g34) & (!g36) & (!reset) & (g580) & (g1592)) + ((g34) & (g36) & (!reset) & (g580) & (!g1592)) + ((g34) & (g36) & (!reset) & (g580) & (g1592)));
	assign g7642 = (((!g832) & (g3049) & (!g1594)) + ((!g832) & (g3049) & (g1594)) + ((g832) & (!g3049) & (g1594)) + ((g832) & (g3049) & (g1594)));
	assign g1595 = (((!g34) & (!g36) & (!reset) & (g582) & (!g1594)) + ((!g34) & (!g36) & (!reset) & (g582) & (g1594)) + ((!g34) & (g36) & (!reset) & (!g582) & (g1594)) + ((!g34) & (g36) & (!reset) & (g582) & (g1594)) + ((g34) & (!g36) & (!reset) & (g582) & (!g1594)) + ((g34) & (!g36) & (!reset) & (g582) & (g1594)) + ((g34) & (g36) & (!reset) & (g582) & (!g1594)) + ((g34) & (g36) & (!reset) & (g582) & (g1594)));
	assign g7643 = (((!g832) & (g3052) & (!g1596)) + ((!g832) & (g3052) & (g1596)) + ((g832) & (!g3052) & (g1596)) + ((g832) & (g3052) & (g1596)));
	assign g1597 = (((!g34) & (!g36) & (!reset) & (g583) & (!g1596)) + ((!g34) & (!g36) & (!reset) & (g583) & (g1596)) + ((!g34) & (g36) & (!reset) & (!g583) & (g1596)) + ((!g34) & (g36) & (!reset) & (g583) & (g1596)) + ((g34) & (!g36) & (!reset) & (g583) & (!g1596)) + ((g34) & (!g36) & (!reset) & (g583) & (g1596)) + ((g34) & (g36) & (!reset) & (g583) & (!g1596)) + ((g34) & (g36) & (!reset) & (g583) & (g1596)));
	assign g7644 = (((!g832) & (g3055) & (!g1598)) + ((!g832) & (g3055) & (g1598)) + ((g832) & (!g3055) & (g1598)) + ((g832) & (g3055) & (g1598)));
	assign g1599 = (((!g34) & (!g36) & (!reset) & (g584) & (!g1598)) + ((!g34) & (!g36) & (!reset) & (g584) & (g1598)) + ((!g34) & (g36) & (!reset) & (!g584) & (g1598)) + ((!g34) & (g36) & (!reset) & (g584) & (g1598)) + ((g34) & (!g36) & (!reset) & (g584) & (!g1598)) + ((g34) & (!g36) & (!reset) & (g584) & (g1598)) + ((g34) & (g36) & (!reset) & (g584) & (!g1598)) + ((g34) & (g36) & (!reset) & (g584) & (g1598)));
	assign g7645 = (((!g832) & (g3058) & (!g1600)) + ((!g832) & (g3058) & (g1600)) + ((g832) & (!g3058) & (g1600)) + ((g832) & (g3058) & (g1600)));
	assign g1601 = (((!g34) & (!g36) & (!reset) & (g585) & (!g1600)) + ((!g34) & (!g36) & (!reset) & (g585) & (g1600)) + ((!g34) & (g36) & (!reset) & (!g585) & (g1600)) + ((!g34) & (g36) & (!reset) & (g585) & (g1600)) + ((g34) & (!g36) & (!reset) & (g585) & (!g1600)) + ((g34) & (!g36) & (!reset) & (g585) & (g1600)) + ((g34) & (g36) & (!reset) & (g585) & (!g1600)) + ((g34) & (g36) & (!reset) & (g585) & (g1600)));
	assign g7646 = (((!g832) & (g3060) & (!g1602)) + ((!g832) & (g3060) & (g1602)) + ((g832) & (!g3060) & (g1602)) + ((g832) & (g3060) & (g1602)));
	assign g1603 = (((!g34) & (!g36) & (!reset) & (g587) & (!g1602)) + ((!g34) & (!g36) & (!reset) & (g587) & (g1602)) + ((!g34) & (g36) & (!reset) & (!g587) & (g1602)) + ((!g34) & (g36) & (!reset) & (g587) & (g1602)) + ((g34) & (!g36) & (!reset) & (g587) & (!g1602)) + ((g34) & (!g36) & (!reset) & (g587) & (g1602)) + ((g34) & (g36) & (!reset) & (g587) & (!g1602)) + ((g34) & (g36) & (!reset) & (g587) & (g1602)));
	assign g7647 = (((!g832) & (g3063) & (!g1604)) + ((!g832) & (g3063) & (g1604)) + ((g832) & (!g3063) & (g1604)) + ((g832) & (g3063) & (g1604)));
	assign g1605 = (((!g34) & (!g36) & (!reset) & (g588) & (!g1604)) + ((!g34) & (!g36) & (!reset) & (g588) & (g1604)) + ((!g34) & (g36) & (!reset) & (!g588) & (g1604)) + ((!g34) & (g36) & (!reset) & (g588) & (g1604)) + ((g34) & (!g36) & (!reset) & (g588) & (!g1604)) + ((g34) & (!g36) & (!reset) & (g588) & (g1604)) + ((g34) & (g36) & (!reset) & (g588) & (!g1604)) + ((g34) & (g36) & (!reset) & (g588) & (g1604)));
	assign g7648 = (((!g832) & (g3066) & (!g1606)) + ((!g832) & (g3066) & (g1606)) + ((g832) & (!g3066) & (g1606)) + ((g832) & (g3066) & (g1606)));
	assign g1607 = (((!g34) & (!g36) & (!reset) & (g589) & (!g1606)) + ((!g34) & (!g36) & (!reset) & (g589) & (g1606)) + ((!g34) & (g36) & (!reset) & (!g589) & (g1606)) + ((!g34) & (g36) & (!reset) & (g589) & (g1606)) + ((g34) & (!g36) & (!reset) & (g589) & (!g1606)) + ((g34) & (!g36) & (!reset) & (g589) & (g1606)) + ((g34) & (g36) & (!reset) & (g589) & (!g1606)) + ((g34) & (g36) & (!reset) & (g589) & (g1606)));
	assign g7649 = (((!g832) & (g3069) & (!g1608)) + ((!g832) & (g3069) & (g1608)) + ((g832) & (!g3069) & (g1608)) + ((g832) & (g3069) & (g1608)));
	assign g1609 = (((!g34) & (!g36) & (!reset) & (g590) & (!g1608)) + ((!g34) & (!g36) & (!reset) & (g590) & (g1608)) + ((!g34) & (g36) & (!reset) & (!g590) & (g1608)) + ((!g34) & (g36) & (!reset) & (g590) & (g1608)) + ((g34) & (!g36) & (!reset) & (g590) & (!g1608)) + ((g34) & (!g36) & (!reset) & (g590) & (g1608)) + ((g34) & (g36) & (!reset) & (g590) & (!g1608)) + ((g34) & (g36) & (!reset) & (g590) & (g1608)));
	assign g7650 = (((!g2017) & (g3072) & (!g1610)) + ((!g2017) & (g3072) & (g1610)) + ((g2017) & (!g3072) & (g1610)) + ((g2017) & (g3072) & (g1610)));
	assign g1611 = (((!g547) & (!g570) & (!g1540) & (!g1577) & (!g1542) & (!g1543)) + ((!g547) & (!g570) & (!g1540) & (!g1577) & (!g1542) & (g1543)) + ((!g547) & (!g570) & (!g1540) & (!g1577) & (g1542) & (!g1543)) + ((!g547) & (!g570) & (!g1540) & (!g1577) & (g1542) & (g1543)) + ((!g547) & (!g570) & (!g1540) & (g1577) & (!g1542) & (!g1543)) + ((!g547) & (!g570) & (!g1540) & (g1577) & (!g1542) & (g1543)) + ((!g547) & (!g570) & (!g1540) & (g1577) & (g1542) & (!g1543)) + ((!g547) & (!g570) & (!g1540) & (g1577) & (g1542) & (g1543)) + ((!g547) & (!g570) & (g1540) & (!g1577) & (!g1542) & (!g1543)) + ((!g547) & (!g570) & (g1540) & (!g1577) & (!g1542) & (g1543)) + ((!g547) & (!g570) & (g1540) & (!g1577) & (g1542) & (!g1543)) + ((!g547) & (!g570) & (g1540) & (!g1577) & (g1542) & (g1543)) + ((!g547) & (!g570) & (g1540) & (g1577) & (!g1542) & (!g1543)) + ((!g547) & (g570) & (!g1540) & (!g1577) & (!g1542) & (!g1543)) + ((!g547) & (g570) & (!g1540) & (!g1577) & (!g1542) & (g1543)) + ((!g547) & (g570) & (!g1540) & (!g1577) & (g1542) & (!g1543)) + ((!g547) & (g570) & (!g1540) & (!g1577) & (g1542) & (g1543)) + ((!g547) & (g570) & (g1540) & (!g1577) & (!g1542) & (!g1543)) + ((g547) & (!g570) & (!g1540) & (!g1577) & (!g1542) & (!g1543)) + ((g547) & (!g570) & (!g1540) & (!g1577) & (!g1542) & (g1543)) + ((g547) & (!g570) & (!g1540) & (!g1577) & (g1542) & (!g1543)) + ((g547) & (!g570) & (!g1540) & (!g1577) & (g1542) & (g1543)) + ((g547) & (!g570) & (!g1540) & (g1577) & (!g1542) & (!g1543)) + ((g547) & (!g570) & (g1540) & (!g1577) & (!g1542) & (!g1543)) + ((g547) & (!g570) & (g1540) & (!g1577) & (!g1542) & (g1543)) + ((g547) & (!g570) & (g1540) & (!g1577) & (g1542) & (!g1543)) + ((g547) & (!g570) & (g1540) & (!g1577) & (g1542) & (g1543)) + ((g547) & (g570) & (!g1540) & (!g1577) & (!g1542) & (!g1543)));
	assign g1612 = (((!g827) & (!g593) & (g1610) & (!g1611)) + ((!g827) & (!g593) & (g1610) & (g1611)) + ((!g827) & (g593) & (g1610) & (!g1611)) + ((!g827) & (g593) & (g1610) & (g1611)) + ((g827) & (!g593) & (!g1610) & (!g1611)) + ((g827) & (!g593) & (g1610) & (g1611)) + ((g827) & (g593) & (!g1610) & (g1611)) + ((g827) & (g593) & (g1610) & (!g1611)));
	assign g1613 = (((!g34) & (!g36) & (!reset) & (g595) & (!g616)) + ((!g34) & (!g36) & (!reset) & (g595) & (g616)) + ((!g34) & (g36) & (!reset) & (!g595) & (g616)) + ((!g34) & (g36) & (!reset) & (g595) & (g616)) + ((g34) & (!g36) & (!reset) & (g595) & (!g616)) + ((g34) & (!g36) & (!reset) & (g595) & (g616)) + ((g34) & (g36) & (!reset) & (g595) & (!g616)) + ((g34) & (g36) & (!reset) & (g595) & (g616)));
	assign g7651 = (((!g832) & (g3073) & (!g1614)) + ((!g832) & (g3073) & (g1614)) + ((g832) & (!g3073) & (g1614)) + ((g832) & (g3073) & (g1614)));
	assign g1615 = (((!g34) & (!g36) & (!reset) & (g596) & (!g1614)) + ((!g34) & (!g36) & (!reset) & (g596) & (g1614)) + ((!g34) & (g36) & (!reset) & (!g596) & (g1614)) + ((!g34) & (g36) & (!reset) & (g596) & (g1614)) + ((g34) & (!g36) & (!reset) & (g596) & (!g1614)) + ((g34) & (!g36) & (!reset) & (g596) & (g1614)) + ((g34) & (g36) & (!reset) & (g596) & (!g1614)) + ((g34) & (g36) & (!reset) & (g596) & (g1614)));
	assign g7652 = (((!g832) & (g3075) & (!g1616)) + ((!g832) & (g3075) & (g1616)) + ((g832) & (!g3075) & (g1616)) + ((g832) & (g3075) & (g1616)));
	assign g1617 = (((!g34) & (!g36) & (!reset) & (g597) & (!g1616)) + ((!g34) & (!g36) & (!reset) & (g597) & (g1616)) + ((!g34) & (g36) & (!reset) & (!g597) & (g1616)) + ((!g34) & (g36) & (!reset) & (g597) & (g1616)) + ((g34) & (!g36) & (!reset) & (g597) & (!g1616)) + ((g34) & (!g36) & (!reset) & (g597) & (g1616)) + ((g34) & (g36) & (!reset) & (g597) & (!g1616)) + ((g34) & (g36) & (!reset) & (g597) & (g1616)));
	assign g7653 = (((!g832) & (g3076) & (!g1618)) + ((!g832) & (g3076) & (g1618)) + ((g832) & (!g3076) & (g1618)) + ((g832) & (g3076) & (g1618)));
	assign g1619 = (((!g34) & (!g36) & (!reset) & (g598) & (!g1618)) + ((!g34) & (!g36) & (!reset) & (g598) & (g1618)) + ((!g34) & (g36) & (!reset) & (!g598) & (g1618)) + ((!g34) & (g36) & (!reset) & (g598) & (g1618)) + ((g34) & (!g36) & (!reset) & (g598) & (!g1618)) + ((g34) & (!g36) & (!reset) & (g598) & (g1618)) + ((g34) & (g36) & (!reset) & (g598) & (!g1618)) + ((g34) & (g36) & (!reset) & (g598) & (g1618)));
	assign g7654 = (((!g832) & (g3077) & (!g1620)) + ((!g832) & (g3077) & (g1620)) + ((g832) & (!g3077) & (g1620)) + ((g832) & (g3077) & (g1620)));
	assign g1621 = (((!g34) & (!g36) & (!reset) & (g600) & (!g1620)) + ((!g34) & (!g36) & (!reset) & (g600) & (g1620)) + ((!g34) & (g36) & (!reset) & (!g600) & (g1620)) + ((!g34) & (g36) & (!reset) & (g600) & (g1620)) + ((g34) & (!g36) & (!reset) & (g600) & (!g1620)) + ((g34) & (!g36) & (!reset) & (g600) & (g1620)) + ((g34) & (g36) & (!reset) & (g600) & (!g1620)) + ((g34) & (g36) & (!reset) & (g600) & (g1620)));
	assign g7655 = (((!g832) & (g3079) & (!g1622)) + ((!g832) & (g3079) & (g1622)) + ((g832) & (!g3079) & (g1622)) + ((g832) & (g3079) & (g1622)));
	assign g1623 = (((!g34) & (!g36) & (!reset) & (g601) & (!g1622)) + ((!g34) & (!g36) & (!reset) & (g601) & (g1622)) + ((!g34) & (g36) & (!reset) & (!g601) & (g1622)) + ((!g34) & (g36) & (!reset) & (g601) & (g1622)) + ((g34) & (!g36) & (!reset) & (g601) & (!g1622)) + ((g34) & (!g36) & (!reset) & (g601) & (g1622)) + ((g34) & (g36) & (!reset) & (g601) & (!g1622)) + ((g34) & (g36) & (!reset) & (g601) & (g1622)));
	assign g7656 = (((!g832) & (g3081) & (!g1624)) + ((!g832) & (g3081) & (g1624)) + ((g832) & (!g3081) & (g1624)) + ((g832) & (g3081) & (g1624)));
	assign g1625 = (((!g34) & (!g36) & (!reset) & (g602) & (!g1624)) + ((!g34) & (!g36) & (!reset) & (g602) & (g1624)) + ((!g34) & (g36) & (!reset) & (!g602) & (g1624)) + ((!g34) & (g36) & (!reset) & (g602) & (g1624)) + ((g34) & (!g36) & (!reset) & (g602) & (!g1624)) + ((g34) & (!g36) & (!reset) & (g602) & (g1624)) + ((g34) & (g36) & (!reset) & (g602) & (!g1624)) + ((g34) & (g36) & (!reset) & (g602) & (g1624)));
	assign g7657 = (((!g832) & (g3083) & (!g1626)) + ((!g832) & (g3083) & (g1626)) + ((g832) & (!g3083) & (g1626)) + ((g832) & (g3083) & (g1626)));
	assign g1627 = (((!g34) & (!g36) & (!reset) & (g603) & (!g1626)) + ((!g34) & (!g36) & (!reset) & (g603) & (g1626)) + ((!g34) & (g36) & (!reset) & (!g603) & (g1626)) + ((!g34) & (g36) & (!reset) & (g603) & (g1626)) + ((g34) & (!g36) & (!reset) & (g603) & (!g1626)) + ((g34) & (!g36) & (!reset) & (g603) & (g1626)) + ((g34) & (g36) & (!reset) & (g603) & (!g1626)) + ((g34) & (g36) & (!reset) & (g603) & (g1626)));
	assign g7658 = (((!g832) & (g3085) & (!g1628)) + ((!g832) & (g3085) & (g1628)) + ((g832) & (!g3085) & (g1628)) + ((g832) & (g3085) & (g1628)));
	assign g1629 = (((!g34) & (!g36) & (!reset) & (g605) & (!g1628)) + ((!g34) & (!g36) & (!reset) & (g605) & (g1628)) + ((!g34) & (g36) & (!reset) & (!g605) & (g1628)) + ((!g34) & (g36) & (!reset) & (g605) & (g1628)) + ((g34) & (!g36) & (!reset) & (g605) & (!g1628)) + ((g34) & (!g36) & (!reset) & (g605) & (g1628)) + ((g34) & (g36) & (!reset) & (g605) & (!g1628)) + ((g34) & (g36) & (!reset) & (g605) & (g1628)));
	assign g7659 = (((!g832) & (g3087) & (!g1630)) + ((!g832) & (g3087) & (g1630)) + ((g832) & (!g3087) & (g1630)) + ((g832) & (g3087) & (g1630)));
	assign g1631 = (((!g34) & (!g36) & (!reset) & (g606) & (!g1630)) + ((!g34) & (!g36) & (!reset) & (g606) & (g1630)) + ((!g34) & (g36) & (!reset) & (!g606) & (g1630)) + ((!g34) & (g36) & (!reset) & (g606) & (g1630)) + ((g34) & (!g36) & (!reset) & (g606) & (!g1630)) + ((g34) & (!g36) & (!reset) & (g606) & (g1630)) + ((g34) & (g36) & (!reset) & (g606) & (!g1630)) + ((g34) & (g36) & (!reset) & (g606) & (g1630)));
	assign g7660 = (((!g832) & (g3089) & (!g1632)) + ((!g832) & (g3089) & (g1632)) + ((g832) & (!g3089) & (g1632)) + ((g832) & (g3089) & (g1632)));
	assign g1633 = (((!g34) & (!g36) & (!reset) & (g607) & (!g1632)) + ((!g34) & (!g36) & (!reset) & (g607) & (g1632)) + ((!g34) & (g36) & (!reset) & (!g607) & (g1632)) + ((!g34) & (g36) & (!reset) & (g607) & (g1632)) + ((g34) & (!g36) & (!reset) & (g607) & (!g1632)) + ((g34) & (!g36) & (!reset) & (g607) & (g1632)) + ((g34) & (g36) & (!reset) & (g607) & (!g1632)) + ((g34) & (g36) & (!reset) & (g607) & (g1632)));
	assign g7661 = (((!g832) & (g3091) & (!g1634)) + ((!g832) & (g3091) & (g1634)) + ((g832) & (!g3091) & (g1634)) + ((g832) & (g3091) & (g1634)));
	assign g1635 = (((!g34) & (!g36) & (!reset) & (g608) & (!g1634)) + ((!g34) & (!g36) & (!reset) & (g608) & (g1634)) + ((!g34) & (g36) & (!reset) & (!g608) & (g1634)) + ((!g34) & (g36) & (!reset) & (g608) & (g1634)) + ((g34) & (!g36) & (!reset) & (g608) & (!g1634)) + ((g34) & (!g36) & (!reset) & (g608) & (g1634)) + ((g34) & (g36) & (!reset) & (g608) & (!g1634)) + ((g34) & (g36) & (!reset) & (g608) & (g1634)));
	assign g7662 = (((!g832) & (g3092) & (!g1636)) + ((!g832) & (g3092) & (g1636)) + ((g832) & (!g3092) & (g1636)) + ((g832) & (g3092) & (g1636)));
	assign g1637 = (((!g34) & (!g36) & (!reset) & (g610) & (!g1636)) + ((!g34) & (!g36) & (!reset) & (g610) & (g1636)) + ((!g34) & (g36) & (!reset) & (!g610) & (g1636)) + ((!g34) & (g36) & (!reset) & (g610) & (g1636)) + ((g34) & (!g36) & (!reset) & (g610) & (!g1636)) + ((g34) & (!g36) & (!reset) & (g610) & (g1636)) + ((g34) & (g36) & (!reset) & (g610) & (!g1636)) + ((g34) & (g36) & (!reset) & (g610) & (g1636)));
	assign g7663 = (((!g832) & (g3094) & (!g1638)) + ((!g832) & (g3094) & (g1638)) + ((g832) & (!g3094) & (g1638)) + ((g832) & (g3094) & (g1638)));
	assign g1639 = (((!g34) & (!g36) & (!reset) & (g611) & (!g1638)) + ((!g34) & (!g36) & (!reset) & (g611) & (g1638)) + ((!g34) & (g36) & (!reset) & (!g611) & (g1638)) + ((!g34) & (g36) & (!reset) & (g611) & (g1638)) + ((g34) & (!g36) & (!reset) & (g611) & (!g1638)) + ((g34) & (!g36) & (!reset) & (g611) & (g1638)) + ((g34) & (g36) & (!reset) & (g611) & (!g1638)) + ((g34) & (g36) & (!reset) & (g611) & (g1638)));
	assign g7664 = (((!g832) & (g3096) & (!g1640)) + ((!g832) & (g3096) & (g1640)) + ((g832) & (!g3096) & (g1640)) + ((g832) & (g3096) & (g1640)));
	assign g1641 = (((!g34) & (!g36) & (!reset) & (g612) & (!g1640)) + ((!g34) & (!g36) & (!reset) & (g612) & (g1640)) + ((!g34) & (g36) & (!reset) & (!g612) & (g1640)) + ((!g34) & (g36) & (!reset) & (g612) & (g1640)) + ((g34) & (!g36) & (!reset) & (g612) & (!g1640)) + ((g34) & (!g36) & (!reset) & (g612) & (g1640)) + ((g34) & (g36) & (!reset) & (g612) & (!g1640)) + ((g34) & (g36) & (!reset) & (g612) & (g1640)));
	assign g7665 = (((!g832) & (g3098) & (!g1642)) + ((!g832) & (g3098) & (g1642)) + ((g832) & (!g3098) & (g1642)) + ((g832) & (g3098) & (g1642)));
	assign g1643 = (((!g34) & (!g36) & (!reset) & (g613) & (!g1642)) + ((!g34) & (!g36) & (!reset) & (g613) & (g1642)) + ((!g34) & (g36) & (!reset) & (!g613) & (g1642)) + ((!g34) & (g36) & (!reset) & (g613) & (g1642)) + ((g34) & (!g36) & (!reset) & (g613) & (!g1642)) + ((g34) & (!g36) & (!reset) & (g613) & (g1642)) + ((g34) & (g36) & (!reset) & (g613) & (!g1642)) + ((g34) & (g36) & (!reset) & (g613) & (g1642)));
	assign g7666 = (((!g2017) & (g3103) & (!g1644)) + ((!g2017) & (g3103) & (g1644)) + ((g2017) & (!g3103) & (g1644)) + ((g2017) & (g3103) & (g1644)));
	assign g1645 = (((!g827) & (!g593) & (!g616) & (!g1610) & (g1644) & (!g1611)) + ((!g827) & (!g593) & (!g616) & (!g1610) & (g1644) & (g1611)) + ((!g827) & (!g593) & (!g616) & (g1610) & (g1644) & (!g1611)) + ((!g827) & (!g593) & (!g616) & (g1610) & (g1644) & (g1611)) + ((!g827) & (!g593) & (g616) & (!g1610) & (g1644) & (!g1611)) + ((!g827) & (!g593) & (g616) & (!g1610) & (g1644) & (g1611)) + ((!g827) & (!g593) & (g616) & (g1610) & (g1644) & (!g1611)) + ((!g827) & (!g593) & (g616) & (g1610) & (g1644) & (g1611)) + ((!g827) & (g593) & (!g616) & (!g1610) & (g1644) & (!g1611)) + ((!g827) & (g593) & (!g616) & (!g1610) & (g1644) & (g1611)) + ((!g827) & (g593) & (!g616) & (g1610) & (g1644) & (!g1611)) + ((!g827) & (g593) & (!g616) & (g1610) & (g1644) & (g1611)) + ((!g827) & (g593) & (g616) & (!g1610) & (g1644) & (!g1611)) + ((!g827) & (g593) & (g616) & (!g1610) & (g1644) & (g1611)) + ((!g827) & (g593) & (g616) & (g1610) & (g1644) & (!g1611)) + ((!g827) & (g593) & (g616) & (g1610) & (g1644) & (g1611)) + ((g827) & (!g593) & (!g616) & (!g1610) & (g1644) & (!g1611)) + ((g827) & (!g593) & (!g616) & (!g1610) & (g1644) & (g1611)) + ((g827) & (!g593) & (!g616) & (g1610) & (!g1644) & (!g1611)) + ((g827) & (!g593) & (!g616) & (g1610) & (g1644) & (g1611)) + ((g827) & (!g593) & (g616) & (!g1610) & (!g1644) & (!g1611)) + ((g827) & (!g593) & (g616) & (!g1610) & (!g1644) & (g1611)) + ((g827) & (!g593) & (g616) & (g1610) & (!g1644) & (g1611)) + ((g827) & (!g593) & (g616) & (g1610) & (g1644) & (!g1611)) + ((g827) & (g593) & (!g616) & (!g1610) & (!g1644) & (!g1611)) + ((g827) & (g593) & (!g616) & (!g1610) & (g1644) & (g1611)) + ((g827) & (g593) & (!g616) & (g1610) & (!g1644) & (!g1611)) + ((g827) & (g593) & (!g616) & (g1610) & (!g1644) & (g1611)) + ((g827) & (g593) & (g616) & (!g1610) & (!g1644) & (g1611)) + ((g827) & (g593) & (g616) & (!g1610) & (g1644) & (!g1611)) + ((g827) & (g593) & (g616) & (g1610) & (g1644) & (!g1611)) + ((g827) & (g593) & (g616) & (g1610) & (g1644) & (g1611)));
	assign g1646 = (((!g34) & (!g36) & (!reset) & (g618) & (!g639)) + ((!g34) & (!g36) & (!reset) & (g618) & (g639)) + ((!g34) & (g36) & (!reset) & (!g618) & (g639)) + ((!g34) & (g36) & (!reset) & (g618) & (g639)) + ((g34) & (!g36) & (!reset) & (g618) & (!g639)) + ((g34) & (!g36) & (!reset) & (g618) & (g639)) + ((g34) & (g36) & (!reset) & (g618) & (!g639)) + ((g34) & (g36) & (!reset) & (g618) & (g639)));
	assign g7667 = (((!g832) & (g3105) & (!g1647)) + ((!g832) & (g3105) & (g1647)) + ((g832) & (!g3105) & (g1647)) + ((g832) & (g3105) & (g1647)));
	assign g1648 = (((!g34) & (!g36) & (!reset) & (g619) & (!g1647)) + ((!g34) & (!g36) & (!reset) & (g619) & (g1647)) + ((!g34) & (g36) & (!reset) & (!g619) & (g1647)) + ((!g34) & (g36) & (!reset) & (g619) & (g1647)) + ((g34) & (!g36) & (!reset) & (g619) & (!g1647)) + ((g34) & (!g36) & (!reset) & (g619) & (g1647)) + ((g34) & (g36) & (!reset) & (g619) & (!g1647)) + ((g34) & (g36) & (!reset) & (g619) & (g1647)));
	assign g7668 = (((!g832) & (g3108) & (!g1649)) + ((!g832) & (g3108) & (g1649)) + ((g832) & (!g3108) & (g1649)) + ((g832) & (g3108) & (g1649)));
	assign g1650 = (((!g34) & (!g36) & (!reset) & (g620) & (!g1649)) + ((!g34) & (!g36) & (!reset) & (g620) & (g1649)) + ((!g34) & (g36) & (!reset) & (!g620) & (g1649)) + ((!g34) & (g36) & (!reset) & (g620) & (g1649)) + ((g34) & (!g36) & (!reset) & (g620) & (!g1649)) + ((g34) & (!g36) & (!reset) & (g620) & (g1649)) + ((g34) & (g36) & (!reset) & (g620) & (!g1649)) + ((g34) & (g36) & (!reset) & (g620) & (g1649)));
	assign g7669 = (((!g832) & (g3110) & (!g1651)) + ((!g832) & (g3110) & (g1651)) + ((g832) & (!g3110) & (g1651)) + ((g832) & (g3110) & (g1651)));
	assign g1652 = (((!g34) & (!g36) & (!reset) & (g621) & (!g1651)) + ((!g34) & (!g36) & (!reset) & (g621) & (g1651)) + ((!g34) & (g36) & (!reset) & (!g621) & (g1651)) + ((!g34) & (g36) & (!reset) & (g621) & (g1651)) + ((g34) & (!g36) & (!reset) & (g621) & (!g1651)) + ((g34) & (!g36) & (!reset) & (g621) & (g1651)) + ((g34) & (g36) & (!reset) & (g621) & (!g1651)) + ((g34) & (g36) & (!reset) & (g621) & (g1651)));
	assign g7670 = (((!g832) & (g3112) & (!g1653)) + ((!g832) & (g3112) & (g1653)) + ((g832) & (!g3112) & (g1653)) + ((g832) & (g3112) & (g1653)));
	assign g1654 = (((!g34) & (!g36) & (!reset) & (g623) & (!g1653)) + ((!g34) & (!g36) & (!reset) & (g623) & (g1653)) + ((!g34) & (g36) & (!reset) & (!g623) & (g1653)) + ((!g34) & (g36) & (!reset) & (g623) & (g1653)) + ((g34) & (!g36) & (!reset) & (g623) & (!g1653)) + ((g34) & (!g36) & (!reset) & (g623) & (g1653)) + ((g34) & (g36) & (!reset) & (g623) & (!g1653)) + ((g34) & (g36) & (!reset) & (g623) & (g1653)));
	assign g7671 = (((!g832) & (g3115) & (!g1655)) + ((!g832) & (g3115) & (g1655)) + ((g832) & (!g3115) & (g1655)) + ((g832) & (g3115) & (g1655)));
	assign g1656 = (((!g34) & (!g36) & (!reset) & (g624) & (!g1655)) + ((!g34) & (!g36) & (!reset) & (g624) & (g1655)) + ((!g34) & (g36) & (!reset) & (!g624) & (g1655)) + ((!g34) & (g36) & (!reset) & (g624) & (g1655)) + ((g34) & (!g36) & (!reset) & (g624) & (!g1655)) + ((g34) & (!g36) & (!reset) & (g624) & (g1655)) + ((g34) & (g36) & (!reset) & (g624) & (!g1655)) + ((g34) & (g36) & (!reset) & (g624) & (g1655)));
	assign g7672 = (((!g832) & (g3118) & (!g1657)) + ((!g832) & (g3118) & (g1657)) + ((g832) & (!g3118) & (g1657)) + ((g832) & (g3118) & (g1657)));
	assign g1658 = (((!g34) & (!g36) & (!reset) & (g625) & (!g1657)) + ((!g34) & (!g36) & (!reset) & (g625) & (g1657)) + ((!g34) & (g36) & (!reset) & (!g625) & (g1657)) + ((!g34) & (g36) & (!reset) & (g625) & (g1657)) + ((g34) & (!g36) & (!reset) & (g625) & (!g1657)) + ((g34) & (!g36) & (!reset) & (g625) & (g1657)) + ((g34) & (g36) & (!reset) & (g625) & (!g1657)) + ((g34) & (g36) & (!reset) & (g625) & (g1657)));
	assign g7673 = (((!g832) & (g3121) & (!g1659)) + ((!g832) & (g3121) & (g1659)) + ((g832) & (!g3121) & (g1659)) + ((g832) & (g3121) & (g1659)));
	assign g1660 = (((!g34) & (!g36) & (!reset) & (g626) & (!g1659)) + ((!g34) & (!g36) & (!reset) & (g626) & (g1659)) + ((!g34) & (g36) & (!reset) & (!g626) & (g1659)) + ((!g34) & (g36) & (!reset) & (g626) & (g1659)) + ((g34) & (!g36) & (!reset) & (g626) & (!g1659)) + ((g34) & (!g36) & (!reset) & (g626) & (g1659)) + ((g34) & (g36) & (!reset) & (g626) & (!g1659)) + ((g34) & (g36) & (!reset) & (g626) & (g1659)));
	assign g7674 = (((!g832) & (g3124) & (!g1661)) + ((!g832) & (g3124) & (g1661)) + ((g832) & (!g3124) & (g1661)) + ((g832) & (g3124) & (g1661)));
	assign g1662 = (((!g34) & (!g36) & (!reset) & (g628) & (!g1661)) + ((!g34) & (!g36) & (!reset) & (g628) & (g1661)) + ((!g34) & (g36) & (!reset) & (!g628) & (g1661)) + ((!g34) & (g36) & (!reset) & (g628) & (g1661)) + ((g34) & (!g36) & (!reset) & (g628) & (!g1661)) + ((g34) & (!g36) & (!reset) & (g628) & (g1661)) + ((g34) & (g36) & (!reset) & (g628) & (!g1661)) + ((g34) & (g36) & (!reset) & (g628) & (g1661)));
	assign g7675 = (((!g832) & (g3127) & (!g1663)) + ((!g832) & (g3127) & (g1663)) + ((g832) & (!g3127) & (g1663)) + ((g832) & (g3127) & (g1663)));
	assign g1664 = (((!g34) & (!g36) & (!reset) & (g629) & (!g1663)) + ((!g34) & (!g36) & (!reset) & (g629) & (g1663)) + ((!g34) & (g36) & (!reset) & (!g629) & (g1663)) + ((!g34) & (g36) & (!reset) & (g629) & (g1663)) + ((g34) & (!g36) & (!reset) & (g629) & (!g1663)) + ((g34) & (!g36) & (!reset) & (g629) & (g1663)) + ((g34) & (g36) & (!reset) & (g629) & (!g1663)) + ((g34) & (g36) & (!reset) & (g629) & (g1663)));
	assign g7676 = (((!g832) & (g3130) & (!g1665)) + ((!g832) & (g3130) & (g1665)) + ((g832) & (!g3130) & (g1665)) + ((g832) & (g3130) & (g1665)));
	assign g1666 = (((!g34) & (!g36) & (!reset) & (g630) & (!g1665)) + ((!g34) & (!g36) & (!reset) & (g630) & (g1665)) + ((!g34) & (g36) & (!reset) & (!g630) & (g1665)) + ((!g34) & (g36) & (!reset) & (g630) & (g1665)) + ((g34) & (!g36) & (!reset) & (g630) & (!g1665)) + ((g34) & (!g36) & (!reset) & (g630) & (g1665)) + ((g34) & (g36) & (!reset) & (g630) & (!g1665)) + ((g34) & (g36) & (!reset) & (g630) & (g1665)));
	assign g7677 = (((!g832) & (g3133) & (!g1667)) + ((!g832) & (g3133) & (g1667)) + ((g832) & (!g3133) & (g1667)) + ((g832) & (g3133) & (g1667)));
	assign g1668 = (((!g34) & (!g36) & (!reset) & (g631) & (!g1667)) + ((!g34) & (!g36) & (!reset) & (g631) & (g1667)) + ((!g34) & (g36) & (!reset) & (!g631) & (g1667)) + ((!g34) & (g36) & (!reset) & (g631) & (g1667)) + ((g34) & (!g36) & (!reset) & (g631) & (!g1667)) + ((g34) & (!g36) & (!reset) & (g631) & (g1667)) + ((g34) & (g36) & (!reset) & (g631) & (!g1667)) + ((g34) & (g36) & (!reset) & (g631) & (g1667)));
	assign g7678 = (((!g832) & (g3135) & (!g1669)) + ((!g832) & (g3135) & (g1669)) + ((g832) & (!g3135) & (g1669)) + ((g832) & (g3135) & (g1669)));
	assign g1670 = (((!g34) & (!g36) & (!reset) & (g633) & (!g1669)) + ((!g34) & (!g36) & (!reset) & (g633) & (g1669)) + ((!g34) & (g36) & (!reset) & (!g633) & (g1669)) + ((!g34) & (g36) & (!reset) & (g633) & (g1669)) + ((g34) & (!g36) & (!reset) & (g633) & (!g1669)) + ((g34) & (!g36) & (!reset) & (g633) & (g1669)) + ((g34) & (g36) & (!reset) & (g633) & (!g1669)) + ((g34) & (g36) & (!reset) & (g633) & (g1669)));
	assign g7679 = (((!g832) & (g3138) & (!g1671)) + ((!g832) & (g3138) & (g1671)) + ((g832) & (!g3138) & (g1671)) + ((g832) & (g3138) & (g1671)));
	assign g1672 = (((!g34) & (!g36) & (!reset) & (g634) & (!g1671)) + ((!g34) & (!g36) & (!reset) & (g634) & (g1671)) + ((!g34) & (g36) & (!reset) & (!g634) & (g1671)) + ((!g34) & (g36) & (!reset) & (g634) & (g1671)) + ((g34) & (!g36) & (!reset) & (g634) & (!g1671)) + ((g34) & (!g36) & (!reset) & (g634) & (g1671)) + ((g34) & (g36) & (!reset) & (g634) & (!g1671)) + ((g34) & (g36) & (!reset) & (g634) & (g1671)));
	assign g7680 = (((!g832) & (g3141) & (!g1673)) + ((!g832) & (g3141) & (g1673)) + ((g832) & (!g3141) & (g1673)) + ((g832) & (g3141) & (g1673)));
	assign g1674 = (((!g34) & (!g36) & (!reset) & (g635) & (!g1673)) + ((!g34) & (!g36) & (!reset) & (g635) & (g1673)) + ((!g34) & (g36) & (!reset) & (!g635) & (g1673)) + ((!g34) & (g36) & (!reset) & (g635) & (g1673)) + ((g34) & (!g36) & (!reset) & (g635) & (!g1673)) + ((g34) & (!g36) & (!reset) & (g635) & (g1673)) + ((g34) & (g36) & (!reset) & (g635) & (!g1673)) + ((g34) & (g36) & (!reset) & (g635) & (g1673)));
	assign g7681 = (((!g832) & (g3144) & (!g1675)) + ((!g832) & (g3144) & (g1675)) + ((g832) & (!g3144) & (g1675)) + ((g832) & (g3144) & (g1675)));
	assign g1676 = (((!g34) & (!g36) & (!reset) & (g636) & (!g1675)) + ((!g34) & (!g36) & (!reset) & (g636) & (g1675)) + ((!g34) & (g36) & (!reset) & (!g636) & (g1675)) + ((!g34) & (g36) & (!reset) & (g636) & (g1675)) + ((g34) & (!g36) & (!reset) & (g636) & (!g1675)) + ((g34) & (!g36) & (!reset) & (g636) & (g1675)) + ((g34) & (g36) & (!reset) & (g636) & (!g1675)) + ((g34) & (g36) & (!reset) & (g636) & (g1675)));
	assign g7682 = (((!g2017) & (g3147) & (!g1677)) + ((!g2017) & (g3147) & (g1677)) + ((g2017) & (!g3147) & (g1677)) + ((g2017) & (g3147) & (g1677)));
	assign g1678 = (((!g593) & (!g616) & (g1610) & (g1644) & (!g1611)) + ((!g593) & (g616) & (!g1610) & (g1644) & (!g1611)) + ((!g593) & (g616) & (!g1610) & (g1644) & (g1611)) + ((!g593) & (g616) & (g1610) & (!g1644) & (!g1611)) + ((!g593) & (g616) & (g1610) & (g1644) & (!g1611)) + ((!g593) & (g616) & (g1610) & (g1644) & (g1611)) + ((g593) & (!g616) & (!g1610) & (g1644) & (!g1611)) + ((g593) & (!g616) & (g1610) & (g1644) & (!g1611)) + ((g593) & (!g616) & (g1610) & (g1644) & (g1611)) + ((g593) & (g616) & (!g1610) & (!g1644) & (!g1611)) + ((g593) & (g616) & (!g1610) & (g1644) & (!g1611)) + ((g593) & (g616) & (!g1610) & (g1644) & (g1611)) + ((g593) & (g616) & (g1610) & (!g1644) & (!g1611)) + ((g593) & (g616) & (g1610) & (!g1644) & (g1611)) + ((g593) & (g616) & (g1610) & (g1644) & (!g1611)) + ((g593) & (g616) & (g1610) & (g1644) & (g1611)));
	assign g1679 = (((!g827) & (!g639) & (g1677) & (!g1678)) + ((!g827) & (!g639) & (g1677) & (g1678)) + ((!g827) & (g639) & (g1677) & (!g1678)) + ((!g827) & (g639) & (g1677) & (g1678)) + ((g827) & (!g639) & (!g1677) & (g1678)) + ((g827) & (!g639) & (g1677) & (!g1678)) + ((g827) & (g639) & (!g1677) & (!g1678)) + ((g827) & (g639) & (g1677) & (g1678)));
	assign g1680 = (((!g34) & (!g36) & (!reset) & (g641) & (!g662)) + ((!g34) & (!g36) & (!reset) & (g641) & (g662)) + ((!g34) & (g36) & (!reset) & (!g641) & (g662)) + ((!g34) & (g36) & (!reset) & (g641) & (g662)) + ((g34) & (!g36) & (!reset) & (g641) & (!g662)) + ((g34) & (!g36) & (!reset) & (g641) & (g662)) + ((g34) & (g36) & (!reset) & (g641) & (!g662)) + ((g34) & (g36) & (!reset) & (g641) & (g662)));
	assign g7683 = (((!g832) & (g3148) & (!g1681)) + ((!g832) & (g3148) & (g1681)) + ((g832) & (!g3148) & (g1681)) + ((g832) & (g3148) & (g1681)));
	assign g1682 = (((!g34) & (!g36) & (!reset) & (g642) & (!g1681)) + ((!g34) & (!g36) & (!reset) & (g642) & (g1681)) + ((!g34) & (g36) & (!reset) & (!g642) & (g1681)) + ((!g34) & (g36) & (!reset) & (g642) & (g1681)) + ((g34) & (!g36) & (!reset) & (g642) & (!g1681)) + ((g34) & (!g36) & (!reset) & (g642) & (g1681)) + ((g34) & (g36) & (!reset) & (g642) & (!g1681)) + ((g34) & (g36) & (!reset) & (g642) & (g1681)));
	assign g7684 = (((!g832) & (g3150) & (!g1683)) + ((!g832) & (g3150) & (g1683)) + ((g832) & (!g3150) & (g1683)) + ((g832) & (g3150) & (g1683)));
	assign g1684 = (((!g34) & (!g36) & (!reset) & (g643) & (!g1683)) + ((!g34) & (!g36) & (!reset) & (g643) & (g1683)) + ((!g34) & (g36) & (!reset) & (!g643) & (g1683)) + ((!g34) & (g36) & (!reset) & (g643) & (g1683)) + ((g34) & (!g36) & (!reset) & (g643) & (!g1683)) + ((g34) & (!g36) & (!reset) & (g643) & (g1683)) + ((g34) & (g36) & (!reset) & (g643) & (!g1683)) + ((g34) & (g36) & (!reset) & (g643) & (g1683)));
	assign g7685 = (((!g832) & (g3151) & (!g1685)) + ((!g832) & (g3151) & (g1685)) + ((g832) & (!g3151) & (g1685)) + ((g832) & (g3151) & (g1685)));
	assign g1686 = (((!g34) & (!g36) & (!reset) & (g644) & (!g1685)) + ((!g34) & (!g36) & (!reset) & (g644) & (g1685)) + ((!g34) & (g36) & (!reset) & (!g644) & (g1685)) + ((!g34) & (g36) & (!reset) & (g644) & (g1685)) + ((g34) & (!g36) & (!reset) & (g644) & (!g1685)) + ((g34) & (!g36) & (!reset) & (g644) & (g1685)) + ((g34) & (g36) & (!reset) & (g644) & (!g1685)) + ((g34) & (g36) & (!reset) & (g644) & (g1685)));
	assign g7686 = (((!g832) & (g3152) & (!g1687)) + ((!g832) & (g3152) & (g1687)) + ((g832) & (!g3152) & (g1687)) + ((g832) & (g3152) & (g1687)));
	assign g1688 = (((!g34) & (!g36) & (!reset) & (g646) & (!g1687)) + ((!g34) & (!g36) & (!reset) & (g646) & (g1687)) + ((!g34) & (g36) & (!reset) & (!g646) & (g1687)) + ((!g34) & (g36) & (!reset) & (g646) & (g1687)) + ((g34) & (!g36) & (!reset) & (g646) & (!g1687)) + ((g34) & (!g36) & (!reset) & (g646) & (g1687)) + ((g34) & (g36) & (!reset) & (g646) & (!g1687)) + ((g34) & (g36) & (!reset) & (g646) & (g1687)));
	assign g7687 = (((!g832) & (g3154) & (!g1689)) + ((!g832) & (g3154) & (g1689)) + ((g832) & (!g3154) & (g1689)) + ((g832) & (g3154) & (g1689)));
	assign g1690 = (((!g34) & (!g36) & (!reset) & (g647) & (!g1689)) + ((!g34) & (!g36) & (!reset) & (g647) & (g1689)) + ((!g34) & (g36) & (!reset) & (!g647) & (g1689)) + ((!g34) & (g36) & (!reset) & (g647) & (g1689)) + ((g34) & (!g36) & (!reset) & (g647) & (!g1689)) + ((g34) & (!g36) & (!reset) & (g647) & (g1689)) + ((g34) & (g36) & (!reset) & (g647) & (!g1689)) + ((g34) & (g36) & (!reset) & (g647) & (g1689)));
	assign g7688 = (((!g832) & (g3156) & (!g1691)) + ((!g832) & (g3156) & (g1691)) + ((g832) & (!g3156) & (g1691)) + ((g832) & (g3156) & (g1691)));
	assign g1692 = (((!g34) & (!g36) & (!reset) & (g648) & (!g1691)) + ((!g34) & (!g36) & (!reset) & (g648) & (g1691)) + ((!g34) & (g36) & (!reset) & (!g648) & (g1691)) + ((!g34) & (g36) & (!reset) & (g648) & (g1691)) + ((g34) & (!g36) & (!reset) & (g648) & (!g1691)) + ((g34) & (!g36) & (!reset) & (g648) & (g1691)) + ((g34) & (g36) & (!reset) & (g648) & (!g1691)) + ((g34) & (g36) & (!reset) & (g648) & (g1691)));
	assign g7689 = (((!g832) & (g3158) & (!g1693)) + ((!g832) & (g3158) & (g1693)) + ((g832) & (!g3158) & (g1693)) + ((g832) & (g3158) & (g1693)));
	assign g1694 = (((!g34) & (!g36) & (!reset) & (g649) & (!g1693)) + ((!g34) & (!g36) & (!reset) & (g649) & (g1693)) + ((!g34) & (g36) & (!reset) & (!g649) & (g1693)) + ((!g34) & (g36) & (!reset) & (g649) & (g1693)) + ((g34) & (!g36) & (!reset) & (g649) & (!g1693)) + ((g34) & (!g36) & (!reset) & (g649) & (g1693)) + ((g34) & (g36) & (!reset) & (g649) & (!g1693)) + ((g34) & (g36) & (!reset) & (g649) & (g1693)));
	assign g7690 = (((!g832) & (g3160) & (!g1695)) + ((!g832) & (g3160) & (g1695)) + ((g832) & (!g3160) & (g1695)) + ((g832) & (g3160) & (g1695)));
	assign g1696 = (((!g34) & (!g36) & (!reset) & (g651) & (!g1695)) + ((!g34) & (!g36) & (!reset) & (g651) & (g1695)) + ((!g34) & (g36) & (!reset) & (!g651) & (g1695)) + ((!g34) & (g36) & (!reset) & (g651) & (g1695)) + ((g34) & (!g36) & (!reset) & (g651) & (!g1695)) + ((g34) & (!g36) & (!reset) & (g651) & (g1695)) + ((g34) & (g36) & (!reset) & (g651) & (!g1695)) + ((g34) & (g36) & (!reset) & (g651) & (g1695)));
	assign g7691 = (((!g832) & (g3162) & (!g1697)) + ((!g832) & (g3162) & (g1697)) + ((g832) & (!g3162) & (g1697)) + ((g832) & (g3162) & (g1697)));
	assign g1698 = (((!g34) & (!g36) & (!reset) & (g652) & (!g1697)) + ((!g34) & (!g36) & (!reset) & (g652) & (g1697)) + ((!g34) & (g36) & (!reset) & (!g652) & (g1697)) + ((!g34) & (g36) & (!reset) & (g652) & (g1697)) + ((g34) & (!g36) & (!reset) & (g652) & (!g1697)) + ((g34) & (!g36) & (!reset) & (g652) & (g1697)) + ((g34) & (g36) & (!reset) & (g652) & (!g1697)) + ((g34) & (g36) & (!reset) & (g652) & (g1697)));
	assign g7692 = (((!g832) & (g3164) & (!g1699)) + ((!g832) & (g3164) & (g1699)) + ((g832) & (!g3164) & (g1699)) + ((g832) & (g3164) & (g1699)));
	assign g1700 = (((!g34) & (!g36) & (!reset) & (g653) & (!g1699)) + ((!g34) & (!g36) & (!reset) & (g653) & (g1699)) + ((!g34) & (g36) & (!reset) & (!g653) & (g1699)) + ((!g34) & (g36) & (!reset) & (g653) & (g1699)) + ((g34) & (!g36) & (!reset) & (g653) & (!g1699)) + ((g34) & (!g36) & (!reset) & (g653) & (g1699)) + ((g34) & (g36) & (!reset) & (g653) & (!g1699)) + ((g34) & (g36) & (!reset) & (g653) & (g1699)));
	assign g7693 = (((!g832) & (g3166) & (!g1701)) + ((!g832) & (g3166) & (g1701)) + ((g832) & (!g3166) & (g1701)) + ((g832) & (g3166) & (g1701)));
	assign g1702 = (((!g34) & (!g36) & (!reset) & (g654) & (!g1701)) + ((!g34) & (!g36) & (!reset) & (g654) & (g1701)) + ((!g34) & (g36) & (!reset) & (!g654) & (g1701)) + ((!g34) & (g36) & (!reset) & (g654) & (g1701)) + ((g34) & (!g36) & (!reset) & (g654) & (!g1701)) + ((g34) & (!g36) & (!reset) & (g654) & (g1701)) + ((g34) & (g36) & (!reset) & (g654) & (!g1701)) + ((g34) & (g36) & (!reset) & (g654) & (g1701)));
	assign g7694 = (((!g832) & (g3167) & (!g1703)) + ((!g832) & (g3167) & (g1703)) + ((g832) & (!g3167) & (g1703)) + ((g832) & (g3167) & (g1703)));
	assign g1704 = (((!g34) & (!g36) & (!reset) & (g656) & (!g1703)) + ((!g34) & (!g36) & (!reset) & (g656) & (g1703)) + ((!g34) & (g36) & (!reset) & (!g656) & (g1703)) + ((!g34) & (g36) & (!reset) & (g656) & (g1703)) + ((g34) & (!g36) & (!reset) & (g656) & (!g1703)) + ((g34) & (!g36) & (!reset) & (g656) & (g1703)) + ((g34) & (g36) & (!reset) & (g656) & (!g1703)) + ((g34) & (g36) & (!reset) & (g656) & (g1703)));
	assign g7695 = (((!g832) & (g3169) & (!g1705)) + ((!g832) & (g3169) & (g1705)) + ((g832) & (!g3169) & (g1705)) + ((g832) & (g3169) & (g1705)));
	assign g1706 = (((!g34) & (!g36) & (!reset) & (g657) & (!g1705)) + ((!g34) & (!g36) & (!reset) & (g657) & (g1705)) + ((!g34) & (g36) & (!reset) & (!g657) & (g1705)) + ((!g34) & (g36) & (!reset) & (g657) & (g1705)) + ((g34) & (!g36) & (!reset) & (g657) & (!g1705)) + ((g34) & (!g36) & (!reset) & (g657) & (g1705)) + ((g34) & (g36) & (!reset) & (g657) & (!g1705)) + ((g34) & (g36) & (!reset) & (g657) & (g1705)));
	assign g7696 = (((!g832) & (g3171) & (!g1707)) + ((!g832) & (g3171) & (g1707)) + ((g832) & (!g3171) & (g1707)) + ((g832) & (g3171) & (g1707)));
	assign g1708 = (((!g34) & (!g36) & (!reset) & (g658) & (!g1707)) + ((!g34) & (!g36) & (!reset) & (g658) & (g1707)) + ((!g34) & (g36) & (!reset) & (!g658) & (g1707)) + ((!g34) & (g36) & (!reset) & (g658) & (g1707)) + ((g34) & (!g36) & (!reset) & (g658) & (!g1707)) + ((g34) & (!g36) & (!reset) & (g658) & (g1707)) + ((g34) & (g36) & (!reset) & (g658) & (!g1707)) + ((g34) & (g36) & (!reset) & (g658) & (g1707)));
	assign g7697 = (((!g832) & (g3173) & (!g1709)) + ((!g832) & (g3173) & (g1709)) + ((g832) & (!g3173) & (g1709)) + ((g832) & (g3173) & (g1709)));
	assign g1710 = (((!g34) & (!g36) & (!reset) & (g659) & (!g1709)) + ((!g34) & (!g36) & (!reset) & (g659) & (g1709)) + ((!g34) & (g36) & (!reset) & (!g659) & (g1709)) + ((!g34) & (g36) & (!reset) & (g659) & (g1709)) + ((g34) & (!g36) & (!reset) & (g659) & (!g1709)) + ((g34) & (!g36) & (!reset) & (g659) & (g1709)) + ((g34) & (g36) & (!reset) & (g659) & (!g1709)) + ((g34) & (g36) & (!reset) & (g659) & (g1709)));
	assign g7698 = (((!g2017) & (g7101) & (!g1711)) + ((!g2017) & (g7101) & (g1711)) + ((g2017) & (!g7101) & (g1711)) + ((g2017) & (g7101) & (g1711)));
	assign g1712 = (((!g827) & (!g639) & (!g662) & (!g1677) & (g1711) & (!g1678)) + ((!g827) & (!g639) & (!g662) & (!g1677) & (g1711) & (g1678)) + ((!g827) & (!g639) & (!g662) & (g1677) & (g1711) & (!g1678)) + ((!g827) & (!g639) & (!g662) & (g1677) & (g1711) & (g1678)) + ((!g827) & (!g639) & (g662) & (!g1677) & (g1711) & (!g1678)) + ((!g827) & (!g639) & (g662) & (!g1677) & (g1711) & (g1678)) + ((!g827) & (!g639) & (g662) & (g1677) & (g1711) & (!g1678)) + ((!g827) & (!g639) & (g662) & (g1677) & (g1711) & (g1678)) + ((!g827) & (g639) & (!g662) & (!g1677) & (g1711) & (!g1678)) + ((!g827) & (g639) & (!g662) & (!g1677) & (g1711) & (g1678)) + ((!g827) & (g639) & (!g662) & (g1677) & (g1711) & (!g1678)) + ((!g827) & (g639) & (!g662) & (g1677) & (g1711) & (g1678)) + ((!g827) & (g639) & (g662) & (!g1677) & (g1711) & (!g1678)) + ((!g827) & (g639) & (g662) & (!g1677) & (g1711) & (g1678)) + ((!g827) & (g639) & (g662) & (g1677) & (g1711) & (!g1678)) + ((!g827) & (g639) & (g662) & (g1677) & (g1711) & (g1678)) + ((g827) & (!g639) & (!g662) & (!g1677) & (g1711) & (!g1678)) + ((g827) & (!g639) & (!g662) & (!g1677) & (g1711) & (g1678)) + ((g827) & (!g639) & (!g662) & (g1677) & (!g1711) & (g1678)) + ((g827) & (!g639) & (!g662) & (g1677) & (g1711) & (!g1678)) + ((g827) & (!g639) & (g662) & (!g1677) & (!g1711) & (!g1678)) + ((g827) & (!g639) & (g662) & (!g1677) & (!g1711) & (g1678)) + ((g827) & (!g639) & (g662) & (g1677) & (!g1711) & (!g1678)) + ((g827) & (!g639) & (g662) & (g1677) & (g1711) & (g1678)) + ((g827) & (g639) & (!g662) & (!g1677) & (!g1711) & (g1678)) + ((g827) & (g639) & (!g662) & (!g1677) & (g1711) & (!g1678)) + ((g827) & (g639) & (!g662) & (g1677) & (!g1711) & (!g1678)) + ((g827) & (g639) & (!g662) & (g1677) & (!g1711) & (g1678)) + ((g827) & (g639) & (g662) & (!g1677) & (!g1711) & (!g1678)) + ((g827) & (g639) & (g662) & (!g1677) & (g1711) & (g1678)) + ((g827) & (g639) & (g662) & (g1677) & (g1711) & (!g1678)) + ((g827) & (g639) & (g662) & (g1677) & (g1711) & (g1678)));
	assign g1713 = (((!g34) & (!g36) & (!reset) & (g664) & (!g685)) + ((!g34) & (!g36) & (!reset) & (g664) & (g685)) + ((!g34) & (g36) & (!reset) & (!g664) & (g685)) + ((!g34) & (g36) & (!reset) & (g664) & (g685)) + ((g34) & (!g36) & (!reset) & (g664) & (!g685)) + ((g34) & (!g36) & (!reset) & (g664) & (g685)) + ((g34) & (g36) & (!reset) & (g664) & (!g685)) + ((g34) & (g36) & (!reset) & (g664) & (g685)));
	assign g7699 = (((!g832) & (g3176) & (!g1714)) + ((!g832) & (g3176) & (g1714)) + ((g832) & (!g3176) & (g1714)) + ((g832) & (g3176) & (g1714)));
	assign g1715 = (((!g34) & (!g36) & (!reset) & (g665) & (!g1714)) + ((!g34) & (!g36) & (!reset) & (g665) & (g1714)) + ((!g34) & (g36) & (!reset) & (!g665) & (g1714)) + ((!g34) & (g36) & (!reset) & (g665) & (g1714)) + ((g34) & (!g36) & (!reset) & (g665) & (!g1714)) + ((g34) & (!g36) & (!reset) & (g665) & (g1714)) + ((g34) & (g36) & (!reset) & (g665) & (!g1714)) + ((g34) & (g36) & (!reset) & (g665) & (g1714)));
	assign g7700 = (((!g832) & (g3179) & (!g1716)) + ((!g832) & (g3179) & (g1716)) + ((g832) & (!g3179) & (g1716)) + ((g832) & (g3179) & (g1716)));
	assign g1717 = (((!g34) & (!g36) & (!reset) & (g666) & (!g1716)) + ((!g34) & (!g36) & (!reset) & (g666) & (g1716)) + ((!g34) & (g36) & (!reset) & (!g666) & (g1716)) + ((!g34) & (g36) & (!reset) & (g666) & (g1716)) + ((g34) & (!g36) & (!reset) & (g666) & (!g1716)) + ((g34) & (!g36) & (!reset) & (g666) & (g1716)) + ((g34) & (g36) & (!reset) & (g666) & (!g1716)) + ((g34) & (g36) & (!reset) & (g666) & (g1716)));
	assign g7701 = (((!g832) & (g3181) & (!g1718)) + ((!g832) & (g3181) & (g1718)) + ((g832) & (!g3181) & (g1718)) + ((g832) & (g3181) & (g1718)));
	assign g1719 = (((!g34) & (!g36) & (!reset) & (g667) & (!g1718)) + ((!g34) & (!g36) & (!reset) & (g667) & (g1718)) + ((!g34) & (g36) & (!reset) & (!g667) & (g1718)) + ((!g34) & (g36) & (!reset) & (g667) & (g1718)) + ((g34) & (!g36) & (!reset) & (g667) & (!g1718)) + ((g34) & (!g36) & (!reset) & (g667) & (g1718)) + ((g34) & (g36) & (!reset) & (g667) & (!g1718)) + ((g34) & (g36) & (!reset) & (g667) & (g1718)));
	assign g7702 = (((!g832) & (g3183) & (!g1720)) + ((!g832) & (g3183) & (g1720)) + ((g832) & (!g3183) & (g1720)) + ((g832) & (g3183) & (g1720)));
	assign g1721 = (((!g34) & (!g36) & (!reset) & (g669) & (!g1720)) + ((!g34) & (!g36) & (!reset) & (g669) & (g1720)) + ((!g34) & (g36) & (!reset) & (!g669) & (g1720)) + ((!g34) & (g36) & (!reset) & (g669) & (g1720)) + ((g34) & (!g36) & (!reset) & (g669) & (!g1720)) + ((g34) & (!g36) & (!reset) & (g669) & (g1720)) + ((g34) & (g36) & (!reset) & (g669) & (!g1720)) + ((g34) & (g36) & (!reset) & (g669) & (g1720)));
	assign g7703 = (((!g832) & (g3186) & (!g1722)) + ((!g832) & (g3186) & (g1722)) + ((g832) & (!g3186) & (g1722)) + ((g832) & (g3186) & (g1722)));
	assign g1723 = (((!g34) & (!g36) & (!reset) & (g670) & (!g1722)) + ((!g34) & (!g36) & (!reset) & (g670) & (g1722)) + ((!g34) & (g36) & (!reset) & (!g670) & (g1722)) + ((!g34) & (g36) & (!reset) & (g670) & (g1722)) + ((g34) & (!g36) & (!reset) & (g670) & (!g1722)) + ((g34) & (!g36) & (!reset) & (g670) & (g1722)) + ((g34) & (g36) & (!reset) & (g670) & (!g1722)) + ((g34) & (g36) & (!reset) & (g670) & (g1722)));
	assign g7704 = (((!g832) & (g3189) & (!g1724)) + ((!g832) & (g3189) & (g1724)) + ((g832) & (!g3189) & (g1724)) + ((g832) & (g3189) & (g1724)));
	assign g1725 = (((!g34) & (!g36) & (!reset) & (g671) & (!g1724)) + ((!g34) & (!g36) & (!reset) & (g671) & (g1724)) + ((!g34) & (g36) & (!reset) & (!g671) & (g1724)) + ((!g34) & (g36) & (!reset) & (g671) & (g1724)) + ((g34) & (!g36) & (!reset) & (g671) & (!g1724)) + ((g34) & (!g36) & (!reset) & (g671) & (g1724)) + ((g34) & (g36) & (!reset) & (g671) & (!g1724)) + ((g34) & (g36) & (!reset) & (g671) & (g1724)));
	assign g7705 = (((!g832) & (g3192) & (!g1726)) + ((!g832) & (g3192) & (g1726)) + ((g832) & (!g3192) & (g1726)) + ((g832) & (g3192) & (g1726)));
	assign g1727 = (((!g34) & (!g36) & (!reset) & (g672) & (!g1726)) + ((!g34) & (!g36) & (!reset) & (g672) & (g1726)) + ((!g34) & (g36) & (!reset) & (!g672) & (g1726)) + ((!g34) & (g36) & (!reset) & (g672) & (g1726)) + ((g34) & (!g36) & (!reset) & (g672) & (!g1726)) + ((g34) & (!g36) & (!reset) & (g672) & (g1726)) + ((g34) & (g36) & (!reset) & (g672) & (!g1726)) + ((g34) & (g36) & (!reset) & (g672) & (g1726)));
	assign g7706 = (((!g832) & (g3195) & (!g1728)) + ((!g832) & (g3195) & (g1728)) + ((g832) & (!g3195) & (g1728)) + ((g832) & (g3195) & (g1728)));
	assign g1729 = (((!g34) & (!g36) & (!reset) & (g674) & (!g1728)) + ((!g34) & (!g36) & (!reset) & (g674) & (g1728)) + ((!g34) & (g36) & (!reset) & (!g674) & (g1728)) + ((!g34) & (g36) & (!reset) & (g674) & (g1728)) + ((g34) & (!g36) & (!reset) & (g674) & (!g1728)) + ((g34) & (!g36) & (!reset) & (g674) & (g1728)) + ((g34) & (g36) & (!reset) & (g674) & (!g1728)) + ((g34) & (g36) & (!reset) & (g674) & (g1728)));
	assign g7707 = (((!g832) & (g3198) & (!g1730)) + ((!g832) & (g3198) & (g1730)) + ((g832) & (!g3198) & (g1730)) + ((g832) & (g3198) & (g1730)));
	assign g1731 = (((!g34) & (!g36) & (!reset) & (g675) & (!g1730)) + ((!g34) & (!g36) & (!reset) & (g675) & (g1730)) + ((!g34) & (g36) & (!reset) & (!g675) & (g1730)) + ((!g34) & (g36) & (!reset) & (g675) & (g1730)) + ((g34) & (!g36) & (!reset) & (g675) & (!g1730)) + ((g34) & (!g36) & (!reset) & (g675) & (g1730)) + ((g34) & (g36) & (!reset) & (g675) & (!g1730)) + ((g34) & (g36) & (!reset) & (g675) & (g1730)));
	assign g7708 = (((!g832) & (g3201) & (!g1732)) + ((!g832) & (g3201) & (g1732)) + ((g832) & (!g3201) & (g1732)) + ((g832) & (g3201) & (g1732)));
	assign g1733 = (((!g34) & (!g36) & (!reset) & (g676) & (!g1732)) + ((!g34) & (!g36) & (!reset) & (g676) & (g1732)) + ((!g34) & (g36) & (!reset) & (!g676) & (g1732)) + ((!g34) & (g36) & (!reset) & (g676) & (g1732)) + ((g34) & (!g36) & (!reset) & (g676) & (!g1732)) + ((g34) & (!g36) & (!reset) & (g676) & (g1732)) + ((g34) & (g36) & (!reset) & (g676) & (!g1732)) + ((g34) & (g36) & (!reset) & (g676) & (g1732)));
	assign g7709 = (((!g832) & (g3204) & (!g1734)) + ((!g832) & (g3204) & (g1734)) + ((g832) & (!g3204) & (g1734)) + ((g832) & (g3204) & (g1734)));
	assign g1735 = (((!g34) & (!g36) & (!reset) & (g677) & (!g1734)) + ((!g34) & (!g36) & (!reset) & (g677) & (g1734)) + ((!g34) & (g36) & (!reset) & (!g677) & (g1734)) + ((!g34) & (g36) & (!reset) & (g677) & (g1734)) + ((g34) & (!g36) & (!reset) & (g677) & (!g1734)) + ((g34) & (!g36) & (!reset) & (g677) & (g1734)) + ((g34) & (g36) & (!reset) & (g677) & (!g1734)) + ((g34) & (g36) & (!reset) & (g677) & (g1734)));
	assign g7710 = (((!g832) & (g3206) & (!g1736)) + ((!g832) & (g3206) & (g1736)) + ((g832) & (!g3206) & (g1736)) + ((g832) & (g3206) & (g1736)));
	assign g1737 = (((!g34) & (!g36) & (!reset) & (g679) & (!g1736)) + ((!g34) & (!g36) & (!reset) & (g679) & (g1736)) + ((!g34) & (g36) & (!reset) & (!g679) & (g1736)) + ((!g34) & (g36) & (!reset) & (g679) & (g1736)) + ((g34) & (!g36) & (!reset) & (g679) & (!g1736)) + ((g34) & (!g36) & (!reset) & (g679) & (g1736)) + ((g34) & (g36) & (!reset) & (g679) & (!g1736)) + ((g34) & (g36) & (!reset) & (g679) & (g1736)));
	assign g7711 = (((!g832) & (g3209) & (!g1738)) + ((!g832) & (g3209) & (g1738)) + ((g832) & (!g3209) & (g1738)) + ((g832) & (g3209) & (g1738)));
	assign g1739 = (((!g34) & (!g36) & (!reset) & (g680) & (!g1738)) + ((!g34) & (!g36) & (!reset) & (g680) & (g1738)) + ((!g34) & (g36) & (!reset) & (!g680) & (g1738)) + ((!g34) & (g36) & (!reset) & (g680) & (g1738)) + ((g34) & (!g36) & (!reset) & (g680) & (!g1738)) + ((g34) & (!g36) & (!reset) & (g680) & (g1738)) + ((g34) & (g36) & (!reset) & (g680) & (!g1738)) + ((g34) & (g36) & (!reset) & (g680) & (g1738)));
	assign g7712 = (((!g832) & (g3212) & (!g1740)) + ((!g832) & (g3212) & (g1740)) + ((g832) & (!g3212) & (g1740)) + ((g832) & (g3212) & (g1740)));
	assign g1741 = (((!g34) & (!g36) & (!reset) & (g681) & (!g1740)) + ((!g34) & (!g36) & (!reset) & (g681) & (g1740)) + ((!g34) & (g36) & (!reset) & (!g681) & (g1740)) + ((!g34) & (g36) & (!reset) & (g681) & (g1740)) + ((g34) & (!g36) & (!reset) & (g681) & (!g1740)) + ((g34) & (!g36) & (!reset) & (g681) & (g1740)) + ((g34) & (g36) & (!reset) & (g681) & (!g1740)) + ((g34) & (g36) & (!reset) & (g681) & (g1740)));
	assign g7713 = (((!g832) & (g3215) & (!g1742)) + ((!g832) & (g3215) & (g1742)) + ((g832) & (!g3215) & (g1742)) + ((g832) & (g3215) & (g1742)));
	assign g1743 = (((!g34) & (!g36) & (!reset) & (g682) & (!g1742)) + ((!g34) & (!g36) & (!reset) & (g682) & (g1742)) + ((!g34) & (g36) & (!reset) & (!g682) & (g1742)) + ((!g34) & (g36) & (!reset) & (g682) & (g1742)) + ((g34) & (!g36) & (!reset) & (g682) & (!g1742)) + ((g34) & (!g36) & (!reset) & (g682) & (g1742)) + ((g34) & (g36) & (!reset) & (g682) & (!g1742)) + ((g34) & (g36) & (!reset) & (g682) & (g1742)));
	assign g7714 = (((!g2017) & (g7095) & (!g1744)) + ((!g2017) & (g7095) & (g1744)) + ((g2017) & (!g7095) & (g1744)) + ((g2017) & (g7095) & (g1744)));
	assign g1745 = (((!g639) & (!g662) & (g1677) & (g1711) & (g1678)) + ((!g639) & (g662) & (!g1677) & (g1711) & (!g1678)) + ((!g639) & (g662) & (!g1677) & (g1711) & (g1678)) + ((!g639) & (g662) & (g1677) & (!g1711) & (g1678)) + ((!g639) & (g662) & (g1677) & (g1711) & (!g1678)) + ((!g639) & (g662) & (g1677) & (g1711) & (g1678)) + ((g639) & (!g662) & (!g1677) & (g1711) & (g1678)) + ((g639) & (!g662) & (g1677) & (g1711) & (!g1678)) + ((g639) & (!g662) & (g1677) & (g1711) & (g1678)) + ((g639) & (g662) & (!g1677) & (!g1711) & (g1678)) + ((g639) & (g662) & (!g1677) & (g1711) & (!g1678)) + ((g639) & (g662) & (!g1677) & (g1711) & (g1678)) + ((g639) & (g662) & (g1677) & (!g1711) & (!g1678)) + ((g639) & (g662) & (g1677) & (!g1711) & (g1678)) + ((g639) & (g662) & (g1677) & (g1711) & (!g1678)) + ((g639) & (g662) & (g1677) & (g1711) & (g1678)));
	assign g1746 = (((!g827) & (!g685) & (g1744) & (!g1745)) + ((!g827) & (!g685) & (g1744) & (g1745)) + ((!g827) & (g685) & (g1744) & (!g1745)) + ((!g827) & (g685) & (g1744) & (g1745)) + ((g827) & (!g685) & (!g1744) & (g1745)) + ((g827) & (!g685) & (g1744) & (!g1745)) + ((g827) & (g685) & (!g1744) & (!g1745)) + ((g827) & (g685) & (g1744) & (g1745)));
	assign g1747 = (((!g34) & (!g36) & (!reset) & (g687) & (!g708)) + ((!g34) & (!g36) & (!reset) & (g687) & (g708)) + ((!g34) & (g36) & (!reset) & (!g687) & (g708)) + ((!g34) & (g36) & (!reset) & (g687) & (g708)) + ((g34) & (!g36) & (!reset) & (g687) & (!g708)) + ((g34) & (!g36) & (!reset) & (g687) & (g708)) + ((g34) & (g36) & (!reset) & (g687) & (!g708)) + ((g34) & (g36) & (!reset) & (g687) & (g708)));
	assign g7715 = (((!g832) & (g3221) & (!g1748)) + ((!g832) & (g3221) & (g1748)) + ((g832) & (!g3221) & (g1748)) + ((g832) & (g3221) & (g1748)));
	assign g1749 = (((!g34) & (!g36) & (!reset) & (g688) & (!g1748)) + ((!g34) & (!g36) & (!reset) & (g688) & (g1748)) + ((!g34) & (g36) & (!reset) & (!g688) & (g1748)) + ((!g34) & (g36) & (!reset) & (g688) & (g1748)) + ((g34) & (!g36) & (!reset) & (g688) & (!g1748)) + ((g34) & (!g36) & (!reset) & (g688) & (g1748)) + ((g34) & (g36) & (!reset) & (g688) & (!g1748)) + ((g34) & (g36) & (!reset) & (g688) & (g1748)));
	assign g7716 = (((!g832) & (g3226) & (!g1750)) + ((!g832) & (g3226) & (g1750)) + ((g832) & (!g3226) & (g1750)) + ((g832) & (g3226) & (g1750)));
	assign g1751 = (((!g34) & (!g36) & (!reset) & (g689) & (!g1750)) + ((!g34) & (!g36) & (!reset) & (g689) & (g1750)) + ((!g34) & (g36) & (!reset) & (!g689) & (g1750)) + ((!g34) & (g36) & (!reset) & (g689) & (g1750)) + ((g34) & (!g36) & (!reset) & (g689) & (!g1750)) + ((g34) & (!g36) & (!reset) & (g689) & (g1750)) + ((g34) & (g36) & (!reset) & (g689) & (!g1750)) + ((g34) & (g36) & (!reset) & (g689) & (g1750)));
	assign g7717 = (((!g832) & (g3230) & (!g1752)) + ((!g832) & (g3230) & (g1752)) + ((g832) & (!g3230) & (g1752)) + ((g832) & (g3230) & (g1752)));
	assign g1753 = (((!g34) & (!g36) & (!reset) & (g690) & (!g1752)) + ((!g34) & (!g36) & (!reset) & (g690) & (g1752)) + ((!g34) & (g36) & (!reset) & (!g690) & (g1752)) + ((!g34) & (g36) & (!reset) & (g690) & (g1752)) + ((g34) & (!g36) & (!reset) & (g690) & (!g1752)) + ((g34) & (!g36) & (!reset) & (g690) & (g1752)) + ((g34) & (g36) & (!reset) & (g690) & (!g1752)) + ((g34) & (g36) & (!reset) & (g690) & (g1752)));
	assign g7718 = (((!g832) & (g3234) & (!g1754)) + ((!g832) & (g3234) & (g1754)) + ((g832) & (!g3234) & (g1754)) + ((g832) & (g3234) & (g1754)));
	assign g1755 = (((!g34) & (!g36) & (!reset) & (g692) & (!g1754)) + ((!g34) & (!g36) & (!reset) & (g692) & (g1754)) + ((!g34) & (g36) & (!reset) & (!g692) & (g1754)) + ((!g34) & (g36) & (!reset) & (g692) & (g1754)) + ((g34) & (!g36) & (!reset) & (g692) & (!g1754)) + ((g34) & (!g36) & (!reset) & (g692) & (g1754)) + ((g34) & (g36) & (!reset) & (g692) & (!g1754)) + ((g34) & (g36) & (!reset) & (g692) & (g1754)));
	assign g7719 = (((!g832) & (g3239) & (!g1756)) + ((!g832) & (g3239) & (g1756)) + ((g832) & (!g3239) & (g1756)) + ((g832) & (g3239) & (g1756)));
	assign g1757 = (((!g34) & (!g36) & (!reset) & (g693) & (!g1756)) + ((!g34) & (!g36) & (!reset) & (g693) & (g1756)) + ((!g34) & (g36) & (!reset) & (!g693) & (g1756)) + ((!g34) & (g36) & (!reset) & (g693) & (g1756)) + ((g34) & (!g36) & (!reset) & (g693) & (!g1756)) + ((g34) & (!g36) & (!reset) & (g693) & (g1756)) + ((g34) & (g36) & (!reset) & (g693) & (!g1756)) + ((g34) & (g36) & (!reset) & (g693) & (g1756)));
	assign g7720 = (((!g832) & (g3244) & (!g1758)) + ((!g832) & (g3244) & (g1758)) + ((g832) & (!g3244) & (g1758)) + ((g832) & (g3244) & (g1758)));
	assign g1759 = (((!g34) & (!g36) & (!reset) & (g694) & (!g1758)) + ((!g34) & (!g36) & (!reset) & (g694) & (g1758)) + ((!g34) & (g36) & (!reset) & (!g694) & (g1758)) + ((!g34) & (g36) & (!reset) & (g694) & (g1758)) + ((g34) & (!g36) & (!reset) & (g694) & (!g1758)) + ((g34) & (!g36) & (!reset) & (g694) & (g1758)) + ((g34) & (g36) & (!reset) & (g694) & (!g1758)) + ((g34) & (g36) & (!reset) & (g694) & (g1758)));
	assign g7721 = (((!g832) & (g3249) & (!g1760)) + ((!g832) & (g3249) & (g1760)) + ((g832) & (!g3249) & (g1760)) + ((g832) & (g3249) & (g1760)));
	assign g1761 = (((!g34) & (!g36) & (!reset) & (g695) & (!g1760)) + ((!g34) & (!g36) & (!reset) & (g695) & (g1760)) + ((!g34) & (g36) & (!reset) & (!g695) & (g1760)) + ((!g34) & (g36) & (!reset) & (g695) & (g1760)) + ((g34) & (!g36) & (!reset) & (g695) & (!g1760)) + ((g34) & (!g36) & (!reset) & (g695) & (g1760)) + ((g34) & (g36) & (!reset) & (g695) & (!g1760)) + ((g34) & (g36) & (!reset) & (g695) & (g1760)));
	assign g7722 = (((!g832) & (g3254) & (!g1762)) + ((!g832) & (g3254) & (g1762)) + ((g832) & (!g3254) & (g1762)) + ((g832) & (g3254) & (g1762)));
	assign g1763 = (((!g34) & (!g36) & (!reset) & (g697) & (!g1762)) + ((!g34) & (!g36) & (!reset) & (g697) & (g1762)) + ((!g34) & (g36) & (!reset) & (!g697) & (g1762)) + ((!g34) & (g36) & (!reset) & (g697) & (g1762)) + ((g34) & (!g36) & (!reset) & (g697) & (!g1762)) + ((g34) & (!g36) & (!reset) & (g697) & (g1762)) + ((g34) & (g36) & (!reset) & (g697) & (!g1762)) + ((g34) & (g36) & (!reset) & (g697) & (g1762)));
	assign g7723 = (((!g832) & (g3259) & (!g1764)) + ((!g832) & (g3259) & (g1764)) + ((g832) & (!g3259) & (g1764)) + ((g832) & (g3259) & (g1764)));
	assign g1765 = (((!g34) & (!g36) & (!reset) & (g698) & (!g1764)) + ((!g34) & (!g36) & (!reset) & (g698) & (g1764)) + ((!g34) & (g36) & (!reset) & (!g698) & (g1764)) + ((!g34) & (g36) & (!reset) & (g698) & (g1764)) + ((g34) & (!g36) & (!reset) & (g698) & (!g1764)) + ((g34) & (!g36) & (!reset) & (g698) & (g1764)) + ((g34) & (g36) & (!reset) & (g698) & (!g1764)) + ((g34) & (g36) & (!reset) & (g698) & (g1764)));
	assign g7724 = (((!g832) & (g3264) & (!g1766)) + ((!g832) & (g3264) & (g1766)) + ((g832) & (!g3264) & (g1766)) + ((g832) & (g3264) & (g1766)));
	assign g1767 = (((!g34) & (!g36) & (!reset) & (g699) & (!g1766)) + ((!g34) & (!g36) & (!reset) & (g699) & (g1766)) + ((!g34) & (g36) & (!reset) & (!g699) & (g1766)) + ((!g34) & (g36) & (!reset) & (g699) & (g1766)) + ((g34) & (!g36) & (!reset) & (g699) & (!g1766)) + ((g34) & (!g36) & (!reset) & (g699) & (g1766)) + ((g34) & (g36) & (!reset) & (g699) & (!g1766)) + ((g34) & (g36) & (!reset) & (g699) & (g1766)));
	assign g7725 = (((!g832) & (g3269) & (!g1768)) + ((!g832) & (g3269) & (g1768)) + ((g832) & (!g3269) & (g1768)) + ((g832) & (g3269) & (g1768)));
	assign g1769 = (((!g34) & (!g36) & (!reset) & (g700) & (!g1768)) + ((!g34) & (!g36) & (!reset) & (g700) & (g1768)) + ((!g34) & (g36) & (!reset) & (!g700) & (g1768)) + ((!g34) & (g36) & (!reset) & (g700) & (g1768)) + ((g34) & (!g36) & (!reset) & (g700) & (!g1768)) + ((g34) & (!g36) & (!reset) & (g700) & (g1768)) + ((g34) & (g36) & (!reset) & (g700) & (!g1768)) + ((g34) & (g36) & (!reset) & (g700) & (g1768)));
	assign g7726 = (((!g832) & (g3273) & (!g1770)) + ((!g832) & (g3273) & (g1770)) + ((g832) & (!g3273) & (g1770)) + ((g832) & (g3273) & (g1770)));
	assign g1771 = (((!g34) & (!g36) & (!reset) & (g702) & (!g1770)) + ((!g34) & (!g36) & (!reset) & (g702) & (g1770)) + ((!g34) & (g36) & (!reset) & (!g702) & (g1770)) + ((!g34) & (g36) & (!reset) & (g702) & (g1770)) + ((g34) & (!g36) & (!reset) & (g702) & (!g1770)) + ((g34) & (!g36) & (!reset) & (g702) & (g1770)) + ((g34) & (g36) & (!reset) & (g702) & (!g1770)) + ((g34) & (g36) & (!reset) & (g702) & (g1770)));
	assign g7727 = (((!g832) & (g3278) & (!g1772)) + ((!g832) & (g3278) & (g1772)) + ((g832) & (!g3278) & (g1772)) + ((g832) & (g3278) & (g1772)));
	assign g1773 = (((!g34) & (!g36) & (!reset) & (g703) & (!g1772)) + ((!g34) & (!g36) & (!reset) & (g703) & (g1772)) + ((!g34) & (g36) & (!reset) & (!g703) & (g1772)) + ((!g34) & (g36) & (!reset) & (g703) & (g1772)) + ((g34) & (!g36) & (!reset) & (g703) & (!g1772)) + ((g34) & (!g36) & (!reset) & (g703) & (g1772)) + ((g34) & (g36) & (!reset) & (g703) & (!g1772)) + ((g34) & (g36) & (!reset) & (g703) & (g1772)));
	assign g7728 = (((!g832) & (g3283) & (!g1774)) + ((!g832) & (g3283) & (g1774)) + ((g832) & (!g3283) & (g1774)) + ((g832) & (g3283) & (g1774)));
	assign g1775 = (((!g34) & (!g36) & (!reset) & (g704) & (!g1774)) + ((!g34) & (!g36) & (!reset) & (g704) & (g1774)) + ((!g34) & (g36) & (!reset) & (!g704) & (g1774)) + ((!g34) & (g36) & (!reset) & (g704) & (g1774)) + ((g34) & (!g36) & (!reset) & (g704) & (!g1774)) + ((g34) & (!g36) & (!reset) & (g704) & (g1774)) + ((g34) & (g36) & (!reset) & (g704) & (!g1774)) + ((g34) & (g36) & (!reset) & (g704) & (g1774)));
	assign g7729 = (((!g832) & (g3288) & (!g1776)) + ((!g832) & (g3288) & (g1776)) + ((g832) & (!g3288) & (g1776)) + ((g832) & (g3288) & (g1776)));
	assign g1777 = (((!g34) & (!g36) & (!reset) & (g705) & (!g1776)) + ((!g34) & (!g36) & (!reset) & (g705) & (g1776)) + ((!g34) & (g36) & (!reset) & (!g705) & (g1776)) + ((!g34) & (g36) & (!reset) & (g705) & (g1776)) + ((g34) & (!g36) & (!reset) & (g705) & (!g1776)) + ((g34) & (!g36) & (!reset) & (g705) & (g1776)) + ((g34) & (g36) & (!reset) & (g705) & (!g1776)) + ((g34) & (g36) & (!reset) & (g705) & (g1776)));
	assign g7730 = (((!g2017) & (g7089) & (!g1778)) + ((!g2017) & (g7089) & (g1778)) + ((g2017) & (!g7089) & (g1778)) + ((g2017) & (g7089) & (g1778)));
	assign g1779 = (((!g685) & (g1744)) + ((g685) & (!g1744)));
	assign g1780 = (((!g639) & (!g662) & (g1677) & (g1711) & (g1678) & (g1779)) + ((!g639) & (g662) & (!g1677) & (g1711) & (!g1678) & (g1779)) + ((!g639) & (g662) & (!g1677) & (g1711) & (g1678) & (g1779)) + ((!g639) & (g662) & (g1677) & (!g1711) & (g1678) & (g1779)) + ((!g639) & (g662) & (g1677) & (g1711) & (!g1678) & (g1779)) + ((!g639) & (g662) & (g1677) & (g1711) & (g1678) & (g1779)) + ((g639) & (!g662) & (!g1677) & (g1711) & (g1678) & (g1779)) + ((g639) & (!g662) & (g1677) & (g1711) & (!g1678) & (g1779)) + ((g639) & (!g662) & (g1677) & (g1711) & (g1678) & (g1779)) + ((g639) & (g662) & (!g1677) & (!g1711) & (g1678) & (g1779)) + ((g639) & (g662) & (!g1677) & (g1711) & (!g1678) & (g1779)) + ((g639) & (g662) & (!g1677) & (g1711) & (g1678) & (g1779)) + ((g639) & (g662) & (g1677) & (!g1711) & (!g1678) & (g1779)) + ((g639) & (g662) & (g1677) & (!g1711) & (g1678) & (g1779)) + ((g639) & (g662) & (g1677) & (g1711) & (!g1678) & (g1779)) + ((g639) & (g662) & (g1677) & (g1711) & (g1678) & (g1779)));
	assign g1781 = (((g685) & (g1744)));
	assign g1782 = (((!g827) & (!g708) & (g1778) & (!g1780) & (!g1781)) + ((!g827) & (!g708) & (g1778) & (!g1780) & (g1781)) + ((!g827) & (!g708) & (g1778) & (g1780) & (!g1781)) + ((!g827) & (!g708) & (g1778) & (g1780) & (g1781)) + ((!g827) & (g708) & (g1778) & (!g1780) & (!g1781)) + ((!g827) & (g708) & (g1778) & (!g1780) & (g1781)) + ((!g827) & (g708) & (g1778) & (g1780) & (!g1781)) + ((!g827) & (g708) & (g1778) & (g1780) & (g1781)) + ((g827) & (!g708) & (!g1778) & (!g1780) & (g1781)) + ((g827) & (!g708) & (!g1778) & (g1780) & (!g1781)) + ((g827) & (!g708) & (!g1778) & (g1780) & (g1781)) + ((g827) & (!g708) & (g1778) & (!g1780) & (!g1781)) + ((g827) & (g708) & (!g1778) & (!g1780) & (!g1781)) + ((g827) & (g708) & (g1778) & (!g1780) & (g1781)) + ((g827) & (g708) & (g1778) & (g1780) & (!g1781)) + ((g827) & (g708) & (g1778) & (g1780) & (g1781)));
	assign g1783 = (((!g34) & (!g36) & (!reset) & (g710) & (!g731)) + ((!g34) & (!g36) & (!reset) & (g710) & (g731)) + ((!g34) & (g36) & (!reset) & (!g710) & (g731)) + ((!g34) & (g36) & (!reset) & (g710) & (g731)) + ((g34) & (!g36) & (!reset) & (g710) & (!g731)) + ((g34) & (!g36) & (!reset) & (g710) & (g731)) + ((g34) & (g36) & (!reset) & (g710) & (!g731)) + ((g34) & (g36) & (!reset) & (g710) & (g731)));
	assign g7731 = (((!g832) & (g3290) & (!g1784)) + ((!g832) & (g3290) & (g1784)) + ((g832) & (!g3290) & (g1784)) + ((g832) & (g3290) & (g1784)));
	assign g1785 = (((!g34) & (!g36) & (!reset) & (g711) & (!g1784)) + ((!g34) & (!g36) & (!reset) & (g711) & (g1784)) + ((!g34) & (g36) & (!reset) & (!g711) & (g1784)) + ((!g34) & (g36) & (!reset) & (g711) & (g1784)) + ((g34) & (!g36) & (!reset) & (g711) & (!g1784)) + ((g34) & (!g36) & (!reset) & (g711) & (g1784)) + ((g34) & (g36) & (!reset) & (g711) & (!g1784)) + ((g34) & (g36) & (!reset) & (g711) & (g1784)));
	assign g7732 = (((!g832) & (g3292) & (!g1786)) + ((!g832) & (g3292) & (g1786)) + ((g832) & (!g3292) & (g1786)) + ((g832) & (g3292) & (g1786)));
	assign g1787 = (((!g34) & (!g36) & (!reset) & (g712) & (!g1786)) + ((!g34) & (!g36) & (!reset) & (g712) & (g1786)) + ((!g34) & (g36) & (!reset) & (!g712) & (g1786)) + ((!g34) & (g36) & (!reset) & (g712) & (g1786)) + ((g34) & (!g36) & (!reset) & (g712) & (!g1786)) + ((g34) & (!g36) & (!reset) & (g712) & (g1786)) + ((g34) & (g36) & (!reset) & (g712) & (!g1786)) + ((g34) & (g36) & (!reset) & (g712) & (g1786)));
	assign g7733 = (((!g832) & (g3293) & (!g1788)) + ((!g832) & (g3293) & (g1788)) + ((g832) & (!g3293) & (g1788)) + ((g832) & (g3293) & (g1788)));
	assign g1789 = (((!g34) & (!g36) & (!reset) & (g713) & (!g1788)) + ((!g34) & (!g36) & (!reset) & (g713) & (g1788)) + ((!g34) & (g36) & (!reset) & (!g713) & (g1788)) + ((!g34) & (g36) & (!reset) & (g713) & (g1788)) + ((g34) & (!g36) & (!reset) & (g713) & (!g1788)) + ((g34) & (!g36) & (!reset) & (g713) & (g1788)) + ((g34) & (g36) & (!reset) & (g713) & (!g1788)) + ((g34) & (g36) & (!reset) & (g713) & (g1788)));
	assign g7734 = (((!g832) & (g3294) & (!g1790)) + ((!g832) & (g3294) & (g1790)) + ((g832) & (!g3294) & (g1790)) + ((g832) & (g3294) & (g1790)));
	assign g1791 = (((!g34) & (!g36) & (!reset) & (g715) & (!g1790)) + ((!g34) & (!g36) & (!reset) & (g715) & (g1790)) + ((!g34) & (g36) & (!reset) & (!g715) & (g1790)) + ((!g34) & (g36) & (!reset) & (g715) & (g1790)) + ((g34) & (!g36) & (!reset) & (g715) & (!g1790)) + ((g34) & (!g36) & (!reset) & (g715) & (g1790)) + ((g34) & (g36) & (!reset) & (g715) & (!g1790)) + ((g34) & (g36) & (!reset) & (g715) & (g1790)));
	assign g7735 = (((!g832) & (g3296) & (!g1792)) + ((!g832) & (g3296) & (g1792)) + ((g832) & (!g3296) & (g1792)) + ((g832) & (g3296) & (g1792)));
	assign g1793 = (((!g34) & (!g36) & (!reset) & (g716) & (!g1792)) + ((!g34) & (!g36) & (!reset) & (g716) & (g1792)) + ((!g34) & (g36) & (!reset) & (!g716) & (g1792)) + ((!g34) & (g36) & (!reset) & (g716) & (g1792)) + ((g34) & (!g36) & (!reset) & (g716) & (!g1792)) + ((g34) & (!g36) & (!reset) & (g716) & (g1792)) + ((g34) & (g36) & (!reset) & (g716) & (!g1792)) + ((g34) & (g36) & (!reset) & (g716) & (g1792)));
	assign g7736 = (((!g832) & (g3298) & (!g1794)) + ((!g832) & (g3298) & (g1794)) + ((g832) & (!g3298) & (g1794)) + ((g832) & (g3298) & (g1794)));
	assign g1795 = (((!g34) & (!g36) & (!reset) & (g717) & (!g1794)) + ((!g34) & (!g36) & (!reset) & (g717) & (g1794)) + ((!g34) & (g36) & (!reset) & (!g717) & (g1794)) + ((!g34) & (g36) & (!reset) & (g717) & (g1794)) + ((g34) & (!g36) & (!reset) & (g717) & (!g1794)) + ((g34) & (!g36) & (!reset) & (g717) & (g1794)) + ((g34) & (g36) & (!reset) & (g717) & (!g1794)) + ((g34) & (g36) & (!reset) & (g717) & (g1794)));
	assign g7737 = (((!g832) & (g3300) & (!g1796)) + ((!g832) & (g3300) & (g1796)) + ((g832) & (!g3300) & (g1796)) + ((g832) & (g3300) & (g1796)));
	assign g1797 = (((!g34) & (!g36) & (!reset) & (g718) & (!g1796)) + ((!g34) & (!g36) & (!reset) & (g718) & (g1796)) + ((!g34) & (g36) & (!reset) & (!g718) & (g1796)) + ((!g34) & (g36) & (!reset) & (g718) & (g1796)) + ((g34) & (!g36) & (!reset) & (g718) & (!g1796)) + ((g34) & (!g36) & (!reset) & (g718) & (g1796)) + ((g34) & (g36) & (!reset) & (g718) & (!g1796)) + ((g34) & (g36) & (!reset) & (g718) & (g1796)));
	assign g7738 = (((!g832) & (g3302) & (!g1798)) + ((!g832) & (g3302) & (g1798)) + ((g832) & (!g3302) & (g1798)) + ((g832) & (g3302) & (g1798)));
	assign g1799 = (((!g34) & (!g36) & (!reset) & (g720) & (!g1798)) + ((!g34) & (!g36) & (!reset) & (g720) & (g1798)) + ((!g34) & (g36) & (!reset) & (!g720) & (g1798)) + ((!g34) & (g36) & (!reset) & (g720) & (g1798)) + ((g34) & (!g36) & (!reset) & (g720) & (!g1798)) + ((g34) & (!g36) & (!reset) & (g720) & (g1798)) + ((g34) & (g36) & (!reset) & (g720) & (!g1798)) + ((g34) & (g36) & (!reset) & (g720) & (g1798)));
	assign g7739 = (((!g832) & (g3304) & (!g1800)) + ((!g832) & (g3304) & (g1800)) + ((g832) & (!g3304) & (g1800)) + ((g832) & (g3304) & (g1800)));
	assign g1801 = (((!g34) & (!g36) & (!reset) & (g721) & (!g1800)) + ((!g34) & (!g36) & (!reset) & (g721) & (g1800)) + ((!g34) & (g36) & (!reset) & (!g721) & (g1800)) + ((!g34) & (g36) & (!reset) & (g721) & (g1800)) + ((g34) & (!g36) & (!reset) & (g721) & (!g1800)) + ((g34) & (!g36) & (!reset) & (g721) & (g1800)) + ((g34) & (g36) & (!reset) & (g721) & (!g1800)) + ((g34) & (g36) & (!reset) & (g721) & (g1800)));
	assign g7740 = (((!g832) & (g3306) & (!g1802)) + ((!g832) & (g3306) & (g1802)) + ((g832) & (!g3306) & (g1802)) + ((g832) & (g3306) & (g1802)));
	assign g1803 = (((!g34) & (!g36) & (!reset) & (g722) & (!g1802)) + ((!g34) & (!g36) & (!reset) & (g722) & (g1802)) + ((!g34) & (g36) & (!reset) & (!g722) & (g1802)) + ((!g34) & (g36) & (!reset) & (g722) & (g1802)) + ((g34) & (!g36) & (!reset) & (g722) & (!g1802)) + ((g34) & (!g36) & (!reset) & (g722) & (g1802)) + ((g34) & (g36) & (!reset) & (g722) & (!g1802)) + ((g34) & (g36) & (!reset) & (g722) & (g1802)));
	assign g7741 = (((!g832) & (g3308) & (!g1804)) + ((!g832) & (g3308) & (g1804)) + ((g832) & (!g3308) & (g1804)) + ((g832) & (g3308) & (g1804)));
	assign g1805 = (((!g34) & (!g36) & (!reset) & (g723) & (!g1804)) + ((!g34) & (!g36) & (!reset) & (g723) & (g1804)) + ((!g34) & (g36) & (!reset) & (!g723) & (g1804)) + ((!g34) & (g36) & (!reset) & (g723) & (g1804)) + ((g34) & (!g36) & (!reset) & (g723) & (!g1804)) + ((g34) & (!g36) & (!reset) & (g723) & (g1804)) + ((g34) & (g36) & (!reset) & (g723) & (!g1804)) + ((g34) & (g36) & (!reset) & (g723) & (g1804)));
	assign g7742 = (((!g832) & (g3309) & (!g1806)) + ((!g832) & (g3309) & (g1806)) + ((g832) & (!g3309) & (g1806)) + ((g832) & (g3309) & (g1806)));
	assign g1807 = (((!g34) & (!g36) & (!reset) & (g725) & (!g1806)) + ((!g34) & (!g36) & (!reset) & (g725) & (g1806)) + ((!g34) & (g36) & (!reset) & (!g725) & (g1806)) + ((!g34) & (g36) & (!reset) & (g725) & (g1806)) + ((g34) & (!g36) & (!reset) & (g725) & (!g1806)) + ((g34) & (!g36) & (!reset) & (g725) & (g1806)) + ((g34) & (g36) & (!reset) & (g725) & (!g1806)) + ((g34) & (g36) & (!reset) & (g725) & (g1806)));
	assign g7743 = (((!g832) & (g3311) & (!g1808)) + ((!g832) & (g3311) & (g1808)) + ((g832) & (!g3311) & (g1808)) + ((g832) & (g3311) & (g1808)));
	assign g1809 = (((!g34) & (!g36) & (!reset) & (g726) & (!g1808)) + ((!g34) & (!g36) & (!reset) & (g726) & (g1808)) + ((!g34) & (g36) & (!reset) & (!g726) & (g1808)) + ((!g34) & (g36) & (!reset) & (g726) & (g1808)) + ((g34) & (!g36) & (!reset) & (g726) & (!g1808)) + ((g34) & (!g36) & (!reset) & (g726) & (g1808)) + ((g34) & (g36) & (!reset) & (g726) & (!g1808)) + ((g34) & (g36) & (!reset) & (g726) & (g1808)));
	assign g7744 = (((!g832) & (g3313) & (!g1810)) + ((!g832) & (g3313) & (g1810)) + ((g832) & (!g3313) & (g1810)) + ((g832) & (g3313) & (g1810)));
	assign g1811 = (((!g34) & (!g36) & (!reset) & (g727) & (!g1810)) + ((!g34) & (!g36) & (!reset) & (g727) & (g1810)) + ((!g34) & (g36) & (!reset) & (!g727) & (g1810)) + ((!g34) & (g36) & (!reset) & (g727) & (g1810)) + ((g34) & (!g36) & (!reset) & (g727) & (!g1810)) + ((g34) & (!g36) & (!reset) & (g727) & (g1810)) + ((g34) & (g36) & (!reset) & (g727) & (!g1810)) + ((g34) & (g36) & (!reset) & (g727) & (g1810)));
	assign g7745 = (((!g832) & (g3315) & (!g1812)) + ((!g832) & (g3315) & (g1812)) + ((g832) & (!g3315) & (g1812)) + ((g832) & (g3315) & (g1812)));
	assign g1813 = (((!g34) & (!g36) & (!reset) & (g728) & (!g1812)) + ((!g34) & (!g36) & (!reset) & (g728) & (g1812)) + ((!g34) & (g36) & (!reset) & (!g728) & (g1812)) + ((!g34) & (g36) & (!reset) & (g728) & (g1812)) + ((g34) & (!g36) & (!reset) & (g728) & (!g1812)) + ((g34) & (!g36) & (!reset) & (g728) & (g1812)) + ((g34) & (g36) & (!reset) & (g728) & (!g1812)) + ((g34) & (g36) & (!reset) & (g728) & (g1812)));
	assign g7746 = (((!g2017) & (g3320) & (!g1814)) + ((!g2017) & (g3320) & (g1814)) + ((g2017) & (!g3320) & (g1814)) + ((g2017) & (g3320) & (g1814)));
	assign g1815 = (((!g827) & (!g708) & (!g1778) & (!g1780) & (!g1781) & (g5648)) + ((!g827) & (!g708) & (!g1778) & (!g1780) & (g1781) & (g5648)) + ((!g827) & (!g708) & (!g1778) & (g1780) & (!g1781) & (g5648)) + ((!g827) & (!g708) & (!g1778) & (g1780) & (g1781) & (g5648)) + ((!g827) & (!g708) & (g1778) & (!g1780) & (!g1781) & (g5648)) + ((!g827) & (!g708) & (g1778) & (!g1780) & (g1781) & (g5648)) + ((!g827) & (!g708) & (g1778) & (g1780) & (!g1781) & (g5648)) + ((!g827) & (!g708) & (g1778) & (g1780) & (g1781) & (g5648)) + ((!g827) & (g708) & (!g1778) & (!g1780) & (!g1781) & (g5648)) + ((!g827) & (g708) & (!g1778) & (!g1780) & (g1781) & (g5648)) + ((!g827) & (g708) & (!g1778) & (g1780) & (!g1781) & (g5648)) + ((!g827) & (g708) & (!g1778) & (g1780) & (g1781) & (g5648)) + ((!g827) & (g708) & (g1778) & (!g1780) & (!g1781) & (g5648)) + ((!g827) & (g708) & (g1778) & (!g1780) & (g1781) & (g5648)) + ((!g827) & (g708) & (g1778) & (g1780) & (!g1781) & (g5648)) + ((!g827) & (g708) & (g1778) & (g1780) & (g1781) & (g5648)) + ((g827) & (!g708) & (!g1778) & (!g1780) & (!g1781) & (!g5648)) + ((g827) & (!g708) & (!g1778) & (!g1780) & (g1781) & (!g5648)) + ((g827) & (!g708) & (!g1778) & (g1780) & (!g1781) & (!g5648)) + ((g827) & (!g708) & (!g1778) & (g1780) & (g1781) & (!g5648)) + ((g827) & (!g708) & (g1778) & (!g1780) & (!g1781) & (!g5648)) + ((g827) & (!g708) & (g1778) & (!g1780) & (g1781) & (g5648)) + ((g827) & (!g708) & (g1778) & (g1780) & (!g1781) & (g5648)) + ((g827) & (!g708) & (g1778) & (g1780) & (g1781) & (g5648)) + ((g827) & (g708) & (!g1778) & (!g1780) & (!g1781) & (!g5648)) + ((g827) & (g708) & (!g1778) & (!g1780) & (g1781) & (g5648)) + ((g827) & (g708) & (!g1778) & (g1780) & (!g1781) & (g5648)) + ((g827) & (g708) & (!g1778) & (g1780) & (g1781) & (g5648)) + ((g827) & (g708) & (g1778) & (!g1780) & (!g1781) & (g5648)) + ((g827) & (g708) & (g1778) & (!g1780) & (g1781) & (g5648)) + ((g827) & (g708) & (g1778) & (g1780) & (!g1781) & (g5648)) + ((g827) & (g708) & (g1778) & (g1780) & (g1781) & (g5648)));
	assign g1816 = (((!g34) & (!g36) & (!reset) & (g733) & (!g754)) + ((!g34) & (!g36) & (!reset) & (g733) & (g754)) + ((!g34) & (g36) & (!reset) & (!g733) & (g754)) + ((!g34) & (g36) & (!reset) & (g733) & (g754)) + ((g34) & (!g36) & (!reset) & (g733) & (!g754)) + ((g34) & (!g36) & (!reset) & (g733) & (g754)) + ((g34) & (g36) & (!reset) & (g733) & (!g754)) + ((g34) & (g36) & (!reset) & (g733) & (g754)));
	assign g7747 = (((!g832) & (g3322) & (!g1817)) + ((!g832) & (g3322) & (g1817)) + ((g832) & (!g3322) & (g1817)) + ((g832) & (g3322) & (g1817)));
	assign g1818 = (((!g34) & (!g36) & (!reset) & (g734) & (!g1817)) + ((!g34) & (!g36) & (!reset) & (g734) & (g1817)) + ((!g34) & (g36) & (!reset) & (!g734) & (g1817)) + ((!g34) & (g36) & (!reset) & (g734) & (g1817)) + ((g34) & (!g36) & (!reset) & (g734) & (!g1817)) + ((g34) & (!g36) & (!reset) & (g734) & (g1817)) + ((g34) & (g36) & (!reset) & (g734) & (!g1817)) + ((g34) & (g36) & (!reset) & (g734) & (g1817)));
	assign g7748 = (((!g832) & (g3325) & (!g1819)) + ((!g832) & (g3325) & (g1819)) + ((g832) & (!g3325) & (g1819)) + ((g832) & (g3325) & (g1819)));
	assign g1820 = (((!g34) & (!g36) & (!reset) & (g735) & (!g1819)) + ((!g34) & (!g36) & (!reset) & (g735) & (g1819)) + ((!g34) & (g36) & (!reset) & (!g735) & (g1819)) + ((!g34) & (g36) & (!reset) & (g735) & (g1819)) + ((g34) & (!g36) & (!reset) & (g735) & (!g1819)) + ((g34) & (!g36) & (!reset) & (g735) & (g1819)) + ((g34) & (g36) & (!reset) & (g735) & (!g1819)) + ((g34) & (g36) & (!reset) & (g735) & (g1819)));
	assign g7749 = (((!g832) & (g3327) & (!g1821)) + ((!g832) & (g3327) & (g1821)) + ((g832) & (!g3327) & (g1821)) + ((g832) & (g3327) & (g1821)));
	assign g1822 = (((!g34) & (!g36) & (!reset) & (g736) & (!g1821)) + ((!g34) & (!g36) & (!reset) & (g736) & (g1821)) + ((!g34) & (g36) & (!reset) & (!g736) & (g1821)) + ((!g34) & (g36) & (!reset) & (g736) & (g1821)) + ((g34) & (!g36) & (!reset) & (g736) & (!g1821)) + ((g34) & (!g36) & (!reset) & (g736) & (g1821)) + ((g34) & (g36) & (!reset) & (g736) & (!g1821)) + ((g34) & (g36) & (!reset) & (g736) & (g1821)));
	assign g7750 = (((!g832) & (g3329) & (!g1823)) + ((!g832) & (g3329) & (g1823)) + ((g832) & (!g3329) & (g1823)) + ((g832) & (g3329) & (g1823)));
	assign g1824 = (((!g34) & (!g36) & (!reset) & (g738) & (!g1823)) + ((!g34) & (!g36) & (!reset) & (g738) & (g1823)) + ((!g34) & (g36) & (!reset) & (!g738) & (g1823)) + ((!g34) & (g36) & (!reset) & (g738) & (g1823)) + ((g34) & (!g36) & (!reset) & (g738) & (!g1823)) + ((g34) & (!g36) & (!reset) & (g738) & (g1823)) + ((g34) & (g36) & (!reset) & (g738) & (!g1823)) + ((g34) & (g36) & (!reset) & (g738) & (g1823)));
	assign g7751 = (((!g832) & (g3332) & (!g1825)) + ((!g832) & (g3332) & (g1825)) + ((g832) & (!g3332) & (g1825)) + ((g832) & (g3332) & (g1825)));
	assign g1826 = (((!g34) & (!g36) & (!reset) & (g739) & (!g1825)) + ((!g34) & (!g36) & (!reset) & (g739) & (g1825)) + ((!g34) & (g36) & (!reset) & (!g739) & (g1825)) + ((!g34) & (g36) & (!reset) & (g739) & (g1825)) + ((g34) & (!g36) & (!reset) & (g739) & (!g1825)) + ((g34) & (!g36) & (!reset) & (g739) & (g1825)) + ((g34) & (g36) & (!reset) & (g739) & (!g1825)) + ((g34) & (g36) & (!reset) & (g739) & (g1825)));
	assign g7752 = (((!g832) & (g3335) & (!g1827)) + ((!g832) & (g3335) & (g1827)) + ((g832) & (!g3335) & (g1827)) + ((g832) & (g3335) & (g1827)));
	assign g1828 = (((!g34) & (!g36) & (!reset) & (g740) & (!g1827)) + ((!g34) & (!g36) & (!reset) & (g740) & (g1827)) + ((!g34) & (g36) & (!reset) & (!g740) & (g1827)) + ((!g34) & (g36) & (!reset) & (g740) & (g1827)) + ((g34) & (!g36) & (!reset) & (g740) & (!g1827)) + ((g34) & (!g36) & (!reset) & (g740) & (g1827)) + ((g34) & (g36) & (!reset) & (g740) & (!g1827)) + ((g34) & (g36) & (!reset) & (g740) & (g1827)));
	assign g7753 = (((!g832) & (g3338) & (!g1829)) + ((!g832) & (g3338) & (g1829)) + ((g832) & (!g3338) & (g1829)) + ((g832) & (g3338) & (g1829)));
	assign g1830 = (((!g34) & (!g36) & (!reset) & (g741) & (!g1829)) + ((!g34) & (!g36) & (!reset) & (g741) & (g1829)) + ((!g34) & (g36) & (!reset) & (!g741) & (g1829)) + ((!g34) & (g36) & (!reset) & (g741) & (g1829)) + ((g34) & (!g36) & (!reset) & (g741) & (!g1829)) + ((g34) & (!g36) & (!reset) & (g741) & (g1829)) + ((g34) & (g36) & (!reset) & (g741) & (!g1829)) + ((g34) & (g36) & (!reset) & (g741) & (g1829)));
	assign g7754 = (((!g832) & (g3341) & (!g1831)) + ((!g832) & (g3341) & (g1831)) + ((g832) & (!g3341) & (g1831)) + ((g832) & (g3341) & (g1831)));
	assign g1832 = (((!g34) & (!g36) & (!reset) & (g743) & (!g1831)) + ((!g34) & (!g36) & (!reset) & (g743) & (g1831)) + ((!g34) & (g36) & (!reset) & (!g743) & (g1831)) + ((!g34) & (g36) & (!reset) & (g743) & (g1831)) + ((g34) & (!g36) & (!reset) & (g743) & (!g1831)) + ((g34) & (!g36) & (!reset) & (g743) & (g1831)) + ((g34) & (g36) & (!reset) & (g743) & (!g1831)) + ((g34) & (g36) & (!reset) & (g743) & (g1831)));
	assign g7755 = (((!g832) & (g3344) & (!g1833)) + ((!g832) & (g3344) & (g1833)) + ((g832) & (!g3344) & (g1833)) + ((g832) & (g3344) & (g1833)));
	assign g1834 = (((!g34) & (!g36) & (!reset) & (g744) & (!g1833)) + ((!g34) & (!g36) & (!reset) & (g744) & (g1833)) + ((!g34) & (g36) & (!reset) & (!g744) & (g1833)) + ((!g34) & (g36) & (!reset) & (g744) & (g1833)) + ((g34) & (!g36) & (!reset) & (g744) & (!g1833)) + ((g34) & (!g36) & (!reset) & (g744) & (g1833)) + ((g34) & (g36) & (!reset) & (g744) & (!g1833)) + ((g34) & (g36) & (!reset) & (g744) & (g1833)));
	assign g7756 = (((!g832) & (g3347) & (!g1835)) + ((!g832) & (g3347) & (g1835)) + ((g832) & (!g3347) & (g1835)) + ((g832) & (g3347) & (g1835)));
	assign g1836 = (((!g34) & (!g36) & (!reset) & (g745) & (!g1835)) + ((!g34) & (!g36) & (!reset) & (g745) & (g1835)) + ((!g34) & (g36) & (!reset) & (!g745) & (g1835)) + ((!g34) & (g36) & (!reset) & (g745) & (g1835)) + ((g34) & (!g36) & (!reset) & (g745) & (!g1835)) + ((g34) & (!g36) & (!reset) & (g745) & (g1835)) + ((g34) & (g36) & (!reset) & (g745) & (!g1835)) + ((g34) & (g36) & (!reset) & (g745) & (g1835)));
	assign g7757 = (((!g832) & (g3350) & (!g1837)) + ((!g832) & (g3350) & (g1837)) + ((g832) & (!g3350) & (g1837)) + ((g832) & (g3350) & (g1837)));
	assign g1838 = (((!g34) & (!g36) & (!reset) & (g746) & (!g1837)) + ((!g34) & (!g36) & (!reset) & (g746) & (g1837)) + ((!g34) & (g36) & (!reset) & (!g746) & (g1837)) + ((!g34) & (g36) & (!reset) & (g746) & (g1837)) + ((g34) & (!g36) & (!reset) & (g746) & (!g1837)) + ((g34) & (!g36) & (!reset) & (g746) & (g1837)) + ((g34) & (g36) & (!reset) & (g746) & (!g1837)) + ((g34) & (g36) & (!reset) & (g746) & (g1837)));
	assign g7758 = (((!g832) & (g3352) & (!g1839)) + ((!g832) & (g3352) & (g1839)) + ((g832) & (!g3352) & (g1839)) + ((g832) & (g3352) & (g1839)));
	assign g1840 = (((!g34) & (!g36) & (!reset) & (g748) & (!g1839)) + ((!g34) & (!g36) & (!reset) & (g748) & (g1839)) + ((!g34) & (g36) & (!reset) & (!g748) & (g1839)) + ((!g34) & (g36) & (!reset) & (g748) & (g1839)) + ((g34) & (!g36) & (!reset) & (g748) & (!g1839)) + ((g34) & (!g36) & (!reset) & (g748) & (g1839)) + ((g34) & (g36) & (!reset) & (g748) & (!g1839)) + ((g34) & (g36) & (!reset) & (g748) & (g1839)));
	assign g7759 = (((!g832) & (g3355) & (!g1841)) + ((!g832) & (g3355) & (g1841)) + ((g832) & (!g3355) & (g1841)) + ((g832) & (g3355) & (g1841)));
	assign g1842 = (((!g34) & (!g36) & (!reset) & (g749) & (!g1841)) + ((!g34) & (!g36) & (!reset) & (g749) & (g1841)) + ((!g34) & (g36) & (!reset) & (!g749) & (g1841)) + ((!g34) & (g36) & (!reset) & (g749) & (g1841)) + ((g34) & (!g36) & (!reset) & (g749) & (!g1841)) + ((g34) & (!g36) & (!reset) & (g749) & (g1841)) + ((g34) & (g36) & (!reset) & (g749) & (!g1841)) + ((g34) & (g36) & (!reset) & (g749) & (g1841)));
	assign g7760 = (((!g832) & (g3358) & (!g1843)) + ((!g832) & (g3358) & (g1843)) + ((g832) & (!g3358) & (g1843)) + ((g832) & (g3358) & (g1843)));
	assign g1844 = (((!g34) & (!g36) & (!reset) & (g750) & (!g1843)) + ((!g34) & (!g36) & (!reset) & (g750) & (g1843)) + ((!g34) & (g36) & (!reset) & (!g750) & (g1843)) + ((!g34) & (g36) & (!reset) & (g750) & (g1843)) + ((g34) & (!g36) & (!reset) & (g750) & (!g1843)) + ((g34) & (!g36) & (!reset) & (g750) & (g1843)) + ((g34) & (g36) & (!reset) & (g750) & (!g1843)) + ((g34) & (g36) & (!reset) & (g750) & (g1843)));
	assign g7761 = (((!g832) & (g3361) & (!g1845)) + ((!g832) & (g3361) & (g1845)) + ((g832) & (!g3361) & (g1845)) + ((g832) & (g3361) & (g1845)));
	assign g1846 = (((!g34) & (!g36) & (!reset) & (g751) & (!g1845)) + ((!g34) & (!g36) & (!reset) & (g751) & (g1845)) + ((!g34) & (g36) & (!reset) & (!g751) & (g1845)) + ((!g34) & (g36) & (!reset) & (g751) & (g1845)) + ((g34) & (!g36) & (!reset) & (g751) & (!g1845)) + ((g34) & (!g36) & (!reset) & (g751) & (g1845)) + ((g34) & (g36) & (!reset) & (g751) & (!g1845)) + ((g34) & (g36) & (!reset) & (g751) & (g1845)));
	assign g7762 = (((!g2017) & (g3364) & (!g1847)) + ((!g2017) & (g3364) & (g1847)) + ((g2017) & (!g3364) & (g1847)) + ((g2017) & (g3364) & (g1847)));
	assign g1848 = (((!g708) & (!g731) & (!g1778) & (!g1814) & (!g1780) & (!g1781)) + ((!g708) & (!g731) & (!g1778) & (!g1814) & (!g1780) & (g1781)) + ((!g708) & (!g731) & (!g1778) & (!g1814) & (g1780) & (!g1781)) + ((!g708) & (!g731) & (!g1778) & (!g1814) & (g1780) & (g1781)) + ((!g708) & (!g731) & (!g1778) & (g1814) & (!g1780) & (!g1781)) + ((!g708) & (!g731) & (!g1778) & (g1814) & (!g1780) & (g1781)) + ((!g708) & (!g731) & (!g1778) & (g1814) & (g1780) & (!g1781)) + ((!g708) & (!g731) & (!g1778) & (g1814) & (g1780) & (g1781)) + ((!g708) & (!g731) & (g1778) & (!g1814) & (!g1780) & (!g1781)) + ((!g708) & (!g731) & (g1778) & (!g1814) & (!g1780) & (g1781)) + ((!g708) & (!g731) & (g1778) & (!g1814) & (g1780) & (!g1781)) + ((!g708) & (!g731) & (g1778) & (!g1814) & (g1780) & (g1781)) + ((!g708) & (!g731) & (g1778) & (g1814) & (!g1780) & (!g1781)) + ((!g708) & (g731) & (!g1778) & (!g1814) & (!g1780) & (!g1781)) + ((!g708) & (g731) & (!g1778) & (!g1814) & (!g1780) & (g1781)) + ((!g708) & (g731) & (!g1778) & (!g1814) & (g1780) & (!g1781)) + ((!g708) & (g731) & (!g1778) & (!g1814) & (g1780) & (g1781)) + ((!g708) & (g731) & (g1778) & (!g1814) & (!g1780) & (!g1781)) + ((g708) & (!g731) & (!g1778) & (!g1814) & (!g1780) & (!g1781)) + ((g708) & (!g731) & (!g1778) & (!g1814) & (!g1780) & (g1781)) + ((g708) & (!g731) & (!g1778) & (!g1814) & (g1780) & (!g1781)) + ((g708) & (!g731) & (!g1778) & (!g1814) & (g1780) & (g1781)) + ((g708) & (!g731) & (!g1778) & (g1814) & (!g1780) & (!g1781)) + ((g708) & (!g731) & (g1778) & (!g1814) & (!g1780) & (!g1781)) + ((g708) & (!g731) & (g1778) & (!g1814) & (!g1780) & (g1781)) + ((g708) & (!g731) & (g1778) & (!g1814) & (g1780) & (!g1781)) + ((g708) & (!g731) & (g1778) & (!g1814) & (g1780) & (g1781)) + ((g708) & (g731) & (!g1778) & (!g1814) & (!g1780) & (!g1781)));
	assign g1849 = (((!g827) & (!g754) & (g1847) & (!g1848)) + ((!g827) & (!g754) & (g1847) & (g1848)) + ((!g827) & (g754) & (g1847) & (!g1848)) + ((!g827) & (g754) & (g1847) & (g1848)) + ((g827) & (!g754) & (!g1847) & (!g1848)) + ((g827) & (!g754) & (g1847) & (g1848)) + ((g827) & (g754) & (!g1847) & (g1848)) + ((g827) & (g754) & (g1847) & (!g1848)));
	assign g1850 = (((!g34) & (!g36) & (!reset) & (g756) & (!g777)) + ((!g34) & (!g36) & (!reset) & (g756) & (g777)) + ((!g34) & (g36) & (!reset) & (!g756) & (g777)) + ((!g34) & (g36) & (!reset) & (g756) & (g777)) + ((g34) & (!g36) & (!reset) & (g756) & (!g777)) + ((g34) & (!g36) & (!reset) & (g756) & (g777)) + ((g34) & (g36) & (!reset) & (g756) & (!g777)) + ((g34) & (g36) & (!reset) & (g756) & (g777)));
	assign g7763 = (((!g832) & (g3365) & (!g1851)) + ((!g832) & (g3365) & (g1851)) + ((g832) & (!g3365) & (g1851)) + ((g832) & (g3365) & (g1851)));
	assign g1852 = (((!g34) & (!g36) & (!reset) & (g757) & (!g1851)) + ((!g34) & (!g36) & (!reset) & (g757) & (g1851)) + ((!g34) & (g36) & (!reset) & (!g757) & (g1851)) + ((!g34) & (g36) & (!reset) & (g757) & (g1851)) + ((g34) & (!g36) & (!reset) & (g757) & (!g1851)) + ((g34) & (!g36) & (!reset) & (g757) & (g1851)) + ((g34) & (g36) & (!reset) & (g757) & (!g1851)) + ((g34) & (g36) & (!reset) & (g757) & (g1851)));
	assign g7764 = (((!g832) & (g3367) & (!g1853)) + ((!g832) & (g3367) & (g1853)) + ((g832) & (!g3367) & (g1853)) + ((g832) & (g3367) & (g1853)));
	assign g1854 = (((!g34) & (!g36) & (!reset) & (g758) & (!g1853)) + ((!g34) & (!g36) & (!reset) & (g758) & (g1853)) + ((!g34) & (g36) & (!reset) & (!g758) & (g1853)) + ((!g34) & (g36) & (!reset) & (g758) & (g1853)) + ((g34) & (!g36) & (!reset) & (g758) & (!g1853)) + ((g34) & (!g36) & (!reset) & (g758) & (g1853)) + ((g34) & (g36) & (!reset) & (g758) & (!g1853)) + ((g34) & (g36) & (!reset) & (g758) & (g1853)));
	assign g7765 = (((!g832) & (g3368) & (!g1855)) + ((!g832) & (g3368) & (g1855)) + ((g832) & (!g3368) & (g1855)) + ((g832) & (g3368) & (g1855)));
	assign g1856 = (((!g34) & (!g36) & (!reset) & (g759) & (!g1855)) + ((!g34) & (!g36) & (!reset) & (g759) & (g1855)) + ((!g34) & (g36) & (!reset) & (!g759) & (g1855)) + ((!g34) & (g36) & (!reset) & (g759) & (g1855)) + ((g34) & (!g36) & (!reset) & (g759) & (!g1855)) + ((g34) & (!g36) & (!reset) & (g759) & (g1855)) + ((g34) & (g36) & (!reset) & (g759) & (!g1855)) + ((g34) & (g36) & (!reset) & (g759) & (g1855)));
	assign g7766 = (((!g832) & (g3369) & (!g1857)) + ((!g832) & (g3369) & (g1857)) + ((g832) & (!g3369) & (g1857)) + ((g832) & (g3369) & (g1857)));
	assign g1858 = (((!g34) & (!g36) & (!reset) & (g761) & (!g1857)) + ((!g34) & (!g36) & (!reset) & (g761) & (g1857)) + ((!g34) & (g36) & (!reset) & (!g761) & (g1857)) + ((!g34) & (g36) & (!reset) & (g761) & (g1857)) + ((g34) & (!g36) & (!reset) & (g761) & (!g1857)) + ((g34) & (!g36) & (!reset) & (g761) & (g1857)) + ((g34) & (g36) & (!reset) & (g761) & (!g1857)) + ((g34) & (g36) & (!reset) & (g761) & (g1857)));
	assign g7767 = (((!g832) & (g3371) & (!g1859)) + ((!g832) & (g3371) & (g1859)) + ((g832) & (!g3371) & (g1859)) + ((g832) & (g3371) & (g1859)));
	assign g1860 = (((!g34) & (!g36) & (!reset) & (g762) & (!g1859)) + ((!g34) & (!g36) & (!reset) & (g762) & (g1859)) + ((!g34) & (g36) & (!reset) & (!g762) & (g1859)) + ((!g34) & (g36) & (!reset) & (g762) & (g1859)) + ((g34) & (!g36) & (!reset) & (g762) & (!g1859)) + ((g34) & (!g36) & (!reset) & (g762) & (g1859)) + ((g34) & (g36) & (!reset) & (g762) & (!g1859)) + ((g34) & (g36) & (!reset) & (g762) & (g1859)));
	assign g7768 = (((!g832) & (g3373) & (!g1861)) + ((!g832) & (g3373) & (g1861)) + ((g832) & (!g3373) & (g1861)) + ((g832) & (g3373) & (g1861)));
	assign g1862 = (((!g34) & (!g36) & (!reset) & (g763) & (!g1861)) + ((!g34) & (!g36) & (!reset) & (g763) & (g1861)) + ((!g34) & (g36) & (!reset) & (!g763) & (g1861)) + ((!g34) & (g36) & (!reset) & (g763) & (g1861)) + ((g34) & (!g36) & (!reset) & (g763) & (!g1861)) + ((g34) & (!g36) & (!reset) & (g763) & (g1861)) + ((g34) & (g36) & (!reset) & (g763) & (!g1861)) + ((g34) & (g36) & (!reset) & (g763) & (g1861)));
	assign g7769 = (((!g832) & (g3375) & (!g1863)) + ((!g832) & (g3375) & (g1863)) + ((g832) & (!g3375) & (g1863)) + ((g832) & (g3375) & (g1863)));
	assign g1864 = (((!g34) & (!g36) & (!reset) & (g764) & (!g1863)) + ((!g34) & (!g36) & (!reset) & (g764) & (g1863)) + ((!g34) & (g36) & (!reset) & (!g764) & (g1863)) + ((!g34) & (g36) & (!reset) & (g764) & (g1863)) + ((g34) & (!g36) & (!reset) & (g764) & (!g1863)) + ((g34) & (!g36) & (!reset) & (g764) & (g1863)) + ((g34) & (g36) & (!reset) & (g764) & (!g1863)) + ((g34) & (g36) & (!reset) & (g764) & (g1863)));
	assign g7770 = (((!g832) & (g3377) & (!g1865)) + ((!g832) & (g3377) & (g1865)) + ((g832) & (!g3377) & (g1865)) + ((g832) & (g3377) & (g1865)));
	assign g1866 = (((!g34) & (!g36) & (!reset) & (g766) & (!g1865)) + ((!g34) & (!g36) & (!reset) & (g766) & (g1865)) + ((!g34) & (g36) & (!reset) & (!g766) & (g1865)) + ((!g34) & (g36) & (!reset) & (g766) & (g1865)) + ((g34) & (!g36) & (!reset) & (g766) & (!g1865)) + ((g34) & (!g36) & (!reset) & (g766) & (g1865)) + ((g34) & (g36) & (!reset) & (g766) & (!g1865)) + ((g34) & (g36) & (!reset) & (g766) & (g1865)));
	assign g7771 = (((!g832) & (g3379) & (!g1867)) + ((!g832) & (g3379) & (g1867)) + ((g832) & (!g3379) & (g1867)) + ((g832) & (g3379) & (g1867)));
	assign g1868 = (((!g34) & (!g36) & (!reset) & (g767) & (!g1867)) + ((!g34) & (!g36) & (!reset) & (g767) & (g1867)) + ((!g34) & (g36) & (!reset) & (!g767) & (g1867)) + ((!g34) & (g36) & (!reset) & (g767) & (g1867)) + ((g34) & (!g36) & (!reset) & (g767) & (!g1867)) + ((g34) & (!g36) & (!reset) & (g767) & (g1867)) + ((g34) & (g36) & (!reset) & (g767) & (!g1867)) + ((g34) & (g36) & (!reset) & (g767) & (g1867)));
	assign g7772 = (((!g832) & (g3381) & (!g1869)) + ((!g832) & (g3381) & (g1869)) + ((g832) & (!g3381) & (g1869)) + ((g832) & (g3381) & (g1869)));
	assign g1870 = (((!g34) & (!g36) & (!reset) & (g768) & (!g1869)) + ((!g34) & (!g36) & (!reset) & (g768) & (g1869)) + ((!g34) & (g36) & (!reset) & (!g768) & (g1869)) + ((!g34) & (g36) & (!reset) & (g768) & (g1869)) + ((g34) & (!g36) & (!reset) & (g768) & (!g1869)) + ((g34) & (!g36) & (!reset) & (g768) & (g1869)) + ((g34) & (g36) & (!reset) & (g768) & (!g1869)) + ((g34) & (g36) & (!reset) & (g768) & (g1869)));
	assign g7773 = (((!g832) & (g3383) & (!g1871)) + ((!g832) & (g3383) & (g1871)) + ((g832) & (!g3383) & (g1871)) + ((g832) & (g3383) & (g1871)));
	assign g1872 = (((!g34) & (!g36) & (!reset) & (g769) & (!g1871)) + ((!g34) & (!g36) & (!reset) & (g769) & (g1871)) + ((!g34) & (g36) & (!reset) & (!g769) & (g1871)) + ((!g34) & (g36) & (!reset) & (g769) & (g1871)) + ((g34) & (!g36) & (!reset) & (g769) & (!g1871)) + ((g34) & (!g36) & (!reset) & (g769) & (g1871)) + ((g34) & (g36) & (!reset) & (g769) & (!g1871)) + ((g34) & (g36) & (!reset) & (g769) & (g1871)));
	assign g7774 = (((!g832) & (g3384) & (!g1873)) + ((!g832) & (g3384) & (g1873)) + ((g832) & (!g3384) & (g1873)) + ((g832) & (g3384) & (g1873)));
	assign g1874 = (((!g34) & (!g36) & (!reset) & (g771) & (!g1873)) + ((!g34) & (!g36) & (!reset) & (g771) & (g1873)) + ((!g34) & (g36) & (!reset) & (!g771) & (g1873)) + ((!g34) & (g36) & (!reset) & (g771) & (g1873)) + ((g34) & (!g36) & (!reset) & (g771) & (!g1873)) + ((g34) & (!g36) & (!reset) & (g771) & (g1873)) + ((g34) & (g36) & (!reset) & (g771) & (!g1873)) + ((g34) & (g36) & (!reset) & (g771) & (g1873)));
	assign g7775 = (((!g832) & (g3386) & (!g1875)) + ((!g832) & (g3386) & (g1875)) + ((g832) & (!g3386) & (g1875)) + ((g832) & (g3386) & (g1875)));
	assign g1876 = (((!g34) & (!g36) & (!reset) & (g772) & (!g1875)) + ((!g34) & (!g36) & (!reset) & (g772) & (g1875)) + ((!g34) & (g36) & (!reset) & (!g772) & (g1875)) + ((!g34) & (g36) & (!reset) & (g772) & (g1875)) + ((g34) & (!g36) & (!reset) & (g772) & (!g1875)) + ((g34) & (!g36) & (!reset) & (g772) & (g1875)) + ((g34) & (g36) & (!reset) & (g772) & (!g1875)) + ((g34) & (g36) & (!reset) & (g772) & (g1875)));
	assign g7776 = (((!g832) & (g3388) & (!g1877)) + ((!g832) & (g3388) & (g1877)) + ((g832) & (!g3388) & (g1877)) + ((g832) & (g3388) & (g1877)));
	assign g1878 = (((!g34) & (!g36) & (!reset) & (g773) & (!g1877)) + ((!g34) & (!g36) & (!reset) & (g773) & (g1877)) + ((!g34) & (g36) & (!reset) & (!g773) & (g1877)) + ((!g34) & (g36) & (!reset) & (g773) & (g1877)) + ((g34) & (!g36) & (!reset) & (g773) & (!g1877)) + ((g34) & (!g36) & (!reset) & (g773) & (g1877)) + ((g34) & (g36) & (!reset) & (g773) & (!g1877)) + ((g34) & (g36) & (!reset) & (g773) & (g1877)));
	assign g7777 = (((!g832) & (g3390) & (!g1879)) + ((!g832) & (g3390) & (g1879)) + ((g832) & (!g3390) & (g1879)) + ((g832) & (g3390) & (g1879)));
	assign g1880 = (((!g34) & (!g36) & (!reset) & (g774) & (!g1879)) + ((!g34) & (!g36) & (!reset) & (g774) & (g1879)) + ((!g34) & (g36) & (!reset) & (!g774) & (g1879)) + ((!g34) & (g36) & (!reset) & (g774) & (g1879)) + ((g34) & (!g36) & (!reset) & (g774) & (!g1879)) + ((g34) & (!g36) & (!reset) & (g774) & (g1879)) + ((g34) & (g36) & (!reset) & (g774) & (!g1879)) + ((g34) & (g36) & (!reset) & (g774) & (g1879)));
	assign g7778 = (((!g2017) & (g7083) & (!g1881)) + ((!g2017) & (g7083) & (g1881)) + ((g2017) & (!g7083) & (g1881)) + ((g2017) & (g7083) & (g1881)));
	assign g1882 = (((!g827) & (!g754) & (!g777) & (!g1847) & (g1881) & (!g1848)) + ((!g827) & (!g754) & (!g777) & (!g1847) & (g1881) & (g1848)) + ((!g827) & (!g754) & (!g777) & (g1847) & (g1881) & (!g1848)) + ((!g827) & (!g754) & (!g777) & (g1847) & (g1881) & (g1848)) + ((!g827) & (!g754) & (g777) & (!g1847) & (g1881) & (!g1848)) + ((!g827) & (!g754) & (g777) & (!g1847) & (g1881) & (g1848)) + ((!g827) & (!g754) & (g777) & (g1847) & (g1881) & (!g1848)) + ((!g827) & (!g754) & (g777) & (g1847) & (g1881) & (g1848)) + ((!g827) & (g754) & (!g777) & (!g1847) & (g1881) & (!g1848)) + ((!g827) & (g754) & (!g777) & (!g1847) & (g1881) & (g1848)) + ((!g827) & (g754) & (!g777) & (g1847) & (g1881) & (!g1848)) + ((!g827) & (g754) & (!g777) & (g1847) & (g1881) & (g1848)) + ((!g827) & (g754) & (g777) & (!g1847) & (g1881) & (!g1848)) + ((!g827) & (g754) & (g777) & (!g1847) & (g1881) & (g1848)) + ((!g827) & (g754) & (g777) & (g1847) & (g1881) & (!g1848)) + ((!g827) & (g754) & (g777) & (g1847) & (g1881) & (g1848)) + ((g827) & (!g754) & (!g777) & (!g1847) & (g1881) & (!g1848)) + ((g827) & (!g754) & (!g777) & (!g1847) & (g1881) & (g1848)) + ((g827) & (!g754) & (!g777) & (g1847) & (!g1881) & (!g1848)) + ((g827) & (!g754) & (!g777) & (g1847) & (g1881) & (g1848)) + ((g827) & (!g754) & (g777) & (!g1847) & (!g1881) & (!g1848)) + ((g827) & (!g754) & (g777) & (!g1847) & (!g1881) & (g1848)) + ((g827) & (!g754) & (g777) & (g1847) & (!g1881) & (g1848)) + ((g827) & (!g754) & (g777) & (g1847) & (g1881) & (!g1848)) + ((g827) & (g754) & (!g777) & (!g1847) & (!g1881) & (!g1848)) + ((g827) & (g754) & (!g777) & (!g1847) & (g1881) & (g1848)) + ((g827) & (g754) & (!g777) & (g1847) & (!g1881) & (!g1848)) + ((g827) & (g754) & (!g777) & (g1847) & (!g1881) & (g1848)) + ((g827) & (g754) & (g777) & (!g1847) & (!g1881) & (g1848)) + ((g827) & (g754) & (g777) & (!g1847) & (g1881) & (!g1848)) + ((g827) & (g754) & (g777) & (g1847) & (g1881) & (!g1848)) + ((g827) & (g754) & (g777) & (g1847) & (g1881) & (g1848)));
	assign g1883 = (((!reset) & (!g779) & (!g827) & (!g830) & (!g831)) + ((!reset) & (!g779) & (!g827) & (!g830) & (g831)) + ((!reset) & (g779) & (!g827) & (!g830) & (!g831)) + ((!reset) & (g779) & (!g827) & (!g830) & (g831)) + ((!reset) & (g779) & (!g827) & (g830) & (!g831)) + ((!reset) & (g779) & (!g827) & (g830) & (g831)) + ((!reset) & (g779) & (g827) & (!g830) & (g831)) + ((!reset) & (g779) & (g827) & (g830) & (!g831)) + ((!reset) & (g779) & (g827) & (g830) & (g831)) + ((reset) & (!g779) & (!g827) & (!g830) & (!g831)) + ((reset) & (!g779) & (!g827) & (!g830) & (g831)) + ((reset) & (!g779) & (!g827) & (g830) & (!g831)) + ((reset) & (!g779) & (!g827) & (g830) & (g831)) + ((reset) & (!g779) & (g827) & (!g830) & (!g831)) + ((reset) & (!g779) & (g827) & (!g830) & (g831)) + ((reset) & (!g779) & (g827) & (g830) & (!g831)) + ((reset) & (!g779) & (g827) & (g830) & (g831)) + ((reset) & (g779) & (!g827) & (!g830) & (!g831)) + ((reset) & (g779) & (!g827) & (!g830) & (g831)) + ((reset) & (g779) & (!g827) & (g830) & (!g831)) + ((reset) & (g779) & (!g827) & (g830) & (g831)) + ((reset) & (g779) & (g827) & (!g830) & (!g831)) + ((reset) & (g779) & (g827) & (!g830) & (g831)) + ((reset) & (g779) & (g827) & (g830) & (!g831)) + ((reset) & (g779) & (g827) & (g830) & (g831)));
	assign g7779 = (((!g3429) & (g3428) & (!g1884)) + ((!g3429) & (g3428) & (g1884)) + ((g3429) & (!g3428) & (g1884)) + ((g3429) & (g3428) & (g1884)));
	assign g1885 = (((!g790) & (!g827) & (g1884)) + ((!g790) & (g827) & (g1884)) + ((g790) & (!g827) & (g1884)) + ((g790) & (g827) & (!g1884)));
	assign g7780 = (((!g3464) & (g3462) & (!g1886)) + ((!g3464) & (g3462) & (g1886)) + ((g3464) & (!g3462) & (g1886)) + ((g3464) & (g3462) & (g1886)));
	assign g1887 = (((!g792) & (!g827) & (g1886)) + ((!g792) & (g827) & (g1886)) + ((g792) & (!g827) & (g1886)) + ((g792) & (g827) & (!g1886)));
	assign g7781 = (((!g3499) & (g3498) & (!g1888)) + ((!g3499) & (g3498) & (g1888)) + ((g3499) & (!g3498) & (g1888)) + ((g3499) & (g3498) & (g1888)));
	assign g1889 = (((!g794) & (!g827) & (g1888)) + ((!g794) & (g827) & (g1888)) + ((g794) & (!g827) & (g1888)) + ((g794) & (g827) & (!g1888)));
	assign g7782 = (((!g3429) & (g3534) & (!g1890)) + ((!g3429) & (g3534) & (g1890)) + ((g3429) & (!g3534) & (g1890)) + ((g3429) & (g3534) & (g1890)));
	assign g1891 = (((!g800) & (!g827) & (g1890)) + ((!g800) & (g827) & (g1890)) + ((g800) & (!g827) & (g1890)) + ((g800) & (g827) & (!g1890)));
	assign g7783 = (((!g2017) & (g7053) & (!g1892)) + ((!g2017) & (g7053) & (g1892)) + ((g2017) & (!g7053) & (g1892)) + ((g2017) & (g7053) & (g1892)));
	assign g1893 = (((!g802) & (!g827) & (g1892)) + ((!g802) & (g827) & (g1892)) + ((g802) & (!g827) & (g1892)) + ((g802) & (g827) & (!g1892)));
	assign g7784 = (((!g3499) & (g3587) & (!g1894)) + ((!g3499) & (g3587) & (g1894)) + ((g3499) & (!g3587) & (g1894)) + ((g3499) & (g3587) & (g1894)));
	assign g1895 = (((!g804) & (!g827) & (g1894)) + ((!g804) & (g827) & (g1894)) + ((g804) & (!g827) & (g1894)) + ((g804) & (g827) & (!g1894)));
	assign g7785 = (((!g3464) & (g3620) & (!g1896)) + ((!g3464) & (g3620) & (g1896)) + ((g3464) & (!g3620) & (g1896)) + ((g3464) & (g3620) & (g1896)));
	assign g1897 = (((!g806) & (!g827) & (g1896)) + ((!g806) & (g827) & (g1896)) + ((g806) & (!g827) & (g1896)) + ((g806) & (g827) & (!g1896)));
	assign g7786 = (((!g3499) & (g3653) & (!g1898)) + ((!g3499) & (g3653) & (g1898)) + ((g3499) & (!g3653) & (g1898)) + ((g3499) & (g3653) & (g1898)));
	assign g1899 = (((!g808) & (!g827) & (g1898)) + ((!g808) & (g827) & (g1898)) + ((g808) & (!g827) & (g1898)) + ((g808) & (g827) & (!g1898)));
	assign g7787 = (((!g3464) & (g3688) & (!g1900)) + ((!g3464) & (g3688) & (g1900)) + ((g3464) & (!g3688) & (g1900)) + ((g3464) & (g3688) & (g1900)));
	assign g1901 = (((!g810) & (!g827) & (g1900)) + ((!g810) & (g827) & (g1900)) + ((g810) & (!g827) & (g1900)) + ((g810) & (g827) & (!g1900)));
	assign g7788 = (((!g2017) & (g7012) & (!g1902)) + ((!g2017) & (g7012) & (g1902)) + ((g2017) & (!g7012) & (g1902)) + ((g2017) & (g7012) & (g1902)));
	assign g1903 = (((!g812) & (!g827) & (g1902)) + ((!g812) & (g827) & (g1902)) + ((g812) & (!g827) & (g1902)) + ((g812) & (g827) & (!g1902)));
	assign g7789 = (((!g3429) & (g3744) & (!g1904)) + ((!g3429) & (g3744) & (g1904)) + ((g3429) & (!g3744) & (g1904)) + ((g3429) & (g3744) & (g1904)));
	assign g1905 = (((!g814) & (!g827) & (g1904)) + ((!g814) & (g827) & (g1904)) + ((g814) & (!g827) & (g1904)) + ((g814) & (g827) & (!g1904)));
	assign g7790 = (((!g3464) & (g3777) & (!g1906)) + ((!g3464) & (g3777) & (g1906)) + ((g3464) & (!g3777) & (g1906)) + ((g3464) & (g3777) & (g1906)));
	assign g1907 = (((!g816) & (!g827) & (g1906)) + ((!g816) & (g827) & (g1906)) + ((g816) & (!g827) & (g1906)) + ((g816) & (g827) & (!g1906)));
	assign g7791 = (((!g3499) & (g3810) & (!g1908)) + ((!g3499) & (g3810) & (g1908)) + ((g3499) & (!g3810) & (g1908)) + ((g3499) & (g3810) & (g1908)));
	assign g1909 = (((!g818) & (!g827) & (g1908)) + ((!g818) & (g827) & (g1908)) + ((g818) & (!g827) & (g1908)) + ((g818) & (g827) & (!g1908)));
	assign g7792 = (((!g3429) & (g3845) & (!g1910)) + ((!g3429) & (g3845) & (g1910)) + ((g3429) & (!g3845) & (g1910)) + ((g3429) & (g3845) & (g1910)));
	assign g1911 = (((!g820) & (!g827) & (g1910)) + ((!g820) & (g827) & (g1910)) + ((g820) & (!g827) & (g1910)) + ((g820) & (g827) & (!g1910)));
	assign g7793 = (((!g2017) & (g6982) & (!g1912)) + ((!g2017) & (g6982) & (g1912)) + ((g2017) & (!g6982) & (g1912)) + ((g2017) & (g6982) & (g1912)));
	assign g1913 = (((!g822) & (!g827) & (g1912)) + ((!g822) & (g827) & (g1912)) + ((g822) & (!g827) & (g1912)) + ((g822) & (g827) & (!g1912)));
	assign g7794 = (((!g3869) & (!g3868) & (g1914)) + ((!g3869) & (g3868) & (g1914)) + ((g3869) & (g3868) & (!g1914)) + ((g3869) & (g3868) & (g1914)));
	assign g7795 = (((!g3869) & (!g3872) & (g1915)) + ((!g3869) & (g3872) & (g1915)) + ((g3869) & (g3872) & (!g1915)) + ((g3869) & (g3872) & (g1915)));
	assign g7796 = (((!g3869) & (!g3873) & (g1916)) + ((!g3869) & (g3873) & (g1916)) + ((g3869) & (g3873) & (!g1916)) + ((g3869) & (g3873) & (g1916)));
	assign g7797 = (((!g3869) & (!g3874) & (g1917)) + ((!g3869) & (g3874) & (g1917)) + ((g3869) & (g3874) & (!g1917)) + ((g3869) & (g3874) & (g1917)));
	assign g7798 = (((!g3869) & (!g3875) & (g1918)) + ((!g3869) & (g3875) & (g1918)) + ((g3869) & (g3875) & (!g1918)) + ((g3869) & (g3875) & (g1918)));
	assign g7799 = (((!g3869) & (!g3876) & (g1919)) + ((!g3869) & (g3876) & (g1919)) + ((g3869) & (g3876) & (!g1919)) + ((g3869) & (g3876) & (g1919)));
	assign g7800 = (((!g3869) & (!g3877) & (g1920)) + ((!g3869) & (g3877) & (g1920)) + ((g3869) & (g3877) & (!g1920)) + ((g3869) & (g3877) & (g1920)));
	assign g1921 = (((!g1915) & (!g1916) & (!g1917) & (!g1918) & (!g1919) & (g1920)));
	assign g7801 = (((!g3869) & (!g3878) & (g1922)) + ((!g3869) & (g3878) & (g1922)) + ((g3869) & (g3878) & (!g1922)) + ((g3869) & (g3878) & (g1922)));
	assign g1923 = (((g1914) & (g1921) & (g1922)));
	assign g7802 = (((!g3880) & (g3879) & (!g1924)) + ((!g3880) & (g3879) & (g1924)) + ((g3880) & (!g3879) & (g1924)) + ((g3880) & (g3879) & (g1924)));
	assign g7803 = (((!g3880) & (g3881) & (!g1925)) + ((!g3880) & (g3881) & (g1925)) + ((g3880) & (!g3881) & (g1925)) + ((g3880) & (g3881) & (g1925)));
	assign g7804 = (((!g3880) & (g3884) & (!g1926)) + ((!g3880) & (g3884) & (g1926)) + ((g3880) & (!g3884) & (g1926)) + ((g3880) & (g3884) & (g1926)));
	assign g7805 = (((!g3880) & (g3885) & (!g1927)) + ((!g3880) & (g3885) & (g1927)) + ((g3880) & (!g3885) & (g1927)) + ((g3880) & (g3885) & (g1927)));
	assign g7806 = (((!g3880) & (g3886) & (!g1928)) + ((!g3880) & (g3886) & (g1928)) + ((g3880) & (!g3886) & (g1928)) + ((g3880) & (g3886) & (g1928)));
	assign g7807 = (((!g3880) & (g3887) & (!g1929)) + ((!g3880) & (g3887) & (g1929)) + ((g3880) & (!g3887) & (g1929)) + ((g3880) & (g3887) & (g1929)));
	assign g1930 = (((g1924) & (!g1925) & (!g1926) & (!g1927) & (!g1928) & (!g1929)));
	assign g7808 = (((!g3880) & (g3888) & (!g1931)) + ((!g3880) & (g3888) & (g1931)) + ((g3880) & (!g3888) & (g1931)) + ((g3880) & (g3888) & (g1931)));
	assign g7809 = (((!g3880) & (g3889) & (!g1932)) + ((!g3880) & (g3889) & (g1932)) + ((g3880) & (!g3889) & (g1932)) + ((g3880) & (g3889) & (g1932)));
	assign g1933 = (((!g1931) & (g1932)));
	assign g1934 = (((g1930) & (g1933)));
	assign g7810 = (((!reset) & (g3890) & (!g1935)) + ((!reset) & (g3890) & (g1935)) + ((reset) & (!g3890) & (g1935)) + ((reset) & (g3890) & (g1935)));
	assign g1936 = (((!g827) & (!g831) & (!g1935) & (!start)) + ((!g827) & (!g831) & (g1935) & (!start)) + ((g827) & (g831) & (!g1935) & (!start)) + ((g827) & (g831) & (!g1935) & (start)));
	assign g1937 = (((!reset) & (!g827) & (g830) & (g1923) & (g1934) & (!g1936)) + ((!reset) & (!g827) & (g830) & (g1923) & (g1934) & (g1936)) + ((!reset) & (g827) & (!g830) & (!g1923) & (!g1934) & (g1936)) + ((!reset) & (g827) & (!g830) & (!g1923) & (g1934) & (g1936)) + ((!reset) & (g827) & (!g830) & (g1923) & (!g1934) & (g1936)) + ((!reset) & (g827) & (!g830) & (g1923) & (g1934) & (g1936)) + ((!reset) & (g827) & (g830) & (!g1923) & (!g1934) & (!g1936)) + ((!reset) & (g827) & (g830) & (!g1923) & (!g1934) & (g1936)) + ((!reset) & (g827) & (g830) & (!g1923) & (g1934) & (!g1936)) + ((!reset) & (g827) & (g830) & (!g1923) & (g1934) & (g1936)) + ((!reset) & (g827) & (g830) & (g1923) & (!g1934) & (!g1936)) + ((!reset) & (g827) & (g830) & (g1923) & (!g1934) & (g1936)) + ((!reset) & (g827) & (g830) & (g1923) & (g1934) & (!g1936)) + ((!reset) & (g827) & (g830) & (g1923) & (g1934) & (g1936)));
	assign g1938 = (((!reset) & (!g831)));
	assign g7811 = (((!g3429) & (g3895) & (!g1939)) + ((!g3429) & (g3895) & (g1939)) + ((g3429) & (!g3895) & (g1939)) + ((g3429) & (g3895) & (g1939)));
	assign g7812 = (((!g3464) & (g3901) & (!g1940)) + ((!g3464) & (g3901) & (g1940)) + ((g3464) & (!g3901) & (g1940)) + ((g3464) & (g3901) & (g1940)));
	assign g7813 = (((!g3429) & (g3904) & (!g1941)) + ((!g3429) & (g3904) & (g1941)) + ((g3429) & (!g3904) & (g1941)) + ((g3429) & (g3904) & (g1941)));
	assign g7814 = (((!g3464) & (g3911) & (!g1942)) + ((!g3464) & (g3911) & (g1942)) + ((g3464) & (!g3911) & (g1942)) + ((g3464) & (g3911) & (g1942)));
	assign g1943 = (((!g1890) & (!g1906) & (!g1939) & (!g1940) & (g1941) & (g1942)) + ((!g1890) & (!g1906) & (!g1939) & (g1940) & (g1941) & (g1942)) + ((!g1890) & (!g1906) & (g1939) & (!g1940) & (g1941) & (g1942)) + ((!g1890) & (!g1906) & (g1939) & (g1940) & (!g1941) & (g1942)) + ((!g1890) & (!g1906) & (g1939) & (g1940) & (g1941) & (!g1942)) + ((!g1890) & (!g1906) & (g1939) & (g1940) & (g1941) & (g1942)) + ((!g1890) & (g1906) & (!g1939) & (!g1940) & (g1941) & (g1942)) + ((!g1890) & (g1906) & (!g1939) & (g1940) & (g1941) & (g1942)) + ((!g1890) & (g1906) & (g1939) & (!g1940) & (g1941) & (g1942)) + ((!g1890) & (g1906) & (g1939) & (g1940) & (!g1941) & (g1942)) + ((!g1890) & (g1906) & (g1939) & (g1940) & (g1941) & (!g1942)) + ((!g1890) & (g1906) & (g1939) & (g1940) & (g1941) & (g1942)) + ((g1890) & (!g1906) & (!g1939) & (!g1940) & (g1941) & (g1942)) + ((g1890) & (!g1906) & (!g1939) & (g1940) & (g1941) & (g1942)) + ((g1890) & (!g1906) & (g1939) & (!g1940) & (g1941) & (g1942)) + ((g1890) & (!g1906) & (g1939) & (g1940) & (!g1941) & (g1942)) + ((g1890) & (!g1906) & (g1939) & (g1940) & (g1941) & (!g1942)) + ((g1890) & (!g1906) & (g1939) & (g1940) & (g1941) & (g1942)) + ((g1890) & (g1906) & (!g1939) & (!g1940) & (g1941) & (g1942)) + ((g1890) & (g1906) & (!g1939) & (g1940) & (!g1941) & (g1942)) + ((g1890) & (g1906) & (!g1939) & (g1940) & (g1941) & (!g1942)) + ((g1890) & (g1906) & (!g1939) & (g1940) & (g1941) & (g1942)) + ((g1890) & (g1906) & (g1939) & (!g1940) & (!g1941) & (g1942)) + ((g1890) & (g1906) & (g1939) & (!g1940) & (g1941) & (!g1942)) + ((g1890) & (g1906) & (g1939) & (!g1940) & (g1941) & (g1942)) + ((g1890) & (g1906) & (g1939) & (g1940) & (!g1941) & (g1942)) + ((g1890) & (g1906) & (g1939) & (g1940) & (g1941) & (!g1942)) + ((g1890) & (g1906) & (g1939) & (g1940) & (g1941) & (g1942)));
	assign g7815 = (((!g3429) & (g3920) & (!g1944)) + ((!g3429) & (g3920) & (g1944)) + ((g3429) & (!g3920) & (g1944)) + ((g3429) & (g3920) & (g1944)));
	assign g7816 = (((!g3464) & (g3924) & (!g1945)) + ((!g3464) & (g3924) & (g1945)) + ((g3464) & (!g3924) & (g1945)) + ((g3464) & (g3924) & (g1945)));
	assign g7817 = (((!g3429) & (g3929) & (!g1946)) + ((!g3429) & (g3929) & (g1946)) + ((g3429) & (!g3929) & (g1946)) + ((g3429) & (g3929) & (g1946)));
	assign g7818 = (((!g3464) & (g3933) & (!g1947)) + ((!g3464) & (g3933) & (g1947)) + ((g3464) & (!g3933) & (g1947)) + ((g3464) & (g3933) & (g1947)));
	assign g7819 = (((!g3429) & (g3938) & (!g1948)) + ((!g3429) & (g3938) & (g1948)) + ((g3429) & (!g3938) & (g1948)) + ((g3429) & (g3938) & (g1948)));
	assign g7820 = (((!g3464) & (g3941) & (!g1949)) + ((!g3464) & (g3941) & (g1949)) + ((g3464) & (!g3941) & (g1949)) + ((g3464) & (g3941) & (g1949)));
	assign g1950 = (((!g1948) & (g1949)) + ((g1948) & (!g1949)));
	assign g1951 = (((!g1943) & (!g1944) & (!g1945) & (g1946) & (g1947) & (g1950)) + ((!g1943) & (!g1944) & (g1945) & (g1946) & (g1947) & (g1950)) + ((!g1943) & (g1944) & (!g1945) & (g1946) & (g1947) & (g1950)) + ((!g1943) & (g1944) & (g1945) & (!g1946) & (g1947) & (g1950)) + ((!g1943) & (g1944) & (g1945) & (g1946) & (!g1947) & (g1950)) + ((!g1943) & (g1944) & (g1945) & (g1946) & (g1947) & (g1950)) + ((g1943) & (!g1944) & (!g1945) & (g1946) & (g1947) & (g1950)) + ((g1943) & (!g1944) & (g1945) & (!g1946) & (g1947) & (g1950)) + ((g1943) & (!g1944) & (g1945) & (g1946) & (!g1947) & (g1950)) + ((g1943) & (!g1944) & (g1945) & (g1946) & (g1947) & (g1950)) + ((g1943) & (g1944) & (!g1945) & (!g1946) & (g1947) & (g1950)) + ((g1943) & (g1944) & (!g1945) & (g1946) & (!g1947) & (g1950)) + ((g1943) & (g1944) & (!g1945) & (g1946) & (g1947) & (g1950)) + ((g1943) & (g1944) & (g1945) & (!g1946) & (g1947) & (g1950)) + ((g1943) & (g1944) & (g1945) & (g1946) & (!g1947) & (g1950)) + ((g1943) & (g1944) & (g1945) & (g1946) & (g1947) & (g1950)));
	assign g1952 = (((g1948) & (g1949)));
	assign g7821 = (((!g3429) & (g3944) & (!g1953)) + ((!g3429) & (g3944) & (g1953)) + ((g3429) & (!g3944) & (g1953)) + ((g3429) & (g3944) & (g1953)));
	assign g7822 = (((!g3464) & (g3947) & (!g1954)) + ((!g3464) & (g3947) & (g1954)) + ((g3464) & (!g3947) & (g1954)) + ((g3464) & (g3947) & (g1954)));
	assign g7823 = (((!g3429) & (g3950) & (!g1955)) + ((!g3429) & (g3950) & (g1955)) + ((g3429) & (!g3950) & (g1955)) + ((g3429) & (g3950) & (g1955)));
	assign g7824 = (((!g3464) & (g6971) & (!g1956)) + ((!g3464) & (g6971) & (g1956)) + ((g3464) & (!g6971) & (g1956)) + ((g3464) & (g6971) & (g1956)));
	assign g1957 = (((!g1951) & (!g1952) & (!g1953) & (!g1954) & (g1955) & (g1956)) + ((!g1951) & (!g1952) & (!g1953) & (g1954) & (g1955) & (g1956)) + ((!g1951) & (!g1952) & (g1953) & (!g1954) & (g1955) & (g1956)) + ((!g1951) & (!g1952) & (g1953) & (g1954) & (!g1955) & (g1956)) + ((!g1951) & (!g1952) & (g1953) & (g1954) & (g1955) & (!g1956)) + ((!g1951) & (!g1952) & (g1953) & (g1954) & (g1955) & (g1956)) + ((!g1951) & (g1952) & (!g1953) & (!g1954) & (g1955) & (g1956)) + ((!g1951) & (g1952) & (!g1953) & (g1954) & (!g1955) & (g1956)) + ((!g1951) & (g1952) & (!g1953) & (g1954) & (g1955) & (!g1956)) + ((!g1951) & (g1952) & (!g1953) & (g1954) & (g1955) & (g1956)) + ((!g1951) & (g1952) & (g1953) & (!g1954) & (!g1955) & (g1956)) + ((!g1951) & (g1952) & (g1953) & (!g1954) & (g1955) & (!g1956)) + ((!g1951) & (g1952) & (g1953) & (!g1954) & (g1955) & (g1956)) + ((!g1951) & (g1952) & (g1953) & (g1954) & (!g1955) & (g1956)) + ((!g1951) & (g1952) & (g1953) & (g1954) & (g1955) & (!g1956)) + ((!g1951) & (g1952) & (g1953) & (g1954) & (g1955) & (g1956)) + ((g1951) & (!g1952) & (!g1953) & (!g1954) & (g1955) & (g1956)) + ((g1951) & (!g1952) & (!g1953) & (g1954) & (!g1955) & (g1956)) + ((g1951) & (!g1952) & (!g1953) & (g1954) & (g1955) & (!g1956)) + ((g1951) & (!g1952) & (!g1953) & (g1954) & (g1955) & (g1956)) + ((g1951) & (!g1952) & (g1953) & (!g1954) & (!g1955) & (g1956)) + ((g1951) & (!g1952) & (g1953) & (!g1954) & (g1955) & (!g1956)) + ((g1951) & (!g1952) & (g1953) & (!g1954) & (g1955) & (g1956)) + ((g1951) & (!g1952) & (g1953) & (g1954) & (!g1955) & (g1956)) + ((g1951) & (!g1952) & (g1953) & (g1954) & (g1955) & (!g1956)) + ((g1951) & (!g1952) & (g1953) & (g1954) & (g1955) & (g1956)) + ((g1951) & (g1952) & (!g1953) & (!g1954) & (g1955) & (g1956)) + ((g1951) & (g1952) & (!g1953) & (g1954) & (!g1955) & (g1956)) + ((g1951) & (g1952) & (!g1953) & (g1954) & (g1955) & (!g1956)) + ((g1951) & (g1952) & (!g1953) & (g1954) & (g1955) & (g1956)) + ((g1951) & (g1952) & (g1953) & (!g1954) & (!g1955) & (g1956)) + ((g1951) & (g1952) & (g1953) & (!g1954) & (g1955) & (!g1956)) + ((g1951) & (g1952) & (g1953) & (!g1954) & (g1955) & (g1956)) + ((g1951) & (g1952) & (g1953) & (g1954) & (!g1955) & (g1956)) + ((g1951) & (g1952) & (g1953) & (g1954) & (g1955) & (!g1956)) + ((g1951) & (g1952) & (g1953) & (g1954) & (g1955) & (g1956)));
	assign g7825 = (((!g3429) & (g3957) & (!g1958)) + ((!g3429) & (g3957) & (g1958)) + ((g3429) & (!g3957) & (g1958)) + ((g3429) & (g3957) & (g1958)));
	assign g7826 = (((!g3464) & (g3961) & (!g1959)) + ((!g3464) & (g3961) & (g1959)) + ((g3464) & (!g3961) & (g1959)) + ((g3464) & (g3961) & (g1959)));
	assign g7827 = (((!g3429) & (g3963) & (!g1960)) + ((!g3429) & (g3963) & (g1960)) + ((g3429) & (!g3963) & (g1960)) + ((g3429) & (g3963) & (g1960)));
	assign g7828 = (((!g3464) & (g3967) & (!g1961)) + ((!g3464) & (g3967) & (g1961)) + ((g3464) & (!g3967) & (g1961)) + ((g3464) & (g3967) & (g1961)));
	assign g7829 = (((!g3429) & (g3970) & (!g1962)) + ((!g3429) & (g3970) & (g1962)) + ((g3429) & (!g3970) & (g1962)) + ((g3429) & (g3970) & (g1962)));
	assign g7830 = (((!g3464) & (g3973) & (!g1963)) + ((!g3464) & (g3973) & (g1963)) + ((g3464) & (!g3973) & (g1963)) + ((g3464) & (g3973) & (g1963)));
	assign g1964 = (((!g1962) & (g1963)) + ((g1962) & (!g1963)));
	assign g1965 = (((!g1957) & (!g1958) & (!g1959) & (g1960) & (g1961) & (g1964)) + ((!g1957) & (!g1958) & (g1959) & (g1960) & (g1961) & (g1964)) + ((!g1957) & (g1958) & (!g1959) & (g1960) & (g1961) & (g1964)) + ((!g1957) & (g1958) & (g1959) & (!g1960) & (g1961) & (g1964)) + ((!g1957) & (g1958) & (g1959) & (g1960) & (!g1961) & (g1964)) + ((!g1957) & (g1958) & (g1959) & (g1960) & (g1961) & (g1964)) + ((g1957) & (!g1958) & (!g1959) & (g1960) & (g1961) & (g1964)) + ((g1957) & (!g1958) & (g1959) & (!g1960) & (g1961) & (g1964)) + ((g1957) & (!g1958) & (g1959) & (g1960) & (!g1961) & (g1964)) + ((g1957) & (!g1958) & (g1959) & (g1960) & (g1961) & (g1964)) + ((g1957) & (g1958) & (!g1959) & (!g1960) & (g1961) & (g1964)) + ((g1957) & (g1958) & (!g1959) & (g1960) & (!g1961) & (g1964)) + ((g1957) & (g1958) & (!g1959) & (g1960) & (g1961) & (g1964)) + ((g1957) & (g1958) & (g1959) & (!g1960) & (g1961) & (g1964)) + ((g1957) & (g1958) & (g1959) & (g1960) & (!g1961) & (g1964)) + ((g1957) & (g1958) & (g1959) & (g1960) & (g1961) & (g1964)));
	assign g1966 = (((g1962) & (g1963)));
	assign g7831 = (((!g3429) & (g3978) & (!g1967)) + ((!g3429) & (g3978) & (g1967)) + ((g3429) & (!g3978) & (g1967)) + ((g3429) & (g3978) & (g1967)));
	assign g7832 = (((!g3464) & (g3981) & (!g1968)) + ((!g3464) & (g3981) & (g1968)) + ((g3464) & (!g3981) & (g1968)) + ((g3464) & (g3981) & (g1968)));
	assign g7833 = (((!g3429) & (g3984) & (!g1969)) + ((!g3429) & (g3984) & (g1969)) + ((g3429) & (!g3984) & (g1969)) + ((g3429) & (g3984) & (g1969)));
	assign g7834 = (((!g3464) & (g6961) & (!g1970)) + ((!g3464) & (g6961) & (g1970)) + ((g3464) & (!g6961) & (g1970)) + ((g3464) & (g6961) & (g1970)));
	assign g1971 = (((!g1965) & (!g1966) & (!g1967) & (!g1968) & (g1969) & (g1970)) + ((!g1965) & (!g1966) & (!g1967) & (g1968) & (g1969) & (g1970)) + ((!g1965) & (!g1966) & (g1967) & (!g1968) & (g1969) & (g1970)) + ((!g1965) & (!g1966) & (g1967) & (g1968) & (!g1969) & (g1970)) + ((!g1965) & (!g1966) & (g1967) & (g1968) & (g1969) & (!g1970)) + ((!g1965) & (!g1966) & (g1967) & (g1968) & (g1969) & (g1970)) + ((!g1965) & (g1966) & (!g1967) & (!g1968) & (g1969) & (g1970)) + ((!g1965) & (g1966) & (!g1967) & (g1968) & (!g1969) & (g1970)) + ((!g1965) & (g1966) & (!g1967) & (g1968) & (g1969) & (!g1970)) + ((!g1965) & (g1966) & (!g1967) & (g1968) & (g1969) & (g1970)) + ((!g1965) & (g1966) & (g1967) & (!g1968) & (!g1969) & (g1970)) + ((!g1965) & (g1966) & (g1967) & (!g1968) & (g1969) & (!g1970)) + ((!g1965) & (g1966) & (g1967) & (!g1968) & (g1969) & (g1970)) + ((!g1965) & (g1966) & (g1967) & (g1968) & (!g1969) & (g1970)) + ((!g1965) & (g1966) & (g1967) & (g1968) & (g1969) & (!g1970)) + ((!g1965) & (g1966) & (g1967) & (g1968) & (g1969) & (g1970)) + ((g1965) & (!g1966) & (!g1967) & (!g1968) & (g1969) & (g1970)) + ((g1965) & (!g1966) & (!g1967) & (g1968) & (!g1969) & (g1970)) + ((g1965) & (!g1966) & (!g1967) & (g1968) & (g1969) & (!g1970)) + ((g1965) & (!g1966) & (!g1967) & (g1968) & (g1969) & (g1970)) + ((g1965) & (!g1966) & (g1967) & (!g1968) & (!g1969) & (g1970)) + ((g1965) & (!g1966) & (g1967) & (!g1968) & (g1969) & (!g1970)) + ((g1965) & (!g1966) & (g1967) & (!g1968) & (g1969) & (g1970)) + ((g1965) & (!g1966) & (g1967) & (g1968) & (!g1969) & (g1970)) + ((g1965) & (!g1966) & (g1967) & (g1968) & (g1969) & (!g1970)) + ((g1965) & (!g1966) & (g1967) & (g1968) & (g1969) & (g1970)) + ((g1965) & (g1966) & (!g1967) & (!g1968) & (g1969) & (g1970)) + ((g1965) & (g1966) & (!g1967) & (g1968) & (!g1969) & (g1970)) + ((g1965) & (g1966) & (!g1967) & (g1968) & (g1969) & (!g1970)) + ((g1965) & (g1966) & (!g1967) & (g1968) & (g1969) & (g1970)) + ((g1965) & (g1966) & (g1967) & (!g1968) & (!g1969) & (g1970)) + ((g1965) & (g1966) & (g1967) & (!g1968) & (g1969) & (!g1970)) + ((g1965) & (g1966) & (g1967) & (!g1968) & (g1969) & (g1970)) + ((g1965) & (g1966) & (g1967) & (g1968) & (!g1969) & (g1970)) + ((g1965) & (g1966) & (g1967) & (g1968) & (g1969) & (!g1970)) + ((g1965) & (g1966) & (g1967) & (g1968) & (g1969) & (g1970)));
	assign g7835 = (((!g3429) & (g3989) & (!g1972)) + ((!g3429) & (g3989) & (g1972)) + ((g3429) & (!g3989) & (g1972)) + ((g3429) & (g3989) & (g1972)));
	assign g7836 = (((!g3464) & (g3992) & (!g1973)) + ((!g3464) & (g3992) & (g1973)) + ((g3464) & (!g3992) & (g1973)) + ((g3464) & (g3992) & (g1973)));
	assign g1974 = (((!g1971) & (g1972) & (g1973)) + ((g1971) & (!g1972) & (g1973)) + ((g1971) & (g1972) & (!g1973)) + ((g1971) & (g1972) & (g1973)));
	assign g7837 = (((!g3429) & (g3995) & (!g1975)) + ((!g3429) & (g3995) & (g1975)) + ((g3429) & (!g3995) & (g1975)) + ((g3429) & (g3995) & (g1975)));
	assign g7838 = (((!g3464) & (g3997) & (!g1976)) + ((!g3464) & (g3997) & (g1976)) + ((g3464) & (!g3997) & (g1976)) + ((g3464) & (g3997) & (g1976)));
	assign g7839 = (((!g3429) & (g4001) & (!g1977)) + ((!g3429) & (g4001) & (g1977)) + ((g3429) & (!g4001) & (g1977)) + ((g3429) & (g4001) & (g1977)));
	assign g7840 = (((!g3499) & (g4007) & (!g1978)) + ((!g3499) & (g4007) & (g1978)) + ((g3499) & (!g4007) & (g1978)) + ((g3499) & (g4007) & (g1978)));
	assign g7841 = (((!g3429) & (g4011) & (!g1979)) + ((!g3429) & (g4011) & (g1979)) + ((g3429) & (!g4011) & (g1979)) + ((g3429) & (g4011) & (g1979)));
	assign g7842 = (((!g3499) & (g4018) & (!g1980)) + ((!g3499) & (g4018) & (g1980)) + ((g3499) & (!g4018) & (g1980)) + ((g3499) & (g4018) & (g1980)));
	assign g1981 = (((!g1884) & (!g1888) & (!g1977) & (!g1978) & (g1979) & (g1980)) + ((!g1884) & (!g1888) & (!g1977) & (g1978) & (g1979) & (g1980)) + ((!g1884) & (!g1888) & (g1977) & (!g1978) & (g1979) & (g1980)) + ((!g1884) & (!g1888) & (g1977) & (g1978) & (!g1979) & (g1980)) + ((!g1884) & (!g1888) & (g1977) & (g1978) & (g1979) & (!g1980)) + ((!g1884) & (!g1888) & (g1977) & (g1978) & (g1979) & (g1980)) + ((!g1884) & (g1888) & (!g1977) & (!g1978) & (g1979) & (g1980)) + ((!g1884) & (g1888) & (!g1977) & (g1978) & (g1979) & (g1980)) + ((!g1884) & (g1888) & (g1977) & (!g1978) & (g1979) & (g1980)) + ((!g1884) & (g1888) & (g1977) & (g1978) & (!g1979) & (g1980)) + ((!g1884) & (g1888) & (g1977) & (g1978) & (g1979) & (!g1980)) + ((!g1884) & (g1888) & (g1977) & (g1978) & (g1979) & (g1980)) + ((g1884) & (!g1888) & (!g1977) & (!g1978) & (g1979) & (g1980)) + ((g1884) & (!g1888) & (!g1977) & (g1978) & (g1979) & (g1980)) + ((g1884) & (!g1888) & (g1977) & (!g1978) & (g1979) & (g1980)) + ((g1884) & (!g1888) & (g1977) & (g1978) & (!g1979) & (g1980)) + ((g1884) & (!g1888) & (g1977) & (g1978) & (g1979) & (!g1980)) + ((g1884) & (!g1888) & (g1977) & (g1978) & (g1979) & (g1980)) + ((g1884) & (g1888) & (!g1977) & (!g1978) & (g1979) & (g1980)) + ((g1884) & (g1888) & (!g1977) & (g1978) & (!g1979) & (g1980)) + ((g1884) & (g1888) & (!g1977) & (g1978) & (g1979) & (!g1980)) + ((g1884) & (g1888) & (!g1977) & (g1978) & (g1979) & (g1980)) + ((g1884) & (g1888) & (g1977) & (!g1978) & (!g1979) & (g1980)) + ((g1884) & (g1888) & (g1977) & (!g1978) & (g1979) & (!g1980)) + ((g1884) & (g1888) & (g1977) & (!g1978) & (g1979) & (g1980)) + ((g1884) & (g1888) & (g1977) & (g1978) & (!g1979) & (g1980)) + ((g1884) & (g1888) & (g1977) & (g1978) & (g1979) & (!g1980)) + ((g1884) & (g1888) & (g1977) & (g1978) & (g1979) & (g1980)));
	assign g7843 = (((!g3429) & (g4028) & (!g1982)) + ((!g3429) & (g4028) & (g1982)) + ((g3429) & (!g4028) & (g1982)) + ((g3429) & (g4028) & (g1982)));
	assign g7844 = (((!g3499) & (g4032) & (!g1983)) + ((!g3499) & (g4032) & (g1983)) + ((g3499) & (!g4032) & (g1983)) + ((g3499) & (g4032) & (g1983)));
	assign g7845 = (((!g3429) & (g4037) & (!g1984)) + ((!g3429) & (g4037) & (g1984)) + ((g3429) & (!g4037) & (g1984)) + ((g3429) & (g4037) & (g1984)));
	assign g7846 = (((!g3499) & (g4041) & (!g1985)) + ((!g3499) & (g4041) & (g1985)) + ((g3499) & (!g4041) & (g1985)) + ((g3499) & (g4041) & (g1985)));
	assign g7847 = (((!g3429) & (g4047) & (!g1986)) + ((!g3429) & (g4047) & (g1986)) + ((g3429) & (!g4047) & (g1986)) + ((g3429) & (g4047) & (g1986)));
	assign g7848 = (((!g3499) & (g4050) & (!g1987)) + ((!g3499) & (g4050) & (g1987)) + ((g3499) & (!g4050) & (g1987)) + ((g3499) & (g4050) & (g1987)));
	assign g1988 = (((!g1986) & (g1987)) + ((g1986) & (!g1987)));
	assign g1989 = (((!g1981) & (!g1982) & (!g1983) & (g1984) & (g1985) & (g1988)) + ((!g1981) & (!g1982) & (g1983) & (g1984) & (g1985) & (g1988)) + ((!g1981) & (g1982) & (!g1983) & (g1984) & (g1985) & (g1988)) + ((!g1981) & (g1982) & (g1983) & (!g1984) & (g1985) & (g1988)) + ((!g1981) & (g1982) & (g1983) & (g1984) & (!g1985) & (g1988)) + ((!g1981) & (g1982) & (g1983) & (g1984) & (g1985) & (g1988)) + ((g1981) & (!g1982) & (!g1983) & (g1984) & (g1985) & (g1988)) + ((g1981) & (!g1982) & (g1983) & (!g1984) & (g1985) & (g1988)) + ((g1981) & (!g1982) & (g1983) & (g1984) & (!g1985) & (g1988)) + ((g1981) & (!g1982) & (g1983) & (g1984) & (g1985) & (g1988)) + ((g1981) & (g1982) & (!g1983) & (!g1984) & (g1985) & (g1988)) + ((g1981) & (g1982) & (!g1983) & (g1984) & (!g1985) & (g1988)) + ((g1981) & (g1982) & (!g1983) & (g1984) & (g1985) & (g1988)) + ((g1981) & (g1982) & (g1983) & (!g1984) & (g1985) & (g1988)) + ((g1981) & (g1982) & (g1983) & (g1984) & (!g1985) & (g1988)) + ((g1981) & (g1982) & (g1983) & (g1984) & (g1985) & (g1988)));
	assign g1990 = (((g1986) & (g1987)));
	assign g7849 = (((!g3429) & (g4054) & (!g1991)) + ((!g3429) & (g4054) & (g1991)) + ((g3429) & (!g4054) & (g1991)) + ((g3429) & (g4054) & (g1991)));
	assign g7850 = (((!g3499) & (g4057) & (!g1992)) + ((!g3499) & (g4057) & (g1992)) + ((g3499) & (!g4057) & (g1992)) + ((g3499) & (g4057) & (g1992)));
	assign g7851 = (((!g3429) & (g4061) & (!g1993)) + ((!g3429) & (g4061) & (g1993)) + ((g3429) & (!g4061) & (g1993)) + ((g3429) & (g4061) & (g1993)));
	assign g7852 = (((!g3499) & (g6926) & (!g1994)) + ((!g3499) & (g6926) & (g1994)) + ((g3499) & (!g6926) & (g1994)) + ((g3499) & (g6926) & (g1994)));
	assign g1995 = (((!g1989) & (!g1990) & (!g1991) & (!g1992) & (!g1993) & (!g1994)) + ((!g1989) & (!g1990) & (!g1991) & (!g1992) & (!g1993) & (g1994)) + ((!g1989) & (!g1990) & (!g1991) & (!g1992) & (g1993) & (!g1994)) + ((!g1989) & (!g1990) & (!g1991) & (g1992) & (!g1993) & (!g1994)) + ((!g1989) & (!g1990) & (!g1991) & (g1992) & (!g1993) & (g1994)) + ((!g1989) & (!g1990) & (!g1991) & (g1992) & (g1993) & (!g1994)) + ((!g1989) & (!g1990) & (g1991) & (!g1992) & (!g1993) & (!g1994)) + ((!g1989) & (!g1990) & (g1991) & (!g1992) & (!g1993) & (g1994)) + ((!g1989) & (!g1990) & (g1991) & (!g1992) & (g1993) & (!g1994)) + ((!g1989) & (!g1990) & (g1991) & (g1992) & (!g1993) & (!g1994)) + ((!g1989) & (g1990) & (!g1991) & (!g1992) & (!g1993) & (!g1994)) + ((!g1989) & (g1990) & (!g1991) & (!g1992) & (!g1993) & (g1994)) + ((!g1989) & (g1990) & (!g1991) & (!g1992) & (g1993) & (!g1994)) + ((!g1989) & (g1990) & (!g1991) & (g1992) & (!g1993) & (!g1994)) + ((!g1989) & (g1990) & (g1991) & (!g1992) & (!g1993) & (!g1994)) + ((!g1989) & (g1990) & (g1991) & (g1992) & (!g1993) & (!g1994)) + ((g1989) & (!g1990) & (!g1991) & (!g1992) & (!g1993) & (!g1994)) + ((g1989) & (!g1990) & (!g1991) & (!g1992) & (!g1993) & (g1994)) + ((g1989) & (!g1990) & (!g1991) & (!g1992) & (g1993) & (!g1994)) + ((g1989) & (!g1990) & (!g1991) & (g1992) & (!g1993) & (!g1994)) + ((g1989) & (!g1990) & (g1991) & (!g1992) & (!g1993) & (!g1994)) + ((g1989) & (!g1990) & (g1991) & (g1992) & (!g1993) & (!g1994)) + ((g1989) & (g1990) & (!g1991) & (!g1992) & (!g1993) & (!g1994)) + ((g1989) & (g1990) & (!g1991) & (!g1992) & (!g1993) & (g1994)) + ((g1989) & (g1990) & (!g1991) & (!g1992) & (g1993) & (!g1994)) + ((g1989) & (g1990) & (!g1991) & (g1992) & (!g1993) & (!g1994)) + ((g1989) & (g1990) & (g1991) & (!g1992) & (!g1993) & (!g1994)) + ((g1989) & (g1990) & (g1991) & (g1992) & (!g1993) & (!g1994)));
	assign g7853 = (((!g3429) & (g4069) & (!g1996)) + ((!g3429) & (g4069) & (g1996)) + ((g3429) & (!g4069) & (g1996)) + ((g3429) & (g4069) & (g1996)));
	assign g7854 = (((!g3499) & (g4073) & (!g1997)) + ((!g3499) & (g4073) & (g1997)) + ((g3499) & (!g4073) & (g1997)) + ((g3499) & (g4073) & (g1997)));
	assign g7855 = (((!g3429) & (g4076) & (!g1998)) + ((!g3429) & (g4076) & (g1998)) + ((g3429) & (!g4076) & (g1998)) + ((g3429) & (g4076) & (g1998)));
	assign g7856 = (((!g3499) & (g4080) & (!g1999)) + ((!g3499) & (g4080) & (g1999)) + ((g3499) & (!g4080) & (g1999)) + ((g3499) & (g4080) & (g1999)));
	assign g2000 = (((!g1995) & (!g1996) & (!g1997) & (g1998) & (g1999)) + ((!g1995) & (!g1996) & (g1997) & (!g1998) & (g1999)) + ((!g1995) & (!g1996) & (g1997) & (g1998) & (!g1999)) + ((!g1995) & (!g1996) & (g1997) & (g1998) & (g1999)) + ((!g1995) & (g1996) & (!g1997) & (!g1998) & (g1999)) + ((!g1995) & (g1996) & (!g1997) & (g1998) & (!g1999)) + ((!g1995) & (g1996) & (!g1997) & (g1998) & (g1999)) + ((!g1995) & (g1996) & (g1997) & (!g1998) & (g1999)) + ((!g1995) & (g1996) & (g1997) & (g1998) & (!g1999)) + ((!g1995) & (g1996) & (g1997) & (g1998) & (g1999)) + ((g1995) & (!g1996) & (!g1997) & (g1998) & (g1999)) + ((g1995) & (!g1996) & (g1997) & (g1998) & (g1999)) + ((g1995) & (g1996) & (!g1997) & (g1998) & (g1999)) + ((g1995) & (g1996) & (g1997) & (!g1998) & (g1999)) + ((g1995) & (g1996) & (g1997) & (g1998) & (!g1999)) + ((g1995) & (g1996) & (g1997) & (g1998) & (g1999)));
	assign g7857 = (((!g3429) & (g4084) & (!g2001)) + ((!g3429) & (g4084) & (g2001)) + ((g3429) & (!g4084) & (g2001)) + ((g3429) & (g4084) & (g2001)));
	assign g7858 = (((!g3499) & (g4087) & (!g2002)) + ((!g3499) & (g4087) & (g2002)) + ((g3499) & (!g4087) & (g2002)) + ((g3499) & (g4087) & (g2002)));
	assign g7859 = (((!g3429) & (g4092) & (!g2003)) + ((!g3429) & (g4092) & (g2003)) + ((g3429) & (!g4092) & (g2003)) + ((g3429) & (g4092) & (g2003)));
	assign g7860 = (((!g3499) & (g4095) & (!g2004)) + ((!g3499) & (g4095) & (g2004)) + ((g3499) & (!g4095) & (g2004)) + ((g3499) & (g4095) & (g2004)));
	assign g7861 = (((!g3429) & (g4099) & (!g2005)) + ((!g3429) & (g4099) & (g2005)) + ((g3429) & (!g4099) & (g2005)) + ((g3429) & (g4099) & (g2005)));
	assign g7862 = (((!g3499) & (g6916) & (!g2006)) + ((!g3499) & (g6916) & (g2006)) + ((g3499) & (!g6916) & (g2006)) + ((g3499) & (g6916) & (g2006)));
	assign g2007 = (((!g2005) & (g2006)) + ((g2005) & (!g2006)));
	assign g2008 = (((!g2000) & (!g2001) & (!g2002) & (g2003) & (g2004) & (g2007)) + ((!g2000) & (!g2001) & (g2002) & (g2003) & (g2004) & (g2007)) + ((!g2000) & (g2001) & (!g2002) & (g2003) & (g2004) & (g2007)) + ((!g2000) & (g2001) & (g2002) & (!g2003) & (g2004) & (g2007)) + ((!g2000) & (g2001) & (g2002) & (g2003) & (!g2004) & (g2007)) + ((!g2000) & (g2001) & (g2002) & (g2003) & (g2004) & (g2007)) + ((g2000) & (!g2001) & (!g2002) & (g2003) & (g2004) & (g2007)) + ((g2000) & (!g2001) & (g2002) & (!g2003) & (g2004) & (g2007)) + ((g2000) & (!g2001) & (g2002) & (g2003) & (!g2004) & (g2007)) + ((g2000) & (!g2001) & (g2002) & (g2003) & (g2004) & (g2007)) + ((g2000) & (g2001) & (!g2002) & (!g2003) & (g2004) & (g2007)) + ((g2000) & (g2001) & (!g2002) & (g2003) & (!g2004) & (g2007)) + ((g2000) & (g2001) & (!g2002) & (g2003) & (g2004) & (g2007)) + ((g2000) & (g2001) & (g2002) & (!g2003) & (g2004) & (g2007)) + ((g2000) & (g2001) & (g2002) & (g2003) & (!g2004) & (g2007)) + ((g2000) & (g2001) & (g2002) & (g2003) & (g2004) & (g2007)));
	assign g2009 = (((g2005) & (g2006)));
	assign g2010 = (((!g2008) & (!g2009)));
	assign g7863 = (((!g3429) & (g4105) & (!g2011)) + ((!g3429) & (g4105) & (g2011)) + ((g3429) & (!g4105) & (g2011)) + ((g3429) & (g4105) & (g2011)));
	assign g7864 = (((!g3499) & (g4108) & (!g2012)) + ((!g3499) & (g4108) & (g2012)) + ((g3499) & (!g4108) & (g2012)) + ((g3499) & (g4108) & (g2012)));
	assign g7865 = (((!g3429) & (g4111) & (!g2013)) + ((!g3429) & (g4111) & (g2013)) + ((g3429) & (!g4111) & (g2013)) + ((g3429) & (g4111) & (g2013)));
	assign g7866 = (((!g3499) & (g4113) & (!g2014)) + ((!g3499) & (g4113) & (g2014)) + ((g3499) & (!g4113) & (g2014)) + ((g3499) & (g4113) & (g2014)));
	assign g2015 = (((!g2010) & (!g2011) & (!g2012) & (!g2013) & (g2014)) + ((!g2010) & (!g2011) & (!g2012) & (g2013) & (!g2014)) + ((!g2010) & (!g2011) & (g2012) & (!g2013) & (!g2014)) + ((!g2010) & (!g2011) & (g2012) & (g2013) & (g2014)) + ((!g2010) & (g2011) & (!g2012) & (!g2013) & (!g2014)) + ((!g2010) & (g2011) & (!g2012) & (g2013) & (g2014)) + ((!g2010) & (g2011) & (g2012) & (!g2013) & (!g2014)) + ((!g2010) & (g2011) & (g2012) & (g2013) & (g2014)) + ((g2010) & (!g2011) & (!g2012) & (!g2013) & (g2014)) + ((g2010) & (!g2011) & (!g2012) & (g2013) & (!g2014)) + ((g2010) & (!g2011) & (g2012) & (!g2013) & (g2014)) + ((g2010) & (!g2011) & (g2012) & (g2013) & (!g2014)) + ((g2010) & (g2011) & (!g2012) & (!g2013) & (g2014)) + ((g2010) & (g2011) & (!g2012) & (g2013) & (!g2014)) + ((g2010) & (g2011) & (g2012) & (!g2013) & (!g2014)) + ((g2010) & (g2011) & (g2012) & (g2013) & (g2014)));
	assign g2016 = (((!g827) & (g831)));
	assign g2017 = (((!reset) & (!g830) & (!g1921) & (!g1922) & (!g2016)) + ((!reset) & (!g830) & (!g1921) & (g1922) & (!g2016)) + ((!reset) & (!g830) & (g1921) & (!g1922) & (!g2016)) + ((!reset) & (!g830) & (g1921) & (g1922) & (!g2016)) + ((!reset) & (g830) & (!g1921) & (!g1922) & (!g2016)) + ((!reset) & (g830) & (!g1921) & (!g1922) & (g2016)) + ((!reset) & (g830) & (!g1921) & (g1922) & (!g2016)) + ((!reset) & (g830) & (!g1921) & (g1922) & (g2016)) + ((!reset) & (g830) & (g1921) & (!g1922) & (!g2016)) + ((!reset) & (g830) & (g1921) & (!g1922) & (g2016)) + ((!reset) & (g830) & (g1921) & (g1922) & (!g2016)) + ((reset) & (!g830) & (!g1921) & (!g1922) & (!g2016)) + ((reset) & (!g830) & (!g1921) & (!g1922) & (g2016)) + ((reset) & (!g830) & (!g1921) & (g1922) & (!g2016)) + ((reset) & (!g830) & (!g1921) & (g1922) & (g2016)) + ((reset) & (!g830) & (g1921) & (!g1922) & (!g2016)) + ((reset) & (!g830) & (g1921) & (!g1922) & (g2016)) + ((reset) & (!g830) & (g1921) & (g1922) & (!g2016)) + ((reset) & (!g830) & (g1921) & (g1922) & (g2016)) + ((reset) & (g830) & (!g1921) & (!g1922) & (!g2016)) + ((reset) & (g830) & (!g1921) & (!g1922) & (g2016)) + ((reset) & (g830) & (!g1921) & (g1922) & (!g2016)) + ((reset) & (g830) & (!g1921) & (g1922) & (g2016)) + ((reset) & (g830) & (g1921) & (!g1922) & (!g2016)) + ((reset) & (g830) & (g1921) & (!g1922) & (g2016)) + ((reset) & (g830) & (g1921) & (g1922) & (!g2016)) + ((reset) & (g830) & (g1921) & (g1922) & (g2016)));
	assign g2018 = (((!reset) & (!g830) & (g2016) & (!g1923) & (!g1934)) + ((!reset) & (!g830) & (g2016) & (!g1923) & (g1934)) + ((!reset) & (!g830) & (g2016) & (g1923) & (!g1934)) + ((!reset) & (!g830) & (g2016) & (g1923) & (g1934)) + ((!reset) & (g830) & (!g2016) & (!g1923) & (!g1934)) + ((!reset) & (g830) & (!g2016) & (!g1923) & (g1934)) + ((!reset) & (g830) & (!g2016) & (g1923) & (!g1934)) + ((!reset) & (g830) & (!g2016) & (g1923) & (g1934)) + ((!reset) & (g830) & (g2016) & (!g1923) & (!g1934)) + ((!reset) & (g830) & (g2016) & (!g1923) & (g1934)) + ((!reset) & (g830) & (g2016) & (g1923) & (!g1934)));
	assign g2019 = (((g1923) & (g1934)));
	assign g2020 = (((!reset) & (!g827) & (!g830) & (!g831) & (!g2019) & (!g1936)) + ((!reset) & (!g827) & (!g830) & (!g831) & (g2019) & (!g1936)) + ((!reset) & (!g827) & (!g830) & (g831) & (!g2019) & (g1936)) + ((!reset) & (!g827) & (!g830) & (g831) & (g2019) & (g1936)) + ((!reset) & (!g827) & (g830) & (!g831) & (!g2019) & (!g1936)) + ((!reset) & (!g827) & (g830) & (!g831) & (!g2019) & (g1936)) + ((!reset) & (!g827) & (g830) & (!g831) & (g2019) & (!g1936)) + ((!reset) & (!g827) & (g830) & (!g831) & (g2019) & (g1936)) + ((!reset) & (!g827) & (g830) & (g831) & (!g2019) & (!g1936)) + ((!reset) & (!g827) & (g830) & (g831) & (!g2019) & (g1936)) + ((!reset) & (g827) & (!g830) & (!g831) & (!g2019) & (!g1936)) + ((!reset) & (g827) & (!g830) & (!g831) & (g2019) & (!g1936)) + ((!reset) & (g827) & (!g830) & (g831) & (!g2019) & (!g1936)) + ((!reset) & (g827) & (!g830) & (g831) & (!g2019) & (g1936)) + ((!reset) & (g827) & (!g830) & (g831) & (g2019) & (!g1936)) + ((!reset) & (g827) & (!g830) & (g831) & (g2019) & (g1936)) + ((!reset) & (g827) & (g830) & (g831) & (!g2019) & (!g1936)) + ((!reset) & (g827) & (g830) & (g831) & (!g2019) & (g1936)) + ((!reset) & (g827) & (g830) & (g831) & (g2019) & (!g1936)) + ((!reset) & (g827) & (g830) & (g831) & (g2019) & (g1936)));
	assign g2021 = (((!g800) & (!g827) & (!g834) & (!g1890) & (g1939)) + ((!g800) & (!g827) & (!g834) & (g1890) & (g1939)) + ((!g800) & (!g827) & (g834) & (!g1890) & (g1939)) + ((!g800) & (!g827) & (g834) & (g1890) & (g1939)) + ((!g800) & (g827) & (!g834) & (!g1890) & (g1939)) + ((!g800) & (g827) & (!g834) & (g1890) & (g1939)) + ((!g800) & (g827) & (g834) & (!g1890) & (!g1939)) + ((!g800) & (g827) & (g834) & (g1890) & (!g1939)) + ((g800) & (!g827) & (!g834) & (!g1890) & (g1939)) + ((g800) & (!g827) & (!g834) & (g1890) & (g1939)) + ((g800) & (!g827) & (g834) & (!g1890) & (g1939)) + ((g800) & (!g827) & (g834) & (g1890) & (g1939)) + ((g800) & (g827) & (!g834) & (!g1890) & (g1939)) + ((g800) & (g827) & (!g834) & (g1890) & (!g1939)) + ((g800) & (g827) & (g834) & (!g1890) & (!g1939)) + ((g800) & (g827) & (g834) & (g1890) & (g1939)));
	assign g7867 = (((!g3499) & (g4119) & (!g2022)) + ((!g3499) & (g4119) & (g2022)) + ((g3499) & (!g4119) & (g2022)) + ((g3499) & (g4119) & (g2022)));
	assign g2023 = (((!g808) & (!g827) & (!g836) & (!g1898) & (g2022)) + ((!g808) & (!g827) & (!g836) & (g1898) & (g2022)) + ((!g808) & (!g827) & (g836) & (!g1898) & (g2022)) + ((!g808) & (!g827) & (g836) & (g1898) & (g2022)) + ((!g808) & (g827) & (!g836) & (!g1898) & (g2022)) + ((!g808) & (g827) & (!g836) & (g1898) & (g2022)) + ((!g808) & (g827) & (g836) & (!g1898) & (!g2022)) + ((!g808) & (g827) & (g836) & (g1898) & (!g2022)) + ((g808) & (!g827) & (!g836) & (!g1898) & (g2022)) + ((g808) & (!g827) & (!g836) & (g1898) & (g2022)) + ((g808) & (!g827) & (g836) & (!g1898) & (g2022)) + ((g808) & (!g827) & (g836) & (g1898) & (g2022)) + ((g808) & (g827) & (!g836) & (!g1898) & (g2022)) + ((g808) & (g827) & (!g836) & (g1898) & (!g2022)) + ((g808) & (g827) & (g836) & (!g1898) & (!g2022)) + ((g808) & (g827) & (g836) & (g1898) & (g2022)));
	assign g2024 = (((!g816) & (!g827) & (!g838) & (!g1906) & (g1940)) + ((!g816) & (!g827) & (!g838) & (g1906) & (g1940)) + ((!g816) & (!g827) & (g838) & (!g1906) & (g1940)) + ((!g816) & (!g827) & (g838) & (g1906) & (g1940)) + ((!g816) & (g827) & (!g838) & (!g1906) & (g1940)) + ((!g816) & (g827) & (!g838) & (g1906) & (g1940)) + ((!g816) & (g827) & (g838) & (!g1906) & (!g1940)) + ((!g816) & (g827) & (g838) & (g1906) & (!g1940)) + ((g816) & (!g827) & (!g838) & (!g1906) & (g1940)) + ((g816) & (!g827) & (!g838) & (g1906) & (g1940)) + ((g816) & (!g827) & (g838) & (!g1906) & (g1940)) + ((g816) & (!g827) & (g838) & (g1906) & (g1940)) + ((g816) & (g827) & (!g838) & (!g1906) & (g1940)) + ((g816) & (g827) & (!g838) & (g1906) & (!g1940)) + ((g816) & (g827) & (g838) & (!g1906) & (!g1940)) + ((g816) & (g827) & (g838) & (g1906) & (g1940)));
	assign g2025 = (((!g790) & (!g827) & (!g840) & (!g1884) & (g1977)) + ((!g790) & (!g827) & (!g840) & (g1884) & (g1977)) + ((!g790) & (!g827) & (g840) & (!g1884) & (g1977)) + ((!g790) & (!g827) & (g840) & (g1884) & (g1977)) + ((!g790) & (g827) & (!g840) & (!g1884) & (g1977)) + ((!g790) & (g827) & (!g840) & (g1884) & (g1977)) + ((!g790) & (g827) & (g840) & (!g1884) & (!g1977)) + ((!g790) & (g827) & (g840) & (g1884) & (!g1977)) + ((g790) & (!g827) & (!g840) & (!g1884) & (g1977)) + ((g790) & (!g827) & (!g840) & (g1884) & (g1977)) + ((g790) & (!g827) & (g840) & (!g1884) & (g1977)) + ((g790) & (!g827) & (g840) & (g1884) & (g1977)) + ((g790) & (g827) & (!g840) & (!g1884) & (g1977)) + ((g790) & (g827) & (!g840) & (g1884) & (!g1977)) + ((g790) & (g827) & (g840) & (!g1884) & (!g1977)) + ((g790) & (g827) & (g840) & (g1884) & (g1977)));
	assign g7868 = (((!g2017) & (g6887) & (!g2026)) + ((!g2017) & (g6887) & (g2026)) + ((g2017) & (!g6887) & (g2026)) + ((g2017) & (g6887) & (g2026)));
	assign g2027 = (((!g802) & (!g827) & (!g842) & (!g1892) & (g2026)) + ((!g802) & (!g827) & (!g842) & (g1892) & (g2026)) + ((!g802) & (!g827) & (g842) & (!g1892) & (g2026)) + ((!g802) & (!g827) & (g842) & (g1892) & (g2026)) + ((!g802) & (g827) & (!g842) & (!g1892) & (g2026)) + ((!g802) & (g827) & (!g842) & (g1892) & (g2026)) + ((!g802) & (g827) & (g842) & (!g1892) & (!g2026)) + ((!g802) & (g827) & (g842) & (g1892) & (!g2026)) + ((g802) & (!g827) & (!g842) & (!g1892) & (g2026)) + ((g802) & (!g827) & (!g842) & (g1892) & (g2026)) + ((g802) & (!g827) & (g842) & (!g1892) & (g2026)) + ((g802) & (!g827) & (g842) & (g1892) & (g2026)) + ((g802) & (g827) & (!g842) & (!g1892) & (g2026)) + ((g802) & (g827) & (!g842) & (g1892) & (!g2026)) + ((g802) & (g827) & (g842) & (!g1892) & (!g2026)) + ((g802) & (g827) & (g842) & (g1892) & (g2026)));
	assign g7869 = (((!g3464) & (g4128) & (!g2028)) + ((!g3464) & (g4128) & (g2028)) + ((g3464) & (!g4128) & (g2028)) + ((g3464) & (g4128) & (g2028)));
	assign g2029 = (((!g810) & (!g827) & (!g844) & (!g1900) & (g2028)) + ((!g810) & (!g827) & (!g844) & (g1900) & (g2028)) + ((!g810) & (!g827) & (g844) & (!g1900) & (g2028)) + ((!g810) & (!g827) & (g844) & (g1900) & (g2028)) + ((!g810) & (g827) & (!g844) & (!g1900) & (g2028)) + ((!g810) & (g827) & (!g844) & (g1900) & (g2028)) + ((!g810) & (g827) & (g844) & (!g1900) & (!g2028)) + ((!g810) & (g827) & (g844) & (g1900) & (!g2028)) + ((g810) & (!g827) & (!g844) & (!g1900) & (g2028)) + ((g810) & (!g827) & (!g844) & (g1900) & (g2028)) + ((g810) & (!g827) & (g844) & (!g1900) & (g2028)) + ((g810) & (!g827) & (g844) & (g1900) & (g2028)) + ((g810) & (g827) & (!g844) & (!g1900) & (g2028)) + ((g810) & (g827) & (!g844) & (g1900) & (!g2028)) + ((g810) & (g827) & (g844) & (!g1900) & (!g2028)) + ((g810) & (g827) & (g844) & (g1900) & (g2028)));
	assign g7870 = (((!g3499) & (g4134) & (!g2030)) + ((!g3499) & (g4134) & (g2030)) + ((g3499) & (!g4134) & (g2030)) + ((g3499) & (g4134) & (g2030)));
	assign g2031 = (((!g818) & (!g827) & (!g846) & (!g1908) & (g2030)) + ((!g818) & (!g827) & (!g846) & (g1908) & (g2030)) + ((!g818) & (!g827) & (g846) & (!g1908) & (g2030)) + ((!g818) & (!g827) & (g846) & (g1908) & (g2030)) + ((!g818) & (g827) & (!g846) & (!g1908) & (g2030)) + ((!g818) & (g827) & (!g846) & (g1908) & (g2030)) + ((!g818) & (g827) & (g846) & (!g1908) & (!g2030)) + ((!g818) & (g827) & (g846) & (g1908) & (!g2030)) + ((g818) & (!g827) & (!g846) & (!g1908) & (g2030)) + ((g818) & (!g827) & (!g846) & (g1908) & (g2030)) + ((g818) & (!g827) & (g846) & (!g1908) & (g2030)) + ((g818) & (!g827) & (g846) & (g1908) & (g2030)) + ((g818) & (g827) & (!g846) & (!g1908) & (g2030)) + ((g818) & (g827) & (!g846) & (g1908) & (!g2030)) + ((g818) & (g827) & (g846) & (!g1908) & (!g2030)) + ((g818) & (g827) & (g846) & (g1908) & (g2030)));
	assign g7871 = (((!g3464) & (g4140) & (!g2032)) + ((!g3464) & (g4140) & (g2032)) + ((g3464) & (!g4140) & (g2032)) + ((g3464) & (g4140) & (g2032)));
	assign g2033 = (((!g792) & (!g827) & (!g848) & (!g1886) & (g2032)) + ((!g792) & (!g827) & (!g848) & (g1886) & (g2032)) + ((!g792) & (!g827) & (g848) & (!g1886) & (g2032)) + ((!g792) & (!g827) & (g848) & (g1886) & (g2032)) + ((!g792) & (g827) & (!g848) & (!g1886) & (g2032)) + ((!g792) & (g827) & (!g848) & (g1886) & (g2032)) + ((!g792) & (g827) & (g848) & (!g1886) & (!g2032)) + ((!g792) & (g827) & (g848) & (g1886) & (!g2032)) + ((g792) & (!g827) & (!g848) & (!g1886) & (g2032)) + ((g792) & (!g827) & (!g848) & (g1886) & (g2032)) + ((g792) & (!g827) & (g848) & (!g1886) & (g2032)) + ((g792) & (!g827) & (g848) & (g1886) & (g2032)) + ((g792) & (g827) & (!g848) & (!g1886) & (g2032)) + ((g792) & (g827) & (!g848) & (g1886) & (!g2032)) + ((g792) & (g827) & (g848) & (!g1886) & (!g2032)) + ((g792) & (g827) & (g848) & (g1886) & (g2032)));
	assign g7872 = (((!g3499) & (g4146) & (!g2034)) + ((!g3499) & (g4146) & (g2034)) + ((g3499) & (!g4146) & (g2034)) + ((g3499) & (g4146) & (g2034)));
	assign g2035 = (((!g804) & (!g827) & (!g850) & (!g1894) & (g2034)) + ((!g804) & (!g827) & (!g850) & (g1894) & (g2034)) + ((!g804) & (!g827) & (g850) & (!g1894) & (g2034)) + ((!g804) & (!g827) & (g850) & (g1894) & (g2034)) + ((!g804) & (g827) & (!g850) & (!g1894) & (g2034)) + ((!g804) & (g827) & (!g850) & (g1894) & (g2034)) + ((!g804) & (g827) & (g850) & (!g1894) & (!g2034)) + ((!g804) & (g827) & (g850) & (g1894) & (!g2034)) + ((g804) & (!g827) & (!g850) & (!g1894) & (g2034)) + ((g804) & (!g827) & (!g850) & (g1894) & (g2034)) + ((g804) & (!g827) & (g850) & (!g1894) & (g2034)) + ((g804) & (!g827) & (g850) & (g1894) & (g2034)) + ((g804) & (g827) & (!g850) & (!g1894) & (g2034)) + ((g804) & (g827) & (!g850) & (g1894) & (!g2034)) + ((g804) & (g827) & (g850) & (!g1894) & (!g2034)) + ((g804) & (g827) & (g850) & (g1894) & (g2034)));
	assign g7873 = (((!g2017) & (g6880) & (!g2036)) + ((!g2017) & (g6880) & (g2036)) + ((g2017) & (!g6880) & (g2036)) + ((g2017) & (g6880) & (g2036)));
	assign g2037 = (((!g812) & (!g827) & (!g852) & (!g1902) & (g2036)) + ((!g812) & (!g827) & (!g852) & (g1902) & (g2036)) + ((!g812) & (!g827) & (g852) & (!g1902) & (g2036)) + ((!g812) & (!g827) & (g852) & (g1902) & (g2036)) + ((!g812) & (g827) & (!g852) & (!g1902) & (g2036)) + ((!g812) & (g827) & (!g852) & (g1902) & (g2036)) + ((!g812) & (g827) & (g852) & (!g1902) & (!g2036)) + ((!g812) & (g827) & (g852) & (g1902) & (!g2036)) + ((g812) & (!g827) & (!g852) & (!g1902) & (g2036)) + ((g812) & (!g827) & (!g852) & (g1902) & (g2036)) + ((g812) & (!g827) & (g852) & (!g1902) & (g2036)) + ((g812) & (!g827) & (g852) & (g1902) & (g2036)) + ((g812) & (g827) & (!g852) & (!g1902) & (g2036)) + ((g812) & (g827) & (!g852) & (g1902) & (!g2036)) + ((g812) & (g827) & (g852) & (!g1902) & (!g2036)) + ((g812) & (g827) & (g852) & (g1902) & (g2036)));
	assign g7874 = (((!g3429) & (g4153) & (!g2038)) + ((!g3429) & (g4153) & (g2038)) + ((g3429) & (!g4153) & (g2038)) + ((g3429) & (g4153) & (g2038)));
	assign g2039 = (((!g820) & (!g827) & (!g854) & (!g1910) & (g2038)) + ((!g820) & (!g827) & (!g854) & (g1910) & (g2038)) + ((!g820) & (!g827) & (g854) & (!g1910) & (g2038)) + ((!g820) & (!g827) & (g854) & (g1910) & (g2038)) + ((!g820) & (g827) & (!g854) & (!g1910) & (g2038)) + ((!g820) & (g827) & (!g854) & (g1910) & (g2038)) + ((!g820) & (g827) & (g854) & (!g1910) & (!g2038)) + ((!g820) & (g827) & (g854) & (g1910) & (!g2038)) + ((g820) & (!g827) & (!g854) & (!g1910) & (g2038)) + ((g820) & (!g827) & (!g854) & (g1910) & (g2038)) + ((g820) & (!g827) & (g854) & (!g1910) & (g2038)) + ((g820) & (!g827) & (g854) & (g1910) & (g2038)) + ((g820) & (g827) & (!g854) & (!g1910) & (g2038)) + ((g820) & (g827) & (!g854) & (g1910) & (!g2038)) + ((g820) & (g827) & (g854) & (!g1910) & (!g2038)) + ((g820) & (g827) & (g854) & (g1910) & (g2038)));
	assign g2040 = (((!g794) & (!g827) & (!g856) & (!g1888) & (g1978)) + ((!g794) & (!g827) & (!g856) & (g1888) & (g1978)) + ((!g794) & (!g827) & (g856) & (!g1888) & (g1978)) + ((!g794) & (!g827) & (g856) & (g1888) & (g1978)) + ((!g794) & (g827) & (!g856) & (!g1888) & (g1978)) + ((!g794) & (g827) & (!g856) & (g1888) & (g1978)) + ((!g794) & (g827) & (g856) & (!g1888) & (!g1978)) + ((!g794) & (g827) & (g856) & (g1888) & (!g1978)) + ((g794) & (!g827) & (!g856) & (!g1888) & (g1978)) + ((g794) & (!g827) & (!g856) & (g1888) & (g1978)) + ((g794) & (!g827) & (g856) & (!g1888) & (g1978)) + ((g794) & (!g827) & (g856) & (g1888) & (g1978)) + ((g794) & (g827) & (!g856) & (!g1888) & (g1978)) + ((g794) & (g827) & (!g856) & (g1888) & (!g1978)) + ((g794) & (g827) & (g856) & (!g1888) & (!g1978)) + ((g794) & (g827) & (g856) & (g1888) & (g1978)));
	assign g7875 = (((!g3464) & (g4159) & (!g2041)) + ((!g3464) & (g4159) & (g2041)) + ((g3464) & (!g4159) & (g2041)) + ((g3464) & (g4159) & (g2041)));
	assign g2042 = (((!g806) & (!g827) & (!g858) & (!g1896) & (g2041)) + ((!g806) & (!g827) & (!g858) & (g1896) & (g2041)) + ((!g806) & (!g827) & (g858) & (!g1896) & (g2041)) + ((!g806) & (!g827) & (g858) & (g1896) & (g2041)) + ((!g806) & (g827) & (!g858) & (!g1896) & (g2041)) + ((!g806) & (g827) & (!g858) & (g1896) & (g2041)) + ((!g806) & (g827) & (g858) & (!g1896) & (!g2041)) + ((!g806) & (g827) & (g858) & (g1896) & (!g2041)) + ((g806) & (!g827) & (!g858) & (!g1896) & (g2041)) + ((g806) & (!g827) & (!g858) & (g1896) & (g2041)) + ((g806) & (!g827) & (g858) & (!g1896) & (g2041)) + ((g806) & (!g827) & (g858) & (g1896) & (g2041)) + ((g806) & (g827) & (!g858) & (!g1896) & (g2041)) + ((g806) & (g827) & (!g858) & (g1896) & (!g2041)) + ((g806) & (g827) & (g858) & (!g1896) & (!g2041)) + ((g806) & (g827) & (g858) & (g1896) & (g2041)));
	assign g7876 = (((!g3429) & (g4164) & (!g2043)) + ((!g3429) & (g4164) & (g2043)) + ((g3429) & (!g4164) & (g2043)) + ((g3429) & (g4164) & (g2043)));
	assign g2044 = (((!g814) & (!g827) & (!g860) & (!g1904) & (g2043)) + ((!g814) & (!g827) & (!g860) & (g1904) & (g2043)) + ((!g814) & (!g827) & (g860) & (!g1904) & (g2043)) + ((!g814) & (!g827) & (g860) & (g1904) & (g2043)) + ((!g814) & (g827) & (!g860) & (!g1904) & (g2043)) + ((!g814) & (g827) & (!g860) & (g1904) & (g2043)) + ((!g814) & (g827) & (g860) & (!g1904) & (!g2043)) + ((!g814) & (g827) & (g860) & (g1904) & (!g2043)) + ((g814) & (!g827) & (!g860) & (!g1904) & (g2043)) + ((g814) & (!g827) & (!g860) & (g1904) & (g2043)) + ((g814) & (!g827) & (g860) & (!g1904) & (g2043)) + ((g814) & (!g827) & (g860) & (g1904) & (g2043)) + ((g814) & (g827) & (!g860) & (!g1904) & (g2043)) + ((g814) & (g827) & (!g860) & (g1904) & (!g2043)) + ((g814) & (g827) & (g860) & (!g1904) & (!g2043)) + ((g814) & (g827) & (g860) & (g1904) & (g2043)));
	assign g7877 = (((!g2017) & (g6874) & (!g2045)) + ((!g2017) & (g6874) & (g2045)) + ((g2017) & (!g6874) & (g2045)) + ((g2017) & (g6874) & (g2045)));
	assign g2046 = (((!g822) & (!g827) & (!g862) & (!g1912) & (g2045)) + ((!g822) & (!g827) & (!g862) & (g1912) & (g2045)) + ((!g822) & (!g827) & (g862) & (!g1912) & (g2045)) + ((!g822) & (!g827) & (g862) & (g1912) & (g2045)) + ((!g822) & (g827) & (!g862) & (!g1912) & (g2045)) + ((!g822) & (g827) & (!g862) & (g1912) & (g2045)) + ((!g822) & (g827) & (g862) & (!g1912) & (!g2045)) + ((!g822) & (g827) & (g862) & (g1912) & (!g2045)) + ((g822) & (!g827) & (!g862) & (!g1912) & (g2045)) + ((g822) & (!g827) & (!g862) & (g1912) & (g2045)) + ((g822) & (!g827) & (g862) & (!g1912) & (g2045)) + ((g822) & (!g827) & (g862) & (g1912) & (g2045)) + ((g822) & (g827) & (!g862) & (!g1912) & (g2045)) + ((g822) & (g827) & (!g862) & (g1912) & (!g2045)) + ((g822) & (g827) & (g862) & (!g1912) & (!g2045)) + ((g822) & (g827) & (g862) & (g1912) & (g2045)));
	assign g7878 = (((!g3429) & (g4171) & (!g2047)) + ((!g3429) & (g4171) & (g2047)) + ((g3429) & (!g4171) & (g2047)) + ((g3429) & (g4171) & (g2047)));
	assign g7879 = (((!g3464) & (g4174) & (!g2048)) + ((!g3464) & (g4174) & (g2048)) + ((g3464) & (!g4174) & (g2048)) + ((g3464) & (g4174) & (g2048)));
	assign g2049 = (((!g1974) & (!g1975) & (!g1976) & (!g2047) & (g2048)) + ((!g1974) & (!g1975) & (!g1976) & (g2047) & (!g2048)) + ((!g1974) & (!g1975) & (g1976) & (!g2047) & (g2048)) + ((!g1974) & (!g1975) & (g1976) & (g2047) & (!g2048)) + ((!g1974) & (g1975) & (!g1976) & (!g2047) & (g2048)) + ((!g1974) & (g1975) & (!g1976) & (g2047) & (!g2048)) + ((!g1974) & (g1975) & (g1976) & (!g2047) & (!g2048)) + ((!g1974) & (g1975) & (g1976) & (g2047) & (g2048)) + ((g1974) & (!g1975) & (!g1976) & (!g2047) & (g2048)) + ((g1974) & (!g1975) & (!g1976) & (g2047) & (!g2048)) + ((g1974) & (!g1975) & (g1976) & (!g2047) & (!g2048)) + ((g1974) & (!g1975) & (g1976) & (g2047) & (g2048)) + ((g1974) & (g1975) & (!g1976) & (!g2047) & (!g2048)) + ((g1974) & (g1975) & (!g1976) & (g2047) & (g2048)) + ((g1974) & (g1975) & (g1976) & (!g2047) & (!g2048)) + ((g1974) & (g1975) & (g1976) & (g2047) & (g2048)));
	assign g2050 = (((!g2008) & (!g2009) & (!g2011) & (!g2012) & (g2013) & (g2014)) + ((!g2008) & (!g2009) & (!g2011) & (g2012) & (g2013) & (g2014)) + ((!g2008) & (!g2009) & (g2011) & (!g2012) & (g2013) & (g2014)) + ((!g2008) & (!g2009) & (g2011) & (g2012) & (!g2013) & (g2014)) + ((!g2008) & (!g2009) & (g2011) & (g2012) & (g2013) & (!g2014)) + ((!g2008) & (!g2009) & (g2011) & (g2012) & (g2013) & (g2014)) + ((!g2008) & (g2009) & (!g2011) & (!g2012) & (g2013) & (g2014)) + ((!g2008) & (g2009) & (!g2011) & (g2012) & (!g2013) & (g2014)) + ((!g2008) & (g2009) & (!g2011) & (g2012) & (g2013) & (!g2014)) + ((!g2008) & (g2009) & (!g2011) & (g2012) & (g2013) & (g2014)) + ((!g2008) & (g2009) & (g2011) & (!g2012) & (!g2013) & (g2014)) + ((!g2008) & (g2009) & (g2011) & (!g2012) & (g2013) & (!g2014)) + ((!g2008) & (g2009) & (g2011) & (!g2012) & (g2013) & (g2014)) + ((!g2008) & (g2009) & (g2011) & (g2012) & (!g2013) & (g2014)) + ((!g2008) & (g2009) & (g2011) & (g2012) & (g2013) & (!g2014)) + ((!g2008) & (g2009) & (g2011) & (g2012) & (g2013) & (g2014)) + ((g2008) & (!g2009) & (!g2011) & (!g2012) & (g2013) & (g2014)) + ((g2008) & (!g2009) & (!g2011) & (g2012) & (!g2013) & (g2014)) + ((g2008) & (!g2009) & (!g2011) & (g2012) & (g2013) & (!g2014)) + ((g2008) & (!g2009) & (!g2011) & (g2012) & (g2013) & (g2014)) + ((g2008) & (!g2009) & (g2011) & (!g2012) & (!g2013) & (g2014)) + ((g2008) & (!g2009) & (g2011) & (!g2012) & (g2013) & (!g2014)) + ((g2008) & (!g2009) & (g2011) & (!g2012) & (g2013) & (g2014)) + ((g2008) & (!g2009) & (g2011) & (g2012) & (!g2013) & (g2014)) + ((g2008) & (!g2009) & (g2011) & (g2012) & (g2013) & (!g2014)) + ((g2008) & (!g2009) & (g2011) & (g2012) & (g2013) & (g2014)) + ((g2008) & (g2009) & (!g2011) & (!g2012) & (g2013) & (g2014)) + ((g2008) & (g2009) & (!g2011) & (g2012) & (!g2013) & (g2014)) + ((g2008) & (g2009) & (!g2011) & (g2012) & (g2013) & (!g2014)) + ((g2008) & (g2009) & (!g2011) & (g2012) & (g2013) & (g2014)) + ((g2008) & (g2009) & (g2011) & (!g2012) & (!g2013) & (g2014)) + ((g2008) & (g2009) & (g2011) & (!g2012) & (g2013) & (!g2014)) + ((g2008) & (g2009) & (g2011) & (!g2012) & (g2013) & (g2014)) + ((g2008) & (g2009) & (g2011) & (g2012) & (!g2013) & (g2014)) + ((g2008) & (g2009) & (g2011) & (g2012) & (g2013) & (!g2014)) + ((g2008) & (g2009) & (g2011) & (g2012) & (g2013) & (g2014)));
	assign g7880 = (((!g3429) & (g4178) & (!g2051)) + ((!g3429) & (g4178) & (g2051)) + ((g3429) & (!g4178) & (g2051)) + ((g3429) & (g4178) & (g2051)));
	assign g7881 = (((!g3499) & (g4181) & (!g2052)) + ((!g3499) & (g4181) & (g2052)) + ((g3499) & (!g4181) & (g2052)) + ((g3499) & (g4181) & (g2052)));
	assign g2053 = (((!g790) & (g840) & (!g1884) & (g1977)) + ((!g790) & (g840) & (g1884) & (g1977)) + ((g790) & (!g840) & (g1884) & (g1977)) + ((g790) & (g840) & (!g1884) & (g1977)) + ((g790) & (g840) & (g1884) & (!g1977)) + ((g790) & (g840) & (g1884) & (g1977)));
	assign g2054 = (((!g827) & (!g867) & (g1979) & (!g2053)) + ((!g827) & (!g867) & (g1979) & (g2053)) + ((!g827) & (g867) & (g1979) & (!g2053)) + ((!g827) & (g867) & (g1979) & (g2053)) + ((g827) & (!g867) & (!g1979) & (g2053)) + ((g827) & (!g867) & (g1979) & (!g2053)) + ((g827) & (g867) & (!g1979) & (!g2053)) + ((g827) & (g867) & (g1979) & (g2053)));
	assign g7882 = (((!g3464) & (g4188) & (!g2055)) + ((!g3464) & (g4188) & (g2055)) + ((g3464) & (!g4188) & (g2055)) + ((g3464) & (g4188) & (g2055)));
	assign g2056 = (((!g792) & (g848) & (!g1886) & (g2032)) + ((!g792) & (g848) & (g1886) & (g2032)) + ((g792) & (!g848) & (g1886) & (g2032)) + ((g792) & (g848) & (!g1886) & (g2032)) + ((g792) & (g848) & (g1886) & (!g2032)) + ((g792) & (g848) & (g1886) & (g2032)));
	assign g2057 = (((!g827) & (!g869) & (g2055) & (!g2056)) + ((!g827) & (!g869) & (g2055) & (g2056)) + ((!g827) & (g869) & (g2055) & (!g2056)) + ((!g827) & (g869) & (g2055) & (g2056)) + ((g827) & (!g869) & (!g2055) & (g2056)) + ((g827) & (!g869) & (g2055) & (!g2056)) + ((g827) & (g869) & (!g2055) & (!g2056)) + ((g827) & (g869) & (g2055) & (g2056)));
	assign g2058 = (((!g794) & (g856) & (!g1888) & (g1978)) + ((!g794) & (g856) & (g1888) & (g1978)) + ((g794) & (!g856) & (g1888) & (g1978)) + ((g794) & (g856) & (!g1888) & (g1978)) + ((g794) & (g856) & (g1888) & (!g1978)) + ((g794) & (g856) & (g1888) & (g1978)));
	assign g2059 = (((!g827) & (!g871) & (g1980) & (!g2058)) + ((!g827) & (!g871) & (g1980) & (g2058)) + ((!g827) & (g871) & (g1980) & (!g2058)) + ((!g827) & (g871) & (g1980) & (g2058)) + ((g827) & (!g871) & (!g1980) & (g2058)) + ((g827) & (!g871) & (g1980) & (!g2058)) + ((g827) & (g871) & (!g1980) & (!g2058)) + ((g827) & (g871) & (g1980) & (g2058)));
	assign g2060 = (((!g800) & (g834) & (!g1890) & (g1939)) + ((!g800) & (g834) & (g1890) & (g1939)) + ((g800) & (!g834) & (g1890) & (g1939)) + ((g800) & (g834) & (!g1890) & (g1939)) + ((g800) & (g834) & (g1890) & (!g1939)) + ((g800) & (g834) & (g1890) & (g1939)));
	assign g2061 = (((!g827) & (!g873) & (g1941) & (!g2060)) + ((!g827) & (!g873) & (g1941) & (g2060)) + ((!g827) & (g873) & (g1941) & (!g2060)) + ((!g827) & (g873) & (g1941) & (g2060)) + ((g827) & (!g873) & (!g1941) & (g2060)) + ((g827) & (!g873) & (g1941) & (!g2060)) + ((g827) & (g873) & (!g1941) & (!g2060)) + ((g827) & (g873) & (g1941) & (g2060)));
	assign g7883 = (((!g2017) & (g6855) & (!g2062)) + ((!g2017) & (g6855) & (g2062)) + ((g2017) & (!g6855) & (g2062)) + ((g2017) & (g6855) & (g2062)));
	assign g2063 = (((!g802) & (g842) & (!g1892) & (g2026)) + ((!g802) & (g842) & (g1892) & (g2026)) + ((g802) & (!g842) & (g1892) & (g2026)) + ((g802) & (g842) & (!g1892) & (g2026)) + ((g802) & (g842) & (g1892) & (!g2026)) + ((g802) & (g842) & (g1892) & (g2026)));
	assign g2064 = (((!g827) & (!g875) & (g2062) & (!g2063)) + ((!g827) & (!g875) & (g2062) & (g2063)) + ((!g827) & (g875) & (g2062) & (!g2063)) + ((!g827) & (g875) & (g2062) & (g2063)) + ((g827) & (!g875) & (!g2062) & (g2063)) + ((g827) & (!g875) & (g2062) & (!g2063)) + ((g827) & (g875) & (!g2062) & (!g2063)) + ((g827) & (g875) & (g2062) & (g2063)));
	assign g7884 = (((!g3499) & (g4200) & (!g2065)) + ((!g3499) & (g4200) & (g2065)) + ((g3499) & (!g4200) & (g2065)) + ((g3499) & (g4200) & (g2065)));
	assign g2066 = (((!g804) & (g850) & (!g1894) & (g2034)) + ((!g804) & (g850) & (g1894) & (g2034)) + ((g804) & (!g850) & (g1894) & (g2034)) + ((g804) & (g850) & (!g1894) & (g2034)) + ((g804) & (g850) & (g1894) & (!g2034)) + ((g804) & (g850) & (g1894) & (g2034)));
	assign g2067 = (((!g827) & (!g877) & (g2065) & (!g2066)) + ((!g827) & (!g877) & (g2065) & (g2066)) + ((!g827) & (g877) & (g2065) & (!g2066)) + ((!g827) & (g877) & (g2065) & (g2066)) + ((g827) & (!g877) & (!g2065) & (g2066)) + ((g827) & (!g877) & (g2065) & (!g2066)) + ((g827) & (g877) & (!g2065) & (!g2066)) + ((g827) & (g877) & (g2065) & (g2066)));
	assign g7885 = (((!g3464) & (g4207) & (!g2068)) + ((!g3464) & (g4207) & (g2068)) + ((g3464) & (!g4207) & (g2068)) + ((g3464) & (g4207) & (g2068)));
	assign g2069 = (((!g806) & (g858) & (!g1896) & (g2041)) + ((!g806) & (g858) & (g1896) & (g2041)) + ((g806) & (!g858) & (g1896) & (g2041)) + ((g806) & (g858) & (!g1896) & (g2041)) + ((g806) & (g858) & (g1896) & (!g2041)) + ((g806) & (g858) & (g1896) & (g2041)));
	assign g2070 = (((!g827) & (!g879) & (g2068) & (!g2069)) + ((!g827) & (!g879) & (g2068) & (g2069)) + ((!g827) & (g879) & (g2068) & (!g2069)) + ((!g827) & (g879) & (g2068) & (g2069)) + ((g827) & (!g879) & (!g2068) & (g2069)) + ((g827) & (!g879) & (g2068) & (!g2069)) + ((g827) & (g879) & (!g2068) & (!g2069)) + ((g827) & (g879) & (g2068) & (g2069)));
	assign g7886 = (((!g3499) & (g4214) & (!g2071)) + ((!g3499) & (g4214) & (g2071)) + ((g3499) & (!g4214) & (g2071)) + ((g3499) & (g4214) & (g2071)));
	assign g2072 = (((!g808) & (g836) & (!g1898) & (g2022)) + ((!g808) & (g836) & (g1898) & (g2022)) + ((g808) & (!g836) & (g1898) & (g2022)) + ((g808) & (g836) & (!g1898) & (g2022)) + ((g808) & (g836) & (g1898) & (!g2022)) + ((g808) & (g836) & (g1898) & (g2022)));
	assign g2073 = (((!g827) & (!g881) & (g2071) & (!g2072)) + ((!g827) & (!g881) & (g2071) & (g2072)) + ((!g827) & (g881) & (g2071) & (!g2072)) + ((!g827) & (g881) & (g2071) & (g2072)) + ((g827) & (!g881) & (!g2071) & (g2072)) + ((g827) & (!g881) & (g2071) & (!g2072)) + ((g827) & (g881) & (!g2071) & (!g2072)) + ((g827) & (g881) & (g2071) & (g2072)));
	assign g7887 = (((!g3464) & (g4222) & (!g2074)) + ((!g3464) & (g4222) & (g2074)) + ((g3464) & (!g4222) & (g2074)) + ((g3464) & (g4222) & (g2074)));
	assign g2075 = (((!g810) & (g844) & (!g1900) & (g2028)) + ((!g810) & (g844) & (g1900) & (g2028)) + ((g810) & (!g844) & (g1900) & (g2028)) + ((g810) & (g844) & (!g1900) & (g2028)) + ((g810) & (g844) & (g1900) & (!g2028)) + ((g810) & (g844) & (g1900) & (g2028)));
	assign g2076 = (((!g827) & (!g883) & (g2074) & (!g2075)) + ((!g827) & (!g883) & (g2074) & (g2075)) + ((!g827) & (g883) & (g2074) & (!g2075)) + ((!g827) & (g883) & (g2074) & (g2075)) + ((g827) & (!g883) & (!g2074) & (g2075)) + ((g827) & (!g883) & (g2074) & (!g2075)) + ((g827) & (g883) & (!g2074) & (!g2075)) + ((g827) & (g883) & (g2074) & (g2075)));
	assign g7888 = (((!g2017) & (g6848) & (!g2077)) + ((!g2017) & (g6848) & (g2077)) + ((g2017) & (!g6848) & (g2077)) + ((g2017) & (g6848) & (g2077)));
	assign g2078 = (((!g812) & (g852) & (!g1902) & (g2036)) + ((!g812) & (g852) & (g1902) & (g2036)) + ((g812) & (!g852) & (g1902) & (g2036)) + ((g812) & (g852) & (!g1902) & (g2036)) + ((g812) & (g852) & (g1902) & (!g2036)) + ((g812) & (g852) & (g1902) & (g2036)));
	assign g2079 = (((!g827) & (!g885) & (g2077) & (!g2078)) + ((!g827) & (!g885) & (g2077) & (g2078)) + ((!g827) & (g885) & (g2077) & (!g2078)) + ((!g827) & (g885) & (g2077) & (g2078)) + ((g827) & (!g885) & (!g2077) & (g2078)) + ((g827) & (!g885) & (g2077) & (!g2078)) + ((g827) & (g885) & (!g2077) & (!g2078)) + ((g827) & (g885) & (g2077) & (g2078)));
	assign g7889 = (((!g3429) & (g4229) & (!g2080)) + ((!g3429) & (g4229) & (g2080)) + ((g3429) & (!g4229) & (g2080)) + ((g3429) & (g4229) & (g2080)));
	assign g2081 = (((!g814) & (g860) & (!g1904) & (g2043)) + ((!g814) & (g860) & (g1904) & (g2043)) + ((g814) & (!g860) & (g1904) & (g2043)) + ((g814) & (g860) & (!g1904) & (g2043)) + ((g814) & (g860) & (g1904) & (!g2043)) + ((g814) & (g860) & (g1904) & (g2043)));
	assign g2082 = (((!g827) & (!g887) & (g2080) & (!g2081)) + ((!g827) & (!g887) & (g2080) & (g2081)) + ((!g827) & (g887) & (g2080) & (!g2081)) + ((!g827) & (g887) & (g2080) & (g2081)) + ((g827) & (!g887) & (!g2080) & (g2081)) + ((g827) & (!g887) & (g2080) & (!g2081)) + ((g827) & (g887) & (!g2080) & (!g2081)) + ((g827) & (g887) & (g2080) & (g2081)));
	assign g2083 = (((!g816) & (g838) & (!g1906) & (g1940)) + ((!g816) & (g838) & (g1906) & (g1940)) + ((g816) & (!g838) & (g1906) & (g1940)) + ((g816) & (g838) & (!g1906) & (g1940)) + ((g816) & (g838) & (g1906) & (!g1940)) + ((g816) & (g838) & (g1906) & (g1940)));
	assign g2084 = (((!g827) & (!g889) & (g1942) & (!g2083)) + ((!g827) & (!g889) & (g1942) & (g2083)) + ((!g827) & (g889) & (g1942) & (!g2083)) + ((!g827) & (g889) & (g1942) & (g2083)) + ((g827) & (!g889) & (!g1942) & (g2083)) + ((g827) & (!g889) & (g1942) & (!g2083)) + ((g827) & (g889) & (!g1942) & (!g2083)) + ((g827) & (g889) & (g1942) & (g2083)));
	assign g7890 = (((!g3499) & (g4236) & (!g2085)) + ((!g3499) & (g4236) & (g2085)) + ((g3499) & (!g4236) & (g2085)) + ((g3499) & (g4236) & (g2085)));
	assign g2086 = (((!g818) & (g846) & (!g1908) & (g2030)) + ((!g818) & (g846) & (g1908) & (g2030)) + ((g818) & (!g846) & (g1908) & (g2030)) + ((g818) & (g846) & (!g1908) & (g2030)) + ((g818) & (g846) & (g1908) & (!g2030)) + ((g818) & (g846) & (g1908) & (g2030)));
	assign g2087 = (((!g827) & (!g891) & (g2085) & (!g2086)) + ((!g827) & (!g891) & (g2085) & (g2086)) + ((!g827) & (g891) & (g2085) & (!g2086)) + ((!g827) & (g891) & (g2085) & (g2086)) + ((g827) & (!g891) & (!g2085) & (g2086)) + ((g827) & (!g891) & (g2085) & (!g2086)) + ((g827) & (g891) & (!g2085) & (!g2086)) + ((g827) & (g891) & (g2085) & (g2086)));
	assign g7891 = (((!g3429) & (g4239) & (!g2088)) + ((!g3429) & (g4239) & (g2088)) + ((g3429) & (!g4239) & (g2088)) + ((g3429) & (g4239) & (g2088)));
	assign g2089 = (((!g820) & (g854) & (!g1910) & (g2038)) + ((!g820) & (g854) & (g1910) & (g2038)) + ((g820) & (!g854) & (g1910) & (g2038)) + ((g820) & (g854) & (!g1910) & (g2038)) + ((g820) & (g854) & (g1910) & (!g2038)) + ((g820) & (g854) & (g1910) & (g2038)));
	assign g2090 = (((!g827) & (!g893) & (g2088) & (!g2089)) + ((!g827) & (!g893) & (g2088) & (g2089)) + ((!g827) & (g893) & (g2088) & (!g2089)) + ((!g827) & (g893) & (g2088) & (g2089)) + ((g827) & (!g893) & (!g2088) & (g2089)) + ((g827) & (!g893) & (g2088) & (!g2089)) + ((g827) & (g893) & (!g2088) & (!g2089)) + ((g827) & (g893) & (g2088) & (g2089)));
	assign g7892 = (((!g2017) & (g6841) & (!g2091)) + ((!g2017) & (g6841) & (g2091)) + ((g2017) & (!g6841) & (g2091)) + ((g2017) & (g6841) & (g2091)));
	assign g2092 = (((!g822) & (g862) & (!g1912) & (g2045)) + ((!g822) & (g862) & (g1912) & (g2045)) + ((g822) & (!g862) & (g1912) & (g2045)) + ((g822) & (g862) & (!g1912) & (g2045)) + ((g822) & (g862) & (g1912) & (!g2045)) + ((g822) & (g862) & (g1912) & (g2045)));
	assign g2093 = (((!g827) & (!g895) & (g2091) & (!g2092)) + ((!g827) & (!g895) & (g2091) & (g2092)) + ((!g827) & (g895) & (g2091) & (!g2092)) + ((!g827) & (g895) & (g2091) & (g2092)) + ((g827) & (!g895) & (!g2091) & (g2092)) + ((g827) & (!g895) & (g2091) & (!g2092)) + ((g827) & (g895) & (!g2091) & (!g2092)) + ((g827) & (g895) & (g2091) & (g2092)));
	assign g2094 = (((!g2047) & (g2048)) + ((g2047) & (!g2048)));
	assign g2095 = (((!g1971) & (!g1972) & (!g1973) & (g1975) & (g1976) & (g2094)) + ((!g1971) & (!g1972) & (g1973) & (g1975) & (g1976) & (g2094)) + ((!g1971) & (g1972) & (!g1973) & (g1975) & (g1976) & (g2094)) + ((!g1971) & (g1972) & (g1973) & (!g1975) & (g1976) & (g2094)) + ((!g1971) & (g1972) & (g1973) & (g1975) & (!g1976) & (g2094)) + ((!g1971) & (g1972) & (g1973) & (g1975) & (g1976) & (g2094)) + ((g1971) & (!g1972) & (!g1973) & (g1975) & (g1976) & (g2094)) + ((g1971) & (!g1972) & (g1973) & (!g1975) & (g1976) & (g2094)) + ((g1971) & (!g1972) & (g1973) & (g1975) & (!g1976) & (g2094)) + ((g1971) & (!g1972) & (g1973) & (g1975) & (g1976) & (g2094)) + ((g1971) & (g1972) & (!g1973) & (!g1975) & (g1976) & (g2094)) + ((g1971) & (g1972) & (!g1973) & (g1975) & (!g1976) & (g2094)) + ((g1971) & (g1972) & (!g1973) & (g1975) & (g1976) & (g2094)) + ((g1971) & (g1972) & (g1973) & (!g1975) & (g1976) & (g2094)) + ((g1971) & (g1972) & (g1973) & (g1975) & (!g1976) & (g2094)) + ((g1971) & (g1972) & (g1973) & (g1975) & (g1976) & (g2094)));
	assign g2096 = (((g2047) & (g2048)));
	assign g2097 = (((!g2095) & (g2096)) + ((g2095) & (!g2096)) + ((g2095) & (g2096)));
	assign g7893 = (((!g3429) & (g4246) & (!g2098)) + ((!g3429) & (g4246) & (g2098)) + ((g3429) & (!g4246) & (g2098)) + ((g3429) & (g4246) & (g2098)));
	assign g7894 = (((!g3464) & (g4250) & (!g2099)) + ((!g3464) & (g4250) & (g2099)) + ((g3464) & (!g4250) & (g2099)) + ((g3464) & (g4250) & (g2099)));
	assign g7895 = (((!g3429) & (g4253) & (!g2100)) + ((!g3429) & (g4253) & (g2100)) + ((g3429) & (!g4253) & (g2100)) + ((g3429) & (g4253) & (g2100)));
	assign g7896 = (((!g3499) & (g4257) & (!g2101)) + ((!g3499) & (g4257) & (g2101)) + ((g3499) & (!g4257) & (g2101)) + ((g3499) & (g4257) & (g2101)));
	assign g2102 = (((!g2050) & (!g2051) & (!g2052) & (!g2100) & (g2101)) + ((!g2050) & (!g2051) & (!g2052) & (g2100) & (!g2101)) + ((!g2050) & (!g2051) & (g2052) & (!g2100) & (g2101)) + ((!g2050) & (!g2051) & (g2052) & (g2100) & (!g2101)) + ((!g2050) & (g2051) & (!g2052) & (!g2100) & (g2101)) + ((!g2050) & (g2051) & (!g2052) & (g2100) & (!g2101)) + ((!g2050) & (g2051) & (g2052) & (!g2100) & (!g2101)) + ((!g2050) & (g2051) & (g2052) & (g2100) & (g2101)) + ((g2050) & (!g2051) & (!g2052) & (!g2100) & (g2101)) + ((g2050) & (!g2051) & (!g2052) & (g2100) & (!g2101)) + ((g2050) & (!g2051) & (g2052) & (!g2100) & (!g2101)) + ((g2050) & (!g2051) & (g2052) & (g2100) & (g2101)) + ((g2050) & (g2051) & (!g2052) & (!g2100) & (!g2101)) + ((g2050) & (g2051) & (!g2052) & (g2100) & (g2101)) + ((g2050) & (g2051) & (g2052) & (!g2100) & (!g2101)) + ((g2050) & (g2051) & (g2052) & (g2100) & (g2101)));
	assign g2103 = (((!g827) & (!g873) & (!g901) & (!g1941) & (g1944) & (!g2060)) + ((!g827) & (!g873) & (!g901) & (!g1941) & (g1944) & (g2060)) + ((!g827) & (!g873) & (!g901) & (g1941) & (g1944) & (!g2060)) + ((!g827) & (!g873) & (!g901) & (g1941) & (g1944) & (g2060)) + ((!g827) & (!g873) & (g901) & (!g1941) & (g1944) & (!g2060)) + ((!g827) & (!g873) & (g901) & (!g1941) & (g1944) & (g2060)) + ((!g827) & (!g873) & (g901) & (g1941) & (g1944) & (!g2060)) + ((!g827) & (!g873) & (g901) & (g1941) & (g1944) & (g2060)) + ((!g827) & (g873) & (!g901) & (!g1941) & (g1944) & (!g2060)) + ((!g827) & (g873) & (!g901) & (!g1941) & (g1944) & (g2060)) + ((!g827) & (g873) & (!g901) & (g1941) & (g1944) & (!g2060)) + ((!g827) & (g873) & (!g901) & (g1941) & (g1944) & (g2060)) + ((!g827) & (g873) & (g901) & (!g1941) & (g1944) & (!g2060)) + ((!g827) & (g873) & (g901) & (!g1941) & (g1944) & (g2060)) + ((!g827) & (g873) & (g901) & (g1941) & (g1944) & (!g2060)) + ((!g827) & (g873) & (g901) & (g1941) & (g1944) & (g2060)) + ((g827) & (!g873) & (!g901) & (!g1941) & (g1944) & (!g2060)) + ((g827) & (!g873) & (!g901) & (!g1941) & (g1944) & (g2060)) + ((g827) & (!g873) & (!g901) & (g1941) & (!g1944) & (g2060)) + ((g827) & (!g873) & (!g901) & (g1941) & (g1944) & (!g2060)) + ((g827) & (!g873) & (g901) & (!g1941) & (!g1944) & (!g2060)) + ((g827) & (!g873) & (g901) & (!g1941) & (!g1944) & (g2060)) + ((g827) & (!g873) & (g901) & (g1941) & (!g1944) & (!g2060)) + ((g827) & (!g873) & (g901) & (g1941) & (g1944) & (g2060)) + ((g827) & (g873) & (!g901) & (!g1941) & (!g1944) & (g2060)) + ((g827) & (g873) & (!g901) & (!g1941) & (g1944) & (!g2060)) + ((g827) & (g873) & (!g901) & (g1941) & (!g1944) & (!g2060)) + ((g827) & (g873) & (!g901) & (g1941) & (!g1944) & (g2060)) + ((g827) & (g873) & (g901) & (!g1941) & (!g1944) & (!g2060)) + ((g827) & (g873) & (g901) & (!g1941) & (g1944) & (g2060)) + ((g827) & (g873) & (g901) & (g1941) & (g1944) & (!g2060)) + ((g827) & (g873) & (g901) & (g1941) & (g1944) & (g2060)));
	assign g7897 = (((!g3499) & (g4261) & (!g2104)) + ((!g3499) & (g4261) & (g2104)) + ((g3499) & (!g4261) & (g2104)) + ((g3499) & (g4261) & (g2104)));
	assign g2105 = (((!g827) & (!g881) & (!g903) & (!g2071) & (g2104) & (!g2072)) + ((!g827) & (!g881) & (!g903) & (!g2071) & (g2104) & (g2072)) + ((!g827) & (!g881) & (!g903) & (g2071) & (g2104) & (!g2072)) + ((!g827) & (!g881) & (!g903) & (g2071) & (g2104) & (g2072)) + ((!g827) & (!g881) & (g903) & (!g2071) & (g2104) & (!g2072)) + ((!g827) & (!g881) & (g903) & (!g2071) & (g2104) & (g2072)) + ((!g827) & (!g881) & (g903) & (g2071) & (g2104) & (!g2072)) + ((!g827) & (!g881) & (g903) & (g2071) & (g2104) & (g2072)) + ((!g827) & (g881) & (!g903) & (!g2071) & (g2104) & (!g2072)) + ((!g827) & (g881) & (!g903) & (!g2071) & (g2104) & (g2072)) + ((!g827) & (g881) & (!g903) & (g2071) & (g2104) & (!g2072)) + ((!g827) & (g881) & (!g903) & (g2071) & (g2104) & (g2072)) + ((!g827) & (g881) & (g903) & (!g2071) & (g2104) & (!g2072)) + ((!g827) & (g881) & (g903) & (!g2071) & (g2104) & (g2072)) + ((!g827) & (g881) & (g903) & (g2071) & (g2104) & (!g2072)) + ((!g827) & (g881) & (g903) & (g2071) & (g2104) & (g2072)) + ((g827) & (!g881) & (!g903) & (!g2071) & (g2104) & (!g2072)) + ((g827) & (!g881) & (!g903) & (!g2071) & (g2104) & (g2072)) + ((g827) & (!g881) & (!g903) & (g2071) & (!g2104) & (g2072)) + ((g827) & (!g881) & (!g903) & (g2071) & (g2104) & (!g2072)) + ((g827) & (!g881) & (g903) & (!g2071) & (!g2104) & (!g2072)) + ((g827) & (!g881) & (g903) & (!g2071) & (!g2104) & (g2072)) + ((g827) & (!g881) & (g903) & (g2071) & (!g2104) & (!g2072)) + ((g827) & (!g881) & (g903) & (g2071) & (g2104) & (g2072)) + ((g827) & (g881) & (!g903) & (!g2071) & (!g2104) & (g2072)) + ((g827) & (g881) & (!g903) & (!g2071) & (g2104) & (!g2072)) + ((g827) & (g881) & (!g903) & (g2071) & (!g2104) & (!g2072)) + ((g827) & (g881) & (!g903) & (g2071) & (!g2104) & (g2072)) + ((g827) & (g881) & (g903) & (!g2071) & (!g2104) & (!g2072)) + ((g827) & (g881) & (g903) & (!g2071) & (g2104) & (g2072)) + ((g827) & (g881) & (g903) & (g2071) & (g2104) & (!g2072)) + ((g827) & (g881) & (g903) & (g2071) & (g2104) & (g2072)));
	assign g2106 = (((!g827) & (!g889) & (!g905) & (!g1942) & (g1945) & (!g2083)) + ((!g827) & (!g889) & (!g905) & (!g1942) & (g1945) & (g2083)) + ((!g827) & (!g889) & (!g905) & (g1942) & (g1945) & (!g2083)) + ((!g827) & (!g889) & (!g905) & (g1942) & (g1945) & (g2083)) + ((!g827) & (!g889) & (g905) & (!g1942) & (g1945) & (!g2083)) + ((!g827) & (!g889) & (g905) & (!g1942) & (g1945) & (g2083)) + ((!g827) & (!g889) & (g905) & (g1942) & (g1945) & (!g2083)) + ((!g827) & (!g889) & (g905) & (g1942) & (g1945) & (g2083)) + ((!g827) & (g889) & (!g905) & (!g1942) & (g1945) & (!g2083)) + ((!g827) & (g889) & (!g905) & (!g1942) & (g1945) & (g2083)) + ((!g827) & (g889) & (!g905) & (g1942) & (g1945) & (!g2083)) + ((!g827) & (g889) & (!g905) & (g1942) & (g1945) & (g2083)) + ((!g827) & (g889) & (g905) & (!g1942) & (g1945) & (!g2083)) + ((!g827) & (g889) & (g905) & (!g1942) & (g1945) & (g2083)) + ((!g827) & (g889) & (g905) & (g1942) & (g1945) & (!g2083)) + ((!g827) & (g889) & (g905) & (g1942) & (g1945) & (g2083)) + ((g827) & (!g889) & (!g905) & (!g1942) & (g1945) & (!g2083)) + ((g827) & (!g889) & (!g905) & (!g1942) & (g1945) & (g2083)) + ((g827) & (!g889) & (!g905) & (g1942) & (!g1945) & (g2083)) + ((g827) & (!g889) & (!g905) & (g1942) & (g1945) & (!g2083)) + ((g827) & (!g889) & (g905) & (!g1942) & (!g1945) & (!g2083)) + ((g827) & (!g889) & (g905) & (!g1942) & (!g1945) & (g2083)) + ((g827) & (!g889) & (g905) & (g1942) & (!g1945) & (!g2083)) + ((g827) & (!g889) & (g905) & (g1942) & (g1945) & (g2083)) + ((g827) & (g889) & (!g905) & (!g1942) & (!g1945) & (g2083)) + ((g827) & (g889) & (!g905) & (!g1942) & (g1945) & (!g2083)) + ((g827) & (g889) & (!g905) & (g1942) & (!g1945) & (!g2083)) + ((g827) & (g889) & (!g905) & (g1942) & (!g1945) & (g2083)) + ((g827) & (g889) & (g905) & (!g1942) & (!g1945) & (!g2083)) + ((g827) & (g889) & (g905) & (!g1942) & (g1945) & (g2083)) + ((g827) & (g889) & (g905) & (g1942) & (g1945) & (!g2083)) + ((g827) & (g889) & (g905) & (g1942) & (g1945) & (g2083)));
	assign g2107 = (((!g827) & (!g867) & (!g907) & (!g1979) & (g1982) & (!g2053)) + ((!g827) & (!g867) & (!g907) & (!g1979) & (g1982) & (g2053)) + ((!g827) & (!g867) & (!g907) & (g1979) & (g1982) & (!g2053)) + ((!g827) & (!g867) & (!g907) & (g1979) & (g1982) & (g2053)) + ((!g827) & (!g867) & (g907) & (!g1979) & (g1982) & (!g2053)) + ((!g827) & (!g867) & (g907) & (!g1979) & (g1982) & (g2053)) + ((!g827) & (!g867) & (g907) & (g1979) & (g1982) & (!g2053)) + ((!g827) & (!g867) & (g907) & (g1979) & (g1982) & (g2053)) + ((!g827) & (g867) & (!g907) & (!g1979) & (g1982) & (!g2053)) + ((!g827) & (g867) & (!g907) & (!g1979) & (g1982) & (g2053)) + ((!g827) & (g867) & (!g907) & (g1979) & (g1982) & (!g2053)) + ((!g827) & (g867) & (!g907) & (g1979) & (g1982) & (g2053)) + ((!g827) & (g867) & (g907) & (!g1979) & (g1982) & (!g2053)) + ((!g827) & (g867) & (g907) & (!g1979) & (g1982) & (g2053)) + ((!g827) & (g867) & (g907) & (g1979) & (g1982) & (!g2053)) + ((!g827) & (g867) & (g907) & (g1979) & (g1982) & (g2053)) + ((g827) & (!g867) & (!g907) & (!g1979) & (g1982) & (!g2053)) + ((g827) & (!g867) & (!g907) & (!g1979) & (g1982) & (g2053)) + ((g827) & (!g867) & (!g907) & (g1979) & (!g1982) & (g2053)) + ((g827) & (!g867) & (!g907) & (g1979) & (g1982) & (!g2053)) + ((g827) & (!g867) & (g907) & (!g1979) & (!g1982) & (!g2053)) + ((g827) & (!g867) & (g907) & (!g1979) & (!g1982) & (g2053)) + ((g827) & (!g867) & (g907) & (g1979) & (!g1982) & (!g2053)) + ((g827) & (!g867) & (g907) & (g1979) & (g1982) & (g2053)) + ((g827) & (g867) & (!g907) & (!g1979) & (!g1982) & (g2053)) + ((g827) & (g867) & (!g907) & (!g1979) & (g1982) & (!g2053)) + ((g827) & (g867) & (!g907) & (g1979) & (!g1982) & (!g2053)) + ((g827) & (g867) & (!g907) & (g1979) & (!g1982) & (g2053)) + ((g827) & (g867) & (g907) & (!g1979) & (!g1982) & (!g2053)) + ((g827) & (g867) & (g907) & (!g1979) & (g1982) & (g2053)) + ((g827) & (g867) & (g907) & (g1979) & (g1982) & (!g2053)) + ((g827) & (g867) & (g907) & (g1979) & (g1982) & (g2053)));
	assign g7898 = (((!g2017) & (g6824) & (!g2108)) + ((!g2017) & (g6824) & (g2108)) + ((g2017) & (!g6824) & (g2108)) + ((g2017) & (g6824) & (g2108)));
	assign g2109 = (((!g827) & (!g875) & (!g909) & (!g2062) & (g2108) & (!g2063)) + ((!g827) & (!g875) & (!g909) & (!g2062) & (g2108) & (g2063)) + ((!g827) & (!g875) & (!g909) & (g2062) & (g2108) & (!g2063)) + ((!g827) & (!g875) & (!g909) & (g2062) & (g2108) & (g2063)) + ((!g827) & (!g875) & (g909) & (!g2062) & (g2108) & (!g2063)) + ((!g827) & (!g875) & (g909) & (!g2062) & (g2108) & (g2063)) + ((!g827) & (!g875) & (g909) & (g2062) & (g2108) & (!g2063)) + ((!g827) & (!g875) & (g909) & (g2062) & (g2108) & (g2063)) + ((!g827) & (g875) & (!g909) & (!g2062) & (g2108) & (!g2063)) + ((!g827) & (g875) & (!g909) & (!g2062) & (g2108) & (g2063)) + ((!g827) & (g875) & (!g909) & (g2062) & (g2108) & (!g2063)) + ((!g827) & (g875) & (!g909) & (g2062) & (g2108) & (g2063)) + ((!g827) & (g875) & (g909) & (!g2062) & (g2108) & (!g2063)) + ((!g827) & (g875) & (g909) & (!g2062) & (g2108) & (g2063)) + ((!g827) & (g875) & (g909) & (g2062) & (g2108) & (!g2063)) + ((!g827) & (g875) & (g909) & (g2062) & (g2108) & (g2063)) + ((g827) & (!g875) & (!g909) & (!g2062) & (g2108) & (!g2063)) + ((g827) & (!g875) & (!g909) & (!g2062) & (g2108) & (g2063)) + ((g827) & (!g875) & (!g909) & (g2062) & (!g2108) & (g2063)) + ((g827) & (!g875) & (!g909) & (g2062) & (g2108) & (!g2063)) + ((g827) & (!g875) & (g909) & (!g2062) & (!g2108) & (!g2063)) + ((g827) & (!g875) & (g909) & (!g2062) & (!g2108) & (g2063)) + ((g827) & (!g875) & (g909) & (g2062) & (!g2108) & (!g2063)) + ((g827) & (!g875) & (g909) & (g2062) & (g2108) & (g2063)) + ((g827) & (g875) & (!g909) & (!g2062) & (!g2108) & (g2063)) + ((g827) & (g875) & (!g909) & (!g2062) & (g2108) & (!g2063)) + ((g827) & (g875) & (!g909) & (g2062) & (!g2108) & (!g2063)) + ((g827) & (g875) & (!g909) & (g2062) & (!g2108) & (g2063)) + ((g827) & (g875) & (g909) & (!g2062) & (!g2108) & (!g2063)) + ((g827) & (g875) & (g909) & (!g2062) & (g2108) & (g2063)) + ((g827) & (g875) & (g909) & (g2062) & (g2108) & (!g2063)) + ((g827) & (g875) & (g909) & (g2062) & (g2108) & (g2063)));
	assign g7899 = (((!g3464) & (g4268) & (!g2110)) + ((!g3464) & (g4268) & (g2110)) + ((g3464) & (!g4268) & (g2110)) + ((g3464) & (g4268) & (g2110)));
	assign g2111 = (((!g827) & (!g883) & (!g911) & (!g2074) & (g2110) & (!g2075)) + ((!g827) & (!g883) & (!g911) & (!g2074) & (g2110) & (g2075)) + ((!g827) & (!g883) & (!g911) & (g2074) & (g2110) & (!g2075)) + ((!g827) & (!g883) & (!g911) & (g2074) & (g2110) & (g2075)) + ((!g827) & (!g883) & (g911) & (!g2074) & (g2110) & (!g2075)) + ((!g827) & (!g883) & (g911) & (!g2074) & (g2110) & (g2075)) + ((!g827) & (!g883) & (g911) & (g2074) & (g2110) & (!g2075)) + ((!g827) & (!g883) & (g911) & (g2074) & (g2110) & (g2075)) + ((!g827) & (g883) & (!g911) & (!g2074) & (g2110) & (!g2075)) + ((!g827) & (g883) & (!g911) & (!g2074) & (g2110) & (g2075)) + ((!g827) & (g883) & (!g911) & (g2074) & (g2110) & (!g2075)) + ((!g827) & (g883) & (!g911) & (g2074) & (g2110) & (g2075)) + ((!g827) & (g883) & (g911) & (!g2074) & (g2110) & (!g2075)) + ((!g827) & (g883) & (g911) & (!g2074) & (g2110) & (g2075)) + ((!g827) & (g883) & (g911) & (g2074) & (g2110) & (!g2075)) + ((!g827) & (g883) & (g911) & (g2074) & (g2110) & (g2075)) + ((g827) & (!g883) & (!g911) & (!g2074) & (g2110) & (!g2075)) + ((g827) & (!g883) & (!g911) & (!g2074) & (g2110) & (g2075)) + ((g827) & (!g883) & (!g911) & (g2074) & (!g2110) & (g2075)) + ((g827) & (!g883) & (!g911) & (g2074) & (g2110) & (!g2075)) + ((g827) & (!g883) & (g911) & (!g2074) & (!g2110) & (!g2075)) + ((g827) & (!g883) & (g911) & (!g2074) & (!g2110) & (g2075)) + ((g827) & (!g883) & (g911) & (g2074) & (!g2110) & (!g2075)) + ((g827) & (!g883) & (g911) & (g2074) & (g2110) & (g2075)) + ((g827) & (g883) & (!g911) & (!g2074) & (!g2110) & (g2075)) + ((g827) & (g883) & (!g911) & (!g2074) & (g2110) & (!g2075)) + ((g827) & (g883) & (!g911) & (g2074) & (!g2110) & (!g2075)) + ((g827) & (g883) & (!g911) & (g2074) & (!g2110) & (g2075)) + ((g827) & (g883) & (g911) & (!g2074) & (!g2110) & (!g2075)) + ((g827) & (g883) & (g911) & (!g2074) & (g2110) & (g2075)) + ((g827) & (g883) & (g911) & (g2074) & (g2110) & (!g2075)) + ((g827) & (g883) & (g911) & (g2074) & (g2110) & (g2075)));
	assign g7900 = (((!g3499) & (g4272) & (!g2112)) + ((!g3499) & (g4272) & (g2112)) + ((g3499) & (!g4272) & (g2112)) + ((g3499) & (g4272) & (g2112)));
	assign g2113 = (((!g827) & (!g891) & (!g913) & (!g2085) & (g2112) & (!g2086)) + ((!g827) & (!g891) & (!g913) & (!g2085) & (g2112) & (g2086)) + ((!g827) & (!g891) & (!g913) & (g2085) & (g2112) & (!g2086)) + ((!g827) & (!g891) & (!g913) & (g2085) & (g2112) & (g2086)) + ((!g827) & (!g891) & (g913) & (!g2085) & (g2112) & (!g2086)) + ((!g827) & (!g891) & (g913) & (!g2085) & (g2112) & (g2086)) + ((!g827) & (!g891) & (g913) & (g2085) & (g2112) & (!g2086)) + ((!g827) & (!g891) & (g913) & (g2085) & (g2112) & (g2086)) + ((!g827) & (g891) & (!g913) & (!g2085) & (g2112) & (!g2086)) + ((!g827) & (g891) & (!g913) & (!g2085) & (g2112) & (g2086)) + ((!g827) & (g891) & (!g913) & (g2085) & (g2112) & (!g2086)) + ((!g827) & (g891) & (!g913) & (g2085) & (g2112) & (g2086)) + ((!g827) & (g891) & (g913) & (!g2085) & (g2112) & (!g2086)) + ((!g827) & (g891) & (g913) & (!g2085) & (g2112) & (g2086)) + ((!g827) & (g891) & (g913) & (g2085) & (g2112) & (!g2086)) + ((!g827) & (g891) & (g913) & (g2085) & (g2112) & (g2086)) + ((g827) & (!g891) & (!g913) & (!g2085) & (g2112) & (!g2086)) + ((g827) & (!g891) & (!g913) & (!g2085) & (g2112) & (g2086)) + ((g827) & (!g891) & (!g913) & (g2085) & (!g2112) & (g2086)) + ((g827) & (!g891) & (!g913) & (g2085) & (g2112) & (!g2086)) + ((g827) & (!g891) & (g913) & (!g2085) & (!g2112) & (!g2086)) + ((g827) & (!g891) & (g913) & (!g2085) & (!g2112) & (g2086)) + ((g827) & (!g891) & (g913) & (g2085) & (!g2112) & (!g2086)) + ((g827) & (!g891) & (g913) & (g2085) & (g2112) & (g2086)) + ((g827) & (g891) & (!g913) & (!g2085) & (!g2112) & (g2086)) + ((g827) & (g891) & (!g913) & (!g2085) & (g2112) & (!g2086)) + ((g827) & (g891) & (!g913) & (g2085) & (!g2112) & (!g2086)) + ((g827) & (g891) & (!g913) & (g2085) & (!g2112) & (g2086)) + ((g827) & (g891) & (g913) & (!g2085) & (!g2112) & (!g2086)) + ((g827) & (g891) & (g913) & (!g2085) & (g2112) & (g2086)) + ((g827) & (g891) & (g913) & (g2085) & (g2112) & (!g2086)) + ((g827) & (g891) & (g913) & (g2085) & (g2112) & (g2086)));
	assign g7901 = (((!g3464) & (g4276) & (!g2114)) + ((!g3464) & (g4276) & (g2114)) + ((g3464) & (!g4276) & (g2114)) + ((g3464) & (g4276) & (g2114)));
	assign g2115 = (((!g827) & (!g869) & (!g915) & (!g2055) & (g2114) & (!g2056)) + ((!g827) & (!g869) & (!g915) & (!g2055) & (g2114) & (g2056)) + ((!g827) & (!g869) & (!g915) & (g2055) & (g2114) & (!g2056)) + ((!g827) & (!g869) & (!g915) & (g2055) & (g2114) & (g2056)) + ((!g827) & (!g869) & (g915) & (!g2055) & (g2114) & (!g2056)) + ((!g827) & (!g869) & (g915) & (!g2055) & (g2114) & (g2056)) + ((!g827) & (!g869) & (g915) & (g2055) & (g2114) & (!g2056)) + ((!g827) & (!g869) & (g915) & (g2055) & (g2114) & (g2056)) + ((!g827) & (g869) & (!g915) & (!g2055) & (g2114) & (!g2056)) + ((!g827) & (g869) & (!g915) & (!g2055) & (g2114) & (g2056)) + ((!g827) & (g869) & (!g915) & (g2055) & (g2114) & (!g2056)) + ((!g827) & (g869) & (!g915) & (g2055) & (g2114) & (g2056)) + ((!g827) & (g869) & (g915) & (!g2055) & (g2114) & (!g2056)) + ((!g827) & (g869) & (g915) & (!g2055) & (g2114) & (g2056)) + ((!g827) & (g869) & (g915) & (g2055) & (g2114) & (!g2056)) + ((!g827) & (g869) & (g915) & (g2055) & (g2114) & (g2056)) + ((g827) & (!g869) & (!g915) & (!g2055) & (g2114) & (!g2056)) + ((g827) & (!g869) & (!g915) & (!g2055) & (g2114) & (g2056)) + ((g827) & (!g869) & (!g915) & (g2055) & (!g2114) & (g2056)) + ((g827) & (!g869) & (!g915) & (g2055) & (g2114) & (!g2056)) + ((g827) & (!g869) & (g915) & (!g2055) & (!g2114) & (!g2056)) + ((g827) & (!g869) & (g915) & (!g2055) & (!g2114) & (g2056)) + ((g827) & (!g869) & (g915) & (g2055) & (!g2114) & (!g2056)) + ((g827) & (!g869) & (g915) & (g2055) & (g2114) & (g2056)) + ((g827) & (g869) & (!g915) & (!g2055) & (!g2114) & (g2056)) + ((g827) & (g869) & (!g915) & (!g2055) & (g2114) & (!g2056)) + ((g827) & (g869) & (!g915) & (g2055) & (!g2114) & (!g2056)) + ((g827) & (g869) & (!g915) & (g2055) & (!g2114) & (g2056)) + ((g827) & (g869) & (g915) & (!g2055) & (!g2114) & (!g2056)) + ((g827) & (g869) & (g915) & (!g2055) & (g2114) & (g2056)) + ((g827) & (g869) & (g915) & (g2055) & (g2114) & (!g2056)) + ((g827) & (g869) & (g915) & (g2055) & (g2114) & (g2056)));
	assign g7902 = (((!g3499) & (g4280) & (!g2116)) + ((!g3499) & (g4280) & (g2116)) + ((g3499) & (!g4280) & (g2116)) + ((g3499) & (g4280) & (g2116)));
	assign g2117 = (((!g827) & (!g877) & (!g917) & (!g2065) & (g2116) & (!g2066)) + ((!g827) & (!g877) & (!g917) & (!g2065) & (g2116) & (g2066)) + ((!g827) & (!g877) & (!g917) & (g2065) & (g2116) & (!g2066)) + ((!g827) & (!g877) & (!g917) & (g2065) & (g2116) & (g2066)) + ((!g827) & (!g877) & (g917) & (!g2065) & (g2116) & (!g2066)) + ((!g827) & (!g877) & (g917) & (!g2065) & (g2116) & (g2066)) + ((!g827) & (!g877) & (g917) & (g2065) & (g2116) & (!g2066)) + ((!g827) & (!g877) & (g917) & (g2065) & (g2116) & (g2066)) + ((!g827) & (g877) & (!g917) & (!g2065) & (g2116) & (!g2066)) + ((!g827) & (g877) & (!g917) & (!g2065) & (g2116) & (g2066)) + ((!g827) & (g877) & (!g917) & (g2065) & (g2116) & (!g2066)) + ((!g827) & (g877) & (!g917) & (g2065) & (g2116) & (g2066)) + ((!g827) & (g877) & (g917) & (!g2065) & (g2116) & (!g2066)) + ((!g827) & (g877) & (g917) & (!g2065) & (g2116) & (g2066)) + ((!g827) & (g877) & (g917) & (g2065) & (g2116) & (!g2066)) + ((!g827) & (g877) & (g917) & (g2065) & (g2116) & (g2066)) + ((g827) & (!g877) & (!g917) & (!g2065) & (g2116) & (!g2066)) + ((g827) & (!g877) & (!g917) & (!g2065) & (g2116) & (g2066)) + ((g827) & (!g877) & (!g917) & (g2065) & (!g2116) & (g2066)) + ((g827) & (!g877) & (!g917) & (g2065) & (g2116) & (!g2066)) + ((g827) & (!g877) & (g917) & (!g2065) & (!g2116) & (!g2066)) + ((g827) & (!g877) & (g917) & (!g2065) & (!g2116) & (g2066)) + ((g827) & (!g877) & (g917) & (g2065) & (!g2116) & (!g2066)) + ((g827) & (!g877) & (g917) & (g2065) & (g2116) & (g2066)) + ((g827) & (g877) & (!g917) & (!g2065) & (!g2116) & (g2066)) + ((g827) & (g877) & (!g917) & (!g2065) & (g2116) & (!g2066)) + ((g827) & (g877) & (!g917) & (g2065) & (!g2116) & (!g2066)) + ((g827) & (g877) & (!g917) & (g2065) & (!g2116) & (g2066)) + ((g827) & (g877) & (g917) & (!g2065) & (!g2116) & (!g2066)) + ((g827) & (g877) & (g917) & (!g2065) & (g2116) & (g2066)) + ((g827) & (g877) & (g917) & (g2065) & (g2116) & (!g2066)) + ((g827) & (g877) & (g917) & (g2065) & (g2116) & (g2066)));
	assign g7903 = (((!g2017) & (g6817) & (!g2118)) + ((!g2017) & (g6817) & (g2118)) + ((g2017) & (!g6817) & (g2118)) + ((g2017) & (g6817) & (g2118)));
	assign g2119 = (((!g827) & (!g885) & (!g919) & (!g2077) & (g2118) & (!g2078)) + ((!g827) & (!g885) & (!g919) & (!g2077) & (g2118) & (g2078)) + ((!g827) & (!g885) & (!g919) & (g2077) & (g2118) & (!g2078)) + ((!g827) & (!g885) & (!g919) & (g2077) & (g2118) & (g2078)) + ((!g827) & (!g885) & (g919) & (!g2077) & (g2118) & (!g2078)) + ((!g827) & (!g885) & (g919) & (!g2077) & (g2118) & (g2078)) + ((!g827) & (!g885) & (g919) & (g2077) & (g2118) & (!g2078)) + ((!g827) & (!g885) & (g919) & (g2077) & (g2118) & (g2078)) + ((!g827) & (g885) & (!g919) & (!g2077) & (g2118) & (!g2078)) + ((!g827) & (g885) & (!g919) & (!g2077) & (g2118) & (g2078)) + ((!g827) & (g885) & (!g919) & (g2077) & (g2118) & (!g2078)) + ((!g827) & (g885) & (!g919) & (g2077) & (g2118) & (g2078)) + ((!g827) & (g885) & (g919) & (!g2077) & (g2118) & (!g2078)) + ((!g827) & (g885) & (g919) & (!g2077) & (g2118) & (g2078)) + ((!g827) & (g885) & (g919) & (g2077) & (g2118) & (!g2078)) + ((!g827) & (g885) & (g919) & (g2077) & (g2118) & (g2078)) + ((g827) & (!g885) & (!g919) & (!g2077) & (g2118) & (!g2078)) + ((g827) & (!g885) & (!g919) & (!g2077) & (g2118) & (g2078)) + ((g827) & (!g885) & (!g919) & (g2077) & (!g2118) & (g2078)) + ((g827) & (!g885) & (!g919) & (g2077) & (g2118) & (!g2078)) + ((g827) & (!g885) & (g919) & (!g2077) & (!g2118) & (!g2078)) + ((g827) & (!g885) & (g919) & (!g2077) & (!g2118) & (g2078)) + ((g827) & (!g885) & (g919) & (g2077) & (!g2118) & (!g2078)) + ((g827) & (!g885) & (g919) & (g2077) & (g2118) & (g2078)) + ((g827) & (g885) & (!g919) & (!g2077) & (!g2118) & (g2078)) + ((g827) & (g885) & (!g919) & (!g2077) & (g2118) & (!g2078)) + ((g827) & (g885) & (!g919) & (g2077) & (!g2118) & (!g2078)) + ((g827) & (g885) & (!g919) & (g2077) & (!g2118) & (g2078)) + ((g827) & (g885) & (g919) & (!g2077) & (!g2118) & (!g2078)) + ((g827) & (g885) & (g919) & (!g2077) & (g2118) & (g2078)) + ((g827) & (g885) & (g919) & (g2077) & (g2118) & (!g2078)) + ((g827) & (g885) & (g919) & (g2077) & (g2118) & (g2078)));
	assign g7904 = (((!g3429) & (g4291) & (!g2120)) + ((!g3429) & (g4291) & (g2120)) + ((g3429) & (!g4291) & (g2120)) + ((g3429) & (g4291) & (g2120)));
	assign g2121 = (((!g827) & (!g893) & (!g921) & (!g2088) & (g2120) & (!g2089)) + ((!g827) & (!g893) & (!g921) & (!g2088) & (g2120) & (g2089)) + ((!g827) & (!g893) & (!g921) & (g2088) & (g2120) & (!g2089)) + ((!g827) & (!g893) & (!g921) & (g2088) & (g2120) & (g2089)) + ((!g827) & (!g893) & (g921) & (!g2088) & (g2120) & (!g2089)) + ((!g827) & (!g893) & (g921) & (!g2088) & (g2120) & (g2089)) + ((!g827) & (!g893) & (g921) & (g2088) & (g2120) & (!g2089)) + ((!g827) & (!g893) & (g921) & (g2088) & (g2120) & (g2089)) + ((!g827) & (g893) & (!g921) & (!g2088) & (g2120) & (!g2089)) + ((!g827) & (g893) & (!g921) & (!g2088) & (g2120) & (g2089)) + ((!g827) & (g893) & (!g921) & (g2088) & (g2120) & (!g2089)) + ((!g827) & (g893) & (!g921) & (g2088) & (g2120) & (g2089)) + ((!g827) & (g893) & (g921) & (!g2088) & (g2120) & (!g2089)) + ((!g827) & (g893) & (g921) & (!g2088) & (g2120) & (g2089)) + ((!g827) & (g893) & (g921) & (g2088) & (g2120) & (!g2089)) + ((!g827) & (g893) & (g921) & (g2088) & (g2120) & (g2089)) + ((g827) & (!g893) & (!g921) & (!g2088) & (g2120) & (!g2089)) + ((g827) & (!g893) & (!g921) & (!g2088) & (g2120) & (g2089)) + ((g827) & (!g893) & (!g921) & (g2088) & (!g2120) & (g2089)) + ((g827) & (!g893) & (!g921) & (g2088) & (g2120) & (!g2089)) + ((g827) & (!g893) & (g921) & (!g2088) & (!g2120) & (!g2089)) + ((g827) & (!g893) & (g921) & (!g2088) & (!g2120) & (g2089)) + ((g827) & (!g893) & (g921) & (g2088) & (!g2120) & (!g2089)) + ((g827) & (!g893) & (g921) & (g2088) & (g2120) & (g2089)) + ((g827) & (g893) & (!g921) & (!g2088) & (!g2120) & (g2089)) + ((g827) & (g893) & (!g921) & (!g2088) & (g2120) & (!g2089)) + ((g827) & (g893) & (!g921) & (g2088) & (!g2120) & (!g2089)) + ((g827) & (g893) & (!g921) & (g2088) & (!g2120) & (g2089)) + ((g827) & (g893) & (g921) & (!g2088) & (!g2120) & (!g2089)) + ((g827) & (g893) & (g921) & (!g2088) & (g2120) & (g2089)) + ((g827) & (g893) & (g921) & (g2088) & (g2120) & (!g2089)) + ((g827) & (g893) & (g921) & (g2088) & (g2120) & (g2089)));
	assign g2122 = (((!g827) & (!g871) & (!g923) & (!g1980) & (g1983) & (!g2058)) + ((!g827) & (!g871) & (!g923) & (!g1980) & (g1983) & (g2058)) + ((!g827) & (!g871) & (!g923) & (g1980) & (g1983) & (!g2058)) + ((!g827) & (!g871) & (!g923) & (g1980) & (g1983) & (g2058)) + ((!g827) & (!g871) & (g923) & (!g1980) & (g1983) & (!g2058)) + ((!g827) & (!g871) & (g923) & (!g1980) & (g1983) & (g2058)) + ((!g827) & (!g871) & (g923) & (g1980) & (g1983) & (!g2058)) + ((!g827) & (!g871) & (g923) & (g1980) & (g1983) & (g2058)) + ((!g827) & (g871) & (!g923) & (!g1980) & (g1983) & (!g2058)) + ((!g827) & (g871) & (!g923) & (!g1980) & (g1983) & (g2058)) + ((!g827) & (g871) & (!g923) & (g1980) & (g1983) & (!g2058)) + ((!g827) & (g871) & (!g923) & (g1980) & (g1983) & (g2058)) + ((!g827) & (g871) & (g923) & (!g1980) & (g1983) & (!g2058)) + ((!g827) & (g871) & (g923) & (!g1980) & (g1983) & (g2058)) + ((!g827) & (g871) & (g923) & (g1980) & (g1983) & (!g2058)) + ((!g827) & (g871) & (g923) & (g1980) & (g1983) & (g2058)) + ((g827) & (!g871) & (!g923) & (!g1980) & (g1983) & (!g2058)) + ((g827) & (!g871) & (!g923) & (!g1980) & (g1983) & (g2058)) + ((g827) & (!g871) & (!g923) & (g1980) & (!g1983) & (g2058)) + ((g827) & (!g871) & (!g923) & (g1980) & (g1983) & (!g2058)) + ((g827) & (!g871) & (g923) & (!g1980) & (!g1983) & (!g2058)) + ((g827) & (!g871) & (g923) & (!g1980) & (!g1983) & (g2058)) + ((g827) & (!g871) & (g923) & (g1980) & (!g1983) & (!g2058)) + ((g827) & (!g871) & (g923) & (g1980) & (g1983) & (g2058)) + ((g827) & (g871) & (!g923) & (!g1980) & (!g1983) & (g2058)) + ((g827) & (g871) & (!g923) & (!g1980) & (g1983) & (!g2058)) + ((g827) & (g871) & (!g923) & (g1980) & (!g1983) & (!g2058)) + ((g827) & (g871) & (!g923) & (g1980) & (!g1983) & (g2058)) + ((g827) & (g871) & (g923) & (!g1980) & (!g1983) & (!g2058)) + ((g827) & (g871) & (g923) & (!g1980) & (g1983) & (g2058)) + ((g827) & (g871) & (g923) & (g1980) & (g1983) & (!g2058)) + ((g827) & (g871) & (g923) & (g1980) & (g1983) & (g2058)));
	assign g7905 = (((!g3464) & (g4295) & (!g2123)) + ((!g3464) & (g4295) & (g2123)) + ((g3464) & (!g4295) & (g2123)) + ((g3464) & (g4295) & (g2123)));
	assign g2124 = (((!g827) & (!g879) & (!g925) & (!g2068) & (g2123) & (!g2069)) + ((!g827) & (!g879) & (!g925) & (!g2068) & (g2123) & (g2069)) + ((!g827) & (!g879) & (!g925) & (g2068) & (g2123) & (!g2069)) + ((!g827) & (!g879) & (!g925) & (g2068) & (g2123) & (g2069)) + ((!g827) & (!g879) & (g925) & (!g2068) & (g2123) & (!g2069)) + ((!g827) & (!g879) & (g925) & (!g2068) & (g2123) & (g2069)) + ((!g827) & (!g879) & (g925) & (g2068) & (g2123) & (!g2069)) + ((!g827) & (!g879) & (g925) & (g2068) & (g2123) & (g2069)) + ((!g827) & (g879) & (!g925) & (!g2068) & (g2123) & (!g2069)) + ((!g827) & (g879) & (!g925) & (!g2068) & (g2123) & (g2069)) + ((!g827) & (g879) & (!g925) & (g2068) & (g2123) & (!g2069)) + ((!g827) & (g879) & (!g925) & (g2068) & (g2123) & (g2069)) + ((!g827) & (g879) & (g925) & (!g2068) & (g2123) & (!g2069)) + ((!g827) & (g879) & (g925) & (!g2068) & (g2123) & (g2069)) + ((!g827) & (g879) & (g925) & (g2068) & (g2123) & (!g2069)) + ((!g827) & (g879) & (g925) & (g2068) & (g2123) & (g2069)) + ((g827) & (!g879) & (!g925) & (!g2068) & (g2123) & (!g2069)) + ((g827) & (!g879) & (!g925) & (!g2068) & (g2123) & (g2069)) + ((g827) & (!g879) & (!g925) & (g2068) & (!g2123) & (g2069)) + ((g827) & (!g879) & (!g925) & (g2068) & (g2123) & (!g2069)) + ((g827) & (!g879) & (g925) & (!g2068) & (!g2123) & (!g2069)) + ((g827) & (!g879) & (g925) & (!g2068) & (!g2123) & (g2069)) + ((g827) & (!g879) & (g925) & (g2068) & (!g2123) & (!g2069)) + ((g827) & (!g879) & (g925) & (g2068) & (g2123) & (g2069)) + ((g827) & (g879) & (!g925) & (!g2068) & (!g2123) & (g2069)) + ((g827) & (g879) & (!g925) & (!g2068) & (g2123) & (!g2069)) + ((g827) & (g879) & (!g925) & (g2068) & (!g2123) & (!g2069)) + ((g827) & (g879) & (!g925) & (g2068) & (!g2123) & (g2069)) + ((g827) & (g879) & (g925) & (!g2068) & (!g2123) & (!g2069)) + ((g827) & (g879) & (g925) & (!g2068) & (g2123) & (g2069)) + ((g827) & (g879) & (g925) & (g2068) & (g2123) & (!g2069)) + ((g827) & (g879) & (g925) & (g2068) & (g2123) & (g2069)));
	assign g7906 = (((!g3429) & (g4304) & (!g2125)) + ((!g3429) & (g4304) & (g2125)) + ((g3429) & (!g4304) & (g2125)) + ((g3429) & (g4304) & (g2125)));
	assign g2126 = (((!g827) & (!g887) & (!g927) & (!g2080) & (g2125) & (!g2081)) + ((!g827) & (!g887) & (!g927) & (!g2080) & (g2125) & (g2081)) + ((!g827) & (!g887) & (!g927) & (g2080) & (g2125) & (!g2081)) + ((!g827) & (!g887) & (!g927) & (g2080) & (g2125) & (g2081)) + ((!g827) & (!g887) & (g927) & (!g2080) & (g2125) & (!g2081)) + ((!g827) & (!g887) & (g927) & (!g2080) & (g2125) & (g2081)) + ((!g827) & (!g887) & (g927) & (g2080) & (g2125) & (!g2081)) + ((!g827) & (!g887) & (g927) & (g2080) & (g2125) & (g2081)) + ((!g827) & (g887) & (!g927) & (!g2080) & (g2125) & (!g2081)) + ((!g827) & (g887) & (!g927) & (!g2080) & (g2125) & (g2081)) + ((!g827) & (g887) & (!g927) & (g2080) & (g2125) & (!g2081)) + ((!g827) & (g887) & (!g927) & (g2080) & (g2125) & (g2081)) + ((!g827) & (g887) & (g927) & (!g2080) & (g2125) & (!g2081)) + ((!g827) & (g887) & (g927) & (!g2080) & (g2125) & (g2081)) + ((!g827) & (g887) & (g927) & (g2080) & (g2125) & (!g2081)) + ((!g827) & (g887) & (g927) & (g2080) & (g2125) & (g2081)) + ((g827) & (!g887) & (!g927) & (!g2080) & (g2125) & (!g2081)) + ((g827) & (!g887) & (!g927) & (!g2080) & (g2125) & (g2081)) + ((g827) & (!g887) & (!g927) & (g2080) & (!g2125) & (g2081)) + ((g827) & (!g887) & (!g927) & (g2080) & (g2125) & (!g2081)) + ((g827) & (!g887) & (g927) & (!g2080) & (!g2125) & (!g2081)) + ((g827) & (!g887) & (g927) & (!g2080) & (!g2125) & (g2081)) + ((g827) & (!g887) & (g927) & (g2080) & (!g2125) & (!g2081)) + ((g827) & (!g887) & (g927) & (g2080) & (g2125) & (g2081)) + ((g827) & (g887) & (!g927) & (!g2080) & (!g2125) & (g2081)) + ((g827) & (g887) & (!g927) & (!g2080) & (g2125) & (!g2081)) + ((g827) & (g887) & (!g927) & (g2080) & (!g2125) & (!g2081)) + ((g827) & (g887) & (!g927) & (g2080) & (!g2125) & (g2081)) + ((g827) & (g887) & (g927) & (!g2080) & (!g2125) & (!g2081)) + ((g827) & (g887) & (g927) & (!g2080) & (g2125) & (g2081)) + ((g827) & (g887) & (g927) & (g2080) & (g2125) & (!g2081)) + ((g827) & (g887) & (g927) & (g2080) & (g2125) & (g2081)));
	assign g7907 = (((!g2017) & (g6811) & (!g2127)) + ((!g2017) & (g6811) & (g2127)) + ((g2017) & (!g6811) & (g2127)) + ((g2017) & (g6811) & (g2127)));
	assign g2128 = (((!g827) & (!g895) & (!g929) & (!g2091) & (g2127) & (!g2092)) + ((!g827) & (!g895) & (!g929) & (!g2091) & (g2127) & (g2092)) + ((!g827) & (!g895) & (!g929) & (g2091) & (g2127) & (!g2092)) + ((!g827) & (!g895) & (!g929) & (g2091) & (g2127) & (g2092)) + ((!g827) & (!g895) & (g929) & (!g2091) & (g2127) & (!g2092)) + ((!g827) & (!g895) & (g929) & (!g2091) & (g2127) & (g2092)) + ((!g827) & (!g895) & (g929) & (g2091) & (g2127) & (!g2092)) + ((!g827) & (!g895) & (g929) & (g2091) & (g2127) & (g2092)) + ((!g827) & (g895) & (!g929) & (!g2091) & (g2127) & (!g2092)) + ((!g827) & (g895) & (!g929) & (!g2091) & (g2127) & (g2092)) + ((!g827) & (g895) & (!g929) & (g2091) & (g2127) & (!g2092)) + ((!g827) & (g895) & (!g929) & (g2091) & (g2127) & (g2092)) + ((!g827) & (g895) & (g929) & (!g2091) & (g2127) & (!g2092)) + ((!g827) & (g895) & (g929) & (!g2091) & (g2127) & (g2092)) + ((!g827) & (g895) & (g929) & (g2091) & (g2127) & (!g2092)) + ((!g827) & (g895) & (g929) & (g2091) & (g2127) & (g2092)) + ((g827) & (!g895) & (!g929) & (!g2091) & (g2127) & (!g2092)) + ((g827) & (!g895) & (!g929) & (!g2091) & (g2127) & (g2092)) + ((g827) & (!g895) & (!g929) & (g2091) & (!g2127) & (g2092)) + ((g827) & (!g895) & (!g929) & (g2091) & (g2127) & (!g2092)) + ((g827) & (!g895) & (g929) & (!g2091) & (!g2127) & (!g2092)) + ((g827) & (!g895) & (g929) & (!g2091) & (!g2127) & (g2092)) + ((g827) & (!g895) & (g929) & (g2091) & (!g2127) & (!g2092)) + ((g827) & (!g895) & (g929) & (g2091) & (g2127) & (g2092)) + ((g827) & (g895) & (!g929) & (!g2091) & (!g2127) & (g2092)) + ((g827) & (g895) & (!g929) & (!g2091) & (g2127) & (!g2092)) + ((g827) & (g895) & (!g929) & (g2091) & (!g2127) & (!g2092)) + ((g827) & (g895) & (!g929) & (g2091) & (!g2127) & (g2092)) + ((g827) & (g895) & (g929) & (!g2091) & (!g2127) & (!g2092)) + ((g827) & (g895) & (g929) & (!g2091) & (g2127) & (g2092)) + ((g827) & (g895) & (g929) & (g2091) & (g2127) & (!g2092)) + ((g827) & (g895) & (g929) & (g2091) & (g2127) & (g2092)));
	assign g7908 = (((!g3429) & (g4309) & (!g2129)) + ((!g3429) & (g4309) & (g2129)) + ((g3429) & (!g4309) & (g2129)) + ((g3429) & (g4309) & (g2129)));
	assign g7909 = (((!g3464) & (g4312) & (!g2130)) + ((!g3464) & (g4312) & (g2130)) + ((g3464) & (!g4312) & (g2130)) + ((g3464) & (g4312) & (g2130)));
	assign g2131 = (((!g2097) & (!g2098) & (!g2099) & (!g2129) & (g2130)) + ((!g2097) & (!g2098) & (!g2099) & (g2129) & (!g2130)) + ((!g2097) & (!g2098) & (g2099) & (!g2129) & (g2130)) + ((!g2097) & (!g2098) & (g2099) & (g2129) & (!g2130)) + ((!g2097) & (g2098) & (!g2099) & (!g2129) & (g2130)) + ((!g2097) & (g2098) & (!g2099) & (g2129) & (!g2130)) + ((!g2097) & (g2098) & (g2099) & (!g2129) & (!g2130)) + ((!g2097) & (g2098) & (g2099) & (g2129) & (g2130)) + ((g2097) & (!g2098) & (!g2099) & (!g2129) & (g2130)) + ((g2097) & (!g2098) & (!g2099) & (g2129) & (!g2130)) + ((g2097) & (!g2098) & (g2099) & (!g2129) & (!g2130)) + ((g2097) & (!g2098) & (g2099) & (g2129) & (g2130)) + ((g2097) & (g2098) & (!g2099) & (!g2129) & (!g2130)) + ((g2097) & (g2098) & (!g2099) & (g2129) & (g2130)) + ((g2097) & (g2098) & (g2099) & (!g2129) & (!g2130)) + ((g2097) & (g2098) & (g2099) & (g2129) & (g2130)));
	assign g2132 = (((!g2050) & (!g2051) & (!g2052) & (g2100) & (g2101)) + ((!g2050) & (!g2051) & (g2052) & (g2100) & (g2101)) + ((!g2050) & (g2051) & (!g2052) & (g2100) & (g2101)) + ((!g2050) & (g2051) & (g2052) & (!g2100) & (g2101)) + ((!g2050) & (g2051) & (g2052) & (g2100) & (!g2101)) + ((!g2050) & (g2051) & (g2052) & (g2100) & (g2101)) + ((g2050) & (!g2051) & (!g2052) & (g2100) & (g2101)) + ((g2050) & (!g2051) & (g2052) & (!g2100) & (g2101)) + ((g2050) & (!g2051) & (g2052) & (g2100) & (!g2101)) + ((g2050) & (!g2051) & (g2052) & (g2100) & (g2101)) + ((g2050) & (g2051) & (!g2052) & (!g2100) & (g2101)) + ((g2050) & (g2051) & (!g2052) & (g2100) & (!g2101)) + ((g2050) & (g2051) & (!g2052) & (g2100) & (g2101)) + ((g2050) & (g2051) & (g2052) & (!g2100) & (g2101)) + ((g2050) & (g2051) & (g2052) & (g2100) & (!g2101)) + ((g2050) & (g2051) & (g2052) & (g2100) & (g2101)));
	assign g7910 = (((!g3429) & (g4316) & (!g2133)) + ((!g3429) & (g4316) & (g2133)) + ((g3429) & (!g4316) & (g2133)) + ((g3429) & (g4316) & (g2133)));
	assign g7911 = (((!g3499) & (g4319) & (!g2134)) + ((!g3499) & (g4319) & (g2134)) + ((g3499) & (!g4319) & (g2134)) + ((g3499) & (g4319) & (g2134)));
	assign g2135 = (((!g867) & (!g907) & (g1979) & (g1982) & (g2053)) + ((!g867) & (g907) & (!g1979) & (g1982) & (!g2053)) + ((!g867) & (g907) & (!g1979) & (g1982) & (g2053)) + ((!g867) & (g907) & (g1979) & (!g1982) & (g2053)) + ((!g867) & (g907) & (g1979) & (g1982) & (!g2053)) + ((!g867) & (g907) & (g1979) & (g1982) & (g2053)) + ((g867) & (!g907) & (!g1979) & (g1982) & (g2053)) + ((g867) & (!g907) & (g1979) & (g1982) & (!g2053)) + ((g867) & (!g907) & (g1979) & (g1982) & (g2053)) + ((g867) & (g907) & (!g1979) & (!g1982) & (g2053)) + ((g867) & (g907) & (!g1979) & (g1982) & (!g2053)) + ((g867) & (g907) & (!g1979) & (g1982) & (g2053)) + ((g867) & (g907) & (g1979) & (!g1982) & (!g2053)) + ((g867) & (g907) & (g1979) & (!g1982) & (g2053)) + ((g867) & (g907) & (g1979) & (g1982) & (!g2053)) + ((g867) & (g907) & (g1979) & (g1982) & (g2053)));
	assign g2136 = (((!g827) & (!g934) & (g1984) & (!g2135)) + ((!g827) & (!g934) & (g1984) & (g2135)) + ((!g827) & (g934) & (g1984) & (!g2135)) + ((!g827) & (g934) & (g1984) & (g2135)) + ((g827) & (!g934) & (!g1984) & (g2135)) + ((g827) & (!g934) & (g1984) & (!g2135)) + ((g827) & (g934) & (!g1984) & (!g2135)) + ((g827) & (g934) & (g1984) & (g2135)));
	assign g7912 = (((!g3464) & (g4323) & (!g2137)) + ((!g3464) & (g4323) & (g2137)) + ((g3464) & (!g4323) & (g2137)) + ((g3464) & (g4323) & (g2137)));
	assign g2138 = (((!g869) & (!g915) & (g2055) & (g2114) & (g2056)) + ((!g869) & (g915) & (!g2055) & (g2114) & (!g2056)) + ((!g869) & (g915) & (!g2055) & (g2114) & (g2056)) + ((!g869) & (g915) & (g2055) & (!g2114) & (g2056)) + ((!g869) & (g915) & (g2055) & (g2114) & (!g2056)) + ((!g869) & (g915) & (g2055) & (g2114) & (g2056)) + ((g869) & (!g915) & (!g2055) & (g2114) & (g2056)) + ((g869) & (!g915) & (g2055) & (g2114) & (!g2056)) + ((g869) & (!g915) & (g2055) & (g2114) & (g2056)) + ((g869) & (g915) & (!g2055) & (!g2114) & (g2056)) + ((g869) & (g915) & (!g2055) & (g2114) & (!g2056)) + ((g869) & (g915) & (!g2055) & (g2114) & (g2056)) + ((g869) & (g915) & (g2055) & (!g2114) & (!g2056)) + ((g869) & (g915) & (g2055) & (!g2114) & (g2056)) + ((g869) & (g915) & (g2055) & (g2114) & (!g2056)) + ((g869) & (g915) & (g2055) & (g2114) & (g2056)));
	assign g2139 = (((!g827) & (!g936) & (g2137) & (!g2138)) + ((!g827) & (!g936) & (g2137) & (g2138)) + ((!g827) & (g936) & (g2137) & (!g2138)) + ((!g827) & (g936) & (g2137) & (g2138)) + ((g827) & (!g936) & (!g2137) & (g2138)) + ((g827) & (!g936) & (g2137) & (!g2138)) + ((g827) & (g936) & (!g2137) & (!g2138)) + ((g827) & (g936) & (g2137) & (g2138)));
	assign g2140 = (((!g871) & (!g923) & (g1980) & (g1983) & (g2058)) + ((!g871) & (g923) & (!g1980) & (g1983) & (!g2058)) + ((!g871) & (g923) & (!g1980) & (g1983) & (g2058)) + ((!g871) & (g923) & (g1980) & (!g1983) & (g2058)) + ((!g871) & (g923) & (g1980) & (g1983) & (!g2058)) + ((!g871) & (g923) & (g1980) & (g1983) & (g2058)) + ((g871) & (!g923) & (!g1980) & (g1983) & (g2058)) + ((g871) & (!g923) & (g1980) & (g1983) & (!g2058)) + ((g871) & (!g923) & (g1980) & (g1983) & (g2058)) + ((g871) & (g923) & (!g1980) & (!g1983) & (g2058)) + ((g871) & (g923) & (!g1980) & (g1983) & (!g2058)) + ((g871) & (g923) & (!g1980) & (g1983) & (g2058)) + ((g871) & (g923) & (g1980) & (!g1983) & (!g2058)) + ((g871) & (g923) & (g1980) & (!g1983) & (g2058)) + ((g871) & (g923) & (g1980) & (g1983) & (!g2058)) + ((g871) & (g923) & (g1980) & (g1983) & (g2058)));
	assign g2141 = (((!g827) & (!g938) & (g1985) & (!g2140)) + ((!g827) & (!g938) & (g1985) & (g2140)) + ((!g827) & (g938) & (g1985) & (!g2140)) + ((!g827) & (g938) & (g1985) & (g2140)) + ((g827) & (!g938) & (!g1985) & (g2140)) + ((g827) & (!g938) & (g1985) & (!g2140)) + ((g827) & (g938) & (!g1985) & (!g2140)) + ((g827) & (g938) & (g1985) & (g2140)));
	assign g2142 = (((!g873) & (!g901) & (g1941) & (g1944) & (g2060)) + ((!g873) & (g901) & (!g1941) & (g1944) & (!g2060)) + ((!g873) & (g901) & (!g1941) & (g1944) & (g2060)) + ((!g873) & (g901) & (g1941) & (!g1944) & (g2060)) + ((!g873) & (g901) & (g1941) & (g1944) & (!g2060)) + ((!g873) & (g901) & (g1941) & (g1944) & (g2060)) + ((g873) & (!g901) & (!g1941) & (g1944) & (g2060)) + ((g873) & (!g901) & (g1941) & (g1944) & (!g2060)) + ((g873) & (!g901) & (g1941) & (g1944) & (g2060)) + ((g873) & (g901) & (!g1941) & (!g1944) & (g2060)) + ((g873) & (g901) & (!g1941) & (g1944) & (!g2060)) + ((g873) & (g901) & (!g1941) & (g1944) & (g2060)) + ((g873) & (g901) & (g1941) & (!g1944) & (!g2060)) + ((g873) & (g901) & (g1941) & (!g1944) & (g2060)) + ((g873) & (g901) & (g1941) & (g1944) & (!g2060)) + ((g873) & (g901) & (g1941) & (g1944) & (g2060)));
	assign g2143 = (((!g827) & (!g940) & (g1946) & (!g2142)) + ((!g827) & (!g940) & (g1946) & (g2142)) + ((!g827) & (g940) & (g1946) & (!g2142)) + ((!g827) & (g940) & (g1946) & (g2142)) + ((g827) & (!g940) & (!g1946) & (g2142)) + ((g827) & (!g940) & (g1946) & (!g2142)) + ((g827) & (g940) & (!g1946) & (!g2142)) + ((g827) & (g940) & (g1946) & (g2142)));
	assign g7913 = (((!g2017) & (g6782) & (!g2144)) + ((!g2017) & (g6782) & (g2144)) + ((g2017) & (!g6782) & (g2144)) + ((g2017) & (g6782) & (g2144)));
	assign g2145 = (((!g875) & (!g909) & (g2062) & (g2108) & (g2063)) + ((!g875) & (g909) & (!g2062) & (g2108) & (!g2063)) + ((!g875) & (g909) & (!g2062) & (g2108) & (g2063)) + ((!g875) & (g909) & (g2062) & (!g2108) & (g2063)) + ((!g875) & (g909) & (g2062) & (g2108) & (!g2063)) + ((!g875) & (g909) & (g2062) & (g2108) & (g2063)) + ((g875) & (!g909) & (!g2062) & (g2108) & (g2063)) + ((g875) & (!g909) & (g2062) & (g2108) & (!g2063)) + ((g875) & (!g909) & (g2062) & (g2108) & (g2063)) + ((g875) & (g909) & (!g2062) & (!g2108) & (g2063)) + ((g875) & (g909) & (!g2062) & (g2108) & (!g2063)) + ((g875) & (g909) & (!g2062) & (g2108) & (g2063)) + ((g875) & (g909) & (g2062) & (!g2108) & (!g2063)) + ((g875) & (g909) & (g2062) & (!g2108) & (g2063)) + ((g875) & (g909) & (g2062) & (g2108) & (!g2063)) + ((g875) & (g909) & (g2062) & (g2108) & (g2063)));
	assign g2146 = (((!g827) & (!g942) & (g2144) & (!g2145)) + ((!g827) & (!g942) & (g2144) & (g2145)) + ((!g827) & (g942) & (g2144) & (!g2145)) + ((!g827) & (g942) & (g2144) & (g2145)) + ((g827) & (!g942) & (!g2144) & (g2145)) + ((g827) & (!g942) & (g2144) & (!g2145)) + ((g827) & (g942) & (!g2144) & (!g2145)) + ((g827) & (g942) & (g2144) & (g2145)));
	assign g7914 = (((!g3499) & (g4330) & (!g2147)) + ((!g3499) & (g4330) & (g2147)) + ((g3499) & (!g4330) & (g2147)) + ((g3499) & (g4330) & (g2147)));
	assign g2148 = (((!g877) & (!g917) & (g2065) & (g2116) & (g2066)) + ((!g877) & (g917) & (!g2065) & (g2116) & (!g2066)) + ((!g877) & (g917) & (!g2065) & (g2116) & (g2066)) + ((!g877) & (g917) & (g2065) & (!g2116) & (g2066)) + ((!g877) & (g917) & (g2065) & (g2116) & (!g2066)) + ((!g877) & (g917) & (g2065) & (g2116) & (g2066)) + ((g877) & (!g917) & (!g2065) & (g2116) & (g2066)) + ((g877) & (!g917) & (g2065) & (g2116) & (!g2066)) + ((g877) & (!g917) & (g2065) & (g2116) & (g2066)) + ((g877) & (g917) & (!g2065) & (!g2116) & (g2066)) + ((g877) & (g917) & (!g2065) & (g2116) & (!g2066)) + ((g877) & (g917) & (!g2065) & (g2116) & (g2066)) + ((g877) & (g917) & (g2065) & (!g2116) & (!g2066)) + ((g877) & (g917) & (g2065) & (!g2116) & (g2066)) + ((g877) & (g917) & (g2065) & (g2116) & (!g2066)) + ((g877) & (g917) & (g2065) & (g2116) & (g2066)));
	assign g2149 = (((!g827) & (!g944) & (g2147) & (!g2148)) + ((!g827) & (!g944) & (g2147) & (g2148)) + ((!g827) & (g944) & (g2147) & (!g2148)) + ((!g827) & (g944) & (g2147) & (g2148)) + ((g827) & (!g944) & (!g2147) & (g2148)) + ((g827) & (!g944) & (g2147) & (!g2148)) + ((g827) & (g944) & (!g2147) & (!g2148)) + ((g827) & (g944) & (g2147) & (g2148)));
	assign g7915 = (((!g3464) & (g4334) & (!g2150)) + ((!g3464) & (g4334) & (g2150)) + ((g3464) & (!g4334) & (g2150)) + ((g3464) & (g4334) & (g2150)));
	assign g2151 = (((!g879) & (!g925) & (g2068) & (g2123) & (g2069)) + ((!g879) & (g925) & (!g2068) & (g2123) & (!g2069)) + ((!g879) & (g925) & (!g2068) & (g2123) & (g2069)) + ((!g879) & (g925) & (g2068) & (!g2123) & (g2069)) + ((!g879) & (g925) & (g2068) & (g2123) & (!g2069)) + ((!g879) & (g925) & (g2068) & (g2123) & (g2069)) + ((g879) & (!g925) & (!g2068) & (g2123) & (g2069)) + ((g879) & (!g925) & (g2068) & (g2123) & (!g2069)) + ((g879) & (!g925) & (g2068) & (g2123) & (g2069)) + ((g879) & (g925) & (!g2068) & (!g2123) & (g2069)) + ((g879) & (g925) & (!g2068) & (g2123) & (!g2069)) + ((g879) & (g925) & (!g2068) & (g2123) & (g2069)) + ((g879) & (g925) & (g2068) & (!g2123) & (!g2069)) + ((g879) & (g925) & (g2068) & (!g2123) & (g2069)) + ((g879) & (g925) & (g2068) & (g2123) & (!g2069)) + ((g879) & (g925) & (g2068) & (g2123) & (g2069)));
	assign g2152 = (((!g827) & (!g946) & (g2150) & (!g2151)) + ((!g827) & (!g946) & (g2150) & (g2151)) + ((!g827) & (g946) & (g2150) & (!g2151)) + ((!g827) & (g946) & (g2150) & (g2151)) + ((g827) & (!g946) & (!g2150) & (g2151)) + ((g827) & (!g946) & (g2150) & (!g2151)) + ((g827) & (g946) & (!g2150) & (!g2151)) + ((g827) & (g946) & (g2150) & (g2151)));
	assign g7916 = (((!g3499) & (g4338) & (!g2153)) + ((!g3499) & (g4338) & (g2153)) + ((g3499) & (!g4338) & (g2153)) + ((g3499) & (g4338) & (g2153)));
	assign g2154 = (((!g881) & (!g903) & (g2071) & (g2104) & (g2072)) + ((!g881) & (g903) & (!g2071) & (g2104) & (!g2072)) + ((!g881) & (g903) & (!g2071) & (g2104) & (g2072)) + ((!g881) & (g903) & (g2071) & (!g2104) & (g2072)) + ((!g881) & (g903) & (g2071) & (g2104) & (!g2072)) + ((!g881) & (g903) & (g2071) & (g2104) & (g2072)) + ((g881) & (!g903) & (!g2071) & (g2104) & (g2072)) + ((g881) & (!g903) & (g2071) & (g2104) & (!g2072)) + ((g881) & (!g903) & (g2071) & (g2104) & (g2072)) + ((g881) & (g903) & (!g2071) & (!g2104) & (g2072)) + ((g881) & (g903) & (!g2071) & (g2104) & (!g2072)) + ((g881) & (g903) & (!g2071) & (g2104) & (g2072)) + ((g881) & (g903) & (g2071) & (!g2104) & (!g2072)) + ((g881) & (g903) & (g2071) & (!g2104) & (g2072)) + ((g881) & (g903) & (g2071) & (g2104) & (!g2072)) + ((g881) & (g903) & (g2071) & (g2104) & (g2072)));
	assign g2155 = (((!g827) & (!g948) & (g2153) & (!g2154)) + ((!g827) & (!g948) & (g2153) & (g2154)) + ((!g827) & (g948) & (g2153) & (!g2154)) + ((!g827) & (g948) & (g2153) & (g2154)) + ((g827) & (!g948) & (!g2153) & (g2154)) + ((g827) & (!g948) & (g2153) & (!g2154)) + ((g827) & (g948) & (!g2153) & (!g2154)) + ((g827) & (g948) & (g2153) & (g2154)));
	assign g7917 = (((!g3464) & (g4343) & (!g2156)) + ((!g3464) & (g4343) & (g2156)) + ((g3464) & (!g4343) & (g2156)) + ((g3464) & (g4343) & (g2156)));
	assign g2157 = (((!g883) & (!g911) & (g2074) & (g2110) & (g2075)) + ((!g883) & (g911) & (!g2074) & (g2110) & (!g2075)) + ((!g883) & (g911) & (!g2074) & (g2110) & (g2075)) + ((!g883) & (g911) & (g2074) & (!g2110) & (g2075)) + ((!g883) & (g911) & (g2074) & (g2110) & (!g2075)) + ((!g883) & (g911) & (g2074) & (g2110) & (g2075)) + ((g883) & (!g911) & (!g2074) & (g2110) & (g2075)) + ((g883) & (!g911) & (g2074) & (g2110) & (!g2075)) + ((g883) & (!g911) & (g2074) & (g2110) & (g2075)) + ((g883) & (g911) & (!g2074) & (!g2110) & (g2075)) + ((g883) & (g911) & (!g2074) & (g2110) & (!g2075)) + ((g883) & (g911) & (!g2074) & (g2110) & (g2075)) + ((g883) & (g911) & (g2074) & (!g2110) & (!g2075)) + ((g883) & (g911) & (g2074) & (!g2110) & (g2075)) + ((g883) & (g911) & (g2074) & (g2110) & (!g2075)) + ((g883) & (g911) & (g2074) & (g2110) & (g2075)));
	assign g2158 = (((!g827) & (!g950) & (g2156) & (!g2157)) + ((!g827) & (!g950) & (g2156) & (g2157)) + ((!g827) & (g950) & (g2156) & (!g2157)) + ((!g827) & (g950) & (g2156) & (g2157)) + ((g827) & (!g950) & (!g2156) & (g2157)) + ((g827) & (!g950) & (g2156) & (!g2157)) + ((g827) & (g950) & (!g2156) & (!g2157)) + ((g827) & (g950) & (g2156) & (g2157)));
	assign g7918 = (((!g2017) & (g6776) & (!g2159)) + ((!g2017) & (g6776) & (g2159)) + ((g2017) & (!g6776) & (g2159)) + ((g2017) & (g6776) & (g2159)));
	assign g2160 = (((!g885) & (!g919) & (g2077) & (g2118) & (g2078)) + ((!g885) & (g919) & (!g2077) & (g2118) & (!g2078)) + ((!g885) & (g919) & (!g2077) & (g2118) & (g2078)) + ((!g885) & (g919) & (g2077) & (!g2118) & (g2078)) + ((!g885) & (g919) & (g2077) & (g2118) & (!g2078)) + ((!g885) & (g919) & (g2077) & (g2118) & (g2078)) + ((g885) & (!g919) & (!g2077) & (g2118) & (g2078)) + ((g885) & (!g919) & (g2077) & (g2118) & (!g2078)) + ((g885) & (!g919) & (g2077) & (g2118) & (g2078)) + ((g885) & (g919) & (!g2077) & (!g2118) & (g2078)) + ((g885) & (g919) & (!g2077) & (g2118) & (!g2078)) + ((g885) & (g919) & (!g2077) & (g2118) & (g2078)) + ((g885) & (g919) & (g2077) & (!g2118) & (!g2078)) + ((g885) & (g919) & (g2077) & (!g2118) & (g2078)) + ((g885) & (g919) & (g2077) & (g2118) & (!g2078)) + ((g885) & (g919) & (g2077) & (g2118) & (g2078)));
	assign g2161 = (((!g827) & (!g952) & (g2159) & (!g2160)) + ((!g827) & (!g952) & (g2159) & (g2160)) + ((!g827) & (g952) & (g2159) & (!g2160)) + ((!g827) & (g952) & (g2159) & (g2160)) + ((g827) & (!g952) & (!g2159) & (g2160)) + ((g827) & (!g952) & (g2159) & (!g2160)) + ((g827) & (g952) & (!g2159) & (!g2160)) + ((g827) & (g952) & (g2159) & (g2160)));
	assign g7919 = (((!g3429) & (g4351) & (!g2162)) + ((!g3429) & (g4351) & (g2162)) + ((g3429) & (!g4351) & (g2162)) + ((g3429) & (g4351) & (g2162)));
	assign g2163 = (((!g887) & (!g927) & (g2080) & (g2125) & (g2081)) + ((!g887) & (g927) & (!g2080) & (g2125) & (!g2081)) + ((!g887) & (g927) & (!g2080) & (g2125) & (g2081)) + ((!g887) & (g927) & (g2080) & (!g2125) & (g2081)) + ((!g887) & (g927) & (g2080) & (g2125) & (!g2081)) + ((!g887) & (g927) & (g2080) & (g2125) & (g2081)) + ((g887) & (!g927) & (!g2080) & (g2125) & (g2081)) + ((g887) & (!g927) & (g2080) & (g2125) & (!g2081)) + ((g887) & (!g927) & (g2080) & (g2125) & (g2081)) + ((g887) & (g927) & (!g2080) & (!g2125) & (g2081)) + ((g887) & (g927) & (!g2080) & (g2125) & (!g2081)) + ((g887) & (g927) & (!g2080) & (g2125) & (g2081)) + ((g887) & (g927) & (g2080) & (!g2125) & (!g2081)) + ((g887) & (g927) & (g2080) & (!g2125) & (g2081)) + ((g887) & (g927) & (g2080) & (g2125) & (!g2081)) + ((g887) & (g927) & (g2080) & (g2125) & (g2081)));
	assign g2164 = (((!g827) & (!g954) & (g2162) & (!g2163)) + ((!g827) & (!g954) & (g2162) & (g2163)) + ((!g827) & (g954) & (g2162) & (!g2163)) + ((!g827) & (g954) & (g2162) & (g2163)) + ((g827) & (!g954) & (!g2162) & (g2163)) + ((g827) & (!g954) & (g2162) & (!g2163)) + ((g827) & (g954) & (!g2162) & (!g2163)) + ((g827) & (g954) & (g2162) & (g2163)));
	assign g2165 = (((!g889) & (!g905) & (g1942) & (g1945) & (g2083)) + ((!g889) & (g905) & (!g1942) & (g1945) & (!g2083)) + ((!g889) & (g905) & (!g1942) & (g1945) & (g2083)) + ((!g889) & (g905) & (g1942) & (!g1945) & (g2083)) + ((!g889) & (g905) & (g1942) & (g1945) & (!g2083)) + ((!g889) & (g905) & (g1942) & (g1945) & (g2083)) + ((g889) & (!g905) & (!g1942) & (g1945) & (g2083)) + ((g889) & (!g905) & (g1942) & (g1945) & (!g2083)) + ((g889) & (!g905) & (g1942) & (g1945) & (g2083)) + ((g889) & (g905) & (!g1942) & (!g1945) & (g2083)) + ((g889) & (g905) & (!g1942) & (g1945) & (!g2083)) + ((g889) & (g905) & (!g1942) & (g1945) & (g2083)) + ((g889) & (g905) & (g1942) & (!g1945) & (!g2083)) + ((g889) & (g905) & (g1942) & (!g1945) & (g2083)) + ((g889) & (g905) & (g1942) & (g1945) & (!g2083)) + ((g889) & (g905) & (g1942) & (g1945) & (g2083)));
	assign g2166 = (((!g827) & (!g956) & (g1947) & (!g2165)) + ((!g827) & (!g956) & (g1947) & (g2165)) + ((!g827) & (g956) & (g1947) & (!g2165)) + ((!g827) & (g956) & (g1947) & (g2165)) + ((g827) & (!g956) & (!g1947) & (g2165)) + ((g827) & (!g956) & (g1947) & (!g2165)) + ((g827) & (g956) & (!g1947) & (!g2165)) + ((g827) & (g956) & (g1947) & (g2165)));
	assign g7920 = (((!g3499) & (g4355) & (!g2167)) + ((!g3499) & (g4355) & (g2167)) + ((g3499) & (!g4355) & (g2167)) + ((g3499) & (g4355) & (g2167)));
	assign g2168 = (((!g891) & (!g913) & (g2085) & (g2112) & (g2086)) + ((!g891) & (g913) & (!g2085) & (g2112) & (!g2086)) + ((!g891) & (g913) & (!g2085) & (g2112) & (g2086)) + ((!g891) & (g913) & (g2085) & (!g2112) & (g2086)) + ((!g891) & (g913) & (g2085) & (g2112) & (!g2086)) + ((!g891) & (g913) & (g2085) & (g2112) & (g2086)) + ((g891) & (!g913) & (!g2085) & (g2112) & (g2086)) + ((g891) & (!g913) & (g2085) & (g2112) & (!g2086)) + ((g891) & (!g913) & (g2085) & (g2112) & (g2086)) + ((g891) & (g913) & (!g2085) & (!g2112) & (g2086)) + ((g891) & (g913) & (!g2085) & (g2112) & (!g2086)) + ((g891) & (g913) & (!g2085) & (g2112) & (g2086)) + ((g891) & (g913) & (g2085) & (!g2112) & (!g2086)) + ((g891) & (g913) & (g2085) & (!g2112) & (g2086)) + ((g891) & (g913) & (g2085) & (g2112) & (!g2086)) + ((g891) & (g913) & (g2085) & (g2112) & (g2086)));
	assign g2169 = (((!g827) & (!g958) & (g2167) & (!g2168)) + ((!g827) & (!g958) & (g2167) & (g2168)) + ((!g827) & (g958) & (g2167) & (!g2168)) + ((!g827) & (g958) & (g2167) & (g2168)) + ((g827) & (!g958) & (!g2167) & (g2168)) + ((g827) & (!g958) & (g2167) & (!g2168)) + ((g827) & (g958) & (!g2167) & (!g2168)) + ((g827) & (g958) & (g2167) & (g2168)));
	assign g7921 = (((!g3429) & (g4360) & (!g2170)) + ((!g3429) & (g4360) & (g2170)) + ((g3429) & (!g4360) & (g2170)) + ((g3429) & (g4360) & (g2170)));
	assign g2171 = (((!g893) & (!g921) & (g2088) & (g2120) & (g2089)) + ((!g893) & (g921) & (!g2088) & (g2120) & (!g2089)) + ((!g893) & (g921) & (!g2088) & (g2120) & (g2089)) + ((!g893) & (g921) & (g2088) & (!g2120) & (g2089)) + ((!g893) & (g921) & (g2088) & (g2120) & (!g2089)) + ((!g893) & (g921) & (g2088) & (g2120) & (g2089)) + ((g893) & (!g921) & (!g2088) & (g2120) & (g2089)) + ((g893) & (!g921) & (g2088) & (g2120) & (!g2089)) + ((g893) & (!g921) & (g2088) & (g2120) & (g2089)) + ((g893) & (g921) & (!g2088) & (!g2120) & (g2089)) + ((g893) & (g921) & (!g2088) & (g2120) & (!g2089)) + ((g893) & (g921) & (!g2088) & (g2120) & (g2089)) + ((g893) & (g921) & (g2088) & (!g2120) & (!g2089)) + ((g893) & (g921) & (g2088) & (!g2120) & (g2089)) + ((g893) & (g921) & (g2088) & (g2120) & (!g2089)) + ((g893) & (g921) & (g2088) & (g2120) & (g2089)));
	assign g2172 = (((!g827) & (!g960) & (g2170) & (!g2171)) + ((!g827) & (!g960) & (g2170) & (g2171)) + ((!g827) & (g960) & (g2170) & (!g2171)) + ((!g827) & (g960) & (g2170) & (g2171)) + ((g827) & (!g960) & (!g2170) & (g2171)) + ((g827) & (!g960) & (g2170) & (!g2171)) + ((g827) & (g960) & (!g2170) & (!g2171)) + ((g827) & (g960) & (g2170) & (g2171)));
	assign g7922 = (((!g2017) & (g6769) & (!g2173)) + ((!g2017) & (g6769) & (g2173)) + ((g2017) & (!g6769) & (g2173)) + ((g2017) & (g6769) & (g2173)));
	assign g2174 = (((!g895) & (!g929) & (g2091) & (g2127) & (g2092)) + ((!g895) & (g929) & (!g2091) & (g2127) & (!g2092)) + ((!g895) & (g929) & (!g2091) & (g2127) & (g2092)) + ((!g895) & (g929) & (g2091) & (!g2127) & (g2092)) + ((!g895) & (g929) & (g2091) & (g2127) & (!g2092)) + ((!g895) & (g929) & (g2091) & (g2127) & (g2092)) + ((g895) & (!g929) & (!g2091) & (g2127) & (g2092)) + ((g895) & (!g929) & (g2091) & (g2127) & (!g2092)) + ((g895) & (!g929) & (g2091) & (g2127) & (g2092)) + ((g895) & (g929) & (!g2091) & (!g2127) & (g2092)) + ((g895) & (g929) & (!g2091) & (g2127) & (!g2092)) + ((g895) & (g929) & (!g2091) & (g2127) & (g2092)) + ((g895) & (g929) & (g2091) & (!g2127) & (!g2092)) + ((g895) & (g929) & (g2091) & (!g2127) & (g2092)) + ((g895) & (g929) & (g2091) & (g2127) & (!g2092)) + ((g895) & (g929) & (g2091) & (g2127) & (g2092)));
	assign g2175 = (((!g827) & (!g962) & (g2173) & (!g2174)) + ((!g827) & (!g962) & (g2173) & (g2174)) + ((!g827) & (g962) & (g2173) & (!g2174)) + ((!g827) & (g962) & (g2173) & (g2174)) + ((g827) & (!g962) & (!g2173) & (g2174)) + ((g827) & (!g962) & (g2173) & (!g2174)) + ((g827) & (g962) & (!g2173) & (!g2174)) + ((g827) & (g962) & (g2173) & (g2174)));
	assign g2176 = (((!g2095) & (!g2096) & (!g2098) & (!g2099) & (g2129) & (g2130)) + ((!g2095) & (!g2096) & (!g2098) & (g2099) & (g2129) & (g2130)) + ((!g2095) & (!g2096) & (g2098) & (!g2099) & (g2129) & (g2130)) + ((!g2095) & (!g2096) & (g2098) & (g2099) & (!g2129) & (g2130)) + ((!g2095) & (!g2096) & (g2098) & (g2099) & (g2129) & (!g2130)) + ((!g2095) & (!g2096) & (g2098) & (g2099) & (g2129) & (g2130)) + ((!g2095) & (g2096) & (!g2098) & (!g2099) & (g2129) & (g2130)) + ((!g2095) & (g2096) & (!g2098) & (g2099) & (!g2129) & (g2130)) + ((!g2095) & (g2096) & (!g2098) & (g2099) & (g2129) & (!g2130)) + ((!g2095) & (g2096) & (!g2098) & (g2099) & (g2129) & (g2130)) + ((!g2095) & (g2096) & (g2098) & (!g2099) & (!g2129) & (g2130)) + ((!g2095) & (g2096) & (g2098) & (!g2099) & (g2129) & (!g2130)) + ((!g2095) & (g2096) & (g2098) & (!g2099) & (g2129) & (g2130)) + ((!g2095) & (g2096) & (g2098) & (g2099) & (!g2129) & (g2130)) + ((!g2095) & (g2096) & (g2098) & (g2099) & (g2129) & (!g2130)) + ((!g2095) & (g2096) & (g2098) & (g2099) & (g2129) & (g2130)) + ((g2095) & (!g2096) & (!g2098) & (!g2099) & (g2129) & (g2130)) + ((g2095) & (!g2096) & (!g2098) & (g2099) & (!g2129) & (g2130)) + ((g2095) & (!g2096) & (!g2098) & (g2099) & (g2129) & (!g2130)) + ((g2095) & (!g2096) & (!g2098) & (g2099) & (g2129) & (g2130)) + ((g2095) & (!g2096) & (g2098) & (!g2099) & (!g2129) & (g2130)) + ((g2095) & (!g2096) & (g2098) & (!g2099) & (g2129) & (!g2130)) + ((g2095) & (!g2096) & (g2098) & (!g2099) & (g2129) & (g2130)) + ((g2095) & (!g2096) & (g2098) & (g2099) & (!g2129) & (g2130)) + ((g2095) & (!g2096) & (g2098) & (g2099) & (g2129) & (!g2130)) + ((g2095) & (!g2096) & (g2098) & (g2099) & (g2129) & (g2130)) + ((g2095) & (g2096) & (!g2098) & (!g2099) & (g2129) & (g2130)) + ((g2095) & (g2096) & (!g2098) & (g2099) & (!g2129) & (g2130)) + ((g2095) & (g2096) & (!g2098) & (g2099) & (g2129) & (!g2130)) + ((g2095) & (g2096) & (!g2098) & (g2099) & (g2129) & (g2130)) + ((g2095) & (g2096) & (g2098) & (!g2099) & (!g2129) & (g2130)) + ((g2095) & (g2096) & (g2098) & (!g2099) & (g2129) & (!g2130)) + ((g2095) & (g2096) & (g2098) & (!g2099) & (g2129) & (g2130)) + ((g2095) & (g2096) & (g2098) & (g2099) & (!g2129) & (g2130)) + ((g2095) & (g2096) & (g2098) & (g2099) & (g2129) & (!g2130)) + ((g2095) & (g2096) & (g2098) & (g2099) & (g2129) & (g2130)));
	assign g7923 = (((!g3429) & (g4368) & (!g2177)) + ((!g3429) & (g4368) & (g2177)) + ((g3429) & (!g4368) & (g2177)) + ((g3429) & (g4368) & (g2177)));
	assign g7924 = (((!g3464) & (g4372) & (!g2178)) + ((!g3464) & (g4372) & (g2178)) + ((g3464) & (!g4372) & (g2178)) + ((g3464) & (g4372) & (g2178)));
	assign g2179 = (((!g2132) & (g2133) & (g2134)) + ((g2132) & (!g2133) & (g2134)) + ((g2132) & (g2133) & (!g2134)) + ((g2132) & (g2133) & (g2134)));
	assign g7925 = (((!g3429) & (g4378) & (!g2180)) + ((!g3429) & (g4378) & (g2180)) + ((g3429) & (!g4378) & (g2180)) + ((g3429) & (g4378) & (g2180)));
	assign g7926 = (((!g3499) & (g4382) & (!g2181)) + ((!g3499) & (g4382) & (g2181)) + ((g3499) & (!g4382) & (g2181)) + ((g3499) & (g4382) & (g2181)));
	assign g2182 = (((!g2179) & (!g2180) & (g2181)) + ((!g2179) & (g2180) & (!g2181)) + ((g2179) & (!g2180) & (!g2181)) + ((g2179) & (g2180) & (g2181)));
	assign g2183 = (((!g827) & (!g940) & (!g968) & (!g1946) & (g1948) & (!g2142)) + ((!g827) & (!g940) & (!g968) & (!g1946) & (g1948) & (g2142)) + ((!g827) & (!g940) & (!g968) & (g1946) & (g1948) & (!g2142)) + ((!g827) & (!g940) & (!g968) & (g1946) & (g1948) & (g2142)) + ((!g827) & (!g940) & (g968) & (!g1946) & (g1948) & (!g2142)) + ((!g827) & (!g940) & (g968) & (!g1946) & (g1948) & (g2142)) + ((!g827) & (!g940) & (g968) & (g1946) & (g1948) & (!g2142)) + ((!g827) & (!g940) & (g968) & (g1946) & (g1948) & (g2142)) + ((!g827) & (g940) & (!g968) & (!g1946) & (g1948) & (!g2142)) + ((!g827) & (g940) & (!g968) & (!g1946) & (g1948) & (g2142)) + ((!g827) & (g940) & (!g968) & (g1946) & (g1948) & (!g2142)) + ((!g827) & (g940) & (!g968) & (g1946) & (g1948) & (g2142)) + ((!g827) & (g940) & (g968) & (!g1946) & (g1948) & (!g2142)) + ((!g827) & (g940) & (g968) & (!g1946) & (g1948) & (g2142)) + ((!g827) & (g940) & (g968) & (g1946) & (g1948) & (!g2142)) + ((!g827) & (g940) & (g968) & (g1946) & (g1948) & (g2142)) + ((g827) & (!g940) & (!g968) & (!g1946) & (g1948) & (!g2142)) + ((g827) & (!g940) & (!g968) & (!g1946) & (g1948) & (g2142)) + ((g827) & (!g940) & (!g968) & (g1946) & (!g1948) & (g2142)) + ((g827) & (!g940) & (!g968) & (g1946) & (g1948) & (!g2142)) + ((g827) & (!g940) & (g968) & (!g1946) & (!g1948) & (!g2142)) + ((g827) & (!g940) & (g968) & (!g1946) & (!g1948) & (g2142)) + ((g827) & (!g940) & (g968) & (g1946) & (!g1948) & (!g2142)) + ((g827) & (!g940) & (g968) & (g1946) & (g1948) & (g2142)) + ((g827) & (g940) & (!g968) & (!g1946) & (!g1948) & (g2142)) + ((g827) & (g940) & (!g968) & (!g1946) & (g1948) & (!g2142)) + ((g827) & (g940) & (!g968) & (g1946) & (!g1948) & (!g2142)) + ((g827) & (g940) & (!g968) & (g1946) & (!g1948) & (g2142)) + ((g827) & (g940) & (g968) & (!g1946) & (!g1948) & (!g2142)) + ((g827) & (g940) & (g968) & (!g1946) & (g1948) & (g2142)) + ((g827) & (g940) & (g968) & (g1946) & (g1948) & (!g2142)) + ((g827) & (g940) & (g968) & (g1946) & (g1948) & (g2142)));
	assign g7927 = (((!g3499) & (g4385) & (!g2184)) + ((!g3499) & (g4385) & (g2184)) + ((g3499) & (!g4385) & (g2184)) + ((g3499) & (g4385) & (g2184)));
	assign g2185 = (((!g827) & (!g948) & (!g970) & (!g2153) & (g2184) & (!g2154)) + ((!g827) & (!g948) & (!g970) & (!g2153) & (g2184) & (g2154)) + ((!g827) & (!g948) & (!g970) & (g2153) & (g2184) & (!g2154)) + ((!g827) & (!g948) & (!g970) & (g2153) & (g2184) & (g2154)) + ((!g827) & (!g948) & (g970) & (!g2153) & (g2184) & (!g2154)) + ((!g827) & (!g948) & (g970) & (!g2153) & (g2184) & (g2154)) + ((!g827) & (!g948) & (g970) & (g2153) & (g2184) & (!g2154)) + ((!g827) & (!g948) & (g970) & (g2153) & (g2184) & (g2154)) + ((!g827) & (g948) & (!g970) & (!g2153) & (g2184) & (!g2154)) + ((!g827) & (g948) & (!g970) & (!g2153) & (g2184) & (g2154)) + ((!g827) & (g948) & (!g970) & (g2153) & (g2184) & (!g2154)) + ((!g827) & (g948) & (!g970) & (g2153) & (g2184) & (g2154)) + ((!g827) & (g948) & (g970) & (!g2153) & (g2184) & (!g2154)) + ((!g827) & (g948) & (g970) & (!g2153) & (g2184) & (g2154)) + ((!g827) & (g948) & (g970) & (g2153) & (g2184) & (!g2154)) + ((!g827) & (g948) & (g970) & (g2153) & (g2184) & (g2154)) + ((g827) & (!g948) & (!g970) & (!g2153) & (g2184) & (!g2154)) + ((g827) & (!g948) & (!g970) & (!g2153) & (g2184) & (g2154)) + ((g827) & (!g948) & (!g970) & (g2153) & (!g2184) & (g2154)) + ((g827) & (!g948) & (!g970) & (g2153) & (g2184) & (!g2154)) + ((g827) & (!g948) & (g970) & (!g2153) & (!g2184) & (!g2154)) + ((g827) & (!g948) & (g970) & (!g2153) & (!g2184) & (g2154)) + ((g827) & (!g948) & (g970) & (g2153) & (!g2184) & (!g2154)) + ((g827) & (!g948) & (g970) & (g2153) & (g2184) & (g2154)) + ((g827) & (g948) & (!g970) & (!g2153) & (!g2184) & (g2154)) + ((g827) & (g948) & (!g970) & (!g2153) & (g2184) & (!g2154)) + ((g827) & (g948) & (!g970) & (g2153) & (!g2184) & (!g2154)) + ((g827) & (g948) & (!g970) & (g2153) & (!g2184) & (g2154)) + ((g827) & (g948) & (g970) & (!g2153) & (!g2184) & (!g2154)) + ((g827) & (g948) & (g970) & (!g2153) & (g2184) & (g2154)) + ((g827) & (g948) & (g970) & (g2153) & (g2184) & (!g2154)) + ((g827) & (g948) & (g970) & (g2153) & (g2184) & (g2154)));
	assign g2186 = (((!g827) & (!g956) & (!g972) & (!g1947) & (g1949) & (!g2165)) + ((!g827) & (!g956) & (!g972) & (!g1947) & (g1949) & (g2165)) + ((!g827) & (!g956) & (!g972) & (g1947) & (g1949) & (!g2165)) + ((!g827) & (!g956) & (!g972) & (g1947) & (g1949) & (g2165)) + ((!g827) & (!g956) & (g972) & (!g1947) & (g1949) & (!g2165)) + ((!g827) & (!g956) & (g972) & (!g1947) & (g1949) & (g2165)) + ((!g827) & (!g956) & (g972) & (g1947) & (g1949) & (!g2165)) + ((!g827) & (!g956) & (g972) & (g1947) & (g1949) & (g2165)) + ((!g827) & (g956) & (!g972) & (!g1947) & (g1949) & (!g2165)) + ((!g827) & (g956) & (!g972) & (!g1947) & (g1949) & (g2165)) + ((!g827) & (g956) & (!g972) & (g1947) & (g1949) & (!g2165)) + ((!g827) & (g956) & (!g972) & (g1947) & (g1949) & (g2165)) + ((!g827) & (g956) & (g972) & (!g1947) & (g1949) & (!g2165)) + ((!g827) & (g956) & (g972) & (!g1947) & (g1949) & (g2165)) + ((!g827) & (g956) & (g972) & (g1947) & (g1949) & (!g2165)) + ((!g827) & (g956) & (g972) & (g1947) & (g1949) & (g2165)) + ((g827) & (!g956) & (!g972) & (!g1947) & (g1949) & (!g2165)) + ((g827) & (!g956) & (!g972) & (!g1947) & (g1949) & (g2165)) + ((g827) & (!g956) & (!g972) & (g1947) & (!g1949) & (g2165)) + ((g827) & (!g956) & (!g972) & (g1947) & (g1949) & (!g2165)) + ((g827) & (!g956) & (g972) & (!g1947) & (!g1949) & (!g2165)) + ((g827) & (!g956) & (g972) & (!g1947) & (!g1949) & (g2165)) + ((g827) & (!g956) & (g972) & (g1947) & (!g1949) & (!g2165)) + ((g827) & (!g956) & (g972) & (g1947) & (g1949) & (g2165)) + ((g827) & (g956) & (!g972) & (!g1947) & (!g1949) & (g2165)) + ((g827) & (g956) & (!g972) & (!g1947) & (g1949) & (!g2165)) + ((g827) & (g956) & (!g972) & (g1947) & (!g1949) & (!g2165)) + ((g827) & (g956) & (!g972) & (g1947) & (!g1949) & (g2165)) + ((g827) & (g956) & (g972) & (!g1947) & (!g1949) & (!g2165)) + ((g827) & (g956) & (g972) & (!g1947) & (g1949) & (g2165)) + ((g827) & (g956) & (g972) & (g1947) & (g1949) & (!g2165)) + ((g827) & (g956) & (g972) & (g1947) & (g1949) & (g2165)));
	assign g2187 = (((!g827) & (!g934) & (!g974) & (!g1984) & (g1986) & (!g2135)) + ((!g827) & (!g934) & (!g974) & (!g1984) & (g1986) & (g2135)) + ((!g827) & (!g934) & (!g974) & (g1984) & (g1986) & (!g2135)) + ((!g827) & (!g934) & (!g974) & (g1984) & (g1986) & (g2135)) + ((!g827) & (!g934) & (g974) & (!g1984) & (g1986) & (!g2135)) + ((!g827) & (!g934) & (g974) & (!g1984) & (g1986) & (g2135)) + ((!g827) & (!g934) & (g974) & (g1984) & (g1986) & (!g2135)) + ((!g827) & (!g934) & (g974) & (g1984) & (g1986) & (g2135)) + ((!g827) & (g934) & (!g974) & (!g1984) & (g1986) & (!g2135)) + ((!g827) & (g934) & (!g974) & (!g1984) & (g1986) & (g2135)) + ((!g827) & (g934) & (!g974) & (g1984) & (g1986) & (!g2135)) + ((!g827) & (g934) & (!g974) & (g1984) & (g1986) & (g2135)) + ((!g827) & (g934) & (g974) & (!g1984) & (g1986) & (!g2135)) + ((!g827) & (g934) & (g974) & (!g1984) & (g1986) & (g2135)) + ((!g827) & (g934) & (g974) & (g1984) & (g1986) & (!g2135)) + ((!g827) & (g934) & (g974) & (g1984) & (g1986) & (g2135)) + ((g827) & (!g934) & (!g974) & (!g1984) & (g1986) & (!g2135)) + ((g827) & (!g934) & (!g974) & (!g1984) & (g1986) & (g2135)) + ((g827) & (!g934) & (!g974) & (g1984) & (!g1986) & (g2135)) + ((g827) & (!g934) & (!g974) & (g1984) & (g1986) & (!g2135)) + ((g827) & (!g934) & (g974) & (!g1984) & (!g1986) & (!g2135)) + ((g827) & (!g934) & (g974) & (!g1984) & (!g1986) & (g2135)) + ((g827) & (!g934) & (g974) & (g1984) & (!g1986) & (!g2135)) + ((g827) & (!g934) & (g974) & (g1984) & (g1986) & (g2135)) + ((g827) & (g934) & (!g974) & (!g1984) & (!g1986) & (g2135)) + ((g827) & (g934) & (!g974) & (!g1984) & (g1986) & (!g2135)) + ((g827) & (g934) & (!g974) & (g1984) & (!g1986) & (!g2135)) + ((g827) & (g934) & (!g974) & (g1984) & (!g1986) & (g2135)) + ((g827) & (g934) & (g974) & (!g1984) & (!g1986) & (!g2135)) + ((g827) & (g934) & (g974) & (!g1984) & (g1986) & (g2135)) + ((g827) & (g934) & (g974) & (g1984) & (g1986) & (!g2135)) + ((g827) & (g934) & (g974) & (g1984) & (g1986) & (g2135)));
	assign g7928 = (((!g2017) & (g6762) & (!g2188)) + ((!g2017) & (g6762) & (g2188)) + ((g2017) & (!g6762) & (g2188)) + ((g2017) & (g6762) & (g2188)));
	assign g2189 = (((!g827) & (!g942) & (!g976) & (!g2144) & (g2188) & (!g2145)) + ((!g827) & (!g942) & (!g976) & (!g2144) & (g2188) & (g2145)) + ((!g827) & (!g942) & (!g976) & (g2144) & (g2188) & (!g2145)) + ((!g827) & (!g942) & (!g976) & (g2144) & (g2188) & (g2145)) + ((!g827) & (!g942) & (g976) & (!g2144) & (g2188) & (!g2145)) + ((!g827) & (!g942) & (g976) & (!g2144) & (g2188) & (g2145)) + ((!g827) & (!g942) & (g976) & (g2144) & (g2188) & (!g2145)) + ((!g827) & (!g942) & (g976) & (g2144) & (g2188) & (g2145)) + ((!g827) & (g942) & (!g976) & (!g2144) & (g2188) & (!g2145)) + ((!g827) & (g942) & (!g976) & (!g2144) & (g2188) & (g2145)) + ((!g827) & (g942) & (!g976) & (g2144) & (g2188) & (!g2145)) + ((!g827) & (g942) & (!g976) & (g2144) & (g2188) & (g2145)) + ((!g827) & (g942) & (g976) & (!g2144) & (g2188) & (!g2145)) + ((!g827) & (g942) & (g976) & (!g2144) & (g2188) & (g2145)) + ((!g827) & (g942) & (g976) & (g2144) & (g2188) & (!g2145)) + ((!g827) & (g942) & (g976) & (g2144) & (g2188) & (g2145)) + ((g827) & (!g942) & (!g976) & (!g2144) & (g2188) & (!g2145)) + ((g827) & (!g942) & (!g976) & (!g2144) & (g2188) & (g2145)) + ((g827) & (!g942) & (!g976) & (g2144) & (!g2188) & (g2145)) + ((g827) & (!g942) & (!g976) & (g2144) & (g2188) & (!g2145)) + ((g827) & (!g942) & (g976) & (!g2144) & (!g2188) & (!g2145)) + ((g827) & (!g942) & (g976) & (!g2144) & (!g2188) & (g2145)) + ((g827) & (!g942) & (g976) & (g2144) & (!g2188) & (!g2145)) + ((g827) & (!g942) & (g976) & (g2144) & (g2188) & (g2145)) + ((g827) & (g942) & (!g976) & (!g2144) & (!g2188) & (g2145)) + ((g827) & (g942) & (!g976) & (!g2144) & (g2188) & (!g2145)) + ((g827) & (g942) & (!g976) & (g2144) & (!g2188) & (!g2145)) + ((g827) & (g942) & (!g976) & (g2144) & (!g2188) & (g2145)) + ((g827) & (g942) & (g976) & (!g2144) & (!g2188) & (!g2145)) + ((g827) & (g942) & (g976) & (!g2144) & (g2188) & (g2145)) + ((g827) & (g942) & (g976) & (g2144) & (g2188) & (!g2145)) + ((g827) & (g942) & (g976) & (g2144) & (g2188) & (g2145)));
	assign g7929 = (((!g3464) & (g4391) & (!g2190)) + ((!g3464) & (g4391) & (g2190)) + ((g3464) & (!g4391) & (g2190)) + ((g3464) & (g4391) & (g2190)));
	assign g2191 = (((!g827) & (!g950) & (!g978) & (!g2156) & (g2190) & (!g2157)) + ((!g827) & (!g950) & (!g978) & (!g2156) & (g2190) & (g2157)) + ((!g827) & (!g950) & (!g978) & (g2156) & (g2190) & (!g2157)) + ((!g827) & (!g950) & (!g978) & (g2156) & (g2190) & (g2157)) + ((!g827) & (!g950) & (g978) & (!g2156) & (g2190) & (!g2157)) + ((!g827) & (!g950) & (g978) & (!g2156) & (g2190) & (g2157)) + ((!g827) & (!g950) & (g978) & (g2156) & (g2190) & (!g2157)) + ((!g827) & (!g950) & (g978) & (g2156) & (g2190) & (g2157)) + ((!g827) & (g950) & (!g978) & (!g2156) & (g2190) & (!g2157)) + ((!g827) & (g950) & (!g978) & (!g2156) & (g2190) & (g2157)) + ((!g827) & (g950) & (!g978) & (g2156) & (g2190) & (!g2157)) + ((!g827) & (g950) & (!g978) & (g2156) & (g2190) & (g2157)) + ((!g827) & (g950) & (g978) & (!g2156) & (g2190) & (!g2157)) + ((!g827) & (g950) & (g978) & (!g2156) & (g2190) & (g2157)) + ((!g827) & (g950) & (g978) & (g2156) & (g2190) & (!g2157)) + ((!g827) & (g950) & (g978) & (g2156) & (g2190) & (g2157)) + ((g827) & (!g950) & (!g978) & (!g2156) & (g2190) & (!g2157)) + ((g827) & (!g950) & (!g978) & (!g2156) & (g2190) & (g2157)) + ((g827) & (!g950) & (!g978) & (g2156) & (!g2190) & (g2157)) + ((g827) & (!g950) & (!g978) & (g2156) & (g2190) & (!g2157)) + ((g827) & (!g950) & (g978) & (!g2156) & (!g2190) & (!g2157)) + ((g827) & (!g950) & (g978) & (!g2156) & (!g2190) & (g2157)) + ((g827) & (!g950) & (g978) & (g2156) & (!g2190) & (!g2157)) + ((g827) & (!g950) & (g978) & (g2156) & (g2190) & (g2157)) + ((g827) & (g950) & (!g978) & (!g2156) & (!g2190) & (g2157)) + ((g827) & (g950) & (!g978) & (!g2156) & (g2190) & (!g2157)) + ((g827) & (g950) & (!g978) & (g2156) & (!g2190) & (!g2157)) + ((g827) & (g950) & (!g978) & (g2156) & (!g2190) & (g2157)) + ((g827) & (g950) & (g978) & (!g2156) & (!g2190) & (!g2157)) + ((g827) & (g950) & (g978) & (!g2156) & (g2190) & (g2157)) + ((g827) & (g950) & (g978) & (g2156) & (g2190) & (!g2157)) + ((g827) & (g950) & (g978) & (g2156) & (g2190) & (g2157)));
	assign g7930 = (((!g3499) & (g4394) & (!g2192)) + ((!g3499) & (g4394) & (g2192)) + ((g3499) & (!g4394) & (g2192)) + ((g3499) & (g4394) & (g2192)));
	assign g2193 = (((!g827) & (!g958) & (!g980) & (!g2167) & (g2192) & (!g2168)) + ((!g827) & (!g958) & (!g980) & (!g2167) & (g2192) & (g2168)) + ((!g827) & (!g958) & (!g980) & (g2167) & (g2192) & (!g2168)) + ((!g827) & (!g958) & (!g980) & (g2167) & (g2192) & (g2168)) + ((!g827) & (!g958) & (g980) & (!g2167) & (g2192) & (!g2168)) + ((!g827) & (!g958) & (g980) & (!g2167) & (g2192) & (g2168)) + ((!g827) & (!g958) & (g980) & (g2167) & (g2192) & (!g2168)) + ((!g827) & (!g958) & (g980) & (g2167) & (g2192) & (g2168)) + ((!g827) & (g958) & (!g980) & (!g2167) & (g2192) & (!g2168)) + ((!g827) & (g958) & (!g980) & (!g2167) & (g2192) & (g2168)) + ((!g827) & (g958) & (!g980) & (g2167) & (g2192) & (!g2168)) + ((!g827) & (g958) & (!g980) & (g2167) & (g2192) & (g2168)) + ((!g827) & (g958) & (g980) & (!g2167) & (g2192) & (!g2168)) + ((!g827) & (g958) & (g980) & (!g2167) & (g2192) & (g2168)) + ((!g827) & (g958) & (g980) & (g2167) & (g2192) & (!g2168)) + ((!g827) & (g958) & (g980) & (g2167) & (g2192) & (g2168)) + ((g827) & (!g958) & (!g980) & (!g2167) & (g2192) & (!g2168)) + ((g827) & (!g958) & (!g980) & (!g2167) & (g2192) & (g2168)) + ((g827) & (!g958) & (!g980) & (g2167) & (!g2192) & (g2168)) + ((g827) & (!g958) & (!g980) & (g2167) & (g2192) & (!g2168)) + ((g827) & (!g958) & (g980) & (!g2167) & (!g2192) & (!g2168)) + ((g827) & (!g958) & (g980) & (!g2167) & (!g2192) & (g2168)) + ((g827) & (!g958) & (g980) & (g2167) & (!g2192) & (!g2168)) + ((g827) & (!g958) & (g980) & (g2167) & (g2192) & (g2168)) + ((g827) & (g958) & (!g980) & (!g2167) & (!g2192) & (g2168)) + ((g827) & (g958) & (!g980) & (!g2167) & (g2192) & (!g2168)) + ((g827) & (g958) & (!g980) & (g2167) & (!g2192) & (!g2168)) + ((g827) & (g958) & (!g980) & (g2167) & (!g2192) & (g2168)) + ((g827) & (g958) & (g980) & (!g2167) & (!g2192) & (!g2168)) + ((g827) & (g958) & (g980) & (!g2167) & (g2192) & (g2168)) + ((g827) & (g958) & (g980) & (g2167) & (g2192) & (!g2168)) + ((g827) & (g958) & (g980) & (g2167) & (g2192) & (g2168)));
	assign g7931 = (((!g3464) & (g4397) & (!g2194)) + ((!g3464) & (g4397) & (g2194)) + ((g3464) & (!g4397) & (g2194)) + ((g3464) & (g4397) & (g2194)));
	assign g2195 = (((!g827) & (!g936) & (!g982) & (!g2137) & (g2194) & (!g2138)) + ((!g827) & (!g936) & (!g982) & (!g2137) & (g2194) & (g2138)) + ((!g827) & (!g936) & (!g982) & (g2137) & (g2194) & (!g2138)) + ((!g827) & (!g936) & (!g982) & (g2137) & (g2194) & (g2138)) + ((!g827) & (!g936) & (g982) & (!g2137) & (g2194) & (!g2138)) + ((!g827) & (!g936) & (g982) & (!g2137) & (g2194) & (g2138)) + ((!g827) & (!g936) & (g982) & (g2137) & (g2194) & (!g2138)) + ((!g827) & (!g936) & (g982) & (g2137) & (g2194) & (g2138)) + ((!g827) & (g936) & (!g982) & (!g2137) & (g2194) & (!g2138)) + ((!g827) & (g936) & (!g982) & (!g2137) & (g2194) & (g2138)) + ((!g827) & (g936) & (!g982) & (g2137) & (g2194) & (!g2138)) + ((!g827) & (g936) & (!g982) & (g2137) & (g2194) & (g2138)) + ((!g827) & (g936) & (g982) & (!g2137) & (g2194) & (!g2138)) + ((!g827) & (g936) & (g982) & (!g2137) & (g2194) & (g2138)) + ((!g827) & (g936) & (g982) & (g2137) & (g2194) & (!g2138)) + ((!g827) & (g936) & (g982) & (g2137) & (g2194) & (g2138)) + ((g827) & (!g936) & (!g982) & (!g2137) & (g2194) & (!g2138)) + ((g827) & (!g936) & (!g982) & (!g2137) & (g2194) & (g2138)) + ((g827) & (!g936) & (!g982) & (g2137) & (!g2194) & (g2138)) + ((g827) & (!g936) & (!g982) & (g2137) & (g2194) & (!g2138)) + ((g827) & (!g936) & (g982) & (!g2137) & (!g2194) & (!g2138)) + ((g827) & (!g936) & (g982) & (!g2137) & (!g2194) & (g2138)) + ((g827) & (!g936) & (g982) & (g2137) & (!g2194) & (!g2138)) + ((g827) & (!g936) & (g982) & (g2137) & (g2194) & (g2138)) + ((g827) & (g936) & (!g982) & (!g2137) & (!g2194) & (g2138)) + ((g827) & (g936) & (!g982) & (!g2137) & (g2194) & (!g2138)) + ((g827) & (g936) & (!g982) & (g2137) & (!g2194) & (!g2138)) + ((g827) & (g936) & (!g982) & (g2137) & (!g2194) & (g2138)) + ((g827) & (g936) & (g982) & (!g2137) & (!g2194) & (!g2138)) + ((g827) & (g936) & (g982) & (!g2137) & (g2194) & (g2138)) + ((g827) & (g936) & (g982) & (g2137) & (g2194) & (!g2138)) + ((g827) & (g936) & (g982) & (g2137) & (g2194) & (g2138)));
	assign g7932 = (((!g3499) & (g4400) & (!g2196)) + ((!g3499) & (g4400) & (g2196)) + ((g3499) & (!g4400) & (g2196)) + ((g3499) & (g4400) & (g2196)));
	assign g2197 = (((!g827) & (!g944) & (!g984) & (!g2147) & (g2196) & (!g2148)) + ((!g827) & (!g944) & (!g984) & (!g2147) & (g2196) & (g2148)) + ((!g827) & (!g944) & (!g984) & (g2147) & (g2196) & (!g2148)) + ((!g827) & (!g944) & (!g984) & (g2147) & (g2196) & (g2148)) + ((!g827) & (!g944) & (g984) & (!g2147) & (g2196) & (!g2148)) + ((!g827) & (!g944) & (g984) & (!g2147) & (g2196) & (g2148)) + ((!g827) & (!g944) & (g984) & (g2147) & (g2196) & (!g2148)) + ((!g827) & (!g944) & (g984) & (g2147) & (g2196) & (g2148)) + ((!g827) & (g944) & (!g984) & (!g2147) & (g2196) & (!g2148)) + ((!g827) & (g944) & (!g984) & (!g2147) & (g2196) & (g2148)) + ((!g827) & (g944) & (!g984) & (g2147) & (g2196) & (!g2148)) + ((!g827) & (g944) & (!g984) & (g2147) & (g2196) & (g2148)) + ((!g827) & (g944) & (g984) & (!g2147) & (g2196) & (!g2148)) + ((!g827) & (g944) & (g984) & (!g2147) & (g2196) & (g2148)) + ((!g827) & (g944) & (g984) & (g2147) & (g2196) & (!g2148)) + ((!g827) & (g944) & (g984) & (g2147) & (g2196) & (g2148)) + ((g827) & (!g944) & (!g984) & (!g2147) & (g2196) & (!g2148)) + ((g827) & (!g944) & (!g984) & (!g2147) & (g2196) & (g2148)) + ((g827) & (!g944) & (!g984) & (g2147) & (!g2196) & (g2148)) + ((g827) & (!g944) & (!g984) & (g2147) & (g2196) & (!g2148)) + ((g827) & (!g944) & (g984) & (!g2147) & (!g2196) & (!g2148)) + ((g827) & (!g944) & (g984) & (!g2147) & (!g2196) & (g2148)) + ((g827) & (!g944) & (g984) & (g2147) & (!g2196) & (!g2148)) + ((g827) & (!g944) & (g984) & (g2147) & (g2196) & (g2148)) + ((g827) & (g944) & (!g984) & (!g2147) & (!g2196) & (g2148)) + ((g827) & (g944) & (!g984) & (!g2147) & (g2196) & (!g2148)) + ((g827) & (g944) & (!g984) & (g2147) & (!g2196) & (!g2148)) + ((g827) & (g944) & (!g984) & (g2147) & (!g2196) & (g2148)) + ((g827) & (g944) & (g984) & (!g2147) & (!g2196) & (!g2148)) + ((g827) & (g944) & (g984) & (!g2147) & (g2196) & (g2148)) + ((g827) & (g944) & (g984) & (g2147) & (g2196) & (!g2148)) + ((g827) & (g944) & (g984) & (g2147) & (g2196) & (g2148)));
	assign g7933 = (((!g2017) & (g6755) & (!g2198)) + ((!g2017) & (g6755) & (g2198)) + ((g2017) & (!g6755) & (g2198)) + ((g2017) & (g6755) & (g2198)));
	assign g2199 = (((!g827) & (!g952) & (!g986) & (!g2159) & (g2198) & (!g2160)) + ((!g827) & (!g952) & (!g986) & (!g2159) & (g2198) & (g2160)) + ((!g827) & (!g952) & (!g986) & (g2159) & (g2198) & (!g2160)) + ((!g827) & (!g952) & (!g986) & (g2159) & (g2198) & (g2160)) + ((!g827) & (!g952) & (g986) & (!g2159) & (g2198) & (!g2160)) + ((!g827) & (!g952) & (g986) & (!g2159) & (g2198) & (g2160)) + ((!g827) & (!g952) & (g986) & (g2159) & (g2198) & (!g2160)) + ((!g827) & (!g952) & (g986) & (g2159) & (g2198) & (g2160)) + ((!g827) & (g952) & (!g986) & (!g2159) & (g2198) & (!g2160)) + ((!g827) & (g952) & (!g986) & (!g2159) & (g2198) & (g2160)) + ((!g827) & (g952) & (!g986) & (g2159) & (g2198) & (!g2160)) + ((!g827) & (g952) & (!g986) & (g2159) & (g2198) & (g2160)) + ((!g827) & (g952) & (g986) & (!g2159) & (g2198) & (!g2160)) + ((!g827) & (g952) & (g986) & (!g2159) & (g2198) & (g2160)) + ((!g827) & (g952) & (g986) & (g2159) & (g2198) & (!g2160)) + ((!g827) & (g952) & (g986) & (g2159) & (g2198) & (g2160)) + ((g827) & (!g952) & (!g986) & (!g2159) & (g2198) & (!g2160)) + ((g827) & (!g952) & (!g986) & (!g2159) & (g2198) & (g2160)) + ((g827) & (!g952) & (!g986) & (g2159) & (!g2198) & (g2160)) + ((g827) & (!g952) & (!g986) & (g2159) & (g2198) & (!g2160)) + ((g827) & (!g952) & (g986) & (!g2159) & (!g2198) & (!g2160)) + ((g827) & (!g952) & (g986) & (!g2159) & (!g2198) & (g2160)) + ((g827) & (!g952) & (g986) & (g2159) & (!g2198) & (!g2160)) + ((g827) & (!g952) & (g986) & (g2159) & (g2198) & (g2160)) + ((g827) & (g952) & (!g986) & (!g2159) & (!g2198) & (g2160)) + ((g827) & (g952) & (!g986) & (!g2159) & (g2198) & (!g2160)) + ((g827) & (g952) & (!g986) & (g2159) & (!g2198) & (!g2160)) + ((g827) & (g952) & (!g986) & (g2159) & (!g2198) & (g2160)) + ((g827) & (g952) & (g986) & (!g2159) & (!g2198) & (!g2160)) + ((g827) & (g952) & (g986) & (!g2159) & (g2198) & (g2160)) + ((g827) & (g952) & (g986) & (g2159) & (g2198) & (!g2160)) + ((g827) & (g952) & (g986) & (g2159) & (g2198) & (g2160)));
	assign g7934 = (((!g3429) & (g4407) & (!g2200)) + ((!g3429) & (g4407) & (g2200)) + ((g3429) & (!g4407) & (g2200)) + ((g3429) & (g4407) & (g2200)));
	assign g2201 = (((!g827) & (!g960) & (!g988) & (!g2170) & (g2200) & (!g2171)) + ((!g827) & (!g960) & (!g988) & (!g2170) & (g2200) & (g2171)) + ((!g827) & (!g960) & (!g988) & (g2170) & (g2200) & (!g2171)) + ((!g827) & (!g960) & (!g988) & (g2170) & (g2200) & (g2171)) + ((!g827) & (!g960) & (g988) & (!g2170) & (g2200) & (!g2171)) + ((!g827) & (!g960) & (g988) & (!g2170) & (g2200) & (g2171)) + ((!g827) & (!g960) & (g988) & (g2170) & (g2200) & (!g2171)) + ((!g827) & (!g960) & (g988) & (g2170) & (g2200) & (g2171)) + ((!g827) & (g960) & (!g988) & (!g2170) & (g2200) & (!g2171)) + ((!g827) & (g960) & (!g988) & (!g2170) & (g2200) & (g2171)) + ((!g827) & (g960) & (!g988) & (g2170) & (g2200) & (!g2171)) + ((!g827) & (g960) & (!g988) & (g2170) & (g2200) & (g2171)) + ((!g827) & (g960) & (g988) & (!g2170) & (g2200) & (!g2171)) + ((!g827) & (g960) & (g988) & (!g2170) & (g2200) & (g2171)) + ((!g827) & (g960) & (g988) & (g2170) & (g2200) & (!g2171)) + ((!g827) & (g960) & (g988) & (g2170) & (g2200) & (g2171)) + ((g827) & (!g960) & (!g988) & (!g2170) & (g2200) & (!g2171)) + ((g827) & (!g960) & (!g988) & (!g2170) & (g2200) & (g2171)) + ((g827) & (!g960) & (!g988) & (g2170) & (!g2200) & (g2171)) + ((g827) & (!g960) & (!g988) & (g2170) & (g2200) & (!g2171)) + ((g827) & (!g960) & (g988) & (!g2170) & (!g2200) & (!g2171)) + ((g827) & (!g960) & (g988) & (!g2170) & (!g2200) & (g2171)) + ((g827) & (!g960) & (g988) & (g2170) & (!g2200) & (!g2171)) + ((g827) & (!g960) & (g988) & (g2170) & (g2200) & (g2171)) + ((g827) & (g960) & (!g988) & (!g2170) & (!g2200) & (g2171)) + ((g827) & (g960) & (!g988) & (!g2170) & (g2200) & (!g2171)) + ((g827) & (g960) & (!g988) & (g2170) & (!g2200) & (!g2171)) + ((g827) & (g960) & (!g988) & (g2170) & (!g2200) & (g2171)) + ((g827) & (g960) & (g988) & (!g2170) & (!g2200) & (!g2171)) + ((g827) & (g960) & (g988) & (!g2170) & (g2200) & (g2171)) + ((g827) & (g960) & (g988) & (g2170) & (g2200) & (!g2171)) + ((g827) & (g960) & (g988) & (g2170) & (g2200) & (g2171)));
	assign g2202 = (((!g827) & (!g938) & (!g990) & (!g1985) & (g1987) & (!g2140)) + ((!g827) & (!g938) & (!g990) & (!g1985) & (g1987) & (g2140)) + ((!g827) & (!g938) & (!g990) & (g1985) & (g1987) & (!g2140)) + ((!g827) & (!g938) & (!g990) & (g1985) & (g1987) & (g2140)) + ((!g827) & (!g938) & (g990) & (!g1985) & (g1987) & (!g2140)) + ((!g827) & (!g938) & (g990) & (!g1985) & (g1987) & (g2140)) + ((!g827) & (!g938) & (g990) & (g1985) & (g1987) & (!g2140)) + ((!g827) & (!g938) & (g990) & (g1985) & (g1987) & (g2140)) + ((!g827) & (g938) & (!g990) & (!g1985) & (g1987) & (!g2140)) + ((!g827) & (g938) & (!g990) & (!g1985) & (g1987) & (g2140)) + ((!g827) & (g938) & (!g990) & (g1985) & (g1987) & (!g2140)) + ((!g827) & (g938) & (!g990) & (g1985) & (g1987) & (g2140)) + ((!g827) & (g938) & (g990) & (!g1985) & (g1987) & (!g2140)) + ((!g827) & (g938) & (g990) & (!g1985) & (g1987) & (g2140)) + ((!g827) & (g938) & (g990) & (g1985) & (g1987) & (!g2140)) + ((!g827) & (g938) & (g990) & (g1985) & (g1987) & (g2140)) + ((g827) & (!g938) & (!g990) & (!g1985) & (g1987) & (!g2140)) + ((g827) & (!g938) & (!g990) & (!g1985) & (g1987) & (g2140)) + ((g827) & (!g938) & (!g990) & (g1985) & (!g1987) & (g2140)) + ((g827) & (!g938) & (!g990) & (g1985) & (g1987) & (!g2140)) + ((g827) & (!g938) & (g990) & (!g1985) & (!g1987) & (!g2140)) + ((g827) & (!g938) & (g990) & (!g1985) & (!g1987) & (g2140)) + ((g827) & (!g938) & (g990) & (g1985) & (!g1987) & (!g2140)) + ((g827) & (!g938) & (g990) & (g1985) & (g1987) & (g2140)) + ((g827) & (g938) & (!g990) & (!g1985) & (!g1987) & (g2140)) + ((g827) & (g938) & (!g990) & (!g1985) & (g1987) & (!g2140)) + ((g827) & (g938) & (!g990) & (g1985) & (!g1987) & (!g2140)) + ((g827) & (g938) & (!g990) & (g1985) & (!g1987) & (g2140)) + ((g827) & (g938) & (g990) & (!g1985) & (!g1987) & (!g2140)) + ((g827) & (g938) & (g990) & (!g1985) & (g1987) & (g2140)) + ((g827) & (g938) & (g990) & (g1985) & (g1987) & (!g2140)) + ((g827) & (g938) & (g990) & (g1985) & (g1987) & (g2140)));
	assign g7935 = (((!g3464) & (g4410) & (!g2203)) + ((!g3464) & (g4410) & (g2203)) + ((g3464) & (!g4410) & (g2203)) + ((g3464) & (g4410) & (g2203)));
	assign g2204 = (((!g827) & (!g946) & (!g992) & (!g2150) & (g2203) & (!g2151)) + ((!g827) & (!g946) & (!g992) & (!g2150) & (g2203) & (g2151)) + ((!g827) & (!g946) & (!g992) & (g2150) & (g2203) & (!g2151)) + ((!g827) & (!g946) & (!g992) & (g2150) & (g2203) & (g2151)) + ((!g827) & (!g946) & (g992) & (!g2150) & (g2203) & (!g2151)) + ((!g827) & (!g946) & (g992) & (!g2150) & (g2203) & (g2151)) + ((!g827) & (!g946) & (g992) & (g2150) & (g2203) & (!g2151)) + ((!g827) & (!g946) & (g992) & (g2150) & (g2203) & (g2151)) + ((!g827) & (g946) & (!g992) & (!g2150) & (g2203) & (!g2151)) + ((!g827) & (g946) & (!g992) & (!g2150) & (g2203) & (g2151)) + ((!g827) & (g946) & (!g992) & (g2150) & (g2203) & (!g2151)) + ((!g827) & (g946) & (!g992) & (g2150) & (g2203) & (g2151)) + ((!g827) & (g946) & (g992) & (!g2150) & (g2203) & (!g2151)) + ((!g827) & (g946) & (g992) & (!g2150) & (g2203) & (g2151)) + ((!g827) & (g946) & (g992) & (g2150) & (g2203) & (!g2151)) + ((!g827) & (g946) & (g992) & (g2150) & (g2203) & (g2151)) + ((g827) & (!g946) & (!g992) & (!g2150) & (g2203) & (!g2151)) + ((g827) & (!g946) & (!g992) & (!g2150) & (g2203) & (g2151)) + ((g827) & (!g946) & (!g992) & (g2150) & (!g2203) & (g2151)) + ((g827) & (!g946) & (!g992) & (g2150) & (g2203) & (!g2151)) + ((g827) & (!g946) & (g992) & (!g2150) & (!g2203) & (!g2151)) + ((g827) & (!g946) & (g992) & (!g2150) & (!g2203) & (g2151)) + ((g827) & (!g946) & (g992) & (g2150) & (!g2203) & (!g2151)) + ((g827) & (!g946) & (g992) & (g2150) & (g2203) & (g2151)) + ((g827) & (g946) & (!g992) & (!g2150) & (!g2203) & (g2151)) + ((g827) & (g946) & (!g992) & (!g2150) & (g2203) & (!g2151)) + ((g827) & (g946) & (!g992) & (g2150) & (!g2203) & (!g2151)) + ((g827) & (g946) & (!g992) & (g2150) & (!g2203) & (g2151)) + ((g827) & (g946) & (g992) & (!g2150) & (!g2203) & (!g2151)) + ((g827) & (g946) & (g992) & (!g2150) & (g2203) & (g2151)) + ((g827) & (g946) & (g992) & (g2150) & (g2203) & (!g2151)) + ((g827) & (g946) & (g992) & (g2150) & (g2203) & (g2151)));
	assign g7936 = (((!g3429) & (g4415) & (!g2205)) + ((!g3429) & (g4415) & (g2205)) + ((g3429) & (!g4415) & (g2205)) + ((g3429) & (g4415) & (g2205)));
	assign g2206 = (((!g827) & (!g954) & (!g994) & (!g2162) & (g2205) & (!g2163)) + ((!g827) & (!g954) & (!g994) & (!g2162) & (g2205) & (g2163)) + ((!g827) & (!g954) & (!g994) & (g2162) & (g2205) & (!g2163)) + ((!g827) & (!g954) & (!g994) & (g2162) & (g2205) & (g2163)) + ((!g827) & (!g954) & (g994) & (!g2162) & (g2205) & (!g2163)) + ((!g827) & (!g954) & (g994) & (!g2162) & (g2205) & (g2163)) + ((!g827) & (!g954) & (g994) & (g2162) & (g2205) & (!g2163)) + ((!g827) & (!g954) & (g994) & (g2162) & (g2205) & (g2163)) + ((!g827) & (g954) & (!g994) & (!g2162) & (g2205) & (!g2163)) + ((!g827) & (g954) & (!g994) & (!g2162) & (g2205) & (g2163)) + ((!g827) & (g954) & (!g994) & (g2162) & (g2205) & (!g2163)) + ((!g827) & (g954) & (!g994) & (g2162) & (g2205) & (g2163)) + ((!g827) & (g954) & (g994) & (!g2162) & (g2205) & (!g2163)) + ((!g827) & (g954) & (g994) & (!g2162) & (g2205) & (g2163)) + ((!g827) & (g954) & (g994) & (g2162) & (g2205) & (!g2163)) + ((!g827) & (g954) & (g994) & (g2162) & (g2205) & (g2163)) + ((g827) & (!g954) & (!g994) & (!g2162) & (g2205) & (!g2163)) + ((g827) & (!g954) & (!g994) & (!g2162) & (g2205) & (g2163)) + ((g827) & (!g954) & (!g994) & (g2162) & (!g2205) & (g2163)) + ((g827) & (!g954) & (!g994) & (g2162) & (g2205) & (!g2163)) + ((g827) & (!g954) & (g994) & (!g2162) & (!g2205) & (!g2163)) + ((g827) & (!g954) & (g994) & (!g2162) & (!g2205) & (g2163)) + ((g827) & (!g954) & (g994) & (g2162) & (!g2205) & (!g2163)) + ((g827) & (!g954) & (g994) & (g2162) & (g2205) & (g2163)) + ((g827) & (g954) & (!g994) & (!g2162) & (!g2205) & (g2163)) + ((g827) & (g954) & (!g994) & (!g2162) & (g2205) & (!g2163)) + ((g827) & (g954) & (!g994) & (g2162) & (!g2205) & (!g2163)) + ((g827) & (g954) & (!g994) & (g2162) & (!g2205) & (g2163)) + ((g827) & (g954) & (g994) & (!g2162) & (!g2205) & (!g2163)) + ((g827) & (g954) & (g994) & (!g2162) & (g2205) & (g2163)) + ((g827) & (g954) & (g994) & (g2162) & (g2205) & (!g2163)) + ((g827) & (g954) & (g994) & (g2162) & (g2205) & (g2163)));
	assign g7937 = (((!g2017) & (g6748) & (!g2207)) + ((!g2017) & (g6748) & (g2207)) + ((g2017) & (!g6748) & (g2207)) + ((g2017) & (g6748) & (g2207)));
	assign g2208 = (((!g827) & (!g962) & (!g996) & (!g2173) & (g2207) & (!g2174)) + ((!g827) & (!g962) & (!g996) & (!g2173) & (g2207) & (g2174)) + ((!g827) & (!g962) & (!g996) & (g2173) & (g2207) & (!g2174)) + ((!g827) & (!g962) & (!g996) & (g2173) & (g2207) & (g2174)) + ((!g827) & (!g962) & (g996) & (!g2173) & (g2207) & (!g2174)) + ((!g827) & (!g962) & (g996) & (!g2173) & (g2207) & (g2174)) + ((!g827) & (!g962) & (g996) & (g2173) & (g2207) & (!g2174)) + ((!g827) & (!g962) & (g996) & (g2173) & (g2207) & (g2174)) + ((!g827) & (g962) & (!g996) & (!g2173) & (g2207) & (!g2174)) + ((!g827) & (g962) & (!g996) & (!g2173) & (g2207) & (g2174)) + ((!g827) & (g962) & (!g996) & (g2173) & (g2207) & (!g2174)) + ((!g827) & (g962) & (!g996) & (g2173) & (g2207) & (g2174)) + ((!g827) & (g962) & (g996) & (!g2173) & (g2207) & (!g2174)) + ((!g827) & (g962) & (g996) & (!g2173) & (g2207) & (g2174)) + ((!g827) & (g962) & (g996) & (g2173) & (g2207) & (!g2174)) + ((!g827) & (g962) & (g996) & (g2173) & (g2207) & (g2174)) + ((g827) & (!g962) & (!g996) & (!g2173) & (g2207) & (!g2174)) + ((g827) & (!g962) & (!g996) & (!g2173) & (g2207) & (g2174)) + ((g827) & (!g962) & (!g996) & (g2173) & (!g2207) & (g2174)) + ((g827) & (!g962) & (!g996) & (g2173) & (g2207) & (!g2174)) + ((g827) & (!g962) & (g996) & (!g2173) & (!g2207) & (!g2174)) + ((g827) & (!g962) & (g996) & (!g2173) & (!g2207) & (g2174)) + ((g827) & (!g962) & (g996) & (g2173) & (!g2207) & (!g2174)) + ((g827) & (!g962) & (g996) & (g2173) & (g2207) & (g2174)) + ((g827) & (g962) & (!g996) & (!g2173) & (!g2207) & (g2174)) + ((g827) & (g962) & (!g996) & (!g2173) & (g2207) & (!g2174)) + ((g827) & (g962) & (!g996) & (g2173) & (!g2207) & (!g2174)) + ((g827) & (g962) & (!g996) & (g2173) & (!g2207) & (g2174)) + ((g827) & (g962) & (g996) & (!g2173) & (!g2207) & (!g2174)) + ((g827) & (g962) & (g996) & (!g2173) & (g2207) & (g2174)) + ((g827) & (g962) & (g996) & (g2173) & (g2207) & (!g2174)) + ((g827) & (g962) & (g996) & (g2173) & (g2207) & (g2174)));
	assign g2209 = (((!g2176) & (g2177) & (g2178)) + ((g2176) & (!g2177) & (g2178)) + ((g2176) & (g2177) & (!g2178)) + ((g2176) & (g2177) & (g2178)));
	assign g7938 = (((!g3429) & (g4420) & (!g2210)) + ((!g3429) & (g4420) & (g2210)) + ((g3429) & (!g4420) & (g2210)) + ((g3429) & (g4420) & (g2210)));
	assign g7939 = (((!g3464) & (g4424) & (!g2211)) + ((!g3464) & (g4424) & (g2211)) + ((g3464) & (!g4424) & (g2211)) + ((g3464) & (g4424) & (g2211)));
	assign g7940 = (((!g3429) & (g4427) & (!g2212)) + ((!g3429) & (g4427) & (g2212)) + ((g3429) & (!g4427) & (g2212)) + ((g3429) & (g4427) & (g2212)));
	assign g7941 = (((!g3499) & (g4431) & (!g2213)) + ((!g3499) & (g4431) & (g2213)) + ((g3499) & (!g4431) & (g2213)) + ((g3499) & (g4431) & (g2213)));
	assign g2214 = (((!g2179) & (!g2180) & (!g2181) & (!g2212) & (g2213)) + ((!g2179) & (!g2180) & (!g2181) & (g2212) & (!g2213)) + ((!g2179) & (!g2180) & (g2181) & (!g2212) & (g2213)) + ((!g2179) & (!g2180) & (g2181) & (g2212) & (!g2213)) + ((!g2179) & (g2180) & (!g2181) & (!g2212) & (g2213)) + ((!g2179) & (g2180) & (!g2181) & (g2212) & (!g2213)) + ((!g2179) & (g2180) & (g2181) & (!g2212) & (!g2213)) + ((!g2179) & (g2180) & (g2181) & (g2212) & (g2213)) + ((g2179) & (!g2180) & (!g2181) & (!g2212) & (g2213)) + ((g2179) & (!g2180) & (!g2181) & (g2212) & (!g2213)) + ((g2179) & (!g2180) & (g2181) & (!g2212) & (!g2213)) + ((g2179) & (!g2180) & (g2181) & (g2212) & (g2213)) + ((g2179) & (g2180) & (!g2181) & (!g2212) & (!g2213)) + ((g2179) & (g2180) & (!g2181) & (g2212) & (g2213)) + ((g2179) & (g2180) & (g2181) & (!g2212) & (!g2213)) + ((g2179) & (g2180) & (g2181) & (g2212) & (g2213)));
	assign g2215 = (((!g934) & (!g974) & (g1984) & (g1986) & (g2135)) + ((!g934) & (g974) & (!g1984) & (g1986) & (!g2135)) + ((!g934) & (g974) & (!g1984) & (g1986) & (g2135)) + ((!g934) & (g974) & (g1984) & (!g1986) & (g2135)) + ((!g934) & (g974) & (g1984) & (g1986) & (!g2135)) + ((!g934) & (g974) & (g1984) & (g1986) & (g2135)) + ((g934) & (!g974) & (!g1984) & (g1986) & (g2135)) + ((g934) & (!g974) & (g1984) & (g1986) & (!g2135)) + ((g934) & (!g974) & (g1984) & (g1986) & (g2135)) + ((g934) & (g974) & (!g1984) & (!g1986) & (g2135)) + ((g934) & (g974) & (!g1984) & (g1986) & (!g2135)) + ((g934) & (g974) & (!g1984) & (g1986) & (g2135)) + ((g934) & (g974) & (g1984) & (!g1986) & (!g2135)) + ((g934) & (g974) & (g1984) & (!g1986) & (g2135)) + ((g934) & (g974) & (g1984) & (g1986) & (!g2135)) + ((g934) & (g974) & (g1984) & (g1986) & (g2135)));
	assign g2216 = (((!g827) & (!g1001) & (g1991) & (!g2215)) + ((!g827) & (!g1001) & (g1991) & (g2215)) + ((!g827) & (g1001) & (g1991) & (!g2215)) + ((!g827) & (g1001) & (g1991) & (g2215)) + ((g827) & (!g1001) & (!g1991) & (g2215)) + ((g827) & (!g1001) & (g1991) & (!g2215)) + ((g827) & (g1001) & (!g1991) & (!g2215)) + ((g827) & (g1001) & (g1991) & (g2215)));
	assign g7942 = (((!g3464) & (g4434) & (!g2217)) + ((!g3464) & (g4434) & (g2217)) + ((g3464) & (!g4434) & (g2217)) + ((g3464) & (g4434) & (g2217)));
	assign g2218 = (((!g936) & (!g982) & (g2137) & (g2194) & (g2138)) + ((!g936) & (g982) & (!g2137) & (g2194) & (!g2138)) + ((!g936) & (g982) & (!g2137) & (g2194) & (g2138)) + ((!g936) & (g982) & (g2137) & (!g2194) & (g2138)) + ((!g936) & (g982) & (g2137) & (g2194) & (!g2138)) + ((!g936) & (g982) & (g2137) & (g2194) & (g2138)) + ((g936) & (!g982) & (!g2137) & (g2194) & (g2138)) + ((g936) & (!g982) & (g2137) & (g2194) & (!g2138)) + ((g936) & (!g982) & (g2137) & (g2194) & (g2138)) + ((g936) & (g982) & (!g2137) & (!g2194) & (g2138)) + ((g936) & (g982) & (!g2137) & (g2194) & (!g2138)) + ((g936) & (g982) & (!g2137) & (g2194) & (g2138)) + ((g936) & (g982) & (g2137) & (!g2194) & (!g2138)) + ((g936) & (g982) & (g2137) & (!g2194) & (g2138)) + ((g936) & (g982) & (g2137) & (g2194) & (!g2138)) + ((g936) & (g982) & (g2137) & (g2194) & (g2138)));
	assign g2219 = (((!g827) & (!g1003) & (g2217) & (!g2218)) + ((!g827) & (!g1003) & (g2217) & (g2218)) + ((!g827) & (g1003) & (g2217) & (!g2218)) + ((!g827) & (g1003) & (g2217) & (g2218)) + ((g827) & (!g1003) & (!g2217) & (g2218)) + ((g827) & (!g1003) & (g2217) & (!g2218)) + ((g827) & (g1003) & (!g2217) & (!g2218)) + ((g827) & (g1003) & (g2217) & (g2218)));
	assign g2220 = (((!g938) & (!g990) & (g1985) & (g1987) & (g2140)) + ((!g938) & (g990) & (!g1985) & (g1987) & (!g2140)) + ((!g938) & (g990) & (!g1985) & (g1987) & (g2140)) + ((!g938) & (g990) & (g1985) & (!g1987) & (g2140)) + ((!g938) & (g990) & (g1985) & (g1987) & (!g2140)) + ((!g938) & (g990) & (g1985) & (g1987) & (g2140)) + ((g938) & (!g990) & (!g1985) & (g1987) & (g2140)) + ((g938) & (!g990) & (g1985) & (g1987) & (!g2140)) + ((g938) & (!g990) & (g1985) & (g1987) & (g2140)) + ((g938) & (g990) & (!g1985) & (!g1987) & (g2140)) + ((g938) & (g990) & (!g1985) & (g1987) & (!g2140)) + ((g938) & (g990) & (!g1985) & (g1987) & (g2140)) + ((g938) & (g990) & (g1985) & (!g1987) & (!g2140)) + ((g938) & (g990) & (g1985) & (!g1987) & (g2140)) + ((g938) & (g990) & (g1985) & (g1987) & (!g2140)) + ((g938) & (g990) & (g1985) & (g1987) & (g2140)));
	assign g2221 = (((!g827) & (!g1005) & (g1992) & (!g2220)) + ((!g827) & (!g1005) & (g1992) & (g2220)) + ((!g827) & (g1005) & (g1992) & (!g2220)) + ((!g827) & (g1005) & (g1992) & (g2220)) + ((g827) & (!g1005) & (!g1992) & (g2220)) + ((g827) & (!g1005) & (g1992) & (!g2220)) + ((g827) & (g1005) & (!g1992) & (!g2220)) + ((g827) & (g1005) & (g1992) & (g2220)));
	assign g2222 = (((!g940) & (!g968) & (g1946) & (g1948) & (g2142)) + ((!g940) & (g968) & (!g1946) & (g1948) & (!g2142)) + ((!g940) & (g968) & (!g1946) & (g1948) & (g2142)) + ((!g940) & (g968) & (g1946) & (!g1948) & (g2142)) + ((!g940) & (g968) & (g1946) & (g1948) & (!g2142)) + ((!g940) & (g968) & (g1946) & (g1948) & (g2142)) + ((g940) & (!g968) & (!g1946) & (g1948) & (g2142)) + ((g940) & (!g968) & (g1946) & (g1948) & (!g2142)) + ((g940) & (!g968) & (g1946) & (g1948) & (g2142)) + ((g940) & (g968) & (!g1946) & (!g1948) & (g2142)) + ((g940) & (g968) & (!g1946) & (g1948) & (!g2142)) + ((g940) & (g968) & (!g1946) & (g1948) & (g2142)) + ((g940) & (g968) & (g1946) & (!g1948) & (!g2142)) + ((g940) & (g968) & (g1946) & (!g1948) & (g2142)) + ((g940) & (g968) & (g1946) & (g1948) & (!g2142)) + ((g940) & (g968) & (g1946) & (g1948) & (g2142)));
	assign g2223 = (((!g827) & (!g1007) & (g1953) & (!g2222)) + ((!g827) & (!g1007) & (g1953) & (g2222)) + ((!g827) & (g1007) & (g1953) & (!g2222)) + ((!g827) & (g1007) & (g1953) & (g2222)) + ((g827) & (!g1007) & (!g1953) & (g2222)) + ((g827) & (!g1007) & (g1953) & (!g2222)) + ((g827) & (g1007) & (!g1953) & (!g2222)) + ((g827) & (g1007) & (g1953) & (g2222)));
	assign g7943 = (((!g2017) & (g4439) & (!g2224)) + ((!g2017) & (g4439) & (g2224)) + ((g2017) & (!g4439) & (g2224)) + ((g2017) & (g4439) & (g2224)));
	assign g2225 = (((!g942) & (!g976) & (g2144) & (g2188) & (g2145)) + ((!g942) & (g976) & (!g2144) & (g2188) & (!g2145)) + ((!g942) & (g976) & (!g2144) & (g2188) & (g2145)) + ((!g942) & (g976) & (g2144) & (!g2188) & (g2145)) + ((!g942) & (g976) & (g2144) & (g2188) & (!g2145)) + ((!g942) & (g976) & (g2144) & (g2188) & (g2145)) + ((g942) & (!g976) & (!g2144) & (g2188) & (g2145)) + ((g942) & (!g976) & (g2144) & (g2188) & (!g2145)) + ((g942) & (!g976) & (g2144) & (g2188) & (g2145)) + ((g942) & (g976) & (!g2144) & (!g2188) & (g2145)) + ((g942) & (g976) & (!g2144) & (g2188) & (!g2145)) + ((g942) & (g976) & (!g2144) & (g2188) & (g2145)) + ((g942) & (g976) & (g2144) & (!g2188) & (!g2145)) + ((g942) & (g976) & (g2144) & (!g2188) & (g2145)) + ((g942) & (g976) & (g2144) & (g2188) & (!g2145)) + ((g942) & (g976) & (g2144) & (g2188) & (g2145)));
	assign g2226 = (((!g827) & (!g1009) & (g2224) & (!g2225)) + ((!g827) & (!g1009) & (g2224) & (g2225)) + ((!g827) & (g1009) & (g2224) & (!g2225)) + ((!g827) & (g1009) & (g2224) & (g2225)) + ((g827) & (!g1009) & (!g2224) & (g2225)) + ((g827) & (!g1009) & (g2224) & (!g2225)) + ((g827) & (g1009) & (!g2224) & (!g2225)) + ((g827) & (g1009) & (g2224) & (g2225)));
	assign g7944 = (((!g3499) & (g4442) & (!g2227)) + ((!g3499) & (g4442) & (g2227)) + ((g3499) & (!g4442) & (g2227)) + ((g3499) & (g4442) & (g2227)));
	assign g2228 = (((!g944) & (!g984) & (g2147) & (g2196) & (g2148)) + ((!g944) & (g984) & (!g2147) & (g2196) & (!g2148)) + ((!g944) & (g984) & (!g2147) & (g2196) & (g2148)) + ((!g944) & (g984) & (g2147) & (!g2196) & (g2148)) + ((!g944) & (g984) & (g2147) & (g2196) & (!g2148)) + ((!g944) & (g984) & (g2147) & (g2196) & (g2148)) + ((g944) & (!g984) & (!g2147) & (g2196) & (g2148)) + ((g944) & (!g984) & (g2147) & (g2196) & (!g2148)) + ((g944) & (!g984) & (g2147) & (g2196) & (g2148)) + ((g944) & (g984) & (!g2147) & (!g2196) & (g2148)) + ((g944) & (g984) & (!g2147) & (g2196) & (!g2148)) + ((g944) & (g984) & (!g2147) & (g2196) & (g2148)) + ((g944) & (g984) & (g2147) & (!g2196) & (!g2148)) + ((g944) & (g984) & (g2147) & (!g2196) & (g2148)) + ((g944) & (g984) & (g2147) & (g2196) & (!g2148)) + ((g944) & (g984) & (g2147) & (g2196) & (g2148)));
	assign g2229 = (((!g827) & (!g1011) & (g2227) & (!g2228)) + ((!g827) & (!g1011) & (g2227) & (g2228)) + ((!g827) & (g1011) & (g2227) & (!g2228)) + ((!g827) & (g1011) & (g2227) & (g2228)) + ((g827) & (!g1011) & (!g2227) & (g2228)) + ((g827) & (!g1011) & (g2227) & (!g2228)) + ((g827) & (g1011) & (!g2227) & (!g2228)) + ((g827) & (g1011) & (g2227) & (g2228)));
	assign g7945 = (((!g3464) & (g4445) & (!g2230)) + ((!g3464) & (g4445) & (g2230)) + ((g3464) & (!g4445) & (g2230)) + ((g3464) & (g4445) & (g2230)));
	assign g2231 = (((!g946) & (!g992) & (g2150) & (g2203) & (g2151)) + ((!g946) & (g992) & (!g2150) & (g2203) & (!g2151)) + ((!g946) & (g992) & (!g2150) & (g2203) & (g2151)) + ((!g946) & (g992) & (g2150) & (!g2203) & (g2151)) + ((!g946) & (g992) & (g2150) & (g2203) & (!g2151)) + ((!g946) & (g992) & (g2150) & (g2203) & (g2151)) + ((g946) & (!g992) & (!g2150) & (g2203) & (g2151)) + ((g946) & (!g992) & (g2150) & (g2203) & (!g2151)) + ((g946) & (!g992) & (g2150) & (g2203) & (g2151)) + ((g946) & (g992) & (!g2150) & (!g2203) & (g2151)) + ((g946) & (g992) & (!g2150) & (g2203) & (!g2151)) + ((g946) & (g992) & (!g2150) & (g2203) & (g2151)) + ((g946) & (g992) & (g2150) & (!g2203) & (!g2151)) + ((g946) & (g992) & (g2150) & (!g2203) & (g2151)) + ((g946) & (g992) & (g2150) & (g2203) & (!g2151)) + ((g946) & (g992) & (g2150) & (g2203) & (g2151)));
	assign g2232 = (((!g827) & (!g1013) & (g2230) & (!g2231)) + ((!g827) & (!g1013) & (g2230) & (g2231)) + ((!g827) & (g1013) & (g2230) & (!g2231)) + ((!g827) & (g1013) & (g2230) & (g2231)) + ((g827) & (!g1013) & (!g2230) & (g2231)) + ((g827) & (!g1013) & (g2230) & (!g2231)) + ((g827) & (g1013) & (!g2230) & (!g2231)) + ((g827) & (g1013) & (g2230) & (g2231)));
	assign g7946 = (((!g3499) & (g4448) & (!g2233)) + ((!g3499) & (g4448) & (g2233)) + ((g3499) & (!g4448) & (g2233)) + ((g3499) & (g4448) & (g2233)));
	assign g2234 = (((!g948) & (!g970) & (g2153) & (g2184) & (g2154)) + ((!g948) & (g970) & (!g2153) & (g2184) & (!g2154)) + ((!g948) & (g970) & (!g2153) & (g2184) & (g2154)) + ((!g948) & (g970) & (g2153) & (!g2184) & (g2154)) + ((!g948) & (g970) & (g2153) & (g2184) & (!g2154)) + ((!g948) & (g970) & (g2153) & (g2184) & (g2154)) + ((g948) & (!g970) & (!g2153) & (g2184) & (g2154)) + ((g948) & (!g970) & (g2153) & (g2184) & (!g2154)) + ((g948) & (!g970) & (g2153) & (g2184) & (g2154)) + ((g948) & (g970) & (!g2153) & (!g2184) & (g2154)) + ((g948) & (g970) & (!g2153) & (g2184) & (!g2154)) + ((g948) & (g970) & (!g2153) & (g2184) & (g2154)) + ((g948) & (g970) & (g2153) & (!g2184) & (!g2154)) + ((g948) & (g970) & (g2153) & (!g2184) & (g2154)) + ((g948) & (g970) & (g2153) & (g2184) & (!g2154)) + ((g948) & (g970) & (g2153) & (g2184) & (g2154)));
	assign g2235 = (((!g827) & (!g1015) & (g2233) & (!g2234)) + ((!g827) & (!g1015) & (g2233) & (g2234)) + ((!g827) & (g1015) & (g2233) & (!g2234)) + ((!g827) & (g1015) & (g2233) & (g2234)) + ((g827) & (!g1015) & (!g2233) & (g2234)) + ((g827) & (!g1015) & (g2233) & (!g2234)) + ((g827) & (g1015) & (!g2233) & (!g2234)) + ((g827) & (g1015) & (g2233) & (g2234)));
	assign g7947 = (((!g3464) & (g4452) & (!g2236)) + ((!g3464) & (g4452) & (g2236)) + ((g3464) & (!g4452) & (g2236)) + ((g3464) & (g4452) & (g2236)));
	assign g2237 = (((!g950) & (!g978) & (g2156) & (g2190) & (g2157)) + ((!g950) & (g978) & (!g2156) & (g2190) & (!g2157)) + ((!g950) & (g978) & (!g2156) & (g2190) & (g2157)) + ((!g950) & (g978) & (g2156) & (!g2190) & (g2157)) + ((!g950) & (g978) & (g2156) & (g2190) & (!g2157)) + ((!g950) & (g978) & (g2156) & (g2190) & (g2157)) + ((g950) & (!g978) & (!g2156) & (g2190) & (g2157)) + ((g950) & (!g978) & (g2156) & (g2190) & (!g2157)) + ((g950) & (!g978) & (g2156) & (g2190) & (g2157)) + ((g950) & (g978) & (!g2156) & (!g2190) & (g2157)) + ((g950) & (g978) & (!g2156) & (g2190) & (!g2157)) + ((g950) & (g978) & (!g2156) & (g2190) & (g2157)) + ((g950) & (g978) & (g2156) & (!g2190) & (!g2157)) + ((g950) & (g978) & (g2156) & (!g2190) & (g2157)) + ((g950) & (g978) & (g2156) & (g2190) & (!g2157)) + ((g950) & (g978) & (g2156) & (g2190) & (g2157)));
	assign g2238 = (((!g827) & (!g1017) & (g2236) & (!g2237)) + ((!g827) & (!g1017) & (g2236) & (g2237)) + ((!g827) & (g1017) & (g2236) & (!g2237)) + ((!g827) & (g1017) & (g2236) & (g2237)) + ((g827) & (!g1017) & (!g2236) & (g2237)) + ((g827) & (!g1017) & (g2236) & (!g2237)) + ((g827) & (g1017) & (!g2236) & (!g2237)) + ((g827) & (g1017) & (g2236) & (g2237)));
	assign g7948 = (((!g2017) & (g4457) & (!g2239)) + ((!g2017) & (g4457) & (g2239)) + ((g2017) & (!g4457) & (g2239)) + ((g2017) & (g4457) & (g2239)));
	assign g2240 = (((!g952) & (!g986) & (g2159) & (g2198) & (g2160)) + ((!g952) & (g986) & (!g2159) & (g2198) & (!g2160)) + ((!g952) & (g986) & (!g2159) & (g2198) & (g2160)) + ((!g952) & (g986) & (g2159) & (!g2198) & (g2160)) + ((!g952) & (g986) & (g2159) & (g2198) & (!g2160)) + ((!g952) & (g986) & (g2159) & (g2198) & (g2160)) + ((g952) & (!g986) & (!g2159) & (g2198) & (g2160)) + ((g952) & (!g986) & (g2159) & (g2198) & (!g2160)) + ((g952) & (!g986) & (g2159) & (g2198) & (g2160)) + ((g952) & (g986) & (!g2159) & (!g2198) & (g2160)) + ((g952) & (g986) & (!g2159) & (g2198) & (!g2160)) + ((g952) & (g986) & (!g2159) & (g2198) & (g2160)) + ((g952) & (g986) & (g2159) & (!g2198) & (!g2160)) + ((g952) & (g986) & (g2159) & (!g2198) & (g2160)) + ((g952) & (g986) & (g2159) & (g2198) & (!g2160)) + ((g952) & (g986) & (g2159) & (g2198) & (g2160)));
	assign g2241 = (((!g827) & (!g1019) & (g2239) & (!g2240)) + ((!g827) & (!g1019) & (g2239) & (g2240)) + ((!g827) & (g1019) & (g2239) & (!g2240)) + ((!g827) & (g1019) & (g2239) & (g2240)) + ((g827) & (!g1019) & (!g2239) & (g2240)) + ((g827) & (!g1019) & (g2239) & (!g2240)) + ((g827) & (g1019) & (!g2239) & (!g2240)) + ((g827) & (g1019) & (g2239) & (g2240)));
	assign g7949 = (((!g3429) & (g4460) & (!g2242)) + ((!g3429) & (g4460) & (g2242)) + ((g3429) & (!g4460) & (g2242)) + ((g3429) & (g4460) & (g2242)));
	assign g2243 = (((!g954) & (!g994) & (g2162) & (g2205) & (g2163)) + ((!g954) & (g994) & (!g2162) & (g2205) & (!g2163)) + ((!g954) & (g994) & (!g2162) & (g2205) & (g2163)) + ((!g954) & (g994) & (g2162) & (!g2205) & (g2163)) + ((!g954) & (g994) & (g2162) & (g2205) & (!g2163)) + ((!g954) & (g994) & (g2162) & (g2205) & (g2163)) + ((g954) & (!g994) & (!g2162) & (g2205) & (g2163)) + ((g954) & (!g994) & (g2162) & (g2205) & (!g2163)) + ((g954) & (!g994) & (g2162) & (g2205) & (g2163)) + ((g954) & (g994) & (!g2162) & (!g2205) & (g2163)) + ((g954) & (g994) & (!g2162) & (g2205) & (!g2163)) + ((g954) & (g994) & (!g2162) & (g2205) & (g2163)) + ((g954) & (g994) & (g2162) & (!g2205) & (!g2163)) + ((g954) & (g994) & (g2162) & (!g2205) & (g2163)) + ((g954) & (g994) & (g2162) & (g2205) & (!g2163)) + ((g954) & (g994) & (g2162) & (g2205) & (g2163)));
	assign g2244 = (((!g827) & (!g1021) & (g2242) & (!g2243)) + ((!g827) & (!g1021) & (g2242) & (g2243)) + ((!g827) & (g1021) & (g2242) & (!g2243)) + ((!g827) & (g1021) & (g2242) & (g2243)) + ((g827) & (!g1021) & (!g2242) & (g2243)) + ((g827) & (!g1021) & (g2242) & (!g2243)) + ((g827) & (g1021) & (!g2242) & (!g2243)) + ((g827) & (g1021) & (g2242) & (g2243)));
	assign g2245 = (((!g956) & (!g972) & (g1947) & (g1949) & (g2165)) + ((!g956) & (g972) & (!g1947) & (g1949) & (!g2165)) + ((!g956) & (g972) & (!g1947) & (g1949) & (g2165)) + ((!g956) & (g972) & (g1947) & (!g1949) & (g2165)) + ((!g956) & (g972) & (g1947) & (g1949) & (!g2165)) + ((!g956) & (g972) & (g1947) & (g1949) & (g2165)) + ((g956) & (!g972) & (!g1947) & (g1949) & (g2165)) + ((g956) & (!g972) & (g1947) & (g1949) & (!g2165)) + ((g956) & (!g972) & (g1947) & (g1949) & (g2165)) + ((g956) & (g972) & (!g1947) & (!g1949) & (g2165)) + ((g956) & (g972) & (!g1947) & (g1949) & (!g2165)) + ((g956) & (g972) & (!g1947) & (g1949) & (g2165)) + ((g956) & (g972) & (g1947) & (!g1949) & (!g2165)) + ((g956) & (g972) & (g1947) & (!g1949) & (g2165)) + ((g956) & (g972) & (g1947) & (g1949) & (!g2165)) + ((g956) & (g972) & (g1947) & (g1949) & (g2165)));
	assign g2246 = (((!g827) & (!g1023) & (g1954) & (!g2245)) + ((!g827) & (!g1023) & (g1954) & (g2245)) + ((!g827) & (g1023) & (g1954) & (!g2245)) + ((!g827) & (g1023) & (g1954) & (g2245)) + ((g827) & (!g1023) & (!g1954) & (g2245)) + ((g827) & (!g1023) & (g1954) & (!g2245)) + ((g827) & (g1023) & (!g1954) & (!g2245)) + ((g827) & (g1023) & (g1954) & (g2245)));
	assign g7950 = (((!g3499) & (g4463) & (!g2247)) + ((!g3499) & (g4463) & (g2247)) + ((g3499) & (!g4463) & (g2247)) + ((g3499) & (g4463) & (g2247)));
	assign g2248 = (((!g958) & (!g980) & (g2167) & (g2192) & (g2168)) + ((!g958) & (g980) & (!g2167) & (g2192) & (!g2168)) + ((!g958) & (g980) & (!g2167) & (g2192) & (g2168)) + ((!g958) & (g980) & (g2167) & (!g2192) & (g2168)) + ((!g958) & (g980) & (g2167) & (g2192) & (!g2168)) + ((!g958) & (g980) & (g2167) & (g2192) & (g2168)) + ((g958) & (!g980) & (!g2167) & (g2192) & (g2168)) + ((g958) & (!g980) & (g2167) & (g2192) & (!g2168)) + ((g958) & (!g980) & (g2167) & (g2192) & (g2168)) + ((g958) & (g980) & (!g2167) & (!g2192) & (g2168)) + ((g958) & (g980) & (!g2167) & (g2192) & (!g2168)) + ((g958) & (g980) & (!g2167) & (g2192) & (g2168)) + ((g958) & (g980) & (g2167) & (!g2192) & (!g2168)) + ((g958) & (g980) & (g2167) & (!g2192) & (g2168)) + ((g958) & (g980) & (g2167) & (g2192) & (!g2168)) + ((g958) & (g980) & (g2167) & (g2192) & (g2168)));
	assign g2249 = (((!g827) & (!g1025) & (g2247) & (!g2248)) + ((!g827) & (!g1025) & (g2247) & (g2248)) + ((!g827) & (g1025) & (g2247) & (!g2248)) + ((!g827) & (g1025) & (g2247) & (g2248)) + ((g827) & (!g1025) & (!g2247) & (g2248)) + ((g827) & (!g1025) & (g2247) & (!g2248)) + ((g827) & (g1025) & (!g2247) & (!g2248)) + ((g827) & (g1025) & (g2247) & (g2248)));
	assign g7951 = (((!g3429) & (g4466) & (!g2250)) + ((!g3429) & (g4466) & (g2250)) + ((g3429) & (!g4466) & (g2250)) + ((g3429) & (g4466) & (g2250)));
	assign g2251 = (((!g960) & (!g988) & (g2170) & (g2200) & (g2171)) + ((!g960) & (g988) & (!g2170) & (g2200) & (!g2171)) + ((!g960) & (g988) & (!g2170) & (g2200) & (g2171)) + ((!g960) & (g988) & (g2170) & (!g2200) & (g2171)) + ((!g960) & (g988) & (g2170) & (g2200) & (!g2171)) + ((!g960) & (g988) & (g2170) & (g2200) & (g2171)) + ((g960) & (!g988) & (!g2170) & (g2200) & (g2171)) + ((g960) & (!g988) & (g2170) & (g2200) & (!g2171)) + ((g960) & (!g988) & (g2170) & (g2200) & (g2171)) + ((g960) & (g988) & (!g2170) & (!g2200) & (g2171)) + ((g960) & (g988) & (!g2170) & (g2200) & (!g2171)) + ((g960) & (g988) & (!g2170) & (g2200) & (g2171)) + ((g960) & (g988) & (g2170) & (!g2200) & (!g2171)) + ((g960) & (g988) & (g2170) & (!g2200) & (g2171)) + ((g960) & (g988) & (g2170) & (g2200) & (!g2171)) + ((g960) & (g988) & (g2170) & (g2200) & (g2171)));
	assign g2252 = (((!g827) & (!g1027) & (g2250) & (!g2251)) + ((!g827) & (!g1027) & (g2250) & (g2251)) + ((!g827) & (g1027) & (g2250) & (!g2251)) + ((!g827) & (g1027) & (g2250) & (g2251)) + ((g827) & (!g1027) & (!g2250) & (g2251)) + ((g827) & (!g1027) & (g2250) & (!g2251)) + ((g827) & (g1027) & (!g2250) & (!g2251)) + ((g827) & (g1027) & (g2250) & (g2251)));
	assign g7952 = (((!g2017) & (g4471) & (!g2253)) + ((!g2017) & (g4471) & (g2253)) + ((g2017) & (!g4471) & (g2253)) + ((g2017) & (g4471) & (g2253)));
	assign g2254 = (((!g962) & (!g996) & (g2173) & (g2207) & (g2174)) + ((!g962) & (g996) & (!g2173) & (g2207) & (!g2174)) + ((!g962) & (g996) & (!g2173) & (g2207) & (g2174)) + ((!g962) & (g996) & (g2173) & (!g2207) & (g2174)) + ((!g962) & (g996) & (g2173) & (g2207) & (!g2174)) + ((!g962) & (g996) & (g2173) & (g2207) & (g2174)) + ((g962) & (!g996) & (!g2173) & (g2207) & (g2174)) + ((g962) & (!g996) & (g2173) & (g2207) & (!g2174)) + ((g962) & (!g996) & (g2173) & (g2207) & (g2174)) + ((g962) & (g996) & (!g2173) & (!g2207) & (g2174)) + ((g962) & (g996) & (!g2173) & (g2207) & (!g2174)) + ((g962) & (g996) & (!g2173) & (g2207) & (g2174)) + ((g962) & (g996) & (g2173) & (!g2207) & (!g2174)) + ((g962) & (g996) & (g2173) & (!g2207) & (g2174)) + ((g962) & (g996) & (g2173) & (g2207) & (!g2174)) + ((g962) & (g996) & (g2173) & (g2207) & (g2174)));
	assign g2255 = (((!g827) & (!g1029) & (g2253) & (!g2254)) + ((!g827) & (!g1029) & (g2253) & (g2254)) + ((!g827) & (g1029) & (g2253) & (!g2254)) + ((!g827) & (g1029) & (g2253) & (g2254)) + ((g827) & (!g1029) & (!g2253) & (g2254)) + ((g827) & (!g1029) & (g2253) & (!g2254)) + ((g827) & (g1029) & (!g2253) & (!g2254)) + ((g827) & (g1029) & (g2253) & (g2254)));
	assign g7953 = (((!g3429) & (g4476) & (!g2256)) + ((!g3429) & (g4476) & (g2256)) + ((g3429) & (!g4476) & (g2256)) + ((g3429) & (g4476) & (g2256)));
	assign g7954 = (((!g3464) & (g4479) & (!g2257)) + ((!g3464) & (g4479) & (g2257)) + ((g3464) & (!g4479) & (g2257)) + ((g3464) & (g4479) & (g2257)));
	assign g2258 = (((!g2209) & (!g2210) & (!g2211) & (!g2256) & (g2257)) + ((!g2209) & (!g2210) & (!g2211) & (g2256) & (!g2257)) + ((!g2209) & (!g2210) & (g2211) & (!g2256) & (g2257)) + ((!g2209) & (!g2210) & (g2211) & (g2256) & (!g2257)) + ((!g2209) & (g2210) & (!g2211) & (!g2256) & (g2257)) + ((!g2209) & (g2210) & (!g2211) & (g2256) & (!g2257)) + ((!g2209) & (g2210) & (g2211) & (!g2256) & (!g2257)) + ((!g2209) & (g2210) & (g2211) & (g2256) & (g2257)) + ((g2209) & (!g2210) & (!g2211) & (!g2256) & (g2257)) + ((g2209) & (!g2210) & (!g2211) & (g2256) & (!g2257)) + ((g2209) & (!g2210) & (g2211) & (!g2256) & (!g2257)) + ((g2209) & (!g2210) & (g2211) & (g2256) & (g2257)) + ((g2209) & (g2210) & (!g2211) & (!g2256) & (!g2257)) + ((g2209) & (g2210) & (!g2211) & (g2256) & (g2257)) + ((g2209) & (g2210) & (g2211) & (!g2256) & (!g2257)) + ((g2209) & (g2210) & (g2211) & (g2256) & (g2257)));
	assign g2259 = (((!g2212) & (g2213)) + ((g2212) & (!g2213)));
	assign g2260 = (((!g2132) & (!g2133) & (!g2134) & (g2180) & (g2181) & (g2259)) + ((!g2132) & (!g2133) & (g2134) & (g2180) & (g2181) & (g2259)) + ((!g2132) & (g2133) & (!g2134) & (g2180) & (g2181) & (g2259)) + ((!g2132) & (g2133) & (g2134) & (!g2180) & (g2181) & (g2259)) + ((!g2132) & (g2133) & (g2134) & (g2180) & (!g2181) & (g2259)) + ((!g2132) & (g2133) & (g2134) & (g2180) & (g2181) & (g2259)) + ((g2132) & (!g2133) & (!g2134) & (g2180) & (g2181) & (g2259)) + ((g2132) & (!g2133) & (g2134) & (!g2180) & (g2181) & (g2259)) + ((g2132) & (!g2133) & (g2134) & (g2180) & (!g2181) & (g2259)) + ((g2132) & (!g2133) & (g2134) & (g2180) & (g2181) & (g2259)) + ((g2132) & (g2133) & (!g2134) & (!g2180) & (g2181) & (g2259)) + ((g2132) & (g2133) & (!g2134) & (g2180) & (!g2181) & (g2259)) + ((g2132) & (g2133) & (!g2134) & (g2180) & (g2181) & (g2259)) + ((g2132) & (g2133) & (g2134) & (!g2180) & (g2181) & (g2259)) + ((g2132) & (g2133) & (g2134) & (g2180) & (!g2181) & (g2259)) + ((g2132) & (g2133) & (g2134) & (g2180) & (g2181) & (g2259)));
	assign g2261 = (((g2212) & (g2213)));
	assign g7955 = (((!g3429) & (g4483) & (!g2262)) + ((!g3429) & (g4483) & (g2262)) + ((g3429) & (!g4483) & (g2262)) + ((g3429) & (g4483) & (g2262)));
	assign g7956 = (((!g3499) & (g4486) & (!g2263)) + ((!g3499) & (g4486) & (g2263)) + ((g3499) & (!g4486) & (g2263)) + ((g3499) & (g4486) & (g2263)));
	assign g2264 = (((!g2260) & (!g2261) & (!g2262) & (g2263)) + ((!g2260) & (!g2261) & (g2262) & (!g2263)) + ((!g2260) & (g2261) & (!g2262) & (!g2263)) + ((!g2260) & (g2261) & (g2262) & (g2263)) + ((g2260) & (!g2261) & (!g2262) & (!g2263)) + ((g2260) & (!g2261) & (g2262) & (g2263)) + ((g2260) & (g2261) & (!g2262) & (!g2263)) + ((g2260) & (g2261) & (g2262) & (g2263)));
	assign g2265 = (((!g830) & (!g1914) & (!g2258) & (!g2264) & (!g1031)) + ((!g830) & (!g1914) & (!g2258) & (!g2264) & (g1031)) + ((!g830) & (!g1914) & (!g2258) & (g2264) & (!g1031)) + ((!g830) & (!g1914) & (!g2258) & (g2264) & (g1031)) + ((!g830) & (!g1914) & (g2258) & (!g2264) & (!g1031)) + ((!g830) & (!g1914) & (g2258) & (!g2264) & (g1031)) + ((!g830) & (!g1914) & (g2258) & (g2264) & (!g1031)) + ((!g830) & (!g1914) & (g2258) & (g2264) & (g1031)) + ((!g830) & (g1914) & (!g2258) & (!g2264) & (!g1031)) + ((!g830) & (g1914) & (!g2258) & (!g2264) & (g1031)) + ((!g830) & (g1914) & (!g2258) & (g2264) & (!g1031)) + ((!g830) & (g1914) & (!g2258) & (g2264) & (g1031)) + ((!g830) & (g1914) & (g2258) & (!g2264) & (!g1031)) + ((!g830) & (g1914) & (g2258) & (!g2264) & (g1031)) + ((!g830) & (g1914) & (g2258) & (g2264) & (!g1031)) + ((!g830) & (g1914) & (g2258) & (g2264) & (g1031)) + ((g830) & (!g1914) & (!g2258) & (!g2264) & (g1031)) + ((g830) & (!g1914) & (!g2258) & (g2264) & (!g1031)) + ((g830) & (!g1914) & (g2258) & (!g2264) & (g1031)) + ((g830) & (!g1914) & (g2258) & (g2264) & (!g1031)) + ((g830) & (g1914) & (!g2258) & (!g2264) & (g1031)) + ((g830) & (g1914) & (!g2258) & (g2264) & (g1031)) + ((g830) & (g1914) & (g2258) & (!g2264) & (!g1031)) + ((g830) & (g1914) & (g2258) & (g2264) & (!g1031)));
	assign g2266 = (((!g827) & (!g1007) & (!g1035) & (!g1953) & (g1955) & (!g2222)) + ((!g827) & (!g1007) & (!g1035) & (!g1953) & (g1955) & (g2222)) + ((!g827) & (!g1007) & (!g1035) & (g1953) & (g1955) & (!g2222)) + ((!g827) & (!g1007) & (!g1035) & (g1953) & (g1955) & (g2222)) + ((!g827) & (!g1007) & (g1035) & (!g1953) & (g1955) & (!g2222)) + ((!g827) & (!g1007) & (g1035) & (!g1953) & (g1955) & (g2222)) + ((!g827) & (!g1007) & (g1035) & (g1953) & (g1955) & (!g2222)) + ((!g827) & (!g1007) & (g1035) & (g1953) & (g1955) & (g2222)) + ((!g827) & (g1007) & (!g1035) & (!g1953) & (g1955) & (!g2222)) + ((!g827) & (g1007) & (!g1035) & (!g1953) & (g1955) & (g2222)) + ((!g827) & (g1007) & (!g1035) & (g1953) & (g1955) & (!g2222)) + ((!g827) & (g1007) & (!g1035) & (g1953) & (g1955) & (g2222)) + ((!g827) & (g1007) & (g1035) & (!g1953) & (g1955) & (!g2222)) + ((!g827) & (g1007) & (g1035) & (!g1953) & (g1955) & (g2222)) + ((!g827) & (g1007) & (g1035) & (g1953) & (g1955) & (!g2222)) + ((!g827) & (g1007) & (g1035) & (g1953) & (g1955) & (g2222)) + ((g827) & (!g1007) & (!g1035) & (!g1953) & (g1955) & (!g2222)) + ((g827) & (!g1007) & (!g1035) & (!g1953) & (g1955) & (g2222)) + ((g827) & (!g1007) & (!g1035) & (g1953) & (!g1955) & (g2222)) + ((g827) & (!g1007) & (!g1035) & (g1953) & (g1955) & (!g2222)) + ((g827) & (!g1007) & (g1035) & (!g1953) & (!g1955) & (!g2222)) + ((g827) & (!g1007) & (g1035) & (!g1953) & (!g1955) & (g2222)) + ((g827) & (!g1007) & (g1035) & (g1953) & (!g1955) & (!g2222)) + ((g827) & (!g1007) & (g1035) & (g1953) & (g1955) & (g2222)) + ((g827) & (g1007) & (!g1035) & (!g1953) & (!g1955) & (g2222)) + ((g827) & (g1007) & (!g1035) & (!g1953) & (g1955) & (!g2222)) + ((g827) & (g1007) & (!g1035) & (g1953) & (!g1955) & (!g2222)) + ((g827) & (g1007) & (!g1035) & (g1953) & (!g1955) & (g2222)) + ((g827) & (g1007) & (g1035) & (!g1953) & (!g1955) & (!g2222)) + ((g827) & (g1007) & (g1035) & (!g1953) & (g1955) & (g2222)) + ((g827) & (g1007) & (g1035) & (g1953) & (g1955) & (!g2222)) + ((g827) & (g1007) & (g1035) & (g1953) & (g1955) & (g2222)));
	assign g7957 = (((!g3499) & (g6713) & (!g2267)) + ((!g3499) & (g6713) & (g2267)) + ((g3499) & (!g6713) & (g2267)) + ((g3499) & (g6713) & (g2267)));
	assign g2268 = (((!g827) & (!g1015) & (!g1037) & (!g2233) & (g2267) & (!g2234)) + ((!g827) & (!g1015) & (!g1037) & (!g2233) & (g2267) & (g2234)) + ((!g827) & (!g1015) & (!g1037) & (g2233) & (g2267) & (!g2234)) + ((!g827) & (!g1015) & (!g1037) & (g2233) & (g2267) & (g2234)) + ((!g827) & (!g1015) & (g1037) & (!g2233) & (g2267) & (!g2234)) + ((!g827) & (!g1015) & (g1037) & (!g2233) & (g2267) & (g2234)) + ((!g827) & (!g1015) & (g1037) & (g2233) & (g2267) & (!g2234)) + ((!g827) & (!g1015) & (g1037) & (g2233) & (g2267) & (g2234)) + ((!g827) & (g1015) & (!g1037) & (!g2233) & (g2267) & (!g2234)) + ((!g827) & (g1015) & (!g1037) & (!g2233) & (g2267) & (g2234)) + ((!g827) & (g1015) & (!g1037) & (g2233) & (g2267) & (!g2234)) + ((!g827) & (g1015) & (!g1037) & (g2233) & (g2267) & (g2234)) + ((!g827) & (g1015) & (g1037) & (!g2233) & (g2267) & (!g2234)) + ((!g827) & (g1015) & (g1037) & (!g2233) & (g2267) & (g2234)) + ((!g827) & (g1015) & (g1037) & (g2233) & (g2267) & (!g2234)) + ((!g827) & (g1015) & (g1037) & (g2233) & (g2267) & (g2234)) + ((g827) & (!g1015) & (!g1037) & (!g2233) & (g2267) & (!g2234)) + ((g827) & (!g1015) & (!g1037) & (!g2233) & (g2267) & (g2234)) + ((g827) & (!g1015) & (!g1037) & (g2233) & (!g2267) & (g2234)) + ((g827) & (!g1015) & (!g1037) & (g2233) & (g2267) & (!g2234)) + ((g827) & (!g1015) & (g1037) & (!g2233) & (!g2267) & (!g2234)) + ((g827) & (!g1015) & (g1037) & (!g2233) & (!g2267) & (g2234)) + ((g827) & (!g1015) & (g1037) & (g2233) & (!g2267) & (!g2234)) + ((g827) & (!g1015) & (g1037) & (g2233) & (g2267) & (g2234)) + ((g827) & (g1015) & (!g1037) & (!g2233) & (!g2267) & (g2234)) + ((g827) & (g1015) & (!g1037) & (!g2233) & (g2267) & (!g2234)) + ((g827) & (g1015) & (!g1037) & (g2233) & (!g2267) & (!g2234)) + ((g827) & (g1015) & (!g1037) & (g2233) & (!g2267) & (g2234)) + ((g827) & (g1015) & (g1037) & (!g2233) & (!g2267) & (!g2234)) + ((g827) & (g1015) & (g1037) & (!g2233) & (g2267) & (g2234)) + ((g827) & (g1015) & (g1037) & (g2233) & (g2267) & (!g2234)) + ((g827) & (g1015) & (g1037) & (g2233) & (g2267) & (g2234)));
	assign g2269 = (((!g827) & (!g1023) & (!g1039) & (!g1954) & (g1956) & (!g2245)) + ((!g827) & (!g1023) & (!g1039) & (!g1954) & (g1956) & (g2245)) + ((!g827) & (!g1023) & (!g1039) & (g1954) & (g1956) & (!g2245)) + ((!g827) & (!g1023) & (!g1039) & (g1954) & (g1956) & (g2245)) + ((!g827) & (!g1023) & (g1039) & (!g1954) & (g1956) & (!g2245)) + ((!g827) & (!g1023) & (g1039) & (!g1954) & (g1956) & (g2245)) + ((!g827) & (!g1023) & (g1039) & (g1954) & (g1956) & (!g2245)) + ((!g827) & (!g1023) & (g1039) & (g1954) & (g1956) & (g2245)) + ((!g827) & (g1023) & (!g1039) & (!g1954) & (g1956) & (!g2245)) + ((!g827) & (g1023) & (!g1039) & (!g1954) & (g1956) & (g2245)) + ((!g827) & (g1023) & (!g1039) & (g1954) & (g1956) & (!g2245)) + ((!g827) & (g1023) & (!g1039) & (g1954) & (g1956) & (g2245)) + ((!g827) & (g1023) & (g1039) & (!g1954) & (g1956) & (!g2245)) + ((!g827) & (g1023) & (g1039) & (!g1954) & (g1956) & (g2245)) + ((!g827) & (g1023) & (g1039) & (g1954) & (g1956) & (!g2245)) + ((!g827) & (g1023) & (g1039) & (g1954) & (g1956) & (g2245)) + ((g827) & (!g1023) & (!g1039) & (!g1954) & (g1956) & (!g2245)) + ((g827) & (!g1023) & (!g1039) & (!g1954) & (g1956) & (g2245)) + ((g827) & (!g1023) & (!g1039) & (g1954) & (!g1956) & (g2245)) + ((g827) & (!g1023) & (!g1039) & (g1954) & (g1956) & (!g2245)) + ((g827) & (!g1023) & (g1039) & (!g1954) & (!g1956) & (!g2245)) + ((g827) & (!g1023) & (g1039) & (!g1954) & (!g1956) & (g2245)) + ((g827) & (!g1023) & (g1039) & (g1954) & (!g1956) & (!g2245)) + ((g827) & (!g1023) & (g1039) & (g1954) & (g1956) & (g2245)) + ((g827) & (g1023) & (!g1039) & (!g1954) & (!g1956) & (g2245)) + ((g827) & (g1023) & (!g1039) & (!g1954) & (g1956) & (!g2245)) + ((g827) & (g1023) & (!g1039) & (g1954) & (!g1956) & (!g2245)) + ((g827) & (g1023) & (!g1039) & (g1954) & (!g1956) & (g2245)) + ((g827) & (g1023) & (g1039) & (!g1954) & (!g1956) & (!g2245)) + ((g827) & (g1023) & (g1039) & (!g1954) & (g1956) & (g2245)) + ((g827) & (g1023) & (g1039) & (g1954) & (g1956) & (!g2245)) + ((g827) & (g1023) & (g1039) & (g1954) & (g1956) & (g2245)));
	assign g2270 = (((!g827) & (!g1001) & (!g1041) & (!g1991) & (g1993) & (!g2215)) + ((!g827) & (!g1001) & (!g1041) & (!g1991) & (g1993) & (g2215)) + ((!g827) & (!g1001) & (!g1041) & (g1991) & (g1993) & (!g2215)) + ((!g827) & (!g1001) & (!g1041) & (g1991) & (g1993) & (g2215)) + ((!g827) & (!g1001) & (g1041) & (!g1991) & (g1993) & (!g2215)) + ((!g827) & (!g1001) & (g1041) & (!g1991) & (g1993) & (g2215)) + ((!g827) & (!g1001) & (g1041) & (g1991) & (g1993) & (!g2215)) + ((!g827) & (!g1001) & (g1041) & (g1991) & (g1993) & (g2215)) + ((!g827) & (g1001) & (!g1041) & (!g1991) & (g1993) & (!g2215)) + ((!g827) & (g1001) & (!g1041) & (!g1991) & (g1993) & (g2215)) + ((!g827) & (g1001) & (!g1041) & (g1991) & (g1993) & (!g2215)) + ((!g827) & (g1001) & (!g1041) & (g1991) & (g1993) & (g2215)) + ((!g827) & (g1001) & (g1041) & (!g1991) & (g1993) & (!g2215)) + ((!g827) & (g1001) & (g1041) & (!g1991) & (g1993) & (g2215)) + ((!g827) & (g1001) & (g1041) & (g1991) & (g1993) & (!g2215)) + ((!g827) & (g1001) & (g1041) & (g1991) & (g1993) & (g2215)) + ((g827) & (!g1001) & (!g1041) & (!g1991) & (g1993) & (!g2215)) + ((g827) & (!g1001) & (!g1041) & (!g1991) & (g1993) & (g2215)) + ((g827) & (!g1001) & (!g1041) & (g1991) & (!g1993) & (g2215)) + ((g827) & (!g1001) & (!g1041) & (g1991) & (g1993) & (!g2215)) + ((g827) & (!g1001) & (g1041) & (!g1991) & (!g1993) & (!g2215)) + ((g827) & (!g1001) & (g1041) & (!g1991) & (!g1993) & (g2215)) + ((g827) & (!g1001) & (g1041) & (g1991) & (!g1993) & (!g2215)) + ((g827) & (!g1001) & (g1041) & (g1991) & (g1993) & (g2215)) + ((g827) & (g1001) & (!g1041) & (!g1991) & (!g1993) & (g2215)) + ((g827) & (g1001) & (!g1041) & (!g1991) & (g1993) & (!g2215)) + ((g827) & (g1001) & (!g1041) & (g1991) & (!g1993) & (!g2215)) + ((g827) & (g1001) & (!g1041) & (g1991) & (!g1993) & (g2215)) + ((g827) & (g1001) & (g1041) & (!g1991) & (!g1993) & (!g2215)) + ((g827) & (g1001) & (g1041) & (!g1991) & (g1993) & (g2215)) + ((g827) & (g1001) & (g1041) & (g1991) & (g1993) & (!g2215)) + ((g827) & (g1001) & (g1041) & (g1991) & (g1993) & (g2215)));
	assign g7958 = (((!g2017) & (g4496) & (!g2271)) + ((!g2017) & (g4496) & (g2271)) + ((g2017) & (!g4496) & (g2271)) + ((g2017) & (g4496) & (g2271)));
	assign g2272 = (((!g827) & (!g1009) & (!g1043) & (!g2224) & (g2271) & (!g2225)) + ((!g827) & (!g1009) & (!g1043) & (!g2224) & (g2271) & (g2225)) + ((!g827) & (!g1009) & (!g1043) & (g2224) & (g2271) & (!g2225)) + ((!g827) & (!g1009) & (!g1043) & (g2224) & (g2271) & (g2225)) + ((!g827) & (!g1009) & (g1043) & (!g2224) & (g2271) & (!g2225)) + ((!g827) & (!g1009) & (g1043) & (!g2224) & (g2271) & (g2225)) + ((!g827) & (!g1009) & (g1043) & (g2224) & (g2271) & (!g2225)) + ((!g827) & (!g1009) & (g1043) & (g2224) & (g2271) & (g2225)) + ((!g827) & (g1009) & (!g1043) & (!g2224) & (g2271) & (!g2225)) + ((!g827) & (g1009) & (!g1043) & (!g2224) & (g2271) & (g2225)) + ((!g827) & (g1009) & (!g1043) & (g2224) & (g2271) & (!g2225)) + ((!g827) & (g1009) & (!g1043) & (g2224) & (g2271) & (g2225)) + ((!g827) & (g1009) & (g1043) & (!g2224) & (g2271) & (!g2225)) + ((!g827) & (g1009) & (g1043) & (!g2224) & (g2271) & (g2225)) + ((!g827) & (g1009) & (g1043) & (g2224) & (g2271) & (!g2225)) + ((!g827) & (g1009) & (g1043) & (g2224) & (g2271) & (g2225)) + ((g827) & (!g1009) & (!g1043) & (!g2224) & (g2271) & (!g2225)) + ((g827) & (!g1009) & (!g1043) & (!g2224) & (g2271) & (g2225)) + ((g827) & (!g1009) & (!g1043) & (g2224) & (!g2271) & (g2225)) + ((g827) & (!g1009) & (!g1043) & (g2224) & (g2271) & (!g2225)) + ((g827) & (!g1009) & (g1043) & (!g2224) & (!g2271) & (!g2225)) + ((g827) & (!g1009) & (g1043) & (!g2224) & (!g2271) & (g2225)) + ((g827) & (!g1009) & (g1043) & (g2224) & (!g2271) & (!g2225)) + ((g827) & (!g1009) & (g1043) & (g2224) & (g2271) & (g2225)) + ((g827) & (g1009) & (!g1043) & (!g2224) & (!g2271) & (g2225)) + ((g827) & (g1009) & (!g1043) & (!g2224) & (g2271) & (!g2225)) + ((g827) & (g1009) & (!g1043) & (g2224) & (!g2271) & (!g2225)) + ((g827) & (g1009) & (!g1043) & (g2224) & (!g2271) & (g2225)) + ((g827) & (g1009) & (g1043) & (!g2224) & (!g2271) & (!g2225)) + ((g827) & (g1009) & (g1043) & (!g2224) & (g2271) & (g2225)) + ((g827) & (g1009) & (g1043) & (g2224) & (g2271) & (!g2225)) + ((g827) & (g1009) & (g1043) & (g2224) & (g2271) & (g2225)));
	assign g7959 = (((!g3464) & (g6702) & (!g2273)) + ((!g3464) & (g6702) & (g2273)) + ((g3464) & (!g6702) & (g2273)) + ((g3464) & (g6702) & (g2273)));
	assign g2274 = (((!g827) & (!g1017) & (!g1045) & (!g2236) & (g2273) & (!g2237)) + ((!g827) & (!g1017) & (!g1045) & (!g2236) & (g2273) & (g2237)) + ((!g827) & (!g1017) & (!g1045) & (g2236) & (g2273) & (!g2237)) + ((!g827) & (!g1017) & (!g1045) & (g2236) & (g2273) & (g2237)) + ((!g827) & (!g1017) & (g1045) & (!g2236) & (g2273) & (!g2237)) + ((!g827) & (!g1017) & (g1045) & (!g2236) & (g2273) & (g2237)) + ((!g827) & (!g1017) & (g1045) & (g2236) & (g2273) & (!g2237)) + ((!g827) & (!g1017) & (g1045) & (g2236) & (g2273) & (g2237)) + ((!g827) & (g1017) & (!g1045) & (!g2236) & (g2273) & (!g2237)) + ((!g827) & (g1017) & (!g1045) & (!g2236) & (g2273) & (g2237)) + ((!g827) & (g1017) & (!g1045) & (g2236) & (g2273) & (!g2237)) + ((!g827) & (g1017) & (!g1045) & (g2236) & (g2273) & (g2237)) + ((!g827) & (g1017) & (g1045) & (!g2236) & (g2273) & (!g2237)) + ((!g827) & (g1017) & (g1045) & (!g2236) & (g2273) & (g2237)) + ((!g827) & (g1017) & (g1045) & (g2236) & (g2273) & (!g2237)) + ((!g827) & (g1017) & (g1045) & (g2236) & (g2273) & (g2237)) + ((g827) & (!g1017) & (!g1045) & (!g2236) & (g2273) & (!g2237)) + ((g827) & (!g1017) & (!g1045) & (!g2236) & (g2273) & (g2237)) + ((g827) & (!g1017) & (!g1045) & (g2236) & (!g2273) & (g2237)) + ((g827) & (!g1017) & (!g1045) & (g2236) & (g2273) & (!g2237)) + ((g827) & (!g1017) & (g1045) & (!g2236) & (!g2273) & (!g2237)) + ((g827) & (!g1017) & (g1045) & (!g2236) & (!g2273) & (g2237)) + ((g827) & (!g1017) & (g1045) & (g2236) & (!g2273) & (!g2237)) + ((g827) & (!g1017) & (g1045) & (g2236) & (g2273) & (g2237)) + ((g827) & (g1017) & (!g1045) & (!g2236) & (!g2273) & (g2237)) + ((g827) & (g1017) & (!g1045) & (!g2236) & (g2273) & (!g2237)) + ((g827) & (g1017) & (!g1045) & (g2236) & (!g2273) & (!g2237)) + ((g827) & (g1017) & (!g1045) & (g2236) & (!g2273) & (g2237)) + ((g827) & (g1017) & (g1045) & (!g2236) & (!g2273) & (!g2237)) + ((g827) & (g1017) & (g1045) & (!g2236) & (g2273) & (g2237)) + ((g827) & (g1017) & (g1045) & (g2236) & (g2273) & (!g2237)) + ((g827) & (g1017) & (g1045) & (g2236) & (g2273) & (g2237)));
	assign g7960 = (((!g3499) & (g6691) & (!g2275)) + ((!g3499) & (g6691) & (g2275)) + ((g3499) & (!g6691) & (g2275)) + ((g3499) & (g6691) & (g2275)));
	assign g2276 = (((!g827) & (!g1025) & (!g1047) & (!g2247) & (g2275) & (!g2248)) + ((!g827) & (!g1025) & (!g1047) & (!g2247) & (g2275) & (g2248)) + ((!g827) & (!g1025) & (!g1047) & (g2247) & (g2275) & (!g2248)) + ((!g827) & (!g1025) & (!g1047) & (g2247) & (g2275) & (g2248)) + ((!g827) & (!g1025) & (g1047) & (!g2247) & (g2275) & (!g2248)) + ((!g827) & (!g1025) & (g1047) & (!g2247) & (g2275) & (g2248)) + ((!g827) & (!g1025) & (g1047) & (g2247) & (g2275) & (!g2248)) + ((!g827) & (!g1025) & (g1047) & (g2247) & (g2275) & (g2248)) + ((!g827) & (g1025) & (!g1047) & (!g2247) & (g2275) & (!g2248)) + ((!g827) & (g1025) & (!g1047) & (!g2247) & (g2275) & (g2248)) + ((!g827) & (g1025) & (!g1047) & (g2247) & (g2275) & (!g2248)) + ((!g827) & (g1025) & (!g1047) & (g2247) & (g2275) & (g2248)) + ((!g827) & (g1025) & (g1047) & (!g2247) & (g2275) & (!g2248)) + ((!g827) & (g1025) & (g1047) & (!g2247) & (g2275) & (g2248)) + ((!g827) & (g1025) & (g1047) & (g2247) & (g2275) & (!g2248)) + ((!g827) & (g1025) & (g1047) & (g2247) & (g2275) & (g2248)) + ((g827) & (!g1025) & (!g1047) & (!g2247) & (g2275) & (!g2248)) + ((g827) & (!g1025) & (!g1047) & (!g2247) & (g2275) & (g2248)) + ((g827) & (!g1025) & (!g1047) & (g2247) & (!g2275) & (g2248)) + ((g827) & (!g1025) & (!g1047) & (g2247) & (g2275) & (!g2248)) + ((g827) & (!g1025) & (g1047) & (!g2247) & (!g2275) & (!g2248)) + ((g827) & (!g1025) & (g1047) & (!g2247) & (!g2275) & (g2248)) + ((g827) & (!g1025) & (g1047) & (g2247) & (!g2275) & (!g2248)) + ((g827) & (!g1025) & (g1047) & (g2247) & (g2275) & (g2248)) + ((g827) & (g1025) & (!g1047) & (!g2247) & (!g2275) & (g2248)) + ((g827) & (g1025) & (!g1047) & (!g2247) & (g2275) & (!g2248)) + ((g827) & (g1025) & (!g1047) & (g2247) & (!g2275) & (!g2248)) + ((g827) & (g1025) & (!g1047) & (g2247) & (!g2275) & (g2248)) + ((g827) & (g1025) & (g1047) & (!g2247) & (!g2275) & (!g2248)) + ((g827) & (g1025) & (g1047) & (!g2247) & (g2275) & (g2248)) + ((g827) & (g1025) & (g1047) & (g2247) & (g2275) & (!g2248)) + ((g827) & (g1025) & (g1047) & (g2247) & (g2275) & (g2248)));
	assign g7961 = (((!g3464) & (g6680) & (!g2277)) + ((!g3464) & (g6680) & (g2277)) + ((g3464) & (!g6680) & (g2277)) + ((g3464) & (g6680) & (g2277)));
	assign g2278 = (((!g827) & (!g1003) & (!g1049) & (!g2217) & (g2277) & (!g2218)) + ((!g827) & (!g1003) & (!g1049) & (!g2217) & (g2277) & (g2218)) + ((!g827) & (!g1003) & (!g1049) & (g2217) & (g2277) & (!g2218)) + ((!g827) & (!g1003) & (!g1049) & (g2217) & (g2277) & (g2218)) + ((!g827) & (!g1003) & (g1049) & (!g2217) & (g2277) & (!g2218)) + ((!g827) & (!g1003) & (g1049) & (!g2217) & (g2277) & (g2218)) + ((!g827) & (!g1003) & (g1049) & (g2217) & (g2277) & (!g2218)) + ((!g827) & (!g1003) & (g1049) & (g2217) & (g2277) & (g2218)) + ((!g827) & (g1003) & (!g1049) & (!g2217) & (g2277) & (!g2218)) + ((!g827) & (g1003) & (!g1049) & (!g2217) & (g2277) & (g2218)) + ((!g827) & (g1003) & (!g1049) & (g2217) & (g2277) & (!g2218)) + ((!g827) & (g1003) & (!g1049) & (g2217) & (g2277) & (g2218)) + ((!g827) & (g1003) & (g1049) & (!g2217) & (g2277) & (!g2218)) + ((!g827) & (g1003) & (g1049) & (!g2217) & (g2277) & (g2218)) + ((!g827) & (g1003) & (g1049) & (g2217) & (g2277) & (!g2218)) + ((!g827) & (g1003) & (g1049) & (g2217) & (g2277) & (g2218)) + ((g827) & (!g1003) & (!g1049) & (!g2217) & (g2277) & (!g2218)) + ((g827) & (!g1003) & (!g1049) & (!g2217) & (g2277) & (g2218)) + ((g827) & (!g1003) & (!g1049) & (g2217) & (!g2277) & (g2218)) + ((g827) & (!g1003) & (!g1049) & (g2217) & (g2277) & (!g2218)) + ((g827) & (!g1003) & (g1049) & (!g2217) & (!g2277) & (!g2218)) + ((g827) & (!g1003) & (g1049) & (!g2217) & (!g2277) & (g2218)) + ((g827) & (!g1003) & (g1049) & (g2217) & (!g2277) & (!g2218)) + ((g827) & (!g1003) & (g1049) & (g2217) & (g2277) & (g2218)) + ((g827) & (g1003) & (!g1049) & (!g2217) & (!g2277) & (g2218)) + ((g827) & (g1003) & (!g1049) & (!g2217) & (g2277) & (!g2218)) + ((g827) & (g1003) & (!g1049) & (g2217) & (!g2277) & (!g2218)) + ((g827) & (g1003) & (!g1049) & (g2217) & (!g2277) & (g2218)) + ((g827) & (g1003) & (g1049) & (!g2217) & (!g2277) & (!g2218)) + ((g827) & (g1003) & (g1049) & (!g2217) & (g2277) & (g2218)) + ((g827) & (g1003) & (g1049) & (g2217) & (g2277) & (!g2218)) + ((g827) & (g1003) & (g1049) & (g2217) & (g2277) & (g2218)));
	assign g7962 = (((!g3499) & (g6669) & (!g2279)) + ((!g3499) & (g6669) & (g2279)) + ((g3499) & (!g6669) & (g2279)) + ((g3499) & (g6669) & (g2279)));
	assign g2280 = (((!g827) & (!g1011) & (!g1051) & (!g2227) & (g2279) & (!g2228)) + ((!g827) & (!g1011) & (!g1051) & (!g2227) & (g2279) & (g2228)) + ((!g827) & (!g1011) & (!g1051) & (g2227) & (g2279) & (!g2228)) + ((!g827) & (!g1011) & (!g1051) & (g2227) & (g2279) & (g2228)) + ((!g827) & (!g1011) & (g1051) & (!g2227) & (g2279) & (!g2228)) + ((!g827) & (!g1011) & (g1051) & (!g2227) & (g2279) & (g2228)) + ((!g827) & (!g1011) & (g1051) & (g2227) & (g2279) & (!g2228)) + ((!g827) & (!g1011) & (g1051) & (g2227) & (g2279) & (g2228)) + ((!g827) & (g1011) & (!g1051) & (!g2227) & (g2279) & (!g2228)) + ((!g827) & (g1011) & (!g1051) & (!g2227) & (g2279) & (g2228)) + ((!g827) & (g1011) & (!g1051) & (g2227) & (g2279) & (!g2228)) + ((!g827) & (g1011) & (!g1051) & (g2227) & (g2279) & (g2228)) + ((!g827) & (g1011) & (g1051) & (!g2227) & (g2279) & (!g2228)) + ((!g827) & (g1011) & (g1051) & (!g2227) & (g2279) & (g2228)) + ((!g827) & (g1011) & (g1051) & (g2227) & (g2279) & (!g2228)) + ((!g827) & (g1011) & (g1051) & (g2227) & (g2279) & (g2228)) + ((g827) & (!g1011) & (!g1051) & (!g2227) & (g2279) & (!g2228)) + ((g827) & (!g1011) & (!g1051) & (!g2227) & (g2279) & (g2228)) + ((g827) & (!g1011) & (!g1051) & (g2227) & (!g2279) & (g2228)) + ((g827) & (!g1011) & (!g1051) & (g2227) & (g2279) & (!g2228)) + ((g827) & (!g1011) & (g1051) & (!g2227) & (!g2279) & (!g2228)) + ((g827) & (!g1011) & (g1051) & (!g2227) & (!g2279) & (g2228)) + ((g827) & (!g1011) & (g1051) & (g2227) & (!g2279) & (!g2228)) + ((g827) & (!g1011) & (g1051) & (g2227) & (g2279) & (g2228)) + ((g827) & (g1011) & (!g1051) & (!g2227) & (!g2279) & (g2228)) + ((g827) & (g1011) & (!g1051) & (!g2227) & (g2279) & (!g2228)) + ((g827) & (g1011) & (!g1051) & (g2227) & (!g2279) & (!g2228)) + ((g827) & (g1011) & (!g1051) & (g2227) & (!g2279) & (g2228)) + ((g827) & (g1011) & (g1051) & (!g2227) & (!g2279) & (!g2228)) + ((g827) & (g1011) & (g1051) & (!g2227) & (g2279) & (g2228)) + ((g827) & (g1011) & (g1051) & (g2227) & (g2279) & (!g2228)) + ((g827) & (g1011) & (g1051) & (g2227) & (g2279) & (g2228)));
	assign g7963 = (((!g2017) & (g4519) & (!g2281)) + ((!g2017) & (g4519) & (g2281)) + ((g2017) & (!g4519) & (g2281)) + ((g2017) & (g4519) & (g2281)));
	assign g2282 = (((!g827) & (!g1019) & (!g1053) & (!g2239) & (g2281) & (!g2240)) + ((!g827) & (!g1019) & (!g1053) & (!g2239) & (g2281) & (g2240)) + ((!g827) & (!g1019) & (!g1053) & (g2239) & (g2281) & (!g2240)) + ((!g827) & (!g1019) & (!g1053) & (g2239) & (g2281) & (g2240)) + ((!g827) & (!g1019) & (g1053) & (!g2239) & (g2281) & (!g2240)) + ((!g827) & (!g1019) & (g1053) & (!g2239) & (g2281) & (g2240)) + ((!g827) & (!g1019) & (g1053) & (g2239) & (g2281) & (!g2240)) + ((!g827) & (!g1019) & (g1053) & (g2239) & (g2281) & (g2240)) + ((!g827) & (g1019) & (!g1053) & (!g2239) & (g2281) & (!g2240)) + ((!g827) & (g1019) & (!g1053) & (!g2239) & (g2281) & (g2240)) + ((!g827) & (g1019) & (!g1053) & (g2239) & (g2281) & (!g2240)) + ((!g827) & (g1019) & (!g1053) & (g2239) & (g2281) & (g2240)) + ((!g827) & (g1019) & (g1053) & (!g2239) & (g2281) & (!g2240)) + ((!g827) & (g1019) & (g1053) & (!g2239) & (g2281) & (g2240)) + ((!g827) & (g1019) & (g1053) & (g2239) & (g2281) & (!g2240)) + ((!g827) & (g1019) & (g1053) & (g2239) & (g2281) & (g2240)) + ((g827) & (!g1019) & (!g1053) & (!g2239) & (g2281) & (!g2240)) + ((g827) & (!g1019) & (!g1053) & (!g2239) & (g2281) & (g2240)) + ((g827) & (!g1019) & (!g1053) & (g2239) & (!g2281) & (g2240)) + ((g827) & (!g1019) & (!g1053) & (g2239) & (g2281) & (!g2240)) + ((g827) & (!g1019) & (g1053) & (!g2239) & (!g2281) & (!g2240)) + ((g827) & (!g1019) & (g1053) & (!g2239) & (!g2281) & (g2240)) + ((g827) & (!g1019) & (g1053) & (g2239) & (!g2281) & (!g2240)) + ((g827) & (!g1019) & (g1053) & (g2239) & (g2281) & (g2240)) + ((g827) & (g1019) & (!g1053) & (!g2239) & (!g2281) & (g2240)) + ((g827) & (g1019) & (!g1053) & (!g2239) & (g2281) & (!g2240)) + ((g827) & (g1019) & (!g1053) & (g2239) & (!g2281) & (!g2240)) + ((g827) & (g1019) & (!g1053) & (g2239) & (!g2281) & (g2240)) + ((g827) & (g1019) & (g1053) & (!g2239) & (!g2281) & (!g2240)) + ((g827) & (g1019) & (g1053) & (!g2239) & (g2281) & (g2240)) + ((g827) & (g1019) & (g1053) & (g2239) & (g2281) & (!g2240)) + ((g827) & (g1019) & (g1053) & (g2239) & (g2281) & (g2240)));
	assign g7964 = (((!g3429) & (g4522) & (!g2283)) + ((!g3429) & (g4522) & (g2283)) + ((g3429) & (!g4522) & (g2283)) + ((g3429) & (g4522) & (g2283)));
	assign g2284 = (((!g827) & (!g1027) & (!g1055) & (!g2250) & (g2283) & (!g2251)) + ((!g827) & (!g1027) & (!g1055) & (!g2250) & (g2283) & (g2251)) + ((!g827) & (!g1027) & (!g1055) & (g2250) & (g2283) & (!g2251)) + ((!g827) & (!g1027) & (!g1055) & (g2250) & (g2283) & (g2251)) + ((!g827) & (!g1027) & (g1055) & (!g2250) & (g2283) & (!g2251)) + ((!g827) & (!g1027) & (g1055) & (!g2250) & (g2283) & (g2251)) + ((!g827) & (!g1027) & (g1055) & (g2250) & (g2283) & (!g2251)) + ((!g827) & (!g1027) & (g1055) & (g2250) & (g2283) & (g2251)) + ((!g827) & (g1027) & (!g1055) & (!g2250) & (g2283) & (!g2251)) + ((!g827) & (g1027) & (!g1055) & (!g2250) & (g2283) & (g2251)) + ((!g827) & (g1027) & (!g1055) & (g2250) & (g2283) & (!g2251)) + ((!g827) & (g1027) & (!g1055) & (g2250) & (g2283) & (g2251)) + ((!g827) & (g1027) & (g1055) & (!g2250) & (g2283) & (!g2251)) + ((!g827) & (g1027) & (g1055) & (!g2250) & (g2283) & (g2251)) + ((!g827) & (g1027) & (g1055) & (g2250) & (g2283) & (!g2251)) + ((!g827) & (g1027) & (g1055) & (g2250) & (g2283) & (g2251)) + ((g827) & (!g1027) & (!g1055) & (!g2250) & (g2283) & (!g2251)) + ((g827) & (!g1027) & (!g1055) & (!g2250) & (g2283) & (g2251)) + ((g827) & (!g1027) & (!g1055) & (g2250) & (!g2283) & (g2251)) + ((g827) & (!g1027) & (!g1055) & (g2250) & (g2283) & (!g2251)) + ((g827) & (!g1027) & (g1055) & (!g2250) & (!g2283) & (!g2251)) + ((g827) & (!g1027) & (g1055) & (!g2250) & (!g2283) & (g2251)) + ((g827) & (!g1027) & (g1055) & (g2250) & (!g2283) & (!g2251)) + ((g827) & (!g1027) & (g1055) & (g2250) & (g2283) & (g2251)) + ((g827) & (g1027) & (!g1055) & (!g2250) & (!g2283) & (g2251)) + ((g827) & (g1027) & (!g1055) & (!g2250) & (g2283) & (!g2251)) + ((g827) & (g1027) & (!g1055) & (g2250) & (!g2283) & (!g2251)) + ((g827) & (g1027) & (!g1055) & (g2250) & (!g2283) & (g2251)) + ((g827) & (g1027) & (g1055) & (!g2250) & (!g2283) & (!g2251)) + ((g827) & (g1027) & (g1055) & (!g2250) & (g2283) & (g2251)) + ((g827) & (g1027) & (g1055) & (g2250) & (g2283) & (!g2251)) + ((g827) & (g1027) & (g1055) & (g2250) & (g2283) & (g2251)));
	assign g2285 = (((!g827) & (!g1005) & (!g1057) & (!g1992) & (g1994) & (!g2220)) + ((!g827) & (!g1005) & (!g1057) & (!g1992) & (g1994) & (g2220)) + ((!g827) & (!g1005) & (!g1057) & (g1992) & (g1994) & (!g2220)) + ((!g827) & (!g1005) & (!g1057) & (g1992) & (g1994) & (g2220)) + ((!g827) & (!g1005) & (g1057) & (!g1992) & (g1994) & (!g2220)) + ((!g827) & (!g1005) & (g1057) & (!g1992) & (g1994) & (g2220)) + ((!g827) & (!g1005) & (g1057) & (g1992) & (g1994) & (!g2220)) + ((!g827) & (!g1005) & (g1057) & (g1992) & (g1994) & (g2220)) + ((!g827) & (g1005) & (!g1057) & (!g1992) & (g1994) & (!g2220)) + ((!g827) & (g1005) & (!g1057) & (!g1992) & (g1994) & (g2220)) + ((!g827) & (g1005) & (!g1057) & (g1992) & (g1994) & (!g2220)) + ((!g827) & (g1005) & (!g1057) & (g1992) & (g1994) & (g2220)) + ((!g827) & (g1005) & (g1057) & (!g1992) & (g1994) & (!g2220)) + ((!g827) & (g1005) & (g1057) & (!g1992) & (g1994) & (g2220)) + ((!g827) & (g1005) & (g1057) & (g1992) & (g1994) & (!g2220)) + ((!g827) & (g1005) & (g1057) & (g1992) & (g1994) & (g2220)) + ((g827) & (!g1005) & (!g1057) & (!g1992) & (g1994) & (!g2220)) + ((g827) & (!g1005) & (!g1057) & (!g1992) & (g1994) & (g2220)) + ((g827) & (!g1005) & (!g1057) & (g1992) & (!g1994) & (g2220)) + ((g827) & (!g1005) & (!g1057) & (g1992) & (g1994) & (!g2220)) + ((g827) & (!g1005) & (g1057) & (!g1992) & (!g1994) & (!g2220)) + ((g827) & (!g1005) & (g1057) & (!g1992) & (!g1994) & (g2220)) + ((g827) & (!g1005) & (g1057) & (g1992) & (!g1994) & (!g2220)) + ((g827) & (!g1005) & (g1057) & (g1992) & (g1994) & (g2220)) + ((g827) & (g1005) & (!g1057) & (!g1992) & (!g1994) & (g2220)) + ((g827) & (g1005) & (!g1057) & (!g1992) & (g1994) & (!g2220)) + ((g827) & (g1005) & (!g1057) & (g1992) & (!g1994) & (!g2220)) + ((g827) & (g1005) & (!g1057) & (g1992) & (!g1994) & (g2220)) + ((g827) & (g1005) & (g1057) & (!g1992) & (!g1994) & (!g2220)) + ((g827) & (g1005) & (g1057) & (!g1992) & (g1994) & (g2220)) + ((g827) & (g1005) & (g1057) & (g1992) & (g1994) & (!g2220)) + ((g827) & (g1005) & (g1057) & (g1992) & (g1994) & (g2220)));
	assign g7965 = (((!g3464) & (g6658) & (!g2286)) + ((!g3464) & (g6658) & (g2286)) + ((g3464) & (!g6658) & (g2286)) + ((g3464) & (g6658) & (g2286)));
	assign g2287 = (((!g827) & (!g1013) & (!g1059) & (!g2230) & (g2286) & (!g2231)) + ((!g827) & (!g1013) & (!g1059) & (!g2230) & (g2286) & (g2231)) + ((!g827) & (!g1013) & (!g1059) & (g2230) & (g2286) & (!g2231)) + ((!g827) & (!g1013) & (!g1059) & (g2230) & (g2286) & (g2231)) + ((!g827) & (!g1013) & (g1059) & (!g2230) & (g2286) & (!g2231)) + ((!g827) & (!g1013) & (g1059) & (!g2230) & (g2286) & (g2231)) + ((!g827) & (!g1013) & (g1059) & (g2230) & (g2286) & (!g2231)) + ((!g827) & (!g1013) & (g1059) & (g2230) & (g2286) & (g2231)) + ((!g827) & (g1013) & (!g1059) & (!g2230) & (g2286) & (!g2231)) + ((!g827) & (g1013) & (!g1059) & (!g2230) & (g2286) & (g2231)) + ((!g827) & (g1013) & (!g1059) & (g2230) & (g2286) & (!g2231)) + ((!g827) & (g1013) & (!g1059) & (g2230) & (g2286) & (g2231)) + ((!g827) & (g1013) & (g1059) & (!g2230) & (g2286) & (!g2231)) + ((!g827) & (g1013) & (g1059) & (!g2230) & (g2286) & (g2231)) + ((!g827) & (g1013) & (g1059) & (g2230) & (g2286) & (!g2231)) + ((!g827) & (g1013) & (g1059) & (g2230) & (g2286) & (g2231)) + ((g827) & (!g1013) & (!g1059) & (!g2230) & (g2286) & (!g2231)) + ((g827) & (!g1013) & (!g1059) & (!g2230) & (g2286) & (g2231)) + ((g827) & (!g1013) & (!g1059) & (g2230) & (!g2286) & (g2231)) + ((g827) & (!g1013) & (!g1059) & (g2230) & (g2286) & (!g2231)) + ((g827) & (!g1013) & (g1059) & (!g2230) & (!g2286) & (!g2231)) + ((g827) & (!g1013) & (g1059) & (!g2230) & (!g2286) & (g2231)) + ((g827) & (!g1013) & (g1059) & (g2230) & (!g2286) & (!g2231)) + ((g827) & (!g1013) & (g1059) & (g2230) & (g2286) & (g2231)) + ((g827) & (g1013) & (!g1059) & (!g2230) & (!g2286) & (g2231)) + ((g827) & (g1013) & (!g1059) & (!g2230) & (g2286) & (!g2231)) + ((g827) & (g1013) & (!g1059) & (g2230) & (!g2286) & (!g2231)) + ((g827) & (g1013) & (!g1059) & (g2230) & (!g2286) & (g2231)) + ((g827) & (g1013) & (g1059) & (!g2230) & (!g2286) & (!g2231)) + ((g827) & (g1013) & (g1059) & (!g2230) & (g2286) & (g2231)) + ((g827) & (g1013) & (g1059) & (g2230) & (g2286) & (!g2231)) + ((g827) & (g1013) & (g1059) & (g2230) & (g2286) & (g2231)));
	assign g7966 = (((!g3429) & (g4529) & (!g2288)) + ((!g3429) & (g4529) & (g2288)) + ((g3429) & (!g4529) & (g2288)) + ((g3429) & (g4529) & (g2288)));
	assign g2289 = (((!g827) & (!g1021) & (!g1061) & (!g2242) & (g2288) & (!g2243)) + ((!g827) & (!g1021) & (!g1061) & (!g2242) & (g2288) & (g2243)) + ((!g827) & (!g1021) & (!g1061) & (g2242) & (g2288) & (!g2243)) + ((!g827) & (!g1021) & (!g1061) & (g2242) & (g2288) & (g2243)) + ((!g827) & (!g1021) & (g1061) & (!g2242) & (g2288) & (!g2243)) + ((!g827) & (!g1021) & (g1061) & (!g2242) & (g2288) & (g2243)) + ((!g827) & (!g1021) & (g1061) & (g2242) & (g2288) & (!g2243)) + ((!g827) & (!g1021) & (g1061) & (g2242) & (g2288) & (g2243)) + ((!g827) & (g1021) & (!g1061) & (!g2242) & (g2288) & (!g2243)) + ((!g827) & (g1021) & (!g1061) & (!g2242) & (g2288) & (g2243)) + ((!g827) & (g1021) & (!g1061) & (g2242) & (g2288) & (!g2243)) + ((!g827) & (g1021) & (!g1061) & (g2242) & (g2288) & (g2243)) + ((!g827) & (g1021) & (g1061) & (!g2242) & (g2288) & (!g2243)) + ((!g827) & (g1021) & (g1061) & (!g2242) & (g2288) & (g2243)) + ((!g827) & (g1021) & (g1061) & (g2242) & (g2288) & (!g2243)) + ((!g827) & (g1021) & (g1061) & (g2242) & (g2288) & (g2243)) + ((g827) & (!g1021) & (!g1061) & (!g2242) & (g2288) & (!g2243)) + ((g827) & (!g1021) & (!g1061) & (!g2242) & (g2288) & (g2243)) + ((g827) & (!g1021) & (!g1061) & (g2242) & (!g2288) & (g2243)) + ((g827) & (!g1021) & (!g1061) & (g2242) & (g2288) & (!g2243)) + ((g827) & (!g1021) & (g1061) & (!g2242) & (!g2288) & (!g2243)) + ((g827) & (!g1021) & (g1061) & (!g2242) & (!g2288) & (g2243)) + ((g827) & (!g1021) & (g1061) & (g2242) & (!g2288) & (!g2243)) + ((g827) & (!g1021) & (g1061) & (g2242) & (g2288) & (g2243)) + ((g827) & (g1021) & (!g1061) & (!g2242) & (!g2288) & (g2243)) + ((g827) & (g1021) & (!g1061) & (!g2242) & (g2288) & (!g2243)) + ((g827) & (g1021) & (!g1061) & (g2242) & (!g2288) & (!g2243)) + ((g827) & (g1021) & (!g1061) & (g2242) & (!g2288) & (g2243)) + ((g827) & (g1021) & (g1061) & (!g2242) & (!g2288) & (!g2243)) + ((g827) & (g1021) & (g1061) & (!g2242) & (g2288) & (g2243)) + ((g827) & (g1021) & (g1061) & (g2242) & (g2288) & (!g2243)) + ((g827) & (g1021) & (g1061) & (g2242) & (g2288) & (g2243)));
	assign g7967 = (((!g2017) & (g4535) & (!g2290)) + ((!g2017) & (g4535) & (g2290)) + ((g2017) & (!g4535) & (g2290)) + ((g2017) & (g4535) & (g2290)));
	assign g2291 = (((!g827) & (!g1029) & (!g1063) & (!g2253) & (g2290) & (!g2254)) + ((!g827) & (!g1029) & (!g1063) & (!g2253) & (g2290) & (g2254)) + ((!g827) & (!g1029) & (!g1063) & (g2253) & (g2290) & (!g2254)) + ((!g827) & (!g1029) & (!g1063) & (g2253) & (g2290) & (g2254)) + ((!g827) & (!g1029) & (g1063) & (!g2253) & (g2290) & (!g2254)) + ((!g827) & (!g1029) & (g1063) & (!g2253) & (g2290) & (g2254)) + ((!g827) & (!g1029) & (g1063) & (g2253) & (g2290) & (!g2254)) + ((!g827) & (!g1029) & (g1063) & (g2253) & (g2290) & (g2254)) + ((!g827) & (g1029) & (!g1063) & (!g2253) & (g2290) & (!g2254)) + ((!g827) & (g1029) & (!g1063) & (!g2253) & (g2290) & (g2254)) + ((!g827) & (g1029) & (!g1063) & (g2253) & (g2290) & (!g2254)) + ((!g827) & (g1029) & (!g1063) & (g2253) & (g2290) & (g2254)) + ((!g827) & (g1029) & (g1063) & (!g2253) & (g2290) & (!g2254)) + ((!g827) & (g1029) & (g1063) & (!g2253) & (g2290) & (g2254)) + ((!g827) & (g1029) & (g1063) & (g2253) & (g2290) & (!g2254)) + ((!g827) & (g1029) & (g1063) & (g2253) & (g2290) & (g2254)) + ((g827) & (!g1029) & (!g1063) & (!g2253) & (g2290) & (!g2254)) + ((g827) & (!g1029) & (!g1063) & (!g2253) & (g2290) & (g2254)) + ((g827) & (!g1029) & (!g1063) & (g2253) & (!g2290) & (g2254)) + ((g827) & (!g1029) & (!g1063) & (g2253) & (g2290) & (!g2254)) + ((g827) & (!g1029) & (g1063) & (!g2253) & (!g2290) & (!g2254)) + ((g827) & (!g1029) & (g1063) & (!g2253) & (!g2290) & (g2254)) + ((g827) & (!g1029) & (g1063) & (g2253) & (!g2290) & (!g2254)) + ((g827) & (!g1029) & (g1063) & (g2253) & (g2290) & (g2254)) + ((g827) & (g1029) & (!g1063) & (!g2253) & (!g2290) & (g2254)) + ((g827) & (g1029) & (!g1063) & (!g2253) & (g2290) & (!g2254)) + ((g827) & (g1029) & (!g1063) & (g2253) & (!g2290) & (!g2254)) + ((g827) & (g1029) & (!g1063) & (g2253) & (!g2290) & (g2254)) + ((g827) & (g1029) & (g1063) & (!g2253) & (!g2290) & (!g2254)) + ((g827) & (g1029) & (g1063) & (!g2253) & (g2290) & (g2254)) + ((g827) & (g1029) & (g1063) & (g2253) & (g2290) & (!g2254)) + ((g827) & (g1029) & (g1063) & (g2253) & (g2290) & (g2254)));
	assign g2292 = (((!g2256) & (g2257)) + ((g2256) & (!g2257)));
	assign g2293 = (((!g2176) & (!g2177) & (!g2178) & (g2210) & (g2211) & (g2292)) + ((!g2176) & (!g2177) & (g2178) & (g2210) & (g2211) & (g2292)) + ((!g2176) & (g2177) & (!g2178) & (g2210) & (g2211) & (g2292)) + ((!g2176) & (g2177) & (g2178) & (!g2210) & (g2211) & (g2292)) + ((!g2176) & (g2177) & (g2178) & (g2210) & (!g2211) & (g2292)) + ((!g2176) & (g2177) & (g2178) & (g2210) & (g2211) & (g2292)) + ((g2176) & (!g2177) & (!g2178) & (g2210) & (g2211) & (g2292)) + ((g2176) & (!g2177) & (g2178) & (!g2210) & (g2211) & (g2292)) + ((g2176) & (!g2177) & (g2178) & (g2210) & (!g2211) & (g2292)) + ((g2176) & (!g2177) & (g2178) & (g2210) & (g2211) & (g2292)) + ((g2176) & (g2177) & (!g2178) & (!g2210) & (g2211) & (g2292)) + ((g2176) & (g2177) & (!g2178) & (g2210) & (!g2211) & (g2292)) + ((g2176) & (g2177) & (!g2178) & (g2210) & (g2211) & (g2292)) + ((g2176) & (g2177) & (g2178) & (!g2210) & (g2211) & (g2292)) + ((g2176) & (g2177) & (g2178) & (g2210) & (!g2211) & (g2292)) + ((g2176) & (g2177) & (g2178) & (g2210) & (g2211) & (g2292)));
	assign g2294 = (((g2256) & (g2257)));
	assign g7968 = (((!g3429) & (g4538) & (!g2295)) + ((!g3429) & (g4538) & (g2295)) + ((g3429) & (!g4538) & (g2295)) + ((g3429) & (g4538) & (g2295)));
	assign g7969 = (((!g3464) & (g4542) & (!g2296)) + ((!g3464) & (g4542) & (g2296)) + ((g3464) & (!g4542) & (g2296)) + ((g3464) & (g4542) & (g2296)));
	assign g2297 = (((!g2293) & (!g2294) & (!g2295) & (g2296)) + ((!g2293) & (!g2294) & (g2295) & (!g2296)) + ((!g2293) & (g2294) & (!g2295) & (!g2296)) + ((!g2293) & (g2294) & (g2295) & (g2296)) + ((g2293) & (!g2294) & (!g2295) & (!g2296)) + ((g2293) & (!g2294) & (g2295) & (g2296)) + ((g2293) & (g2294) & (!g2295) & (!g2296)) + ((g2293) & (g2294) & (g2295) & (g2296)));
	assign g7970 = (((!g3429) & (g4546) & (!g2298)) + ((!g3429) & (g4546) & (g2298)) + ((g3429) & (!g4546) & (g2298)) + ((g3429) & (g4546) & (g2298)));
	assign g7971 = (((!g3499) & (g4550) & (!g2299)) + ((!g3499) & (g4550) & (g2299)) + ((g3499) & (!g4550) & (g2299)) + ((g3499) & (g4550) & (g2299)));
	assign g2300 = (((!g2260) & (!g2261) & (!g2262) & (!g2263) & (!g2298) & (g2299)) + ((!g2260) & (!g2261) & (!g2262) & (!g2263) & (g2298) & (!g2299)) + ((!g2260) & (!g2261) & (!g2262) & (g2263) & (!g2298) & (g2299)) + ((!g2260) & (!g2261) & (!g2262) & (g2263) & (g2298) & (!g2299)) + ((!g2260) & (!g2261) & (g2262) & (!g2263) & (!g2298) & (g2299)) + ((!g2260) & (!g2261) & (g2262) & (!g2263) & (g2298) & (!g2299)) + ((!g2260) & (!g2261) & (g2262) & (g2263) & (!g2298) & (!g2299)) + ((!g2260) & (!g2261) & (g2262) & (g2263) & (g2298) & (g2299)) + ((!g2260) & (g2261) & (!g2262) & (!g2263) & (!g2298) & (g2299)) + ((!g2260) & (g2261) & (!g2262) & (!g2263) & (g2298) & (!g2299)) + ((!g2260) & (g2261) & (!g2262) & (g2263) & (!g2298) & (!g2299)) + ((!g2260) & (g2261) & (!g2262) & (g2263) & (g2298) & (g2299)) + ((!g2260) & (g2261) & (g2262) & (!g2263) & (!g2298) & (!g2299)) + ((!g2260) & (g2261) & (g2262) & (!g2263) & (g2298) & (g2299)) + ((!g2260) & (g2261) & (g2262) & (g2263) & (!g2298) & (!g2299)) + ((!g2260) & (g2261) & (g2262) & (g2263) & (g2298) & (g2299)) + ((g2260) & (!g2261) & (!g2262) & (!g2263) & (!g2298) & (g2299)) + ((g2260) & (!g2261) & (!g2262) & (!g2263) & (g2298) & (!g2299)) + ((g2260) & (!g2261) & (!g2262) & (g2263) & (!g2298) & (!g2299)) + ((g2260) & (!g2261) & (!g2262) & (g2263) & (g2298) & (g2299)) + ((g2260) & (!g2261) & (g2262) & (!g2263) & (!g2298) & (!g2299)) + ((g2260) & (!g2261) & (g2262) & (!g2263) & (g2298) & (g2299)) + ((g2260) & (!g2261) & (g2262) & (g2263) & (!g2298) & (!g2299)) + ((g2260) & (!g2261) & (g2262) & (g2263) & (g2298) & (g2299)) + ((g2260) & (g2261) & (!g2262) & (!g2263) & (!g2298) & (g2299)) + ((g2260) & (g2261) & (!g2262) & (!g2263) & (g2298) & (!g2299)) + ((g2260) & (g2261) & (!g2262) & (g2263) & (!g2298) & (!g2299)) + ((g2260) & (g2261) & (!g2262) & (g2263) & (g2298) & (g2299)) + ((g2260) & (g2261) & (g2262) & (!g2263) & (!g2298) & (!g2299)) + ((g2260) & (g2261) & (g2262) & (!g2263) & (g2298) & (g2299)) + ((g2260) & (g2261) & (g2262) & (g2263) & (!g2298) & (!g2299)) + ((g2260) & (g2261) & (g2262) & (g2263) & (g2298) & (g2299)));
	assign g2301 = (((g830) & (!g1914) & (!g2297) & (!g2300) & (g1065)) + ((g830) & (!g1914) & (!g2297) & (g2300) & (!g1065)) + ((g830) & (!g1914) & (g2297) & (!g2300) & (g1065)) + ((g830) & (!g1914) & (g2297) & (g2300) & (!g1065)) + ((g830) & (g1914) & (!g2297) & (!g2300) & (g1065)) + ((g830) & (g1914) & (!g2297) & (g2300) & (g1065)) + ((g830) & (g1914) & (g2297) & (!g2300) & (!g1065)) + ((g830) & (g1914) & (g2297) & (g2300) & (!g1065)));
	assign g2302 = (((!g1001) & (!g1041) & (g1991) & (g1993) & (g2215)) + ((!g1001) & (g1041) & (!g1991) & (g1993) & (!g2215)) + ((!g1001) & (g1041) & (!g1991) & (g1993) & (g2215)) + ((!g1001) & (g1041) & (g1991) & (!g1993) & (g2215)) + ((!g1001) & (g1041) & (g1991) & (g1993) & (!g2215)) + ((!g1001) & (g1041) & (g1991) & (g1993) & (g2215)) + ((g1001) & (!g1041) & (!g1991) & (g1993) & (g2215)) + ((g1001) & (!g1041) & (g1991) & (g1993) & (!g2215)) + ((g1001) & (!g1041) & (g1991) & (g1993) & (g2215)) + ((g1001) & (g1041) & (!g1991) & (!g1993) & (g2215)) + ((g1001) & (g1041) & (!g1991) & (g1993) & (!g2215)) + ((g1001) & (g1041) & (!g1991) & (g1993) & (g2215)) + ((g1001) & (g1041) & (g1991) & (!g1993) & (!g2215)) + ((g1001) & (g1041) & (g1991) & (!g1993) & (g2215)) + ((g1001) & (g1041) & (g1991) & (g1993) & (!g2215)) + ((g1001) & (g1041) & (g1991) & (g1993) & (g2215)));
	assign g2303 = (((!g827) & (!g1068) & (g1996) & (!g2302)) + ((!g827) & (!g1068) & (g1996) & (g2302)) + ((!g827) & (g1068) & (g1996) & (!g2302)) + ((!g827) & (g1068) & (g1996) & (g2302)) + ((g827) & (!g1068) & (!g1996) & (g2302)) + ((g827) & (!g1068) & (g1996) & (!g2302)) + ((g827) & (g1068) & (!g1996) & (!g2302)) + ((g827) & (g1068) & (g1996) & (g2302)));
	assign g7972 = (((!g3464) & (g4554) & (!g2304)) + ((!g3464) & (g4554) & (g2304)) + ((g3464) & (!g4554) & (g2304)) + ((g3464) & (g4554) & (g2304)));
	assign g2305 = (((!g1003) & (!g1049) & (g2217) & (g2277) & (g2218)) + ((!g1003) & (g1049) & (!g2217) & (g2277) & (!g2218)) + ((!g1003) & (g1049) & (!g2217) & (g2277) & (g2218)) + ((!g1003) & (g1049) & (g2217) & (!g2277) & (g2218)) + ((!g1003) & (g1049) & (g2217) & (g2277) & (!g2218)) + ((!g1003) & (g1049) & (g2217) & (g2277) & (g2218)) + ((g1003) & (!g1049) & (!g2217) & (g2277) & (g2218)) + ((g1003) & (!g1049) & (g2217) & (g2277) & (!g2218)) + ((g1003) & (!g1049) & (g2217) & (g2277) & (g2218)) + ((g1003) & (g1049) & (!g2217) & (!g2277) & (g2218)) + ((g1003) & (g1049) & (!g2217) & (g2277) & (!g2218)) + ((g1003) & (g1049) & (!g2217) & (g2277) & (g2218)) + ((g1003) & (g1049) & (g2217) & (!g2277) & (!g2218)) + ((g1003) & (g1049) & (g2217) & (!g2277) & (g2218)) + ((g1003) & (g1049) & (g2217) & (g2277) & (!g2218)) + ((g1003) & (g1049) & (g2217) & (g2277) & (g2218)));
	assign g2306 = (((!g827) & (!g1070) & (g2304) & (!g2305)) + ((!g827) & (!g1070) & (g2304) & (g2305)) + ((!g827) & (g1070) & (g2304) & (!g2305)) + ((!g827) & (g1070) & (g2304) & (g2305)) + ((g827) & (!g1070) & (!g2304) & (g2305)) + ((g827) & (!g1070) & (g2304) & (!g2305)) + ((g827) & (g1070) & (!g2304) & (!g2305)) + ((g827) & (g1070) & (g2304) & (g2305)));
	assign g2307 = (((!g1005) & (!g1057) & (g1992) & (g1994) & (g2220)) + ((!g1005) & (g1057) & (!g1992) & (g1994) & (!g2220)) + ((!g1005) & (g1057) & (!g1992) & (g1994) & (g2220)) + ((!g1005) & (g1057) & (g1992) & (!g1994) & (g2220)) + ((!g1005) & (g1057) & (g1992) & (g1994) & (!g2220)) + ((!g1005) & (g1057) & (g1992) & (g1994) & (g2220)) + ((g1005) & (!g1057) & (!g1992) & (g1994) & (g2220)) + ((g1005) & (!g1057) & (g1992) & (g1994) & (!g2220)) + ((g1005) & (!g1057) & (g1992) & (g1994) & (g2220)) + ((g1005) & (g1057) & (!g1992) & (!g1994) & (g2220)) + ((g1005) & (g1057) & (!g1992) & (g1994) & (!g2220)) + ((g1005) & (g1057) & (!g1992) & (g1994) & (g2220)) + ((g1005) & (g1057) & (g1992) & (!g1994) & (!g2220)) + ((g1005) & (g1057) & (g1992) & (!g1994) & (g2220)) + ((g1005) & (g1057) & (g1992) & (g1994) & (!g2220)) + ((g1005) & (g1057) & (g1992) & (g1994) & (g2220)));
	assign g2308 = (((!g827) & (!g1072) & (g1997) & (!g2307)) + ((!g827) & (!g1072) & (g1997) & (g2307)) + ((!g827) & (g1072) & (g1997) & (!g2307)) + ((!g827) & (g1072) & (g1997) & (g2307)) + ((g827) & (!g1072) & (!g1997) & (g2307)) + ((g827) & (!g1072) & (g1997) & (!g2307)) + ((g827) & (g1072) & (!g1997) & (!g2307)) + ((g827) & (g1072) & (g1997) & (g2307)));
	assign g2309 = (((!g1007) & (!g1035) & (g1953) & (g1955) & (g2222)) + ((!g1007) & (g1035) & (!g1953) & (g1955) & (!g2222)) + ((!g1007) & (g1035) & (!g1953) & (g1955) & (g2222)) + ((!g1007) & (g1035) & (g1953) & (!g1955) & (g2222)) + ((!g1007) & (g1035) & (g1953) & (g1955) & (!g2222)) + ((!g1007) & (g1035) & (g1953) & (g1955) & (g2222)) + ((g1007) & (!g1035) & (!g1953) & (g1955) & (g2222)) + ((g1007) & (!g1035) & (g1953) & (g1955) & (!g2222)) + ((g1007) & (!g1035) & (g1953) & (g1955) & (g2222)) + ((g1007) & (g1035) & (!g1953) & (!g1955) & (g2222)) + ((g1007) & (g1035) & (!g1953) & (g1955) & (!g2222)) + ((g1007) & (g1035) & (!g1953) & (g1955) & (g2222)) + ((g1007) & (g1035) & (g1953) & (!g1955) & (!g2222)) + ((g1007) & (g1035) & (g1953) & (!g1955) & (g2222)) + ((g1007) & (g1035) & (g1953) & (g1955) & (!g2222)) + ((g1007) & (g1035) & (g1953) & (g1955) & (g2222)));
	assign g2310 = (((!g827) & (!g1074) & (g1958) & (!g2309)) + ((!g827) & (!g1074) & (g1958) & (g2309)) + ((!g827) & (g1074) & (g1958) & (!g2309)) + ((!g827) & (g1074) & (g1958) & (g2309)) + ((g827) & (!g1074) & (!g1958) & (g2309)) + ((g827) & (!g1074) & (g1958) & (!g2309)) + ((g827) & (g1074) & (!g1958) & (!g2309)) + ((g827) & (g1074) & (g1958) & (g2309)));
	assign g7973 = (((!g2017) & (g6651) & (!g2311)) + ((!g2017) & (g6651) & (g2311)) + ((g2017) & (!g6651) & (g2311)) + ((g2017) & (g6651) & (g2311)));
	assign g2312 = (((!g1009) & (!g1043) & (g2224) & (g2271) & (g2225)) + ((!g1009) & (g1043) & (!g2224) & (g2271) & (!g2225)) + ((!g1009) & (g1043) & (!g2224) & (g2271) & (g2225)) + ((!g1009) & (g1043) & (g2224) & (!g2271) & (g2225)) + ((!g1009) & (g1043) & (g2224) & (g2271) & (!g2225)) + ((!g1009) & (g1043) & (g2224) & (g2271) & (g2225)) + ((g1009) & (!g1043) & (!g2224) & (g2271) & (g2225)) + ((g1009) & (!g1043) & (g2224) & (g2271) & (!g2225)) + ((g1009) & (!g1043) & (g2224) & (g2271) & (g2225)) + ((g1009) & (g1043) & (!g2224) & (!g2271) & (g2225)) + ((g1009) & (g1043) & (!g2224) & (g2271) & (!g2225)) + ((g1009) & (g1043) & (!g2224) & (g2271) & (g2225)) + ((g1009) & (g1043) & (g2224) & (!g2271) & (!g2225)) + ((g1009) & (g1043) & (g2224) & (!g2271) & (g2225)) + ((g1009) & (g1043) & (g2224) & (g2271) & (!g2225)) + ((g1009) & (g1043) & (g2224) & (g2271) & (g2225)));
	assign g2313 = (((!g827) & (!g1076) & (g2311) & (!g2312)) + ((!g827) & (!g1076) & (g2311) & (g2312)) + ((!g827) & (g1076) & (g2311) & (!g2312)) + ((!g827) & (g1076) & (g2311) & (g2312)) + ((g827) & (!g1076) & (!g2311) & (g2312)) + ((g827) & (!g1076) & (g2311) & (!g2312)) + ((g827) & (g1076) & (!g2311) & (!g2312)) + ((g827) & (g1076) & (g2311) & (g2312)));
	assign g7974 = (((!g3499) & (g4560) & (!g2314)) + ((!g3499) & (g4560) & (g2314)) + ((g3499) & (!g4560) & (g2314)) + ((g3499) & (g4560) & (g2314)));
	assign g2315 = (((!g1011) & (!g1051) & (g2227) & (g2279) & (g2228)) + ((!g1011) & (g1051) & (!g2227) & (g2279) & (!g2228)) + ((!g1011) & (g1051) & (!g2227) & (g2279) & (g2228)) + ((!g1011) & (g1051) & (g2227) & (!g2279) & (g2228)) + ((!g1011) & (g1051) & (g2227) & (g2279) & (!g2228)) + ((!g1011) & (g1051) & (g2227) & (g2279) & (g2228)) + ((g1011) & (!g1051) & (!g2227) & (g2279) & (g2228)) + ((g1011) & (!g1051) & (g2227) & (g2279) & (!g2228)) + ((g1011) & (!g1051) & (g2227) & (g2279) & (g2228)) + ((g1011) & (g1051) & (!g2227) & (!g2279) & (g2228)) + ((g1011) & (g1051) & (!g2227) & (g2279) & (!g2228)) + ((g1011) & (g1051) & (!g2227) & (g2279) & (g2228)) + ((g1011) & (g1051) & (g2227) & (!g2279) & (!g2228)) + ((g1011) & (g1051) & (g2227) & (!g2279) & (g2228)) + ((g1011) & (g1051) & (g2227) & (g2279) & (!g2228)) + ((g1011) & (g1051) & (g2227) & (g2279) & (g2228)));
	assign g2316 = (((!g827) & (!g1078) & (g2314) & (!g2315)) + ((!g827) & (!g1078) & (g2314) & (g2315)) + ((!g827) & (g1078) & (g2314) & (!g2315)) + ((!g827) & (g1078) & (g2314) & (g2315)) + ((g827) & (!g1078) & (!g2314) & (g2315)) + ((g827) & (!g1078) & (g2314) & (!g2315)) + ((g827) & (g1078) & (!g2314) & (!g2315)) + ((g827) & (g1078) & (g2314) & (g2315)));
	assign g7975 = (((!g3464) & (g4564) & (!g2317)) + ((!g3464) & (g4564) & (g2317)) + ((g3464) & (!g4564) & (g2317)) + ((g3464) & (g4564) & (g2317)));
	assign g2318 = (((!g1013) & (!g1059) & (g2230) & (g2286) & (g2231)) + ((!g1013) & (g1059) & (!g2230) & (g2286) & (!g2231)) + ((!g1013) & (g1059) & (!g2230) & (g2286) & (g2231)) + ((!g1013) & (g1059) & (g2230) & (!g2286) & (g2231)) + ((!g1013) & (g1059) & (g2230) & (g2286) & (!g2231)) + ((!g1013) & (g1059) & (g2230) & (g2286) & (g2231)) + ((g1013) & (!g1059) & (!g2230) & (g2286) & (g2231)) + ((g1013) & (!g1059) & (g2230) & (g2286) & (!g2231)) + ((g1013) & (!g1059) & (g2230) & (g2286) & (g2231)) + ((g1013) & (g1059) & (!g2230) & (!g2286) & (g2231)) + ((g1013) & (g1059) & (!g2230) & (g2286) & (!g2231)) + ((g1013) & (g1059) & (!g2230) & (g2286) & (g2231)) + ((g1013) & (g1059) & (g2230) & (!g2286) & (!g2231)) + ((g1013) & (g1059) & (g2230) & (!g2286) & (g2231)) + ((g1013) & (g1059) & (g2230) & (g2286) & (!g2231)) + ((g1013) & (g1059) & (g2230) & (g2286) & (g2231)));
	assign g2319 = (((!g827) & (!g1080) & (g2317) & (!g2318)) + ((!g827) & (!g1080) & (g2317) & (g2318)) + ((!g827) & (g1080) & (g2317) & (!g2318)) + ((!g827) & (g1080) & (g2317) & (g2318)) + ((g827) & (!g1080) & (!g2317) & (g2318)) + ((g827) & (!g1080) & (g2317) & (!g2318)) + ((g827) & (g1080) & (!g2317) & (!g2318)) + ((g827) & (g1080) & (g2317) & (g2318)));
	assign g7976 = (((!g3499) & (g4568) & (!g2320)) + ((!g3499) & (g4568) & (g2320)) + ((g3499) & (!g4568) & (g2320)) + ((g3499) & (g4568) & (g2320)));
	assign g2321 = (((!g1015) & (!g1037) & (g2233) & (g2267) & (g2234)) + ((!g1015) & (g1037) & (!g2233) & (g2267) & (!g2234)) + ((!g1015) & (g1037) & (!g2233) & (g2267) & (g2234)) + ((!g1015) & (g1037) & (g2233) & (!g2267) & (g2234)) + ((!g1015) & (g1037) & (g2233) & (g2267) & (!g2234)) + ((!g1015) & (g1037) & (g2233) & (g2267) & (g2234)) + ((g1015) & (!g1037) & (!g2233) & (g2267) & (g2234)) + ((g1015) & (!g1037) & (g2233) & (g2267) & (!g2234)) + ((g1015) & (!g1037) & (g2233) & (g2267) & (g2234)) + ((g1015) & (g1037) & (!g2233) & (!g2267) & (g2234)) + ((g1015) & (g1037) & (!g2233) & (g2267) & (!g2234)) + ((g1015) & (g1037) & (!g2233) & (g2267) & (g2234)) + ((g1015) & (g1037) & (g2233) & (!g2267) & (!g2234)) + ((g1015) & (g1037) & (g2233) & (!g2267) & (g2234)) + ((g1015) & (g1037) & (g2233) & (g2267) & (!g2234)) + ((g1015) & (g1037) & (g2233) & (g2267) & (g2234)));
	assign g2322 = (((!g827) & (!g1082) & (g2320) & (!g2321)) + ((!g827) & (!g1082) & (g2320) & (g2321)) + ((!g827) & (g1082) & (g2320) & (!g2321)) + ((!g827) & (g1082) & (g2320) & (g2321)) + ((g827) & (!g1082) & (!g2320) & (g2321)) + ((g827) & (!g1082) & (g2320) & (!g2321)) + ((g827) & (g1082) & (!g2320) & (!g2321)) + ((g827) & (g1082) & (g2320) & (g2321)));
	assign g7977 = (((!g3464) & (g4573) & (!g2323)) + ((!g3464) & (g4573) & (g2323)) + ((g3464) & (!g4573) & (g2323)) + ((g3464) & (g4573) & (g2323)));
	assign g2324 = (((!g1017) & (!g1045) & (g2236) & (g2273) & (g2237)) + ((!g1017) & (g1045) & (!g2236) & (g2273) & (!g2237)) + ((!g1017) & (g1045) & (!g2236) & (g2273) & (g2237)) + ((!g1017) & (g1045) & (g2236) & (!g2273) & (g2237)) + ((!g1017) & (g1045) & (g2236) & (g2273) & (!g2237)) + ((!g1017) & (g1045) & (g2236) & (g2273) & (g2237)) + ((g1017) & (!g1045) & (!g2236) & (g2273) & (g2237)) + ((g1017) & (!g1045) & (g2236) & (g2273) & (!g2237)) + ((g1017) & (!g1045) & (g2236) & (g2273) & (g2237)) + ((g1017) & (g1045) & (!g2236) & (!g2273) & (g2237)) + ((g1017) & (g1045) & (!g2236) & (g2273) & (!g2237)) + ((g1017) & (g1045) & (!g2236) & (g2273) & (g2237)) + ((g1017) & (g1045) & (g2236) & (!g2273) & (!g2237)) + ((g1017) & (g1045) & (g2236) & (!g2273) & (g2237)) + ((g1017) & (g1045) & (g2236) & (g2273) & (!g2237)) + ((g1017) & (g1045) & (g2236) & (g2273) & (g2237)));
	assign g2325 = (((!g827) & (!g1084) & (g2323) & (!g2324)) + ((!g827) & (!g1084) & (g2323) & (g2324)) + ((!g827) & (g1084) & (g2323) & (!g2324)) + ((!g827) & (g1084) & (g2323) & (g2324)) + ((g827) & (!g1084) & (!g2323) & (g2324)) + ((g827) & (!g1084) & (g2323) & (!g2324)) + ((g827) & (g1084) & (!g2323) & (!g2324)) + ((g827) & (g1084) & (g2323) & (g2324)));
	assign g7978 = (((!g2017) & (g6645) & (!g2326)) + ((!g2017) & (g6645) & (g2326)) + ((g2017) & (!g6645) & (g2326)) + ((g2017) & (g6645) & (g2326)));
	assign g2327 = (((!g1019) & (!g1053) & (g2239) & (g2281) & (g2240)) + ((!g1019) & (g1053) & (!g2239) & (g2281) & (!g2240)) + ((!g1019) & (g1053) & (!g2239) & (g2281) & (g2240)) + ((!g1019) & (g1053) & (g2239) & (!g2281) & (g2240)) + ((!g1019) & (g1053) & (g2239) & (g2281) & (!g2240)) + ((!g1019) & (g1053) & (g2239) & (g2281) & (g2240)) + ((g1019) & (!g1053) & (!g2239) & (g2281) & (g2240)) + ((g1019) & (!g1053) & (g2239) & (g2281) & (!g2240)) + ((g1019) & (!g1053) & (g2239) & (g2281) & (g2240)) + ((g1019) & (g1053) & (!g2239) & (!g2281) & (g2240)) + ((g1019) & (g1053) & (!g2239) & (g2281) & (!g2240)) + ((g1019) & (g1053) & (!g2239) & (g2281) & (g2240)) + ((g1019) & (g1053) & (g2239) & (!g2281) & (!g2240)) + ((g1019) & (g1053) & (g2239) & (!g2281) & (g2240)) + ((g1019) & (g1053) & (g2239) & (g2281) & (!g2240)) + ((g1019) & (g1053) & (g2239) & (g2281) & (g2240)));
	assign g2328 = (((!g827) & (!g1086) & (g2326) & (!g2327)) + ((!g827) & (!g1086) & (g2326) & (g2327)) + ((!g827) & (g1086) & (g2326) & (!g2327)) + ((!g827) & (g1086) & (g2326) & (g2327)) + ((g827) & (!g1086) & (!g2326) & (g2327)) + ((g827) & (!g1086) & (g2326) & (!g2327)) + ((g827) & (g1086) & (!g2326) & (!g2327)) + ((g827) & (g1086) & (g2326) & (g2327)));
	assign g7979 = (((!g3429) & (g4578) & (!g2329)) + ((!g3429) & (g4578) & (g2329)) + ((g3429) & (!g4578) & (g2329)) + ((g3429) & (g4578) & (g2329)));
	assign g2330 = (((!g1021) & (!g1061) & (g2242) & (g2288) & (g2243)) + ((!g1021) & (g1061) & (!g2242) & (g2288) & (!g2243)) + ((!g1021) & (g1061) & (!g2242) & (g2288) & (g2243)) + ((!g1021) & (g1061) & (g2242) & (!g2288) & (g2243)) + ((!g1021) & (g1061) & (g2242) & (g2288) & (!g2243)) + ((!g1021) & (g1061) & (g2242) & (g2288) & (g2243)) + ((g1021) & (!g1061) & (!g2242) & (g2288) & (g2243)) + ((g1021) & (!g1061) & (g2242) & (g2288) & (!g2243)) + ((g1021) & (!g1061) & (g2242) & (g2288) & (g2243)) + ((g1021) & (g1061) & (!g2242) & (!g2288) & (g2243)) + ((g1021) & (g1061) & (!g2242) & (g2288) & (!g2243)) + ((g1021) & (g1061) & (!g2242) & (g2288) & (g2243)) + ((g1021) & (g1061) & (g2242) & (!g2288) & (!g2243)) + ((g1021) & (g1061) & (g2242) & (!g2288) & (g2243)) + ((g1021) & (g1061) & (g2242) & (g2288) & (!g2243)) + ((g1021) & (g1061) & (g2242) & (g2288) & (g2243)));
	assign g2331 = (((!g827) & (!g1088) & (g2329) & (!g2330)) + ((!g827) & (!g1088) & (g2329) & (g2330)) + ((!g827) & (g1088) & (g2329) & (!g2330)) + ((!g827) & (g1088) & (g2329) & (g2330)) + ((g827) & (!g1088) & (!g2329) & (g2330)) + ((g827) & (!g1088) & (g2329) & (!g2330)) + ((g827) & (g1088) & (!g2329) & (!g2330)) + ((g827) & (g1088) & (g2329) & (g2330)));
	assign g2332 = (((!g1023) & (!g1039) & (g1954) & (g1956) & (g2245)) + ((!g1023) & (g1039) & (!g1954) & (g1956) & (!g2245)) + ((!g1023) & (g1039) & (!g1954) & (g1956) & (g2245)) + ((!g1023) & (g1039) & (g1954) & (!g1956) & (g2245)) + ((!g1023) & (g1039) & (g1954) & (g1956) & (!g2245)) + ((!g1023) & (g1039) & (g1954) & (g1956) & (g2245)) + ((g1023) & (!g1039) & (!g1954) & (g1956) & (g2245)) + ((g1023) & (!g1039) & (g1954) & (g1956) & (!g2245)) + ((g1023) & (!g1039) & (g1954) & (g1956) & (g2245)) + ((g1023) & (g1039) & (!g1954) & (!g1956) & (g2245)) + ((g1023) & (g1039) & (!g1954) & (g1956) & (!g2245)) + ((g1023) & (g1039) & (!g1954) & (g1956) & (g2245)) + ((g1023) & (g1039) & (g1954) & (!g1956) & (!g2245)) + ((g1023) & (g1039) & (g1954) & (!g1956) & (g2245)) + ((g1023) & (g1039) & (g1954) & (g1956) & (!g2245)) + ((g1023) & (g1039) & (g1954) & (g1956) & (g2245)));
	assign g2333 = (((!g827) & (!g1090) & (g1959) & (!g2332)) + ((!g827) & (!g1090) & (g1959) & (g2332)) + ((!g827) & (g1090) & (g1959) & (!g2332)) + ((!g827) & (g1090) & (g1959) & (g2332)) + ((g827) & (!g1090) & (!g1959) & (g2332)) + ((g827) & (!g1090) & (g1959) & (!g2332)) + ((g827) & (g1090) & (!g1959) & (!g2332)) + ((g827) & (g1090) & (g1959) & (g2332)));
	assign g7980 = (((!g3499) & (g4582) & (!g2334)) + ((!g3499) & (g4582) & (g2334)) + ((g3499) & (!g4582) & (g2334)) + ((g3499) & (g4582) & (g2334)));
	assign g2335 = (((!g1025) & (!g1047) & (g2247) & (g2275) & (g2248)) + ((!g1025) & (g1047) & (!g2247) & (g2275) & (!g2248)) + ((!g1025) & (g1047) & (!g2247) & (g2275) & (g2248)) + ((!g1025) & (g1047) & (g2247) & (!g2275) & (g2248)) + ((!g1025) & (g1047) & (g2247) & (g2275) & (!g2248)) + ((!g1025) & (g1047) & (g2247) & (g2275) & (g2248)) + ((g1025) & (!g1047) & (!g2247) & (g2275) & (g2248)) + ((g1025) & (!g1047) & (g2247) & (g2275) & (!g2248)) + ((g1025) & (!g1047) & (g2247) & (g2275) & (g2248)) + ((g1025) & (g1047) & (!g2247) & (!g2275) & (g2248)) + ((g1025) & (g1047) & (!g2247) & (g2275) & (!g2248)) + ((g1025) & (g1047) & (!g2247) & (g2275) & (g2248)) + ((g1025) & (g1047) & (g2247) & (!g2275) & (!g2248)) + ((g1025) & (g1047) & (g2247) & (!g2275) & (g2248)) + ((g1025) & (g1047) & (g2247) & (g2275) & (!g2248)) + ((g1025) & (g1047) & (g2247) & (g2275) & (g2248)));
	assign g2336 = (((!g827) & (!g1092) & (g2334) & (!g2335)) + ((!g827) & (!g1092) & (g2334) & (g2335)) + ((!g827) & (g1092) & (g2334) & (!g2335)) + ((!g827) & (g1092) & (g2334) & (g2335)) + ((g827) & (!g1092) & (!g2334) & (g2335)) + ((g827) & (!g1092) & (g2334) & (!g2335)) + ((g827) & (g1092) & (!g2334) & (!g2335)) + ((g827) & (g1092) & (g2334) & (g2335)));
	assign g7981 = (((!g3429) & (g4585) & (!g2337)) + ((!g3429) & (g4585) & (g2337)) + ((g3429) & (!g4585) & (g2337)) + ((g3429) & (g4585) & (g2337)));
	assign g2338 = (((!g1027) & (!g1055) & (g2250) & (g2283) & (g2251)) + ((!g1027) & (g1055) & (!g2250) & (g2283) & (!g2251)) + ((!g1027) & (g1055) & (!g2250) & (g2283) & (g2251)) + ((!g1027) & (g1055) & (g2250) & (!g2283) & (g2251)) + ((!g1027) & (g1055) & (g2250) & (g2283) & (!g2251)) + ((!g1027) & (g1055) & (g2250) & (g2283) & (g2251)) + ((g1027) & (!g1055) & (!g2250) & (g2283) & (g2251)) + ((g1027) & (!g1055) & (g2250) & (g2283) & (!g2251)) + ((g1027) & (!g1055) & (g2250) & (g2283) & (g2251)) + ((g1027) & (g1055) & (!g2250) & (!g2283) & (g2251)) + ((g1027) & (g1055) & (!g2250) & (g2283) & (!g2251)) + ((g1027) & (g1055) & (!g2250) & (g2283) & (g2251)) + ((g1027) & (g1055) & (g2250) & (!g2283) & (!g2251)) + ((g1027) & (g1055) & (g2250) & (!g2283) & (g2251)) + ((g1027) & (g1055) & (g2250) & (g2283) & (!g2251)) + ((g1027) & (g1055) & (g2250) & (g2283) & (g2251)));
	assign g2339 = (((!g827) & (!g1094) & (g2337) & (!g2338)) + ((!g827) & (!g1094) & (g2337) & (g2338)) + ((!g827) & (g1094) & (g2337) & (!g2338)) + ((!g827) & (g1094) & (g2337) & (g2338)) + ((g827) & (!g1094) & (!g2337) & (g2338)) + ((g827) & (!g1094) & (g2337) & (!g2338)) + ((g827) & (g1094) & (!g2337) & (!g2338)) + ((g827) & (g1094) & (g2337) & (g2338)));
	assign g7982 = (((!g2017) & (g6638) & (!g2340)) + ((!g2017) & (g6638) & (g2340)) + ((g2017) & (!g6638) & (g2340)) + ((g2017) & (g6638) & (g2340)));
	assign g2341 = (((!g1029) & (!g1063) & (g2253) & (g2290) & (g2254)) + ((!g1029) & (g1063) & (!g2253) & (g2290) & (!g2254)) + ((!g1029) & (g1063) & (!g2253) & (g2290) & (g2254)) + ((!g1029) & (g1063) & (g2253) & (!g2290) & (g2254)) + ((!g1029) & (g1063) & (g2253) & (g2290) & (!g2254)) + ((!g1029) & (g1063) & (g2253) & (g2290) & (g2254)) + ((g1029) & (!g1063) & (!g2253) & (g2290) & (g2254)) + ((g1029) & (!g1063) & (g2253) & (g2290) & (!g2254)) + ((g1029) & (!g1063) & (g2253) & (g2290) & (g2254)) + ((g1029) & (g1063) & (!g2253) & (!g2290) & (g2254)) + ((g1029) & (g1063) & (!g2253) & (g2290) & (!g2254)) + ((g1029) & (g1063) & (!g2253) & (g2290) & (g2254)) + ((g1029) & (g1063) & (g2253) & (!g2290) & (!g2254)) + ((g1029) & (g1063) & (g2253) & (!g2290) & (g2254)) + ((g1029) & (g1063) & (g2253) & (g2290) & (!g2254)) + ((g1029) & (g1063) & (g2253) & (g2290) & (g2254)));
	assign g2342 = (((!g827) & (!g1096) & (g2340) & (!g2341)) + ((!g827) & (!g1096) & (g2340) & (g2341)) + ((!g827) & (g1096) & (g2340) & (!g2341)) + ((!g827) & (g1096) & (g2340) & (g2341)) + ((g827) & (!g1096) & (!g2340) & (g2341)) + ((g827) & (!g1096) & (g2340) & (!g2341)) + ((g827) & (g1096) & (!g2340) & (!g2341)) + ((g827) & (g1096) & (g2340) & (g2341)));
	assign g7983 = (((!g3429) & (g4590) & (!g2343)) + ((!g3429) & (g4590) & (g2343)) + ((g3429) & (!g4590) & (g2343)) + ((g3429) & (g4590) & (g2343)));
	assign g7984 = (((!g3464) & (g4593) & (!g2344)) + ((!g3464) & (g4593) & (g2344)) + ((g3464) & (!g4593) & (g2344)) + ((g3464) & (g4593) & (g2344)));
	assign g2345 = (((!g2293) & (!g2294) & (!g2295) & (!g2296) & (!g2343) & (g2344)) + ((!g2293) & (!g2294) & (!g2295) & (!g2296) & (g2343) & (!g2344)) + ((!g2293) & (!g2294) & (!g2295) & (g2296) & (!g2343) & (g2344)) + ((!g2293) & (!g2294) & (!g2295) & (g2296) & (g2343) & (!g2344)) + ((!g2293) & (!g2294) & (g2295) & (!g2296) & (!g2343) & (g2344)) + ((!g2293) & (!g2294) & (g2295) & (!g2296) & (g2343) & (!g2344)) + ((!g2293) & (!g2294) & (g2295) & (g2296) & (!g2343) & (!g2344)) + ((!g2293) & (!g2294) & (g2295) & (g2296) & (g2343) & (g2344)) + ((!g2293) & (g2294) & (!g2295) & (!g2296) & (!g2343) & (g2344)) + ((!g2293) & (g2294) & (!g2295) & (!g2296) & (g2343) & (!g2344)) + ((!g2293) & (g2294) & (!g2295) & (g2296) & (!g2343) & (!g2344)) + ((!g2293) & (g2294) & (!g2295) & (g2296) & (g2343) & (g2344)) + ((!g2293) & (g2294) & (g2295) & (!g2296) & (!g2343) & (!g2344)) + ((!g2293) & (g2294) & (g2295) & (!g2296) & (g2343) & (g2344)) + ((!g2293) & (g2294) & (g2295) & (g2296) & (!g2343) & (!g2344)) + ((!g2293) & (g2294) & (g2295) & (g2296) & (g2343) & (g2344)) + ((g2293) & (!g2294) & (!g2295) & (!g2296) & (!g2343) & (g2344)) + ((g2293) & (!g2294) & (!g2295) & (!g2296) & (g2343) & (!g2344)) + ((g2293) & (!g2294) & (!g2295) & (g2296) & (!g2343) & (!g2344)) + ((g2293) & (!g2294) & (!g2295) & (g2296) & (g2343) & (g2344)) + ((g2293) & (!g2294) & (g2295) & (!g2296) & (!g2343) & (!g2344)) + ((g2293) & (!g2294) & (g2295) & (!g2296) & (g2343) & (g2344)) + ((g2293) & (!g2294) & (g2295) & (g2296) & (!g2343) & (!g2344)) + ((g2293) & (!g2294) & (g2295) & (g2296) & (g2343) & (g2344)) + ((g2293) & (g2294) & (!g2295) & (!g2296) & (!g2343) & (g2344)) + ((g2293) & (g2294) & (!g2295) & (!g2296) & (g2343) & (!g2344)) + ((g2293) & (g2294) & (!g2295) & (g2296) & (!g2343) & (!g2344)) + ((g2293) & (g2294) & (!g2295) & (g2296) & (g2343) & (g2344)) + ((g2293) & (g2294) & (g2295) & (!g2296) & (!g2343) & (!g2344)) + ((g2293) & (g2294) & (g2295) & (!g2296) & (g2343) & (g2344)) + ((g2293) & (g2294) & (g2295) & (g2296) & (!g2343) & (!g2344)) + ((g2293) & (g2294) & (g2295) & (g2296) & (g2343) & (g2344)));
	assign g2346 = (((!g2260) & (!g2261) & (!g2262) & (!g2263) & (g2298) & (g2299)) + ((!g2260) & (!g2261) & (!g2262) & (g2263) & (g2298) & (g2299)) + ((!g2260) & (!g2261) & (g2262) & (!g2263) & (g2298) & (g2299)) + ((!g2260) & (!g2261) & (g2262) & (g2263) & (!g2298) & (g2299)) + ((!g2260) & (!g2261) & (g2262) & (g2263) & (g2298) & (!g2299)) + ((!g2260) & (!g2261) & (g2262) & (g2263) & (g2298) & (g2299)) + ((!g2260) & (g2261) & (!g2262) & (!g2263) & (g2298) & (g2299)) + ((!g2260) & (g2261) & (!g2262) & (g2263) & (!g2298) & (g2299)) + ((!g2260) & (g2261) & (!g2262) & (g2263) & (g2298) & (!g2299)) + ((!g2260) & (g2261) & (!g2262) & (g2263) & (g2298) & (g2299)) + ((!g2260) & (g2261) & (g2262) & (!g2263) & (!g2298) & (g2299)) + ((!g2260) & (g2261) & (g2262) & (!g2263) & (g2298) & (!g2299)) + ((!g2260) & (g2261) & (g2262) & (!g2263) & (g2298) & (g2299)) + ((!g2260) & (g2261) & (g2262) & (g2263) & (!g2298) & (g2299)) + ((!g2260) & (g2261) & (g2262) & (g2263) & (g2298) & (!g2299)) + ((!g2260) & (g2261) & (g2262) & (g2263) & (g2298) & (g2299)) + ((g2260) & (!g2261) & (!g2262) & (!g2263) & (g2298) & (g2299)) + ((g2260) & (!g2261) & (!g2262) & (g2263) & (!g2298) & (g2299)) + ((g2260) & (!g2261) & (!g2262) & (g2263) & (g2298) & (!g2299)) + ((g2260) & (!g2261) & (!g2262) & (g2263) & (g2298) & (g2299)) + ((g2260) & (!g2261) & (g2262) & (!g2263) & (!g2298) & (g2299)) + ((g2260) & (!g2261) & (g2262) & (!g2263) & (g2298) & (!g2299)) + ((g2260) & (!g2261) & (g2262) & (!g2263) & (g2298) & (g2299)) + ((g2260) & (!g2261) & (g2262) & (g2263) & (!g2298) & (g2299)) + ((g2260) & (!g2261) & (g2262) & (g2263) & (g2298) & (!g2299)) + ((g2260) & (!g2261) & (g2262) & (g2263) & (g2298) & (g2299)) + ((g2260) & (g2261) & (!g2262) & (!g2263) & (g2298) & (g2299)) + ((g2260) & (g2261) & (!g2262) & (g2263) & (!g2298) & (g2299)) + ((g2260) & (g2261) & (!g2262) & (g2263) & (g2298) & (!g2299)) + ((g2260) & (g2261) & (!g2262) & (g2263) & (g2298) & (g2299)) + ((g2260) & (g2261) & (g2262) & (!g2263) & (!g2298) & (g2299)) + ((g2260) & (g2261) & (g2262) & (!g2263) & (g2298) & (!g2299)) + ((g2260) & (g2261) & (g2262) & (!g2263) & (g2298) & (g2299)) + ((g2260) & (g2261) & (g2262) & (g2263) & (!g2298) & (g2299)) + ((g2260) & (g2261) & (g2262) & (g2263) & (g2298) & (!g2299)) + ((g2260) & (g2261) & (g2262) & (g2263) & (g2298) & (g2299)));
	assign g7985 = (((!g3429) & (g4597) & (!g2347)) + ((!g3429) & (g4597) & (g2347)) + ((g3429) & (!g4597) & (g2347)) + ((g3429) & (g4597) & (g2347)));
	assign g7986 = (((!g3499) & (g4600) & (!g2348)) + ((!g3499) & (g4600) & (g2348)) + ((g3499) & (!g4600) & (g2348)) + ((g3499) & (g4600) & (g2348)));
	assign g2349 = (((!g827) & (!g1074) & (!g1102) & (!g1958) & (g1960) & (!g2309)) + ((!g827) & (!g1074) & (!g1102) & (!g1958) & (g1960) & (g2309)) + ((!g827) & (!g1074) & (!g1102) & (g1958) & (g1960) & (!g2309)) + ((!g827) & (!g1074) & (!g1102) & (g1958) & (g1960) & (g2309)) + ((!g827) & (!g1074) & (g1102) & (!g1958) & (g1960) & (!g2309)) + ((!g827) & (!g1074) & (g1102) & (!g1958) & (g1960) & (g2309)) + ((!g827) & (!g1074) & (g1102) & (g1958) & (g1960) & (!g2309)) + ((!g827) & (!g1074) & (g1102) & (g1958) & (g1960) & (g2309)) + ((!g827) & (g1074) & (!g1102) & (!g1958) & (g1960) & (!g2309)) + ((!g827) & (g1074) & (!g1102) & (!g1958) & (g1960) & (g2309)) + ((!g827) & (g1074) & (!g1102) & (g1958) & (g1960) & (!g2309)) + ((!g827) & (g1074) & (!g1102) & (g1958) & (g1960) & (g2309)) + ((!g827) & (g1074) & (g1102) & (!g1958) & (g1960) & (!g2309)) + ((!g827) & (g1074) & (g1102) & (!g1958) & (g1960) & (g2309)) + ((!g827) & (g1074) & (g1102) & (g1958) & (g1960) & (!g2309)) + ((!g827) & (g1074) & (g1102) & (g1958) & (g1960) & (g2309)) + ((g827) & (!g1074) & (!g1102) & (!g1958) & (g1960) & (!g2309)) + ((g827) & (!g1074) & (!g1102) & (!g1958) & (g1960) & (g2309)) + ((g827) & (!g1074) & (!g1102) & (g1958) & (!g1960) & (g2309)) + ((g827) & (!g1074) & (!g1102) & (g1958) & (g1960) & (!g2309)) + ((g827) & (!g1074) & (g1102) & (!g1958) & (!g1960) & (!g2309)) + ((g827) & (!g1074) & (g1102) & (!g1958) & (!g1960) & (g2309)) + ((g827) & (!g1074) & (g1102) & (g1958) & (!g1960) & (!g2309)) + ((g827) & (!g1074) & (g1102) & (g1958) & (g1960) & (g2309)) + ((g827) & (g1074) & (!g1102) & (!g1958) & (!g1960) & (g2309)) + ((g827) & (g1074) & (!g1102) & (!g1958) & (g1960) & (!g2309)) + ((g827) & (g1074) & (!g1102) & (g1958) & (!g1960) & (!g2309)) + ((g827) & (g1074) & (!g1102) & (g1958) & (!g1960) & (g2309)) + ((g827) & (g1074) & (g1102) & (!g1958) & (!g1960) & (!g2309)) + ((g827) & (g1074) & (g1102) & (!g1958) & (g1960) & (g2309)) + ((g827) & (g1074) & (g1102) & (g1958) & (g1960) & (!g2309)) + ((g827) & (g1074) & (g1102) & (g1958) & (g1960) & (g2309)));
	assign g7987 = (((!g3499) & (g4604) & (!g2350)) + ((!g3499) & (g4604) & (g2350)) + ((g3499) & (!g4604) & (g2350)) + ((g3499) & (g4604) & (g2350)));
	assign g2351 = (((!g827) & (!g1082) & (!g1104) & (!g2320) & (g2350) & (!g2321)) + ((!g827) & (!g1082) & (!g1104) & (!g2320) & (g2350) & (g2321)) + ((!g827) & (!g1082) & (!g1104) & (g2320) & (g2350) & (!g2321)) + ((!g827) & (!g1082) & (!g1104) & (g2320) & (g2350) & (g2321)) + ((!g827) & (!g1082) & (g1104) & (!g2320) & (g2350) & (!g2321)) + ((!g827) & (!g1082) & (g1104) & (!g2320) & (g2350) & (g2321)) + ((!g827) & (!g1082) & (g1104) & (g2320) & (g2350) & (!g2321)) + ((!g827) & (!g1082) & (g1104) & (g2320) & (g2350) & (g2321)) + ((!g827) & (g1082) & (!g1104) & (!g2320) & (g2350) & (!g2321)) + ((!g827) & (g1082) & (!g1104) & (!g2320) & (g2350) & (g2321)) + ((!g827) & (g1082) & (!g1104) & (g2320) & (g2350) & (!g2321)) + ((!g827) & (g1082) & (!g1104) & (g2320) & (g2350) & (g2321)) + ((!g827) & (g1082) & (g1104) & (!g2320) & (g2350) & (!g2321)) + ((!g827) & (g1082) & (g1104) & (!g2320) & (g2350) & (g2321)) + ((!g827) & (g1082) & (g1104) & (g2320) & (g2350) & (!g2321)) + ((!g827) & (g1082) & (g1104) & (g2320) & (g2350) & (g2321)) + ((g827) & (!g1082) & (!g1104) & (!g2320) & (g2350) & (!g2321)) + ((g827) & (!g1082) & (!g1104) & (!g2320) & (g2350) & (g2321)) + ((g827) & (!g1082) & (!g1104) & (g2320) & (!g2350) & (g2321)) + ((g827) & (!g1082) & (!g1104) & (g2320) & (g2350) & (!g2321)) + ((g827) & (!g1082) & (g1104) & (!g2320) & (!g2350) & (!g2321)) + ((g827) & (!g1082) & (g1104) & (!g2320) & (!g2350) & (g2321)) + ((g827) & (!g1082) & (g1104) & (g2320) & (!g2350) & (!g2321)) + ((g827) & (!g1082) & (g1104) & (g2320) & (g2350) & (g2321)) + ((g827) & (g1082) & (!g1104) & (!g2320) & (!g2350) & (g2321)) + ((g827) & (g1082) & (!g1104) & (!g2320) & (g2350) & (!g2321)) + ((g827) & (g1082) & (!g1104) & (g2320) & (!g2350) & (!g2321)) + ((g827) & (g1082) & (!g1104) & (g2320) & (!g2350) & (g2321)) + ((g827) & (g1082) & (g1104) & (!g2320) & (!g2350) & (!g2321)) + ((g827) & (g1082) & (g1104) & (!g2320) & (g2350) & (g2321)) + ((g827) & (g1082) & (g1104) & (g2320) & (g2350) & (!g2321)) + ((g827) & (g1082) & (g1104) & (g2320) & (g2350) & (g2321)));
	assign g2352 = (((!g827) & (!g1090) & (!g1106) & (!g1959) & (g1961) & (!g2332)) + ((!g827) & (!g1090) & (!g1106) & (!g1959) & (g1961) & (g2332)) + ((!g827) & (!g1090) & (!g1106) & (g1959) & (g1961) & (!g2332)) + ((!g827) & (!g1090) & (!g1106) & (g1959) & (g1961) & (g2332)) + ((!g827) & (!g1090) & (g1106) & (!g1959) & (g1961) & (!g2332)) + ((!g827) & (!g1090) & (g1106) & (!g1959) & (g1961) & (g2332)) + ((!g827) & (!g1090) & (g1106) & (g1959) & (g1961) & (!g2332)) + ((!g827) & (!g1090) & (g1106) & (g1959) & (g1961) & (g2332)) + ((!g827) & (g1090) & (!g1106) & (!g1959) & (g1961) & (!g2332)) + ((!g827) & (g1090) & (!g1106) & (!g1959) & (g1961) & (g2332)) + ((!g827) & (g1090) & (!g1106) & (g1959) & (g1961) & (!g2332)) + ((!g827) & (g1090) & (!g1106) & (g1959) & (g1961) & (g2332)) + ((!g827) & (g1090) & (g1106) & (!g1959) & (g1961) & (!g2332)) + ((!g827) & (g1090) & (g1106) & (!g1959) & (g1961) & (g2332)) + ((!g827) & (g1090) & (g1106) & (g1959) & (g1961) & (!g2332)) + ((!g827) & (g1090) & (g1106) & (g1959) & (g1961) & (g2332)) + ((g827) & (!g1090) & (!g1106) & (!g1959) & (g1961) & (!g2332)) + ((g827) & (!g1090) & (!g1106) & (!g1959) & (g1961) & (g2332)) + ((g827) & (!g1090) & (!g1106) & (g1959) & (!g1961) & (g2332)) + ((g827) & (!g1090) & (!g1106) & (g1959) & (g1961) & (!g2332)) + ((g827) & (!g1090) & (g1106) & (!g1959) & (!g1961) & (!g2332)) + ((g827) & (!g1090) & (g1106) & (!g1959) & (!g1961) & (g2332)) + ((g827) & (!g1090) & (g1106) & (g1959) & (!g1961) & (!g2332)) + ((g827) & (!g1090) & (g1106) & (g1959) & (g1961) & (g2332)) + ((g827) & (g1090) & (!g1106) & (!g1959) & (!g1961) & (g2332)) + ((g827) & (g1090) & (!g1106) & (!g1959) & (g1961) & (!g2332)) + ((g827) & (g1090) & (!g1106) & (g1959) & (!g1961) & (!g2332)) + ((g827) & (g1090) & (!g1106) & (g1959) & (!g1961) & (g2332)) + ((g827) & (g1090) & (g1106) & (!g1959) & (!g1961) & (!g2332)) + ((g827) & (g1090) & (g1106) & (!g1959) & (g1961) & (g2332)) + ((g827) & (g1090) & (g1106) & (g1959) & (g1961) & (!g2332)) + ((g827) & (g1090) & (g1106) & (g1959) & (g1961) & (g2332)));
	assign g2353 = (((!g827) & (!g1068) & (!g1108) & (!g1996) & (g1998) & (!g2302)) + ((!g827) & (!g1068) & (!g1108) & (!g1996) & (g1998) & (g2302)) + ((!g827) & (!g1068) & (!g1108) & (g1996) & (g1998) & (!g2302)) + ((!g827) & (!g1068) & (!g1108) & (g1996) & (g1998) & (g2302)) + ((!g827) & (!g1068) & (g1108) & (!g1996) & (g1998) & (!g2302)) + ((!g827) & (!g1068) & (g1108) & (!g1996) & (g1998) & (g2302)) + ((!g827) & (!g1068) & (g1108) & (g1996) & (g1998) & (!g2302)) + ((!g827) & (!g1068) & (g1108) & (g1996) & (g1998) & (g2302)) + ((!g827) & (g1068) & (!g1108) & (!g1996) & (g1998) & (!g2302)) + ((!g827) & (g1068) & (!g1108) & (!g1996) & (g1998) & (g2302)) + ((!g827) & (g1068) & (!g1108) & (g1996) & (g1998) & (!g2302)) + ((!g827) & (g1068) & (!g1108) & (g1996) & (g1998) & (g2302)) + ((!g827) & (g1068) & (g1108) & (!g1996) & (g1998) & (!g2302)) + ((!g827) & (g1068) & (g1108) & (!g1996) & (g1998) & (g2302)) + ((!g827) & (g1068) & (g1108) & (g1996) & (g1998) & (!g2302)) + ((!g827) & (g1068) & (g1108) & (g1996) & (g1998) & (g2302)) + ((g827) & (!g1068) & (!g1108) & (!g1996) & (g1998) & (!g2302)) + ((g827) & (!g1068) & (!g1108) & (!g1996) & (g1998) & (g2302)) + ((g827) & (!g1068) & (!g1108) & (g1996) & (!g1998) & (g2302)) + ((g827) & (!g1068) & (!g1108) & (g1996) & (g1998) & (!g2302)) + ((g827) & (!g1068) & (g1108) & (!g1996) & (!g1998) & (!g2302)) + ((g827) & (!g1068) & (g1108) & (!g1996) & (!g1998) & (g2302)) + ((g827) & (!g1068) & (g1108) & (g1996) & (!g1998) & (!g2302)) + ((g827) & (!g1068) & (g1108) & (g1996) & (g1998) & (g2302)) + ((g827) & (g1068) & (!g1108) & (!g1996) & (!g1998) & (g2302)) + ((g827) & (g1068) & (!g1108) & (!g1996) & (g1998) & (!g2302)) + ((g827) & (g1068) & (!g1108) & (g1996) & (!g1998) & (!g2302)) + ((g827) & (g1068) & (!g1108) & (g1996) & (!g1998) & (g2302)) + ((g827) & (g1068) & (g1108) & (!g1996) & (!g1998) & (!g2302)) + ((g827) & (g1068) & (g1108) & (!g1996) & (g1998) & (g2302)) + ((g827) & (g1068) & (g1108) & (g1996) & (g1998) & (!g2302)) + ((g827) & (g1068) & (g1108) & (g1996) & (g1998) & (g2302)));
	assign g7988 = (((!g2017) & (g6610) & (!g2354)) + ((!g2017) & (g6610) & (g2354)) + ((g2017) & (!g6610) & (g2354)) + ((g2017) & (g6610) & (g2354)));
	assign g2355 = (((!g827) & (!g1076) & (!g1110) & (!g2311) & (g2354) & (!g2312)) + ((!g827) & (!g1076) & (!g1110) & (!g2311) & (g2354) & (g2312)) + ((!g827) & (!g1076) & (!g1110) & (g2311) & (g2354) & (!g2312)) + ((!g827) & (!g1076) & (!g1110) & (g2311) & (g2354) & (g2312)) + ((!g827) & (!g1076) & (g1110) & (!g2311) & (g2354) & (!g2312)) + ((!g827) & (!g1076) & (g1110) & (!g2311) & (g2354) & (g2312)) + ((!g827) & (!g1076) & (g1110) & (g2311) & (g2354) & (!g2312)) + ((!g827) & (!g1076) & (g1110) & (g2311) & (g2354) & (g2312)) + ((!g827) & (g1076) & (!g1110) & (!g2311) & (g2354) & (!g2312)) + ((!g827) & (g1076) & (!g1110) & (!g2311) & (g2354) & (g2312)) + ((!g827) & (g1076) & (!g1110) & (g2311) & (g2354) & (!g2312)) + ((!g827) & (g1076) & (!g1110) & (g2311) & (g2354) & (g2312)) + ((!g827) & (g1076) & (g1110) & (!g2311) & (g2354) & (!g2312)) + ((!g827) & (g1076) & (g1110) & (!g2311) & (g2354) & (g2312)) + ((!g827) & (g1076) & (g1110) & (g2311) & (g2354) & (!g2312)) + ((!g827) & (g1076) & (g1110) & (g2311) & (g2354) & (g2312)) + ((g827) & (!g1076) & (!g1110) & (!g2311) & (g2354) & (!g2312)) + ((g827) & (!g1076) & (!g1110) & (!g2311) & (g2354) & (g2312)) + ((g827) & (!g1076) & (!g1110) & (g2311) & (!g2354) & (g2312)) + ((g827) & (!g1076) & (!g1110) & (g2311) & (g2354) & (!g2312)) + ((g827) & (!g1076) & (g1110) & (!g2311) & (!g2354) & (!g2312)) + ((g827) & (!g1076) & (g1110) & (!g2311) & (!g2354) & (g2312)) + ((g827) & (!g1076) & (g1110) & (g2311) & (!g2354) & (!g2312)) + ((g827) & (!g1076) & (g1110) & (g2311) & (g2354) & (g2312)) + ((g827) & (g1076) & (!g1110) & (!g2311) & (!g2354) & (g2312)) + ((g827) & (g1076) & (!g1110) & (!g2311) & (g2354) & (!g2312)) + ((g827) & (g1076) & (!g1110) & (g2311) & (!g2354) & (!g2312)) + ((g827) & (g1076) & (!g1110) & (g2311) & (!g2354) & (g2312)) + ((g827) & (g1076) & (g1110) & (!g2311) & (!g2354) & (!g2312)) + ((g827) & (g1076) & (g1110) & (!g2311) & (g2354) & (g2312)) + ((g827) & (g1076) & (g1110) & (g2311) & (g2354) & (!g2312)) + ((g827) & (g1076) & (g1110) & (g2311) & (g2354) & (g2312)));
	assign g7989 = (((!g3464) & (g4611) & (!g2356)) + ((!g3464) & (g4611) & (g2356)) + ((g3464) & (!g4611) & (g2356)) + ((g3464) & (g4611) & (g2356)));
	assign g2357 = (((!g827) & (!g1084) & (!g1112) & (!g2323) & (g2356) & (!g2324)) + ((!g827) & (!g1084) & (!g1112) & (!g2323) & (g2356) & (g2324)) + ((!g827) & (!g1084) & (!g1112) & (g2323) & (g2356) & (!g2324)) + ((!g827) & (!g1084) & (!g1112) & (g2323) & (g2356) & (g2324)) + ((!g827) & (!g1084) & (g1112) & (!g2323) & (g2356) & (!g2324)) + ((!g827) & (!g1084) & (g1112) & (!g2323) & (g2356) & (g2324)) + ((!g827) & (!g1084) & (g1112) & (g2323) & (g2356) & (!g2324)) + ((!g827) & (!g1084) & (g1112) & (g2323) & (g2356) & (g2324)) + ((!g827) & (g1084) & (!g1112) & (!g2323) & (g2356) & (!g2324)) + ((!g827) & (g1084) & (!g1112) & (!g2323) & (g2356) & (g2324)) + ((!g827) & (g1084) & (!g1112) & (g2323) & (g2356) & (!g2324)) + ((!g827) & (g1084) & (!g1112) & (g2323) & (g2356) & (g2324)) + ((!g827) & (g1084) & (g1112) & (!g2323) & (g2356) & (!g2324)) + ((!g827) & (g1084) & (g1112) & (!g2323) & (g2356) & (g2324)) + ((!g827) & (g1084) & (g1112) & (g2323) & (g2356) & (!g2324)) + ((!g827) & (g1084) & (g1112) & (g2323) & (g2356) & (g2324)) + ((g827) & (!g1084) & (!g1112) & (!g2323) & (g2356) & (!g2324)) + ((g827) & (!g1084) & (!g1112) & (!g2323) & (g2356) & (g2324)) + ((g827) & (!g1084) & (!g1112) & (g2323) & (!g2356) & (g2324)) + ((g827) & (!g1084) & (!g1112) & (g2323) & (g2356) & (!g2324)) + ((g827) & (!g1084) & (g1112) & (!g2323) & (!g2356) & (!g2324)) + ((g827) & (!g1084) & (g1112) & (!g2323) & (!g2356) & (g2324)) + ((g827) & (!g1084) & (g1112) & (g2323) & (!g2356) & (!g2324)) + ((g827) & (!g1084) & (g1112) & (g2323) & (g2356) & (g2324)) + ((g827) & (g1084) & (!g1112) & (!g2323) & (!g2356) & (g2324)) + ((g827) & (g1084) & (!g1112) & (!g2323) & (g2356) & (!g2324)) + ((g827) & (g1084) & (!g1112) & (g2323) & (!g2356) & (!g2324)) + ((g827) & (g1084) & (!g1112) & (g2323) & (!g2356) & (g2324)) + ((g827) & (g1084) & (g1112) & (!g2323) & (!g2356) & (!g2324)) + ((g827) & (g1084) & (g1112) & (!g2323) & (g2356) & (g2324)) + ((g827) & (g1084) & (g1112) & (g2323) & (g2356) & (!g2324)) + ((g827) & (g1084) & (g1112) & (g2323) & (g2356) & (g2324)));
	assign g7990 = (((!g3499) & (g4615) & (!g2358)) + ((!g3499) & (g4615) & (g2358)) + ((g3499) & (!g4615) & (g2358)) + ((g3499) & (g4615) & (g2358)));
	assign g2359 = (((!g827) & (!g1092) & (!g1114) & (!g2334) & (g2358) & (!g2335)) + ((!g827) & (!g1092) & (!g1114) & (!g2334) & (g2358) & (g2335)) + ((!g827) & (!g1092) & (!g1114) & (g2334) & (g2358) & (!g2335)) + ((!g827) & (!g1092) & (!g1114) & (g2334) & (g2358) & (g2335)) + ((!g827) & (!g1092) & (g1114) & (!g2334) & (g2358) & (!g2335)) + ((!g827) & (!g1092) & (g1114) & (!g2334) & (g2358) & (g2335)) + ((!g827) & (!g1092) & (g1114) & (g2334) & (g2358) & (!g2335)) + ((!g827) & (!g1092) & (g1114) & (g2334) & (g2358) & (g2335)) + ((!g827) & (g1092) & (!g1114) & (!g2334) & (g2358) & (!g2335)) + ((!g827) & (g1092) & (!g1114) & (!g2334) & (g2358) & (g2335)) + ((!g827) & (g1092) & (!g1114) & (g2334) & (g2358) & (!g2335)) + ((!g827) & (g1092) & (!g1114) & (g2334) & (g2358) & (g2335)) + ((!g827) & (g1092) & (g1114) & (!g2334) & (g2358) & (!g2335)) + ((!g827) & (g1092) & (g1114) & (!g2334) & (g2358) & (g2335)) + ((!g827) & (g1092) & (g1114) & (g2334) & (g2358) & (!g2335)) + ((!g827) & (g1092) & (g1114) & (g2334) & (g2358) & (g2335)) + ((g827) & (!g1092) & (!g1114) & (!g2334) & (g2358) & (!g2335)) + ((g827) & (!g1092) & (!g1114) & (!g2334) & (g2358) & (g2335)) + ((g827) & (!g1092) & (!g1114) & (g2334) & (!g2358) & (g2335)) + ((g827) & (!g1092) & (!g1114) & (g2334) & (g2358) & (!g2335)) + ((g827) & (!g1092) & (g1114) & (!g2334) & (!g2358) & (!g2335)) + ((g827) & (!g1092) & (g1114) & (!g2334) & (!g2358) & (g2335)) + ((g827) & (!g1092) & (g1114) & (g2334) & (!g2358) & (!g2335)) + ((g827) & (!g1092) & (g1114) & (g2334) & (g2358) & (g2335)) + ((g827) & (g1092) & (!g1114) & (!g2334) & (!g2358) & (g2335)) + ((g827) & (g1092) & (!g1114) & (!g2334) & (g2358) & (!g2335)) + ((g827) & (g1092) & (!g1114) & (g2334) & (!g2358) & (!g2335)) + ((g827) & (g1092) & (!g1114) & (g2334) & (!g2358) & (g2335)) + ((g827) & (g1092) & (g1114) & (!g2334) & (!g2358) & (!g2335)) + ((g827) & (g1092) & (g1114) & (!g2334) & (g2358) & (g2335)) + ((g827) & (g1092) & (g1114) & (g2334) & (g2358) & (!g2335)) + ((g827) & (g1092) & (g1114) & (g2334) & (g2358) & (g2335)));
	assign g7991 = (((!g3464) & (g4619) & (!g2360)) + ((!g3464) & (g4619) & (g2360)) + ((g3464) & (!g4619) & (g2360)) + ((g3464) & (g4619) & (g2360)));
	assign g2361 = (((!g827) & (!g1070) & (!g1116) & (!g2304) & (g2360) & (!g2305)) + ((!g827) & (!g1070) & (!g1116) & (!g2304) & (g2360) & (g2305)) + ((!g827) & (!g1070) & (!g1116) & (g2304) & (g2360) & (!g2305)) + ((!g827) & (!g1070) & (!g1116) & (g2304) & (g2360) & (g2305)) + ((!g827) & (!g1070) & (g1116) & (!g2304) & (g2360) & (!g2305)) + ((!g827) & (!g1070) & (g1116) & (!g2304) & (g2360) & (g2305)) + ((!g827) & (!g1070) & (g1116) & (g2304) & (g2360) & (!g2305)) + ((!g827) & (!g1070) & (g1116) & (g2304) & (g2360) & (g2305)) + ((!g827) & (g1070) & (!g1116) & (!g2304) & (g2360) & (!g2305)) + ((!g827) & (g1070) & (!g1116) & (!g2304) & (g2360) & (g2305)) + ((!g827) & (g1070) & (!g1116) & (g2304) & (g2360) & (!g2305)) + ((!g827) & (g1070) & (!g1116) & (g2304) & (g2360) & (g2305)) + ((!g827) & (g1070) & (g1116) & (!g2304) & (g2360) & (!g2305)) + ((!g827) & (g1070) & (g1116) & (!g2304) & (g2360) & (g2305)) + ((!g827) & (g1070) & (g1116) & (g2304) & (g2360) & (!g2305)) + ((!g827) & (g1070) & (g1116) & (g2304) & (g2360) & (g2305)) + ((g827) & (!g1070) & (!g1116) & (!g2304) & (g2360) & (!g2305)) + ((g827) & (!g1070) & (!g1116) & (!g2304) & (g2360) & (g2305)) + ((g827) & (!g1070) & (!g1116) & (g2304) & (!g2360) & (g2305)) + ((g827) & (!g1070) & (!g1116) & (g2304) & (g2360) & (!g2305)) + ((g827) & (!g1070) & (g1116) & (!g2304) & (!g2360) & (!g2305)) + ((g827) & (!g1070) & (g1116) & (!g2304) & (!g2360) & (g2305)) + ((g827) & (!g1070) & (g1116) & (g2304) & (!g2360) & (!g2305)) + ((g827) & (!g1070) & (g1116) & (g2304) & (g2360) & (g2305)) + ((g827) & (g1070) & (!g1116) & (!g2304) & (!g2360) & (g2305)) + ((g827) & (g1070) & (!g1116) & (!g2304) & (g2360) & (!g2305)) + ((g827) & (g1070) & (!g1116) & (g2304) & (!g2360) & (!g2305)) + ((g827) & (g1070) & (!g1116) & (g2304) & (!g2360) & (g2305)) + ((g827) & (g1070) & (g1116) & (!g2304) & (!g2360) & (!g2305)) + ((g827) & (g1070) & (g1116) & (!g2304) & (g2360) & (g2305)) + ((g827) & (g1070) & (g1116) & (g2304) & (g2360) & (!g2305)) + ((g827) & (g1070) & (g1116) & (g2304) & (g2360) & (g2305)));
	assign g7992 = (((!g3499) & (g4623) & (!g2362)) + ((!g3499) & (g4623) & (g2362)) + ((g3499) & (!g4623) & (g2362)) + ((g3499) & (g4623) & (g2362)));
	assign g2363 = (((!g827) & (!g1078) & (!g1118) & (!g2314) & (g2362) & (!g2315)) + ((!g827) & (!g1078) & (!g1118) & (!g2314) & (g2362) & (g2315)) + ((!g827) & (!g1078) & (!g1118) & (g2314) & (g2362) & (!g2315)) + ((!g827) & (!g1078) & (!g1118) & (g2314) & (g2362) & (g2315)) + ((!g827) & (!g1078) & (g1118) & (!g2314) & (g2362) & (!g2315)) + ((!g827) & (!g1078) & (g1118) & (!g2314) & (g2362) & (g2315)) + ((!g827) & (!g1078) & (g1118) & (g2314) & (g2362) & (!g2315)) + ((!g827) & (!g1078) & (g1118) & (g2314) & (g2362) & (g2315)) + ((!g827) & (g1078) & (!g1118) & (!g2314) & (g2362) & (!g2315)) + ((!g827) & (g1078) & (!g1118) & (!g2314) & (g2362) & (g2315)) + ((!g827) & (g1078) & (!g1118) & (g2314) & (g2362) & (!g2315)) + ((!g827) & (g1078) & (!g1118) & (g2314) & (g2362) & (g2315)) + ((!g827) & (g1078) & (g1118) & (!g2314) & (g2362) & (!g2315)) + ((!g827) & (g1078) & (g1118) & (!g2314) & (g2362) & (g2315)) + ((!g827) & (g1078) & (g1118) & (g2314) & (g2362) & (!g2315)) + ((!g827) & (g1078) & (g1118) & (g2314) & (g2362) & (g2315)) + ((g827) & (!g1078) & (!g1118) & (!g2314) & (g2362) & (!g2315)) + ((g827) & (!g1078) & (!g1118) & (!g2314) & (g2362) & (g2315)) + ((g827) & (!g1078) & (!g1118) & (g2314) & (!g2362) & (g2315)) + ((g827) & (!g1078) & (!g1118) & (g2314) & (g2362) & (!g2315)) + ((g827) & (!g1078) & (g1118) & (!g2314) & (!g2362) & (!g2315)) + ((g827) & (!g1078) & (g1118) & (!g2314) & (!g2362) & (g2315)) + ((g827) & (!g1078) & (g1118) & (g2314) & (!g2362) & (!g2315)) + ((g827) & (!g1078) & (g1118) & (g2314) & (g2362) & (g2315)) + ((g827) & (g1078) & (!g1118) & (!g2314) & (!g2362) & (g2315)) + ((g827) & (g1078) & (!g1118) & (!g2314) & (g2362) & (!g2315)) + ((g827) & (g1078) & (!g1118) & (g2314) & (!g2362) & (!g2315)) + ((g827) & (g1078) & (!g1118) & (g2314) & (!g2362) & (g2315)) + ((g827) & (g1078) & (g1118) & (!g2314) & (!g2362) & (!g2315)) + ((g827) & (g1078) & (g1118) & (!g2314) & (g2362) & (g2315)) + ((g827) & (g1078) & (g1118) & (g2314) & (g2362) & (!g2315)) + ((g827) & (g1078) & (g1118) & (g2314) & (g2362) & (g2315)));
	assign g7993 = (((!g2017) & (g6604) & (!g2364)) + ((!g2017) & (g6604) & (g2364)) + ((g2017) & (!g6604) & (g2364)) + ((g2017) & (g6604) & (g2364)));
	assign g2365 = (((!g827) & (!g1086) & (!g1120) & (!g2326) & (g2364) & (!g2327)) + ((!g827) & (!g1086) & (!g1120) & (!g2326) & (g2364) & (g2327)) + ((!g827) & (!g1086) & (!g1120) & (g2326) & (g2364) & (!g2327)) + ((!g827) & (!g1086) & (!g1120) & (g2326) & (g2364) & (g2327)) + ((!g827) & (!g1086) & (g1120) & (!g2326) & (g2364) & (!g2327)) + ((!g827) & (!g1086) & (g1120) & (!g2326) & (g2364) & (g2327)) + ((!g827) & (!g1086) & (g1120) & (g2326) & (g2364) & (!g2327)) + ((!g827) & (!g1086) & (g1120) & (g2326) & (g2364) & (g2327)) + ((!g827) & (g1086) & (!g1120) & (!g2326) & (g2364) & (!g2327)) + ((!g827) & (g1086) & (!g1120) & (!g2326) & (g2364) & (g2327)) + ((!g827) & (g1086) & (!g1120) & (g2326) & (g2364) & (!g2327)) + ((!g827) & (g1086) & (!g1120) & (g2326) & (g2364) & (g2327)) + ((!g827) & (g1086) & (g1120) & (!g2326) & (g2364) & (!g2327)) + ((!g827) & (g1086) & (g1120) & (!g2326) & (g2364) & (g2327)) + ((!g827) & (g1086) & (g1120) & (g2326) & (g2364) & (!g2327)) + ((!g827) & (g1086) & (g1120) & (g2326) & (g2364) & (g2327)) + ((g827) & (!g1086) & (!g1120) & (!g2326) & (g2364) & (!g2327)) + ((g827) & (!g1086) & (!g1120) & (!g2326) & (g2364) & (g2327)) + ((g827) & (!g1086) & (!g1120) & (g2326) & (!g2364) & (g2327)) + ((g827) & (!g1086) & (!g1120) & (g2326) & (g2364) & (!g2327)) + ((g827) & (!g1086) & (g1120) & (!g2326) & (!g2364) & (!g2327)) + ((g827) & (!g1086) & (g1120) & (!g2326) & (!g2364) & (g2327)) + ((g827) & (!g1086) & (g1120) & (g2326) & (!g2364) & (!g2327)) + ((g827) & (!g1086) & (g1120) & (g2326) & (g2364) & (g2327)) + ((g827) & (g1086) & (!g1120) & (!g2326) & (!g2364) & (g2327)) + ((g827) & (g1086) & (!g1120) & (!g2326) & (g2364) & (!g2327)) + ((g827) & (g1086) & (!g1120) & (g2326) & (!g2364) & (!g2327)) + ((g827) & (g1086) & (!g1120) & (g2326) & (!g2364) & (g2327)) + ((g827) & (g1086) & (g1120) & (!g2326) & (!g2364) & (!g2327)) + ((g827) & (g1086) & (g1120) & (!g2326) & (g2364) & (g2327)) + ((g827) & (g1086) & (g1120) & (g2326) & (g2364) & (!g2327)) + ((g827) & (g1086) & (g1120) & (g2326) & (g2364) & (g2327)));
	assign g7994 = (((!g3429) & (g4627) & (!g2366)) + ((!g3429) & (g4627) & (g2366)) + ((g3429) & (!g4627) & (g2366)) + ((g3429) & (g4627) & (g2366)));
	assign g2367 = (((!g827) & (!g1094) & (!g1122) & (!g2337) & (g2366) & (!g2338)) + ((!g827) & (!g1094) & (!g1122) & (!g2337) & (g2366) & (g2338)) + ((!g827) & (!g1094) & (!g1122) & (g2337) & (g2366) & (!g2338)) + ((!g827) & (!g1094) & (!g1122) & (g2337) & (g2366) & (g2338)) + ((!g827) & (!g1094) & (g1122) & (!g2337) & (g2366) & (!g2338)) + ((!g827) & (!g1094) & (g1122) & (!g2337) & (g2366) & (g2338)) + ((!g827) & (!g1094) & (g1122) & (g2337) & (g2366) & (!g2338)) + ((!g827) & (!g1094) & (g1122) & (g2337) & (g2366) & (g2338)) + ((!g827) & (g1094) & (!g1122) & (!g2337) & (g2366) & (!g2338)) + ((!g827) & (g1094) & (!g1122) & (!g2337) & (g2366) & (g2338)) + ((!g827) & (g1094) & (!g1122) & (g2337) & (g2366) & (!g2338)) + ((!g827) & (g1094) & (!g1122) & (g2337) & (g2366) & (g2338)) + ((!g827) & (g1094) & (g1122) & (!g2337) & (g2366) & (!g2338)) + ((!g827) & (g1094) & (g1122) & (!g2337) & (g2366) & (g2338)) + ((!g827) & (g1094) & (g1122) & (g2337) & (g2366) & (!g2338)) + ((!g827) & (g1094) & (g1122) & (g2337) & (g2366) & (g2338)) + ((g827) & (!g1094) & (!g1122) & (!g2337) & (g2366) & (!g2338)) + ((g827) & (!g1094) & (!g1122) & (!g2337) & (g2366) & (g2338)) + ((g827) & (!g1094) & (!g1122) & (g2337) & (!g2366) & (g2338)) + ((g827) & (!g1094) & (!g1122) & (g2337) & (g2366) & (!g2338)) + ((g827) & (!g1094) & (g1122) & (!g2337) & (!g2366) & (!g2338)) + ((g827) & (!g1094) & (g1122) & (!g2337) & (!g2366) & (g2338)) + ((g827) & (!g1094) & (g1122) & (g2337) & (!g2366) & (!g2338)) + ((g827) & (!g1094) & (g1122) & (g2337) & (g2366) & (g2338)) + ((g827) & (g1094) & (!g1122) & (!g2337) & (!g2366) & (g2338)) + ((g827) & (g1094) & (!g1122) & (!g2337) & (g2366) & (!g2338)) + ((g827) & (g1094) & (!g1122) & (g2337) & (!g2366) & (!g2338)) + ((g827) & (g1094) & (!g1122) & (g2337) & (!g2366) & (g2338)) + ((g827) & (g1094) & (g1122) & (!g2337) & (!g2366) & (!g2338)) + ((g827) & (g1094) & (g1122) & (!g2337) & (g2366) & (g2338)) + ((g827) & (g1094) & (g1122) & (g2337) & (g2366) & (!g2338)) + ((g827) & (g1094) & (g1122) & (g2337) & (g2366) & (g2338)));
	assign g2368 = (((!g827) & (!g1072) & (!g1124) & (!g1997) & (g1999) & (!g2307)) + ((!g827) & (!g1072) & (!g1124) & (!g1997) & (g1999) & (g2307)) + ((!g827) & (!g1072) & (!g1124) & (g1997) & (g1999) & (!g2307)) + ((!g827) & (!g1072) & (!g1124) & (g1997) & (g1999) & (g2307)) + ((!g827) & (!g1072) & (g1124) & (!g1997) & (g1999) & (!g2307)) + ((!g827) & (!g1072) & (g1124) & (!g1997) & (g1999) & (g2307)) + ((!g827) & (!g1072) & (g1124) & (g1997) & (g1999) & (!g2307)) + ((!g827) & (!g1072) & (g1124) & (g1997) & (g1999) & (g2307)) + ((!g827) & (g1072) & (!g1124) & (!g1997) & (g1999) & (!g2307)) + ((!g827) & (g1072) & (!g1124) & (!g1997) & (g1999) & (g2307)) + ((!g827) & (g1072) & (!g1124) & (g1997) & (g1999) & (!g2307)) + ((!g827) & (g1072) & (!g1124) & (g1997) & (g1999) & (g2307)) + ((!g827) & (g1072) & (g1124) & (!g1997) & (g1999) & (!g2307)) + ((!g827) & (g1072) & (g1124) & (!g1997) & (g1999) & (g2307)) + ((!g827) & (g1072) & (g1124) & (g1997) & (g1999) & (!g2307)) + ((!g827) & (g1072) & (g1124) & (g1997) & (g1999) & (g2307)) + ((g827) & (!g1072) & (!g1124) & (!g1997) & (g1999) & (!g2307)) + ((g827) & (!g1072) & (!g1124) & (!g1997) & (g1999) & (g2307)) + ((g827) & (!g1072) & (!g1124) & (g1997) & (!g1999) & (g2307)) + ((g827) & (!g1072) & (!g1124) & (g1997) & (g1999) & (!g2307)) + ((g827) & (!g1072) & (g1124) & (!g1997) & (!g1999) & (!g2307)) + ((g827) & (!g1072) & (g1124) & (!g1997) & (!g1999) & (g2307)) + ((g827) & (!g1072) & (g1124) & (g1997) & (!g1999) & (!g2307)) + ((g827) & (!g1072) & (g1124) & (g1997) & (g1999) & (g2307)) + ((g827) & (g1072) & (!g1124) & (!g1997) & (!g1999) & (g2307)) + ((g827) & (g1072) & (!g1124) & (!g1997) & (g1999) & (!g2307)) + ((g827) & (g1072) & (!g1124) & (g1997) & (!g1999) & (!g2307)) + ((g827) & (g1072) & (!g1124) & (g1997) & (!g1999) & (g2307)) + ((g827) & (g1072) & (g1124) & (!g1997) & (!g1999) & (!g2307)) + ((g827) & (g1072) & (g1124) & (!g1997) & (g1999) & (g2307)) + ((g827) & (g1072) & (g1124) & (g1997) & (g1999) & (!g2307)) + ((g827) & (g1072) & (g1124) & (g1997) & (g1999) & (g2307)));
	assign g7995 = (((!g3464) & (g4631) & (!g2369)) + ((!g3464) & (g4631) & (g2369)) + ((g3464) & (!g4631) & (g2369)) + ((g3464) & (g4631) & (g2369)));
	assign g2370 = (((!g827) & (!g1080) & (!g1126) & (!g2317) & (g2369) & (!g2318)) + ((!g827) & (!g1080) & (!g1126) & (!g2317) & (g2369) & (g2318)) + ((!g827) & (!g1080) & (!g1126) & (g2317) & (g2369) & (!g2318)) + ((!g827) & (!g1080) & (!g1126) & (g2317) & (g2369) & (g2318)) + ((!g827) & (!g1080) & (g1126) & (!g2317) & (g2369) & (!g2318)) + ((!g827) & (!g1080) & (g1126) & (!g2317) & (g2369) & (g2318)) + ((!g827) & (!g1080) & (g1126) & (g2317) & (g2369) & (!g2318)) + ((!g827) & (!g1080) & (g1126) & (g2317) & (g2369) & (g2318)) + ((!g827) & (g1080) & (!g1126) & (!g2317) & (g2369) & (!g2318)) + ((!g827) & (g1080) & (!g1126) & (!g2317) & (g2369) & (g2318)) + ((!g827) & (g1080) & (!g1126) & (g2317) & (g2369) & (!g2318)) + ((!g827) & (g1080) & (!g1126) & (g2317) & (g2369) & (g2318)) + ((!g827) & (g1080) & (g1126) & (!g2317) & (g2369) & (!g2318)) + ((!g827) & (g1080) & (g1126) & (!g2317) & (g2369) & (g2318)) + ((!g827) & (g1080) & (g1126) & (g2317) & (g2369) & (!g2318)) + ((!g827) & (g1080) & (g1126) & (g2317) & (g2369) & (g2318)) + ((g827) & (!g1080) & (!g1126) & (!g2317) & (g2369) & (!g2318)) + ((g827) & (!g1080) & (!g1126) & (!g2317) & (g2369) & (g2318)) + ((g827) & (!g1080) & (!g1126) & (g2317) & (!g2369) & (g2318)) + ((g827) & (!g1080) & (!g1126) & (g2317) & (g2369) & (!g2318)) + ((g827) & (!g1080) & (g1126) & (!g2317) & (!g2369) & (!g2318)) + ((g827) & (!g1080) & (g1126) & (!g2317) & (!g2369) & (g2318)) + ((g827) & (!g1080) & (g1126) & (g2317) & (!g2369) & (!g2318)) + ((g827) & (!g1080) & (g1126) & (g2317) & (g2369) & (g2318)) + ((g827) & (g1080) & (!g1126) & (!g2317) & (!g2369) & (g2318)) + ((g827) & (g1080) & (!g1126) & (!g2317) & (g2369) & (!g2318)) + ((g827) & (g1080) & (!g1126) & (g2317) & (!g2369) & (!g2318)) + ((g827) & (g1080) & (!g1126) & (g2317) & (!g2369) & (g2318)) + ((g827) & (g1080) & (g1126) & (!g2317) & (!g2369) & (!g2318)) + ((g827) & (g1080) & (g1126) & (!g2317) & (g2369) & (g2318)) + ((g827) & (g1080) & (g1126) & (g2317) & (g2369) & (!g2318)) + ((g827) & (g1080) & (g1126) & (g2317) & (g2369) & (g2318)));
	assign g7996 = (((!g3429) & (g4633) & (!g2371)) + ((!g3429) & (g4633) & (g2371)) + ((g3429) & (!g4633) & (g2371)) + ((g3429) & (g4633) & (g2371)));
	assign g2372 = (((!g827) & (!g1088) & (!g1128) & (!g2329) & (g2371) & (!g2330)) + ((!g827) & (!g1088) & (!g1128) & (!g2329) & (g2371) & (g2330)) + ((!g827) & (!g1088) & (!g1128) & (g2329) & (g2371) & (!g2330)) + ((!g827) & (!g1088) & (!g1128) & (g2329) & (g2371) & (g2330)) + ((!g827) & (!g1088) & (g1128) & (!g2329) & (g2371) & (!g2330)) + ((!g827) & (!g1088) & (g1128) & (!g2329) & (g2371) & (g2330)) + ((!g827) & (!g1088) & (g1128) & (g2329) & (g2371) & (!g2330)) + ((!g827) & (!g1088) & (g1128) & (g2329) & (g2371) & (g2330)) + ((!g827) & (g1088) & (!g1128) & (!g2329) & (g2371) & (!g2330)) + ((!g827) & (g1088) & (!g1128) & (!g2329) & (g2371) & (g2330)) + ((!g827) & (g1088) & (!g1128) & (g2329) & (g2371) & (!g2330)) + ((!g827) & (g1088) & (!g1128) & (g2329) & (g2371) & (g2330)) + ((!g827) & (g1088) & (g1128) & (!g2329) & (g2371) & (!g2330)) + ((!g827) & (g1088) & (g1128) & (!g2329) & (g2371) & (g2330)) + ((!g827) & (g1088) & (g1128) & (g2329) & (g2371) & (!g2330)) + ((!g827) & (g1088) & (g1128) & (g2329) & (g2371) & (g2330)) + ((g827) & (!g1088) & (!g1128) & (!g2329) & (g2371) & (!g2330)) + ((g827) & (!g1088) & (!g1128) & (!g2329) & (g2371) & (g2330)) + ((g827) & (!g1088) & (!g1128) & (g2329) & (!g2371) & (g2330)) + ((g827) & (!g1088) & (!g1128) & (g2329) & (g2371) & (!g2330)) + ((g827) & (!g1088) & (g1128) & (!g2329) & (!g2371) & (!g2330)) + ((g827) & (!g1088) & (g1128) & (!g2329) & (!g2371) & (g2330)) + ((g827) & (!g1088) & (g1128) & (g2329) & (!g2371) & (!g2330)) + ((g827) & (!g1088) & (g1128) & (g2329) & (g2371) & (g2330)) + ((g827) & (g1088) & (!g1128) & (!g2329) & (!g2371) & (g2330)) + ((g827) & (g1088) & (!g1128) & (!g2329) & (g2371) & (!g2330)) + ((g827) & (g1088) & (!g1128) & (g2329) & (!g2371) & (!g2330)) + ((g827) & (g1088) & (!g1128) & (g2329) & (!g2371) & (g2330)) + ((g827) & (g1088) & (g1128) & (!g2329) & (!g2371) & (!g2330)) + ((g827) & (g1088) & (g1128) & (!g2329) & (g2371) & (g2330)) + ((g827) & (g1088) & (g1128) & (g2329) & (g2371) & (!g2330)) + ((g827) & (g1088) & (g1128) & (g2329) & (g2371) & (g2330)));
	assign g7997 = (((!g2017) & (g6598) & (!g2373)) + ((!g2017) & (g6598) & (g2373)) + ((g2017) & (!g6598) & (g2373)) + ((g2017) & (g6598) & (g2373)));
	assign g2374 = (((!g827) & (!g1096) & (!g1130) & (!g2340) & (g2373) & (!g2341)) + ((!g827) & (!g1096) & (!g1130) & (!g2340) & (g2373) & (g2341)) + ((!g827) & (!g1096) & (!g1130) & (g2340) & (g2373) & (!g2341)) + ((!g827) & (!g1096) & (!g1130) & (g2340) & (g2373) & (g2341)) + ((!g827) & (!g1096) & (g1130) & (!g2340) & (g2373) & (!g2341)) + ((!g827) & (!g1096) & (g1130) & (!g2340) & (g2373) & (g2341)) + ((!g827) & (!g1096) & (g1130) & (g2340) & (g2373) & (!g2341)) + ((!g827) & (!g1096) & (g1130) & (g2340) & (g2373) & (g2341)) + ((!g827) & (g1096) & (!g1130) & (!g2340) & (g2373) & (!g2341)) + ((!g827) & (g1096) & (!g1130) & (!g2340) & (g2373) & (g2341)) + ((!g827) & (g1096) & (!g1130) & (g2340) & (g2373) & (!g2341)) + ((!g827) & (g1096) & (!g1130) & (g2340) & (g2373) & (g2341)) + ((!g827) & (g1096) & (g1130) & (!g2340) & (g2373) & (!g2341)) + ((!g827) & (g1096) & (g1130) & (!g2340) & (g2373) & (g2341)) + ((!g827) & (g1096) & (g1130) & (g2340) & (g2373) & (!g2341)) + ((!g827) & (g1096) & (g1130) & (g2340) & (g2373) & (g2341)) + ((g827) & (!g1096) & (!g1130) & (!g2340) & (g2373) & (!g2341)) + ((g827) & (!g1096) & (!g1130) & (!g2340) & (g2373) & (g2341)) + ((g827) & (!g1096) & (!g1130) & (g2340) & (!g2373) & (g2341)) + ((g827) & (!g1096) & (!g1130) & (g2340) & (g2373) & (!g2341)) + ((g827) & (!g1096) & (g1130) & (!g2340) & (!g2373) & (!g2341)) + ((g827) & (!g1096) & (g1130) & (!g2340) & (!g2373) & (g2341)) + ((g827) & (!g1096) & (g1130) & (g2340) & (!g2373) & (!g2341)) + ((g827) & (!g1096) & (g1130) & (g2340) & (g2373) & (g2341)) + ((g827) & (g1096) & (!g1130) & (!g2340) & (!g2373) & (g2341)) + ((g827) & (g1096) & (!g1130) & (!g2340) & (g2373) & (!g2341)) + ((g827) & (g1096) & (!g1130) & (g2340) & (!g2373) & (!g2341)) + ((g827) & (g1096) & (!g1130) & (g2340) & (!g2373) & (g2341)) + ((g827) & (g1096) & (g1130) & (!g2340) & (!g2373) & (!g2341)) + ((g827) & (g1096) & (g1130) & (!g2340) & (g2373) & (g2341)) + ((g827) & (g1096) & (g1130) & (g2340) & (g2373) & (!g2341)) + ((g827) & (g1096) & (g1130) & (g2340) & (g2373) & (g2341)));
	assign g2375 = (((!g2293) & (!g2294) & (!g2295) & (!g2296) & (g2343) & (g2344)) + ((!g2293) & (!g2294) & (!g2295) & (g2296) & (g2343) & (g2344)) + ((!g2293) & (!g2294) & (g2295) & (!g2296) & (g2343) & (g2344)) + ((!g2293) & (!g2294) & (g2295) & (g2296) & (!g2343) & (g2344)) + ((!g2293) & (!g2294) & (g2295) & (g2296) & (g2343) & (!g2344)) + ((!g2293) & (!g2294) & (g2295) & (g2296) & (g2343) & (g2344)) + ((!g2293) & (g2294) & (!g2295) & (!g2296) & (g2343) & (g2344)) + ((!g2293) & (g2294) & (!g2295) & (g2296) & (!g2343) & (g2344)) + ((!g2293) & (g2294) & (!g2295) & (g2296) & (g2343) & (!g2344)) + ((!g2293) & (g2294) & (!g2295) & (g2296) & (g2343) & (g2344)) + ((!g2293) & (g2294) & (g2295) & (!g2296) & (!g2343) & (g2344)) + ((!g2293) & (g2294) & (g2295) & (!g2296) & (g2343) & (!g2344)) + ((!g2293) & (g2294) & (g2295) & (!g2296) & (g2343) & (g2344)) + ((!g2293) & (g2294) & (g2295) & (g2296) & (!g2343) & (g2344)) + ((!g2293) & (g2294) & (g2295) & (g2296) & (g2343) & (!g2344)) + ((!g2293) & (g2294) & (g2295) & (g2296) & (g2343) & (g2344)) + ((g2293) & (!g2294) & (!g2295) & (!g2296) & (g2343) & (g2344)) + ((g2293) & (!g2294) & (!g2295) & (g2296) & (!g2343) & (g2344)) + ((g2293) & (!g2294) & (!g2295) & (g2296) & (g2343) & (!g2344)) + ((g2293) & (!g2294) & (!g2295) & (g2296) & (g2343) & (g2344)) + ((g2293) & (!g2294) & (g2295) & (!g2296) & (!g2343) & (g2344)) + ((g2293) & (!g2294) & (g2295) & (!g2296) & (g2343) & (!g2344)) + ((g2293) & (!g2294) & (g2295) & (!g2296) & (g2343) & (g2344)) + ((g2293) & (!g2294) & (g2295) & (g2296) & (!g2343) & (g2344)) + ((g2293) & (!g2294) & (g2295) & (g2296) & (g2343) & (!g2344)) + ((g2293) & (!g2294) & (g2295) & (g2296) & (g2343) & (g2344)) + ((g2293) & (g2294) & (!g2295) & (!g2296) & (g2343) & (g2344)) + ((g2293) & (g2294) & (!g2295) & (g2296) & (!g2343) & (g2344)) + ((g2293) & (g2294) & (!g2295) & (g2296) & (g2343) & (!g2344)) + ((g2293) & (g2294) & (!g2295) & (g2296) & (g2343) & (g2344)) + ((g2293) & (g2294) & (g2295) & (!g2296) & (!g2343) & (g2344)) + ((g2293) & (g2294) & (g2295) & (!g2296) & (g2343) & (!g2344)) + ((g2293) & (g2294) & (g2295) & (!g2296) & (g2343) & (g2344)) + ((g2293) & (g2294) & (g2295) & (g2296) & (!g2343) & (g2344)) + ((g2293) & (g2294) & (g2295) & (g2296) & (g2343) & (!g2344)) + ((g2293) & (g2294) & (g2295) & (g2296) & (g2343) & (g2344)));
	assign g7998 = (((!g3429) & (g4640) & (!g2376)) + ((!g3429) & (g4640) & (g2376)) + ((g3429) & (!g4640) & (g2376)) + ((g3429) & (g4640) & (g2376)));
	assign g7999 = (((!g3464) & (g4644) & (!g2377)) + ((!g3464) & (g4644) & (g2377)) + ((g3464) & (!g4644) & (g2377)) + ((g3464) & (g4644) & (g2377)));
	assign g8000 = (((!g3429) & (g4650) & (!g2378)) + ((!g3429) & (g4650) & (g2378)) + ((g3429) & (!g4650) & (g2378)) + ((g3429) & (g4650) & (g2378)));
	assign g8001 = (((!g3499) & (g4654) & (!g2379)) + ((!g3499) & (g4654) & (g2379)) + ((g3499) & (!g4654) & (g2379)) + ((g3499) & (g4654) & (g2379)));
	assign g2380 = (((!g2346) & (!g2347) & (!g2348) & (!g2378) & (g2379)) + ((!g2346) & (!g2347) & (!g2348) & (g2378) & (!g2379)) + ((!g2346) & (!g2347) & (g2348) & (!g2378) & (g2379)) + ((!g2346) & (!g2347) & (g2348) & (g2378) & (!g2379)) + ((!g2346) & (g2347) & (!g2348) & (!g2378) & (g2379)) + ((!g2346) & (g2347) & (!g2348) & (g2378) & (!g2379)) + ((!g2346) & (g2347) & (g2348) & (!g2378) & (!g2379)) + ((!g2346) & (g2347) & (g2348) & (g2378) & (g2379)) + ((g2346) & (!g2347) & (!g2348) & (!g2378) & (g2379)) + ((g2346) & (!g2347) & (!g2348) & (g2378) & (!g2379)) + ((g2346) & (!g2347) & (g2348) & (!g2378) & (!g2379)) + ((g2346) & (!g2347) & (g2348) & (g2378) & (g2379)) + ((g2346) & (g2347) & (!g2348) & (!g2378) & (!g2379)) + ((g2346) & (g2347) & (!g2348) & (g2378) & (g2379)) + ((g2346) & (g2347) & (g2348) & (!g2378) & (!g2379)) + ((g2346) & (g2347) & (g2348) & (g2378) & (g2379)));
	assign g2381 = (((!g1068) & (!g1108) & (g1996) & (g1998) & (g2302)) + ((!g1068) & (g1108) & (!g1996) & (g1998) & (!g2302)) + ((!g1068) & (g1108) & (!g1996) & (g1998) & (g2302)) + ((!g1068) & (g1108) & (g1996) & (!g1998) & (g2302)) + ((!g1068) & (g1108) & (g1996) & (g1998) & (!g2302)) + ((!g1068) & (g1108) & (g1996) & (g1998) & (g2302)) + ((g1068) & (!g1108) & (!g1996) & (g1998) & (g2302)) + ((g1068) & (!g1108) & (g1996) & (g1998) & (!g2302)) + ((g1068) & (!g1108) & (g1996) & (g1998) & (g2302)) + ((g1068) & (g1108) & (!g1996) & (!g1998) & (g2302)) + ((g1068) & (g1108) & (!g1996) & (g1998) & (!g2302)) + ((g1068) & (g1108) & (!g1996) & (g1998) & (g2302)) + ((g1068) & (g1108) & (g1996) & (!g1998) & (!g2302)) + ((g1068) & (g1108) & (g1996) & (!g1998) & (g2302)) + ((g1068) & (g1108) & (g1996) & (g1998) & (!g2302)) + ((g1068) & (g1108) & (g1996) & (g1998) & (g2302)));
	assign g2382 = (((!g827) & (!g1135) & (g2001) & (!g2381)) + ((!g827) & (!g1135) & (g2001) & (g2381)) + ((!g827) & (g1135) & (g2001) & (!g2381)) + ((!g827) & (g1135) & (g2001) & (g2381)) + ((g827) & (!g1135) & (!g2001) & (g2381)) + ((g827) & (!g1135) & (g2001) & (!g2381)) + ((g827) & (g1135) & (!g2001) & (!g2381)) + ((g827) & (g1135) & (g2001) & (g2381)));
	assign g8002 = (((!g3464) & (g4657) & (!g2383)) + ((!g3464) & (g4657) & (g2383)) + ((g3464) & (!g4657) & (g2383)) + ((g3464) & (g4657) & (g2383)));
	assign g2384 = (((!g1070) & (!g1116) & (g2304) & (g2360) & (g2305)) + ((!g1070) & (g1116) & (!g2304) & (g2360) & (!g2305)) + ((!g1070) & (g1116) & (!g2304) & (g2360) & (g2305)) + ((!g1070) & (g1116) & (g2304) & (!g2360) & (g2305)) + ((!g1070) & (g1116) & (g2304) & (g2360) & (!g2305)) + ((!g1070) & (g1116) & (g2304) & (g2360) & (g2305)) + ((g1070) & (!g1116) & (!g2304) & (g2360) & (g2305)) + ((g1070) & (!g1116) & (g2304) & (g2360) & (!g2305)) + ((g1070) & (!g1116) & (g2304) & (g2360) & (g2305)) + ((g1070) & (g1116) & (!g2304) & (!g2360) & (g2305)) + ((g1070) & (g1116) & (!g2304) & (g2360) & (!g2305)) + ((g1070) & (g1116) & (!g2304) & (g2360) & (g2305)) + ((g1070) & (g1116) & (g2304) & (!g2360) & (!g2305)) + ((g1070) & (g1116) & (g2304) & (!g2360) & (g2305)) + ((g1070) & (g1116) & (g2304) & (g2360) & (!g2305)) + ((g1070) & (g1116) & (g2304) & (g2360) & (g2305)));
	assign g2385 = (((!g827) & (!g1137) & (g2383) & (!g2384)) + ((!g827) & (!g1137) & (g2383) & (g2384)) + ((!g827) & (g1137) & (g2383) & (!g2384)) + ((!g827) & (g1137) & (g2383) & (g2384)) + ((g827) & (!g1137) & (!g2383) & (g2384)) + ((g827) & (!g1137) & (g2383) & (!g2384)) + ((g827) & (g1137) & (!g2383) & (!g2384)) + ((g827) & (g1137) & (g2383) & (g2384)));
	assign g2386 = (((!g1072) & (!g1124) & (g1997) & (g1999) & (g2307)) + ((!g1072) & (g1124) & (!g1997) & (g1999) & (!g2307)) + ((!g1072) & (g1124) & (!g1997) & (g1999) & (g2307)) + ((!g1072) & (g1124) & (g1997) & (!g1999) & (g2307)) + ((!g1072) & (g1124) & (g1997) & (g1999) & (!g2307)) + ((!g1072) & (g1124) & (g1997) & (g1999) & (g2307)) + ((g1072) & (!g1124) & (!g1997) & (g1999) & (g2307)) + ((g1072) & (!g1124) & (g1997) & (g1999) & (!g2307)) + ((g1072) & (!g1124) & (g1997) & (g1999) & (g2307)) + ((g1072) & (g1124) & (!g1997) & (!g1999) & (g2307)) + ((g1072) & (g1124) & (!g1997) & (g1999) & (!g2307)) + ((g1072) & (g1124) & (!g1997) & (g1999) & (g2307)) + ((g1072) & (g1124) & (g1997) & (!g1999) & (!g2307)) + ((g1072) & (g1124) & (g1997) & (!g1999) & (g2307)) + ((g1072) & (g1124) & (g1997) & (g1999) & (!g2307)) + ((g1072) & (g1124) & (g1997) & (g1999) & (g2307)));
	assign g2387 = (((!g827) & (!g1139) & (g2002) & (!g2386)) + ((!g827) & (!g1139) & (g2002) & (g2386)) + ((!g827) & (g1139) & (g2002) & (!g2386)) + ((!g827) & (g1139) & (g2002) & (g2386)) + ((g827) & (!g1139) & (!g2002) & (g2386)) + ((g827) & (!g1139) & (g2002) & (!g2386)) + ((g827) & (g1139) & (!g2002) & (!g2386)) + ((g827) & (g1139) & (g2002) & (g2386)));
	assign g2388 = (((!g1074) & (!g1102) & (g1958) & (g1960) & (g2309)) + ((!g1074) & (g1102) & (!g1958) & (g1960) & (!g2309)) + ((!g1074) & (g1102) & (!g1958) & (g1960) & (g2309)) + ((!g1074) & (g1102) & (g1958) & (!g1960) & (g2309)) + ((!g1074) & (g1102) & (g1958) & (g1960) & (!g2309)) + ((!g1074) & (g1102) & (g1958) & (g1960) & (g2309)) + ((g1074) & (!g1102) & (!g1958) & (g1960) & (g2309)) + ((g1074) & (!g1102) & (g1958) & (g1960) & (!g2309)) + ((g1074) & (!g1102) & (g1958) & (g1960) & (g2309)) + ((g1074) & (g1102) & (!g1958) & (!g1960) & (g2309)) + ((g1074) & (g1102) & (!g1958) & (g1960) & (!g2309)) + ((g1074) & (g1102) & (!g1958) & (g1960) & (g2309)) + ((g1074) & (g1102) & (g1958) & (!g1960) & (!g2309)) + ((g1074) & (g1102) & (g1958) & (!g1960) & (g2309)) + ((g1074) & (g1102) & (g1958) & (g1960) & (!g2309)) + ((g1074) & (g1102) & (g1958) & (g1960) & (g2309)));
	assign g2389 = (((!g827) & (!g1141) & (g1962) & (!g2388)) + ((!g827) & (!g1141) & (g1962) & (g2388)) + ((!g827) & (g1141) & (g1962) & (!g2388)) + ((!g827) & (g1141) & (g1962) & (g2388)) + ((g827) & (!g1141) & (!g1962) & (g2388)) + ((g827) & (!g1141) & (g1962) & (!g2388)) + ((g827) & (g1141) & (!g1962) & (!g2388)) + ((g827) & (g1141) & (g1962) & (g2388)));
	assign g8003 = (((!g2017) & (g6591) & (!g2390)) + ((!g2017) & (g6591) & (g2390)) + ((g2017) & (!g6591) & (g2390)) + ((g2017) & (g6591) & (g2390)));
	assign g2391 = (((!g1076) & (!g1110) & (g2311) & (g2354) & (g2312)) + ((!g1076) & (g1110) & (!g2311) & (g2354) & (!g2312)) + ((!g1076) & (g1110) & (!g2311) & (g2354) & (g2312)) + ((!g1076) & (g1110) & (g2311) & (!g2354) & (g2312)) + ((!g1076) & (g1110) & (g2311) & (g2354) & (!g2312)) + ((!g1076) & (g1110) & (g2311) & (g2354) & (g2312)) + ((g1076) & (!g1110) & (!g2311) & (g2354) & (g2312)) + ((g1076) & (!g1110) & (g2311) & (g2354) & (!g2312)) + ((g1076) & (!g1110) & (g2311) & (g2354) & (g2312)) + ((g1076) & (g1110) & (!g2311) & (!g2354) & (g2312)) + ((g1076) & (g1110) & (!g2311) & (g2354) & (!g2312)) + ((g1076) & (g1110) & (!g2311) & (g2354) & (g2312)) + ((g1076) & (g1110) & (g2311) & (!g2354) & (!g2312)) + ((g1076) & (g1110) & (g2311) & (!g2354) & (g2312)) + ((g1076) & (g1110) & (g2311) & (g2354) & (!g2312)) + ((g1076) & (g1110) & (g2311) & (g2354) & (g2312)));
	assign g2392 = (((!g827) & (!g1143) & (g2390) & (!g2391)) + ((!g827) & (!g1143) & (g2390) & (g2391)) + ((!g827) & (g1143) & (g2390) & (!g2391)) + ((!g827) & (g1143) & (g2390) & (g2391)) + ((g827) & (!g1143) & (!g2390) & (g2391)) + ((g827) & (!g1143) & (g2390) & (!g2391)) + ((g827) & (g1143) & (!g2390) & (!g2391)) + ((g827) & (g1143) & (g2390) & (g2391)));
	assign g8004 = (((!g3499) & (g4663) & (!g2393)) + ((!g3499) & (g4663) & (g2393)) + ((g3499) & (!g4663) & (g2393)) + ((g3499) & (g4663) & (g2393)));
	assign g2394 = (((!g1078) & (!g1118) & (g2314) & (g2362) & (g2315)) + ((!g1078) & (g1118) & (!g2314) & (g2362) & (!g2315)) + ((!g1078) & (g1118) & (!g2314) & (g2362) & (g2315)) + ((!g1078) & (g1118) & (g2314) & (!g2362) & (g2315)) + ((!g1078) & (g1118) & (g2314) & (g2362) & (!g2315)) + ((!g1078) & (g1118) & (g2314) & (g2362) & (g2315)) + ((g1078) & (!g1118) & (!g2314) & (g2362) & (g2315)) + ((g1078) & (!g1118) & (g2314) & (g2362) & (!g2315)) + ((g1078) & (!g1118) & (g2314) & (g2362) & (g2315)) + ((g1078) & (g1118) & (!g2314) & (!g2362) & (g2315)) + ((g1078) & (g1118) & (!g2314) & (g2362) & (!g2315)) + ((g1078) & (g1118) & (!g2314) & (g2362) & (g2315)) + ((g1078) & (g1118) & (g2314) & (!g2362) & (!g2315)) + ((g1078) & (g1118) & (g2314) & (!g2362) & (g2315)) + ((g1078) & (g1118) & (g2314) & (g2362) & (!g2315)) + ((g1078) & (g1118) & (g2314) & (g2362) & (g2315)));
	assign g2395 = (((!g827) & (!g1145) & (g2393) & (!g2394)) + ((!g827) & (!g1145) & (g2393) & (g2394)) + ((!g827) & (g1145) & (g2393) & (!g2394)) + ((!g827) & (g1145) & (g2393) & (g2394)) + ((g827) & (!g1145) & (!g2393) & (g2394)) + ((g827) & (!g1145) & (g2393) & (!g2394)) + ((g827) & (g1145) & (!g2393) & (!g2394)) + ((g827) & (g1145) & (g2393) & (g2394)));
	assign g8005 = (((!g3464) & (g4666) & (!g2396)) + ((!g3464) & (g4666) & (g2396)) + ((g3464) & (!g4666) & (g2396)) + ((g3464) & (g4666) & (g2396)));
	assign g2397 = (((!g1080) & (!g1126) & (g2317) & (g2369) & (g2318)) + ((!g1080) & (g1126) & (!g2317) & (g2369) & (!g2318)) + ((!g1080) & (g1126) & (!g2317) & (g2369) & (g2318)) + ((!g1080) & (g1126) & (g2317) & (!g2369) & (g2318)) + ((!g1080) & (g1126) & (g2317) & (g2369) & (!g2318)) + ((!g1080) & (g1126) & (g2317) & (g2369) & (g2318)) + ((g1080) & (!g1126) & (!g2317) & (g2369) & (g2318)) + ((g1080) & (!g1126) & (g2317) & (g2369) & (!g2318)) + ((g1080) & (!g1126) & (g2317) & (g2369) & (g2318)) + ((g1080) & (g1126) & (!g2317) & (!g2369) & (g2318)) + ((g1080) & (g1126) & (!g2317) & (g2369) & (!g2318)) + ((g1080) & (g1126) & (!g2317) & (g2369) & (g2318)) + ((g1080) & (g1126) & (g2317) & (!g2369) & (!g2318)) + ((g1080) & (g1126) & (g2317) & (!g2369) & (g2318)) + ((g1080) & (g1126) & (g2317) & (g2369) & (!g2318)) + ((g1080) & (g1126) & (g2317) & (g2369) & (g2318)));
	assign g2398 = (((!g827) & (!g1147) & (g2396) & (!g2397)) + ((!g827) & (!g1147) & (g2396) & (g2397)) + ((!g827) & (g1147) & (g2396) & (!g2397)) + ((!g827) & (g1147) & (g2396) & (g2397)) + ((g827) & (!g1147) & (!g2396) & (g2397)) + ((g827) & (!g1147) & (g2396) & (!g2397)) + ((g827) & (g1147) & (!g2396) & (!g2397)) + ((g827) & (g1147) & (g2396) & (g2397)));
	assign g8006 = (((!g3499) & (g4669) & (!g2399)) + ((!g3499) & (g4669) & (g2399)) + ((g3499) & (!g4669) & (g2399)) + ((g3499) & (g4669) & (g2399)));
	assign g2400 = (((!g1082) & (!g1104) & (g2320) & (g2350) & (g2321)) + ((!g1082) & (g1104) & (!g2320) & (g2350) & (!g2321)) + ((!g1082) & (g1104) & (!g2320) & (g2350) & (g2321)) + ((!g1082) & (g1104) & (g2320) & (!g2350) & (g2321)) + ((!g1082) & (g1104) & (g2320) & (g2350) & (!g2321)) + ((!g1082) & (g1104) & (g2320) & (g2350) & (g2321)) + ((g1082) & (!g1104) & (!g2320) & (g2350) & (g2321)) + ((g1082) & (!g1104) & (g2320) & (g2350) & (!g2321)) + ((g1082) & (!g1104) & (g2320) & (g2350) & (g2321)) + ((g1082) & (g1104) & (!g2320) & (!g2350) & (g2321)) + ((g1082) & (g1104) & (!g2320) & (g2350) & (!g2321)) + ((g1082) & (g1104) & (!g2320) & (g2350) & (g2321)) + ((g1082) & (g1104) & (g2320) & (!g2350) & (!g2321)) + ((g1082) & (g1104) & (g2320) & (!g2350) & (g2321)) + ((g1082) & (g1104) & (g2320) & (g2350) & (!g2321)) + ((g1082) & (g1104) & (g2320) & (g2350) & (g2321)));
	assign g2401 = (((!g827) & (!g1149) & (g2399) & (!g2400)) + ((!g827) & (!g1149) & (g2399) & (g2400)) + ((!g827) & (g1149) & (g2399) & (!g2400)) + ((!g827) & (g1149) & (g2399) & (g2400)) + ((g827) & (!g1149) & (!g2399) & (g2400)) + ((g827) & (!g1149) & (g2399) & (!g2400)) + ((g827) & (g1149) & (!g2399) & (!g2400)) + ((g827) & (g1149) & (g2399) & (g2400)));
	assign g8007 = (((!g3464) & (g4673) & (!g2402)) + ((!g3464) & (g4673) & (g2402)) + ((g3464) & (!g4673) & (g2402)) + ((g3464) & (g4673) & (g2402)));
	assign g2403 = (((!g1084) & (!g1112) & (g2323) & (g2356) & (g2324)) + ((!g1084) & (g1112) & (!g2323) & (g2356) & (!g2324)) + ((!g1084) & (g1112) & (!g2323) & (g2356) & (g2324)) + ((!g1084) & (g1112) & (g2323) & (!g2356) & (g2324)) + ((!g1084) & (g1112) & (g2323) & (g2356) & (!g2324)) + ((!g1084) & (g1112) & (g2323) & (g2356) & (g2324)) + ((g1084) & (!g1112) & (!g2323) & (g2356) & (g2324)) + ((g1084) & (!g1112) & (g2323) & (g2356) & (!g2324)) + ((g1084) & (!g1112) & (g2323) & (g2356) & (g2324)) + ((g1084) & (g1112) & (!g2323) & (!g2356) & (g2324)) + ((g1084) & (g1112) & (!g2323) & (g2356) & (!g2324)) + ((g1084) & (g1112) & (!g2323) & (g2356) & (g2324)) + ((g1084) & (g1112) & (g2323) & (!g2356) & (!g2324)) + ((g1084) & (g1112) & (g2323) & (!g2356) & (g2324)) + ((g1084) & (g1112) & (g2323) & (g2356) & (!g2324)) + ((g1084) & (g1112) & (g2323) & (g2356) & (g2324)));
	assign g2404 = (((!g827) & (!g1151) & (g2402) & (!g2403)) + ((!g827) & (!g1151) & (g2402) & (g2403)) + ((!g827) & (g1151) & (g2402) & (!g2403)) + ((!g827) & (g1151) & (g2402) & (g2403)) + ((g827) & (!g1151) & (!g2402) & (g2403)) + ((g827) & (!g1151) & (g2402) & (!g2403)) + ((g827) & (g1151) & (!g2402) & (!g2403)) + ((g827) & (g1151) & (g2402) & (g2403)));
	assign g8008 = (((!g2017) & (g6584) & (!g2405)) + ((!g2017) & (g6584) & (g2405)) + ((g2017) & (!g6584) & (g2405)) + ((g2017) & (g6584) & (g2405)));
	assign g2406 = (((!g1086) & (!g1120) & (g2326) & (g2364) & (g2327)) + ((!g1086) & (g1120) & (!g2326) & (g2364) & (!g2327)) + ((!g1086) & (g1120) & (!g2326) & (g2364) & (g2327)) + ((!g1086) & (g1120) & (g2326) & (!g2364) & (g2327)) + ((!g1086) & (g1120) & (g2326) & (g2364) & (!g2327)) + ((!g1086) & (g1120) & (g2326) & (g2364) & (g2327)) + ((g1086) & (!g1120) & (!g2326) & (g2364) & (g2327)) + ((g1086) & (!g1120) & (g2326) & (g2364) & (!g2327)) + ((g1086) & (!g1120) & (g2326) & (g2364) & (g2327)) + ((g1086) & (g1120) & (!g2326) & (!g2364) & (g2327)) + ((g1086) & (g1120) & (!g2326) & (g2364) & (!g2327)) + ((g1086) & (g1120) & (!g2326) & (g2364) & (g2327)) + ((g1086) & (g1120) & (g2326) & (!g2364) & (!g2327)) + ((g1086) & (g1120) & (g2326) & (!g2364) & (g2327)) + ((g1086) & (g1120) & (g2326) & (g2364) & (!g2327)) + ((g1086) & (g1120) & (g2326) & (g2364) & (g2327)));
	assign g2407 = (((!g827) & (!g1153) & (g2405) & (!g2406)) + ((!g827) & (!g1153) & (g2405) & (g2406)) + ((!g827) & (g1153) & (g2405) & (!g2406)) + ((!g827) & (g1153) & (g2405) & (g2406)) + ((g827) & (!g1153) & (!g2405) & (g2406)) + ((g827) & (!g1153) & (g2405) & (!g2406)) + ((g827) & (g1153) & (!g2405) & (!g2406)) + ((g827) & (g1153) & (g2405) & (g2406)));
	assign g8009 = (((!g3429) & (g4679) & (!g2408)) + ((!g3429) & (g4679) & (g2408)) + ((g3429) & (!g4679) & (g2408)) + ((g3429) & (g4679) & (g2408)));
	assign g2409 = (((!g1088) & (!g1128) & (g2329) & (g2371) & (g2330)) + ((!g1088) & (g1128) & (!g2329) & (g2371) & (!g2330)) + ((!g1088) & (g1128) & (!g2329) & (g2371) & (g2330)) + ((!g1088) & (g1128) & (g2329) & (!g2371) & (g2330)) + ((!g1088) & (g1128) & (g2329) & (g2371) & (!g2330)) + ((!g1088) & (g1128) & (g2329) & (g2371) & (g2330)) + ((g1088) & (!g1128) & (!g2329) & (g2371) & (g2330)) + ((g1088) & (!g1128) & (g2329) & (g2371) & (!g2330)) + ((g1088) & (!g1128) & (g2329) & (g2371) & (g2330)) + ((g1088) & (g1128) & (!g2329) & (!g2371) & (g2330)) + ((g1088) & (g1128) & (!g2329) & (g2371) & (!g2330)) + ((g1088) & (g1128) & (!g2329) & (g2371) & (g2330)) + ((g1088) & (g1128) & (g2329) & (!g2371) & (!g2330)) + ((g1088) & (g1128) & (g2329) & (!g2371) & (g2330)) + ((g1088) & (g1128) & (g2329) & (g2371) & (!g2330)) + ((g1088) & (g1128) & (g2329) & (g2371) & (g2330)));
	assign g2410 = (((!g827) & (!g1155) & (g2408) & (!g2409)) + ((!g827) & (!g1155) & (g2408) & (g2409)) + ((!g827) & (g1155) & (g2408) & (!g2409)) + ((!g827) & (g1155) & (g2408) & (g2409)) + ((g827) & (!g1155) & (!g2408) & (g2409)) + ((g827) & (!g1155) & (g2408) & (!g2409)) + ((g827) & (g1155) & (!g2408) & (!g2409)) + ((g827) & (g1155) & (g2408) & (g2409)));
	assign g2411 = (((!g1090) & (!g1106) & (g1959) & (g1961) & (g2332)) + ((!g1090) & (g1106) & (!g1959) & (g1961) & (!g2332)) + ((!g1090) & (g1106) & (!g1959) & (g1961) & (g2332)) + ((!g1090) & (g1106) & (g1959) & (!g1961) & (g2332)) + ((!g1090) & (g1106) & (g1959) & (g1961) & (!g2332)) + ((!g1090) & (g1106) & (g1959) & (g1961) & (g2332)) + ((g1090) & (!g1106) & (!g1959) & (g1961) & (g2332)) + ((g1090) & (!g1106) & (g1959) & (g1961) & (!g2332)) + ((g1090) & (!g1106) & (g1959) & (g1961) & (g2332)) + ((g1090) & (g1106) & (!g1959) & (!g1961) & (g2332)) + ((g1090) & (g1106) & (!g1959) & (g1961) & (!g2332)) + ((g1090) & (g1106) & (!g1959) & (g1961) & (g2332)) + ((g1090) & (g1106) & (g1959) & (!g1961) & (!g2332)) + ((g1090) & (g1106) & (g1959) & (!g1961) & (g2332)) + ((g1090) & (g1106) & (g1959) & (g1961) & (!g2332)) + ((g1090) & (g1106) & (g1959) & (g1961) & (g2332)));
	assign g2412 = (((!g827) & (!g1157) & (g1963) & (!g2411)) + ((!g827) & (!g1157) & (g1963) & (g2411)) + ((!g827) & (g1157) & (g1963) & (!g2411)) + ((!g827) & (g1157) & (g1963) & (g2411)) + ((g827) & (!g1157) & (!g1963) & (g2411)) + ((g827) & (!g1157) & (g1963) & (!g2411)) + ((g827) & (g1157) & (!g1963) & (!g2411)) + ((g827) & (g1157) & (g1963) & (g2411)));
	assign g8010 = (((!g3499) & (g4682) & (!g2413)) + ((!g3499) & (g4682) & (g2413)) + ((g3499) & (!g4682) & (g2413)) + ((g3499) & (g4682) & (g2413)));
	assign g2414 = (((!g1092) & (!g1114) & (g2334) & (g2358) & (g2335)) + ((!g1092) & (g1114) & (!g2334) & (g2358) & (!g2335)) + ((!g1092) & (g1114) & (!g2334) & (g2358) & (g2335)) + ((!g1092) & (g1114) & (g2334) & (!g2358) & (g2335)) + ((!g1092) & (g1114) & (g2334) & (g2358) & (!g2335)) + ((!g1092) & (g1114) & (g2334) & (g2358) & (g2335)) + ((g1092) & (!g1114) & (!g2334) & (g2358) & (g2335)) + ((g1092) & (!g1114) & (g2334) & (g2358) & (!g2335)) + ((g1092) & (!g1114) & (g2334) & (g2358) & (g2335)) + ((g1092) & (g1114) & (!g2334) & (!g2358) & (g2335)) + ((g1092) & (g1114) & (!g2334) & (g2358) & (!g2335)) + ((g1092) & (g1114) & (!g2334) & (g2358) & (g2335)) + ((g1092) & (g1114) & (g2334) & (!g2358) & (!g2335)) + ((g1092) & (g1114) & (g2334) & (!g2358) & (g2335)) + ((g1092) & (g1114) & (g2334) & (g2358) & (!g2335)) + ((g1092) & (g1114) & (g2334) & (g2358) & (g2335)));
	assign g2415 = (((!g827) & (!g1159) & (g2413) & (!g2414)) + ((!g827) & (!g1159) & (g2413) & (g2414)) + ((!g827) & (g1159) & (g2413) & (!g2414)) + ((!g827) & (g1159) & (g2413) & (g2414)) + ((g827) & (!g1159) & (!g2413) & (g2414)) + ((g827) & (!g1159) & (g2413) & (!g2414)) + ((g827) & (g1159) & (!g2413) & (!g2414)) + ((g827) & (g1159) & (g2413) & (g2414)));
	assign g8011 = (((!g3429) & (g4685) & (!g2416)) + ((!g3429) & (g4685) & (g2416)) + ((g3429) & (!g4685) & (g2416)) + ((g3429) & (g4685) & (g2416)));
	assign g2417 = (((!g1094) & (!g1122) & (g2337) & (g2366) & (g2338)) + ((!g1094) & (g1122) & (!g2337) & (g2366) & (!g2338)) + ((!g1094) & (g1122) & (!g2337) & (g2366) & (g2338)) + ((!g1094) & (g1122) & (g2337) & (!g2366) & (g2338)) + ((!g1094) & (g1122) & (g2337) & (g2366) & (!g2338)) + ((!g1094) & (g1122) & (g2337) & (g2366) & (g2338)) + ((g1094) & (!g1122) & (!g2337) & (g2366) & (g2338)) + ((g1094) & (!g1122) & (g2337) & (g2366) & (!g2338)) + ((g1094) & (!g1122) & (g2337) & (g2366) & (g2338)) + ((g1094) & (g1122) & (!g2337) & (!g2366) & (g2338)) + ((g1094) & (g1122) & (!g2337) & (g2366) & (!g2338)) + ((g1094) & (g1122) & (!g2337) & (g2366) & (g2338)) + ((g1094) & (g1122) & (g2337) & (!g2366) & (!g2338)) + ((g1094) & (g1122) & (g2337) & (!g2366) & (g2338)) + ((g1094) & (g1122) & (g2337) & (g2366) & (!g2338)) + ((g1094) & (g1122) & (g2337) & (g2366) & (g2338)));
	assign g2418 = (((!g827) & (!g1161) & (g2416) & (!g2417)) + ((!g827) & (!g1161) & (g2416) & (g2417)) + ((!g827) & (g1161) & (g2416) & (!g2417)) + ((!g827) & (g1161) & (g2416) & (g2417)) + ((g827) & (!g1161) & (!g2416) & (g2417)) + ((g827) & (!g1161) & (g2416) & (!g2417)) + ((g827) & (g1161) & (!g2416) & (!g2417)) + ((g827) & (g1161) & (g2416) & (g2417)));
	assign g8012 = (((!g2017) & (g6577) & (!g2419)) + ((!g2017) & (g6577) & (g2419)) + ((g2017) & (!g6577) & (g2419)) + ((g2017) & (g6577) & (g2419)));
	assign g2420 = (((!g1096) & (!g1130) & (g2340) & (g2373) & (g2341)) + ((!g1096) & (g1130) & (!g2340) & (g2373) & (!g2341)) + ((!g1096) & (g1130) & (!g2340) & (g2373) & (g2341)) + ((!g1096) & (g1130) & (g2340) & (!g2373) & (g2341)) + ((!g1096) & (g1130) & (g2340) & (g2373) & (!g2341)) + ((!g1096) & (g1130) & (g2340) & (g2373) & (g2341)) + ((g1096) & (!g1130) & (!g2340) & (g2373) & (g2341)) + ((g1096) & (!g1130) & (g2340) & (g2373) & (!g2341)) + ((g1096) & (!g1130) & (g2340) & (g2373) & (g2341)) + ((g1096) & (g1130) & (!g2340) & (!g2373) & (g2341)) + ((g1096) & (g1130) & (!g2340) & (g2373) & (!g2341)) + ((g1096) & (g1130) & (!g2340) & (g2373) & (g2341)) + ((g1096) & (g1130) & (g2340) & (!g2373) & (!g2341)) + ((g1096) & (g1130) & (g2340) & (!g2373) & (g2341)) + ((g1096) & (g1130) & (g2340) & (g2373) & (!g2341)) + ((g1096) & (g1130) & (g2340) & (g2373) & (g2341)));
	assign g2421 = (((!g827) & (!g1163) & (g2419) & (!g2420)) + ((!g827) & (!g1163) & (g2419) & (g2420)) + ((!g827) & (g1163) & (g2419) & (!g2420)) + ((!g827) & (g1163) & (g2419) & (g2420)) + ((g827) & (!g1163) & (!g2419) & (g2420)) + ((g827) & (!g1163) & (g2419) & (!g2420)) + ((g827) & (g1163) & (!g2419) & (!g2420)) + ((g827) & (g1163) & (g2419) & (g2420)));
	assign g2422 = (((!g2375) & (g2376) & (g2377)) + ((g2375) & (!g2376) & (g2377)) + ((g2375) & (g2376) & (!g2377)) + ((g2375) & (g2376) & (g2377)));
	assign g8013 = (((!g3429) & (g4691) & (!g2423)) + ((!g3429) & (g4691) & (g2423)) + ((g3429) & (!g4691) & (g2423)) + ((g3429) & (g4691) & (g2423)));
	assign g8014 = (((!g3464) & (g4694) & (!g2424)) + ((!g3464) & (g4694) & (g2424)) + ((g3464) & (!g4694) & (g2424)) + ((g3464) & (g4694) & (g2424)));
	assign g2425 = (((!g2346) & (!g2347) & (!g2348) & (g2378) & (g2379)) + ((!g2346) & (!g2347) & (g2348) & (g2378) & (g2379)) + ((!g2346) & (g2347) & (!g2348) & (g2378) & (g2379)) + ((!g2346) & (g2347) & (g2348) & (!g2378) & (g2379)) + ((!g2346) & (g2347) & (g2348) & (g2378) & (!g2379)) + ((!g2346) & (g2347) & (g2348) & (g2378) & (g2379)) + ((g2346) & (!g2347) & (!g2348) & (g2378) & (g2379)) + ((g2346) & (!g2347) & (g2348) & (!g2378) & (g2379)) + ((g2346) & (!g2347) & (g2348) & (g2378) & (!g2379)) + ((g2346) & (!g2347) & (g2348) & (g2378) & (g2379)) + ((g2346) & (g2347) & (!g2348) & (!g2378) & (g2379)) + ((g2346) & (g2347) & (!g2348) & (g2378) & (!g2379)) + ((g2346) & (g2347) & (!g2348) & (g2378) & (g2379)) + ((g2346) & (g2347) & (g2348) & (!g2378) & (g2379)) + ((g2346) & (g2347) & (g2348) & (g2378) & (!g2379)) + ((g2346) & (g2347) & (g2348) & (g2378) & (g2379)));
	assign g8015 = (((!g3429) & (g4697) & (!g2426)) + ((!g3429) & (g4697) & (g2426)) + ((g3429) & (!g4697) & (g2426)) + ((g3429) & (g4697) & (g2426)));
	assign g8016 = (((!g3499) & (g4700) & (!g2427)) + ((!g3499) & (g4700) & (g2427)) + ((g3499) & (!g4700) & (g2427)) + ((g3499) & (g4700) & (g2427)));
	assign g2428 = (((!g2425) & (!g2426) & (g2427)) + ((!g2425) & (g2426) & (!g2427)) + ((g2425) & (!g2426) & (!g2427)) + ((g2425) & (g2426) & (g2427)));
	assign g2429 = (((!g1141) & (g1962)) + ((g1141) & (!g1962)));
	assign g2430 = (((!g1074) & (!g1102) & (g1958) & (g1960) & (g2309) & (g2429)) + ((!g1074) & (g1102) & (!g1958) & (g1960) & (!g2309) & (g2429)) + ((!g1074) & (g1102) & (!g1958) & (g1960) & (g2309) & (g2429)) + ((!g1074) & (g1102) & (g1958) & (!g1960) & (g2309) & (g2429)) + ((!g1074) & (g1102) & (g1958) & (g1960) & (!g2309) & (g2429)) + ((!g1074) & (g1102) & (g1958) & (g1960) & (g2309) & (g2429)) + ((g1074) & (!g1102) & (!g1958) & (g1960) & (g2309) & (g2429)) + ((g1074) & (!g1102) & (g1958) & (g1960) & (!g2309) & (g2429)) + ((g1074) & (!g1102) & (g1958) & (g1960) & (g2309) & (g2429)) + ((g1074) & (g1102) & (!g1958) & (!g1960) & (g2309) & (g2429)) + ((g1074) & (g1102) & (!g1958) & (g1960) & (!g2309) & (g2429)) + ((g1074) & (g1102) & (!g1958) & (g1960) & (g2309) & (g2429)) + ((g1074) & (g1102) & (g1958) & (!g1960) & (!g2309) & (g2429)) + ((g1074) & (g1102) & (g1958) & (!g1960) & (g2309) & (g2429)) + ((g1074) & (g1102) & (g1958) & (g1960) & (!g2309) & (g2429)) + ((g1074) & (g1102) & (g1958) & (g1960) & (g2309) & (g2429)));
	assign g2431 = (((g1141) & (g1962)));
	assign g2432 = (((!g2430) & (!g2431)));
	assign g2433 = (((!g827) & (!g1169) & (g1967) & (!g2432)) + ((!g827) & (!g1169) & (g1967) & (g2432)) + ((!g827) & (g1169) & (g1967) & (!g2432)) + ((!g827) & (g1169) & (g1967) & (g2432)) + ((g827) & (!g1169) & (!g1967) & (!g2432)) + ((g827) & (!g1169) & (g1967) & (g2432)) + ((g827) & (g1169) & (!g1967) & (g2432)) + ((g827) & (g1169) & (g1967) & (!g2432)));
	assign g8017 = (((!g3499) & (g4703) & (!g2434)) + ((!g3499) & (g4703) & (g2434)) + ((g3499) & (!g4703) & (g2434)) + ((g3499) & (g4703) & (g2434)));
	assign g2435 = (((!g1149) & (g2399)) + ((g1149) & (!g2399)));
	assign g2436 = (((!g1082) & (!g1104) & (g2320) & (g2350) & (g2321) & (g2435)) + ((!g1082) & (g1104) & (!g2320) & (g2350) & (!g2321) & (g2435)) + ((!g1082) & (g1104) & (!g2320) & (g2350) & (g2321) & (g2435)) + ((!g1082) & (g1104) & (g2320) & (!g2350) & (g2321) & (g2435)) + ((!g1082) & (g1104) & (g2320) & (g2350) & (!g2321) & (g2435)) + ((!g1082) & (g1104) & (g2320) & (g2350) & (g2321) & (g2435)) + ((g1082) & (!g1104) & (!g2320) & (g2350) & (g2321) & (g2435)) + ((g1082) & (!g1104) & (g2320) & (g2350) & (!g2321) & (g2435)) + ((g1082) & (!g1104) & (g2320) & (g2350) & (g2321) & (g2435)) + ((g1082) & (g1104) & (!g2320) & (!g2350) & (g2321) & (g2435)) + ((g1082) & (g1104) & (!g2320) & (g2350) & (!g2321) & (g2435)) + ((g1082) & (g1104) & (!g2320) & (g2350) & (g2321) & (g2435)) + ((g1082) & (g1104) & (g2320) & (!g2350) & (!g2321) & (g2435)) + ((g1082) & (g1104) & (g2320) & (!g2350) & (g2321) & (g2435)) + ((g1082) & (g1104) & (g2320) & (g2350) & (!g2321) & (g2435)) + ((g1082) & (g1104) & (g2320) & (g2350) & (g2321) & (g2435)));
	assign g2437 = (((g1149) & (g2399)));
	assign g2438 = (((!g2436) & (!g2437)));
	assign g2439 = (((!g827) & (!g1171) & (g2434) & (!g2438)) + ((!g827) & (!g1171) & (g2434) & (g2438)) + ((!g827) & (g1171) & (g2434) & (!g2438)) + ((!g827) & (g1171) & (g2434) & (g2438)) + ((g827) & (!g1171) & (!g2434) & (!g2438)) + ((g827) & (!g1171) & (g2434) & (g2438)) + ((g827) & (g1171) & (!g2434) & (g2438)) + ((g827) & (g1171) & (g2434) & (!g2438)));
	assign g2440 = (((!g1157) & (g1963)) + ((g1157) & (!g1963)));
	assign g2441 = (((!g1090) & (!g1106) & (g1959) & (g1961) & (g2332) & (g2440)) + ((!g1090) & (g1106) & (!g1959) & (g1961) & (!g2332) & (g2440)) + ((!g1090) & (g1106) & (!g1959) & (g1961) & (g2332) & (g2440)) + ((!g1090) & (g1106) & (g1959) & (!g1961) & (g2332) & (g2440)) + ((!g1090) & (g1106) & (g1959) & (g1961) & (!g2332) & (g2440)) + ((!g1090) & (g1106) & (g1959) & (g1961) & (g2332) & (g2440)) + ((g1090) & (!g1106) & (!g1959) & (g1961) & (g2332) & (g2440)) + ((g1090) & (!g1106) & (g1959) & (g1961) & (!g2332) & (g2440)) + ((g1090) & (!g1106) & (g1959) & (g1961) & (g2332) & (g2440)) + ((g1090) & (g1106) & (!g1959) & (!g1961) & (g2332) & (g2440)) + ((g1090) & (g1106) & (!g1959) & (g1961) & (!g2332) & (g2440)) + ((g1090) & (g1106) & (!g1959) & (g1961) & (g2332) & (g2440)) + ((g1090) & (g1106) & (g1959) & (!g1961) & (!g2332) & (g2440)) + ((g1090) & (g1106) & (g1959) & (!g1961) & (g2332) & (g2440)) + ((g1090) & (g1106) & (g1959) & (g1961) & (!g2332) & (g2440)) + ((g1090) & (g1106) & (g1959) & (g1961) & (g2332) & (g2440)));
	assign g2442 = (((g1157) & (g1963)));
	assign g2443 = (((!g2441) & (!g2442)));
	assign g2444 = (((!g827) & (!g1173) & (g1968) & (!g2443)) + ((!g827) & (!g1173) & (g1968) & (g2443)) + ((!g827) & (g1173) & (g1968) & (!g2443)) + ((!g827) & (g1173) & (g1968) & (g2443)) + ((g827) & (!g1173) & (!g1968) & (!g2443)) + ((g827) & (!g1173) & (g1968) & (g2443)) + ((g827) & (g1173) & (!g1968) & (g2443)) + ((g827) & (g1173) & (g1968) & (!g2443)));
	assign g2445 = (((!g1135) & (g2001)) + ((g1135) & (!g2001)));
	assign g2446 = (((!g1068) & (!g1108) & (g1996) & (g1998) & (g2302) & (g2445)) + ((!g1068) & (g1108) & (!g1996) & (g1998) & (!g2302) & (g2445)) + ((!g1068) & (g1108) & (!g1996) & (g1998) & (g2302) & (g2445)) + ((!g1068) & (g1108) & (g1996) & (!g1998) & (g2302) & (g2445)) + ((!g1068) & (g1108) & (g1996) & (g1998) & (!g2302) & (g2445)) + ((!g1068) & (g1108) & (g1996) & (g1998) & (g2302) & (g2445)) + ((g1068) & (!g1108) & (!g1996) & (g1998) & (g2302) & (g2445)) + ((g1068) & (!g1108) & (g1996) & (g1998) & (!g2302) & (g2445)) + ((g1068) & (!g1108) & (g1996) & (g1998) & (g2302) & (g2445)) + ((g1068) & (g1108) & (!g1996) & (!g1998) & (g2302) & (g2445)) + ((g1068) & (g1108) & (!g1996) & (g1998) & (!g2302) & (g2445)) + ((g1068) & (g1108) & (!g1996) & (g1998) & (g2302) & (g2445)) + ((g1068) & (g1108) & (g1996) & (!g1998) & (!g2302) & (g2445)) + ((g1068) & (g1108) & (g1996) & (!g1998) & (g2302) & (g2445)) + ((g1068) & (g1108) & (g1996) & (g1998) & (!g2302) & (g2445)) + ((g1068) & (g1108) & (g1996) & (g1998) & (g2302) & (g2445)));
	assign g2447 = (((g1135) & (g2001)));
	assign g2448 = (((!g2446) & (!g2447)));
	assign g2449 = (((!g827) & (!g1175) & (g2003) & (!g2448)) + ((!g827) & (!g1175) & (g2003) & (g2448)) + ((!g827) & (g1175) & (g2003) & (!g2448)) + ((!g827) & (g1175) & (g2003) & (g2448)) + ((g827) & (!g1175) & (!g2003) & (!g2448)) + ((g827) & (!g1175) & (g2003) & (g2448)) + ((g827) & (g1175) & (!g2003) & (g2448)) + ((g827) & (g1175) & (g2003) & (!g2448)));
	assign g8018 = (((!g2017) & (g4706) & (!g2450)) + ((!g2017) & (g4706) & (g2450)) + ((g2017) & (!g4706) & (g2450)) + ((g2017) & (g4706) & (g2450)));
	assign g2451 = (((!g1143) & (g2390)) + ((g1143) & (!g2390)));
	assign g2452 = (((!g1076) & (!g1110) & (g2311) & (g2354) & (g2312) & (g2451)) + ((!g1076) & (g1110) & (!g2311) & (g2354) & (!g2312) & (g2451)) + ((!g1076) & (g1110) & (!g2311) & (g2354) & (g2312) & (g2451)) + ((!g1076) & (g1110) & (g2311) & (!g2354) & (g2312) & (g2451)) + ((!g1076) & (g1110) & (g2311) & (g2354) & (!g2312) & (g2451)) + ((!g1076) & (g1110) & (g2311) & (g2354) & (g2312) & (g2451)) + ((g1076) & (!g1110) & (!g2311) & (g2354) & (g2312) & (g2451)) + ((g1076) & (!g1110) & (g2311) & (g2354) & (!g2312) & (g2451)) + ((g1076) & (!g1110) & (g2311) & (g2354) & (g2312) & (g2451)) + ((g1076) & (g1110) & (!g2311) & (!g2354) & (g2312) & (g2451)) + ((g1076) & (g1110) & (!g2311) & (g2354) & (!g2312) & (g2451)) + ((g1076) & (g1110) & (!g2311) & (g2354) & (g2312) & (g2451)) + ((g1076) & (g1110) & (g2311) & (!g2354) & (!g2312) & (g2451)) + ((g1076) & (g1110) & (g2311) & (!g2354) & (g2312) & (g2451)) + ((g1076) & (g1110) & (g2311) & (g2354) & (!g2312) & (g2451)) + ((g1076) & (g1110) & (g2311) & (g2354) & (g2312) & (g2451)));
	assign g2453 = (((g1143) & (g2390)));
	assign g2454 = (((!g2452) & (!g2453)));
	assign g2455 = (((!g827) & (!g1177) & (g2450) & (!g2454)) + ((!g827) & (!g1177) & (g2450) & (g2454)) + ((!g827) & (g1177) & (g2450) & (!g2454)) + ((!g827) & (g1177) & (g2450) & (g2454)) + ((g827) & (!g1177) & (!g2450) & (!g2454)) + ((g827) & (!g1177) & (g2450) & (g2454)) + ((g827) & (g1177) & (!g2450) & (g2454)) + ((g827) & (g1177) & (g2450) & (!g2454)));
	assign g8019 = (((!g3464) & (g4710) & (!g2456)) + ((!g3464) & (g4710) & (g2456)) + ((g3464) & (!g4710) & (g2456)) + ((g3464) & (g4710) & (g2456)));
	assign g2457 = (((!g1151) & (g2402)) + ((g1151) & (!g2402)));
	assign g2458 = (((!g1084) & (!g1112) & (g2323) & (g2356) & (g2324) & (g2457)) + ((!g1084) & (g1112) & (!g2323) & (g2356) & (!g2324) & (g2457)) + ((!g1084) & (g1112) & (!g2323) & (g2356) & (g2324) & (g2457)) + ((!g1084) & (g1112) & (g2323) & (!g2356) & (g2324) & (g2457)) + ((!g1084) & (g1112) & (g2323) & (g2356) & (!g2324) & (g2457)) + ((!g1084) & (g1112) & (g2323) & (g2356) & (g2324) & (g2457)) + ((g1084) & (!g1112) & (!g2323) & (g2356) & (g2324) & (g2457)) + ((g1084) & (!g1112) & (g2323) & (g2356) & (!g2324) & (g2457)) + ((g1084) & (!g1112) & (g2323) & (g2356) & (g2324) & (g2457)) + ((g1084) & (g1112) & (!g2323) & (!g2356) & (g2324) & (g2457)) + ((g1084) & (g1112) & (!g2323) & (g2356) & (!g2324) & (g2457)) + ((g1084) & (g1112) & (!g2323) & (g2356) & (g2324) & (g2457)) + ((g1084) & (g1112) & (g2323) & (!g2356) & (!g2324) & (g2457)) + ((g1084) & (g1112) & (g2323) & (!g2356) & (g2324) & (g2457)) + ((g1084) & (g1112) & (g2323) & (g2356) & (!g2324) & (g2457)) + ((g1084) & (g1112) & (g2323) & (g2356) & (g2324) & (g2457)));
	assign g2459 = (((g1151) & (g2402)));
	assign g2460 = (((!g2458) & (!g2459)));
	assign g2461 = (((!g827) & (!g1179) & (g2456) & (!g2460)) + ((!g827) & (!g1179) & (g2456) & (g2460)) + ((!g827) & (g1179) & (g2456) & (!g2460)) + ((!g827) & (g1179) & (g2456) & (g2460)) + ((g827) & (!g1179) & (!g2456) & (!g2460)) + ((g827) & (!g1179) & (g2456) & (g2460)) + ((g827) & (g1179) & (!g2456) & (g2460)) + ((g827) & (g1179) & (g2456) & (!g2460)));
	assign g8020 = (((!g3499) & (g4713) & (!g2462)) + ((!g3499) & (g4713) & (g2462)) + ((g3499) & (!g4713) & (g2462)) + ((g3499) & (g4713) & (g2462)));
	assign g2463 = (((!g1159) & (g2413)) + ((g1159) & (!g2413)));
	assign g2464 = (((!g1092) & (!g1114) & (g2334) & (g2358) & (g2335) & (g2463)) + ((!g1092) & (g1114) & (!g2334) & (g2358) & (!g2335) & (g2463)) + ((!g1092) & (g1114) & (!g2334) & (g2358) & (g2335) & (g2463)) + ((!g1092) & (g1114) & (g2334) & (!g2358) & (g2335) & (g2463)) + ((!g1092) & (g1114) & (g2334) & (g2358) & (!g2335) & (g2463)) + ((!g1092) & (g1114) & (g2334) & (g2358) & (g2335) & (g2463)) + ((g1092) & (!g1114) & (!g2334) & (g2358) & (g2335) & (g2463)) + ((g1092) & (!g1114) & (g2334) & (g2358) & (!g2335) & (g2463)) + ((g1092) & (!g1114) & (g2334) & (g2358) & (g2335) & (g2463)) + ((g1092) & (g1114) & (!g2334) & (!g2358) & (g2335) & (g2463)) + ((g1092) & (g1114) & (!g2334) & (g2358) & (!g2335) & (g2463)) + ((g1092) & (g1114) & (!g2334) & (g2358) & (g2335) & (g2463)) + ((g1092) & (g1114) & (g2334) & (!g2358) & (!g2335) & (g2463)) + ((g1092) & (g1114) & (g2334) & (!g2358) & (g2335) & (g2463)) + ((g1092) & (g1114) & (g2334) & (g2358) & (!g2335) & (g2463)) + ((g1092) & (g1114) & (g2334) & (g2358) & (g2335) & (g2463)));
	assign g2465 = (((g1159) & (g2413)));
	assign g2466 = (((!g2464) & (!g2465)));
	assign g2467 = (((!g827) & (!g1181) & (g2462) & (!g2466)) + ((!g827) & (!g1181) & (g2462) & (g2466)) + ((!g827) & (g1181) & (g2462) & (!g2466)) + ((!g827) & (g1181) & (g2462) & (g2466)) + ((g827) & (!g1181) & (!g2462) & (!g2466)) + ((g827) & (!g1181) & (g2462) & (g2466)) + ((g827) & (g1181) & (!g2462) & (g2466)) + ((g827) & (g1181) & (g2462) & (!g2466)));
	assign g8021 = (((!g3464) & (g4716) & (!g2468)) + ((!g3464) & (g4716) & (g2468)) + ((g3464) & (!g4716) & (g2468)) + ((g3464) & (g4716) & (g2468)));
	assign g2469 = (((!g1137) & (g2383)) + ((g1137) & (!g2383)));
	assign g2470 = (((!g1070) & (!g1116) & (g2304) & (g2360) & (g2305) & (g2469)) + ((!g1070) & (g1116) & (!g2304) & (g2360) & (!g2305) & (g2469)) + ((!g1070) & (g1116) & (!g2304) & (g2360) & (g2305) & (g2469)) + ((!g1070) & (g1116) & (g2304) & (!g2360) & (g2305) & (g2469)) + ((!g1070) & (g1116) & (g2304) & (g2360) & (!g2305) & (g2469)) + ((!g1070) & (g1116) & (g2304) & (g2360) & (g2305) & (g2469)) + ((g1070) & (!g1116) & (!g2304) & (g2360) & (g2305) & (g2469)) + ((g1070) & (!g1116) & (g2304) & (g2360) & (!g2305) & (g2469)) + ((g1070) & (!g1116) & (g2304) & (g2360) & (g2305) & (g2469)) + ((g1070) & (g1116) & (!g2304) & (!g2360) & (g2305) & (g2469)) + ((g1070) & (g1116) & (!g2304) & (g2360) & (!g2305) & (g2469)) + ((g1070) & (g1116) & (!g2304) & (g2360) & (g2305) & (g2469)) + ((g1070) & (g1116) & (g2304) & (!g2360) & (!g2305) & (g2469)) + ((g1070) & (g1116) & (g2304) & (!g2360) & (g2305) & (g2469)) + ((g1070) & (g1116) & (g2304) & (g2360) & (!g2305) & (g2469)) + ((g1070) & (g1116) & (g2304) & (g2360) & (g2305) & (g2469)));
	assign g2471 = (((g1137) & (g2383)));
	assign g2472 = (((!g2470) & (!g2471)));
	assign g2473 = (((!g827) & (!g1183) & (g2468) & (!g2472)) + ((!g827) & (!g1183) & (g2468) & (g2472)) + ((!g827) & (g1183) & (g2468) & (!g2472)) + ((!g827) & (g1183) & (g2468) & (g2472)) + ((g827) & (!g1183) & (!g2468) & (!g2472)) + ((g827) & (!g1183) & (g2468) & (g2472)) + ((g827) & (g1183) & (!g2468) & (g2472)) + ((g827) & (g1183) & (g2468) & (!g2472)));
	assign g8022 = (((!g3499) & (g4719) & (!g2474)) + ((!g3499) & (g4719) & (g2474)) + ((g3499) & (!g4719) & (g2474)) + ((g3499) & (g4719) & (g2474)));
	assign g2475 = (((!g1145) & (g2393)) + ((g1145) & (!g2393)));
	assign g2476 = (((!g1078) & (!g1118) & (g2314) & (g2362) & (g2315) & (g2475)) + ((!g1078) & (g1118) & (!g2314) & (g2362) & (!g2315) & (g2475)) + ((!g1078) & (g1118) & (!g2314) & (g2362) & (g2315) & (g2475)) + ((!g1078) & (g1118) & (g2314) & (!g2362) & (g2315) & (g2475)) + ((!g1078) & (g1118) & (g2314) & (g2362) & (!g2315) & (g2475)) + ((!g1078) & (g1118) & (g2314) & (g2362) & (g2315) & (g2475)) + ((g1078) & (!g1118) & (!g2314) & (g2362) & (g2315) & (g2475)) + ((g1078) & (!g1118) & (g2314) & (g2362) & (!g2315) & (g2475)) + ((g1078) & (!g1118) & (g2314) & (g2362) & (g2315) & (g2475)) + ((g1078) & (g1118) & (!g2314) & (!g2362) & (g2315) & (g2475)) + ((g1078) & (g1118) & (!g2314) & (g2362) & (!g2315) & (g2475)) + ((g1078) & (g1118) & (!g2314) & (g2362) & (g2315) & (g2475)) + ((g1078) & (g1118) & (g2314) & (!g2362) & (!g2315) & (g2475)) + ((g1078) & (g1118) & (g2314) & (!g2362) & (g2315) & (g2475)) + ((g1078) & (g1118) & (g2314) & (g2362) & (!g2315) & (g2475)) + ((g1078) & (g1118) & (g2314) & (g2362) & (g2315) & (g2475)));
	assign g2477 = (((g1145) & (g2393)));
	assign g2478 = (((!g2476) & (!g2477)));
	assign g2479 = (((!g827) & (!g1185) & (g2474) & (!g2478)) + ((!g827) & (!g1185) & (g2474) & (g2478)) + ((!g827) & (g1185) & (g2474) & (!g2478)) + ((!g827) & (g1185) & (g2474) & (g2478)) + ((g827) & (!g1185) & (!g2474) & (!g2478)) + ((g827) & (!g1185) & (g2474) & (g2478)) + ((g827) & (g1185) & (!g2474) & (g2478)) + ((g827) & (g1185) & (g2474) & (!g2478)));
	assign g8023 = (((!g2017) & (g4722) & (!g2480)) + ((!g2017) & (g4722) & (g2480)) + ((g2017) & (!g4722) & (g2480)) + ((g2017) & (g4722) & (g2480)));
	assign g2481 = (((!g1153) & (g2405)) + ((g1153) & (!g2405)));
	assign g2482 = (((!g1086) & (!g1120) & (g2326) & (g2364) & (g2327) & (g2481)) + ((!g1086) & (g1120) & (!g2326) & (g2364) & (!g2327) & (g2481)) + ((!g1086) & (g1120) & (!g2326) & (g2364) & (g2327) & (g2481)) + ((!g1086) & (g1120) & (g2326) & (!g2364) & (g2327) & (g2481)) + ((!g1086) & (g1120) & (g2326) & (g2364) & (!g2327) & (g2481)) + ((!g1086) & (g1120) & (g2326) & (g2364) & (g2327) & (g2481)) + ((g1086) & (!g1120) & (!g2326) & (g2364) & (g2327) & (g2481)) + ((g1086) & (!g1120) & (g2326) & (g2364) & (!g2327) & (g2481)) + ((g1086) & (!g1120) & (g2326) & (g2364) & (g2327) & (g2481)) + ((g1086) & (g1120) & (!g2326) & (!g2364) & (g2327) & (g2481)) + ((g1086) & (g1120) & (!g2326) & (g2364) & (!g2327) & (g2481)) + ((g1086) & (g1120) & (!g2326) & (g2364) & (g2327) & (g2481)) + ((g1086) & (g1120) & (g2326) & (!g2364) & (!g2327) & (g2481)) + ((g1086) & (g1120) & (g2326) & (!g2364) & (g2327) & (g2481)) + ((g1086) & (g1120) & (g2326) & (g2364) & (!g2327) & (g2481)) + ((g1086) & (g1120) & (g2326) & (g2364) & (g2327) & (g2481)));
	assign g2483 = (((g1153) & (g2405)));
	assign g2484 = (((!g2482) & (!g2483)));
	assign g2485 = (((!g827) & (!g1187) & (g2480) & (!g2484)) + ((!g827) & (!g1187) & (g2480) & (g2484)) + ((!g827) & (g1187) & (g2480) & (!g2484)) + ((!g827) & (g1187) & (g2480) & (g2484)) + ((g827) & (!g1187) & (!g2480) & (!g2484)) + ((g827) & (!g1187) & (g2480) & (g2484)) + ((g827) & (g1187) & (!g2480) & (g2484)) + ((g827) & (g1187) & (g2480) & (!g2484)));
	assign g8024 = (((!g3429) & (g4727) & (!g2486)) + ((!g3429) & (g4727) & (g2486)) + ((g3429) & (!g4727) & (g2486)) + ((g3429) & (g4727) & (g2486)));
	assign g2487 = (((!g1161) & (g2416)) + ((g1161) & (!g2416)));
	assign g2488 = (((!g1094) & (!g1122) & (g2337) & (g2366) & (g2338) & (g2487)) + ((!g1094) & (g1122) & (!g2337) & (g2366) & (!g2338) & (g2487)) + ((!g1094) & (g1122) & (!g2337) & (g2366) & (g2338) & (g2487)) + ((!g1094) & (g1122) & (g2337) & (!g2366) & (g2338) & (g2487)) + ((!g1094) & (g1122) & (g2337) & (g2366) & (!g2338) & (g2487)) + ((!g1094) & (g1122) & (g2337) & (g2366) & (g2338) & (g2487)) + ((g1094) & (!g1122) & (!g2337) & (g2366) & (g2338) & (g2487)) + ((g1094) & (!g1122) & (g2337) & (g2366) & (!g2338) & (g2487)) + ((g1094) & (!g1122) & (g2337) & (g2366) & (g2338) & (g2487)) + ((g1094) & (g1122) & (!g2337) & (!g2366) & (g2338) & (g2487)) + ((g1094) & (g1122) & (!g2337) & (g2366) & (!g2338) & (g2487)) + ((g1094) & (g1122) & (!g2337) & (g2366) & (g2338) & (g2487)) + ((g1094) & (g1122) & (g2337) & (!g2366) & (!g2338) & (g2487)) + ((g1094) & (g1122) & (g2337) & (!g2366) & (g2338) & (g2487)) + ((g1094) & (g1122) & (g2337) & (g2366) & (!g2338) & (g2487)) + ((g1094) & (g1122) & (g2337) & (g2366) & (g2338) & (g2487)));
	assign g2489 = (((g1161) & (g2416)));
	assign g2490 = (((!g2488) & (!g2489)));
	assign g2491 = (((!g827) & (!g1189) & (g2486) & (!g2490)) + ((!g827) & (!g1189) & (g2486) & (g2490)) + ((!g827) & (g1189) & (g2486) & (!g2490)) + ((!g827) & (g1189) & (g2486) & (g2490)) + ((g827) & (!g1189) & (!g2486) & (!g2490)) + ((g827) & (!g1189) & (g2486) & (g2490)) + ((g827) & (g1189) & (!g2486) & (g2490)) + ((g827) & (g1189) & (g2486) & (!g2490)));
	assign g2492 = (((!g1139) & (g2002)) + ((g1139) & (!g2002)));
	assign g2493 = (((!g1072) & (!g1124) & (g1997) & (g1999) & (g2307) & (g2492)) + ((!g1072) & (g1124) & (!g1997) & (g1999) & (!g2307) & (g2492)) + ((!g1072) & (g1124) & (!g1997) & (g1999) & (g2307) & (g2492)) + ((!g1072) & (g1124) & (g1997) & (!g1999) & (g2307) & (g2492)) + ((!g1072) & (g1124) & (g1997) & (g1999) & (!g2307) & (g2492)) + ((!g1072) & (g1124) & (g1997) & (g1999) & (g2307) & (g2492)) + ((g1072) & (!g1124) & (!g1997) & (g1999) & (g2307) & (g2492)) + ((g1072) & (!g1124) & (g1997) & (g1999) & (!g2307) & (g2492)) + ((g1072) & (!g1124) & (g1997) & (g1999) & (g2307) & (g2492)) + ((g1072) & (g1124) & (!g1997) & (!g1999) & (g2307) & (g2492)) + ((g1072) & (g1124) & (!g1997) & (g1999) & (!g2307) & (g2492)) + ((g1072) & (g1124) & (!g1997) & (g1999) & (g2307) & (g2492)) + ((g1072) & (g1124) & (g1997) & (!g1999) & (!g2307) & (g2492)) + ((g1072) & (g1124) & (g1997) & (!g1999) & (g2307) & (g2492)) + ((g1072) & (g1124) & (g1997) & (g1999) & (!g2307) & (g2492)) + ((g1072) & (g1124) & (g1997) & (g1999) & (g2307) & (g2492)));
	assign g2494 = (((g1139) & (g2002)));
	assign g2495 = (((!g2493) & (!g2494)));
	assign g2496 = (((!g827) & (!g1191) & (g2004) & (!g2495)) + ((!g827) & (!g1191) & (g2004) & (g2495)) + ((!g827) & (g1191) & (g2004) & (!g2495)) + ((!g827) & (g1191) & (g2004) & (g2495)) + ((g827) & (!g1191) & (!g2004) & (!g2495)) + ((g827) & (!g1191) & (g2004) & (g2495)) + ((g827) & (g1191) & (!g2004) & (g2495)) + ((g827) & (g1191) & (g2004) & (!g2495)));
	assign g8025 = (((!g3464) & (g4730) & (!g2497)) + ((!g3464) & (g4730) & (g2497)) + ((g3464) & (!g4730) & (g2497)) + ((g3464) & (g4730) & (g2497)));
	assign g2498 = (((!g1147) & (g2396)) + ((g1147) & (!g2396)));
	assign g2499 = (((!g1080) & (!g1126) & (g2317) & (g2369) & (g2318) & (g2498)) + ((!g1080) & (g1126) & (!g2317) & (g2369) & (!g2318) & (g2498)) + ((!g1080) & (g1126) & (!g2317) & (g2369) & (g2318) & (g2498)) + ((!g1080) & (g1126) & (g2317) & (!g2369) & (g2318) & (g2498)) + ((!g1080) & (g1126) & (g2317) & (g2369) & (!g2318) & (g2498)) + ((!g1080) & (g1126) & (g2317) & (g2369) & (g2318) & (g2498)) + ((g1080) & (!g1126) & (!g2317) & (g2369) & (g2318) & (g2498)) + ((g1080) & (!g1126) & (g2317) & (g2369) & (!g2318) & (g2498)) + ((g1080) & (!g1126) & (g2317) & (g2369) & (g2318) & (g2498)) + ((g1080) & (g1126) & (!g2317) & (!g2369) & (g2318) & (g2498)) + ((g1080) & (g1126) & (!g2317) & (g2369) & (!g2318) & (g2498)) + ((g1080) & (g1126) & (!g2317) & (g2369) & (g2318) & (g2498)) + ((g1080) & (g1126) & (g2317) & (!g2369) & (!g2318) & (g2498)) + ((g1080) & (g1126) & (g2317) & (!g2369) & (g2318) & (g2498)) + ((g1080) & (g1126) & (g2317) & (g2369) & (!g2318) & (g2498)) + ((g1080) & (g1126) & (g2317) & (g2369) & (g2318) & (g2498)));
	assign g2500 = (((g1147) & (g2396)));
	assign g2501 = (((!g2499) & (!g2500)));
	assign g2502 = (((!g827) & (!g1193) & (g2497) & (!g2501)) + ((!g827) & (!g1193) & (g2497) & (g2501)) + ((!g827) & (g1193) & (g2497) & (!g2501)) + ((!g827) & (g1193) & (g2497) & (g2501)) + ((g827) & (!g1193) & (!g2497) & (!g2501)) + ((g827) & (!g1193) & (g2497) & (g2501)) + ((g827) & (g1193) & (!g2497) & (g2501)) + ((g827) & (g1193) & (g2497) & (!g2501)));
	assign g8026 = (((!g3429) & (g4735) & (!g2503)) + ((!g3429) & (g4735) & (g2503)) + ((g3429) & (!g4735) & (g2503)) + ((g3429) & (g4735) & (g2503)));
	assign g2504 = (((!g1155) & (g2408)) + ((g1155) & (!g2408)));
	assign g2505 = (((!g1088) & (!g1128) & (g2329) & (g2371) & (g2330) & (g2504)) + ((!g1088) & (g1128) & (!g2329) & (g2371) & (!g2330) & (g2504)) + ((!g1088) & (g1128) & (!g2329) & (g2371) & (g2330) & (g2504)) + ((!g1088) & (g1128) & (g2329) & (!g2371) & (g2330) & (g2504)) + ((!g1088) & (g1128) & (g2329) & (g2371) & (!g2330) & (g2504)) + ((!g1088) & (g1128) & (g2329) & (g2371) & (g2330) & (g2504)) + ((g1088) & (!g1128) & (!g2329) & (g2371) & (g2330) & (g2504)) + ((g1088) & (!g1128) & (g2329) & (g2371) & (!g2330) & (g2504)) + ((g1088) & (!g1128) & (g2329) & (g2371) & (g2330) & (g2504)) + ((g1088) & (g1128) & (!g2329) & (!g2371) & (g2330) & (g2504)) + ((g1088) & (g1128) & (!g2329) & (g2371) & (!g2330) & (g2504)) + ((g1088) & (g1128) & (!g2329) & (g2371) & (g2330) & (g2504)) + ((g1088) & (g1128) & (g2329) & (!g2371) & (!g2330) & (g2504)) + ((g1088) & (g1128) & (g2329) & (!g2371) & (g2330) & (g2504)) + ((g1088) & (g1128) & (g2329) & (g2371) & (!g2330) & (g2504)) + ((g1088) & (g1128) & (g2329) & (g2371) & (g2330) & (g2504)));
	assign g2506 = (((g1155) & (g2408)));
	assign g2507 = (((!g2505) & (!g2506)));
	assign g2508 = (((!g827) & (!g1195) & (g2503) & (!g2507)) + ((!g827) & (!g1195) & (g2503) & (g2507)) + ((!g827) & (g1195) & (g2503) & (!g2507)) + ((!g827) & (g1195) & (g2503) & (g2507)) + ((g827) & (!g1195) & (!g2503) & (!g2507)) + ((g827) & (!g1195) & (g2503) & (g2507)) + ((g827) & (g1195) & (!g2503) & (g2507)) + ((g827) & (g1195) & (g2503) & (!g2507)));
	assign g8027 = (((!g2017) & (g4738) & (!g2509)) + ((!g2017) & (g4738) & (g2509)) + ((g2017) & (!g4738) & (g2509)) + ((g2017) & (g4738) & (g2509)));
	assign g2510 = (((!g1163) & (g2419)) + ((g1163) & (!g2419)));
	assign g2511 = (((!g1096) & (!g1130) & (g2340) & (g2373) & (g2341) & (g2510)) + ((!g1096) & (g1130) & (!g2340) & (g2373) & (!g2341) & (g2510)) + ((!g1096) & (g1130) & (!g2340) & (g2373) & (g2341) & (g2510)) + ((!g1096) & (g1130) & (g2340) & (!g2373) & (g2341) & (g2510)) + ((!g1096) & (g1130) & (g2340) & (g2373) & (!g2341) & (g2510)) + ((!g1096) & (g1130) & (g2340) & (g2373) & (g2341) & (g2510)) + ((g1096) & (!g1130) & (!g2340) & (g2373) & (g2341) & (g2510)) + ((g1096) & (!g1130) & (g2340) & (g2373) & (!g2341) & (g2510)) + ((g1096) & (!g1130) & (g2340) & (g2373) & (g2341) & (g2510)) + ((g1096) & (g1130) & (!g2340) & (!g2373) & (g2341) & (g2510)) + ((g1096) & (g1130) & (!g2340) & (g2373) & (!g2341) & (g2510)) + ((g1096) & (g1130) & (!g2340) & (g2373) & (g2341) & (g2510)) + ((g1096) & (g1130) & (g2340) & (!g2373) & (!g2341) & (g2510)) + ((g1096) & (g1130) & (g2340) & (!g2373) & (g2341) & (g2510)) + ((g1096) & (g1130) & (g2340) & (g2373) & (!g2341) & (g2510)) + ((g1096) & (g1130) & (g2340) & (g2373) & (g2341) & (g2510)));
	assign g2512 = (((g1163) & (g2419)));
	assign g2513 = (((!g2511) & (!g2512)));
	assign g2514 = (((!g827) & (!g1197) & (g2509) & (!g2513)) + ((!g827) & (!g1197) & (g2509) & (g2513)) + ((!g827) & (g1197) & (g2509) & (!g2513)) + ((!g827) & (g1197) & (g2509) & (g2513)) + ((g827) & (!g1197) & (!g2509) & (!g2513)) + ((g827) & (!g1197) & (g2509) & (g2513)) + ((g827) & (g1197) & (!g2509) & (g2513)) + ((g827) & (g1197) & (g2509) & (!g2513)));
	assign g8028 = (((!g3429) & (g4743) & (!g2515)) + ((!g3429) & (g4743) & (g2515)) + ((g3429) & (!g4743) & (g2515)) + ((g3429) & (g4743) & (g2515)));
	assign g8029 = (((!g3464) & (g4746) & (!g2516)) + ((!g3464) & (g4746) & (g2516)) + ((g3464) & (!g4746) & (g2516)) + ((g3464) & (g4746) & (g2516)));
	assign g2517 = (((!g2422) & (!g2423) & (!g2424) & (!g2515) & (g2516)) + ((!g2422) & (!g2423) & (!g2424) & (g2515) & (!g2516)) + ((!g2422) & (!g2423) & (g2424) & (!g2515) & (g2516)) + ((!g2422) & (!g2423) & (g2424) & (g2515) & (!g2516)) + ((!g2422) & (g2423) & (!g2424) & (!g2515) & (g2516)) + ((!g2422) & (g2423) & (!g2424) & (g2515) & (!g2516)) + ((!g2422) & (g2423) & (g2424) & (!g2515) & (!g2516)) + ((!g2422) & (g2423) & (g2424) & (g2515) & (g2516)) + ((g2422) & (!g2423) & (!g2424) & (!g2515) & (g2516)) + ((g2422) & (!g2423) & (!g2424) & (g2515) & (!g2516)) + ((g2422) & (!g2423) & (g2424) & (!g2515) & (!g2516)) + ((g2422) & (!g2423) & (g2424) & (g2515) & (g2516)) + ((g2422) & (g2423) & (!g2424) & (!g2515) & (!g2516)) + ((g2422) & (g2423) & (!g2424) & (g2515) & (g2516)) + ((g2422) & (g2423) & (g2424) & (!g2515) & (!g2516)) + ((g2422) & (g2423) & (g2424) & (g2515) & (g2516)));
	assign g8030 = (((!g3429) & (g4750) & (!g2518)) + ((!g3429) & (g4750) & (g2518)) + ((g3429) & (!g4750) & (g2518)) + ((g3429) & (g4750) & (g2518)));
	assign g8031 = (((!g3499) & (g4753) & (!g2519)) + ((!g3499) & (g4753) & (g2519)) + ((g3499) & (!g4753) & (g2519)) + ((g3499) & (g4753) & (g2519)));
	assign g2520 = (((!g2425) & (!g2426) & (!g2427) & (!g2518) & (g2519)) + ((!g2425) & (!g2426) & (!g2427) & (g2518) & (!g2519)) + ((!g2425) & (!g2426) & (g2427) & (!g2518) & (g2519)) + ((!g2425) & (!g2426) & (g2427) & (g2518) & (!g2519)) + ((!g2425) & (g2426) & (!g2427) & (!g2518) & (g2519)) + ((!g2425) & (g2426) & (!g2427) & (g2518) & (!g2519)) + ((!g2425) & (g2426) & (g2427) & (!g2518) & (!g2519)) + ((!g2425) & (g2426) & (g2427) & (g2518) & (g2519)) + ((g2425) & (!g2426) & (!g2427) & (!g2518) & (g2519)) + ((g2425) & (!g2426) & (!g2427) & (g2518) & (!g2519)) + ((g2425) & (!g2426) & (g2427) & (!g2518) & (!g2519)) + ((g2425) & (!g2426) & (g2427) & (g2518) & (g2519)) + ((g2425) & (g2426) & (!g2427) & (!g2518) & (!g2519)) + ((g2425) & (g2426) & (!g2427) & (g2518) & (g2519)) + ((g2425) & (g2426) & (g2427) & (!g2518) & (!g2519)) + ((g2425) & (g2426) & (g2427) & (g2518) & (g2519)));
	assign g2521 = (((!g830) & (!g1914) & (!g2517) & (!g2520) & (!g1199)) + ((!g830) & (!g1914) & (!g2517) & (!g2520) & (g1199)) + ((!g830) & (!g1914) & (!g2517) & (g2520) & (!g1199)) + ((!g830) & (!g1914) & (!g2517) & (g2520) & (g1199)) + ((!g830) & (!g1914) & (g2517) & (!g2520) & (!g1199)) + ((!g830) & (!g1914) & (g2517) & (!g2520) & (g1199)) + ((!g830) & (!g1914) & (g2517) & (g2520) & (!g1199)) + ((!g830) & (!g1914) & (g2517) & (g2520) & (g1199)) + ((!g830) & (g1914) & (!g2517) & (!g2520) & (!g1199)) + ((!g830) & (g1914) & (!g2517) & (!g2520) & (g1199)) + ((!g830) & (g1914) & (!g2517) & (g2520) & (!g1199)) + ((!g830) & (g1914) & (!g2517) & (g2520) & (g1199)) + ((!g830) & (g1914) & (g2517) & (!g2520) & (!g1199)) + ((!g830) & (g1914) & (g2517) & (!g2520) & (g1199)) + ((!g830) & (g1914) & (g2517) & (g2520) & (!g1199)) + ((!g830) & (g1914) & (g2517) & (g2520) & (g1199)) + ((g830) & (!g1914) & (!g2517) & (!g2520) & (g1199)) + ((g830) & (!g1914) & (!g2517) & (g2520) & (!g1199)) + ((g830) & (!g1914) & (g2517) & (!g2520) & (g1199)) + ((g830) & (!g1914) & (g2517) & (g2520) & (!g1199)) + ((g830) & (g1914) & (!g2517) & (!g2520) & (g1199)) + ((g830) & (g1914) & (!g2517) & (g2520) & (g1199)) + ((g830) & (g1914) & (g2517) & (!g2520) & (!g1199)) + ((g830) & (g1914) & (g2517) & (g2520) & (!g1199)));
	assign g2522 = (((!g827) & (!g1175) & (!g1206) & (!g2003) & (g2005) & (!g2448)) + ((!g827) & (!g1175) & (!g1206) & (!g2003) & (g2005) & (g2448)) + ((!g827) & (!g1175) & (!g1206) & (g2003) & (g2005) & (!g2448)) + ((!g827) & (!g1175) & (!g1206) & (g2003) & (g2005) & (g2448)) + ((!g827) & (!g1175) & (g1206) & (!g2003) & (g2005) & (!g2448)) + ((!g827) & (!g1175) & (g1206) & (!g2003) & (g2005) & (g2448)) + ((!g827) & (!g1175) & (g1206) & (g2003) & (g2005) & (!g2448)) + ((!g827) & (!g1175) & (g1206) & (g2003) & (g2005) & (g2448)) + ((!g827) & (g1175) & (!g1206) & (!g2003) & (g2005) & (!g2448)) + ((!g827) & (g1175) & (!g1206) & (!g2003) & (g2005) & (g2448)) + ((!g827) & (g1175) & (!g1206) & (g2003) & (g2005) & (!g2448)) + ((!g827) & (g1175) & (!g1206) & (g2003) & (g2005) & (g2448)) + ((!g827) & (g1175) & (g1206) & (!g2003) & (g2005) & (!g2448)) + ((!g827) & (g1175) & (g1206) & (!g2003) & (g2005) & (g2448)) + ((!g827) & (g1175) & (g1206) & (g2003) & (g2005) & (!g2448)) + ((!g827) & (g1175) & (g1206) & (g2003) & (g2005) & (g2448)) + ((g827) & (!g1175) & (!g1206) & (!g2003) & (g2005) & (!g2448)) + ((g827) & (!g1175) & (!g1206) & (!g2003) & (g2005) & (g2448)) + ((g827) & (!g1175) & (!g1206) & (g2003) & (!g2005) & (!g2448)) + ((g827) & (!g1175) & (!g1206) & (g2003) & (g2005) & (g2448)) + ((g827) & (!g1175) & (g1206) & (!g2003) & (!g2005) & (!g2448)) + ((g827) & (!g1175) & (g1206) & (!g2003) & (!g2005) & (g2448)) + ((g827) & (!g1175) & (g1206) & (g2003) & (!g2005) & (g2448)) + ((g827) & (!g1175) & (g1206) & (g2003) & (g2005) & (!g2448)) + ((g827) & (g1175) & (!g1206) & (!g2003) & (!g2005) & (!g2448)) + ((g827) & (g1175) & (!g1206) & (!g2003) & (g2005) & (g2448)) + ((g827) & (g1175) & (!g1206) & (g2003) & (!g2005) & (!g2448)) + ((g827) & (g1175) & (!g1206) & (g2003) & (!g2005) & (g2448)) + ((g827) & (g1175) & (g1206) & (!g2003) & (!g2005) & (g2448)) + ((g827) & (g1175) & (g1206) & (!g2003) & (g2005) & (!g2448)) + ((g827) & (g1175) & (g1206) & (g2003) & (g2005) & (!g2448)) + ((g827) & (g1175) & (g1206) & (g2003) & (g2005) & (g2448)));
	assign g8032 = (((!g3464) & (g6521) & (!g2523)) + ((!g3464) & (g6521) & (g2523)) + ((g3464) & (!g6521) & (g2523)) + ((g3464) & (g6521) & (g2523)));
	assign g2524 = (((!g827) & (!g1183) & (!g1208) & (!g2468) & (g2523) & (!g2472)) + ((!g827) & (!g1183) & (!g1208) & (!g2468) & (g2523) & (g2472)) + ((!g827) & (!g1183) & (!g1208) & (g2468) & (g2523) & (!g2472)) + ((!g827) & (!g1183) & (!g1208) & (g2468) & (g2523) & (g2472)) + ((!g827) & (!g1183) & (g1208) & (!g2468) & (g2523) & (!g2472)) + ((!g827) & (!g1183) & (g1208) & (!g2468) & (g2523) & (g2472)) + ((!g827) & (!g1183) & (g1208) & (g2468) & (g2523) & (!g2472)) + ((!g827) & (!g1183) & (g1208) & (g2468) & (g2523) & (g2472)) + ((!g827) & (g1183) & (!g1208) & (!g2468) & (g2523) & (!g2472)) + ((!g827) & (g1183) & (!g1208) & (!g2468) & (g2523) & (g2472)) + ((!g827) & (g1183) & (!g1208) & (g2468) & (g2523) & (!g2472)) + ((!g827) & (g1183) & (!g1208) & (g2468) & (g2523) & (g2472)) + ((!g827) & (g1183) & (g1208) & (!g2468) & (g2523) & (!g2472)) + ((!g827) & (g1183) & (g1208) & (!g2468) & (g2523) & (g2472)) + ((!g827) & (g1183) & (g1208) & (g2468) & (g2523) & (!g2472)) + ((!g827) & (g1183) & (g1208) & (g2468) & (g2523) & (g2472)) + ((g827) & (!g1183) & (!g1208) & (!g2468) & (g2523) & (!g2472)) + ((g827) & (!g1183) & (!g1208) & (!g2468) & (g2523) & (g2472)) + ((g827) & (!g1183) & (!g1208) & (g2468) & (!g2523) & (!g2472)) + ((g827) & (!g1183) & (!g1208) & (g2468) & (g2523) & (g2472)) + ((g827) & (!g1183) & (g1208) & (!g2468) & (!g2523) & (!g2472)) + ((g827) & (!g1183) & (g1208) & (!g2468) & (!g2523) & (g2472)) + ((g827) & (!g1183) & (g1208) & (g2468) & (!g2523) & (g2472)) + ((g827) & (!g1183) & (g1208) & (g2468) & (g2523) & (!g2472)) + ((g827) & (g1183) & (!g1208) & (!g2468) & (!g2523) & (!g2472)) + ((g827) & (g1183) & (!g1208) & (!g2468) & (g2523) & (g2472)) + ((g827) & (g1183) & (!g1208) & (g2468) & (!g2523) & (!g2472)) + ((g827) & (g1183) & (!g1208) & (g2468) & (!g2523) & (g2472)) + ((g827) & (g1183) & (g1208) & (!g2468) & (!g2523) & (g2472)) + ((g827) & (g1183) & (g1208) & (!g2468) & (g2523) & (!g2472)) + ((g827) & (g1183) & (g1208) & (g2468) & (g2523) & (!g2472)) + ((g827) & (g1183) & (g1208) & (g2468) & (g2523) & (g2472)));
	assign g2525 = (((!g827) & (!g1191) & (!g1210) & (!g2004) & (g2006) & (!g2495)) + ((!g827) & (!g1191) & (!g1210) & (!g2004) & (g2006) & (g2495)) + ((!g827) & (!g1191) & (!g1210) & (g2004) & (g2006) & (!g2495)) + ((!g827) & (!g1191) & (!g1210) & (g2004) & (g2006) & (g2495)) + ((!g827) & (!g1191) & (g1210) & (!g2004) & (g2006) & (!g2495)) + ((!g827) & (!g1191) & (g1210) & (!g2004) & (g2006) & (g2495)) + ((!g827) & (!g1191) & (g1210) & (g2004) & (g2006) & (!g2495)) + ((!g827) & (!g1191) & (g1210) & (g2004) & (g2006) & (g2495)) + ((!g827) & (g1191) & (!g1210) & (!g2004) & (g2006) & (!g2495)) + ((!g827) & (g1191) & (!g1210) & (!g2004) & (g2006) & (g2495)) + ((!g827) & (g1191) & (!g1210) & (g2004) & (g2006) & (!g2495)) + ((!g827) & (g1191) & (!g1210) & (g2004) & (g2006) & (g2495)) + ((!g827) & (g1191) & (g1210) & (!g2004) & (g2006) & (!g2495)) + ((!g827) & (g1191) & (g1210) & (!g2004) & (g2006) & (g2495)) + ((!g827) & (g1191) & (g1210) & (g2004) & (g2006) & (!g2495)) + ((!g827) & (g1191) & (g1210) & (g2004) & (g2006) & (g2495)) + ((g827) & (!g1191) & (!g1210) & (!g2004) & (g2006) & (!g2495)) + ((g827) & (!g1191) & (!g1210) & (!g2004) & (g2006) & (g2495)) + ((g827) & (!g1191) & (!g1210) & (g2004) & (!g2006) & (!g2495)) + ((g827) & (!g1191) & (!g1210) & (g2004) & (g2006) & (g2495)) + ((g827) & (!g1191) & (g1210) & (!g2004) & (!g2006) & (!g2495)) + ((g827) & (!g1191) & (g1210) & (!g2004) & (!g2006) & (g2495)) + ((g827) & (!g1191) & (g1210) & (g2004) & (!g2006) & (g2495)) + ((g827) & (!g1191) & (g1210) & (g2004) & (g2006) & (!g2495)) + ((g827) & (g1191) & (!g1210) & (!g2004) & (!g2006) & (!g2495)) + ((g827) & (g1191) & (!g1210) & (!g2004) & (g2006) & (g2495)) + ((g827) & (g1191) & (!g1210) & (g2004) & (!g2006) & (!g2495)) + ((g827) & (g1191) & (!g1210) & (g2004) & (!g2006) & (g2495)) + ((g827) & (g1191) & (g1210) & (!g2004) & (!g2006) & (g2495)) + ((g827) & (g1191) & (g1210) & (!g2004) & (g2006) & (!g2495)) + ((g827) & (g1191) & (g1210) & (g2004) & (g2006) & (!g2495)) + ((g827) & (g1191) & (g1210) & (g2004) & (g2006) & (g2495)));
	assign g2526 = (((!g827) & (!g1169) & (!g1212) & (!g1967) & (g1969) & (!g2432)) + ((!g827) & (!g1169) & (!g1212) & (!g1967) & (g1969) & (g2432)) + ((!g827) & (!g1169) & (!g1212) & (g1967) & (g1969) & (!g2432)) + ((!g827) & (!g1169) & (!g1212) & (g1967) & (g1969) & (g2432)) + ((!g827) & (!g1169) & (g1212) & (!g1967) & (g1969) & (!g2432)) + ((!g827) & (!g1169) & (g1212) & (!g1967) & (g1969) & (g2432)) + ((!g827) & (!g1169) & (g1212) & (g1967) & (g1969) & (!g2432)) + ((!g827) & (!g1169) & (g1212) & (g1967) & (g1969) & (g2432)) + ((!g827) & (g1169) & (!g1212) & (!g1967) & (g1969) & (!g2432)) + ((!g827) & (g1169) & (!g1212) & (!g1967) & (g1969) & (g2432)) + ((!g827) & (g1169) & (!g1212) & (g1967) & (g1969) & (!g2432)) + ((!g827) & (g1169) & (!g1212) & (g1967) & (g1969) & (g2432)) + ((!g827) & (g1169) & (g1212) & (!g1967) & (g1969) & (!g2432)) + ((!g827) & (g1169) & (g1212) & (!g1967) & (g1969) & (g2432)) + ((!g827) & (g1169) & (g1212) & (g1967) & (g1969) & (!g2432)) + ((!g827) & (g1169) & (g1212) & (g1967) & (g1969) & (g2432)) + ((g827) & (!g1169) & (!g1212) & (!g1967) & (g1969) & (!g2432)) + ((g827) & (!g1169) & (!g1212) & (!g1967) & (g1969) & (g2432)) + ((g827) & (!g1169) & (!g1212) & (g1967) & (!g1969) & (!g2432)) + ((g827) & (!g1169) & (!g1212) & (g1967) & (g1969) & (g2432)) + ((g827) & (!g1169) & (g1212) & (!g1967) & (!g1969) & (!g2432)) + ((g827) & (!g1169) & (g1212) & (!g1967) & (!g1969) & (g2432)) + ((g827) & (!g1169) & (g1212) & (g1967) & (!g1969) & (g2432)) + ((g827) & (!g1169) & (g1212) & (g1967) & (g1969) & (!g2432)) + ((g827) & (g1169) & (!g1212) & (!g1967) & (!g1969) & (!g2432)) + ((g827) & (g1169) & (!g1212) & (!g1967) & (g1969) & (g2432)) + ((g827) & (g1169) & (!g1212) & (g1967) & (!g1969) & (!g2432)) + ((g827) & (g1169) & (!g1212) & (g1967) & (!g1969) & (g2432)) + ((g827) & (g1169) & (g1212) & (!g1967) & (!g1969) & (g2432)) + ((g827) & (g1169) & (g1212) & (!g1967) & (g1969) & (!g2432)) + ((g827) & (g1169) & (g1212) & (g1967) & (g1969) & (!g2432)) + ((g827) & (g1169) & (g1212) & (g1967) & (g1969) & (g2432)));
	assign g8033 = (((!g2017) & (g6515) & (!g2527)) + ((!g2017) & (g6515) & (g2527)) + ((g2017) & (!g6515) & (g2527)) + ((g2017) & (g6515) & (g2527)));
	assign g2528 = (((!g827) & (!g1177) & (!g1214) & (!g2450) & (g2527) & (!g2454)) + ((!g827) & (!g1177) & (!g1214) & (!g2450) & (g2527) & (g2454)) + ((!g827) & (!g1177) & (!g1214) & (g2450) & (g2527) & (!g2454)) + ((!g827) & (!g1177) & (!g1214) & (g2450) & (g2527) & (g2454)) + ((!g827) & (!g1177) & (g1214) & (!g2450) & (g2527) & (!g2454)) + ((!g827) & (!g1177) & (g1214) & (!g2450) & (g2527) & (g2454)) + ((!g827) & (!g1177) & (g1214) & (g2450) & (g2527) & (!g2454)) + ((!g827) & (!g1177) & (g1214) & (g2450) & (g2527) & (g2454)) + ((!g827) & (g1177) & (!g1214) & (!g2450) & (g2527) & (!g2454)) + ((!g827) & (g1177) & (!g1214) & (!g2450) & (g2527) & (g2454)) + ((!g827) & (g1177) & (!g1214) & (g2450) & (g2527) & (!g2454)) + ((!g827) & (g1177) & (!g1214) & (g2450) & (g2527) & (g2454)) + ((!g827) & (g1177) & (g1214) & (!g2450) & (g2527) & (!g2454)) + ((!g827) & (g1177) & (g1214) & (!g2450) & (g2527) & (g2454)) + ((!g827) & (g1177) & (g1214) & (g2450) & (g2527) & (!g2454)) + ((!g827) & (g1177) & (g1214) & (g2450) & (g2527) & (g2454)) + ((g827) & (!g1177) & (!g1214) & (!g2450) & (g2527) & (!g2454)) + ((g827) & (!g1177) & (!g1214) & (!g2450) & (g2527) & (g2454)) + ((g827) & (!g1177) & (!g1214) & (g2450) & (!g2527) & (!g2454)) + ((g827) & (!g1177) & (!g1214) & (g2450) & (g2527) & (g2454)) + ((g827) & (!g1177) & (g1214) & (!g2450) & (!g2527) & (!g2454)) + ((g827) & (!g1177) & (g1214) & (!g2450) & (!g2527) & (g2454)) + ((g827) & (!g1177) & (g1214) & (g2450) & (!g2527) & (g2454)) + ((g827) & (!g1177) & (g1214) & (g2450) & (g2527) & (!g2454)) + ((g827) & (g1177) & (!g1214) & (!g2450) & (!g2527) & (!g2454)) + ((g827) & (g1177) & (!g1214) & (!g2450) & (g2527) & (g2454)) + ((g827) & (g1177) & (!g1214) & (g2450) & (!g2527) & (!g2454)) + ((g827) & (g1177) & (!g1214) & (g2450) & (!g2527) & (g2454)) + ((g827) & (g1177) & (g1214) & (!g2450) & (!g2527) & (g2454)) + ((g827) & (g1177) & (g1214) & (!g2450) & (g2527) & (!g2454)) + ((g827) & (g1177) & (g1214) & (g2450) & (g2527) & (!g2454)) + ((g827) & (g1177) & (g1214) & (g2450) & (g2527) & (g2454)));
	assign g8034 = (((!g3499) & (g6505) & (!g2529)) + ((!g3499) & (g6505) & (g2529)) + ((g3499) & (!g6505) & (g2529)) + ((g3499) & (g6505) & (g2529)));
	assign g2530 = (((!g827) & (!g1185) & (!g1216) & (!g2474) & (g2529) & (!g2478)) + ((!g827) & (!g1185) & (!g1216) & (!g2474) & (g2529) & (g2478)) + ((!g827) & (!g1185) & (!g1216) & (g2474) & (g2529) & (!g2478)) + ((!g827) & (!g1185) & (!g1216) & (g2474) & (g2529) & (g2478)) + ((!g827) & (!g1185) & (g1216) & (!g2474) & (g2529) & (!g2478)) + ((!g827) & (!g1185) & (g1216) & (!g2474) & (g2529) & (g2478)) + ((!g827) & (!g1185) & (g1216) & (g2474) & (g2529) & (!g2478)) + ((!g827) & (!g1185) & (g1216) & (g2474) & (g2529) & (g2478)) + ((!g827) & (g1185) & (!g1216) & (!g2474) & (g2529) & (!g2478)) + ((!g827) & (g1185) & (!g1216) & (!g2474) & (g2529) & (g2478)) + ((!g827) & (g1185) & (!g1216) & (g2474) & (g2529) & (!g2478)) + ((!g827) & (g1185) & (!g1216) & (g2474) & (g2529) & (g2478)) + ((!g827) & (g1185) & (g1216) & (!g2474) & (g2529) & (!g2478)) + ((!g827) & (g1185) & (g1216) & (!g2474) & (g2529) & (g2478)) + ((!g827) & (g1185) & (g1216) & (g2474) & (g2529) & (!g2478)) + ((!g827) & (g1185) & (g1216) & (g2474) & (g2529) & (g2478)) + ((g827) & (!g1185) & (!g1216) & (!g2474) & (g2529) & (!g2478)) + ((g827) & (!g1185) & (!g1216) & (!g2474) & (g2529) & (g2478)) + ((g827) & (!g1185) & (!g1216) & (g2474) & (!g2529) & (!g2478)) + ((g827) & (!g1185) & (!g1216) & (g2474) & (g2529) & (g2478)) + ((g827) & (!g1185) & (g1216) & (!g2474) & (!g2529) & (!g2478)) + ((g827) & (!g1185) & (g1216) & (!g2474) & (!g2529) & (g2478)) + ((g827) & (!g1185) & (g1216) & (g2474) & (!g2529) & (g2478)) + ((g827) & (!g1185) & (g1216) & (g2474) & (g2529) & (!g2478)) + ((g827) & (g1185) & (!g1216) & (!g2474) & (!g2529) & (!g2478)) + ((g827) & (g1185) & (!g1216) & (!g2474) & (g2529) & (g2478)) + ((g827) & (g1185) & (!g1216) & (g2474) & (!g2529) & (!g2478)) + ((g827) & (g1185) & (!g1216) & (g2474) & (!g2529) & (g2478)) + ((g827) & (g1185) & (g1216) & (!g2474) & (!g2529) & (g2478)) + ((g827) & (g1185) & (g1216) & (!g2474) & (g2529) & (!g2478)) + ((g827) & (g1185) & (g1216) & (g2474) & (g2529) & (!g2478)) + ((g827) & (g1185) & (g1216) & (g2474) & (g2529) & (g2478)));
	assign g8035 = (((!g3464) & (g6495) & (!g2531)) + ((!g3464) & (g6495) & (g2531)) + ((g3464) & (!g6495) & (g2531)) + ((g3464) & (g6495) & (g2531)));
	assign g2532 = (((!g827) & (!g1193) & (!g1218) & (!g2497) & (g2531) & (!g2501)) + ((!g827) & (!g1193) & (!g1218) & (!g2497) & (g2531) & (g2501)) + ((!g827) & (!g1193) & (!g1218) & (g2497) & (g2531) & (!g2501)) + ((!g827) & (!g1193) & (!g1218) & (g2497) & (g2531) & (g2501)) + ((!g827) & (!g1193) & (g1218) & (!g2497) & (g2531) & (!g2501)) + ((!g827) & (!g1193) & (g1218) & (!g2497) & (g2531) & (g2501)) + ((!g827) & (!g1193) & (g1218) & (g2497) & (g2531) & (!g2501)) + ((!g827) & (!g1193) & (g1218) & (g2497) & (g2531) & (g2501)) + ((!g827) & (g1193) & (!g1218) & (!g2497) & (g2531) & (!g2501)) + ((!g827) & (g1193) & (!g1218) & (!g2497) & (g2531) & (g2501)) + ((!g827) & (g1193) & (!g1218) & (g2497) & (g2531) & (!g2501)) + ((!g827) & (g1193) & (!g1218) & (g2497) & (g2531) & (g2501)) + ((!g827) & (g1193) & (g1218) & (!g2497) & (g2531) & (!g2501)) + ((!g827) & (g1193) & (g1218) & (!g2497) & (g2531) & (g2501)) + ((!g827) & (g1193) & (g1218) & (g2497) & (g2531) & (!g2501)) + ((!g827) & (g1193) & (g1218) & (g2497) & (g2531) & (g2501)) + ((g827) & (!g1193) & (!g1218) & (!g2497) & (g2531) & (!g2501)) + ((g827) & (!g1193) & (!g1218) & (!g2497) & (g2531) & (g2501)) + ((g827) & (!g1193) & (!g1218) & (g2497) & (!g2531) & (!g2501)) + ((g827) & (!g1193) & (!g1218) & (g2497) & (g2531) & (g2501)) + ((g827) & (!g1193) & (g1218) & (!g2497) & (!g2531) & (!g2501)) + ((g827) & (!g1193) & (g1218) & (!g2497) & (!g2531) & (g2501)) + ((g827) & (!g1193) & (g1218) & (g2497) & (!g2531) & (g2501)) + ((g827) & (!g1193) & (g1218) & (g2497) & (g2531) & (!g2501)) + ((g827) & (g1193) & (!g1218) & (!g2497) & (!g2531) & (!g2501)) + ((g827) & (g1193) & (!g1218) & (!g2497) & (g2531) & (g2501)) + ((g827) & (g1193) & (!g1218) & (g2497) & (!g2531) & (!g2501)) + ((g827) & (g1193) & (!g1218) & (g2497) & (!g2531) & (g2501)) + ((g827) & (g1193) & (g1218) & (!g2497) & (!g2531) & (g2501)) + ((g827) & (g1193) & (g1218) & (!g2497) & (g2531) & (!g2501)) + ((g827) & (g1193) & (g1218) & (g2497) & (g2531) & (!g2501)) + ((g827) & (g1193) & (g1218) & (g2497) & (g2531) & (g2501)));
	assign g8036 = (((!g3499) & (g6485) & (!g2533)) + ((!g3499) & (g6485) & (g2533)) + ((g3499) & (!g6485) & (g2533)) + ((g3499) & (g6485) & (g2533)));
	assign g2534 = (((!g827) & (!g1171) & (!g1220) & (!g2434) & (g2533) & (!g2438)) + ((!g827) & (!g1171) & (!g1220) & (!g2434) & (g2533) & (g2438)) + ((!g827) & (!g1171) & (!g1220) & (g2434) & (g2533) & (!g2438)) + ((!g827) & (!g1171) & (!g1220) & (g2434) & (g2533) & (g2438)) + ((!g827) & (!g1171) & (g1220) & (!g2434) & (g2533) & (!g2438)) + ((!g827) & (!g1171) & (g1220) & (!g2434) & (g2533) & (g2438)) + ((!g827) & (!g1171) & (g1220) & (g2434) & (g2533) & (!g2438)) + ((!g827) & (!g1171) & (g1220) & (g2434) & (g2533) & (g2438)) + ((!g827) & (g1171) & (!g1220) & (!g2434) & (g2533) & (!g2438)) + ((!g827) & (g1171) & (!g1220) & (!g2434) & (g2533) & (g2438)) + ((!g827) & (g1171) & (!g1220) & (g2434) & (g2533) & (!g2438)) + ((!g827) & (g1171) & (!g1220) & (g2434) & (g2533) & (g2438)) + ((!g827) & (g1171) & (g1220) & (!g2434) & (g2533) & (!g2438)) + ((!g827) & (g1171) & (g1220) & (!g2434) & (g2533) & (g2438)) + ((!g827) & (g1171) & (g1220) & (g2434) & (g2533) & (!g2438)) + ((!g827) & (g1171) & (g1220) & (g2434) & (g2533) & (g2438)) + ((g827) & (!g1171) & (!g1220) & (!g2434) & (g2533) & (!g2438)) + ((g827) & (!g1171) & (!g1220) & (!g2434) & (g2533) & (g2438)) + ((g827) & (!g1171) & (!g1220) & (g2434) & (!g2533) & (!g2438)) + ((g827) & (!g1171) & (!g1220) & (g2434) & (g2533) & (g2438)) + ((g827) & (!g1171) & (g1220) & (!g2434) & (!g2533) & (!g2438)) + ((g827) & (!g1171) & (g1220) & (!g2434) & (!g2533) & (g2438)) + ((g827) & (!g1171) & (g1220) & (g2434) & (!g2533) & (g2438)) + ((g827) & (!g1171) & (g1220) & (g2434) & (g2533) & (!g2438)) + ((g827) & (g1171) & (!g1220) & (!g2434) & (!g2533) & (!g2438)) + ((g827) & (g1171) & (!g1220) & (!g2434) & (g2533) & (g2438)) + ((g827) & (g1171) & (!g1220) & (g2434) & (!g2533) & (!g2438)) + ((g827) & (g1171) & (!g1220) & (g2434) & (!g2533) & (g2438)) + ((g827) & (g1171) & (g1220) & (!g2434) & (!g2533) & (g2438)) + ((g827) & (g1171) & (g1220) & (!g2434) & (g2533) & (!g2438)) + ((g827) & (g1171) & (g1220) & (g2434) & (g2533) & (!g2438)) + ((g827) & (g1171) & (g1220) & (g2434) & (g2533) & (g2438)));
	assign g8037 = (((!g3464) & (g6475) & (!g2535)) + ((!g3464) & (g6475) & (g2535)) + ((g3464) & (!g6475) & (g2535)) + ((g3464) & (g6475) & (g2535)));
	assign g2536 = (((!g827) & (!g1179) & (!g1222) & (!g2456) & (g2535) & (!g2460)) + ((!g827) & (!g1179) & (!g1222) & (!g2456) & (g2535) & (g2460)) + ((!g827) & (!g1179) & (!g1222) & (g2456) & (g2535) & (!g2460)) + ((!g827) & (!g1179) & (!g1222) & (g2456) & (g2535) & (g2460)) + ((!g827) & (!g1179) & (g1222) & (!g2456) & (g2535) & (!g2460)) + ((!g827) & (!g1179) & (g1222) & (!g2456) & (g2535) & (g2460)) + ((!g827) & (!g1179) & (g1222) & (g2456) & (g2535) & (!g2460)) + ((!g827) & (!g1179) & (g1222) & (g2456) & (g2535) & (g2460)) + ((!g827) & (g1179) & (!g1222) & (!g2456) & (g2535) & (!g2460)) + ((!g827) & (g1179) & (!g1222) & (!g2456) & (g2535) & (g2460)) + ((!g827) & (g1179) & (!g1222) & (g2456) & (g2535) & (!g2460)) + ((!g827) & (g1179) & (!g1222) & (g2456) & (g2535) & (g2460)) + ((!g827) & (g1179) & (g1222) & (!g2456) & (g2535) & (!g2460)) + ((!g827) & (g1179) & (g1222) & (!g2456) & (g2535) & (g2460)) + ((!g827) & (g1179) & (g1222) & (g2456) & (g2535) & (!g2460)) + ((!g827) & (g1179) & (g1222) & (g2456) & (g2535) & (g2460)) + ((g827) & (!g1179) & (!g1222) & (!g2456) & (g2535) & (!g2460)) + ((g827) & (!g1179) & (!g1222) & (!g2456) & (g2535) & (g2460)) + ((g827) & (!g1179) & (!g1222) & (g2456) & (!g2535) & (!g2460)) + ((g827) & (!g1179) & (!g1222) & (g2456) & (g2535) & (g2460)) + ((g827) & (!g1179) & (g1222) & (!g2456) & (!g2535) & (!g2460)) + ((g827) & (!g1179) & (g1222) & (!g2456) & (!g2535) & (g2460)) + ((g827) & (!g1179) & (g1222) & (g2456) & (!g2535) & (g2460)) + ((g827) & (!g1179) & (g1222) & (g2456) & (g2535) & (!g2460)) + ((g827) & (g1179) & (!g1222) & (!g2456) & (!g2535) & (!g2460)) + ((g827) & (g1179) & (!g1222) & (!g2456) & (g2535) & (g2460)) + ((g827) & (g1179) & (!g1222) & (g2456) & (!g2535) & (!g2460)) + ((g827) & (g1179) & (!g1222) & (g2456) & (!g2535) & (g2460)) + ((g827) & (g1179) & (g1222) & (!g2456) & (!g2535) & (g2460)) + ((g827) & (g1179) & (g1222) & (!g2456) & (g2535) & (!g2460)) + ((g827) & (g1179) & (g1222) & (g2456) & (g2535) & (!g2460)) + ((g827) & (g1179) & (g1222) & (g2456) & (g2535) & (g2460)));
	assign g8038 = (((!g2017) & (g6469) & (!g2537)) + ((!g2017) & (g6469) & (g2537)) + ((g2017) & (!g6469) & (g2537)) + ((g2017) & (g6469) & (g2537)));
	assign g2538 = (((!g827) & (!g1187) & (!g1224) & (!g2480) & (g2537) & (!g2484)) + ((!g827) & (!g1187) & (!g1224) & (!g2480) & (g2537) & (g2484)) + ((!g827) & (!g1187) & (!g1224) & (g2480) & (g2537) & (!g2484)) + ((!g827) & (!g1187) & (!g1224) & (g2480) & (g2537) & (g2484)) + ((!g827) & (!g1187) & (g1224) & (!g2480) & (g2537) & (!g2484)) + ((!g827) & (!g1187) & (g1224) & (!g2480) & (g2537) & (g2484)) + ((!g827) & (!g1187) & (g1224) & (g2480) & (g2537) & (!g2484)) + ((!g827) & (!g1187) & (g1224) & (g2480) & (g2537) & (g2484)) + ((!g827) & (g1187) & (!g1224) & (!g2480) & (g2537) & (!g2484)) + ((!g827) & (g1187) & (!g1224) & (!g2480) & (g2537) & (g2484)) + ((!g827) & (g1187) & (!g1224) & (g2480) & (g2537) & (!g2484)) + ((!g827) & (g1187) & (!g1224) & (g2480) & (g2537) & (g2484)) + ((!g827) & (g1187) & (g1224) & (!g2480) & (g2537) & (!g2484)) + ((!g827) & (g1187) & (g1224) & (!g2480) & (g2537) & (g2484)) + ((!g827) & (g1187) & (g1224) & (g2480) & (g2537) & (!g2484)) + ((!g827) & (g1187) & (g1224) & (g2480) & (g2537) & (g2484)) + ((g827) & (!g1187) & (!g1224) & (!g2480) & (g2537) & (!g2484)) + ((g827) & (!g1187) & (!g1224) & (!g2480) & (g2537) & (g2484)) + ((g827) & (!g1187) & (!g1224) & (g2480) & (!g2537) & (!g2484)) + ((g827) & (!g1187) & (!g1224) & (g2480) & (g2537) & (g2484)) + ((g827) & (!g1187) & (g1224) & (!g2480) & (!g2537) & (!g2484)) + ((g827) & (!g1187) & (g1224) & (!g2480) & (!g2537) & (g2484)) + ((g827) & (!g1187) & (g1224) & (g2480) & (!g2537) & (g2484)) + ((g827) & (!g1187) & (g1224) & (g2480) & (g2537) & (!g2484)) + ((g827) & (g1187) & (!g1224) & (!g2480) & (!g2537) & (!g2484)) + ((g827) & (g1187) & (!g1224) & (!g2480) & (g2537) & (g2484)) + ((g827) & (g1187) & (!g1224) & (g2480) & (!g2537) & (!g2484)) + ((g827) & (g1187) & (!g1224) & (g2480) & (!g2537) & (g2484)) + ((g827) & (g1187) & (g1224) & (!g2480) & (!g2537) & (g2484)) + ((g827) & (g1187) & (g1224) & (!g2480) & (g2537) & (!g2484)) + ((g827) & (g1187) & (g1224) & (g2480) & (g2537) & (!g2484)) + ((g827) & (g1187) & (g1224) & (g2480) & (g2537) & (g2484)));
	assign g8039 = (((!g3429) & (g4767) & (!g2539)) + ((!g3429) & (g4767) & (g2539)) + ((g3429) & (!g4767) & (g2539)) + ((g3429) & (g4767) & (g2539)));
	assign g2540 = (((!g827) & (!g1195) & (!g1226) & (!g2503) & (g2539) & (!g2507)) + ((!g827) & (!g1195) & (!g1226) & (!g2503) & (g2539) & (g2507)) + ((!g827) & (!g1195) & (!g1226) & (g2503) & (g2539) & (!g2507)) + ((!g827) & (!g1195) & (!g1226) & (g2503) & (g2539) & (g2507)) + ((!g827) & (!g1195) & (g1226) & (!g2503) & (g2539) & (!g2507)) + ((!g827) & (!g1195) & (g1226) & (!g2503) & (g2539) & (g2507)) + ((!g827) & (!g1195) & (g1226) & (g2503) & (g2539) & (!g2507)) + ((!g827) & (!g1195) & (g1226) & (g2503) & (g2539) & (g2507)) + ((!g827) & (g1195) & (!g1226) & (!g2503) & (g2539) & (!g2507)) + ((!g827) & (g1195) & (!g1226) & (!g2503) & (g2539) & (g2507)) + ((!g827) & (g1195) & (!g1226) & (g2503) & (g2539) & (!g2507)) + ((!g827) & (g1195) & (!g1226) & (g2503) & (g2539) & (g2507)) + ((!g827) & (g1195) & (g1226) & (!g2503) & (g2539) & (!g2507)) + ((!g827) & (g1195) & (g1226) & (!g2503) & (g2539) & (g2507)) + ((!g827) & (g1195) & (g1226) & (g2503) & (g2539) & (!g2507)) + ((!g827) & (g1195) & (g1226) & (g2503) & (g2539) & (g2507)) + ((g827) & (!g1195) & (!g1226) & (!g2503) & (g2539) & (!g2507)) + ((g827) & (!g1195) & (!g1226) & (!g2503) & (g2539) & (g2507)) + ((g827) & (!g1195) & (!g1226) & (g2503) & (!g2539) & (!g2507)) + ((g827) & (!g1195) & (!g1226) & (g2503) & (g2539) & (g2507)) + ((g827) & (!g1195) & (g1226) & (!g2503) & (!g2539) & (!g2507)) + ((g827) & (!g1195) & (g1226) & (!g2503) & (!g2539) & (g2507)) + ((g827) & (!g1195) & (g1226) & (g2503) & (!g2539) & (g2507)) + ((g827) & (!g1195) & (g1226) & (g2503) & (g2539) & (!g2507)) + ((g827) & (g1195) & (!g1226) & (!g2503) & (!g2539) & (!g2507)) + ((g827) & (g1195) & (!g1226) & (!g2503) & (g2539) & (g2507)) + ((g827) & (g1195) & (!g1226) & (g2503) & (!g2539) & (!g2507)) + ((g827) & (g1195) & (!g1226) & (g2503) & (!g2539) & (g2507)) + ((g827) & (g1195) & (g1226) & (!g2503) & (!g2539) & (g2507)) + ((g827) & (g1195) & (g1226) & (!g2503) & (g2539) & (!g2507)) + ((g827) & (g1195) & (g1226) & (g2503) & (g2539) & (!g2507)) + ((g827) & (g1195) & (g1226) & (g2503) & (g2539) & (g2507)));
	assign g2541 = (((!g827) & (!g1173) & (!g1228) & (!g1968) & (g1970) & (!g2443)) + ((!g827) & (!g1173) & (!g1228) & (!g1968) & (g1970) & (g2443)) + ((!g827) & (!g1173) & (!g1228) & (g1968) & (g1970) & (!g2443)) + ((!g827) & (!g1173) & (!g1228) & (g1968) & (g1970) & (g2443)) + ((!g827) & (!g1173) & (g1228) & (!g1968) & (g1970) & (!g2443)) + ((!g827) & (!g1173) & (g1228) & (!g1968) & (g1970) & (g2443)) + ((!g827) & (!g1173) & (g1228) & (g1968) & (g1970) & (!g2443)) + ((!g827) & (!g1173) & (g1228) & (g1968) & (g1970) & (g2443)) + ((!g827) & (g1173) & (!g1228) & (!g1968) & (g1970) & (!g2443)) + ((!g827) & (g1173) & (!g1228) & (!g1968) & (g1970) & (g2443)) + ((!g827) & (g1173) & (!g1228) & (g1968) & (g1970) & (!g2443)) + ((!g827) & (g1173) & (!g1228) & (g1968) & (g1970) & (g2443)) + ((!g827) & (g1173) & (g1228) & (!g1968) & (g1970) & (!g2443)) + ((!g827) & (g1173) & (g1228) & (!g1968) & (g1970) & (g2443)) + ((!g827) & (g1173) & (g1228) & (g1968) & (g1970) & (!g2443)) + ((!g827) & (g1173) & (g1228) & (g1968) & (g1970) & (g2443)) + ((g827) & (!g1173) & (!g1228) & (!g1968) & (g1970) & (!g2443)) + ((g827) & (!g1173) & (!g1228) & (!g1968) & (g1970) & (g2443)) + ((g827) & (!g1173) & (!g1228) & (g1968) & (!g1970) & (!g2443)) + ((g827) & (!g1173) & (!g1228) & (g1968) & (g1970) & (g2443)) + ((g827) & (!g1173) & (g1228) & (!g1968) & (!g1970) & (!g2443)) + ((g827) & (!g1173) & (g1228) & (!g1968) & (!g1970) & (g2443)) + ((g827) & (!g1173) & (g1228) & (g1968) & (!g1970) & (g2443)) + ((g827) & (!g1173) & (g1228) & (g1968) & (g1970) & (!g2443)) + ((g827) & (g1173) & (!g1228) & (!g1968) & (!g1970) & (!g2443)) + ((g827) & (g1173) & (!g1228) & (!g1968) & (g1970) & (g2443)) + ((g827) & (g1173) & (!g1228) & (g1968) & (!g1970) & (!g2443)) + ((g827) & (g1173) & (!g1228) & (g1968) & (!g1970) & (g2443)) + ((g827) & (g1173) & (g1228) & (!g1968) & (!g1970) & (g2443)) + ((g827) & (g1173) & (g1228) & (!g1968) & (g1970) & (!g2443)) + ((g827) & (g1173) & (g1228) & (g1968) & (g1970) & (!g2443)) + ((g827) & (g1173) & (g1228) & (g1968) & (g1970) & (g2443)));
	assign g8040 = (((!g3499) & (g6459) & (!g2542)) + ((!g3499) & (g6459) & (g2542)) + ((g3499) & (!g6459) & (g2542)) + ((g3499) & (g6459) & (g2542)));
	assign g2543 = (((!g827) & (!g1181) & (!g1230) & (!g2462) & (g2542) & (!g2466)) + ((!g827) & (!g1181) & (!g1230) & (!g2462) & (g2542) & (g2466)) + ((!g827) & (!g1181) & (!g1230) & (g2462) & (g2542) & (!g2466)) + ((!g827) & (!g1181) & (!g1230) & (g2462) & (g2542) & (g2466)) + ((!g827) & (!g1181) & (g1230) & (!g2462) & (g2542) & (!g2466)) + ((!g827) & (!g1181) & (g1230) & (!g2462) & (g2542) & (g2466)) + ((!g827) & (!g1181) & (g1230) & (g2462) & (g2542) & (!g2466)) + ((!g827) & (!g1181) & (g1230) & (g2462) & (g2542) & (g2466)) + ((!g827) & (g1181) & (!g1230) & (!g2462) & (g2542) & (!g2466)) + ((!g827) & (g1181) & (!g1230) & (!g2462) & (g2542) & (g2466)) + ((!g827) & (g1181) & (!g1230) & (g2462) & (g2542) & (!g2466)) + ((!g827) & (g1181) & (!g1230) & (g2462) & (g2542) & (g2466)) + ((!g827) & (g1181) & (g1230) & (!g2462) & (g2542) & (!g2466)) + ((!g827) & (g1181) & (g1230) & (!g2462) & (g2542) & (g2466)) + ((!g827) & (g1181) & (g1230) & (g2462) & (g2542) & (!g2466)) + ((!g827) & (g1181) & (g1230) & (g2462) & (g2542) & (g2466)) + ((g827) & (!g1181) & (!g1230) & (!g2462) & (g2542) & (!g2466)) + ((g827) & (!g1181) & (!g1230) & (!g2462) & (g2542) & (g2466)) + ((g827) & (!g1181) & (!g1230) & (g2462) & (!g2542) & (!g2466)) + ((g827) & (!g1181) & (!g1230) & (g2462) & (g2542) & (g2466)) + ((g827) & (!g1181) & (g1230) & (!g2462) & (!g2542) & (!g2466)) + ((g827) & (!g1181) & (g1230) & (!g2462) & (!g2542) & (g2466)) + ((g827) & (!g1181) & (g1230) & (g2462) & (!g2542) & (g2466)) + ((g827) & (!g1181) & (g1230) & (g2462) & (g2542) & (!g2466)) + ((g827) & (g1181) & (!g1230) & (!g2462) & (!g2542) & (!g2466)) + ((g827) & (g1181) & (!g1230) & (!g2462) & (g2542) & (g2466)) + ((g827) & (g1181) & (!g1230) & (g2462) & (!g2542) & (!g2466)) + ((g827) & (g1181) & (!g1230) & (g2462) & (!g2542) & (g2466)) + ((g827) & (g1181) & (g1230) & (!g2462) & (!g2542) & (g2466)) + ((g827) & (g1181) & (g1230) & (!g2462) & (g2542) & (!g2466)) + ((g827) & (g1181) & (g1230) & (g2462) & (g2542) & (!g2466)) + ((g827) & (g1181) & (g1230) & (g2462) & (g2542) & (g2466)));
	assign g8041 = (((!g3429) & (g4770) & (!g2544)) + ((!g3429) & (g4770) & (g2544)) + ((g3429) & (!g4770) & (g2544)) + ((g3429) & (g4770) & (g2544)));
	assign g2545 = (((!g827) & (!g1189) & (!g1232) & (!g2486) & (g2544) & (!g2490)) + ((!g827) & (!g1189) & (!g1232) & (!g2486) & (g2544) & (g2490)) + ((!g827) & (!g1189) & (!g1232) & (g2486) & (g2544) & (!g2490)) + ((!g827) & (!g1189) & (!g1232) & (g2486) & (g2544) & (g2490)) + ((!g827) & (!g1189) & (g1232) & (!g2486) & (g2544) & (!g2490)) + ((!g827) & (!g1189) & (g1232) & (!g2486) & (g2544) & (g2490)) + ((!g827) & (!g1189) & (g1232) & (g2486) & (g2544) & (!g2490)) + ((!g827) & (!g1189) & (g1232) & (g2486) & (g2544) & (g2490)) + ((!g827) & (g1189) & (!g1232) & (!g2486) & (g2544) & (!g2490)) + ((!g827) & (g1189) & (!g1232) & (!g2486) & (g2544) & (g2490)) + ((!g827) & (g1189) & (!g1232) & (g2486) & (g2544) & (!g2490)) + ((!g827) & (g1189) & (!g1232) & (g2486) & (g2544) & (g2490)) + ((!g827) & (g1189) & (g1232) & (!g2486) & (g2544) & (!g2490)) + ((!g827) & (g1189) & (g1232) & (!g2486) & (g2544) & (g2490)) + ((!g827) & (g1189) & (g1232) & (g2486) & (g2544) & (!g2490)) + ((!g827) & (g1189) & (g1232) & (g2486) & (g2544) & (g2490)) + ((g827) & (!g1189) & (!g1232) & (!g2486) & (g2544) & (!g2490)) + ((g827) & (!g1189) & (!g1232) & (!g2486) & (g2544) & (g2490)) + ((g827) & (!g1189) & (!g1232) & (g2486) & (!g2544) & (!g2490)) + ((g827) & (!g1189) & (!g1232) & (g2486) & (g2544) & (g2490)) + ((g827) & (!g1189) & (g1232) & (!g2486) & (!g2544) & (!g2490)) + ((g827) & (!g1189) & (g1232) & (!g2486) & (!g2544) & (g2490)) + ((g827) & (!g1189) & (g1232) & (g2486) & (!g2544) & (g2490)) + ((g827) & (!g1189) & (g1232) & (g2486) & (g2544) & (!g2490)) + ((g827) & (g1189) & (!g1232) & (!g2486) & (!g2544) & (!g2490)) + ((g827) & (g1189) & (!g1232) & (!g2486) & (g2544) & (g2490)) + ((g827) & (g1189) & (!g1232) & (g2486) & (!g2544) & (!g2490)) + ((g827) & (g1189) & (!g1232) & (g2486) & (!g2544) & (g2490)) + ((g827) & (g1189) & (g1232) & (!g2486) & (!g2544) & (g2490)) + ((g827) & (g1189) & (g1232) & (!g2486) & (g2544) & (!g2490)) + ((g827) & (g1189) & (g1232) & (g2486) & (g2544) & (!g2490)) + ((g827) & (g1189) & (g1232) & (g2486) & (g2544) & (g2490)));
	assign g8042 = (((!g2017) & (g6453) & (!g2546)) + ((!g2017) & (g6453) & (g2546)) + ((g2017) & (!g6453) & (g2546)) + ((g2017) & (g6453) & (g2546)));
	assign g2547 = (((!g827) & (!g1197) & (!g1234) & (!g2509) & (g2546) & (!g2513)) + ((!g827) & (!g1197) & (!g1234) & (!g2509) & (g2546) & (g2513)) + ((!g827) & (!g1197) & (!g1234) & (g2509) & (g2546) & (!g2513)) + ((!g827) & (!g1197) & (!g1234) & (g2509) & (g2546) & (g2513)) + ((!g827) & (!g1197) & (g1234) & (!g2509) & (g2546) & (!g2513)) + ((!g827) & (!g1197) & (g1234) & (!g2509) & (g2546) & (g2513)) + ((!g827) & (!g1197) & (g1234) & (g2509) & (g2546) & (!g2513)) + ((!g827) & (!g1197) & (g1234) & (g2509) & (g2546) & (g2513)) + ((!g827) & (g1197) & (!g1234) & (!g2509) & (g2546) & (!g2513)) + ((!g827) & (g1197) & (!g1234) & (!g2509) & (g2546) & (g2513)) + ((!g827) & (g1197) & (!g1234) & (g2509) & (g2546) & (!g2513)) + ((!g827) & (g1197) & (!g1234) & (g2509) & (g2546) & (g2513)) + ((!g827) & (g1197) & (g1234) & (!g2509) & (g2546) & (!g2513)) + ((!g827) & (g1197) & (g1234) & (!g2509) & (g2546) & (g2513)) + ((!g827) & (g1197) & (g1234) & (g2509) & (g2546) & (!g2513)) + ((!g827) & (g1197) & (g1234) & (g2509) & (g2546) & (g2513)) + ((g827) & (!g1197) & (!g1234) & (!g2509) & (g2546) & (!g2513)) + ((g827) & (!g1197) & (!g1234) & (!g2509) & (g2546) & (g2513)) + ((g827) & (!g1197) & (!g1234) & (g2509) & (!g2546) & (!g2513)) + ((g827) & (!g1197) & (!g1234) & (g2509) & (g2546) & (g2513)) + ((g827) & (!g1197) & (g1234) & (!g2509) & (!g2546) & (!g2513)) + ((g827) & (!g1197) & (g1234) & (!g2509) & (!g2546) & (g2513)) + ((g827) & (!g1197) & (g1234) & (g2509) & (!g2546) & (g2513)) + ((g827) & (!g1197) & (g1234) & (g2509) & (g2546) & (!g2513)) + ((g827) & (g1197) & (!g1234) & (!g2509) & (!g2546) & (!g2513)) + ((g827) & (g1197) & (!g1234) & (!g2509) & (g2546) & (g2513)) + ((g827) & (g1197) & (!g1234) & (g2509) & (!g2546) & (!g2513)) + ((g827) & (g1197) & (!g1234) & (g2509) & (!g2546) & (g2513)) + ((g827) & (g1197) & (g1234) & (!g2509) & (!g2546) & (g2513)) + ((g827) & (g1197) & (g1234) & (!g2509) & (g2546) & (!g2513)) + ((g827) & (g1197) & (g1234) & (g2509) & (g2546) & (!g2513)) + ((g827) & (g1197) & (g1234) & (g2509) & (g2546) & (g2513)));
	assign g2548 = (((!g2515) & (g2516)) + ((g2515) & (!g2516)));
	assign g2549 = (((!g2375) & (!g2376) & (!g2377) & (g2423) & (g2424) & (g2548)) + ((!g2375) & (!g2376) & (g2377) & (g2423) & (g2424) & (g2548)) + ((!g2375) & (g2376) & (!g2377) & (g2423) & (g2424) & (g2548)) + ((!g2375) & (g2376) & (g2377) & (!g2423) & (g2424) & (g2548)) + ((!g2375) & (g2376) & (g2377) & (g2423) & (!g2424) & (g2548)) + ((!g2375) & (g2376) & (g2377) & (g2423) & (g2424) & (g2548)) + ((g2375) & (!g2376) & (!g2377) & (g2423) & (g2424) & (g2548)) + ((g2375) & (!g2376) & (g2377) & (!g2423) & (g2424) & (g2548)) + ((g2375) & (!g2376) & (g2377) & (g2423) & (!g2424) & (g2548)) + ((g2375) & (!g2376) & (g2377) & (g2423) & (g2424) & (g2548)) + ((g2375) & (g2376) & (!g2377) & (!g2423) & (g2424) & (g2548)) + ((g2375) & (g2376) & (!g2377) & (g2423) & (!g2424) & (g2548)) + ((g2375) & (g2376) & (!g2377) & (g2423) & (g2424) & (g2548)) + ((g2375) & (g2376) & (g2377) & (!g2423) & (g2424) & (g2548)) + ((g2375) & (g2376) & (g2377) & (g2423) & (!g2424) & (g2548)) + ((g2375) & (g2376) & (g2377) & (g2423) & (g2424) & (g2548)));
	assign g2550 = (((g2515) & (g2516)));
	assign g8043 = (((!g3429) & (g4778) & (!g2551)) + ((!g3429) & (g4778) & (g2551)) + ((g3429) & (!g4778) & (g2551)) + ((g3429) & (g4778) & (g2551)));
	assign g8044 = (((!g3464) & (g4782) & (!g2552)) + ((!g3464) & (g4782) & (g2552)) + ((g3464) & (!g4782) & (g2552)) + ((g3464) & (g4782) & (g2552)));
	assign g2553 = (((!g2549) & (!g2550) & (!g2551) & (g2552)) + ((!g2549) & (!g2550) & (g2551) & (!g2552)) + ((!g2549) & (g2550) & (!g2551) & (!g2552)) + ((!g2549) & (g2550) & (g2551) & (g2552)) + ((g2549) & (!g2550) & (!g2551) & (!g2552)) + ((g2549) & (!g2550) & (g2551) & (g2552)) + ((g2549) & (g2550) & (!g2551) & (!g2552)) + ((g2549) & (g2550) & (g2551) & (g2552)));
	assign g2554 = (((!g2346) & (!g2347) & (!g2348) & (!g5723) & (!g5724)) + ((!g2346) & (!g2347) & (g2348) & (!g5723) & (!g5724)) + ((!g2346) & (g2347) & (!g2348) & (!g5723) & (!g5724)) + ((!g2346) & (g2347) & (g2348) & (!g5723) & (!g5724)) + ((!g2346) & (g2347) & (g2348) & (!g5723) & (g5724)) + ((g2346) & (!g2347) & (!g2348) & (!g5723) & (!g5724)) + ((g2346) & (!g2347) & (g2348) & (!g5723) & (!g5724)) + ((g2346) & (!g2347) & (g2348) & (!g5723) & (g5724)) + ((g2346) & (g2347) & (!g2348) & (!g5723) & (!g5724)) + ((g2346) & (g2347) & (!g2348) & (!g5723) & (g5724)) + ((g2346) & (g2347) & (g2348) & (!g5723) & (!g5724)) + ((g2346) & (g2347) & (g2348) & (!g5723) & (g5724)));
	assign g8045 = (((!g3429) & (g4785) & (!g2555)) + ((!g3429) & (g4785) & (g2555)) + ((g3429) & (!g4785) & (g2555)) + ((g3429) & (g4785) & (g2555)));
	assign g8046 = (((!g3499) & (g4789) & (!g2556)) + ((!g3499) & (g4789) & (g2556)) + ((g3499) & (!g4789) & (g2556)) + ((g3499) & (g4789) & (g2556)));
	assign g2557 = (((!g1169) & (!g1212) & (!g1967) & (!g1969) & (!g2430) & (!g2431)) + ((!g1169) & (!g1212) & (!g1967) & (!g1969) & (!g2430) & (g2431)) + ((!g1169) & (!g1212) & (!g1967) & (!g1969) & (g2430) & (!g2431)) + ((!g1169) & (!g1212) & (!g1967) & (!g1969) & (g2430) & (g2431)) + ((!g1169) & (!g1212) & (!g1967) & (g1969) & (!g2430) & (!g2431)) + ((!g1169) & (!g1212) & (!g1967) & (g1969) & (!g2430) & (g2431)) + ((!g1169) & (!g1212) & (!g1967) & (g1969) & (g2430) & (!g2431)) + ((!g1169) & (!g1212) & (!g1967) & (g1969) & (g2430) & (g2431)) + ((!g1169) & (!g1212) & (g1967) & (!g1969) & (!g2430) & (!g2431)) + ((!g1169) & (!g1212) & (g1967) & (!g1969) & (!g2430) & (g2431)) + ((!g1169) & (!g1212) & (g1967) & (!g1969) & (g2430) & (!g2431)) + ((!g1169) & (!g1212) & (g1967) & (!g1969) & (g2430) & (g2431)) + ((!g1169) & (!g1212) & (g1967) & (g1969) & (!g2430) & (!g2431)) + ((!g1169) & (g1212) & (!g1967) & (!g1969) & (!g2430) & (!g2431)) + ((!g1169) & (g1212) & (!g1967) & (!g1969) & (!g2430) & (g2431)) + ((!g1169) & (g1212) & (!g1967) & (!g1969) & (g2430) & (!g2431)) + ((!g1169) & (g1212) & (!g1967) & (!g1969) & (g2430) & (g2431)) + ((!g1169) & (g1212) & (g1967) & (!g1969) & (!g2430) & (!g2431)) + ((g1169) & (!g1212) & (!g1967) & (!g1969) & (!g2430) & (!g2431)) + ((g1169) & (!g1212) & (!g1967) & (!g1969) & (!g2430) & (g2431)) + ((g1169) & (!g1212) & (!g1967) & (!g1969) & (g2430) & (!g2431)) + ((g1169) & (!g1212) & (!g1967) & (!g1969) & (g2430) & (g2431)) + ((g1169) & (!g1212) & (!g1967) & (g1969) & (!g2430) & (!g2431)) + ((g1169) & (!g1212) & (g1967) & (!g1969) & (!g2430) & (!g2431)) + ((g1169) & (!g1212) & (g1967) & (!g1969) & (!g2430) & (g2431)) + ((g1169) & (!g1212) & (g1967) & (!g1969) & (g2430) & (!g2431)) + ((g1169) & (!g1212) & (g1967) & (!g1969) & (g2430) & (g2431)) + ((g1169) & (g1212) & (!g1967) & (!g1969) & (!g2430) & (!g2431)));
	assign g2558 = (((!g827) & (!g1239) & (g1972) & (!g2557)) + ((!g827) & (!g1239) & (g1972) & (g2557)) + ((!g827) & (g1239) & (g1972) & (!g2557)) + ((!g827) & (g1239) & (g1972) & (g2557)) + ((g827) & (!g1239) & (!g1972) & (!g2557)) + ((g827) & (!g1239) & (g1972) & (g2557)) + ((g827) & (g1239) & (!g1972) & (g2557)) + ((g827) & (g1239) & (g1972) & (!g2557)));
	assign g8047 = (((!g3499) & (g4792) & (!g2559)) + ((!g3499) & (g4792) & (g2559)) + ((g3499) & (!g4792) & (g2559)) + ((g3499) & (g4792) & (g2559)));
	assign g2560 = (((!g1171) & (!g1220) & (!g2434) & (!g2533) & (!g2436) & (!g2437)) + ((!g1171) & (!g1220) & (!g2434) & (!g2533) & (!g2436) & (g2437)) + ((!g1171) & (!g1220) & (!g2434) & (!g2533) & (g2436) & (!g2437)) + ((!g1171) & (!g1220) & (!g2434) & (!g2533) & (g2436) & (g2437)) + ((!g1171) & (!g1220) & (!g2434) & (g2533) & (!g2436) & (!g2437)) + ((!g1171) & (!g1220) & (!g2434) & (g2533) & (!g2436) & (g2437)) + ((!g1171) & (!g1220) & (!g2434) & (g2533) & (g2436) & (!g2437)) + ((!g1171) & (!g1220) & (!g2434) & (g2533) & (g2436) & (g2437)) + ((!g1171) & (!g1220) & (g2434) & (!g2533) & (!g2436) & (!g2437)) + ((!g1171) & (!g1220) & (g2434) & (!g2533) & (!g2436) & (g2437)) + ((!g1171) & (!g1220) & (g2434) & (!g2533) & (g2436) & (!g2437)) + ((!g1171) & (!g1220) & (g2434) & (!g2533) & (g2436) & (g2437)) + ((!g1171) & (!g1220) & (g2434) & (g2533) & (!g2436) & (!g2437)) + ((!g1171) & (g1220) & (!g2434) & (!g2533) & (!g2436) & (!g2437)) + ((!g1171) & (g1220) & (!g2434) & (!g2533) & (!g2436) & (g2437)) + ((!g1171) & (g1220) & (!g2434) & (!g2533) & (g2436) & (!g2437)) + ((!g1171) & (g1220) & (!g2434) & (!g2533) & (g2436) & (g2437)) + ((!g1171) & (g1220) & (g2434) & (!g2533) & (!g2436) & (!g2437)) + ((g1171) & (!g1220) & (!g2434) & (!g2533) & (!g2436) & (!g2437)) + ((g1171) & (!g1220) & (!g2434) & (!g2533) & (!g2436) & (g2437)) + ((g1171) & (!g1220) & (!g2434) & (!g2533) & (g2436) & (!g2437)) + ((g1171) & (!g1220) & (!g2434) & (!g2533) & (g2436) & (g2437)) + ((g1171) & (!g1220) & (!g2434) & (g2533) & (!g2436) & (!g2437)) + ((g1171) & (!g1220) & (g2434) & (!g2533) & (!g2436) & (!g2437)) + ((g1171) & (!g1220) & (g2434) & (!g2533) & (!g2436) & (g2437)) + ((g1171) & (!g1220) & (g2434) & (!g2533) & (g2436) & (!g2437)) + ((g1171) & (!g1220) & (g2434) & (!g2533) & (g2436) & (g2437)) + ((g1171) & (g1220) & (!g2434) & (!g2533) & (!g2436) & (!g2437)));
	assign g2561 = (((!g827) & (!g1241) & (g2559) & (!g2560)) + ((!g827) & (!g1241) & (g2559) & (g2560)) + ((!g827) & (g1241) & (g2559) & (!g2560)) + ((!g827) & (g1241) & (g2559) & (g2560)) + ((g827) & (!g1241) & (!g2559) & (!g2560)) + ((g827) & (!g1241) & (g2559) & (g2560)) + ((g827) & (g1241) & (!g2559) & (g2560)) + ((g827) & (g1241) & (g2559) & (!g2560)));
	assign g2562 = (((!g1173) & (!g1228) & (!g1968) & (!g1970) & (!g2441) & (!g2442)) + ((!g1173) & (!g1228) & (!g1968) & (!g1970) & (!g2441) & (g2442)) + ((!g1173) & (!g1228) & (!g1968) & (!g1970) & (g2441) & (!g2442)) + ((!g1173) & (!g1228) & (!g1968) & (!g1970) & (g2441) & (g2442)) + ((!g1173) & (!g1228) & (!g1968) & (g1970) & (!g2441) & (!g2442)) + ((!g1173) & (!g1228) & (!g1968) & (g1970) & (!g2441) & (g2442)) + ((!g1173) & (!g1228) & (!g1968) & (g1970) & (g2441) & (!g2442)) + ((!g1173) & (!g1228) & (!g1968) & (g1970) & (g2441) & (g2442)) + ((!g1173) & (!g1228) & (g1968) & (!g1970) & (!g2441) & (!g2442)) + ((!g1173) & (!g1228) & (g1968) & (!g1970) & (!g2441) & (g2442)) + ((!g1173) & (!g1228) & (g1968) & (!g1970) & (g2441) & (!g2442)) + ((!g1173) & (!g1228) & (g1968) & (!g1970) & (g2441) & (g2442)) + ((!g1173) & (!g1228) & (g1968) & (g1970) & (!g2441) & (!g2442)) + ((!g1173) & (g1228) & (!g1968) & (!g1970) & (!g2441) & (!g2442)) + ((!g1173) & (g1228) & (!g1968) & (!g1970) & (!g2441) & (g2442)) + ((!g1173) & (g1228) & (!g1968) & (!g1970) & (g2441) & (!g2442)) + ((!g1173) & (g1228) & (!g1968) & (!g1970) & (g2441) & (g2442)) + ((!g1173) & (g1228) & (g1968) & (!g1970) & (!g2441) & (!g2442)) + ((g1173) & (!g1228) & (!g1968) & (!g1970) & (!g2441) & (!g2442)) + ((g1173) & (!g1228) & (!g1968) & (!g1970) & (!g2441) & (g2442)) + ((g1173) & (!g1228) & (!g1968) & (!g1970) & (g2441) & (!g2442)) + ((g1173) & (!g1228) & (!g1968) & (!g1970) & (g2441) & (g2442)) + ((g1173) & (!g1228) & (!g1968) & (g1970) & (!g2441) & (!g2442)) + ((g1173) & (!g1228) & (g1968) & (!g1970) & (!g2441) & (!g2442)) + ((g1173) & (!g1228) & (g1968) & (!g1970) & (!g2441) & (g2442)) + ((g1173) & (!g1228) & (g1968) & (!g1970) & (g2441) & (!g2442)) + ((g1173) & (!g1228) & (g1968) & (!g1970) & (g2441) & (g2442)) + ((g1173) & (g1228) & (!g1968) & (!g1970) & (!g2441) & (!g2442)));
	assign g2563 = (((!g827) & (!g1243) & (g1973) & (!g2562)) + ((!g827) & (!g1243) & (g1973) & (g2562)) + ((!g827) & (g1243) & (g1973) & (!g2562)) + ((!g827) & (g1243) & (g1973) & (g2562)) + ((g827) & (!g1243) & (!g1973) & (!g2562)) + ((g827) & (!g1243) & (g1973) & (g2562)) + ((g827) & (g1243) & (!g1973) & (g2562)) + ((g827) & (g1243) & (g1973) & (!g2562)));
	assign g2564 = (((!g1175) & (!g1206) & (!g2003) & (!g2005) & (!g2446) & (!g2447)) + ((!g1175) & (!g1206) & (!g2003) & (!g2005) & (!g2446) & (g2447)) + ((!g1175) & (!g1206) & (!g2003) & (!g2005) & (g2446) & (!g2447)) + ((!g1175) & (!g1206) & (!g2003) & (!g2005) & (g2446) & (g2447)) + ((!g1175) & (!g1206) & (!g2003) & (g2005) & (!g2446) & (!g2447)) + ((!g1175) & (!g1206) & (!g2003) & (g2005) & (!g2446) & (g2447)) + ((!g1175) & (!g1206) & (!g2003) & (g2005) & (g2446) & (!g2447)) + ((!g1175) & (!g1206) & (!g2003) & (g2005) & (g2446) & (g2447)) + ((!g1175) & (!g1206) & (g2003) & (!g2005) & (!g2446) & (!g2447)) + ((!g1175) & (!g1206) & (g2003) & (!g2005) & (!g2446) & (g2447)) + ((!g1175) & (!g1206) & (g2003) & (!g2005) & (g2446) & (!g2447)) + ((!g1175) & (!g1206) & (g2003) & (!g2005) & (g2446) & (g2447)) + ((!g1175) & (!g1206) & (g2003) & (g2005) & (!g2446) & (!g2447)) + ((!g1175) & (g1206) & (!g2003) & (!g2005) & (!g2446) & (!g2447)) + ((!g1175) & (g1206) & (!g2003) & (!g2005) & (!g2446) & (g2447)) + ((!g1175) & (g1206) & (!g2003) & (!g2005) & (g2446) & (!g2447)) + ((!g1175) & (g1206) & (!g2003) & (!g2005) & (g2446) & (g2447)) + ((!g1175) & (g1206) & (g2003) & (!g2005) & (!g2446) & (!g2447)) + ((g1175) & (!g1206) & (!g2003) & (!g2005) & (!g2446) & (!g2447)) + ((g1175) & (!g1206) & (!g2003) & (!g2005) & (!g2446) & (g2447)) + ((g1175) & (!g1206) & (!g2003) & (!g2005) & (g2446) & (!g2447)) + ((g1175) & (!g1206) & (!g2003) & (!g2005) & (g2446) & (g2447)) + ((g1175) & (!g1206) & (!g2003) & (g2005) & (!g2446) & (!g2447)) + ((g1175) & (!g1206) & (g2003) & (!g2005) & (!g2446) & (!g2447)) + ((g1175) & (!g1206) & (g2003) & (!g2005) & (!g2446) & (g2447)) + ((g1175) & (!g1206) & (g2003) & (!g2005) & (g2446) & (!g2447)) + ((g1175) & (!g1206) & (g2003) & (!g2005) & (g2446) & (g2447)) + ((g1175) & (g1206) & (!g2003) & (!g2005) & (!g2446) & (!g2447)));
	assign g2565 = (((!g827) & (!g1245) & (g2011) & (!g2564)) + ((!g827) & (!g1245) & (g2011) & (g2564)) + ((!g827) & (g1245) & (g2011) & (!g2564)) + ((!g827) & (g1245) & (g2011) & (g2564)) + ((g827) & (!g1245) & (!g2011) & (!g2564)) + ((g827) & (!g1245) & (g2011) & (g2564)) + ((g827) & (g1245) & (!g2011) & (g2564)) + ((g827) & (g1245) & (g2011) & (!g2564)));
	assign g8048 = (((!g2017) & (g4795) & (!g2566)) + ((!g2017) & (g4795) & (g2566)) + ((g2017) & (!g4795) & (g2566)) + ((g2017) & (g4795) & (g2566)));
	assign g2567 = (((!g1177) & (!g1214) & (!g2450) & (!g2527) & (!g2452) & (!g2453)) + ((!g1177) & (!g1214) & (!g2450) & (!g2527) & (!g2452) & (g2453)) + ((!g1177) & (!g1214) & (!g2450) & (!g2527) & (g2452) & (!g2453)) + ((!g1177) & (!g1214) & (!g2450) & (!g2527) & (g2452) & (g2453)) + ((!g1177) & (!g1214) & (!g2450) & (g2527) & (!g2452) & (!g2453)) + ((!g1177) & (!g1214) & (!g2450) & (g2527) & (!g2452) & (g2453)) + ((!g1177) & (!g1214) & (!g2450) & (g2527) & (g2452) & (!g2453)) + ((!g1177) & (!g1214) & (!g2450) & (g2527) & (g2452) & (g2453)) + ((!g1177) & (!g1214) & (g2450) & (!g2527) & (!g2452) & (!g2453)) + ((!g1177) & (!g1214) & (g2450) & (!g2527) & (!g2452) & (g2453)) + ((!g1177) & (!g1214) & (g2450) & (!g2527) & (g2452) & (!g2453)) + ((!g1177) & (!g1214) & (g2450) & (!g2527) & (g2452) & (g2453)) + ((!g1177) & (!g1214) & (g2450) & (g2527) & (!g2452) & (!g2453)) + ((!g1177) & (g1214) & (!g2450) & (!g2527) & (!g2452) & (!g2453)) + ((!g1177) & (g1214) & (!g2450) & (!g2527) & (!g2452) & (g2453)) + ((!g1177) & (g1214) & (!g2450) & (!g2527) & (g2452) & (!g2453)) + ((!g1177) & (g1214) & (!g2450) & (!g2527) & (g2452) & (g2453)) + ((!g1177) & (g1214) & (g2450) & (!g2527) & (!g2452) & (!g2453)) + ((g1177) & (!g1214) & (!g2450) & (!g2527) & (!g2452) & (!g2453)) + ((g1177) & (!g1214) & (!g2450) & (!g2527) & (!g2452) & (g2453)) + ((g1177) & (!g1214) & (!g2450) & (!g2527) & (g2452) & (!g2453)) + ((g1177) & (!g1214) & (!g2450) & (!g2527) & (g2452) & (g2453)) + ((g1177) & (!g1214) & (!g2450) & (g2527) & (!g2452) & (!g2453)) + ((g1177) & (!g1214) & (g2450) & (!g2527) & (!g2452) & (!g2453)) + ((g1177) & (!g1214) & (g2450) & (!g2527) & (!g2452) & (g2453)) + ((g1177) & (!g1214) & (g2450) & (!g2527) & (g2452) & (!g2453)) + ((g1177) & (!g1214) & (g2450) & (!g2527) & (g2452) & (g2453)) + ((g1177) & (g1214) & (!g2450) & (!g2527) & (!g2452) & (!g2453)));
	assign g2568 = (((!g827) & (!g1247) & (g2566) & (!g2567)) + ((!g827) & (!g1247) & (g2566) & (g2567)) + ((!g827) & (g1247) & (g2566) & (!g2567)) + ((!g827) & (g1247) & (g2566) & (g2567)) + ((g827) & (!g1247) & (!g2566) & (!g2567)) + ((g827) & (!g1247) & (g2566) & (g2567)) + ((g827) & (g1247) & (!g2566) & (g2567)) + ((g827) & (g1247) & (g2566) & (!g2567)));
	assign g8049 = (((!g3464) & (g4799) & (!g2569)) + ((!g3464) & (g4799) & (g2569)) + ((g3464) & (!g4799) & (g2569)) + ((g3464) & (g4799) & (g2569)));
	assign g2570 = (((!g1179) & (!g1222) & (!g2456) & (!g2535) & (!g2458) & (!g2459)) + ((!g1179) & (!g1222) & (!g2456) & (!g2535) & (!g2458) & (g2459)) + ((!g1179) & (!g1222) & (!g2456) & (!g2535) & (g2458) & (!g2459)) + ((!g1179) & (!g1222) & (!g2456) & (!g2535) & (g2458) & (g2459)) + ((!g1179) & (!g1222) & (!g2456) & (g2535) & (!g2458) & (!g2459)) + ((!g1179) & (!g1222) & (!g2456) & (g2535) & (!g2458) & (g2459)) + ((!g1179) & (!g1222) & (!g2456) & (g2535) & (g2458) & (!g2459)) + ((!g1179) & (!g1222) & (!g2456) & (g2535) & (g2458) & (g2459)) + ((!g1179) & (!g1222) & (g2456) & (!g2535) & (!g2458) & (!g2459)) + ((!g1179) & (!g1222) & (g2456) & (!g2535) & (!g2458) & (g2459)) + ((!g1179) & (!g1222) & (g2456) & (!g2535) & (g2458) & (!g2459)) + ((!g1179) & (!g1222) & (g2456) & (!g2535) & (g2458) & (g2459)) + ((!g1179) & (!g1222) & (g2456) & (g2535) & (!g2458) & (!g2459)) + ((!g1179) & (g1222) & (!g2456) & (!g2535) & (!g2458) & (!g2459)) + ((!g1179) & (g1222) & (!g2456) & (!g2535) & (!g2458) & (g2459)) + ((!g1179) & (g1222) & (!g2456) & (!g2535) & (g2458) & (!g2459)) + ((!g1179) & (g1222) & (!g2456) & (!g2535) & (g2458) & (g2459)) + ((!g1179) & (g1222) & (g2456) & (!g2535) & (!g2458) & (!g2459)) + ((g1179) & (!g1222) & (!g2456) & (!g2535) & (!g2458) & (!g2459)) + ((g1179) & (!g1222) & (!g2456) & (!g2535) & (!g2458) & (g2459)) + ((g1179) & (!g1222) & (!g2456) & (!g2535) & (g2458) & (!g2459)) + ((g1179) & (!g1222) & (!g2456) & (!g2535) & (g2458) & (g2459)) + ((g1179) & (!g1222) & (!g2456) & (g2535) & (!g2458) & (!g2459)) + ((g1179) & (!g1222) & (g2456) & (!g2535) & (!g2458) & (!g2459)) + ((g1179) & (!g1222) & (g2456) & (!g2535) & (!g2458) & (g2459)) + ((g1179) & (!g1222) & (g2456) & (!g2535) & (g2458) & (!g2459)) + ((g1179) & (!g1222) & (g2456) & (!g2535) & (g2458) & (g2459)) + ((g1179) & (g1222) & (!g2456) & (!g2535) & (!g2458) & (!g2459)));
	assign g2571 = (((!g827) & (!g1249) & (g2569) & (!g2570)) + ((!g827) & (!g1249) & (g2569) & (g2570)) + ((!g827) & (g1249) & (g2569) & (!g2570)) + ((!g827) & (g1249) & (g2569) & (g2570)) + ((g827) & (!g1249) & (!g2569) & (!g2570)) + ((g827) & (!g1249) & (g2569) & (g2570)) + ((g827) & (g1249) & (!g2569) & (g2570)) + ((g827) & (g1249) & (g2569) & (!g2570)));
	assign g8050 = (((!g3499) & (g4802) & (!g2572)) + ((!g3499) & (g4802) & (g2572)) + ((g3499) & (!g4802) & (g2572)) + ((g3499) & (g4802) & (g2572)));
	assign g2573 = (((!g1181) & (!g1230) & (!g2462) & (!g2542) & (!g2464) & (!g2465)) + ((!g1181) & (!g1230) & (!g2462) & (!g2542) & (!g2464) & (g2465)) + ((!g1181) & (!g1230) & (!g2462) & (!g2542) & (g2464) & (!g2465)) + ((!g1181) & (!g1230) & (!g2462) & (!g2542) & (g2464) & (g2465)) + ((!g1181) & (!g1230) & (!g2462) & (g2542) & (!g2464) & (!g2465)) + ((!g1181) & (!g1230) & (!g2462) & (g2542) & (!g2464) & (g2465)) + ((!g1181) & (!g1230) & (!g2462) & (g2542) & (g2464) & (!g2465)) + ((!g1181) & (!g1230) & (!g2462) & (g2542) & (g2464) & (g2465)) + ((!g1181) & (!g1230) & (g2462) & (!g2542) & (!g2464) & (!g2465)) + ((!g1181) & (!g1230) & (g2462) & (!g2542) & (!g2464) & (g2465)) + ((!g1181) & (!g1230) & (g2462) & (!g2542) & (g2464) & (!g2465)) + ((!g1181) & (!g1230) & (g2462) & (!g2542) & (g2464) & (g2465)) + ((!g1181) & (!g1230) & (g2462) & (g2542) & (!g2464) & (!g2465)) + ((!g1181) & (g1230) & (!g2462) & (!g2542) & (!g2464) & (!g2465)) + ((!g1181) & (g1230) & (!g2462) & (!g2542) & (!g2464) & (g2465)) + ((!g1181) & (g1230) & (!g2462) & (!g2542) & (g2464) & (!g2465)) + ((!g1181) & (g1230) & (!g2462) & (!g2542) & (g2464) & (g2465)) + ((!g1181) & (g1230) & (g2462) & (!g2542) & (!g2464) & (!g2465)) + ((g1181) & (!g1230) & (!g2462) & (!g2542) & (!g2464) & (!g2465)) + ((g1181) & (!g1230) & (!g2462) & (!g2542) & (!g2464) & (g2465)) + ((g1181) & (!g1230) & (!g2462) & (!g2542) & (g2464) & (!g2465)) + ((g1181) & (!g1230) & (!g2462) & (!g2542) & (g2464) & (g2465)) + ((g1181) & (!g1230) & (!g2462) & (g2542) & (!g2464) & (!g2465)) + ((g1181) & (!g1230) & (g2462) & (!g2542) & (!g2464) & (!g2465)) + ((g1181) & (!g1230) & (g2462) & (!g2542) & (!g2464) & (g2465)) + ((g1181) & (!g1230) & (g2462) & (!g2542) & (g2464) & (!g2465)) + ((g1181) & (!g1230) & (g2462) & (!g2542) & (g2464) & (g2465)) + ((g1181) & (g1230) & (!g2462) & (!g2542) & (!g2464) & (!g2465)));
	assign g2574 = (((!g827) & (!g1251) & (g2572) & (!g2573)) + ((!g827) & (!g1251) & (g2572) & (g2573)) + ((!g827) & (g1251) & (g2572) & (!g2573)) + ((!g827) & (g1251) & (g2572) & (g2573)) + ((g827) & (!g1251) & (!g2572) & (!g2573)) + ((g827) & (!g1251) & (g2572) & (g2573)) + ((g827) & (g1251) & (!g2572) & (g2573)) + ((g827) & (g1251) & (g2572) & (!g2573)));
	assign g8051 = (((!g3464) & (g4805) & (!g2575)) + ((!g3464) & (g4805) & (g2575)) + ((g3464) & (!g4805) & (g2575)) + ((g3464) & (g4805) & (g2575)));
	assign g2576 = (((!g1183) & (!g1208) & (!g2468) & (!g2523) & (!g2470) & (!g2471)) + ((!g1183) & (!g1208) & (!g2468) & (!g2523) & (!g2470) & (g2471)) + ((!g1183) & (!g1208) & (!g2468) & (!g2523) & (g2470) & (!g2471)) + ((!g1183) & (!g1208) & (!g2468) & (!g2523) & (g2470) & (g2471)) + ((!g1183) & (!g1208) & (!g2468) & (g2523) & (!g2470) & (!g2471)) + ((!g1183) & (!g1208) & (!g2468) & (g2523) & (!g2470) & (g2471)) + ((!g1183) & (!g1208) & (!g2468) & (g2523) & (g2470) & (!g2471)) + ((!g1183) & (!g1208) & (!g2468) & (g2523) & (g2470) & (g2471)) + ((!g1183) & (!g1208) & (g2468) & (!g2523) & (!g2470) & (!g2471)) + ((!g1183) & (!g1208) & (g2468) & (!g2523) & (!g2470) & (g2471)) + ((!g1183) & (!g1208) & (g2468) & (!g2523) & (g2470) & (!g2471)) + ((!g1183) & (!g1208) & (g2468) & (!g2523) & (g2470) & (g2471)) + ((!g1183) & (!g1208) & (g2468) & (g2523) & (!g2470) & (!g2471)) + ((!g1183) & (g1208) & (!g2468) & (!g2523) & (!g2470) & (!g2471)) + ((!g1183) & (g1208) & (!g2468) & (!g2523) & (!g2470) & (g2471)) + ((!g1183) & (g1208) & (!g2468) & (!g2523) & (g2470) & (!g2471)) + ((!g1183) & (g1208) & (!g2468) & (!g2523) & (g2470) & (g2471)) + ((!g1183) & (g1208) & (g2468) & (!g2523) & (!g2470) & (!g2471)) + ((g1183) & (!g1208) & (!g2468) & (!g2523) & (!g2470) & (!g2471)) + ((g1183) & (!g1208) & (!g2468) & (!g2523) & (!g2470) & (g2471)) + ((g1183) & (!g1208) & (!g2468) & (!g2523) & (g2470) & (!g2471)) + ((g1183) & (!g1208) & (!g2468) & (!g2523) & (g2470) & (g2471)) + ((g1183) & (!g1208) & (!g2468) & (g2523) & (!g2470) & (!g2471)) + ((g1183) & (!g1208) & (g2468) & (!g2523) & (!g2470) & (!g2471)) + ((g1183) & (!g1208) & (g2468) & (!g2523) & (!g2470) & (g2471)) + ((g1183) & (!g1208) & (g2468) & (!g2523) & (g2470) & (!g2471)) + ((g1183) & (!g1208) & (g2468) & (!g2523) & (g2470) & (g2471)) + ((g1183) & (g1208) & (!g2468) & (!g2523) & (!g2470) & (!g2471)));
	assign g2577 = (((!g827) & (!g1253) & (g2575) & (!g2576)) + ((!g827) & (!g1253) & (g2575) & (g2576)) + ((!g827) & (g1253) & (g2575) & (!g2576)) + ((!g827) & (g1253) & (g2575) & (g2576)) + ((g827) & (!g1253) & (!g2575) & (!g2576)) + ((g827) & (!g1253) & (g2575) & (g2576)) + ((g827) & (g1253) & (!g2575) & (g2576)) + ((g827) & (g1253) & (g2575) & (!g2576)));
	assign g8052 = (((!g3499) & (g4808) & (!g2578)) + ((!g3499) & (g4808) & (g2578)) + ((g3499) & (!g4808) & (g2578)) + ((g3499) & (g4808) & (g2578)));
	assign g2579 = (((!g1185) & (!g1216) & (!g2474) & (!g2529) & (!g2476) & (!g2477)) + ((!g1185) & (!g1216) & (!g2474) & (!g2529) & (!g2476) & (g2477)) + ((!g1185) & (!g1216) & (!g2474) & (!g2529) & (g2476) & (!g2477)) + ((!g1185) & (!g1216) & (!g2474) & (!g2529) & (g2476) & (g2477)) + ((!g1185) & (!g1216) & (!g2474) & (g2529) & (!g2476) & (!g2477)) + ((!g1185) & (!g1216) & (!g2474) & (g2529) & (!g2476) & (g2477)) + ((!g1185) & (!g1216) & (!g2474) & (g2529) & (g2476) & (!g2477)) + ((!g1185) & (!g1216) & (!g2474) & (g2529) & (g2476) & (g2477)) + ((!g1185) & (!g1216) & (g2474) & (!g2529) & (!g2476) & (!g2477)) + ((!g1185) & (!g1216) & (g2474) & (!g2529) & (!g2476) & (g2477)) + ((!g1185) & (!g1216) & (g2474) & (!g2529) & (g2476) & (!g2477)) + ((!g1185) & (!g1216) & (g2474) & (!g2529) & (g2476) & (g2477)) + ((!g1185) & (!g1216) & (g2474) & (g2529) & (!g2476) & (!g2477)) + ((!g1185) & (g1216) & (!g2474) & (!g2529) & (!g2476) & (!g2477)) + ((!g1185) & (g1216) & (!g2474) & (!g2529) & (!g2476) & (g2477)) + ((!g1185) & (g1216) & (!g2474) & (!g2529) & (g2476) & (!g2477)) + ((!g1185) & (g1216) & (!g2474) & (!g2529) & (g2476) & (g2477)) + ((!g1185) & (g1216) & (g2474) & (!g2529) & (!g2476) & (!g2477)) + ((g1185) & (!g1216) & (!g2474) & (!g2529) & (!g2476) & (!g2477)) + ((g1185) & (!g1216) & (!g2474) & (!g2529) & (!g2476) & (g2477)) + ((g1185) & (!g1216) & (!g2474) & (!g2529) & (g2476) & (!g2477)) + ((g1185) & (!g1216) & (!g2474) & (!g2529) & (g2476) & (g2477)) + ((g1185) & (!g1216) & (!g2474) & (g2529) & (!g2476) & (!g2477)) + ((g1185) & (!g1216) & (g2474) & (!g2529) & (!g2476) & (!g2477)) + ((g1185) & (!g1216) & (g2474) & (!g2529) & (!g2476) & (g2477)) + ((g1185) & (!g1216) & (g2474) & (!g2529) & (g2476) & (!g2477)) + ((g1185) & (!g1216) & (g2474) & (!g2529) & (g2476) & (g2477)) + ((g1185) & (g1216) & (!g2474) & (!g2529) & (!g2476) & (!g2477)));
	assign g2580 = (((!g827) & (!g1255) & (g2578) & (!g2579)) + ((!g827) & (!g1255) & (g2578) & (g2579)) + ((!g827) & (g1255) & (g2578) & (!g2579)) + ((!g827) & (g1255) & (g2578) & (g2579)) + ((g827) & (!g1255) & (!g2578) & (!g2579)) + ((g827) & (!g1255) & (g2578) & (g2579)) + ((g827) & (g1255) & (!g2578) & (g2579)) + ((g827) & (g1255) & (g2578) & (!g2579)));
	assign g8053 = (((!g2017) & (g4811) & (!g2581)) + ((!g2017) & (g4811) & (g2581)) + ((g2017) & (!g4811) & (g2581)) + ((g2017) & (g4811) & (g2581)));
	assign g2582 = (((!g1187) & (!g1224) & (!g2480) & (!g2537) & (!g2482) & (!g2483)) + ((!g1187) & (!g1224) & (!g2480) & (!g2537) & (!g2482) & (g2483)) + ((!g1187) & (!g1224) & (!g2480) & (!g2537) & (g2482) & (!g2483)) + ((!g1187) & (!g1224) & (!g2480) & (!g2537) & (g2482) & (g2483)) + ((!g1187) & (!g1224) & (!g2480) & (g2537) & (!g2482) & (!g2483)) + ((!g1187) & (!g1224) & (!g2480) & (g2537) & (!g2482) & (g2483)) + ((!g1187) & (!g1224) & (!g2480) & (g2537) & (g2482) & (!g2483)) + ((!g1187) & (!g1224) & (!g2480) & (g2537) & (g2482) & (g2483)) + ((!g1187) & (!g1224) & (g2480) & (!g2537) & (!g2482) & (!g2483)) + ((!g1187) & (!g1224) & (g2480) & (!g2537) & (!g2482) & (g2483)) + ((!g1187) & (!g1224) & (g2480) & (!g2537) & (g2482) & (!g2483)) + ((!g1187) & (!g1224) & (g2480) & (!g2537) & (g2482) & (g2483)) + ((!g1187) & (!g1224) & (g2480) & (g2537) & (!g2482) & (!g2483)) + ((!g1187) & (g1224) & (!g2480) & (!g2537) & (!g2482) & (!g2483)) + ((!g1187) & (g1224) & (!g2480) & (!g2537) & (!g2482) & (g2483)) + ((!g1187) & (g1224) & (!g2480) & (!g2537) & (g2482) & (!g2483)) + ((!g1187) & (g1224) & (!g2480) & (!g2537) & (g2482) & (g2483)) + ((!g1187) & (g1224) & (g2480) & (!g2537) & (!g2482) & (!g2483)) + ((g1187) & (!g1224) & (!g2480) & (!g2537) & (!g2482) & (!g2483)) + ((g1187) & (!g1224) & (!g2480) & (!g2537) & (!g2482) & (g2483)) + ((g1187) & (!g1224) & (!g2480) & (!g2537) & (g2482) & (!g2483)) + ((g1187) & (!g1224) & (!g2480) & (!g2537) & (g2482) & (g2483)) + ((g1187) & (!g1224) & (!g2480) & (g2537) & (!g2482) & (!g2483)) + ((g1187) & (!g1224) & (g2480) & (!g2537) & (!g2482) & (!g2483)) + ((g1187) & (!g1224) & (g2480) & (!g2537) & (!g2482) & (g2483)) + ((g1187) & (!g1224) & (g2480) & (!g2537) & (g2482) & (!g2483)) + ((g1187) & (!g1224) & (g2480) & (!g2537) & (g2482) & (g2483)) + ((g1187) & (g1224) & (!g2480) & (!g2537) & (!g2482) & (!g2483)));
	assign g2583 = (((!g827) & (!g1257) & (g2581) & (!g2582)) + ((!g827) & (!g1257) & (g2581) & (g2582)) + ((!g827) & (g1257) & (g2581) & (!g2582)) + ((!g827) & (g1257) & (g2581) & (g2582)) + ((g827) & (!g1257) & (!g2581) & (!g2582)) + ((g827) & (!g1257) & (g2581) & (g2582)) + ((g827) & (g1257) & (!g2581) & (g2582)) + ((g827) & (g1257) & (g2581) & (!g2582)));
	assign g8054 = (((!g3429) & (g4816) & (!g2584)) + ((!g3429) & (g4816) & (g2584)) + ((g3429) & (!g4816) & (g2584)) + ((g3429) & (g4816) & (g2584)));
	assign g2585 = (((!g1189) & (!g1232) & (!g2486) & (!g2544) & (!g2488) & (!g2489)) + ((!g1189) & (!g1232) & (!g2486) & (!g2544) & (!g2488) & (g2489)) + ((!g1189) & (!g1232) & (!g2486) & (!g2544) & (g2488) & (!g2489)) + ((!g1189) & (!g1232) & (!g2486) & (!g2544) & (g2488) & (g2489)) + ((!g1189) & (!g1232) & (!g2486) & (g2544) & (!g2488) & (!g2489)) + ((!g1189) & (!g1232) & (!g2486) & (g2544) & (!g2488) & (g2489)) + ((!g1189) & (!g1232) & (!g2486) & (g2544) & (g2488) & (!g2489)) + ((!g1189) & (!g1232) & (!g2486) & (g2544) & (g2488) & (g2489)) + ((!g1189) & (!g1232) & (g2486) & (!g2544) & (!g2488) & (!g2489)) + ((!g1189) & (!g1232) & (g2486) & (!g2544) & (!g2488) & (g2489)) + ((!g1189) & (!g1232) & (g2486) & (!g2544) & (g2488) & (!g2489)) + ((!g1189) & (!g1232) & (g2486) & (!g2544) & (g2488) & (g2489)) + ((!g1189) & (!g1232) & (g2486) & (g2544) & (!g2488) & (!g2489)) + ((!g1189) & (g1232) & (!g2486) & (!g2544) & (!g2488) & (!g2489)) + ((!g1189) & (g1232) & (!g2486) & (!g2544) & (!g2488) & (g2489)) + ((!g1189) & (g1232) & (!g2486) & (!g2544) & (g2488) & (!g2489)) + ((!g1189) & (g1232) & (!g2486) & (!g2544) & (g2488) & (g2489)) + ((!g1189) & (g1232) & (g2486) & (!g2544) & (!g2488) & (!g2489)) + ((g1189) & (!g1232) & (!g2486) & (!g2544) & (!g2488) & (!g2489)) + ((g1189) & (!g1232) & (!g2486) & (!g2544) & (!g2488) & (g2489)) + ((g1189) & (!g1232) & (!g2486) & (!g2544) & (g2488) & (!g2489)) + ((g1189) & (!g1232) & (!g2486) & (!g2544) & (g2488) & (g2489)) + ((g1189) & (!g1232) & (!g2486) & (g2544) & (!g2488) & (!g2489)) + ((g1189) & (!g1232) & (g2486) & (!g2544) & (!g2488) & (!g2489)) + ((g1189) & (!g1232) & (g2486) & (!g2544) & (!g2488) & (g2489)) + ((g1189) & (!g1232) & (g2486) & (!g2544) & (g2488) & (!g2489)) + ((g1189) & (!g1232) & (g2486) & (!g2544) & (g2488) & (g2489)) + ((g1189) & (g1232) & (!g2486) & (!g2544) & (!g2488) & (!g2489)));
	assign g2586 = (((!g827) & (!g1259) & (g2584) & (!g2585)) + ((!g827) & (!g1259) & (g2584) & (g2585)) + ((!g827) & (g1259) & (g2584) & (!g2585)) + ((!g827) & (g1259) & (g2584) & (g2585)) + ((g827) & (!g1259) & (!g2584) & (!g2585)) + ((g827) & (!g1259) & (g2584) & (g2585)) + ((g827) & (g1259) & (!g2584) & (g2585)) + ((g827) & (g1259) & (g2584) & (!g2585)));
	assign g2587 = (((!g1191) & (!g1210) & (!g2004) & (!g2006) & (!g2493) & (!g2494)) + ((!g1191) & (!g1210) & (!g2004) & (!g2006) & (!g2493) & (g2494)) + ((!g1191) & (!g1210) & (!g2004) & (!g2006) & (g2493) & (!g2494)) + ((!g1191) & (!g1210) & (!g2004) & (!g2006) & (g2493) & (g2494)) + ((!g1191) & (!g1210) & (!g2004) & (g2006) & (!g2493) & (!g2494)) + ((!g1191) & (!g1210) & (!g2004) & (g2006) & (!g2493) & (g2494)) + ((!g1191) & (!g1210) & (!g2004) & (g2006) & (g2493) & (!g2494)) + ((!g1191) & (!g1210) & (!g2004) & (g2006) & (g2493) & (g2494)) + ((!g1191) & (!g1210) & (g2004) & (!g2006) & (!g2493) & (!g2494)) + ((!g1191) & (!g1210) & (g2004) & (!g2006) & (!g2493) & (g2494)) + ((!g1191) & (!g1210) & (g2004) & (!g2006) & (g2493) & (!g2494)) + ((!g1191) & (!g1210) & (g2004) & (!g2006) & (g2493) & (g2494)) + ((!g1191) & (!g1210) & (g2004) & (g2006) & (!g2493) & (!g2494)) + ((!g1191) & (g1210) & (!g2004) & (!g2006) & (!g2493) & (!g2494)) + ((!g1191) & (g1210) & (!g2004) & (!g2006) & (!g2493) & (g2494)) + ((!g1191) & (g1210) & (!g2004) & (!g2006) & (g2493) & (!g2494)) + ((!g1191) & (g1210) & (!g2004) & (!g2006) & (g2493) & (g2494)) + ((!g1191) & (g1210) & (g2004) & (!g2006) & (!g2493) & (!g2494)) + ((g1191) & (!g1210) & (!g2004) & (!g2006) & (!g2493) & (!g2494)) + ((g1191) & (!g1210) & (!g2004) & (!g2006) & (!g2493) & (g2494)) + ((g1191) & (!g1210) & (!g2004) & (!g2006) & (g2493) & (!g2494)) + ((g1191) & (!g1210) & (!g2004) & (!g2006) & (g2493) & (g2494)) + ((g1191) & (!g1210) & (!g2004) & (g2006) & (!g2493) & (!g2494)) + ((g1191) & (!g1210) & (g2004) & (!g2006) & (!g2493) & (!g2494)) + ((g1191) & (!g1210) & (g2004) & (!g2006) & (!g2493) & (g2494)) + ((g1191) & (!g1210) & (g2004) & (!g2006) & (g2493) & (!g2494)) + ((g1191) & (!g1210) & (g2004) & (!g2006) & (g2493) & (g2494)) + ((g1191) & (g1210) & (!g2004) & (!g2006) & (!g2493) & (!g2494)));
	assign g2588 = (((!g827) & (!g1261) & (g2012) & (!g2587)) + ((!g827) & (!g1261) & (g2012) & (g2587)) + ((!g827) & (g1261) & (g2012) & (!g2587)) + ((!g827) & (g1261) & (g2012) & (g2587)) + ((g827) & (!g1261) & (!g2012) & (!g2587)) + ((g827) & (!g1261) & (g2012) & (g2587)) + ((g827) & (g1261) & (!g2012) & (g2587)) + ((g827) & (g1261) & (g2012) & (!g2587)));
	assign g8055 = (((!g3464) & (g4819) & (!g2589)) + ((!g3464) & (g4819) & (g2589)) + ((g3464) & (!g4819) & (g2589)) + ((g3464) & (g4819) & (g2589)));
	assign g2590 = (((!g1193) & (!g1218) & (!g2497) & (!g2531) & (!g2499) & (!g2500)) + ((!g1193) & (!g1218) & (!g2497) & (!g2531) & (!g2499) & (g2500)) + ((!g1193) & (!g1218) & (!g2497) & (!g2531) & (g2499) & (!g2500)) + ((!g1193) & (!g1218) & (!g2497) & (!g2531) & (g2499) & (g2500)) + ((!g1193) & (!g1218) & (!g2497) & (g2531) & (!g2499) & (!g2500)) + ((!g1193) & (!g1218) & (!g2497) & (g2531) & (!g2499) & (g2500)) + ((!g1193) & (!g1218) & (!g2497) & (g2531) & (g2499) & (!g2500)) + ((!g1193) & (!g1218) & (!g2497) & (g2531) & (g2499) & (g2500)) + ((!g1193) & (!g1218) & (g2497) & (!g2531) & (!g2499) & (!g2500)) + ((!g1193) & (!g1218) & (g2497) & (!g2531) & (!g2499) & (g2500)) + ((!g1193) & (!g1218) & (g2497) & (!g2531) & (g2499) & (!g2500)) + ((!g1193) & (!g1218) & (g2497) & (!g2531) & (g2499) & (g2500)) + ((!g1193) & (!g1218) & (g2497) & (g2531) & (!g2499) & (!g2500)) + ((!g1193) & (g1218) & (!g2497) & (!g2531) & (!g2499) & (!g2500)) + ((!g1193) & (g1218) & (!g2497) & (!g2531) & (!g2499) & (g2500)) + ((!g1193) & (g1218) & (!g2497) & (!g2531) & (g2499) & (!g2500)) + ((!g1193) & (g1218) & (!g2497) & (!g2531) & (g2499) & (g2500)) + ((!g1193) & (g1218) & (g2497) & (!g2531) & (!g2499) & (!g2500)) + ((g1193) & (!g1218) & (!g2497) & (!g2531) & (!g2499) & (!g2500)) + ((g1193) & (!g1218) & (!g2497) & (!g2531) & (!g2499) & (g2500)) + ((g1193) & (!g1218) & (!g2497) & (!g2531) & (g2499) & (!g2500)) + ((g1193) & (!g1218) & (!g2497) & (!g2531) & (g2499) & (g2500)) + ((g1193) & (!g1218) & (!g2497) & (g2531) & (!g2499) & (!g2500)) + ((g1193) & (!g1218) & (g2497) & (!g2531) & (!g2499) & (!g2500)) + ((g1193) & (!g1218) & (g2497) & (!g2531) & (!g2499) & (g2500)) + ((g1193) & (!g1218) & (g2497) & (!g2531) & (g2499) & (!g2500)) + ((g1193) & (!g1218) & (g2497) & (!g2531) & (g2499) & (g2500)) + ((g1193) & (g1218) & (!g2497) & (!g2531) & (!g2499) & (!g2500)));
	assign g2591 = (((!g827) & (!g1263) & (g2589) & (!g2590)) + ((!g827) & (!g1263) & (g2589) & (g2590)) + ((!g827) & (g1263) & (g2589) & (!g2590)) + ((!g827) & (g1263) & (g2589) & (g2590)) + ((g827) & (!g1263) & (!g2589) & (!g2590)) + ((g827) & (!g1263) & (g2589) & (g2590)) + ((g827) & (g1263) & (!g2589) & (g2590)) + ((g827) & (g1263) & (g2589) & (!g2590)));
	assign g8056 = (((!g3429) & (g4824) & (!g2592)) + ((!g3429) & (g4824) & (g2592)) + ((g3429) & (!g4824) & (g2592)) + ((g3429) & (g4824) & (g2592)));
	assign g2593 = (((!g1195) & (!g1226) & (!g2503) & (!g2539) & (!g2505) & (!g2506)) + ((!g1195) & (!g1226) & (!g2503) & (!g2539) & (!g2505) & (g2506)) + ((!g1195) & (!g1226) & (!g2503) & (!g2539) & (g2505) & (!g2506)) + ((!g1195) & (!g1226) & (!g2503) & (!g2539) & (g2505) & (g2506)) + ((!g1195) & (!g1226) & (!g2503) & (g2539) & (!g2505) & (!g2506)) + ((!g1195) & (!g1226) & (!g2503) & (g2539) & (!g2505) & (g2506)) + ((!g1195) & (!g1226) & (!g2503) & (g2539) & (g2505) & (!g2506)) + ((!g1195) & (!g1226) & (!g2503) & (g2539) & (g2505) & (g2506)) + ((!g1195) & (!g1226) & (g2503) & (!g2539) & (!g2505) & (!g2506)) + ((!g1195) & (!g1226) & (g2503) & (!g2539) & (!g2505) & (g2506)) + ((!g1195) & (!g1226) & (g2503) & (!g2539) & (g2505) & (!g2506)) + ((!g1195) & (!g1226) & (g2503) & (!g2539) & (g2505) & (g2506)) + ((!g1195) & (!g1226) & (g2503) & (g2539) & (!g2505) & (!g2506)) + ((!g1195) & (g1226) & (!g2503) & (!g2539) & (!g2505) & (!g2506)) + ((!g1195) & (g1226) & (!g2503) & (!g2539) & (!g2505) & (g2506)) + ((!g1195) & (g1226) & (!g2503) & (!g2539) & (g2505) & (!g2506)) + ((!g1195) & (g1226) & (!g2503) & (!g2539) & (g2505) & (g2506)) + ((!g1195) & (g1226) & (g2503) & (!g2539) & (!g2505) & (!g2506)) + ((g1195) & (!g1226) & (!g2503) & (!g2539) & (!g2505) & (!g2506)) + ((g1195) & (!g1226) & (!g2503) & (!g2539) & (!g2505) & (g2506)) + ((g1195) & (!g1226) & (!g2503) & (!g2539) & (g2505) & (!g2506)) + ((g1195) & (!g1226) & (!g2503) & (!g2539) & (g2505) & (g2506)) + ((g1195) & (!g1226) & (!g2503) & (g2539) & (!g2505) & (!g2506)) + ((g1195) & (!g1226) & (g2503) & (!g2539) & (!g2505) & (!g2506)) + ((g1195) & (!g1226) & (g2503) & (!g2539) & (!g2505) & (g2506)) + ((g1195) & (!g1226) & (g2503) & (!g2539) & (g2505) & (!g2506)) + ((g1195) & (!g1226) & (g2503) & (!g2539) & (g2505) & (g2506)) + ((g1195) & (g1226) & (!g2503) & (!g2539) & (!g2505) & (!g2506)));
	assign g2594 = (((!g827) & (!g1265) & (g2592) & (!g2593)) + ((!g827) & (!g1265) & (g2592) & (g2593)) + ((!g827) & (g1265) & (g2592) & (!g2593)) + ((!g827) & (g1265) & (g2592) & (g2593)) + ((g827) & (!g1265) & (!g2592) & (!g2593)) + ((g827) & (!g1265) & (g2592) & (g2593)) + ((g827) & (g1265) & (!g2592) & (g2593)) + ((g827) & (g1265) & (g2592) & (!g2593)));
	assign g8057 = (((!g2017) & (g4827) & (!g2595)) + ((!g2017) & (g4827) & (g2595)) + ((g2017) & (!g4827) & (g2595)) + ((g2017) & (g4827) & (g2595)));
	assign g2596 = (((!g1197) & (!g1234) & (!g2509) & (!g2546) & (!g2511) & (!g2512)) + ((!g1197) & (!g1234) & (!g2509) & (!g2546) & (!g2511) & (g2512)) + ((!g1197) & (!g1234) & (!g2509) & (!g2546) & (g2511) & (!g2512)) + ((!g1197) & (!g1234) & (!g2509) & (!g2546) & (g2511) & (g2512)) + ((!g1197) & (!g1234) & (!g2509) & (g2546) & (!g2511) & (!g2512)) + ((!g1197) & (!g1234) & (!g2509) & (g2546) & (!g2511) & (g2512)) + ((!g1197) & (!g1234) & (!g2509) & (g2546) & (g2511) & (!g2512)) + ((!g1197) & (!g1234) & (!g2509) & (g2546) & (g2511) & (g2512)) + ((!g1197) & (!g1234) & (g2509) & (!g2546) & (!g2511) & (!g2512)) + ((!g1197) & (!g1234) & (g2509) & (!g2546) & (!g2511) & (g2512)) + ((!g1197) & (!g1234) & (g2509) & (!g2546) & (g2511) & (!g2512)) + ((!g1197) & (!g1234) & (g2509) & (!g2546) & (g2511) & (g2512)) + ((!g1197) & (!g1234) & (g2509) & (g2546) & (!g2511) & (!g2512)) + ((!g1197) & (g1234) & (!g2509) & (!g2546) & (!g2511) & (!g2512)) + ((!g1197) & (g1234) & (!g2509) & (!g2546) & (!g2511) & (g2512)) + ((!g1197) & (g1234) & (!g2509) & (!g2546) & (g2511) & (!g2512)) + ((!g1197) & (g1234) & (!g2509) & (!g2546) & (g2511) & (g2512)) + ((!g1197) & (g1234) & (g2509) & (!g2546) & (!g2511) & (!g2512)) + ((g1197) & (!g1234) & (!g2509) & (!g2546) & (!g2511) & (!g2512)) + ((g1197) & (!g1234) & (!g2509) & (!g2546) & (!g2511) & (g2512)) + ((g1197) & (!g1234) & (!g2509) & (!g2546) & (g2511) & (!g2512)) + ((g1197) & (!g1234) & (!g2509) & (!g2546) & (g2511) & (g2512)) + ((g1197) & (!g1234) & (!g2509) & (g2546) & (!g2511) & (!g2512)) + ((g1197) & (!g1234) & (g2509) & (!g2546) & (!g2511) & (!g2512)) + ((g1197) & (!g1234) & (g2509) & (!g2546) & (!g2511) & (g2512)) + ((g1197) & (!g1234) & (g2509) & (!g2546) & (g2511) & (!g2512)) + ((g1197) & (!g1234) & (g2509) & (!g2546) & (g2511) & (g2512)) + ((g1197) & (g1234) & (!g2509) & (!g2546) & (!g2511) & (!g2512)));
	assign g2597 = (((!g827) & (!g1267) & (g2595) & (!g2596)) + ((!g827) & (!g1267) & (g2595) & (g2596)) + ((!g827) & (g1267) & (g2595) & (!g2596)) + ((!g827) & (g1267) & (g2595) & (g2596)) + ((g827) & (!g1267) & (!g2595) & (!g2596)) + ((g827) & (!g1267) & (g2595) & (g2596)) + ((g827) & (g1267) & (!g2595) & (g2596)) + ((g827) & (g1267) & (g2595) & (!g2596)));
	assign g8058 = (((!g3429) & (g4830) & (!g2598)) + ((!g3429) & (g4830) & (g2598)) + ((g3429) & (!g4830) & (g2598)) + ((g3429) & (g4830) & (g2598)));
	assign g8059 = (((!g3464) & (g4832) & (!g2599)) + ((!g3464) & (g4832) & (g2599)) + ((g3464) & (!g4832) & (g2599)) + ((g3464) & (g4832) & (g2599)));
	assign g2600 = (((!g2549) & (!g2550) & (!g2551) & (!g2552) & (!g2598) & (g2599)) + ((!g2549) & (!g2550) & (!g2551) & (!g2552) & (g2598) & (!g2599)) + ((!g2549) & (!g2550) & (!g2551) & (g2552) & (!g2598) & (g2599)) + ((!g2549) & (!g2550) & (!g2551) & (g2552) & (g2598) & (!g2599)) + ((!g2549) & (!g2550) & (g2551) & (!g2552) & (!g2598) & (g2599)) + ((!g2549) & (!g2550) & (g2551) & (!g2552) & (g2598) & (!g2599)) + ((!g2549) & (!g2550) & (g2551) & (g2552) & (!g2598) & (!g2599)) + ((!g2549) & (!g2550) & (g2551) & (g2552) & (g2598) & (g2599)) + ((!g2549) & (g2550) & (!g2551) & (!g2552) & (!g2598) & (g2599)) + ((!g2549) & (g2550) & (!g2551) & (!g2552) & (g2598) & (!g2599)) + ((!g2549) & (g2550) & (!g2551) & (g2552) & (!g2598) & (!g2599)) + ((!g2549) & (g2550) & (!g2551) & (g2552) & (g2598) & (g2599)) + ((!g2549) & (g2550) & (g2551) & (!g2552) & (!g2598) & (!g2599)) + ((!g2549) & (g2550) & (g2551) & (!g2552) & (g2598) & (g2599)) + ((!g2549) & (g2550) & (g2551) & (g2552) & (!g2598) & (!g2599)) + ((!g2549) & (g2550) & (g2551) & (g2552) & (g2598) & (g2599)) + ((g2549) & (!g2550) & (!g2551) & (!g2552) & (!g2598) & (g2599)) + ((g2549) & (!g2550) & (!g2551) & (!g2552) & (g2598) & (!g2599)) + ((g2549) & (!g2550) & (!g2551) & (g2552) & (!g2598) & (!g2599)) + ((g2549) & (!g2550) & (!g2551) & (g2552) & (g2598) & (g2599)) + ((g2549) & (!g2550) & (g2551) & (!g2552) & (!g2598) & (!g2599)) + ((g2549) & (!g2550) & (g2551) & (!g2552) & (g2598) & (g2599)) + ((g2549) & (!g2550) & (g2551) & (g2552) & (!g2598) & (!g2599)) + ((g2549) & (!g2550) & (g2551) & (g2552) & (g2598) & (g2599)) + ((g2549) & (g2550) & (!g2551) & (!g2552) & (!g2598) & (g2599)) + ((g2549) & (g2550) & (!g2551) & (!g2552) & (g2598) & (!g2599)) + ((g2549) & (g2550) & (!g2551) & (g2552) & (!g2598) & (!g2599)) + ((g2549) & (g2550) & (!g2551) & (g2552) & (g2598) & (g2599)) + ((g2549) & (g2550) & (g2551) & (!g2552) & (!g2598) & (!g2599)) + ((g2549) & (g2550) & (g2551) & (!g2552) & (g2598) & (g2599)) + ((g2549) & (g2550) & (g2551) & (g2552) & (!g2598) & (!g2599)) + ((g2549) & (g2550) & (g2551) & (g2552) & (g2598) & (g2599)));
	assign g8060 = (((!g3429) & (g4836) & (!g2601)) + ((!g3429) & (g4836) & (g2601)) + ((g3429) & (!g4836) & (g2601)) + ((g3429) & (g4836) & (g2601)));
	assign g8061 = (((!g3499) & (g4838) & (!g2602)) + ((!g3499) & (g4838) & (g2602)) + ((g3499) & (!g4838) & (g2602)) + ((g3499) & (g4838) & (g2602)));
	assign g2603 = (((!g2554) & (!g2555) & (!g2556) & (!g2601) & (g2602)) + ((!g2554) & (!g2555) & (!g2556) & (g2601) & (!g2602)) + ((!g2554) & (!g2555) & (g2556) & (!g2601) & (g2602)) + ((!g2554) & (!g2555) & (g2556) & (g2601) & (!g2602)) + ((!g2554) & (g2555) & (!g2556) & (!g2601) & (g2602)) + ((!g2554) & (g2555) & (!g2556) & (g2601) & (!g2602)) + ((!g2554) & (g2555) & (g2556) & (!g2601) & (!g2602)) + ((!g2554) & (g2555) & (g2556) & (g2601) & (g2602)) + ((g2554) & (!g2555) & (!g2556) & (!g2601) & (g2602)) + ((g2554) & (!g2555) & (!g2556) & (g2601) & (!g2602)) + ((g2554) & (!g2555) & (g2556) & (!g2601) & (!g2602)) + ((g2554) & (!g2555) & (g2556) & (g2601) & (g2602)) + ((g2554) & (g2555) & (!g2556) & (!g2601) & (!g2602)) + ((g2554) & (g2555) & (!g2556) & (g2601) & (g2602)) + ((g2554) & (g2555) & (g2556) & (!g2601) & (!g2602)) + ((g2554) & (g2555) & (g2556) & (g2601) & (g2602)));
	assign g2604 = (((!g830) & (!g1914) & (!g2600) & (!g2603) & (!g1269)) + ((!g830) & (!g1914) & (!g2600) & (!g2603) & (g1269)) + ((!g830) & (!g1914) & (!g2600) & (g2603) & (!g1269)) + ((!g830) & (!g1914) & (!g2600) & (g2603) & (g1269)) + ((!g830) & (!g1914) & (g2600) & (!g2603) & (!g1269)) + ((!g830) & (!g1914) & (g2600) & (!g2603) & (g1269)) + ((!g830) & (!g1914) & (g2600) & (g2603) & (!g1269)) + ((!g830) & (!g1914) & (g2600) & (g2603) & (g1269)) + ((!g830) & (g1914) & (!g2600) & (!g2603) & (!g1269)) + ((!g830) & (g1914) & (!g2600) & (!g2603) & (g1269)) + ((!g830) & (g1914) & (!g2600) & (g2603) & (!g1269)) + ((!g830) & (g1914) & (!g2600) & (g2603) & (g1269)) + ((!g830) & (g1914) & (g2600) & (!g2603) & (!g1269)) + ((!g830) & (g1914) & (g2600) & (!g2603) & (g1269)) + ((!g830) & (g1914) & (g2600) & (g2603) & (!g1269)) + ((!g830) & (g1914) & (g2600) & (g2603) & (g1269)) + ((g830) & (!g1914) & (!g2600) & (!g2603) & (g1269)) + ((g830) & (!g1914) & (!g2600) & (g2603) & (!g1269)) + ((g830) & (!g1914) & (g2600) & (!g2603) & (g1269)) + ((g830) & (!g1914) & (g2600) & (g2603) & (!g1269)) + ((g830) & (g1914) & (!g2600) & (!g2603) & (g1269)) + ((g830) & (g1914) & (!g2600) & (g2603) & (g1269)) + ((g830) & (g1914) & (g2600) & (!g2603) & (!g1269)) + ((g830) & (g1914) & (g2600) & (g2603) & (!g1269)));
	assign g2605 = (((!g1245) & (g2011) & (!g2564)) + ((g1245) & (!g2011) & (!g2564)) + ((g1245) & (g2011) & (!g2564)) + ((g1245) & (g2011) & (g2564)));
	assign g2606 = (((!g827) & (!g1273) & (g2013) & (!g2605)) + ((!g827) & (!g1273) & (g2013) & (g2605)) + ((!g827) & (g1273) & (g2013) & (!g2605)) + ((!g827) & (g1273) & (g2013) & (g2605)) + ((g827) & (!g1273) & (!g2013) & (g2605)) + ((g827) & (!g1273) & (g2013) & (!g2605)) + ((g827) & (g1273) & (!g2013) & (!g2605)) + ((g827) & (g1273) & (g2013) & (g2605)));
	assign g8062 = (((!g3464) & (g4840) & (!g2607)) + ((!g3464) & (g4840) & (g2607)) + ((g3464) & (!g4840) & (g2607)) + ((g3464) & (g4840) & (g2607)));
	assign g2608 = (((!g1253) & (g2575) & (!g2576)) + ((g1253) & (!g2575) & (!g2576)) + ((g1253) & (g2575) & (!g2576)) + ((g1253) & (g2575) & (g2576)));
	assign g2609 = (((!g827) & (!g1275) & (g2607) & (!g2608)) + ((!g827) & (!g1275) & (g2607) & (g2608)) + ((!g827) & (g1275) & (g2607) & (!g2608)) + ((!g827) & (g1275) & (g2607) & (g2608)) + ((g827) & (!g1275) & (!g2607) & (g2608)) + ((g827) & (!g1275) & (g2607) & (!g2608)) + ((g827) & (g1275) & (!g2607) & (!g2608)) + ((g827) & (g1275) & (g2607) & (g2608)));
	assign g2610 = (((!g1261) & (g2012) & (!g2587)) + ((g1261) & (!g2012) & (!g2587)) + ((g1261) & (g2012) & (!g2587)) + ((g1261) & (g2012) & (g2587)));
	assign g2611 = (((!g827) & (!g1277) & (g2014) & (!g2610)) + ((!g827) & (!g1277) & (g2014) & (g2610)) + ((!g827) & (g1277) & (g2014) & (!g2610)) + ((!g827) & (g1277) & (g2014) & (g2610)) + ((g827) & (!g1277) & (!g2014) & (g2610)) + ((g827) & (!g1277) & (g2014) & (!g2610)) + ((g827) & (g1277) & (!g2014) & (!g2610)) + ((g827) & (g1277) & (g2014) & (g2610)));
	assign g2612 = (((!g1239) & (g1972) & (!g2557)) + ((g1239) & (!g1972) & (!g2557)) + ((g1239) & (g1972) & (!g2557)) + ((g1239) & (g1972) & (g2557)));
	assign g2613 = (((!g827) & (!g1279) & (g1975) & (!g2612)) + ((!g827) & (!g1279) & (g1975) & (g2612)) + ((!g827) & (g1279) & (g1975) & (!g2612)) + ((!g827) & (g1279) & (g1975) & (g2612)) + ((g827) & (!g1279) & (!g1975) & (g2612)) + ((g827) & (!g1279) & (g1975) & (!g2612)) + ((g827) & (g1279) & (!g1975) & (!g2612)) + ((g827) & (g1279) & (g1975) & (g2612)));
	assign g8063 = (((!g2017) & (g6403) & (!g2614)) + ((!g2017) & (g6403) & (g2614)) + ((g2017) & (!g6403) & (g2614)) + ((g2017) & (g6403) & (g2614)));
	assign g2615 = (((!g1247) & (g2566) & (!g2567)) + ((g1247) & (!g2566) & (!g2567)) + ((g1247) & (g2566) & (!g2567)) + ((g1247) & (g2566) & (g2567)));
	assign g2616 = (((!g827) & (!g1281) & (g2614) & (!g2615)) + ((!g827) & (!g1281) & (g2614) & (g2615)) + ((!g827) & (g1281) & (g2614) & (!g2615)) + ((!g827) & (g1281) & (g2614) & (g2615)) + ((g827) & (!g1281) & (!g2614) & (g2615)) + ((g827) & (!g1281) & (g2614) & (!g2615)) + ((g827) & (g1281) & (!g2614) & (!g2615)) + ((g827) & (g1281) & (g2614) & (g2615)));
	assign g8064 = (((!g3499) & (g4844) & (!g2617)) + ((!g3499) & (g4844) & (g2617)) + ((g3499) & (!g4844) & (g2617)) + ((g3499) & (g4844) & (g2617)));
	assign g2618 = (((!g1255) & (g2578) & (!g2579)) + ((g1255) & (!g2578) & (!g2579)) + ((g1255) & (g2578) & (!g2579)) + ((g1255) & (g2578) & (g2579)));
	assign g2619 = (((!g827) & (!g1283) & (g2617) & (!g2618)) + ((!g827) & (!g1283) & (g2617) & (g2618)) + ((!g827) & (g1283) & (g2617) & (!g2618)) + ((!g827) & (g1283) & (g2617) & (g2618)) + ((g827) & (!g1283) & (!g2617) & (g2618)) + ((g827) & (!g1283) & (g2617) & (!g2618)) + ((g827) & (g1283) & (!g2617) & (!g2618)) + ((g827) & (g1283) & (g2617) & (g2618)));
	assign g8065 = (((!g3464) & (g4846) & (!g2620)) + ((!g3464) & (g4846) & (g2620)) + ((g3464) & (!g4846) & (g2620)) + ((g3464) & (g4846) & (g2620)));
	assign g2621 = (((!g1263) & (g2589) & (!g2590)) + ((g1263) & (!g2589) & (!g2590)) + ((g1263) & (g2589) & (!g2590)) + ((g1263) & (g2589) & (g2590)));
	assign g2622 = (((!g827) & (!g1285) & (g2620) & (!g2621)) + ((!g827) & (!g1285) & (g2620) & (g2621)) + ((!g827) & (g1285) & (g2620) & (!g2621)) + ((!g827) & (g1285) & (g2620) & (g2621)) + ((g827) & (!g1285) & (!g2620) & (g2621)) + ((g827) & (!g1285) & (g2620) & (!g2621)) + ((g827) & (g1285) & (!g2620) & (!g2621)) + ((g827) & (g1285) & (g2620) & (g2621)));
	assign g8066 = (((!g3499) & (g4848) & (!g2623)) + ((!g3499) & (g4848) & (g2623)) + ((g3499) & (!g4848) & (g2623)) + ((g3499) & (g4848) & (g2623)));
	assign g2624 = (((!g1241) & (g2559) & (!g2560)) + ((g1241) & (!g2559) & (!g2560)) + ((g1241) & (g2559) & (!g2560)) + ((g1241) & (g2559) & (g2560)));
	assign g2625 = (((!g827) & (!g1287) & (g2623) & (!g2624)) + ((!g827) & (!g1287) & (g2623) & (g2624)) + ((!g827) & (g1287) & (g2623) & (!g2624)) + ((!g827) & (g1287) & (g2623) & (g2624)) + ((g827) & (!g1287) & (!g2623) & (g2624)) + ((g827) & (!g1287) & (g2623) & (!g2624)) + ((g827) & (g1287) & (!g2623) & (!g2624)) + ((g827) & (g1287) & (g2623) & (g2624)));
	assign g8067 = (((!g3464) & (g4851) & (!g2626)) + ((!g3464) & (g4851) & (g2626)) + ((g3464) & (!g4851) & (g2626)) + ((g3464) & (g4851) & (g2626)));
	assign g2627 = (((!g1249) & (g2569) & (!g2570)) + ((g1249) & (!g2569) & (!g2570)) + ((g1249) & (g2569) & (!g2570)) + ((g1249) & (g2569) & (g2570)));
	assign g2628 = (((!g827) & (!g1289) & (g2626) & (!g2627)) + ((!g827) & (!g1289) & (g2626) & (g2627)) + ((!g827) & (g1289) & (g2626) & (!g2627)) + ((!g827) & (g1289) & (g2626) & (g2627)) + ((g827) & (!g1289) & (!g2626) & (g2627)) + ((g827) & (!g1289) & (g2626) & (!g2627)) + ((g827) & (g1289) & (!g2626) & (!g2627)) + ((g827) & (g1289) & (g2626) & (g2627)));
	assign g8068 = (((!g2017) & (g6352) & (!g2629)) + ((!g2017) & (g6352) & (g2629)) + ((g2017) & (!g6352) & (g2629)) + ((g2017) & (g6352) & (g2629)));
	assign g2630 = (((!g1257) & (g2581) & (!g2582)) + ((g1257) & (!g2581) & (!g2582)) + ((g1257) & (g2581) & (!g2582)) + ((g1257) & (g2581) & (g2582)));
	assign g2631 = (((!g827) & (!g1291) & (g2629) & (!g2630)) + ((!g827) & (!g1291) & (g2629) & (g2630)) + ((!g827) & (g1291) & (g2629) & (!g2630)) + ((!g827) & (g1291) & (g2629) & (g2630)) + ((g827) & (!g1291) & (!g2629) & (g2630)) + ((g827) & (!g1291) & (g2629) & (!g2630)) + ((g827) & (g1291) & (!g2629) & (!g2630)) + ((g827) & (g1291) & (g2629) & (g2630)));
	assign g8069 = (((!g3429) & (g4856) & (!g2632)) + ((!g3429) & (g4856) & (g2632)) + ((g3429) & (!g4856) & (g2632)) + ((g3429) & (g4856) & (g2632)));
	assign g2633 = (((!g1265) & (g2592) & (!g2593)) + ((g1265) & (!g2592) & (!g2593)) + ((g1265) & (g2592) & (!g2593)) + ((g1265) & (g2592) & (g2593)));
	assign g2634 = (((!g827) & (!g1293) & (g2632) & (!g2633)) + ((!g827) & (!g1293) & (g2632) & (g2633)) + ((!g827) & (g1293) & (g2632) & (!g2633)) + ((!g827) & (g1293) & (g2632) & (g2633)) + ((g827) & (!g1293) & (!g2632) & (g2633)) + ((g827) & (!g1293) & (g2632) & (!g2633)) + ((g827) & (g1293) & (!g2632) & (!g2633)) + ((g827) & (g1293) & (g2632) & (g2633)));
	assign g2635 = (((!g1243) & (g1973) & (!g2562)) + ((g1243) & (!g1973) & (!g2562)) + ((g1243) & (g1973) & (!g2562)) + ((g1243) & (g1973) & (g2562)));
	assign g2636 = (((!g827) & (!g1295) & (g1976) & (!g2635)) + ((!g827) & (!g1295) & (g1976) & (g2635)) + ((!g827) & (g1295) & (g1976) & (!g2635)) + ((!g827) & (g1295) & (g1976) & (g2635)) + ((g827) & (!g1295) & (!g1976) & (g2635)) + ((g827) & (!g1295) & (g1976) & (!g2635)) + ((g827) & (g1295) & (!g1976) & (!g2635)) + ((g827) & (g1295) & (g1976) & (g2635)));
	assign g8070 = (((!g3499) & (g4858) & (!g2637)) + ((!g3499) & (g4858) & (g2637)) + ((g3499) & (!g4858) & (g2637)) + ((g3499) & (g4858) & (g2637)));
	assign g2638 = (((!g1251) & (g2572) & (!g2573)) + ((g1251) & (!g2572) & (!g2573)) + ((g1251) & (g2572) & (!g2573)) + ((g1251) & (g2572) & (g2573)));
	assign g2639 = (((!g827) & (!g1297) & (g2637) & (!g2638)) + ((!g827) & (!g1297) & (g2637) & (g2638)) + ((!g827) & (g1297) & (g2637) & (!g2638)) + ((!g827) & (g1297) & (g2637) & (g2638)) + ((g827) & (!g1297) & (!g2637) & (g2638)) + ((g827) & (!g1297) & (g2637) & (!g2638)) + ((g827) & (g1297) & (!g2637) & (!g2638)) + ((g827) & (g1297) & (g2637) & (g2638)));
	assign g8071 = (((!g3429) & (g4861) & (!g2640)) + ((!g3429) & (g4861) & (g2640)) + ((g3429) & (!g4861) & (g2640)) + ((g3429) & (g4861) & (g2640)));
	assign g2641 = (((!g1259) & (g2584) & (!g2585)) + ((g1259) & (!g2584) & (!g2585)) + ((g1259) & (g2584) & (!g2585)) + ((g1259) & (g2584) & (g2585)));
	assign g2642 = (((!g827) & (!g1299) & (g2640) & (!g2641)) + ((!g827) & (!g1299) & (g2640) & (g2641)) + ((!g827) & (g1299) & (g2640) & (!g2641)) + ((!g827) & (g1299) & (g2640) & (g2641)) + ((g827) & (!g1299) & (!g2640) & (g2641)) + ((g827) & (!g1299) & (g2640) & (!g2641)) + ((g827) & (g1299) & (!g2640) & (!g2641)) + ((g827) & (g1299) & (g2640) & (g2641)));
	assign g8072 = (((!g2017) & (g6334) & (!g2643)) + ((!g2017) & (g6334) & (g2643)) + ((g2017) & (!g6334) & (g2643)) + ((g2017) & (g6334) & (g2643)));
	assign g2644 = (((!g1267) & (g2595) & (!g2596)) + ((g1267) & (!g2595) & (!g2596)) + ((g1267) & (g2595) & (!g2596)) + ((g1267) & (g2595) & (g2596)));
	assign g2645 = (((!g827) & (!g1301) & (g2643) & (!g2644)) + ((!g827) & (!g1301) & (g2643) & (g2644)) + ((!g827) & (g1301) & (g2643) & (!g2644)) + ((!g827) & (g1301) & (g2643) & (g2644)) + ((g827) & (!g1301) & (!g2643) & (g2644)) + ((g827) & (!g1301) & (g2643) & (!g2644)) + ((g827) & (g1301) & (!g2643) & (!g2644)) + ((g827) & (g1301) & (g2643) & (g2644)));
	assign g2646 = (((!g2549) & (!g2550) & (!g2551) & (!g2552) & (g2598) & (g2599)) + ((!g2549) & (!g2550) & (!g2551) & (g2552) & (g2598) & (g2599)) + ((!g2549) & (!g2550) & (g2551) & (!g2552) & (g2598) & (g2599)) + ((!g2549) & (!g2550) & (g2551) & (g2552) & (!g2598) & (g2599)) + ((!g2549) & (!g2550) & (g2551) & (g2552) & (g2598) & (!g2599)) + ((!g2549) & (!g2550) & (g2551) & (g2552) & (g2598) & (g2599)) + ((!g2549) & (g2550) & (!g2551) & (!g2552) & (g2598) & (g2599)) + ((!g2549) & (g2550) & (!g2551) & (g2552) & (!g2598) & (g2599)) + ((!g2549) & (g2550) & (!g2551) & (g2552) & (g2598) & (!g2599)) + ((!g2549) & (g2550) & (!g2551) & (g2552) & (g2598) & (g2599)) + ((!g2549) & (g2550) & (g2551) & (!g2552) & (!g2598) & (g2599)) + ((!g2549) & (g2550) & (g2551) & (!g2552) & (g2598) & (!g2599)) + ((!g2549) & (g2550) & (g2551) & (!g2552) & (g2598) & (g2599)) + ((!g2549) & (g2550) & (g2551) & (g2552) & (!g2598) & (g2599)) + ((!g2549) & (g2550) & (g2551) & (g2552) & (g2598) & (!g2599)) + ((!g2549) & (g2550) & (g2551) & (g2552) & (g2598) & (g2599)) + ((g2549) & (!g2550) & (!g2551) & (!g2552) & (g2598) & (g2599)) + ((g2549) & (!g2550) & (!g2551) & (g2552) & (!g2598) & (g2599)) + ((g2549) & (!g2550) & (!g2551) & (g2552) & (g2598) & (!g2599)) + ((g2549) & (!g2550) & (!g2551) & (g2552) & (g2598) & (g2599)) + ((g2549) & (!g2550) & (g2551) & (!g2552) & (!g2598) & (g2599)) + ((g2549) & (!g2550) & (g2551) & (!g2552) & (g2598) & (!g2599)) + ((g2549) & (!g2550) & (g2551) & (!g2552) & (g2598) & (g2599)) + ((g2549) & (!g2550) & (g2551) & (g2552) & (!g2598) & (g2599)) + ((g2549) & (!g2550) & (g2551) & (g2552) & (g2598) & (!g2599)) + ((g2549) & (!g2550) & (g2551) & (g2552) & (g2598) & (g2599)) + ((g2549) & (g2550) & (!g2551) & (!g2552) & (g2598) & (g2599)) + ((g2549) & (g2550) & (!g2551) & (g2552) & (!g2598) & (g2599)) + ((g2549) & (g2550) & (!g2551) & (g2552) & (g2598) & (!g2599)) + ((g2549) & (g2550) & (!g2551) & (g2552) & (g2598) & (g2599)) + ((g2549) & (g2550) & (g2551) & (!g2552) & (!g2598) & (g2599)) + ((g2549) & (g2550) & (g2551) & (!g2552) & (g2598) & (!g2599)) + ((g2549) & (g2550) & (g2551) & (!g2552) & (g2598) & (g2599)) + ((g2549) & (g2550) & (g2551) & (g2552) & (!g2598) & (g2599)) + ((g2549) & (g2550) & (g2551) & (g2552) & (g2598) & (!g2599)) + ((g2549) & (g2550) & (g2551) & (g2552) & (g2598) & (g2599)));
	assign g8073 = (((!g3429) & (g4868) & (!g2647)) + ((!g3429) & (g4868) & (g2647)) + ((g3429) & (!g4868) & (g2647)) + ((g3429) & (g4868) & (g2647)));
	assign g8074 = (((!g3464) & (g4872) & (!g2648)) + ((!g3464) & (g4872) & (g2648)) + ((g3464) & (!g4872) & (g2648)) + ((g3464) & (g4872) & (g2648)));
	assign g8075 = (((!g3429) & (g4878) & (!g2649)) + ((!g3429) & (g4878) & (g2649)) + ((g3429) & (!g4878) & (g2649)) + ((g3429) & (g4878) & (g2649)));
	assign g8076 = (((!g3499) & (g4882) & (!g2650)) + ((!g3499) & (g4882) & (g2650)) + ((g3499) & (!g4882) & (g2650)) + ((g3499) & (g4882) & (g2650)));
	assign g2651 = (((!g2554) & (!g2555) & (!g2556) & (!g2601) & (!g2602) & (!g5684)) + ((!g2554) & (!g2555) & (!g2556) & (!g2601) & (g2602) & (!g5684)) + ((!g2554) & (!g2555) & (!g2556) & (g2601) & (!g2602) & (!g5684)) + ((!g2554) & (!g2555) & (!g2556) & (g2601) & (g2602) & (g5684)) + ((!g2554) & (!g2555) & (g2556) & (!g2601) & (!g2602) & (!g5684)) + ((!g2554) & (!g2555) & (g2556) & (!g2601) & (g2602) & (!g5684)) + ((!g2554) & (!g2555) & (g2556) & (g2601) & (!g2602) & (!g5684)) + ((!g2554) & (!g2555) & (g2556) & (g2601) & (g2602) & (g5684)) + ((!g2554) & (g2555) & (!g2556) & (!g2601) & (!g2602) & (!g5684)) + ((!g2554) & (g2555) & (!g2556) & (!g2601) & (g2602) & (!g5684)) + ((!g2554) & (g2555) & (!g2556) & (g2601) & (!g2602) & (!g5684)) + ((!g2554) & (g2555) & (!g2556) & (g2601) & (g2602) & (g5684)) + ((!g2554) & (g2555) & (g2556) & (!g2601) & (!g2602) & (!g5684)) + ((!g2554) & (g2555) & (g2556) & (!g2601) & (g2602) & (g5684)) + ((!g2554) & (g2555) & (g2556) & (g2601) & (!g2602) & (g5684)) + ((!g2554) & (g2555) & (g2556) & (g2601) & (g2602) & (g5684)) + ((g2554) & (!g2555) & (!g2556) & (!g2601) & (!g2602) & (!g5684)) + ((g2554) & (!g2555) & (!g2556) & (!g2601) & (g2602) & (!g5684)) + ((g2554) & (!g2555) & (!g2556) & (g2601) & (!g2602) & (!g5684)) + ((g2554) & (!g2555) & (!g2556) & (g2601) & (g2602) & (g5684)) + ((g2554) & (!g2555) & (g2556) & (!g2601) & (!g2602) & (!g5684)) + ((g2554) & (!g2555) & (g2556) & (!g2601) & (g2602) & (g5684)) + ((g2554) & (!g2555) & (g2556) & (g2601) & (!g2602) & (g5684)) + ((g2554) & (!g2555) & (g2556) & (g2601) & (g2602) & (g5684)) + ((g2554) & (g2555) & (!g2556) & (!g2601) & (!g2602) & (!g5684)) + ((g2554) & (g2555) & (!g2556) & (!g2601) & (g2602) & (g5684)) + ((g2554) & (g2555) & (!g2556) & (g2601) & (!g2602) & (g5684)) + ((g2554) & (g2555) & (!g2556) & (g2601) & (g2602) & (g5684)) + ((g2554) & (g2555) & (g2556) & (!g2601) & (!g2602) & (!g5684)) + ((g2554) & (g2555) & (g2556) & (!g2601) & (g2602) & (g5684)) + ((g2554) & (g2555) & (g2556) & (g2601) & (!g2602) & (g5684)) + ((g2554) & (g2555) & (g2556) & (g2601) & (g2602) & (g5684)));
	assign g2652 = (((!g827) & (!g1279) & (!g1307) & (!g1975) & (g2047) & (!g2612)) + ((!g827) & (!g1279) & (!g1307) & (!g1975) & (g2047) & (g2612)) + ((!g827) & (!g1279) & (!g1307) & (g1975) & (g2047) & (!g2612)) + ((!g827) & (!g1279) & (!g1307) & (g1975) & (g2047) & (g2612)) + ((!g827) & (!g1279) & (g1307) & (!g1975) & (g2047) & (!g2612)) + ((!g827) & (!g1279) & (g1307) & (!g1975) & (g2047) & (g2612)) + ((!g827) & (!g1279) & (g1307) & (g1975) & (g2047) & (!g2612)) + ((!g827) & (!g1279) & (g1307) & (g1975) & (g2047) & (g2612)) + ((!g827) & (g1279) & (!g1307) & (!g1975) & (g2047) & (!g2612)) + ((!g827) & (g1279) & (!g1307) & (!g1975) & (g2047) & (g2612)) + ((!g827) & (g1279) & (!g1307) & (g1975) & (g2047) & (!g2612)) + ((!g827) & (g1279) & (!g1307) & (g1975) & (g2047) & (g2612)) + ((!g827) & (g1279) & (g1307) & (!g1975) & (g2047) & (!g2612)) + ((!g827) & (g1279) & (g1307) & (!g1975) & (g2047) & (g2612)) + ((!g827) & (g1279) & (g1307) & (g1975) & (g2047) & (!g2612)) + ((!g827) & (g1279) & (g1307) & (g1975) & (g2047) & (g2612)) + ((g827) & (!g1279) & (!g1307) & (!g1975) & (g2047) & (!g2612)) + ((g827) & (!g1279) & (!g1307) & (!g1975) & (g2047) & (g2612)) + ((g827) & (!g1279) & (!g1307) & (g1975) & (!g2047) & (g2612)) + ((g827) & (!g1279) & (!g1307) & (g1975) & (g2047) & (!g2612)) + ((g827) & (!g1279) & (g1307) & (!g1975) & (!g2047) & (!g2612)) + ((g827) & (!g1279) & (g1307) & (!g1975) & (!g2047) & (g2612)) + ((g827) & (!g1279) & (g1307) & (g1975) & (!g2047) & (!g2612)) + ((g827) & (!g1279) & (g1307) & (g1975) & (g2047) & (g2612)) + ((g827) & (g1279) & (!g1307) & (!g1975) & (!g2047) & (g2612)) + ((g827) & (g1279) & (!g1307) & (!g1975) & (g2047) & (!g2612)) + ((g827) & (g1279) & (!g1307) & (g1975) & (!g2047) & (!g2612)) + ((g827) & (g1279) & (!g1307) & (g1975) & (!g2047) & (g2612)) + ((g827) & (g1279) & (g1307) & (!g1975) & (!g2047) & (!g2612)) + ((g827) & (g1279) & (g1307) & (!g1975) & (g2047) & (g2612)) + ((g827) & (g1279) & (g1307) & (g1975) & (g2047) & (!g2612)) + ((g827) & (g1279) & (g1307) & (g1975) & (g2047) & (g2612)));
	assign g8077 = (((!g3499) & (g4885) & (!g2653)) + ((!g3499) & (g4885) & (g2653)) + ((g3499) & (!g4885) & (g2653)) + ((g3499) & (g4885) & (g2653)));
	assign g2654 = (((!g827) & (!g1287) & (!g1309) & (!g2623) & (g2653) & (!g2624)) + ((!g827) & (!g1287) & (!g1309) & (!g2623) & (g2653) & (g2624)) + ((!g827) & (!g1287) & (!g1309) & (g2623) & (g2653) & (!g2624)) + ((!g827) & (!g1287) & (!g1309) & (g2623) & (g2653) & (g2624)) + ((!g827) & (!g1287) & (g1309) & (!g2623) & (g2653) & (!g2624)) + ((!g827) & (!g1287) & (g1309) & (!g2623) & (g2653) & (g2624)) + ((!g827) & (!g1287) & (g1309) & (g2623) & (g2653) & (!g2624)) + ((!g827) & (!g1287) & (g1309) & (g2623) & (g2653) & (g2624)) + ((!g827) & (g1287) & (!g1309) & (!g2623) & (g2653) & (!g2624)) + ((!g827) & (g1287) & (!g1309) & (!g2623) & (g2653) & (g2624)) + ((!g827) & (g1287) & (!g1309) & (g2623) & (g2653) & (!g2624)) + ((!g827) & (g1287) & (!g1309) & (g2623) & (g2653) & (g2624)) + ((!g827) & (g1287) & (g1309) & (!g2623) & (g2653) & (!g2624)) + ((!g827) & (g1287) & (g1309) & (!g2623) & (g2653) & (g2624)) + ((!g827) & (g1287) & (g1309) & (g2623) & (g2653) & (!g2624)) + ((!g827) & (g1287) & (g1309) & (g2623) & (g2653) & (g2624)) + ((g827) & (!g1287) & (!g1309) & (!g2623) & (g2653) & (!g2624)) + ((g827) & (!g1287) & (!g1309) & (!g2623) & (g2653) & (g2624)) + ((g827) & (!g1287) & (!g1309) & (g2623) & (!g2653) & (g2624)) + ((g827) & (!g1287) & (!g1309) & (g2623) & (g2653) & (!g2624)) + ((g827) & (!g1287) & (g1309) & (!g2623) & (!g2653) & (!g2624)) + ((g827) & (!g1287) & (g1309) & (!g2623) & (!g2653) & (g2624)) + ((g827) & (!g1287) & (g1309) & (g2623) & (!g2653) & (!g2624)) + ((g827) & (!g1287) & (g1309) & (g2623) & (g2653) & (g2624)) + ((g827) & (g1287) & (!g1309) & (!g2623) & (!g2653) & (g2624)) + ((g827) & (g1287) & (!g1309) & (!g2623) & (g2653) & (!g2624)) + ((g827) & (g1287) & (!g1309) & (g2623) & (!g2653) & (!g2624)) + ((g827) & (g1287) & (!g1309) & (g2623) & (!g2653) & (g2624)) + ((g827) & (g1287) & (g1309) & (!g2623) & (!g2653) & (!g2624)) + ((g827) & (g1287) & (g1309) & (!g2623) & (g2653) & (g2624)) + ((g827) & (g1287) & (g1309) & (g2623) & (g2653) & (!g2624)) + ((g827) & (g1287) & (g1309) & (g2623) & (g2653) & (g2624)));
	assign g2655 = (((!g827) & (!g1295) & (!g1311) & (!g1976) & (g2048) & (!g2635)) + ((!g827) & (!g1295) & (!g1311) & (!g1976) & (g2048) & (g2635)) + ((!g827) & (!g1295) & (!g1311) & (g1976) & (g2048) & (!g2635)) + ((!g827) & (!g1295) & (!g1311) & (g1976) & (g2048) & (g2635)) + ((!g827) & (!g1295) & (g1311) & (!g1976) & (g2048) & (!g2635)) + ((!g827) & (!g1295) & (g1311) & (!g1976) & (g2048) & (g2635)) + ((!g827) & (!g1295) & (g1311) & (g1976) & (g2048) & (!g2635)) + ((!g827) & (!g1295) & (g1311) & (g1976) & (g2048) & (g2635)) + ((!g827) & (g1295) & (!g1311) & (!g1976) & (g2048) & (!g2635)) + ((!g827) & (g1295) & (!g1311) & (!g1976) & (g2048) & (g2635)) + ((!g827) & (g1295) & (!g1311) & (g1976) & (g2048) & (!g2635)) + ((!g827) & (g1295) & (!g1311) & (g1976) & (g2048) & (g2635)) + ((!g827) & (g1295) & (g1311) & (!g1976) & (g2048) & (!g2635)) + ((!g827) & (g1295) & (g1311) & (!g1976) & (g2048) & (g2635)) + ((!g827) & (g1295) & (g1311) & (g1976) & (g2048) & (!g2635)) + ((!g827) & (g1295) & (g1311) & (g1976) & (g2048) & (g2635)) + ((g827) & (!g1295) & (!g1311) & (!g1976) & (g2048) & (!g2635)) + ((g827) & (!g1295) & (!g1311) & (!g1976) & (g2048) & (g2635)) + ((g827) & (!g1295) & (!g1311) & (g1976) & (!g2048) & (g2635)) + ((g827) & (!g1295) & (!g1311) & (g1976) & (g2048) & (!g2635)) + ((g827) & (!g1295) & (g1311) & (!g1976) & (!g2048) & (!g2635)) + ((g827) & (!g1295) & (g1311) & (!g1976) & (!g2048) & (g2635)) + ((g827) & (!g1295) & (g1311) & (g1976) & (!g2048) & (!g2635)) + ((g827) & (!g1295) & (g1311) & (g1976) & (g2048) & (g2635)) + ((g827) & (g1295) & (!g1311) & (!g1976) & (!g2048) & (g2635)) + ((g827) & (g1295) & (!g1311) & (!g1976) & (g2048) & (!g2635)) + ((g827) & (g1295) & (!g1311) & (g1976) & (!g2048) & (!g2635)) + ((g827) & (g1295) & (!g1311) & (g1976) & (!g2048) & (g2635)) + ((g827) & (g1295) & (g1311) & (!g1976) & (!g2048) & (!g2635)) + ((g827) & (g1295) & (g1311) & (!g1976) & (g2048) & (g2635)) + ((g827) & (g1295) & (g1311) & (g1976) & (g2048) & (!g2635)) + ((g827) & (g1295) & (g1311) & (g1976) & (g2048) & (g2635)));
	assign g2656 = (((!g827) & (!g1273) & (!g1313) & (!g2013) & (g2051) & (!g2605)) + ((!g827) & (!g1273) & (!g1313) & (!g2013) & (g2051) & (g2605)) + ((!g827) & (!g1273) & (!g1313) & (g2013) & (g2051) & (!g2605)) + ((!g827) & (!g1273) & (!g1313) & (g2013) & (g2051) & (g2605)) + ((!g827) & (!g1273) & (g1313) & (!g2013) & (g2051) & (!g2605)) + ((!g827) & (!g1273) & (g1313) & (!g2013) & (g2051) & (g2605)) + ((!g827) & (!g1273) & (g1313) & (g2013) & (g2051) & (!g2605)) + ((!g827) & (!g1273) & (g1313) & (g2013) & (g2051) & (g2605)) + ((!g827) & (g1273) & (!g1313) & (!g2013) & (g2051) & (!g2605)) + ((!g827) & (g1273) & (!g1313) & (!g2013) & (g2051) & (g2605)) + ((!g827) & (g1273) & (!g1313) & (g2013) & (g2051) & (!g2605)) + ((!g827) & (g1273) & (!g1313) & (g2013) & (g2051) & (g2605)) + ((!g827) & (g1273) & (g1313) & (!g2013) & (g2051) & (!g2605)) + ((!g827) & (g1273) & (g1313) & (!g2013) & (g2051) & (g2605)) + ((!g827) & (g1273) & (g1313) & (g2013) & (g2051) & (!g2605)) + ((!g827) & (g1273) & (g1313) & (g2013) & (g2051) & (g2605)) + ((g827) & (!g1273) & (!g1313) & (!g2013) & (g2051) & (!g2605)) + ((g827) & (!g1273) & (!g1313) & (!g2013) & (g2051) & (g2605)) + ((g827) & (!g1273) & (!g1313) & (g2013) & (!g2051) & (g2605)) + ((g827) & (!g1273) & (!g1313) & (g2013) & (g2051) & (!g2605)) + ((g827) & (!g1273) & (g1313) & (!g2013) & (!g2051) & (!g2605)) + ((g827) & (!g1273) & (g1313) & (!g2013) & (!g2051) & (g2605)) + ((g827) & (!g1273) & (g1313) & (g2013) & (!g2051) & (!g2605)) + ((g827) & (!g1273) & (g1313) & (g2013) & (g2051) & (g2605)) + ((g827) & (g1273) & (!g1313) & (!g2013) & (!g2051) & (g2605)) + ((g827) & (g1273) & (!g1313) & (!g2013) & (g2051) & (!g2605)) + ((g827) & (g1273) & (!g1313) & (g2013) & (!g2051) & (!g2605)) + ((g827) & (g1273) & (!g1313) & (g2013) & (!g2051) & (g2605)) + ((g827) & (g1273) & (g1313) & (!g2013) & (!g2051) & (!g2605)) + ((g827) & (g1273) & (g1313) & (!g2013) & (g2051) & (g2605)) + ((g827) & (g1273) & (g1313) & (g2013) & (g2051) & (!g2605)) + ((g827) & (g1273) & (g1313) & (g2013) & (g2051) & (g2605)));
	assign g8078 = (((!g2017) & (g4889) & (!g2657)) + ((!g2017) & (g4889) & (g2657)) + ((g2017) & (!g4889) & (g2657)) + ((g2017) & (g4889) & (g2657)));
	assign g2658 = (((!g827) & (!g1281) & (!g1315) & (!g2614) & (g2657) & (!g2615)) + ((!g827) & (!g1281) & (!g1315) & (!g2614) & (g2657) & (g2615)) + ((!g827) & (!g1281) & (!g1315) & (g2614) & (g2657) & (!g2615)) + ((!g827) & (!g1281) & (!g1315) & (g2614) & (g2657) & (g2615)) + ((!g827) & (!g1281) & (g1315) & (!g2614) & (g2657) & (!g2615)) + ((!g827) & (!g1281) & (g1315) & (!g2614) & (g2657) & (g2615)) + ((!g827) & (!g1281) & (g1315) & (g2614) & (g2657) & (!g2615)) + ((!g827) & (!g1281) & (g1315) & (g2614) & (g2657) & (g2615)) + ((!g827) & (g1281) & (!g1315) & (!g2614) & (g2657) & (!g2615)) + ((!g827) & (g1281) & (!g1315) & (!g2614) & (g2657) & (g2615)) + ((!g827) & (g1281) & (!g1315) & (g2614) & (g2657) & (!g2615)) + ((!g827) & (g1281) & (!g1315) & (g2614) & (g2657) & (g2615)) + ((!g827) & (g1281) & (g1315) & (!g2614) & (g2657) & (!g2615)) + ((!g827) & (g1281) & (g1315) & (!g2614) & (g2657) & (g2615)) + ((!g827) & (g1281) & (g1315) & (g2614) & (g2657) & (!g2615)) + ((!g827) & (g1281) & (g1315) & (g2614) & (g2657) & (g2615)) + ((g827) & (!g1281) & (!g1315) & (!g2614) & (g2657) & (!g2615)) + ((g827) & (!g1281) & (!g1315) & (!g2614) & (g2657) & (g2615)) + ((g827) & (!g1281) & (!g1315) & (g2614) & (!g2657) & (g2615)) + ((g827) & (!g1281) & (!g1315) & (g2614) & (g2657) & (!g2615)) + ((g827) & (!g1281) & (g1315) & (!g2614) & (!g2657) & (!g2615)) + ((g827) & (!g1281) & (g1315) & (!g2614) & (!g2657) & (g2615)) + ((g827) & (!g1281) & (g1315) & (g2614) & (!g2657) & (!g2615)) + ((g827) & (!g1281) & (g1315) & (g2614) & (g2657) & (g2615)) + ((g827) & (g1281) & (!g1315) & (!g2614) & (!g2657) & (g2615)) + ((g827) & (g1281) & (!g1315) & (!g2614) & (g2657) & (!g2615)) + ((g827) & (g1281) & (!g1315) & (g2614) & (!g2657) & (!g2615)) + ((g827) & (g1281) & (!g1315) & (g2614) & (!g2657) & (g2615)) + ((g827) & (g1281) & (g1315) & (!g2614) & (!g2657) & (!g2615)) + ((g827) & (g1281) & (g1315) & (!g2614) & (g2657) & (g2615)) + ((g827) & (g1281) & (g1315) & (g2614) & (g2657) & (!g2615)) + ((g827) & (g1281) & (g1315) & (g2614) & (g2657) & (g2615)));
	assign g8079 = (((!g3464) & (g4893) & (!g2659)) + ((!g3464) & (g4893) & (g2659)) + ((g3464) & (!g4893) & (g2659)) + ((g3464) & (g4893) & (g2659)));
	assign g2660 = (((!g827) & (!g1289) & (!g1317) & (!g2626) & (g2659) & (!g2627)) + ((!g827) & (!g1289) & (!g1317) & (!g2626) & (g2659) & (g2627)) + ((!g827) & (!g1289) & (!g1317) & (g2626) & (g2659) & (!g2627)) + ((!g827) & (!g1289) & (!g1317) & (g2626) & (g2659) & (g2627)) + ((!g827) & (!g1289) & (g1317) & (!g2626) & (g2659) & (!g2627)) + ((!g827) & (!g1289) & (g1317) & (!g2626) & (g2659) & (g2627)) + ((!g827) & (!g1289) & (g1317) & (g2626) & (g2659) & (!g2627)) + ((!g827) & (!g1289) & (g1317) & (g2626) & (g2659) & (g2627)) + ((!g827) & (g1289) & (!g1317) & (!g2626) & (g2659) & (!g2627)) + ((!g827) & (g1289) & (!g1317) & (!g2626) & (g2659) & (g2627)) + ((!g827) & (g1289) & (!g1317) & (g2626) & (g2659) & (!g2627)) + ((!g827) & (g1289) & (!g1317) & (g2626) & (g2659) & (g2627)) + ((!g827) & (g1289) & (g1317) & (!g2626) & (g2659) & (!g2627)) + ((!g827) & (g1289) & (g1317) & (!g2626) & (g2659) & (g2627)) + ((!g827) & (g1289) & (g1317) & (g2626) & (g2659) & (!g2627)) + ((!g827) & (g1289) & (g1317) & (g2626) & (g2659) & (g2627)) + ((g827) & (!g1289) & (!g1317) & (!g2626) & (g2659) & (!g2627)) + ((g827) & (!g1289) & (!g1317) & (!g2626) & (g2659) & (g2627)) + ((g827) & (!g1289) & (!g1317) & (g2626) & (!g2659) & (g2627)) + ((g827) & (!g1289) & (!g1317) & (g2626) & (g2659) & (!g2627)) + ((g827) & (!g1289) & (g1317) & (!g2626) & (!g2659) & (!g2627)) + ((g827) & (!g1289) & (g1317) & (!g2626) & (!g2659) & (g2627)) + ((g827) & (!g1289) & (g1317) & (g2626) & (!g2659) & (!g2627)) + ((g827) & (!g1289) & (g1317) & (g2626) & (g2659) & (g2627)) + ((g827) & (g1289) & (!g1317) & (!g2626) & (!g2659) & (g2627)) + ((g827) & (g1289) & (!g1317) & (!g2626) & (g2659) & (!g2627)) + ((g827) & (g1289) & (!g1317) & (g2626) & (!g2659) & (!g2627)) + ((g827) & (g1289) & (!g1317) & (g2626) & (!g2659) & (g2627)) + ((g827) & (g1289) & (g1317) & (!g2626) & (!g2659) & (!g2627)) + ((g827) & (g1289) & (g1317) & (!g2626) & (g2659) & (g2627)) + ((g827) & (g1289) & (g1317) & (g2626) & (g2659) & (!g2627)) + ((g827) & (g1289) & (g1317) & (g2626) & (g2659) & (g2627)));
	assign g8080 = (((!g3499) & (g4896) & (!g2661)) + ((!g3499) & (g4896) & (g2661)) + ((g3499) & (!g4896) & (g2661)) + ((g3499) & (g4896) & (g2661)));
	assign g2662 = (((!g827) & (!g1297) & (!g1319) & (!g2637) & (g2661) & (!g2638)) + ((!g827) & (!g1297) & (!g1319) & (!g2637) & (g2661) & (g2638)) + ((!g827) & (!g1297) & (!g1319) & (g2637) & (g2661) & (!g2638)) + ((!g827) & (!g1297) & (!g1319) & (g2637) & (g2661) & (g2638)) + ((!g827) & (!g1297) & (g1319) & (!g2637) & (g2661) & (!g2638)) + ((!g827) & (!g1297) & (g1319) & (!g2637) & (g2661) & (g2638)) + ((!g827) & (!g1297) & (g1319) & (g2637) & (g2661) & (!g2638)) + ((!g827) & (!g1297) & (g1319) & (g2637) & (g2661) & (g2638)) + ((!g827) & (g1297) & (!g1319) & (!g2637) & (g2661) & (!g2638)) + ((!g827) & (g1297) & (!g1319) & (!g2637) & (g2661) & (g2638)) + ((!g827) & (g1297) & (!g1319) & (g2637) & (g2661) & (!g2638)) + ((!g827) & (g1297) & (!g1319) & (g2637) & (g2661) & (g2638)) + ((!g827) & (g1297) & (g1319) & (!g2637) & (g2661) & (!g2638)) + ((!g827) & (g1297) & (g1319) & (!g2637) & (g2661) & (g2638)) + ((!g827) & (g1297) & (g1319) & (g2637) & (g2661) & (!g2638)) + ((!g827) & (g1297) & (g1319) & (g2637) & (g2661) & (g2638)) + ((g827) & (!g1297) & (!g1319) & (!g2637) & (g2661) & (!g2638)) + ((g827) & (!g1297) & (!g1319) & (!g2637) & (g2661) & (g2638)) + ((g827) & (!g1297) & (!g1319) & (g2637) & (!g2661) & (g2638)) + ((g827) & (!g1297) & (!g1319) & (g2637) & (g2661) & (!g2638)) + ((g827) & (!g1297) & (g1319) & (!g2637) & (!g2661) & (!g2638)) + ((g827) & (!g1297) & (g1319) & (!g2637) & (!g2661) & (g2638)) + ((g827) & (!g1297) & (g1319) & (g2637) & (!g2661) & (!g2638)) + ((g827) & (!g1297) & (g1319) & (g2637) & (g2661) & (g2638)) + ((g827) & (g1297) & (!g1319) & (!g2637) & (!g2661) & (g2638)) + ((g827) & (g1297) & (!g1319) & (!g2637) & (g2661) & (!g2638)) + ((g827) & (g1297) & (!g1319) & (g2637) & (!g2661) & (!g2638)) + ((g827) & (g1297) & (!g1319) & (g2637) & (!g2661) & (g2638)) + ((g827) & (g1297) & (g1319) & (!g2637) & (!g2661) & (!g2638)) + ((g827) & (g1297) & (g1319) & (!g2637) & (g2661) & (g2638)) + ((g827) & (g1297) & (g1319) & (g2637) & (g2661) & (!g2638)) + ((g827) & (g1297) & (g1319) & (g2637) & (g2661) & (g2638)));
	assign g8081 = (((!g3464) & (g4899) & (!g2663)) + ((!g3464) & (g4899) & (g2663)) + ((g3464) & (!g4899) & (g2663)) + ((g3464) & (g4899) & (g2663)));
	assign g2664 = (((!g827) & (!g1275) & (!g1321) & (!g2607) & (g2663) & (!g2608)) + ((!g827) & (!g1275) & (!g1321) & (!g2607) & (g2663) & (g2608)) + ((!g827) & (!g1275) & (!g1321) & (g2607) & (g2663) & (!g2608)) + ((!g827) & (!g1275) & (!g1321) & (g2607) & (g2663) & (g2608)) + ((!g827) & (!g1275) & (g1321) & (!g2607) & (g2663) & (!g2608)) + ((!g827) & (!g1275) & (g1321) & (!g2607) & (g2663) & (g2608)) + ((!g827) & (!g1275) & (g1321) & (g2607) & (g2663) & (!g2608)) + ((!g827) & (!g1275) & (g1321) & (g2607) & (g2663) & (g2608)) + ((!g827) & (g1275) & (!g1321) & (!g2607) & (g2663) & (!g2608)) + ((!g827) & (g1275) & (!g1321) & (!g2607) & (g2663) & (g2608)) + ((!g827) & (g1275) & (!g1321) & (g2607) & (g2663) & (!g2608)) + ((!g827) & (g1275) & (!g1321) & (g2607) & (g2663) & (g2608)) + ((!g827) & (g1275) & (g1321) & (!g2607) & (g2663) & (!g2608)) + ((!g827) & (g1275) & (g1321) & (!g2607) & (g2663) & (g2608)) + ((!g827) & (g1275) & (g1321) & (g2607) & (g2663) & (!g2608)) + ((!g827) & (g1275) & (g1321) & (g2607) & (g2663) & (g2608)) + ((g827) & (!g1275) & (!g1321) & (!g2607) & (g2663) & (!g2608)) + ((g827) & (!g1275) & (!g1321) & (!g2607) & (g2663) & (g2608)) + ((g827) & (!g1275) & (!g1321) & (g2607) & (!g2663) & (g2608)) + ((g827) & (!g1275) & (!g1321) & (g2607) & (g2663) & (!g2608)) + ((g827) & (!g1275) & (g1321) & (!g2607) & (!g2663) & (!g2608)) + ((g827) & (!g1275) & (g1321) & (!g2607) & (!g2663) & (g2608)) + ((g827) & (!g1275) & (g1321) & (g2607) & (!g2663) & (!g2608)) + ((g827) & (!g1275) & (g1321) & (g2607) & (g2663) & (g2608)) + ((g827) & (g1275) & (!g1321) & (!g2607) & (!g2663) & (g2608)) + ((g827) & (g1275) & (!g1321) & (!g2607) & (g2663) & (!g2608)) + ((g827) & (g1275) & (!g1321) & (g2607) & (!g2663) & (!g2608)) + ((g827) & (g1275) & (!g1321) & (g2607) & (!g2663) & (g2608)) + ((g827) & (g1275) & (g1321) & (!g2607) & (!g2663) & (!g2608)) + ((g827) & (g1275) & (g1321) & (!g2607) & (g2663) & (g2608)) + ((g827) & (g1275) & (g1321) & (g2607) & (g2663) & (!g2608)) + ((g827) & (g1275) & (g1321) & (g2607) & (g2663) & (g2608)));
	assign g8082 = (((!g3499) & (g4902) & (!g2665)) + ((!g3499) & (g4902) & (g2665)) + ((g3499) & (!g4902) & (g2665)) + ((g3499) & (g4902) & (g2665)));
	assign g2666 = (((!g827) & (!g1283) & (!g1323) & (!g2617) & (g2665) & (!g2618)) + ((!g827) & (!g1283) & (!g1323) & (!g2617) & (g2665) & (g2618)) + ((!g827) & (!g1283) & (!g1323) & (g2617) & (g2665) & (!g2618)) + ((!g827) & (!g1283) & (!g1323) & (g2617) & (g2665) & (g2618)) + ((!g827) & (!g1283) & (g1323) & (!g2617) & (g2665) & (!g2618)) + ((!g827) & (!g1283) & (g1323) & (!g2617) & (g2665) & (g2618)) + ((!g827) & (!g1283) & (g1323) & (g2617) & (g2665) & (!g2618)) + ((!g827) & (!g1283) & (g1323) & (g2617) & (g2665) & (g2618)) + ((!g827) & (g1283) & (!g1323) & (!g2617) & (g2665) & (!g2618)) + ((!g827) & (g1283) & (!g1323) & (!g2617) & (g2665) & (g2618)) + ((!g827) & (g1283) & (!g1323) & (g2617) & (g2665) & (!g2618)) + ((!g827) & (g1283) & (!g1323) & (g2617) & (g2665) & (g2618)) + ((!g827) & (g1283) & (g1323) & (!g2617) & (g2665) & (!g2618)) + ((!g827) & (g1283) & (g1323) & (!g2617) & (g2665) & (g2618)) + ((!g827) & (g1283) & (g1323) & (g2617) & (g2665) & (!g2618)) + ((!g827) & (g1283) & (g1323) & (g2617) & (g2665) & (g2618)) + ((g827) & (!g1283) & (!g1323) & (!g2617) & (g2665) & (!g2618)) + ((g827) & (!g1283) & (!g1323) & (!g2617) & (g2665) & (g2618)) + ((g827) & (!g1283) & (!g1323) & (g2617) & (!g2665) & (g2618)) + ((g827) & (!g1283) & (!g1323) & (g2617) & (g2665) & (!g2618)) + ((g827) & (!g1283) & (g1323) & (!g2617) & (!g2665) & (!g2618)) + ((g827) & (!g1283) & (g1323) & (!g2617) & (!g2665) & (g2618)) + ((g827) & (!g1283) & (g1323) & (g2617) & (!g2665) & (!g2618)) + ((g827) & (!g1283) & (g1323) & (g2617) & (g2665) & (g2618)) + ((g827) & (g1283) & (!g1323) & (!g2617) & (!g2665) & (g2618)) + ((g827) & (g1283) & (!g1323) & (!g2617) & (g2665) & (!g2618)) + ((g827) & (g1283) & (!g1323) & (g2617) & (!g2665) & (!g2618)) + ((g827) & (g1283) & (!g1323) & (g2617) & (!g2665) & (g2618)) + ((g827) & (g1283) & (g1323) & (!g2617) & (!g2665) & (!g2618)) + ((g827) & (g1283) & (g1323) & (!g2617) & (g2665) & (g2618)) + ((g827) & (g1283) & (g1323) & (g2617) & (g2665) & (!g2618)) + ((g827) & (g1283) & (g1323) & (g2617) & (g2665) & (g2618)));
	assign g8083 = (((!g2017) & (g4906) & (!g2667)) + ((!g2017) & (g4906) & (g2667)) + ((g2017) & (!g4906) & (g2667)) + ((g2017) & (g4906) & (g2667)));
	assign g2668 = (((!g827) & (!g1291) & (!g1325) & (!g2629) & (g2667) & (!g2630)) + ((!g827) & (!g1291) & (!g1325) & (!g2629) & (g2667) & (g2630)) + ((!g827) & (!g1291) & (!g1325) & (g2629) & (g2667) & (!g2630)) + ((!g827) & (!g1291) & (!g1325) & (g2629) & (g2667) & (g2630)) + ((!g827) & (!g1291) & (g1325) & (!g2629) & (g2667) & (!g2630)) + ((!g827) & (!g1291) & (g1325) & (!g2629) & (g2667) & (g2630)) + ((!g827) & (!g1291) & (g1325) & (g2629) & (g2667) & (!g2630)) + ((!g827) & (!g1291) & (g1325) & (g2629) & (g2667) & (g2630)) + ((!g827) & (g1291) & (!g1325) & (!g2629) & (g2667) & (!g2630)) + ((!g827) & (g1291) & (!g1325) & (!g2629) & (g2667) & (g2630)) + ((!g827) & (g1291) & (!g1325) & (g2629) & (g2667) & (!g2630)) + ((!g827) & (g1291) & (!g1325) & (g2629) & (g2667) & (g2630)) + ((!g827) & (g1291) & (g1325) & (!g2629) & (g2667) & (!g2630)) + ((!g827) & (g1291) & (g1325) & (!g2629) & (g2667) & (g2630)) + ((!g827) & (g1291) & (g1325) & (g2629) & (g2667) & (!g2630)) + ((!g827) & (g1291) & (g1325) & (g2629) & (g2667) & (g2630)) + ((g827) & (!g1291) & (!g1325) & (!g2629) & (g2667) & (!g2630)) + ((g827) & (!g1291) & (!g1325) & (!g2629) & (g2667) & (g2630)) + ((g827) & (!g1291) & (!g1325) & (g2629) & (!g2667) & (g2630)) + ((g827) & (!g1291) & (!g1325) & (g2629) & (g2667) & (!g2630)) + ((g827) & (!g1291) & (g1325) & (!g2629) & (!g2667) & (!g2630)) + ((g827) & (!g1291) & (g1325) & (!g2629) & (!g2667) & (g2630)) + ((g827) & (!g1291) & (g1325) & (g2629) & (!g2667) & (!g2630)) + ((g827) & (!g1291) & (g1325) & (g2629) & (g2667) & (g2630)) + ((g827) & (g1291) & (!g1325) & (!g2629) & (!g2667) & (g2630)) + ((g827) & (g1291) & (!g1325) & (!g2629) & (g2667) & (!g2630)) + ((g827) & (g1291) & (!g1325) & (g2629) & (!g2667) & (!g2630)) + ((g827) & (g1291) & (!g1325) & (g2629) & (!g2667) & (g2630)) + ((g827) & (g1291) & (g1325) & (!g2629) & (!g2667) & (!g2630)) + ((g827) & (g1291) & (g1325) & (!g2629) & (g2667) & (g2630)) + ((g827) & (g1291) & (g1325) & (g2629) & (g2667) & (!g2630)) + ((g827) & (g1291) & (g1325) & (g2629) & (g2667) & (g2630)));
	assign g8084 = (((!g3429) & (g4911) & (!g2669)) + ((!g3429) & (g4911) & (g2669)) + ((g3429) & (!g4911) & (g2669)) + ((g3429) & (g4911) & (g2669)));
	assign g2670 = (((!g827) & (!g1299) & (!g1327) & (!g2640) & (g2669) & (!g2641)) + ((!g827) & (!g1299) & (!g1327) & (!g2640) & (g2669) & (g2641)) + ((!g827) & (!g1299) & (!g1327) & (g2640) & (g2669) & (!g2641)) + ((!g827) & (!g1299) & (!g1327) & (g2640) & (g2669) & (g2641)) + ((!g827) & (!g1299) & (g1327) & (!g2640) & (g2669) & (!g2641)) + ((!g827) & (!g1299) & (g1327) & (!g2640) & (g2669) & (g2641)) + ((!g827) & (!g1299) & (g1327) & (g2640) & (g2669) & (!g2641)) + ((!g827) & (!g1299) & (g1327) & (g2640) & (g2669) & (g2641)) + ((!g827) & (g1299) & (!g1327) & (!g2640) & (g2669) & (!g2641)) + ((!g827) & (g1299) & (!g1327) & (!g2640) & (g2669) & (g2641)) + ((!g827) & (g1299) & (!g1327) & (g2640) & (g2669) & (!g2641)) + ((!g827) & (g1299) & (!g1327) & (g2640) & (g2669) & (g2641)) + ((!g827) & (g1299) & (g1327) & (!g2640) & (g2669) & (!g2641)) + ((!g827) & (g1299) & (g1327) & (!g2640) & (g2669) & (g2641)) + ((!g827) & (g1299) & (g1327) & (g2640) & (g2669) & (!g2641)) + ((!g827) & (g1299) & (g1327) & (g2640) & (g2669) & (g2641)) + ((g827) & (!g1299) & (!g1327) & (!g2640) & (g2669) & (!g2641)) + ((g827) & (!g1299) & (!g1327) & (!g2640) & (g2669) & (g2641)) + ((g827) & (!g1299) & (!g1327) & (g2640) & (!g2669) & (g2641)) + ((g827) & (!g1299) & (!g1327) & (g2640) & (g2669) & (!g2641)) + ((g827) & (!g1299) & (g1327) & (!g2640) & (!g2669) & (!g2641)) + ((g827) & (!g1299) & (g1327) & (!g2640) & (!g2669) & (g2641)) + ((g827) & (!g1299) & (g1327) & (g2640) & (!g2669) & (!g2641)) + ((g827) & (!g1299) & (g1327) & (g2640) & (g2669) & (g2641)) + ((g827) & (g1299) & (!g1327) & (!g2640) & (!g2669) & (g2641)) + ((g827) & (g1299) & (!g1327) & (!g2640) & (g2669) & (!g2641)) + ((g827) & (g1299) & (!g1327) & (g2640) & (!g2669) & (!g2641)) + ((g827) & (g1299) & (!g1327) & (g2640) & (!g2669) & (g2641)) + ((g827) & (g1299) & (g1327) & (!g2640) & (!g2669) & (!g2641)) + ((g827) & (g1299) & (g1327) & (!g2640) & (g2669) & (g2641)) + ((g827) & (g1299) & (g1327) & (g2640) & (g2669) & (!g2641)) + ((g827) & (g1299) & (g1327) & (g2640) & (g2669) & (g2641)));
	assign g2671 = (((!g827) & (!g1277) & (!g1329) & (!g2014) & (g2052) & (!g2610)) + ((!g827) & (!g1277) & (!g1329) & (!g2014) & (g2052) & (g2610)) + ((!g827) & (!g1277) & (!g1329) & (g2014) & (g2052) & (!g2610)) + ((!g827) & (!g1277) & (!g1329) & (g2014) & (g2052) & (g2610)) + ((!g827) & (!g1277) & (g1329) & (!g2014) & (g2052) & (!g2610)) + ((!g827) & (!g1277) & (g1329) & (!g2014) & (g2052) & (g2610)) + ((!g827) & (!g1277) & (g1329) & (g2014) & (g2052) & (!g2610)) + ((!g827) & (!g1277) & (g1329) & (g2014) & (g2052) & (g2610)) + ((!g827) & (g1277) & (!g1329) & (!g2014) & (g2052) & (!g2610)) + ((!g827) & (g1277) & (!g1329) & (!g2014) & (g2052) & (g2610)) + ((!g827) & (g1277) & (!g1329) & (g2014) & (g2052) & (!g2610)) + ((!g827) & (g1277) & (!g1329) & (g2014) & (g2052) & (g2610)) + ((!g827) & (g1277) & (g1329) & (!g2014) & (g2052) & (!g2610)) + ((!g827) & (g1277) & (g1329) & (!g2014) & (g2052) & (g2610)) + ((!g827) & (g1277) & (g1329) & (g2014) & (g2052) & (!g2610)) + ((!g827) & (g1277) & (g1329) & (g2014) & (g2052) & (g2610)) + ((g827) & (!g1277) & (!g1329) & (!g2014) & (g2052) & (!g2610)) + ((g827) & (!g1277) & (!g1329) & (!g2014) & (g2052) & (g2610)) + ((g827) & (!g1277) & (!g1329) & (g2014) & (!g2052) & (g2610)) + ((g827) & (!g1277) & (!g1329) & (g2014) & (g2052) & (!g2610)) + ((g827) & (!g1277) & (g1329) & (!g2014) & (!g2052) & (!g2610)) + ((g827) & (!g1277) & (g1329) & (!g2014) & (!g2052) & (g2610)) + ((g827) & (!g1277) & (g1329) & (g2014) & (!g2052) & (!g2610)) + ((g827) & (!g1277) & (g1329) & (g2014) & (g2052) & (g2610)) + ((g827) & (g1277) & (!g1329) & (!g2014) & (!g2052) & (g2610)) + ((g827) & (g1277) & (!g1329) & (!g2014) & (g2052) & (!g2610)) + ((g827) & (g1277) & (!g1329) & (g2014) & (!g2052) & (!g2610)) + ((g827) & (g1277) & (!g1329) & (g2014) & (!g2052) & (g2610)) + ((g827) & (g1277) & (g1329) & (!g2014) & (!g2052) & (!g2610)) + ((g827) & (g1277) & (g1329) & (!g2014) & (g2052) & (g2610)) + ((g827) & (g1277) & (g1329) & (g2014) & (g2052) & (!g2610)) + ((g827) & (g1277) & (g1329) & (g2014) & (g2052) & (g2610)));
	assign g8085 = (((!g3464) & (g4914) & (!g2672)) + ((!g3464) & (g4914) & (g2672)) + ((g3464) & (!g4914) & (g2672)) + ((g3464) & (g4914) & (g2672)));
	assign g2673 = (((!g827) & (!g1285) & (!g1331) & (!g2620) & (g2672) & (!g2621)) + ((!g827) & (!g1285) & (!g1331) & (!g2620) & (g2672) & (g2621)) + ((!g827) & (!g1285) & (!g1331) & (g2620) & (g2672) & (!g2621)) + ((!g827) & (!g1285) & (!g1331) & (g2620) & (g2672) & (g2621)) + ((!g827) & (!g1285) & (g1331) & (!g2620) & (g2672) & (!g2621)) + ((!g827) & (!g1285) & (g1331) & (!g2620) & (g2672) & (g2621)) + ((!g827) & (!g1285) & (g1331) & (g2620) & (g2672) & (!g2621)) + ((!g827) & (!g1285) & (g1331) & (g2620) & (g2672) & (g2621)) + ((!g827) & (g1285) & (!g1331) & (!g2620) & (g2672) & (!g2621)) + ((!g827) & (g1285) & (!g1331) & (!g2620) & (g2672) & (g2621)) + ((!g827) & (g1285) & (!g1331) & (g2620) & (g2672) & (!g2621)) + ((!g827) & (g1285) & (!g1331) & (g2620) & (g2672) & (g2621)) + ((!g827) & (g1285) & (g1331) & (!g2620) & (g2672) & (!g2621)) + ((!g827) & (g1285) & (g1331) & (!g2620) & (g2672) & (g2621)) + ((!g827) & (g1285) & (g1331) & (g2620) & (g2672) & (!g2621)) + ((!g827) & (g1285) & (g1331) & (g2620) & (g2672) & (g2621)) + ((g827) & (!g1285) & (!g1331) & (!g2620) & (g2672) & (!g2621)) + ((g827) & (!g1285) & (!g1331) & (!g2620) & (g2672) & (g2621)) + ((g827) & (!g1285) & (!g1331) & (g2620) & (!g2672) & (g2621)) + ((g827) & (!g1285) & (!g1331) & (g2620) & (g2672) & (!g2621)) + ((g827) & (!g1285) & (g1331) & (!g2620) & (!g2672) & (!g2621)) + ((g827) & (!g1285) & (g1331) & (!g2620) & (!g2672) & (g2621)) + ((g827) & (!g1285) & (g1331) & (g2620) & (!g2672) & (!g2621)) + ((g827) & (!g1285) & (g1331) & (g2620) & (g2672) & (g2621)) + ((g827) & (g1285) & (!g1331) & (!g2620) & (!g2672) & (g2621)) + ((g827) & (g1285) & (!g1331) & (!g2620) & (g2672) & (!g2621)) + ((g827) & (g1285) & (!g1331) & (g2620) & (!g2672) & (!g2621)) + ((g827) & (g1285) & (!g1331) & (g2620) & (!g2672) & (g2621)) + ((g827) & (g1285) & (g1331) & (!g2620) & (!g2672) & (!g2621)) + ((g827) & (g1285) & (g1331) & (!g2620) & (g2672) & (g2621)) + ((g827) & (g1285) & (g1331) & (g2620) & (g2672) & (!g2621)) + ((g827) & (g1285) & (g1331) & (g2620) & (g2672) & (g2621)));
	assign g8086 = (((!g3429) & (g4919) & (!g2674)) + ((!g3429) & (g4919) & (g2674)) + ((g3429) & (!g4919) & (g2674)) + ((g3429) & (g4919) & (g2674)));
	assign g2675 = (((!g827) & (!g1293) & (!g1333) & (!g2632) & (g2674) & (!g2633)) + ((!g827) & (!g1293) & (!g1333) & (!g2632) & (g2674) & (g2633)) + ((!g827) & (!g1293) & (!g1333) & (g2632) & (g2674) & (!g2633)) + ((!g827) & (!g1293) & (!g1333) & (g2632) & (g2674) & (g2633)) + ((!g827) & (!g1293) & (g1333) & (!g2632) & (g2674) & (!g2633)) + ((!g827) & (!g1293) & (g1333) & (!g2632) & (g2674) & (g2633)) + ((!g827) & (!g1293) & (g1333) & (g2632) & (g2674) & (!g2633)) + ((!g827) & (!g1293) & (g1333) & (g2632) & (g2674) & (g2633)) + ((!g827) & (g1293) & (!g1333) & (!g2632) & (g2674) & (!g2633)) + ((!g827) & (g1293) & (!g1333) & (!g2632) & (g2674) & (g2633)) + ((!g827) & (g1293) & (!g1333) & (g2632) & (g2674) & (!g2633)) + ((!g827) & (g1293) & (!g1333) & (g2632) & (g2674) & (g2633)) + ((!g827) & (g1293) & (g1333) & (!g2632) & (g2674) & (!g2633)) + ((!g827) & (g1293) & (g1333) & (!g2632) & (g2674) & (g2633)) + ((!g827) & (g1293) & (g1333) & (g2632) & (g2674) & (!g2633)) + ((!g827) & (g1293) & (g1333) & (g2632) & (g2674) & (g2633)) + ((g827) & (!g1293) & (!g1333) & (!g2632) & (g2674) & (!g2633)) + ((g827) & (!g1293) & (!g1333) & (!g2632) & (g2674) & (g2633)) + ((g827) & (!g1293) & (!g1333) & (g2632) & (!g2674) & (g2633)) + ((g827) & (!g1293) & (!g1333) & (g2632) & (g2674) & (!g2633)) + ((g827) & (!g1293) & (g1333) & (!g2632) & (!g2674) & (!g2633)) + ((g827) & (!g1293) & (g1333) & (!g2632) & (!g2674) & (g2633)) + ((g827) & (!g1293) & (g1333) & (g2632) & (!g2674) & (!g2633)) + ((g827) & (!g1293) & (g1333) & (g2632) & (g2674) & (g2633)) + ((g827) & (g1293) & (!g1333) & (!g2632) & (!g2674) & (g2633)) + ((g827) & (g1293) & (!g1333) & (!g2632) & (g2674) & (!g2633)) + ((g827) & (g1293) & (!g1333) & (g2632) & (!g2674) & (!g2633)) + ((g827) & (g1293) & (!g1333) & (g2632) & (!g2674) & (g2633)) + ((g827) & (g1293) & (g1333) & (!g2632) & (!g2674) & (!g2633)) + ((g827) & (g1293) & (g1333) & (!g2632) & (g2674) & (g2633)) + ((g827) & (g1293) & (g1333) & (g2632) & (g2674) & (!g2633)) + ((g827) & (g1293) & (g1333) & (g2632) & (g2674) & (g2633)));
	assign g8087 = (((!g2017) & (g4923) & (!g2676)) + ((!g2017) & (g4923) & (g2676)) + ((g2017) & (!g4923) & (g2676)) + ((g2017) & (g4923) & (g2676)));
	assign g2677 = (((!g827) & (!g1301) & (!g1335) & (!g2643) & (g2676) & (!g2644)) + ((!g827) & (!g1301) & (!g1335) & (!g2643) & (g2676) & (g2644)) + ((!g827) & (!g1301) & (!g1335) & (g2643) & (g2676) & (!g2644)) + ((!g827) & (!g1301) & (!g1335) & (g2643) & (g2676) & (g2644)) + ((!g827) & (!g1301) & (g1335) & (!g2643) & (g2676) & (!g2644)) + ((!g827) & (!g1301) & (g1335) & (!g2643) & (g2676) & (g2644)) + ((!g827) & (!g1301) & (g1335) & (g2643) & (g2676) & (!g2644)) + ((!g827) & (!g1301) & (g1335) & (g2643) & (g2676) & (g2644)) + ((!g827) & (g1301) & (!g1335) & (!g2643) & (g2676) & (!g2644)) + ((!g827) & (g1301) & (!g1335) & (!g2643) & (g2676) & (g2644)) + ((!g827) & (g1301) & (!g1335) & (g2643) & (g2676) & (!g2644)) + ((!g827) & (g1301) & (!g1335) & (g2643) & (g2676) & (g2644)) + ((!g827) & (g1301) & (g1335) & (!g2643) & (g2676) & (!g2644)) + ((!g827) & (g1301) & (g1335) & (!g2643) & (g2676) & (g2644)) + ((!g827) & (g1301) & (g1335) & (g2643) & (g2676) & (!g2644)) + ((!g827) & (g1301) & (g1335) & (g2643) & (g2676) & (g2644)) + ((g827) & (!g1301) & (!g1335) & (!g2643) & (g2676) & (!g2644)) + ((g827) & (!g1301) & (!g1335) & (!g2643) & (g2676) & (g2644)) + ((g827) & (!g1301) & (!g1335) & (g2643) & (!g2676) & (g2644)) + ((g827) & (!g1301) & (!g1335) & (g2643) & (g2676) & (!g2644)) + ((g827) & (!g1301) & (g1335) & (!g2643) & (!g2676) & (!g2644)) + ((g827) & (!g1301) & (g1335) & (!g2643) & (!g2676) & (g2644)) + ((g827) & (!g1301) & (g1335) & (g2643) & (!g2676) & (!g2644)) + ((g827) & (!g1301) & (g1335) & (g2643) & (g2676) & (g2644)) + ((g827) & (g1301) & (!g1335) & (!g2643) & (!g2676) & (g2644)) + ((g827) & (g1301) & (!g1335) & (!g2643) & (g2676) & (!g2644)) + ((g827) & (g1301) & (!g1335) & (g2643) & (!g2676) & (!g2644)) + ((g827) & (g1301) & (!g1335) & (g2643) & (!g2676) & (g2644)) + ((g827) & (g1301) & (g1335) & (!g2643) & (!g2676) & (!g2644)) + ((g827) & (g1301) & (g1335) & (!g2643) & (g2676) & (g2644)) + ((g827) & (g1301) & (g1335) & (g2643) & (g2676) & (!g2644)) + ((g827) & (g1301) & (g1335) & (g2643) & (g2676) & (g2644)));
	assign g8088 = (((!g3429) & (g4926) & (!g2678)) + ((!g3429) & (g4926) & (g2678)) + ((g3429) & (!g4926) & (g2678)) + ((g3429) & (g4926) & (g2678)));
	assign g8089 = (((!g3464) & (g4929) & (!g2679)) + ((!g3464) & (g4929) & (g2679)) + ((g3464) & (!g4929) & (g2679)) + ((g3464) & (g4929) & (g2679)));
	assign g2680 = (((!g2649) & (g2650)) + ((g2649) & (!g2650)));
	assign g2681 = (((!g2554) & (!g2555) & (!g2556) & (g2601) & (g2602) & (g2680)) + ((!g2554) & (!g2555) & (g2556) & (g2601) & (g2602) & (g2680)) + ((!g2554) & (g2555) & (!g2556) & (g2601) & (g2602) & (g2680)) + ((!g2554) & (g2555) & (g2556) & (!g2601) & (g2602) & (g2680)) + ((!g2554) & (g2555) & (g2556) & (g2601) & (!g2602) & (g2680)) + ((!g2554) & (g2555) & (g2556) & (g2601) & (g2602) & (g2680)) + ((g2554) & (!g2555) & (!g2556) & (g2601) & (g2602) & (g2680)) + ((g2554) & (!g2555) & (g2556) & (!g2601) & (g2602) & (g2680)) + ((g2554) & (!g2555) & (g2556) & (g2601) & (!g2602) & (g2680)) + ((g2554) & (!g2555) & (g2556) & (g2601) & (g2602) & (g2680)) + ((g2554) & (g2555) & (!g2556) & (!g2601) & (g2602) & (g2680)) + ((g2554) & (g2555) & (!g2556) & (g2601) & (!g2602) & (g2680)) + ((g2554) & (g2555) & (!g2556) & (g2601) & (g2602) & (g2680)) + ((g2554) & (g2555) & (g2556) & (!g2601) & (g2602) & (g2680)) + ((g2554) & (g2555) & (g2556) & (g2601) & (!g2602) & (g2680)) + ((g2554) & (g2555) & (g2556) & (g2601) & (g2602) & (g2680)));
	assign g2682 = (((g2649) & (g2650)));
	assign g8090 = (((!g3429) & (g4932) & (!g2683)) + ((!g3429) & (g4932) & (g2683)) + ((g3429) & (!g4932) & (g2683)) + ((g3429) & (g4932) & (g2683)));
	assign g8091 = (((!g3499) & (g4935) & (!g2684)) + ((!g3499) & (g4935) & (g2684)) + ((g3499) & (!g4935) & (g2684)) + ((g3499) & (g4935) & (g2684)));
	assign g2685 = (((g830) & (!g1914) & (!g2681) & (!g5688) & (g5689) & (!g5690)) + ((g830) & (!g1914) & (!g2681) & (!g5688) & (g5689) & (g5690)) + ((g830) & (!g1914) & (!g2681) & (g5688) & (g5689) & (!g5690)) + ((g830) & (!g1914) & (!g2681) & (g5688) & (g5689) & (g5690)) + ((g830) & (!g1914) & (g2681) & (g5688) & (!g5689) & (!g5690)) + ((g830) & (!g1914) & (g2681) & (g5688) & (!g5689) & (g5690)) + ((g830) & (!g1914) & (g2681) & (g5688) & (g5689) & (!g5690)) + ((g830) & (!g1914) & (g2681) & (g5688) & (g5689) & (g5690)) + ((g830) & (g1914) & (!g2681) & (!g5688) & (!g5689) & (g5690)) + ((g830) & (g1914) & (!g2681) & (!g5688) & (g5689) & (g5690)) + ((g830) & (g1914) & (!g2681) & (g5688) & (!g5689) & (g5690)) + ((g830) & (g1914) & (!g2681) & (g5688) & (g5689) & (g5690)) + ((g830) & (g1914) & (g2681) & (!g5688) & (!g5689) & (g5690)) + ((g830) & (g1914) & (g2681) & (!g5688) & (g5689) & (g5690)) + ((g830) & (g1914) & (g2681) & (g5688) & (!g5689) & (g5690)) + ((g830) & (g1914) & (g2681) & (g5688) & (g5689) & (g5690)));
	assign g2686 = (((!g1175) & (!g2003) & (!g2446) & (!g2447) & (!g5735) & (g5736)) + ((!g1175) & (!g2003) & (!g2446) & (g2447) & (!g5735) & (g5736)) + ((!g1175) & (!g2003) & (g2446) & (!g2447) & (!g5735) & (g5736)) + ((!g1175) & (!g2003) & (g2446) & (g2447) & (!g5735) & (g5736)) + ((!g1175) & (g2003) & (!g2446) & (!g2447) & (!g5735) & (g5736)) + ((!g1175) & (g2003) & (!g2446) & (g2447) & (!g5735) & (g5736)) + ((!g1175) & (g2003) & (!g2446) & (g2447) & (g5735) & (g5736)) + ((!g1175) & (g2003) & (g2446) & (!g2447) & (!g5735) & (g5736)) + ((!g1175) & (g2003) & (g2446) & (!g2447) & (g5735) & (g5736)) + ((!g1175) & (g2003) & (g2446) & (g2447) & (!g5735) & (g5736)) + ((!g1175) & (g2003) & (g2446) & (g2447) & (g5735) & (g5736)) + ((g1175) & (!g2003) & (!g2446) & (!g2447) & (!g5735) & (g5736)) + ((g1175) & (!g2003) & (!g2446) & (g2447) & (!g5735) & (g5736)) + ((g1175) & (!g2003) & (!g2446) & (g2447) & (g5735) & (g5736)) + ((g1175) & (!g2003) & (g2446) & (!g2447) & (!g5735) & (g5736)) + ((g1175) & (!g2003) & (g2446) & (!g2447) & (g5735) & (g5736)) + ((g1175) & (!g2003) & (g2446) & (g2447) & (!g5735) & (g5736)) + ((g1175) & (!g2003) & (g2446) & (g2447) & (g5735) & (g5736)) + ((g1175) & (g2003) & (!g2446) & (!g2447) & (!g5735) & (g5736)) + ((g1175) & (g2003) & (!g2446) & (!g2447) & (g5735) & (g5736)) + ((g1175) & (g2003) & (!g2446) & (g2447) & (!g5735) & (g5736)) + ((g1175) & (g2003) & (!g2446) & (g2447) & (g5735) & (g5736)) + ((g1175) & (g2003) & (g2446) & (!g2447) & (!g5735) & (g5736)) + ((g1175) & (g2003) & (g2446) & (!g2447) & (g5735) & (g5736)) + ((g1175) & (g2003) & (g2446) & (g2447) & (!g5735) & (g5736)) + ((g1175) & (g2003) & (g2446) & (g2447) & (g5735) & (g5736)));
	assign g2687 = (((g1313) & (g2051)));
	assign g2688 = (((!g2686) & (!g2687)));
	assign g2689 = (((!g827) & (!g1340) & (g2100) & (!g2688)) + ((!g827) & (!g1340) & (g2100) & (g2688)) + ((!g827) & (g1340) & (g2100) & (!g2688)) + ((!g827) & (g1340) & (g2100) & (g2688)) + ((g827) & (!g1340) & (!g2100) & (!g2688)) + ((g827) & (!g1340) & (g2100) & (g2688)) + ((g827) & (g1340) & (!g2100) & (g2688)) + ((g827) & (g1340) & (g2100) & (!g2688)));
	assign g8092 = (((!g3464) & (g4939) & (!g2690)) + ((!g3464) & (g4939) & (g2690)) + ((g3464) & (!g4939) & (g2690)) + ((g3464) & (g4939) & (g2690)));
	assign g2691 = (((!g1183) & (!g2468) & (!g2470) & (!g2471) & (!g5747) & (g5748)) + ((!g1183) & (!g2468) & (!g2470) & (g2471) & (!g5747) & (g5748)) + ((!g1183) & (!g2468) & (g2470) & (!g2471) & (!g5747) & (g5748)) + ((!g1183) & (!g2468) & (g2470) & (g2471) & (!g5747) & (g5748)) + ((!g1183) & (g2468) & (!g2470) & (!g2471) & (!g5747) & (g5748)) + ((!g1183) & (g2468) & (!g2470) & (g2471) & (!g5747) & (g5748)) + ((!g1183) & (g2468) & (!g2470) & (g2471) & (g5747) & (g5748)) + ((!g1183) & (g2468) & (g2470) & (!g2471) & (!g5747) & (g5748)) + ((!g1183) & (g2468) & (g2470) & (!g2471) & (g5747) & (g5748)) + ((!g1183) & (g2468) & (g2470) & (g2471) & (!g5747) & (g5748)) + ((!g1183) & (g2468) & (g2470) & (g2471) & (g5747) & (g5748)) + ((g1183) & (!g2468) & (!g2470) & (!g2471) & (!g5747) & (g5748)) + ((g1183) & (!g2468) & (!g2470) & (g2471) & (!g5747) & (g5748)) + ((g1183) & (!g2468) & (!g2470) & (g2471) & (g5747) & (g5748)) + ((g1183) & (!g2468) & (g2470) & (!g2471) & (!g5747) & (g5748)) + ((g1183) & (!g2468) & (g2470) & (!g2471) & (g5747) & (g5748)) + ((g1183) & (!g2468) & (g2470) & (g2471) & (!g5747) & (g5748)) + ((g1183) & (!g2468) & (g2470) & (g2471) & (g5747) & (g5748)) + ((g1183) & (g2468) & (!g2470) & (!g2471) & (!g5747) & (g5748)) + ((g1183) & (g2468) & (!g2470) & (!g2471) & (g5747) & (g5748)) + ((g1183) & (g2468) & (!g2470) & (g2471) & (!g5747) & (g5748)) + ((g1183) & (g2468) & (!g2470) & (g2471) & (g5747) & (g5748)) + ((g1183) & (g2468) & (g2470) & (!g2471) & (!g5747) & (g5748)) + ((g1183) & (g2468) & (g2470) & (!g2471) & (g5747) & (g5748)) + ((g1183) & (g2468) & (g2470) & (g2471) & (!g5747) & (g5748)) + ((g1183) & (g2468) & (g2470) & (g2471) & (g5747) & (g5748)));
	assign g2692 = (((g1321) & (g2663)));
	assign g2693 = (((!g2691) & (!g2692)));
	assign g2694 = (((!g827) & (!g1342) & (g2690) & (!g2693)) + ((!g827) & (!g1342) & (g2690) & (g2693)) + ((!g827) & (g1342) & (g2690) & (!g2693)) + ((!g827) & (g1342) & (g2690) & (g2693)) + ((g827) & (!g1342) & (!g2690) & (!g2693)) + ((g827) & (!g1342) & (g2690) & (g2693)) + ((g827) & (g1342) & (!g2690) & (g2693)) + ((g827) & (g1342) & (g2690) & (!g2693)));
	assign g2695 = (((!g1191) & (!g2004) & (!g2493) & (!g2494) & (!g5759) & (g5760)) + ((!g1191) & (!g2004) & (!g2493) & (g2494) & (!g5759) & (g5760)) + ((!g1191) & (!g2004) & (g2493) & (!g2494) & (!g5759) & (g5760)) + ((!g1191) & (!g2004) & (g2493) & (g2494) & (!g5759) & (g5760)) + ((!g1191) & (g2004) & (!g2493) & (!g2494) & (!g5759) & (g5760)) + ((!g1191) & (g2004) & (!g2493) & (g2494) & (!g5759) & (g5760)) + ((!g1191) & (g2004) & (!g2493) & (g2494) & (g5759) & (g5760)) + ((!g1191) & (g2004) & (g2493) & (!g2494) & (!g5759) & (g5760)) + ((!g1191) & (g2004) & (g2493) & (!g2494) & (g5759) & (g5760)) + ((!g1191) & (g2004) & (g2493) & (g2494) & (!g5759) & (g5760)) + ((!g1191) & (g2004) & (g2493) & (g2494) & (g5759) & (g5760)) + ((g1191) & (!g2004) & (!g2493) & (!g2494) & (!g5759) & (g5760)) + ((g1191) & (!g2004) & (!g2493) & (g2494) & (!g5759) & (g5760)) + ((g1191) & (!g2004) & (!g2493) & (g2494) & (g5759) & (g5760)) + ((g1191) & (!g2004) & (g2493) & (!g2494) & (!g5759) & (g5760)) + ((g1191) & (!g2004) & (g2493) & (!g2494) & (g5759) & (g5760)) + ((g1191) & (!g2004) & (g2493) & (g2494) & (!g5759) & (g5760)) + ((g1191) & (!g2004) & (g2493) & (g2494) & (g5759) & (g5760)) + ((g1191) & (g2004) & (!g2493) & (!g2494) & (!g5759) & (g5760)) + ((g1191) & (g2004) & (!g2493) & (!g2494) & (g5759) & (g5760)) + ((g1191) & (g2004) & (!g2493) & (g2494) & (!g5759) & (g5760)) + ((g1191) & (g2004) & (!g2493) & (g2494) & (g5759) & (g5760)) + ((g1191) & (g2004) & (g2493) & (!g2494) & (!g5759) & (g5760)) + ((g1191) & (g2004) & (g2493) & (!g2494) & (g5759) & (g5760)) + ((g1191) & (g2004) & (g2493) & (g2494) & (!g5759) & (g5760)) + ((g1191) & (g2004) & (g2493) & (g2494) & (g5759) & (g5760)));
	assign g2696 = (((g1329) & (g2052)));
	assign g2697 = (((!g2695) & (!g2696)));
	assign g2698 = (((!g827) & (!g1344) & (g2101) & (!g2697)) + ((!g827) & (!g1344) & (g2101) & (g2697)) + ((!g827) & (g1344) & (g2101) & (!g2697)) + ((!g827) & (g1344) & (g2101) & (g2697)) + ((g827) & (!g1344) & (!g2101) & (!g2697)) + ((g827) & (!g1344) & (g2101) & (g2697)) + ((g827) & (g1344) & (!g2101) & (g2697)) + ((g827) & (g1344) & (g2101) & (!g2697)));
	assign g2699 = (((!g1169) & (!g1967) & (!g2430) & (!g2431) & (!g5726) & (g5727)) + ((!g1169) & (!g1967) & (!g2430) & (g2431) & (!g5726) & (g5727)) + ((!g1169) & (!g1967) & (g2430) & (!g2431) & (!g5726) & (g5727)) + ((!g1169) & (!g1967) & (g2430) & (g2431) & (!g5726) & (g5727)) + ((!g1169) & (g1967) & (!g2430) & (!g2431) & (!g5726) & (g5727)) + ((!g1169) & (g1967) & (!g2430) & (g2431) & (!g5726) & (g5727)) + ((!g1169) & (g1967) & (!g2430) & (g2431) & (g5726) & (g5727)) + ((!g1169) & (g1967) & (g2430) & (!g2431) & (!g5726) & (g5727)) + ((!g1169) & (g1967) & (g2430) & (!g2431) & (g5726) & (g5727)) + ((!g1169) & (g1967) & (g2430) & (g2431) & (!g5726) & (g5727)) + ((!g1169) & (g1967) & (g2430) & (g2431) & (g5726) & (g5727)) + ((g1169) & (!g1967) & (!g2430) & (!g2431) & (!g5726) & (g5727)) + ((g1169) & (!g1967) & (!g2430) & (g2431) & (!g5726) & (g5727)) + ((g1169) & (!g1967) & (!g2430) & (g2431) & (g5726) & (g5727)) + ((g1169) & (!g1967) & (g2430) & (!g2431) & (!g5726) & (g5727)) + ((g1169) & (!g1967) & (g2430) & (!g2431) & (g5726) & (g5727)) + ((g1169) & (!g1967) & (g2430) & (g2431) & (!g5726) & (g5727)) + ((g1169) & (!g1967) & (g2430) & (g2431) & (g5726) & (g5727)) + ((g1169) & (g1967) & (!g2430) & (!g2431) & (!g5726) & (g5727)) + ((g1169) & (g1967) & (!g2430) & (!g2431) & (g5726) & (g5727)) + ((g1169) & (g1967) & (!g2430) & (g2431) & (!g5726) & (g5727)) + ((g1169) & (g1967) & (!g2430) & (g2431) & (g5726) & (g5727)) + ((g1169) & (g1967) & (g2430) & (!g2431) & (!g5726) & (g5727)) + ((g1169) & (g1967) & (g2430) & (!g2431) & (g5726) & (g5727)) + ((g1169) & (g1967) & (g2430) & (g2431) & (!g5726) & (g5727)) + ((g1169) & (g1967) & (g2430) & (g2431) & (g5726) & (g5727)));
	assign g2700 = (((g1307) & (g2047)));
	assign g2701 = (((!g2699) & (!g2700)));
	assign g2702 = (((!g827) & (!g1346) & (g2098) & (!g2701)) + ((!g827) & (!g1346) & (g2098) & (g2701)) + ((!g827) & (g1346) & (g2098) & (!g2701)) + ((!g827) & (g1346) & (g2098) & (g2701)) + ((g827) & (!g1346) & (!g2098) & (!g2701)) + ((g827) & (!g1346) & (g2098) & (g2701)) + ((g827) & (g1346) & (!g2098) & (g2701)) + ((g827) & (g1346) & (g2098) & (!g2701)));
	assign g8093 = (((!g2017) & (g4943) & (!g2703)) + ((!g2017) & (g4943) & (g2703)) + ((g2017) & (!g4943) & (g2703)) + ((g2017) & (g4943) & (g2703)));
	assign g2704 = (((!g1177) & (!g2450) & (!g2452) & (!g2453) & (!g5738) & (g5739)) + ((!g1177) & (!g2450) & (!g2452) & (g2453) & (!g5738) & (g5739)) + ((!g1177) & (!g2450) & (g2452) & (!g2453) & (!g5738) & (g5739)) + ((!g1177) & (!g2450) & (g2452) & (g2453) & (!g5738) & (g5739)) + ((!g1177) & (g2450) & (!g2452) & (!g2453) & (!g5738) & (g5739)) + ((!g1177) & (g2450) & (!g2452) & (g2453) & (!g5738) & (g5739)) + ((!g1177) & (g2450) & (!g2452) & (g2453) & (g5738) & (g5739)) + ((!g1177) & (g2450) & (g2452) & (!g2453) & (!g5738) & (g5739)) + ((!g1177) & (g2450) & (g2452) & (!g2453) & (g5738) & (g5739)) + ((!g1177) & (g2450) & (g2452) & (g2453) & (!g5738) & (g5739)) + ((!g1177) & (g2450) & (g2452) & (g2453) & (g5738) & (g5739)) + ((g1177) & (!g2450) & (!g2452) & (!g2453) & (!g5738) & (g5739)) + ((g1177) & (!g2450) & (!g2452) & (g2453) & (!g5738) & (g5739)) + ((g1177) & (!g2450) & (!g2452) & (g2453) & (g5738) & (g5739)) + ((g1177) & (!g2450) & (g2452) & (!g2453) & (!g5738) & (g5739)) + ((g1177) & (!g2450) & (g2452) & (!g2453) & (g5738) & (g5739)) + ((g1177) & (!g2450) & (g2452) & (g2453) & (!g5738) & (g5739)) + ((g1177) & (!g2450) & (g2452) & (g2453) & (g5738) & (g5739)) + ((g1177) & (g2450) & (!g2452) & (!g2453) & (!g5738) & (g5739)) + ((g1177) & (g2450) & (!g2452) & (!g2453) & (g5738) & (g5739)) + ((g1177) & (g2450) & (!g2452) & (g2453) & (!g5738) & (g5739)) + ((g1177) & (g2450) & (!g2452) & (g2453) & (g5738) & (g5739)) + ((g1177) & (g2450) & (g2452) & (!g2453) & (!g5738) & (g5739)) + ((g1177) & (g2450) & (g2452) & (!g2453) & (g5738) & (g5739)) + ((g1177) & (g2450) & (g2452) & (g2453) & (!g5738) & (g5739)) + ((g1177) & (g2450) & (g2452) & (g2453) & (g5738) & (g5739)));
	assign g2705 = (((g1315) & (g2657)));
	assign g2706 = (((!g2704) & (!g2705)));
	assign g2707 = (((!g827) & (!g1348) & (g2703) & (!g2706)) + ((!g827) & (!g1348) & (g2703) & (g2706)) + ((!g827) & (g1348) & (g2703) & (!g2706)) + ((!g827) & (g1348) & (g2703) & (g2706)) + ((g827) & (!g1348) & (!g2703) & (!g2706)) + ((g827) & (!g1348) & (g2703) & (g2706)) + ((g827) & (g1348) & (!g2703) & (g2706)) + ((g827) & (g1348) & (g2703) & (!g2706)));
	assign g8094 = (((!g3499) & (g4947) & (!g2708)) + ((!g3499) & (g4947) & (g2708)) + ((g3499) & (!g4947) & (g2708)) + ((g3499) & (g4947) & (g2708)));
	assign g2709 = (((!g1185) & (!g2474) & (!g2476) & (!g2477) & (!g5750) & (g5751)) + ((!g1185) & (!g2474) & (!g2476) & (g2477) & (!g5750) & (g5751)) + ((!g1185) & (!g2474) & (g2476) & (!g2477) & (!g5750) & (g5751)) + ((!g1185) & (!g2474) & (g2476) & (g2477) & (!g5750) & (g5751)) + ((!g1185) & (g2474) & (!g2476) & (!g2477) & (!g5750) & (g5751)) + ((!g1185) & (g2474) & (!g2476) & (g2477) & (!g5750) & (g5751)) + ((!g1185) & (g2474) & (!g2476) & (g2477) & (g5750) & (g5751)) + ((!g1185) & (g2474) & (g2476) & (!g2477) & (!g5750) & (g5751)) + ((!g1185) & (g2474) & (g2476) & (!g2477) & (g5750) & (g5751)) + ((!g1185) & (g2474) & (g2476) & (g2477) & (!g5750) & (g5751)) + ((!g1185) & (g2474) & (g2476) & (g2477) & (g5750) & (g5751)) + ((g1185) & (!g2474) & (!g2476) & (!g2477) & (!g5750) & (g5751)) + ((g1185) & (!g2474) & (!g2476) & (g2477) & (!g5750) & (g5751)) + ((g1185) & (!g2474) & (!g2476) & (g2477) & (g5750) & (g5751)) + ((g1185) & (!g2474) & (g2476) & (!g2477) & (!g5750) & (g5751)) + ((g1185) & (!g2474) & (g2476) & (!g2477) & (g5750) & (g5751)) + ((g1185) & (!g2474) & (g2476) & (g2477) & (!g5750) & (g5751)) + ((g1185) & (!g2474) & (g2476) & (g2477) & (g5750) & (g5751)) + ((g1185) & (g2474) & (!g2476) & (!g2477) & (!g5750) & (g5751)) + ((g1185) & (g2474) & (!g2476) & (!g2477) & (g5750) & (g5751)) + ((g1185) & (g2474) & (!g2476) & (g2477) & (!g5750) & (g5751)) + ((g1185) & (g2474) & (!g2476) & (g2477) & (g5750) & (g5751)) + ((g1185) & (g2474) & (g2476) & (!g2477) & (!g5750) & (g5751)) + ((g1185) & (g2474) & (g2476) & (!g2477) & (g5750) & (g5751)) + ((g1185) & (g2474) & (g2476) & (g2477) & (!g5750) & (g5751)) + ((g1185) & (g2474) & (g2476) & (g2477) & (g5750) & (g5751)));
	assign g2710 = (((g1323) & (g2665)));
	assign g2711 = (((!g2709) & (!g2710)));
	assign g2712 = (((!g827) & (!g1350) & (g2708) & (!g2711)) + ((!g827) & (!g1350) & (g2708) & (g2711)) + ((!g827) & (g1350) & (g2708) & (!g2711)) + ((!g827) & (g1350) & (g2708) & (g2711)) + ((g827) & (!g1350) & (!g2708) & (!g2711)) + ((g827) & (!g1350) & (g2708) & (g2711)) + ((g827) & (g1350) & (!g2708) & (g2711)) + ((g827) & (g1350) & (g2708) & (!g2711)));
	assign g8095 = (((!g3464) & (g4951) & (!g2713)) + ((!g3464) & (g4951) & (g2713)) + ((g3464) & (!g4951) & (g2713)) + ((g3464) & (g4951) & (g2713)));
	assign g2714 = (((!g1193) & (!g2497) & (!g2499) & (!g2500) & (!g5762) & (g5763)) + ((!g1193) & (!g2497) & (!g2499) & (g2500) & (!g5762) & (g5763)) + ((!g1193) & (!g2497) & (g2499) & (!g2500) & (!g5762) & (g5763)) + ((!g1193) & (!g2497) & (g2499) & (g2500) & (!g5762) & (g5763)) + ((!g1193) & (g2497) & (!g2499) & (!g2500) & (!g5762) & (g5763)) + ((!g1193) & (g2497) & (!g2499) & (g2500) & (!g5762) & (g5763)) + ((!g1193) & (g2497) & (!g2499) & (g2500) & (g5762) & (g5763)) + ((!g1193) & (g2497) & (g2499) & (!g2500) & (!g5762) & (g5763)) + ((!g1193) & (g2497) & (g2499) & (!g2500) & (g5762) & (g5763)) + ((!g1193) & (g2497) & (g2499) & (g2500) & (!g5762) & (g5763)) + ((!g1193) & (g2497) & (g2499) & (g2500) & (g5762) & (g5763)) + ((g1193) & (!g2497) & (!g2499) & (!g2500) & (!g5762) & (g5763)) + ((g1193) & (!g2497) & (!g2499) & (g2500) & (!g5762) & (g5763)) + ((g1193) & (!g2497) & (!g2499) & (g2500) & (g5762) & (g5763)) + ((g1193) & (!g2497) & (g2499) & (!g2500) & (!g5762) & (g5763)) + ((g1193) & (!g2497) & (g2499) & (!g2500) & (g5762) & (g5763)) + ((g1193) & (!g2497) & (g2499) & (g2500) & (!g5762) & (g5763)) + ((g1193) & (!g2497) & (g2499) & (g2500) & (g5762) & (g5763)) + ((g1193) & (g2497) & (!g2499) & (!g2500) & (!g5762) & (g5763)) + ((g1193) & (g2497) & (!g2499) & (!g2500) & (g5762) & (g5763)) + ((g1193) & (g2497) & (!g2499) & (g2500) & (!g5762) & (g5763)) + ((g1193) & (g2497) & (!g2499) & (g2500) & (g5762) & (g5763)) + ((g1193) & (g2497) & (g2499) & (!g2500) & (!g5762) & (g5763)) + ((g1193) & (g2497) & (g2499) & (!g2500) & (g5762) & (g5763)) + ((g1193) & (g2497) & (g2499) & (g2500) & (!g5762) & (g5763)) + ((g1193) & (g2497) & (g2499) & (g2500) & (g5762) & (g5763)));
	assign g2715 = (((g1331) & (g2672)));
	assign g2716 = (((!g2714) & (!g2715)));
	assign g2717 = (((!g827) & (!g1352) & (g2713) & (!g2716)) + ((!g827) & (!g1352) & (g2713) & (g2716)) + ((!g827) & (g1352) & (g2713) & (!g2716)) + ((!g827) & (g1352) & (g2713) & (g2716)) + ((g827) & (!g1352) & (!g2713) & (!g2716)) + ((g827) & (!g1352) & (g2713) & (g2716)) + ((g827) & (g1352) & (!g2713) & (g2716)) + ((g827) & (g1352) & (g2713) & (!g2716)));
	assign g8096 = (((!g3499) & (g4955) & (!g2718)) + ((!g3499) & (g4955) & (g2718)) + ((g3499) & (!g4955) & (g2718)) + ((g3499) & (g4955) & (g2718)));
	assign g2719 = (((!g1171) & (!g2434) & (!g2436) & (!g2437) & (!g5729) & (g5730)) + ((!g1171) & (!g2434) & (!g2436) & (g2437) & (!g5729) & (g5730)) + ((!g1171) & (!g2434) & (g2436) & (!g2437) & (!g5729) & (g5730)) + ((!g1171) & (!g2434) & (g2436) & (g2437) & (!g5729) & (g5730)) + ((!g1171) & (g2434) & (!g2436) & (!g2437) & (!g5729) & (g5730)) + ((!g1171) & (g2434) & (!g2436) & (g2437) & (!g5729) & (g5730)) + ((!g1171) & (g2434) & (!g2436) & (g2437) & (g5729) & (g5730)) + ((!g1171) & (g2434) & (g2436) & (!g2437) & (!g5729) & (g5730)) + ((!g1171) & (g2434) & (g2436) & (!g2437) & (g5729) & (g5730)) + ((!g1171) & (g2434) & (g2436) & (g2437) & (!g5729) & (g5730)) + ((!g1171) & (g2434) & (g2436) & (g2437) & (g5729) & (g5730)) + ((g1171) & (!g2434) & (!g2436) & (!g2437) & (!g5729) & (g5730)) + ((g1171) & (!g2434) & (!g2436) & (g2437) & (!g5729) & (g5730)) + ((g1171) & (!g2434) & (!g2436) & (g2437) & (g5729) & (g5730)) + ((g1171) & (!g2434) & (g2436) & (!g2437) & (!g5729) & (g5730)) + ((g1171) & (!g2434) & (g2436) & (!g2437) & (g5729) & (g5730)) + ((g1171) & (!g2434) & (g2436) & (g2437) & (!g5729) & (g5730)) + ((g1171) & (!g2434) & (g2436) & (g2437) & (g5729) & (g5730)) + ((g1171) & (g2434) & (!g2436) & (!g2437) & (!g5729) & (g5730)) + ((g1171) & (g2434) & (!g2436) & (!g2437) & (g5729) & (g5730)) + ((g1171) & (g2434) & (!g2436) & (g2437) & (!g5729) & (g5730)) + ((g1171) & (g2434) & (!g2436) & (g2437) & (g5729) & (g5730)) + ((g1171) & (g2434) & (g2436) & (!g2437) & (!g5729) & (g5730)) + ((g1171) & (g2434) & (g2436) & (!g2437) & (g5729) & (g5730)) + ((g1171) & (g2434) & (g2436) & (g2437) & (!g5729) & (g5730)) + ((g1171) & (g2434) & (g2436) & (g2437) & (g5729) & (g5730)));
	assign g2720 = (((g1309) & (g2653)));
	assign g2721 = (((!g2719) & (!g2720)));
	assign g2722 = (((!g827) & (!g1354) & (g2718) & (!g2721)) + ((!g827) & (!g1354) & (g2718) & (g2721)) + ((!g827) & (g1354) & (g2718) & (!g2721)) + ((!g827) & (g1354) & (g2718) & (g2721)) + ((g827) & (!g1354) & (!g2718) & (!g2721)) + ((g827) & (!g1354) & (g2718) & (g2721)) + ((g827) & (g1354) & (!g2718) & (g2721)) + ((g827) & (g1354) & (g2718) & (!g2721)));
	assign g8097 = (((!g3464) & (g4960) & (!g2723)) + ((!g3464) & (g4960) & (g2723)) + ((g3464) & (!g4960) & (g2723)) + ((g3464) & (g4960) & (g2723)));
	assign g2724 = (((!g1179) & (!g2456) & (!g2458) & (!g2459) & (!g5741) & (g5742)) + ((!g1179) & (!g2456) & (!g2458) & (g2459) & (!g5741) & (g5742)) + ((!g1179) & (!g2456) & (g2458) & (!g2459) & (!g5741) & (g5742)) + ((!g1179) & (!g2456) & (g2458) & (g2459) & (!g5741) & (g5742)) + ((!g1179) & (g2456) & (!g2458) & (!g2459) & (!g5741) & (g5742)) + ((!g1179) & (g2456) & (!g2458) & (g2459) & (!g5741) & (g5742)) + ((!g1179) & (g2456) & (!g2458) & (g2459) & (g5741) & (g5742)) + ((!g1179) & (g2456) & (g2458) & (!g2459) & (!g5741) & (g5742)) + ((!g1179) & (g2456) & (g2458) & (!g2459) & (g5741) & (g5742)) + ((!g1179) & (g2456) & (g2458) & (g2459) & (!g5741) & (g5742)) + ((!g1179) & (g2456) & (g2458) & (g2459) & (g5741) & (g5742)) + ((g1179) & (!g2456) & (!g2458) & (!g2459) & (!g5741) & (g5742)) + ((g1179) & (!g2456) & (!g2458) & (g2459) & (!g5741) & (g5742)) + ((g1179) & (!g2456) & (!g2458) & (g2459) & (g5741) & (g5742)) + ((g1179) & (!g2456) & (g2458) & (!g2459) & (!g5741) & (g5742)) + ((g1179) & (!g2456) & (g2458) & (!g2459) & (g5741) & (g5742)) + ((g1179) & (!g2456) & (g2458) & (g2459) & (!g5741) & (g5742)) + ((g1179) & (!g2456) & (g2458) & (g2459) & (g5741) & (g5742)) + ((g1179) & (g2456) & (!g2458) & (!g2459) & (!g5741) & (g5742)) + ((g1179) & (g2456) & (!g2458) & (!g2459) & (g5741) & (g5742)) + ((g1179) & (g2456) & (!g2458) & (g2459) & (!g5741) & (g5742)) + ((g1179) & (g2456) & (!g2458) & (g2459) & (g5741) & (g5742)) + ((g1179) & (g2456) & (g2458) & (!g2459) & (!g5741) & (g5742)) + ((g1179) & (g2456) & (g2458) & (!g2459) & (g5741) & (g5742)) + ((g1179) & (g2456) & (g2458) & (g2459) & (!g5741) & (g5742)) + ((g1179) & (g2456) & (g2458) & (g2459) & (g5741) & (g5742)));
	assign g2725 = (((g1317) & (g2659)));
	assign g2726 = (((!g2724) & (!g2725)));
	assign g2727 = (((!g827) & (!g1356) & (g2723) & (!g2726)) + ((!g827) & (!g1356) & (g2723) & (g2726)) + ((!g827) & (g1356) & (g2723) & (!g2726)) + ((!g827) & (g1356) & (g2723) & (g2726)) + ((g827) & (!g1356) & (!g2723) & (!g2726)) + ((g827) & (!g1356) & (g2723) & (g2726)) + ((g827) & (g1356) & (!g2723) & (g2726)) + ((g827) & (g1356) & (g2723) & (!g2726)));
	assign g8098 = (((!g2017) & (g4964) & (!g2728)) + ((!g2017) & (g4964) & (g2728)) + ((g2017) & (!g4964) & (g2728)) + ((g2017) & (g4964) & (g2728)));
	assign g2729 = (((!g1187) & (!g2480) & (!g2482) & (!g2483) & (!g5753) & (g5754)) + ((!g1187) & (!g2480) & (!g2482) & (g2483) & (!g5753) & (g5754)) + ((!g1187) & (!g2480) & (g2482) & (!g2483) & (!g5753) & (g5754)) + ((!g1187) & (!g2480) & (g2482) & (g2483) & (!g5753) & (g5754)) + ((!g1187) & (g2480) & (!g2482) & (!g2483) & (!g5753) & (g5754)) + ((!g1187) & (g2480) & (!g2482) & (g2483) & (!g5753) & (g5754)) + ((!g1187) & (g2480) & (!g2482) & (g2483) & (g5753) & (g5754)) + ((!g1187) & (g2480) & (g2482) & (!g2483) & (!g5753) & (g5754)) + ((!g1187) & (g2480) & (g2482) & (!g2483) & (g5753) & (g5754)) + ((!g1187) & (g2480) & (g2482) & (g2483) & (!g5753) & (g5754)) + ((!g1187) & (g2480) & (g2482) & (g2483) & (g5753) & (g5754)) + ((g1187) & (!g2480) & (!g2482) & (!g2483) & (!g5753) & (g5754)) + ((g1187) & (!g2480) & (!g2482) & (g2483) & (!g5753) & (g5754)) + ((g1187) & (!g2480) & (!g2482) & (g2483) & (g5753) & (g5754)) + ((g1187) & (!g2480) & (g2482) & (!g2483) & (!g5753) & (g5754)) + ((g1187) & (!g2480) & (g2482) & (!g2483) & (g5753) & (g5754)) + ((g1187) & (!g2480) & (g2482) & (g2483) & (!g5753) & (g5754)) + ((g1187) & (!g2480) & (g2482) & (g2483) & (g5753) & (g5754)) + ((g1187) & (g2480) & (!g2482) & (!g2483) & (!g5753) & (g5754)) + ((g1187) & (g2480) & (!g2482) & (!g2483) & (g5753) & (g5754)) + ((g1187) & (g2480) & (!g2482) & (g2483) & (!g5753) & (g5754)) + ((g1187) & (g2480) & (!g2482) & (g2483) & (g5753) & (g5754)) + ((g1187) & (g2480) & (g2482) & (!g2483) & (!g5753) & (g5754)) + ((g1187) & (g2480) & (g2482) & (!g2483) & (g5753) & (g5754)) + ((g1187) & (g2480) & (g2482) & (g2483) & (!g5753) & (g5754)) + ((g1187) & (g2480) & (g2482) & (g2483) & (g5753) & (g5754)));
	assign g2730 = (((g1325) & (g2667)));
	assign g2731 = (((!g2729) & (!g2730)));
	assign g2732 = (((!g827) & (!g1358) & (g2728) & (!g2731)) + ((!g827) & (!g1358) & (g2728) & (g2731)) + ((!g827) & (g1358) & (g2728) & (!g2731)) + ((!g827) & (g1358) & (g2728) & (g2731)) + ((g827) & (!g1358) & (!g2728) & (!g2731)) + ((g827) & (!g1358) & (g2728) & (g2731)) + ((g827) & (g1358) & (!g2728) & (g2731)) + ((g827) & (g1358) & (g2728) & (!g2731)));
	assign g8099 = (((!g3429) & (g4967) & (!g2733)) + ((!g3429) & (g4967) & (g2733)) + ((g3429) & (!g4967) & (g2733)) + ((g3429) & (g4967) & (g2733)));
	assign g2734 = (((!g1195) & (!g2503) & (!g2505) & (!g2506) & (!g5765) & (g5766)) + ((!g1195) & (!g2503) & (!g2505) & (g2506) & (!g5765) & (g5766)) + ((!g1195) & (!g2503) & (g2505) & (!g2506) & (!g5765) & (g5766)) + ((!g1195) & (!g2503) & (g2505) & (g2506) & (!g5765) & (g5766)) + ((!g1195) & (g2503) & (!g2505) & (!g2506) & (!g5765) & (g5766)) + ((!g1195) & (g2503) & (!g2505) & (g2506) & (!g5765) & (g5766)) + ((!g1195) & (g2503) & (!g2505) & (g2506) & (g5765) & (g5766)) + ((!g1195) & (g2503) & (g2505) & (!g2506) & (!g5765) & (g5766)) + ((!g1195) & (g2503) & (g2505) & (!g2506) & (g5765) & (g5766)) + ((!g1195) & (g2503) & (g2505) & (g2506) & (!g5765) & (g5766)) + ((!g1195) & (g2503) & (g2505) & (g2506) & (g5765) & (g5766)) + ((g1195) & (!g2503) & (!g2505) & (!g2506) & (!g5765) & (g5766)) + ((g1195) & (!g2503) & (!g2505) & (g2506) & (!g5765) & (g5766)) + ((g1195) & (!g2503) & (!g2505) & (g2506) & (g5765) & (g5766)) + ((g1195) & (!g2503) & (g2505) & (!g2506) & (!g5765) & (g5766)) + ((g1195) & (!g2503) & (g2505) & (!g2506) & (g5765) & (g5766)) + ((g1195) & (!g2503) & (g2505) & (g2506) & (!g5765) & (g5766)) + ((g1195) & (!g2503) & (g2505) & (g2506) & (g5765) & (g5766)) + ((g1195) & (g2503) & (!g2505) & (!g2506) & (!g5765) & (g5766)) + ((g1195) & (g2503) & (!g2505) & (!g2506) & (g5765) & (g5766)) + ((g1195) & (g2503) & (!g2505) & (g2506) & (!g5765) & (g5766)) + ((g1195) & (g2503) & (!g2505) & (g2506) & (g5765) & (g5766)) + ((g1195) & (g2503) & (g2505) & (!g2506) & (!g5765) & (g5766)) + ((g1195) & (g2503) & (g2505) & (!g2506) & (g5765) & (g5766)) + ((g1195) & (g2503) & (g2505) & (g2506) & (!g5765) & (g5766)) + ((g1195) & (g2503) & (g2505) & (g2506) & (g5765) & (g5766)));
	assign g2735 = (((g1333) & (g2674)));
	assign g2736 = (((!g2734) & (!g2735)));
	assign g2737 = (((!g827) & (!g1360) & (g2733) & (!g2736)) + ((!g827) & (!g1360) & (g2733) & (g2736)) + ((!g827) & (g1360) & (g2733) & (!g2736)) + ((!g827) & (g1360) & (g2733) & (g2736)) + ((g827) & (!g1360) & (!g2733) & (!g2736)) + ((g827) & (!g1360) & (g2733) & (g2736)) + ((g827) & (g1360) & (!g2733) & (g2736)) + ((g827) & (g1360) & (g2733) & (!g2736)));
	assign g2738 = (((!g1173) & (!g1968) & (!g2441) & (!g2442) & (!g5732) & (g5733)) + ((!g1173) & (!g1968) & (!g2441) & (g2442) & (!g5732) & (g5733)) + ((!g1173) & (!g1968) & (g2441) & (!g2442) & (!g5732) & (g5733)) + ((!g1173) & (!g1968) & (g2441) & (g2442) & (!g5732) & (g5733)) + ((!g1173) & (g1968) & (!g2441) & (!g2442) & (!g5732) & (g5733)) + ((!g1173) & (g1968) & (!g2441) & (g2442) & (!g5732) & (g5733)) + ((!g1173) & (g1968) & (!g2441) & (g2442) & (g5732) & (g5733)) + ((!g1173) & (g1968) & (g2441) & (!g2442) & (!g5732) & (g5733)) + ((!g1173) & (g1968) & (g2441) & (!g2442) & (g5732) & (g5733)) + ((!g1173) & (g1968) & (g2441) & (g2442) & (!g5732) & (g5733)) + ((!g1173) & (g1968) & (g2441) & (g2442) & (g5732) & (g5733)) + ((g1173) & (!g1968) & (!g2441) & (!g2442) & (!g5732) & (g5733)) + ((g1173) & (!g1968) & (!g2441) & (g2442) & (!g5732) & (g5733)) + ((g1173) & (!g1968) & (!g2441) & (g2442) & (g5732) & (g5733)) + ((g1173) & (!g1968) & (g2441) & (!g2442) & (!g5732) & (g5733)) + ((g1173) & (!g1968) & (g2441) & (!g2442) & (g5732) & (g5733)) + ((g1173) & (!g1968) & (g2441) & (g2442) & (!g5732) & (g5733)) + ((g1173) & (!g1968) & (g2441) & (g2442) & (g5732) & (g5733)) + ((g1173) & (g1968) & (!g2441) & (!g2442) & (!g5732) & (g5733)) + ((g1173) & (g1968) & (!g2441) & (!g2442) & (g5732) & (g5733)) + ((g1173) & (g1968) & (!g2441) & (g2442) & (!g5732) & (g5733)) + ((g1173) & (g1968) & (!g2441) & (g2442) & (g5732) & (g5733)) + ((g1173) & (g1968) & (g2441) & (!g2442) & (!g5732) & (g5733)) + ((g1173) & (g1968) & (g2441) & (!g2442) & (g5732) & (g5733)) + ((g1173) & (g1968) & (g2441) & (g2442) & (!g5732) & (g5733)) + ((g1173) & (g1968) & (g2441) & (g2442) & (g5732) & (g5733)));
	assign g2739 = (((g1311) & (g2048)));
	assign g2740 = (((!g2738) & (!g2739)));
	assign g2741 = (((!g827) & (!g1362) & (g2099) & (!g2740)) + ((!g827) & (!g1362) & (g2099) & (g2740)) + ((!g827) & (g1362) & (g2099) & (!g2740)) + ((!g827) & (g1362) & (g2099) & (g2740)) + ((g827) & (!g1362) & (!g2099) & (!g2740)) + ((g827) & (!g1362) & (g2099) & (g2740)) + ((g827) & (g1362) & (!g2099) & (g2740)) + ((g827) & (g1362) & (g2099) & (!g2740)));
	assign g8100 = (((!g3499) & (g4971) & (!g2742)) + ((!g3499) & (g4971) & (g2742)) + ((g3499) & (!g4971) & (g2742)) + ((g3499) & (g4971) & (g2742)));
	assign g2743 = (((!g1181) & (!g2462) & (!g2464) & (!g2465) & (!g5744) & (g5745)) + ((!g1181) & (!g2462) & (!g2464) & (g2465) & (!g5744) & (g5745)) + ((!g1181) & (!g2462) & (g2464) & (!g2465) & (!g5744) & (g5745)) + ((!g1181) & (!g2462) & (g2464) & (g2465) & (!g5744) & (g5745)) + ((!g1181) & (g2462) & (!g2464) & (!g2465) & (!g5744) & (g5745)) + ((!g1181) & (g2462) & (!g2464) & (g2465) & (!g5744) & (g5745)) + ((!g1181) & (g2462) & (!g2464) & (g2465) & (g5744) & (g5745)) + ((!g1181) & (g2462) & (g2464) & (!g2465) & (!g5744) & (g5745)) + ((!g1181) & (g2462) & (g2464) & (!g2465) & (g5744) & (g5745)) + ((!g1181) & (g2462) & (g2464) & (g2465) & (!g5744) & (g5745)) + ((!g1181) & (g2462) & (g2464) & (g2465) & (g5744) & (g5745)) + ((g1181) & (!g2462) & (!g2464) & (!g2465) & (!g5744) & (g5745)) + ((g1181) & (!g2462) & (!g2464) & (g2465) & (!g5744) & (g5745)) + ((g1181) & (!g2462) & (!g2464) & (g2465) & (g5744) & (g5745)) + ((g1181) & (!g2462) & (g2464) & (!g2465) & (!g5744) & (g5745)) + ((g1181) & (!g2462) & (g2464) & (!g2465) & (g5744) & (g5745)) + ((g1181) & (!g2462) & (g2464) & (g2465) & (!g5744) & (g5745)) + ((g1181) & (!g2462) & (g2464) & (g2465) & (g5744) & (g5745)) + ((g1181) & (g2462) & (!g2464) & (!g2465) & (!g5744) & (g5745)) + ((g1181) & (g2462) & (!g2464) & (!g2465) & (g5744) & (g5745)) + ((g1181) & (g2462) & (!g2464) & (g2465) & (!g5744) & (g5745)) + ((g1181) & (g2462) & (!g2464) & (g2465) & (g5744) & (g5745)) + ((g1181) & (g2462) & (g2464) & (!g2465) & (!g5744) & (g5745)) + ((g1181) & (g2462) & (g2464) & (!g2465) & (g5744) & (g5745)) + ((g1181) & (g2462) & (g2464) & (g2465) & (!g5744) & (g5745)) + ((g1181) & (g2462) & (g2464) & (g2465) & (g5744) & (g5745)));
	assign g2744 = (((g1319) & (g2661)));
	assign g2745 = (((!g2743) & (!g2744)));
	assign g2746 = (((!g827) & (!g1364) & (g2742) & (!g2745)) + ((!g827) & (!g1364) & (g2742) & (g2745)) + ((!g827) & (g1364) & (g2742) & (!g2745)) + ((!g827) & (g1364) & (g2742) & (g2745)) + ((g827) & (!g1364) & (!g2742) & (!g2745)) + ((g827) & (!g1364) & (g2742) & (g2745)) + ((g827) & (g1364) & (!g2742) & (g2745)) + ((g827) & (g1364) & (g2742) & (!g2745)));
	assign g8101 = (((!g3429) & (g4974) & (!g2747)) + ((!g3429) & (g4974) & (g2747)) + ((g3429) & (!g4974) & (g2747)) + ((g3429) & (g4974) & (g2747)));
	assign g2748 = (((!g1189) & (!g2486) & (!g2488) & (!g2489) & (!g5756) & (g5757)) + ((!g1189) & (!g2486) & (!g2488) & (g2489) & (!g5756) & (g5757)) + ((!g1189) & (!g2486) & (g2488) & (!g2489) & (!g5756) & (g5757)) + ((!g1189) & (!g2486) & (g2488) & (g2489) & (!g5756) & (g5757)) + ((!g1189) & (g2486) & (!g2488) & (!g2489) & (!g5756) & (g5757)) + ((!g1189) & (g2486) & (!g2488) & (g2489) & (!g5756) & (g5757)) + ((!g1189) & (g2486) & (!g2488) & (g2489) & (g5756) & (g5757)) + ((!g1189) & (g2486) & (g2488) & (!g2489) & (!g5756) & (g5757)) + ((!g1189) & (g2486) & (g2488) & (!g2489) & (g5756) & (g5757)) + ((!g1189) & (g2486) & (g2488) & (g2489) & (!g5756) & (g5757)) + ((!g1189) & (g2486) & (g2488) & (g2489) & (g5756) & (g5757)) + ((g1189) & (!g2486) & (!g2488) & (!g2489) & (!g5756) & (g5757)) + ((g1189) & (!g2486) & (!g2488) & (g2489) & (!g5756) & (g5757)) + ((g1189) & (!g2486) & (!g2488) & (g2489) & (g5756) & (g5757)) + ((g1189) & (!g2486) & (g2488) & (!g2489) & (!g5756) & (g5757)) + ((g1189) & (!g2486) & (g2488) & (!g2489) & (g5756) & (g5757)) + ((g1189) & (!g2486) & (g2488) & (g2489) & (!g5756) & (g5757)) + ((g1189) & (!g2486) & (g2488) & (g2489) & (g5756) & (g5757)) + ((g1189) & (g2486) & (!g2488) & (!g2489) & (!g5756) & (g5757)) + ((g1189) & (g2486) & (!g2488) & (!g2489) & (g5756) & (g5757)) + ((g1189) & (g2486) & (!g2488) & (g2489) & (!g5756) & (g5757)) + ((g1189) & (g2486) & (!g2488) & (g2489) & (g5756) & (g5757)) + ((g1189) & (g2486) & (g2488) & (!g2489) & (!g5756) & (g5757)) + ((g1189) & (g2486) & (g2488) & (!g2489) & (g5756) & (g5757)) + ((g1189) & (g2486) & (g2488) & (g2489) & (!g5756) & (g5757)) + ((g1189) & (g2486) & (g2488) & (g2489) & (g5756) & (g5757)));
	assign g2749 = (((g1327) & (g2669)));
	assign g2750 = (((!g2748) & (!g2749)));
	assign g2751 = (((!g827) & (!g1366) & (g2747) & (!g2750)) + ((!g827) & (!g1366) & (g2747) & (g2750)) + ((!g827) & (g1366) & (g2747) & (!g2750)) + ((!g827) & (g1366) & (g2747) & (g2750)) + ((g827) & (!g1366) & (!g2747) & (!g2750)) + ((g827) & (!g1366) & (g2747) & (g2750)) + ((g827) & (g1366) & (!g2747) & (g2750)) + ((g827) & (g1366) & (g2747) & (!g2750)));
	assign g8102 = (((!g2017) & (g4978) & (!g2752)) + ((!g2017) & (g4978) & (g2752)) + ((g2017) & (!g4978) & (g2752)) + ((g2017) & (g4978) & (g2752)));
	assign g2753 = (((!g1197) & (!g2509) & (!g2511) & (!g2512) & (!g5768) & (g5769)) + ((!g1197) & (!g2509) & (!g2511) & (g2512) & (!g5768) & (g5769)) + ((!g1197) & (!g2509) & (g2511) & (!g2512) & (!g5768) & (g5769)) + ((!g1197) & (!g2509) & (g2511) & (g2512) & (!g5768) & (g5769)) + ((!g1197) & (g2509) & (!g2511) & (!g2512) & (!g5768) & (g5769)) + ((!g1197) & (g2509) & (!g2511) & (g2512) & (!g5768) & (g5769)) + ((!g1197) & (g2509) & (!g2511) & (g2512) & (g5768) & (g5769)) + ((!g1197) & (g2509) & (g2511) & (!g2512) & (!g5768) & (g5769)) + ((!g1197) & (g2509) & (g2511) & (!g2512) & (g5768) & (g5769)) + ((!g1197) & (g2509) & (g2511) & (g2512) & (!g5768) & (g5769)) + ((!g1197) & (g2509) & (g2511) & (g2512) & (g5768) & (g5769)) + ((g1197) & (!g2509) & (!g2511) & (!g2512) & (!g5768) & (g5769)) + ((g1197) & (!g2509) & (!g2511) & (g2512) & (!g5768) & (g5769)) + ((g1197) & (!g2509) & (!g2511) & (g2512) & (g5768) & (g5769)) + ((g1197) & (!g2509) & (g2511) & (!g2512) & (!g5768) & (g5769)) + ((g1197) & (!g2509) & (g2511) & (!g2512) & (g5768) & (g5769)) + ((g1197) & (!g2509) & (g2511) & (g2512) & (!g5768) & (g5769)) + ((g1197) & (!g2509) & (g2511) & (g2512) & (g5768) & (g5769)) + ((g1197) & (g2509) & (!g2511) & (!g2512) & (!g5768) & (g5769)) + ((g1197) & (g2509) & (!g2511) & (!g2512) & (g5768) & (g5769)) + ((g1197) & (g2509) & (!g2511) & (g2512) & (!g5768) & (g5769)) + ((g1197) & (g2509) & (!g2511) & (g2512) & (g5768) & (g5769)) + ((g1197) & (g2509) & (g2511) & (!g2512) & (!g5768) & (g5769)) + ((g1197) & (g2509) & (g2511) & (!g2512) & (g5768) & (g5769)) + ((g1197) & (g2509) & (g2511) & (g2512) & (!g5768) & (g5769)) + ((g1197) & (g2509) & (g2511) & (g2512) & (g5768) & (g5769)));
	assign g2754 = (((g1335) & (g2676)));
	assign g2755 = (((!g2753) & (!g2754)));
	assign g2756 = (((!g827) & (!g1368) & (g2752) & (!g2755)) + ((!g827) & (!g1368) & (g2752) & (g2755)) + ((!g827) & (g1368) & (g2752) & (!g2755)) + ((!g827) & (g1368) & (g2752) & (g2755)) + ((g827) & (!g1368) & (!g2752) & (!g2755)) + ((g827) & (!g1368) & (g2752) & (g2755)) + ((g827) & (g1368) & (!g2752) & (g2755)) + ((g827) & (g1368) & (g2752) & (!g2755)));
	assign g2757 = (((!g2646) & (!g2647) & (!g2648) & (g2678) & (g2679)) + ((!g2646) & (!g2647) & (g2648) & (g2678) & (g2679)) + ((!g2646) & (g2647) & (!g2648) & (g2678) & (g2679)) + ((!g2646) & (g2647) & (g2648) & (!g2678) & (g2679)) + ((!g2646) & (g2647) & (g2648) & (g2678) & (!g2679)) + ((!g2646) & (g2647) & (g2648) & (g2678) & (g2679)) + ((g2646) & (!g2647) & (!g2648) & (g2678) & (g2679)) + ((g2646) & (!g2647) & (g2648) & (!g2678) & (g2679)) + ((g2646) & (!g2647) & (g2648) & (g2678) & (!g2679)) + ((g2646) & (!g2647) & (g2648) & (g2678) & (g2679)) + ((g2646) & (g2647) & (!g2648) & (!g2678) & (g2679)) + ((g2646) & (g2647) & (!g2648) & (g2678) & (!g2679)) + ((g2646) & (g2647) & (!g2648) & (g2678) & (g2679)) + ((g2646) & (g2647) & (g2648) & (!g2678) & (g2679)) + ((g2646) & (g2647) & (g2648) & (g2678) & (!g2679)) + ((g2646) & (g2647) & (g2648) & (g2678) & (g2679)));
	assign g8103 = (((!g3429) & (g4981) & (!g2758)) + ((!g3429) & (g4981) & (g2758)) + ((g3429) & (!g4981) & (g2758)) + ((g3429) & (g4981) & (g2758)));
	assign g8104 = (((!g3464) & (g4984) & (!g2759)) + ((!g3464) & (g4984) & (g2759)) + ((g3464) & (!g4984) & (g2759)) + ((g3464) & (g4984) & (g2759)));
	assign g8105 = (((!g3429) & (g4988) & (!g2760)) + ((!g3429) & (g4988) & (g2760)) + ((g3429) & (!g4988) & (g2760)) + ((g3429) & (g4988) & (g2760)));
	assign g8106 = (((!g3499) & (g4991) & (!g2761)) + ((!g3499) & (g4991) & (g2761)) + ((g3499) & (!g4991) & (g2761)) + ((g3499) & (g4991) & (g2761)));
	assign g2762 = (((g830) & (!g1914) & (!g2681) & (!g2757) & (g5692) & (!g5693)) + ((g830) & (!g1914) & (!g2681) & (!g2757) & (g5692) & (g5693)) + ((g830) & (!g1914) & (!g2681) & (g2757) & (g5692) & (!g5693)) + ((g830) & (!g1914) & (!g2681) & (g2757) & (g5692) & (g5693)) + ((g830) & (!g1914) & (g2681) & (!g2757) & (!g5692) & (g5693)) + ((g830) & (!g1914) & (g2681) & (!g2757) & (g5692) & (g5693)) + ((g830) & (!g1914) & (g2681) & (g2757) & (!g5692) & (g5693)) + ((g830) & (!g1914) & (g2681) & (g2757) & (g5692) & (g5693)) + ((g830) & (g1914) & (!g2681) & (!g2757) & (!g5692) & (!g5693)) + ((g830) & (g1914) & (!g2681) & (!g2757) & (!g5692) & (g5693)) + ((g830) & (g1914) & (!g2681) & (g2757) & (g5692) & (!g5693)) + ((g830) & (g1914) & (!g2681) & (g2757) & (g5692) & (g5693)) + ((g830) & (g1914) & (g2681) & (!g2757) & (!g5692) & (!g5693)) + ((g830) & (g1914) & (g2681) & (!g2757) & (!g5692) & (g5693)) + ((g830) & (g1914) & (g2681) & (g2757) & (g5692) & (!g5693)) + ((g830) & (g1914) & (g2681) & (g2757) & (g5692) & (g5693)));
	assign g2763 = (((!g827) & (!g1346) & (!g1376) & (!g2098) & (g2129) & (!g2701)) + ((!g827) & (!g1346) & (!g1376) & (!g2098) & (g2129) & (g2701)) + ((!g827) & (!g1346) & (!g1376) & (g2098) & (g2129) & (!g2701)) + ((!g827) & (!g1346) & (!g1376) & (g2098) & (g2129) & (g2701)) + ((!g827) & (!g1346) & (g1376) & (!g2098) & (g2129) & (!g2701)) + ((!g827) & (!g1346) & (g1376) & (!g2098) & (g2129) & (g2701)) + ((!g827) & (!g1346) & (g1376) & (g2098) & (g2129) & (!g2701)) + ((!g827) & (!g1346) & (g1376) & (g2098) & (g2129) & (g2701)) + ((!g827) & (g1346) & (!g1376) & (!g2098) & (g2129) & (!g2701)) + ((!g827) & (g1346) & (!g1376) & (!g2098) & (g2129) & (g2701)) + ((!g827) & (g1346) & (!g1376) & (g2098) & (g2129) & (!g2701)) + ((!g827) & (g1346) & (!g1376) & (g2098) & (g2129) & (g2701)) + ((!g827) & (g1346) & (g1376) & (!g2098) & (g2129) & (!g2701)) + ((!g827) & (g1346) & (g1376) & (!g2098) & (g2129) & (g2701)) + ((!g827) & (g1346) & (g1376) & (g2098) & (g2129) & (!g2701)) + ((!g827) & (g1346) & (g1376) & (g2098) & (g2129) & (g2701)) + ((g827) & (!g1346) & (!g1376) & (!g2098) & (g2129) & (!g2701)) + ((g827) & (!g1346) & (!g1376) & (!g2098) & (g2129) & (g2701)) + ((g827) & (!g1346) & (!g1376) & (g2098) & (!g2129) & (!g2701)) + ((g827) & (!g1346) & (!g1376) & (g2098) & (g2129) & (g2701)) + ((g827) & (!g1346) & (g1376) & (!g2098) & (!g2129) & (!g2701)) + ((g827) & (!g1346) & (g1376) & (!g2098) & (!g2129) & (g2701)) + ((g827) & (!g1346) & (g1376) & (g2098) & (!g2129) & (g2701)) + ((g827) & (!g1346) & (g1376) & (g2098) & (g2129) & (!g2701)) + ((g827) & (g1346) & (!g1376) & (!g2098) & (!g2129) & (!g2701)) + ((g827) & (g1346) & (!g1376) & (!g2098) & (g2129) & (g2701)) + ((g827) & (g1346) & (!g1376) & (g2098) & (!g2129) & (!g2701)) + ((g827) & (g1346) & (!g1376) & (g2098) & (!g2129) & (g2701)) + ((g827) & (g1346) & (g1376) & (!g2098) & (!g2129) & (g2701)) + ((g827) & (g1346) & (g1376) & (!g2098) & (g2129) & (!g2701)) + ((g827) & (g1346) & (g1376) & (g2098) & (g2129) & (!g2701)) + ((g827) & (g1346) & (g1376) & (g2098) & (g2129) & (g2701)));
	assign g8107 = (((!g3499) & (g4994) & (!g2764)) + ((!g3499) & (g4994) & (g2764)) + ((g3499) & (!g4994) & (g2764)) + ((g3499) & (g4994) & (g2764)));
	assign g2765 = (((!g827) & (!g1354) & (!g1378) & (!g2718) & (g2764) & (!g2721)) + ((!g827) & (!g1354) & (!g1378) & (!g2718) & (g2764) & (g2721)) + ((!g827) & (!g1354) & (!g1378) & (g2718) & (g2764) & (!g2721)) + ((!g827) & (!g1354) & (!g1378) & (g2718) & (g2764) & (g2721)) + ((!g827) & (!g1354) & (g1378) & (!g2718) & (g2764) & (!g2721)) + ((!g827) & (!g1354) & (g1378) & (!g2718) & (g2764) & (g2721)) + ((!g827) & (!g1354) & (g1378) & (g2718) & (g2764) & (!g2721)) + ((!g827) & (!g1354) & (g1378) & (g2718) & (g2764) & (g2721)) + ((!g827) & (g1354) & (!g1378) & (!g2718) & (g2764) & (!g2721)) + ((!g827) & (g1354) & (!g1378) & (!g2718) & (g2764) & (g2721)) + ((!g827) & (g1354) & (!g1378) & (g2718) & (g2764) & (!g2721)) + ((!g827) & (g1354) & (!g1378) & (g2718) & (g2764) & (g2721)) + ((!g827) & (g1354) & (g1378) & (!g2718) & (g2764) & (!g2721)) + ((!g827) & (g1354) & (g1378) & (!g2718) & (g2764) & (g2721)) + ((!g827) & (g1354) & (g1378) & (g2718) & (g2764) & (!g2721)) + ((!g827) & (g1354) & (g1378) & (g2718) & (g2764) & (g2721)) + ((g827) & (!g1354) & (!g1378) & (!g2718) & (g2764) & (!g2721)) + ((g827) & (!g1354) & (!g1378) & (!g2718) & (g2764) & (g2721)) + ((g827) & (!g1354) & (!g1378) & (g2718) & (!g2764) & (!g2721)) + ((g827) & (!g1354) & (!g1378) & (g2718) & (g2764) & (g2721)) + ((g827) & (!g1354) & (g1378) & (!g2718) & (!g2764) & (!g2721)) + ((g827) & (!g1354) & (g1378) & (!g2718) & (!g2764) & (g2721)) + ((g827) & (!g1354) & (g1378) & (g2718) & (!g2764) & (g2721)) + ((g827) & (!g1354) & (g1378) & (g2718) & (g2764) & (!g2721)) + ((g827) & (g1354) & (!g1378) & (!g2718) & (!g2764) & (!g2721)) + ((g827) & (g1354) & (!g1378) & (!g2718) & (g2764) & (g2721)) + ((g827) & (g1354) & (!g1378) & (g2718) & (!g2764) & (!g2721)) + ((g827) & (g1354) & (!g1378) & (g2718) & (!g2764) & (g2721)) + ((g827) & (g1354) & (g1378) & (!g2718) & (!g2764) & (g2721)) + ((g827) & (g1354) & (g1378) & (!g2718) & (g2764) & (!g2721)) + ((g827) & (g1354) & (g1378) & (g2718) & (g2764) & (!g2721)) + ((g827) & (g1354) & (g1378) & (g2718) & (g2764) & (g2721)));
	assign g2766 = (((!g827) & (!g1362) & (!g1380) & (!g2099) & (g2130) & (!g2740)) + ((!g827) & (!g1362) & (!g1380) & (!g2099) & (g2130) & (g2740)) + ((!g827) & (!g1362) & (!g1380) & (g2099) & (g2130) & (!g2740)) + ((!g827) & (!g1362) & (!g1380) & (g2099) & (g2130) & (g2740)) + ((!g827) & (!g1362) & (g1380) & (!g2099) & (g2130) & (!g2740)) + ((!g827) & (!g1362) & (g1380) & (!g2099) & (g2130) & (g2740)) + ((!g827) & (!g1362) & (g1380) & (g2099) & (g2130) & (!g2740)) + ((!g827) & (!g1362) & (g1380) & (g2099) & (g2130) & (g2740)) + ((!g827) & (g1362) & (!g1380) & (!g2099) & (g2130) & (!g2740)) + ((!g827) & (g1362) & (!g1380) & (!g2099) & (g2130) & (g2740)) + ((!g827) & (g1362) & (!g1380) & (g2099) & (g2130) & (!g2740)) + ((!g827) & (g1362) & (!g1380) & (g2099) & (g2130) & (g2740)) + ((!g827) & (g1362) & (g1380) & (!g2099) & (g2130) & (!g2740)) + ((!g827) & (g1362) & (g1380) & (!g2099) & (g2130) & (g2740)) + ((!g827) & (g1362) & (g1380) & (g2099) & (g2130) & (!g2740)) + ((!g827) & (g1362) & (g1380) & (g2099) & (g2130) & (g2740)) + ((g827) & (!g1362) & (!g1380) & (!g2099) & (g2130) & (!g2740)) + ((g827) & (!g1362) & (!g1380) & (!g2099) & (g2130) & (g2740)) + ((g827) & (!g1362) & (!g1380) & (g2099) & (!g2130) & (!g2740)) + ((g827) & (!g1362) & (!g1380) & (g2099) & (g2130) & (g2740)) + ((g827) & (!g1362) & (g1380) & (!g2099) & (!g2130) & (!g2740)) + ((g827) & (!g1362) & (g1380) & (!g2099) & (!g2130) & (g2740)) + ((g827) & (!g1362) & (g1380) & (g2099) & (!g2130) & (g2740)) + ((g827) & (!g1362) & (g1380) & (g2099) & (g2130) & (!g2740)) + ((g827) & (g1362) & (!g1380) & (!g2099) & (!g2130) & (!g2740)) + ((g827) & (g1362) & (!g1380) & (!g2099) & (g2130) & (g2740)) + ((g827) & (g1362) & (!g1380) & (g2099) & (!g2130) & (!g2740)) + ((g827) & (g1362) & (!g1380) & (g2099) & (!g2130) & (g2740)) + ((g827) & (g1362) & (g1380) & (!g2099) & (!g2130) & (g2740)) + ((g827) & (g1362) & (g1380) & (!g2099) & (g2130) & (!g2740)) + ((g827) & (g1362) & (g1380) & (g2099) & (g2130) & (!g2740)) + ((g827) & (g1362) & (g1380) & (g2099) & (g2130) & (g2740)));
	assign g2767 = (((!g827) & (!g1340) & (!g1382) & (!g2100) & (g2133) & (!g2688)) + ((!g827) & (!g1340) & (!g1382) & (!g2100) & (g2133) & (g2688)) + ((!g827) & (!g1340) & (!g1382) & (g2100) & (g2133) & (!g2688)) + ((!g827) & (!g1340) & (!g1382) & (g2100) & (g2133) & (g2688)) + ((!g827) & (!g1340) & (g1382) & (!g2100) & (g2133) & (!g2688)) + ((!g827) & (!g1340) & (g1382) & (!g2100) & (g2133) & (g2688)) + ((!g827) & (!g1340) & (g1382) & (g2100) & (g2133) & (!g2688)) + ((!g827) & (!g1340) & (g1382) & (g2100) & (g2133) & (g2688)) + ((!g827) & (g1340) & (!g1382) & (!g2100) & (g2133) & (!g2688)) + ((!g827) & (g1340) & (!g1382) & (!g2100) & (g2133) & (g2688)) + ((!g827) & (g1340) & (!g1382) & (g2100) & (g2133) & (!g2688)) + ((!g827) & (g1340) & (!g1382) & (g2100) & (g2133) & (g2688)) + ((!g827) & (g1340) & (g1382) & (!g2100) & (g2133) & (!g2688)) + ((!g827) & (g1340) & (g1382) & (!g2100) & (g2133) & (g2688)) + ((!g827) & (g1340) & (g1382) & (g2100) & (g2133) & (!g2688)) + ((!g827) & (g1340) & (g1382) & (g2100) & (g2133) & (g2688)) + ((g827) & (!g1340) & (!g1382) & (!g2100) & (g2133) & (!g2688)) + ((g827) & (!g1340) & (!g1382) & (!g2100) & (g2133) & (g2688)) + ((g827) & (!g1340) & (!g1382) & (g2100) & (!g2133) & (!g2688)) + ((g827) & (!g1340) & (!g1382) & (g2100) & (g2133) & (g2688)) + ((g827) & (!g1340) & (g1382) & (!g2100) & (!g2133) & (!g2688)) + ((g827) & (!g1340) & (g1382) & (!g2100) & (!g2133) & (g2688)) + ((g827) & (!g1340) & (g1382) & (g2100) & (!g2133) & (g2688)) + ((g827) & (!g1340) & (g1382) & (g2100) & (g2133) & (!g2688)) + ((g827) & (g1340) & (!g1382) & (!g2100) & (!g2133) & (!g2688)) + ((g827) & (g1340) & (!g1382) & (!g2100) & (g2133) & (g2688)) + ((g827) & (g1340) & (!g1382) & (g2100) & (!g2133) & (!g2688)) + ((g827) & (g1340) & (!g1382) & (g2100) & (!g2133) & (g2688)) + ((g827) & (g1340) & (g1382) & (!g2100) & (!g2133) & (g2688)) + ((g827) & (g1340) & (g1382) & (!g2100) & (g2133) & (!g2688)) + ((g827) & (g1340) & (g1382) & (g2100) & (g2133) & (!g2688)) + ((g827) & (g1340) & (g1382) & (g2100) & (g2133) & (g2688)));
	assign g8108 = (((!g2017) & (g6266) & (!g2768)) + ((!g2017) & (g6266) & (g2768)) + ((g2017) & (!g6266) & (g2768)) + ((g2017) & (g6266) & (g2768)));
	assign g2769 = (((!g827) & (!g1348) & (!g1384) & (!g2703) & (g2768) & (!g2706)) + ((!g827) & (!g1348) & (!g1384) & (!g2703) & (g2768) & (g2706)) + ((!g827) & (!g1348) & (!g1384) & (g2703) & (g2768) & (!g2706)) + ((!g827) & (!g1348) & (!g1384) & (g2703) & (g2768) & (g2706)) + ((!g827) & (!g1348) & (g1384) & (!g2703) & (g2768) & (!g2706)) + ((!g827) & (!g1348) & (g1384) & (!g2703) & (g2768) & (g2706)) + ((!g827) & (!g1348) & (g1384) & (g2703) & (g2768) & (!g2706)) + ((!g827) & (!g1348) & (g1384) & (g2703) & (g2768) & (g2706)) + ((!g827) & (g1348) & (!g1384) & (!g2703) & (g2768) & (!g2706)) + ((!g827) & (g1348) & (!g1384) & (!g2703) & (g2768) & (g2706)) + ((!g827) & (g1348) & (!g1384) & (g2703) & (g2768) & (!g2706)) + ((!g827) & (g1348) & (!g1384) & (g2703) & (g2768) & (g2706)) + ((!g827) & (g1348) & (g1384) & (!g2703) & (g2768) & (!g2706)) + ((!g827) & (g1348) & (g1384) & (!g2703) & (g2768) & (g2706)) + ((!g827) & (g1348) & (g1384) & (g2703) & (g2768) & (!g2706)) + ((!g827) & (g1348) & (g1384) & (g2703) & (g2768) & (g2706)) + ((g827) & (!g1348) & (!g1384) & (!g2703) & (g2768) & (!g2706)) + ((g827) & (!g1348) & (!g1384) & (!g2703) & (g2768) & (g2706)) + ((g827) & (!g1348) & (!g1384) & (g2703) & (!g2768) & (!g2706)) + ((g827) & (!g1348) & (!g1384) & (g2703) & (g2768) & (g2706)) + ((g827) & (!g1348) & (g1384) & (!g2703) & (!g2768) & (!g2706)) + ((g827) & (!g1348) & (g1384) & (!g2703) & (!g2768) & (g2706)) + ((g827) & (!g1348) & (g1384) & (g2703) & (!g2768) & (g2706)) + ((g827) & (!g1348) & (g1384) & (g2703) & (g2768) & (!g2706)) + ((g827) & (g1348) & (!g1384) & (!g2703) & (!g2768) & (!g2706)) + ((g827) & (g1348) & (!g1384) & (!g2703) & (g2768) & (g2706)) + ((g827) & (g1348) & (!g1384) & (g2703) & (!g2768) & (!g2706)) + ((g827) & (g1348) & (!g1384) & (g2703) & (!g2768) & (g2706)) + ((g827) & (g1348) & (g1384) & (!g2703) & (!g2768) & (g2706)) + ((g827) & (g1348) & (g1384) & (!g2703) & (g2768) & (!g2706)) + ((g827) & (g1348) & (g1384) & (g2703) & (g2768) & (!g2706)) + ((g827) & (g1348) & (g1384) & (g2703) & (g2768) & (g2706)));
	assign g8109 = (((!g3464) & (g5000) & (!g2770)) + ((!g3464) & (g5000) & (g2770)) + ((g3464) & (!g5000) & (g2770)) + ((g3464) & (g5000) & (g2770)));
	assign g2771 = (((!g827) & (!g1356) & (!g1386) & (!g2723) & (g2770) & (!g2726)) + ((!g827) & (!g1356) & (!g1386) & (!g2723) & (g2770) & (g2726)) + ((!g827) & (!g1356) & (!g1386) & (g2723) & (g2770) & (!g2726)) + ((!g827) & (!g1356) & (!g1386) & (g2723) & (g2770) & (g2726)) + ((!g827) & (!g1356) & (g1386) & (!g2723) & (g2770) & (!g2726)) + ((!g827) & (!g1356) & (g1386) & (!g2723) & (g2770) & (g2726)) + ((!g827) & (!g1356) & (g1386) & (g2723) & (g2770) & (!g2726)) + ((!g827) & (!g1356) & (g1386) & (g2723) & (g2770) & (g2726)) + ((!g827) & (g1356) & (!g1386) & (!g2723) & (g2770) & (!g2726)) + ((!g827) & (g1356) & (!g1386) & (!g2723) & (g2770) & (g2726)) + ((!g827) & (g1356) & (!g1386) & (g2723) & (g2770) & (!g2726)) + ((!g827) & (g1356) & (!g1386) & (g2723) & (g2770) & (g2726)) + ((!g827) & (g1356) & (g1386) & (!g2723) & (g2770) & (!g2726)) + ((!g827) & (g1356) & (g1386) & (!g2723) & (g2770) & (g2726)) + ((!g827) & (g1356) & (g1386) & (g2723) & (g2770) & (!g2726)) + ((!g827) & (g1356) & (g1386) & (g2723) & (g2770) & (g2726)) + ((g827) & (!g1356) & (!g1386) & (!g2723) & (g2770) & (!g2726)) + ((g827) & (!g1356) & (!g1386) & (!g2723) & (g2770) & (g2726)) + ((g827) & (!g1356) & (!g1386) & (g2723) & (!g2770) & (!g2726)) + ((g827) & (!g1356) & (!g1386) & (g2723) & (g2770) & (g2726)) + ((g827) & (!g1356) & (g1386) & (!g2723) & (!g2770) & (!g2726)) + ((g827) & (!g1356) & (g1386) & (!g2723) & (!g2770) & (g2726)) + ((g827) & (!g1356) & (g1386) & (g2723) & (!g2770) & (g2726)) + ((g827) & (!g1356) & (g1386) & (g2723) & (g2770) & (!g2726)) + ((g827) & (g1356) & (!g1386) & (!g2723) & (!g2770) & (!g2726)) + ((g827) & (g1356) & (!g1386) & (!g2723) & (g2770) & (g2726)) + ((g827) & (g1356) & (!g1386) & (g2723) & (!g2770) & (!g2726)) + ((g827) & (g1356) & (!g1386) & (g2723) & (!g2770) & (g2726)) + ((g827) & (g1356) & (g1386) & (!g2723) & (!g2770) & (g2726)) + ((g827) & (g1356) & (g1386) & (!g2723) & (g2770) & (!g2726)) + ((g827) & (g1356) & (g1386) & (g2723) & (g2770) & (!g2726)) + ((g827) & (g1356) & (g1386) & (g2723) & (g2770) & (g2726)));
	assign g8110 = (((!g3499) & (g5003) & (!g2772)) + ((!g3499) & (g5003) & (g2772)) + ((g3499) & (!g5003) & (g2772)) + ((g3499) & (g5003) & (g2772)));
	assign g2773 = (((!g827) & (!g1364) & (!g1388) & (!g2742) & (g2772) & (!g2745)) + ((!g827) & (!g1364) & (!g1388) & (!g2742) & (g2772) & (g2745)) + ((!g827) & (!g1364) & (!g1388) & (g2742) & (g2772) & (!g2745)) + ((!g827) & (!g1364) & (!g1388) & (g2742) & (g2772) & (g2745)) + ((!g827) & (!g1364) & (g1388) & (!g2742) & (g2772) & (!g2745)) + ((!g827) & (!g1364) & (g1388) & (!g2742) & (g2772) & (g2745)) + ((!g827) & (!g1364) & (g1388) & (g2742) & (g2772) & (!g2745)) + ((!g827) & (!g1364) & (g1388) & (g2742) & (g2772) & (g2745)) + ((!g827) & (g1364) & (!g1388) & (!g2742) & (g2772) & (!g2745)) + ((!g827) & (g1364) & (!g1388) & (!g2742) & (g2772) & (g2745)) + ((!g827) & (g1364) & (!g1388) & (g2742) & (g2772) & (!g2745)) + ((!g827) & (g1364) & (!g1388) & (g2742) & (g2772) & (g2745)) + ((!g827) & (g1364) & (g1388) & (!g2742) & (g2772) & (!g2745)) + ((!g827) & (g1364) & (g1388) & (!g2742) & (g2772) & (g2745)) + ((!g827) & (g1364) & (g1388) & (g2742) & (g2772) & (!g2745)) + ((!g827) & (g1364) & (g1388) & (g2742) & (g2772) & (g2745)) + ((g827) & (!g1364) & (!g1388) & (!g2742) & (g2772) & (!g2745)) + ((g827) & (!g1364) & (!g1388) & (!g2742) & (g2772) & (g2745)) + ((g827) & (!g1364) & (!g1388) & (g2742) & (!g2772) & (!g2745)) + ((g827) & (!g1364) & (!g1388) & (g2742) & (g2772) & (g2745)) + ((g827) & (!g1364) & (g1388) & (!g2742) & (!g2772) & (!g2745)) + ((g827) & (!g1364) & (g1388) & (!g2742) & (!g2772) & (g2745)) + ((g827) & (!g1364) & (g1388) & (g2742) & (!g2772) & (g2745)) + ((g827) & (!g1364) & (g1388) & (g2742) & (g2772) & (!g2745)) + ((g827) & (g1364) & (!g1388) & (!g2742) & (!g2772) & (!g2745)) + ((g827) & (g1364) & (!g1388) & (!g2742) & (g2772) & (g2745)) + ((g827) & (g1364) & (!g1388) & (g2742) & (!g2772) & (!g2745)) + ((g827) & (g1364) & (!g1388) & (g2742) & (!g2772) & (g2745)) + ((g827) & (g1364) & (g1388) & (!g2742) & (!g2772) & (g2745)) + ((g827) & (g1364) & (g1388) & (!g2742) & (g2772) & (!g2745)) + ((g827) & (g1364) & (g1388) & (g2742) & (g2772) & (!g2745)) + ((g827) & (g1364) & (g1388) & (g2742) & (g2772) & (g2745)));
	assign g8111 = (((!g3464) & (g5006) & (!g2774)) + ((!g3464) & (g5006) & (g2774)) + ((g3464) & (!g5006) & (g2774)) + ((g3464) & (g5006) & (g2774)));
	assign g2775 = (((!g827) & (!g1342) & (!g1390) & (!g2690) & (g2774) & (!g2693)) + ((!g827) & (!g1342) & (!g1390) & (!g2690) & (g2774) & (g2693)) + ((!g827) & (!g1342) & (!g1390) & (g2690) & (g2774) & (!g2693)) + ((!g827) & (!g1342) & (!g1390) & (g2690) & (g2774) & (g2693)) + ((!g827) & (!g1342) & (g1390) & (!g2690) & (g2774) & (!g2693)) + ((!g827) & (!g1342) & (g1390) & (!g2690) & (g2774) & (g2693)) + ((!g827) & (!g1342) & (g1390) & (g2690) & (g2774) & (!g2693)) + ((!g827) & (!g1342) & (g1390) & (g2690) & (g2774) & (g2693)) + ((!g827) & (g1342) & (!g1390) & (!g2690) & (g2774) & (!g2693)) + ((!g827) & (g1342) & (!g1390) & (!g2690) & (g2774) & (g2693)) + ((!g827) & (g1342) & (!g1390) & (g2690) & (g2774) & (!g2693)) + ((!g827) & (g1342) & (!g1390) & (g2690) & (g2774) & (g2693)) + ((!g827) & (g1342) & (g1390) & (!g2690) & (g2774) & (!g2693)) + ((!g827) & (g1342) & (g1390) & (!g2690) & (g2774) & (g2693)) + ((!g827) & (g1342) & (g1390) & (g2690) & (g2774) & (!g2693)) + ((!g827) & (g1342) & (g1390) & (g2690) & (g2774) & (g2693)) + ((g827) & (!g1342) & (!g1390) & (!g2690) & (g2774) & (!g2693)) + ((g827) & (!g1342) & (!g1390) & (!g2690) & (g2774) & (g2693)) + ((g827) & (!g1342) & (!g1390) & (g2690) & (!g2774) & (!g2693)) + ((g827) & (!g1342) & (!g1390) & (g2690) & (g2774) & (g2693)) + ((g827) & (!g1342) & (g1390) & (!g2690) & (!g2774) & (!g2693)) + ((g827) & (!g1342) & (g1390) & (!g2690) & (!g2774) & (g2693)) + ((g827) & (!g1342) & (g1390) & (g2690) & (!g2774) & (g2693)) + ((g827) & (!g1342) & (g1390) & (g2690) & (g2774) & (!g2693)) + ((g827) & (g1342) & (!g1390) & (!g2690) & (!g2774) & (!g2693)) + ((g827) & (g1342) & (!g1390) & (!g2690) & (g2774) & (g2693)) + ((g827) & (g1342) & (!g1390) & (g2690) & (!g2774) & (!g2693)) + ((g827) & (g1342) & (!g1390) & (g2690) & (!g2774) & (g2693)) + ((g827) & (g1342) & (g1390) & (!g2690) & (!g2774) & (g2693)) + ((g827) & (g1342) & (g1390) & (!g2690) & (g2774) & (!g2693)) + ((g827) & (g1342) & (g1390) & (g2690) & (g2774) & (!g2693)) + ((g827) & (g1342) & (g1390) & (g2690) & (g2774) & (g2693)));
	assign g8112 = (((!g3499) & (g5009) & (!g2776)) + ((!g3499) & (g5009) & (g2776)) + ((g3499) & (!g5009) & (g2776)) + ((g3499) & (g5009) & (g2776)));
	assign g2777 = (((!g827) & (!g1350) & (!g1392) & (!g2708) & (g2776) & (!g2711)) + ((!g827) & (!g1350) & (!g1392) & (!g2708) & (g2776) & (g2711)) + ((!g827) & (!g1350) & (!g1392) & (g2708) & (g2776) & (!g2711)) + ((!g827) & (!g1350) & (!g1392) & (g2708) & (g2776) & (g2711)) + ((!g827) & (!g1350) & (g1392) & (!g2708) & (g2776) & (!g2711)) + ((!g827) & (!g1350) & (g1392) & (!g2708) & (g2776) & (g2711)) + ((!g827) & (!g1350) & (g1392) & (g2708) & (g2776) & (!g2711)) + ((!g827) & (!g1350) & (g1392) & (g2708) & (g2776) & (g2711)) + ((!g827) & (g1350) & (!g1392) & (!g2708) & (g2776) & (!g2711)) + ((!g827) & (g1350) & (!g1392) & (!g2708) & (g2776) & (g2711)) + ((!g827) & (g1350) & (!g1392) & (g2708) & (g2776) & (!g2711)) + ((!g827) & (g1350) & (!g1392) & (g2708) & (g2776) & (g2711)) + ((!g827) & (g1350) & (g1392) & (!g2708) & (g2776) & (!g2711)) + ((!g827) & (g1350) & (g1392) & (!g2708) & (g2776) & (g2711)) + ((!g827) & (g1350) & (g1392) & (g2708) & (g2776) & (!g2711)) + ((!g827) & (g1350) & (g1392) & (g2708) & (g2776) & (g2711)) + ((g827) & (!g1350) & (!g1392) & (!g2708) & (g2776) & (!g2711)) + ((g827) & (!g1350) & (!g1392) & (!g2708) & (g2776) & (g2711)) + ((g827) & (!g1350) & (!g1392) & (g2708) & (!g2776) & (!g2711)) + ((g827) & (!g1350) & (!g1392) & (g2708) & (g2776) & (g2711)) + ((g827) & (!g1350) & (g1392) & (!g2708) & (!g2776) & (!g2711)) + ((g827) & (!g1350) & (g1392) & (!g2708) & (!g2776) & (g2711)) + ((g827) & (!g1350) & (g1392) & (g2708) & (!g2776) & (g2711)) + ((g827) & (!g1350) & (g1392) & (g2708) & (g2776) & (!g2711)) + ((g827) & (g1350) & (!g1392) & (!g2708) & (!g2776) & (!g2711)) + ((g827) & (g1350) & (!g1392) & (!g2708) & (g2776) & (g2711)) + ((g827) & (g1350) & (!g1392) & (g2708) & (!g2776) & (!g2711)) + ((g827) & (g1350) & (!g1392) & (g2708) & (!g2776) & (g2711)) + ((g827) & (g1350) & (g1392) & (!g2708) & (!g2776) & (g2711)) + ((g827) & (g1350) & (g1392) & (!g2708) & (g2776) & (!g2711)) + ((g827) & (g1350) & (g1392) & (g2708) & (g2776) & (!g2711)) + ((g827) & (g1350) & (g1392) & (g2708) & (g2776) & (g2711)));
	assign g8113 = (((!g2017) & (g6216) & (!g2778)) + ((!g2017) & (g6216) & (g2778)) + ((g2017) & (!g6216) & (g2778)) + ((g2017) & (g6216) & (g2778)));
	assign g2779 = (((!g827) & (!g1358) & (!g1394) & (!g2728) & (g2778) & (!g2731)) + ((!g827) & (!g1358) & (!g1394) & (!g2728) & (g2778) & (g2731)) + ((!g827) & (!g1358) & (!g1394) & (g2728) & (g2778) & (!g2731)) + ((!g827) & (!g1358) & (!g1394) & (g2728) & (g2778) & (g2731)) + ((!g827) & (!g1358) & (g1394) & (!g2728) & (g2778) & (!g2731)) + ((!g827) & (!g1358) & (g1394) & (!g2728) & (g2778) & (g2731)) + ((!g827) & (!g1358) & (g1394) & (g2728) & (g2778) & (!g2731)) + ((!g827) & (!g1358) & (g1394) & (g2728) & (g2778) & (g2731)) + ((!g827) & (g1358) & (!g1394) & (!g2728) & (g2778) & (!g2731)) + ((!g827) & (g1358) & (!g1394) & (!g2728) & (g2778) & (g2731)) + ((!g827) & (g1358) & (!g1394) & (g2728) & (g2778) & (!g2731)) + ((!g827) & (g1358) & (!g1394) & (g2728) & (g2778) & (g2731)) + ((!g827) & (g1358) & (g1394) & (!g2728) & (g2778) & (!g2731)) + ((!g827) & (g1358) & (g1394) & (!g2728) & (g2778) & (g2731)) + ((!g827) & (g1358) & (g1394) & (g2728) & (g2778) & (!g2731)) + ((!g827) & (g1358) & (g1394) & (g2728) & (g2778) & (g2731)) + ((g827) & (!g1358) & (!g1394) & (!g2728) & (g2778) & (!g2731)) + ((g827) & (!g1358) & (!g1394) & (!g2728) & (g2778) & (g2731)) + ((g827) & (!g1358) & (!g1394) & (g2728) & (!g2778) & (!g2731)) + ((g827) & (!g1358) & (!g1394) & (g2728) & (g2778) & (g2731)) + ((g827) & (!g1358) & (g1394) & (!g2728) & (!g2778) & (!g2731)) + ((g827) & (!g1358) & (g1394) & (!g2728) & (!g2778) & (g2731)) + ((g827) & (!g1358) & (g1394) & (g2728) & (!g2778) & (g2731)) + ((g827) & (!g1358) & (g1394) & (g2728) & (g2778) & (!g2731)) + ((g827) & (g1358) & (!g1394) & (!g2728) & (!g2778) & (!g2731)) + ((g827) & (g1358) & (!g1394) & (!g2728) & (g2778) & (g2731)) + ((g827) & (g1358) & (!g1394) & (g2728) & (!g2778) & (!g2731)) + ((g827) & (g1358) & (!g1394) & (g2728) & (!g2778) & (g2731)) + ((g827) & (g1358) & (g1394) & (!g2728) & (!g2778) & (g2731)) + ((g827) & (g1358) & (g1394) & (!g2728) & (g2778) & (!g2731)) + ((g827) & (g1358) & (g1394) & (g2728) & (g2778) & (!g2731)) + ((g827) & (g1358) & (g1394) & (g2728) & (g2778) & (g2731)));
	assign g8114 = (((!g3429) & (g5014) & (!g2780)) + ((!g3429) & (g5014) & (g2780)) + ((g3429) & (!g5014) & (g2780)) + ((g3429) & (g5014) & (g2780)));
	assign g2781 = (((!g827) & (!g1366) & (!g1396) & (!g2747) & (g2780) & (!g2750)) + ((!g827) & (!g1366) & (!g1396) & (!g2747) & (g2780) & (g2750)) + ((!g827) & (!g1366) & (!g1396) & (g2747) & (g2780) & (!g2750)) + ((!g827) & (!g1366) & (!g1396) & (g2747) & (g2780) & (g2750)) + ((!g827) & (!g1366) & (g1396) & (!g2747) & (g2780) & (!g2750)) + ((!g827) & (!g1366) & (g1396) & (!g2747) & (g2780) & (g2750)) + ((!g827) & (!g1366) & (g1396) & (g2747) & (g2780) & (!g2750)) + ((!g827) & (!g1366) & (g1396) & (g2747) & (g2780) & (g2750)) + ((!g827) & (g1366) & (!g1396) & (!g2747) & (g2780) & (!g2750)) + ((!g827) & (g1366) & (!g1396) & (!g2747) & (g2780) & (g2750)) + ((!g827) & (g1366) & (!g1396) & (g2747) & (g2780) & (!g2750)) + ((!g827) & (g1366) & (!g1396) & (g2747) & (g2780) & (g2750)) + ((!g827) & (g1366) & (g1396) & (!g2747) & (g2780) & (!g2750)) + ((!g827) & (g1366) & (g1396) & (!g2747) & (g2780) & (g2750)) + ((!g827) & (g1366) & (g1396) & (g2747) & (g2780) & (!g2750)) + ((!g827) & (g1366) & (g1396) & (g2747) & (g2780) & (g2750)) + ((g827) & (!g1366) & (!g1396) & (!g2747) & (g2780) & (!g2750)) + ((g827) & (!g1366) & (!g1396) & (!g2747) & (g2780) & (g2750)) + ((g827) & (!g1366) & (!g1396) & (g2747) & (!g2780) & (!g2750)) + ((g827) & (!g1366) & (!g1396) & (g2747) & (g2780) & (g2750)) + ((g827) & (!g1366) & (g1396) & (!g2747) & (!g2780) & (!g2750)) + ((g827) & (!g1366) & (g1396) & (!g2747) & (!g2780) & (g2750)) + ((g827) & (!g1366) & (g1396) & (g2747) & (!g2780) & (g2750)) + ((g827) & (!g1366) & (g1396) & (g2747) & (g2780) & (!g2750)) + ((g827) & (g1366) & (!g1396) & (!g2747) & (!g2780) & (!g2750)) + ((g827) & (g1366) & (!g1396) & (!g2747) & (g2780) & (g2750)) + ((g827) & (g1366) & (!g1396) & (g2747) & (!g2780) & (!g2750)) + ((g827) & (g1366) & (!g1396) & (g2747) & (!g2780) & (g2750)) + ((g827) & (g1366) & (g1396) & (!g2747) & (!g2780) & (g2750)) + ((g827) & (g1366) & (g1396) & (!g2747) & (g2780) & (!g2750)) + ((g827) & (g1366) & (g1396) & (g2747) & (g2780) & (!g2750)) + ((g827) & (g1366) & (g1396) & (g2747) & (g2780) & (g2750)));
	assign g2782 = (((!g827) & (!g1344) & (!g1398) & (!g2101) & (g2134) & (!g2697)) + ((!g827) & (!g1344) & (!g1398) & (!g2101) & (g2134) & (g2697)) + ((!g827) & (!g1344) & (!g1398) & (g2101) & (g2134) & (!g2697)) + ((!g827) & (!g1344) & (!g1398) & (g2101) & (g2134) & (g2697)) + ((!g827) & (!g1344) & (g1398) & (!g2101) & (g2134) & (!g2697)) + ((!g827) & (!g1344) & (g1398) & (!g2101) & (g2134) & (g2697)) + ((!g827) & (!g1344) & (g1398) & (g2101) & (g2134) & (!g2697)) + ((!g827) & (!g1344) & (g1398) & (g2101) & (g2134) & (g2697)) + ((!g827) & (g1344) & (!g1398) & (!g2101) & (g2134) & (!g2697)) + ((!g827) & (g1344) & (!g1398) & (!g2101) & (g2134) & (g2697)) + ((!g827) & (g1344) & (!g1398) & (g2101) & (g2134) & (!g2697)) + ((!g827) & (g1344) & (!g1398) & (g2101) & (g2134) & (g2697)) + ((!g827) & (g1344) & (g1398) & (!g2101) & (g2134) & (!g2697)) + ((!g827) & (g1344) & (g1398) & (!g2101) & (g2134) & (g2697)) + ((!g827) & (g1344) & (g1398) & (g2101) & (g2134) & (!g2697)) + ((!g827) & (g1344) & (g1398) & (g2101) & (g2134) & (g2697)) + ((g827) & (!g1344) & (!g1398) & (!g2101) & (g2134) & (!g2697)) + ((g827) & (!g1344) & (!g1398) & (!g2101) & (g2134) & (g2697)) + ((g827) & (!g1344) & (!g1398) & (g2101) & (!g2134) & (!g2697)) + ((g827) & (!g1344) & (!g1398) & (g2101) & (g2134) & (g2697)) + ((g827) & (!g1344) & (g1398) & (!g2101) & (!g2134) & (!g2697)) + ((g827) & (!g1344) & (g1398) & (!g2101) & (!g2134) & (g2697)) + ((g827) & (!g1344) & (g1398) & (g2101) & (!g2134) & (g2697)) + ((g827) & (!g1344) & (g1398) & (g2101) & (g2134) & (!g2697)) + ((g827) & (g1344) & (!g1398) & (!g2101) & (!g2134) & (!g2697)) + ((g827) & (g1344) & (!g1398) & (!g2101) & (g2134) & (g2697)) + ((g827) & (g1344) & (!g1398) & (g2101) & (!g2134) & (!g2697)) + ((g827) & (g1344) & (!g1398) & (g2101) & (!g2134) & (g2697)) + ((g827) & (g1344) & (g1398) & (!g2101) & (!g2134) & (g2697)) + ((g827) & (g1344) & (g1398) & (!g2101) & (g2134) & (!g2697)) + ((g827) & (g1344) & (g1398) & (g2101) & (g2134) & (!g2697)) + ((g827) & (g1344) & (g1398) & (g2101) & (g2134) & (g2697)));
	assign g8115 = (((!g3464) & (g5017) & (!g2783)) + ((!g3464) & (g5017) & (g2783)) + ((g3464) & (!g5017) & (g2783)) + ((g3464) & (g5017) & (g2783)));
	assign g2784 = (((!g827) & (!g1352) & (!g1400) & (!g2713) & (g2783) & (!g2716)) + ((!g827) & (!g1352) & (!g1400) & (!g2713) & (g2783) & (g2716)) + ((!g827) & (!g1352) & (!g1400) & (g2713) & (g2783) & (!g2716)) + ((!g827) & (!g1352) & (!g1400) & (g2713) & (g2783) & (g2716)) + ((!g827) & (!g1352) & (g1400) & (!g2713) & (g2783) & (!g2716)) + ((!g827) & (!g1352) & (g1400) & (!g2713) & (g2783) & (g2716)) + ((!g827) & (!g1352) & (g1400) & (g2713) & (g2783) & (!g2716)) + ((!g827) & (!g1352) & (g1400) & (g2713) & (g2783) & (g2716)) + ((!g827) & (g1352) & (!g1400) & (!g2713) & (g2783) & (!g2716)) + ((!g827) & (g1352) & (!g1400) & (!g2713) & (g2783) & (g2716)) + ((!g827) & (g1352) & (!g1400) & (g2713) & (g2783) & (!g2716)) + ((!g827) & (g1352) & (!g1400) & (g2713) & (g2783) & (g2716)) + ((!g827) & (g1352) & (g1400) & (!g2713) & (g2783) & (!g2716)) + ((!g827) & (g1352) & (g1400) & (!g2713) & (g2783) & (g2716)) + ((!g827) & (g1352) & (g1400) & (g2713) & (g2783) & (!g2716)) + ((!g827) & (g1352) & (g1400) & (g2713) & (g2783) & (g2716)) + ((g827) & (!g1352) & (!g1400) & (!g2713) & (g2783) & (!g2716)) + ((g827) & (!g1352) & (!g1400) & (!g2713) & (g2783) & (g2716)) + ((g827) & (!g1352) & (!g1400) & (g2713) & (!g2783) & (!g2716)) + ((g827) & (!g1352) & (!g1400) & (g2713) & (g2783) & (g2716)) + ((g827) & (!g1352) & (g1400) & (!g2713) & (!g2783) & (!g2716)) + ((g827) & (!g1352) & (g1400) & (!g2713) & (!g2783) & (g2716)) + ((g827) & (!g1352) & (g1400) & (g2713) & (!g2783) & (g2716)) + ((g827) & (!g1352) & (g1400) & (g2713) & (g2783) & (!g2716)) + ((g827) & (g1352) & (!g1400) & (!g2713) & (!g2783) & (!g2716)) + ((g827) & (g1352) & (!g1400) & (!g2713) & (g2783) & (g2716)) + ((g827) & (g1352) & (!g1400) & (g2713) & (!g2783) & (!g2716)) + ((g827) & (g1352) & (!g1400) & (g2713) & (!g2783) & (g2716)) + ((g827) & (g1352) & (g1400) & (!g2713) & (!g2783) & (g2716)) + ((g827) & (g1352) & (g1400) & (!g2713) & (g2783) & (!g2716)) + ((g827) & (g1352) & (g1400) & (g2713) & (g2783) & (!g2716)) + ((g827) & (g1352) & (g1400) & (g2713) & (g2783) & (g2716)));
	assign g8116 = (((!g3429) & (g5020) & (!g2785)) + ((!g3429) & (g5020) & (g2785)) + ((g3429) & (!g5020) & (g2785)) + ((g3429) & (g5020) & (g2785)));
	assign g2786 = (((!g827) & (!g1360) & (!g1402) & (!g2733) & (g2785) & (!g2736)) + ((!g827) & (!g1360) & (!g1402) & (!g2733) & (g2785) & (g2736)) + ((!g827) & (!g1360) & (!g1402) & (g2733) & (g2785) & (!g2736)) + ((!g827) & (!g1360) & (!g1402) & (g2733) & (g2785) & (g2736)) + ((!g827) & (!g1360) & (g1402) & (!g2733) & (g2785) & (!g2736)) + ((!g827) & (!g1360) & (g1402) & (!g2733) & (g2785) & (g2736)) + ((!g827) & (!g1360) & (g1402) & (g2733) & (g2785) & (!g2736)) + ((!g827) & (!g1360) & (g1402) & (g2733) & (g2785) & (g2736)) + ((!g827) & (g1360) & (!g1402) & (!g2733) & (g2785) & (!g2736)) + ((!g827) & (g1360) & (!g1402) & (!g2733) & (g2785) & (g2736)) + ((!g827) & (g1360) & (!g1402) & (g2733) & (g2785) & (!g2736)) + ((!g827) & (g1360) & (!g1402) & (g2733) & (g2785) & (g2736)) + ((!g827) & (g1360) & (g1402) & (!g2733) & (g2785) & (!g2736)) + ((!g827) & (g1360) & (g1402) & (!g2733) & (g2785) & (g2736)) + ((!g827) & (g1360) & (g1402) & (g2733) & (g2785) & (!g2736)) + ((!g827) & (g1360) & (g1402) & (g2733) & (g2785) & (g2736)) + ((g827) & (!g1360) & (!g1402) & (!g2733) & (g2785) & (!g2736)) + ((g827) & (!g1360) & (!g1402) & (!g2733) & (g2785) & (g2736)) + ((g827) & (!g1360) & (!g1402) & (g2733) & (!g2785) & (!g2736)) + ((g827) & (!g1360) & (!g1402) & (g2733) & (g2785) & (g2736)) + ((g827) & (!g1360) & (g1402) & (!g2733) & (!g2785) & (!g2736)) + ((g827) & (!g1360) & (g1402) & (!g2733) & (!g2785) & (g2736)) + ((g827) & (!g1360) & (g1402) & (g2733) & (!g2785) & (g2736)) + ((g827) & (!g1360) & (g1402) & (g2733) & (g2785) & (!g2736)) + ((g827) & (g1360) & (!g1402) & (!g2733) & (!g2785) & (!g2736)) + ((g827) & (g1360) & (!g1402) & (!g2733) & (g2785) & (g2736)) + ((g827) & (g1360) & (!g1402) & (g2733) & (!g2785) & (!g2736)) + ((g827) & (g1360) & (!g1402) & (g2733) & (!g2785) & (g2736)) + ((g827) & (g1360) & (g1402) & (!g2733) & (!g2785) & (g2736)) + ((g827) & (g1360) & (g1402) & (!g2733) & (g2785) & (!g2736)) + ((g827) & (g1360) & (g1402) & (g2733) & (g2785) & (!g2736)) + ((g827) & (g1360) & (g1402) & (g2733) & (g2785) & (g2736)));
	assign g8117 = (((!g2017) & (g6199) & (!g2787)) + ((!g2017) & (g6199) & (g2787)) + ((g2017) & (!g6199) & (g2787)) + ((g2017) & (g6199) & (g2787)));
	assign g2788 = (((!g827) & (!g1368) & (!g1404) & (!g2752) & (g2787) & (!g2755)) + ((!g827) & (!g1368) & (!g1404) & (!g2752) & (g2787) & (g2755)) + ((!g827) & (!g1368) & (!g1404) & (g2752) & (g2787) & (!g2755)) + ((!g827) & (!g1368) & (!g1404) & (g2752) & (g2787) & (g2755)) + ((!g827) & (!g1368) & (g1404) & (!g2752) & (g2787) & (!g2755)) + ((!g827) & (!g1368) & (g1404) & (!g2752) & (g2787) & (g2755)) + ((!g827) & (!g1368) & (g1404) & (g2752) & (g2787) & (!g2755)) + ((!g827) & (!g1368) & (g1404) & (g2752) & (g2787) & (g2755)) + ((!g827) & (g1368) & (!g1404) & (!g2752) & (g2787) & (!g2755)) + ((!g827) & (g1368) & (!g1404) & (!g2752) & (g2787) & (g2755)) + ((!g827) & (g1368) & (!g1404) & (g2752) & (g2787) & (!g2755)) + ((!g827) & (g1368) & (!g1404) & (g2752) & (g2787) & (g2755)) + ((!g827) & (g1368) & (g1404) & (!g2752) & (g2787) & (!g2755)) + ((!g827) & (g1368) & (g1404) & (!g2752) & (g2787) & (g2755)) + ((!g827) & (g1368) & (g1404) & (g2752) & (g2787) & (!g2755)) + ((!g827) & (g1368) & (g1404) & (g2752) & (g2787) & (g2755)) + ((g827) & (!g1368) & (!g1404) & (!g2752) & (g2787) & (!g2755)) + ((g827) & (!g1368) & (!g1404) & (!g2752) & (g2787) & (g2755)) + ((g827) & (!g1368) & (!g1404) & (g2752) & (!g2787) & (!g2755)) + ((g827) & (!g1368) & (!g1404) & (g2752) & (g2787) & (g2755)) + ((g827) & (!g1368) & (g1404) & (!g2752) & (!g2787) & (!g2755)) + ((g827) & (!g1368) & (g1404) & (!g2752) & (!g2787) & (g2755)) + ((g827) & (!g1368) & (g1404) & (g2752) & (!g2787) & (g2755)) + ((g827) & (!g1368) & (g1404) & (g2752) & (g2787) & (!g2755)) + ((g827) & (g1368) & (!g1404) & (!g2752) & (!g2787) & (!g2755)) + ((g827) & (g1368) & (!g1404) & (!g2752) & (g2787) & (g2755)) + ((g827) & (g1368) & (!g1404) & (g2752) & (!g2787) & (!g2755)) + ((g827) & (g1368) & (!g1404) & (g2752) & (!g2787) & (g2755)) + ((g827) & (g1368) & (g1404) & (!g2752) & (!g2787) & (g2755)) + ((g827) & (g1368) & (g1404) & (!g2752) & (g2787) & (!g2755)) + ((g827) & (g1368) & (g1404) & (g2752) & (g2787) & (!g2755)) + ((g827) & (g1368) & (g1404) & (g2752) & (g2787) & (g2755)));
	assign g8118 = (((!g3429) & (g5027) & (!g2789)) + ((!g3429) & (g5027) & (g2789)) + ((g3429) & (!g5027) & (g2789)) + ((g3429) & (g5027) & (g2789)));
	assign g8119 = (((!g3464) & (g5030) & (!g2790)) + ((!g3464) & (g5030) & (g2790)) + ((g3464) & (!g5030) & (g2790)) + ((g3464) & (g5030) & (g2790)));
	assign g2791 = (((!g2757) & (!g2758) & (!g2759) & (!g2789) & (g2790)) + ((!g2757) & (!g2758) & (!g2759) & (g2789) & (!g2790)) + ((!g2757) & (!g2758) & (g2759) & (!g2789) & (g2790)) + ((!g2757) & (!g2758) & (g2759) & (g2789) & (!g2790)) + ((!g2757) & (g2758) & (!g2759) & (!g2789) & (g2790)) + ((!g2757) & (g2758) & (!g2759) & (g2789) & (!g2790)) + ((!g2757) & (g2758) & (g2759) & (!g2789) & (!g2790)) + ((!g2757) & (g2758) & (g2759) & (g2789) & (g2790)) + ((g2757) & (!g2758) & (!g2759) & (!g2789) & (g2790)) + ((g2757) & (!g2758) & (!g2759) & (g2789) & (!g2790)) + ((g2757) & (!g2758) & (g2759) & (!g2789) & (!g2790)) + ((g2757) & (!g2758) & (g2759) & (g2789) & (g2790)) + ((g2757) & (g2758) & (!g2759) & (!g2789) & (!g2790)) + ((g2757) & (g2758) & (!g2759) & (g2789) & (g2790)) + ((g2757) & (g2758) & (g2759) & (!g2789) & (!g2790)) + ((g2757) & (g2758) & (g2759) & (g2789) & (g2790)));
	assign g2792 = (((!g2681) & (!g2682) & (!g2683) & (!g2684) & (g2760) & (g2761)) + ((!g2681) & (!g2682) & (!g2683) & (g2684) & (g2760) & (g2761)) + ((!g2681) & (!g2682) & (g2683) & (!g2684) & (g2760) & (g2761)) + ((!g2681) & (!g2682) & (g2683) & (g2684) & (!g2760) & (g2761)) + ((!g2681) & (!g2682) & (g2683) & (g2684) & (g2760) & (!g2761)) + ((!g2681) & (!g2682) & (g2683) & (g2684) & (g2760) & (g2761)) + ((!g2681) & (g2682) & (!g2683) & (!g2684) & (g2760) & (g2761)) + ((!g2681) & (g2682) & (!g2683) & (g2684) & (!g2760) & (g2761)) + ((!g2681) & (g2682) & (!g2683) & (g2684) & (g2760) & (!g2761)) + ((!g2681) & (g2682) & (!g2683) & (g2684) & (g2760) & (g2761)) + ((!g2681) & (g2682) & (g2683) & (!g2684) & (!g2760) & (g2761)) + ((!g2681) & (g2682) & (g2683) & (!g2684) & (g2760) & (!g2761)) + ((!g2681) & (g2682) & (g2683) & (!g2684) & (g2760) & (g2761)) + ((!g2681) & (g2682) & (g2683) & (g2684) & (!g2760) & (g2761)) + ((!g2681) & (g2682) & (g2683) & (g2684) & (g2760) & (!g2761)) + ((!g2681) & (g2682) & (g2683) & (g2684) & (g2760) & (g2761)) + ((g2681) & (!g2682) & (!g2683) & (!g2684) & (g2760) & (g2761)) + ((g2681) & (!g2682) & (!g2683) & (g2684) & (!g2760) & (g2761)) + ((g2681) & (!g2682) & (!g2683) & (g2684) & (g2760) & (!g2761)) + ((g2681) & (!g2682) & (!g2683) & (g2684) & (g2760) & (g2761)) + ((g2681) & (!g2682) & (g2683) & (!g2684) & (!g2760) & (g2761)) + ((g2681) & (!g2682) & (g2683) & (!g2684) & (g2760) & (!g2761)) + ((g2681) & (!g2682) & (g2683) & (!g2684) & (g2760) & (g2761)) + ((g2681) & (!g2682) & (g2683) & (g2684) & (!g2760) & (g2761)) + ((g2681) & (!g2682) & (g2683) & (g2684) & (g2760) & (!g2761)) + ((g2681) & (!g2682) & (g2683) & (g2684) & (g2760) & (g2761)) + ((g2681) & (g2682) & (!g2683) & (!g2684) & (g2760) & (g2761)) + ((g2681) & (g2682) & (!g2683) & (g2684) & (!g2760) & (g2761)) + ((g2681) & (g2682) & (!g2683) & (g2684) & (g2760) & (!g2761)) + ((g2681) & (g2682) & (!g2683) & (g2684) & (g2760) & (g2761)) + ((g2681) & (g2682) & (g2683) & (!g2684) & (!g2760) & (g2761)) + ((g2681) & (g2682) & (g2683) & (!g2684) & (g2760) & (!g2761)) + ((g2681) & (g2682) & (g2683) & (!g2684) & (g2760) & (g2761)) + ((g2681) & (g2682) & (g2683) & (g2684) & (!g2760) & (g2761)) + ((g2681) & (g2682) & (g2683) & (g2684) & (g2760) & (!g2761)) + ((g2681) & (g2682) & (g2683) & (g2684) & (g2760) & (g2761)));
	assign g8120 = (((!g3429) & (g5034) & (!g2793)) + ((!g3429) & (g5034) & (g2793)) + ((g3429) & (!g5034) & (g2793)) + ((g3429) & (g5034) & (g2793)));
	assign g8121 = (((!g3499) & (g5037) & (!g2794)) + ((!g3499) & (g5037) & (g2794)) + ((g3499) & (!g5037) & (g2794)) + ((g3499) & (g5037) & (g2794)));
	assign g2795 = (((!g1340) & (!g1382) & (!g2100) & (!g2133) & (!g2686) & (!g2687)) + ((!g1340) & (!g1382) & (!g2100) & (!g2133) & (!g2686) & (g2687)) + ((!g1340) & (!g1382) & (!g2100) & (!g2133) & (g2686) & (!g2687)) + ((!g1340) & (!g1382) & (!g2100) & (!g2133) & (g2686) & (g2687)) + ((!g1340) & (!g1382) & (!g2100) & (g2133) & (!g2686) & (!g2687)) + ((!g1340) & (!g1382) & (!g2100) & (g2133) & (!g2686) & (g2687)) + ((!g1340) & (!g1382) & (!g2100) & (g2133) & (g2686) & (!g2687)) + ((!g1340) & (!g1382) & (!g2100) & (g2133) & (g2686) & (g2687)) + ((!g1340) & (!g1382) & (g2100) & (!g2133) & (!g2686) & (!g2687)) + ((!g1340) & (!g1382) & (g2100) & (!g2133) & (!g2686) & (g2687)) + ((!g1340) & (!g1382) & (g2100) & (!g2133) & (g2686) & (!g2687)) + ((!g1340) & (!g1382) & (g2100) & (!g2133) & (g2686) & (g2687)) + ((!g1340) & (!g1382) & (g2100) & (g2133) & (!g2686) & (!g2687)) + ((!g1340) & (g1382) & (!g2100) & (!g2133) & (!g2686) & (!g2687)) + ((!g1340) & (g1382) & (!g2100) & (!g2133) & (!g2686) & (g2687)) + ((!g1340) & (g1382) & (!g2100) & (!g2133) & (g2686) & (!g2687)) + ((!g1340) & (g1382) & (!g2100) & (!g2133) & (g2686) & (g2687)) + ((!g1340) & (g1382) & (g2100) & (!g2133) & (!g2686) & (!g2687)) + ((g1340) & (!g1382) & (!g2100) & (!g2133) & (!g2686) & (!g2687)) + ((g1340) & (!g1382) & (!g2100) & (!g2133) & (!g2686) & (g2687)) + ((g1340) & (!g1382) & (!g2100) & (!g2133) & (g2686) & (!g2687)) + ((g1340) & (!g1382) & (!g2100) & (!g2133) & (g2686) & (g2687)) + ((g1340) & (!g1382) & (!g2100) & (g2133) & (!g2686) & (!g2687)) + ((g1340) & (!g1382) & (g2100) & (!g2133) & (!g2686) & (!g2687)) + ((g1340) & (!g1382) & (g2100) & (!g2133) & (!g2686) & (g2687)) + ((g1340) & (!g1382) & (g2100) & (!g2133) & (g2686) & (!g2687)) + ((g1340) & (!g1382) & (g2100) & (!g2133) & (g2686) & (g2687)) + ((g1340) & (g1382) & (!g2100) & (!g2133) & (!g2686) & (!g2687)));
	assign g2796 = (((!g827) & (!g1409) & (g2180) & (!g2795)) + ((!g827) & (!g1409) & (g2180) & (g2795)) + ((!g827) & (g1409) & (g2180) & (!g2795)) + ((!g827) & (g1409) & (g2180) & (g2795)) + ((g827) & (!g1409) & (!g2180) & (!g2795)) + ((g827) & (!g1409) & (g2180) & (g2795)) + ((g827) & (g1409) & (!g2180) & (g2795)) + ((g827) & (g1409) & (g2180) & (!g2795)));
	assign g8122 = (((!g3464) & (g5041) & (!g2797)) + ((!g3464) & (g5041) & (g2797)) + ((g3464) & (!g5041) & (g2797)) + ((g3464) & (g5041) & (g2797)));
	assign g2798 = (((!g1342) & (!g1390) & (!g2690) & (!g2774) & (!g2691) & (!g2692)) + ((!g1342) & (!g1390) & (!g2690) & (!g2774) & (!g2691) & (g2692)) + ((!g1342) & (!g1390) & (!g2690) & (!g2774) & (g2691) & (!g2692)) + ((!g1342) & (!g1390) & (!g2690) & (!g2774) & (g2691) & (g2692)) + ((!g1342) & (!g1390) & (!g2690) & (g2774) & (!g2691) & (!g2692)) + ((!g1342) & (!g1390) & (!g2690) & (g2774) & (!g2691) & (g2692)) + ((!g1342) & (!g1390) & (!g2690) & (g2774) & (g2691) & (!g2692)) + ((!g1342) & (!g1390) & (!g2690) & (g2774) & (g2691) & (g2692)) + ((!g1342) & (!g1390) & (g2690) & (!g2774) & (!g2691) & (!g2692)) + ((!g1342) & (!g1390) & (g2690) & (!g2774) & (!g2691) & (g2692)) + ((!g1342) & (!g1390) & (g2690) & (!g2774) & (g2691) & (!g2692)) + ((!g1342) & (!g1390) & (g2690) & (!g2774) & (g2691) & (g2692)) + ((!g1342) & (!g1390) & (g2690) & (g2774) & (!g2691) & (!g2692)) + ((!g1342) & (g1390) & (!g2690) & (!g2774) & (!g2691) & (!g2692)) + ((!g1342) & (g1390) & (!g2690) & (!g2774) & (!g2691) & (g2692)) + ((!g1342) & (g1390) & (!g2690) & (!g2774) & (g2691) & (!g2692)) + ((!g1342) & (g1390) & (!g2690) & (!g2774) & (g2691) & (g2692)) + ((!g1342) & (g1390) & (g2690) & (!g2774) & (!g2691) & (!g2692)) + ((g1342) & (!g1390) & (!g2690) & (!g2774) & (!g2691) & (!g2692)) + ((g1342) & (!g1390) & (!g2690) & (!g2774) & (!g2691) & (g2692)) + ((g1342) & (!g1390) & (!g2690) & (!g2774) & (g2691) & (!g2692)) + ((g1342) & (!g1390) & (!g2690) & (!g2774) & (g2691) & (g2692)) + ((g1342) & (!g1390) & (!g2690) & (g2774) & (!g2691) & (!g2692)) + ((g1342) & (!g1390) & (g2690) & (!g2774) & (!g2691) & (!g2692)) + ((g1342) & (!g1390) & (g2690) & (!g2774) & (!g2691) & (g2692)) + ((g1342) & (!g1390) & (g2690) & (!g2774) & (g2691) & (!g2692)) + ((g1342) & (!g1390) & (g2690) & (!g2774) & (g2691) & (g2692)) + ((g1342) & (g1390) & (!g2690) & (!g2774) & (!g2691) & (!g2692)));
	assign g2799 = (((!g827) & (!g1411) & (g2797) & (!g2798)) + ((!g827) & (!g1411) & (g2797) & (g2798)) + ((!g827) & (g1411) & (g2797) & (!g2798)) + ((!g827) & (g1411) & (g2797) & (g2798)) + ((g827) & (!g1411) & (!g2797) & (!g2798)) + ((g827) & (!g1411) & (g2797) & (g2798)) + ((g827) & (g1411) & (!g2797) & (g2798)) + ((g827) & (g1411) & (g2797) & (!g2798)));
	assign g2800 = (((!g1344) & (!g1398) & (!g2101) & (!g2134) & (!g2695) & (!g2696)) + ((!g1344) & (!g1398) & (!g2101) & (!g2134) & (!g2695) & (g2696)) + ((!g1344) & (!g1398) & (!g2101) & (!g2134) & (g2695) & (!g2696)) + ((!g1344) & (!g1398) & (!g2101) & (!g2134) & (g2695) & (g2696)) + ((!g1344) & (!g1398) & (!g2101) & (g2134) & (!g2695) & (!g2696)) + ((!g1344) & (!g1398) & (!g2101) & (g2134) & (!g2695) & (g2696)) + ((!g1344) & (!g1398) & (!g2101) & (g2134) & (g2695) & (!g2696)) + ((!g1344) & (!g1398) & (!g2101) & (g2134) & (g2695) & (g2696)) + ((!g1344) & (!g1398) & (g2101) & (!g2134) & (!g2695) & (!g2696)) + ((!g1344) & (!g1398) & (g2101) & (!g2134) & (!g2695) & (g2696)) + ((!g1344) & (!g1398) & (g2101) & (!g2134) & (g2695) & (!g2696)) + ((!g1344) & (!g1398) & (g2101) & (!g2134) & (g2695) & (g2696)) + ((!g1344) & (!g1398) & (g2101) & (g2134) & (!g2695) & (!g2696)) + ((!g1344) & (g1398) & (!g2101) & (!g2134) & (!g2695) & (!g2696)) + ((!g1344) & (g1398) & (!g2101) & (!g2134) & (!g2695) & (g2696)) + ((!g1344) & (g1398) & (!g2101) & (!g2134) & (g2695) & (!g2696)) + ((!g1344) & (g1398) & (!g2101) & (!g2134) & (g2695) & (g2696)) + ((!g1344) & (g1398) & (g2101) & (!g2134) & (!g2695) & (!g2696)) + ((g1344) & (!g1398) & (!g2101) & (!g2134) & (!g2695) & (!g2696)) + ((g1344) & (!g1398) & (!g2101) & (!g2134) & (!g2695) & (g2696)) + ((g1344) & (!g1398) & (!g2101) & (!g2134) & (g2695) & (!g2696)) + ((g1344) & (!g1398) & (!g2101) & (!g2134) & (g2695) & (g2696)) + ((g1344) & (!g1398) & (!g2101) & (g2134) & (!g2695) & (!g2696)) + ((g1344) & (!g1398) & (g2101) & (!g2134) & (!g2695) & (!g2696)) + ((g1344) & (!g1398) & (g2101) & (!g2134) & (!g2695) & (g2696)) + ((g1344) & (!g1398) & (g2101) & (!g2134) & (g2695) & (!g2696)) + ((g1344) & (!g1398) & (g2101) & (!g2134) & (g2695) & (g2696)) + ((g1344) & (g1398) & (!g2101) & (!g2134) & (!g2695) & (!g2696)));
	assign g2801 = (((!g827) & (!g1413) & (g2181) & (!g2800)) + ((!g827) & (!g1413) & (g2181) & (g2800)) + ((!g827) & (g1413) & (g2181) & (!g2800)) + ((!g827) & (g1413) & (g2181) & (g2800)) + ((g827) & (!g1413) & (!g2181) & (!g2800)) + ((g827) & (!g1413) & (g2181) & (g2800)) + ((g827) & (g1413) & (!g2181) & (g2800)) + ((g827) & (g1413) & (g2181) & (!g2800)));
	assign g2802 = (((!g1346) & (!g1376) & (!g2098) & (!g2129) & (!g2699) & (!g2700)) + ((!g1346) & (!g1376) & (!g2098) & (!g2129) & (!g2699) & (g2700)) + ((!g1346) & (!g1376) & (!g2098) & (!g2129) & (g2699) & (!g2700)) + ((!g1346) & (!g1376) & (!g2098) & (!g2129) & (g2699) & (g2700)) + ((!g1346) & (!g1376) & (!g2098) & (g2129) & (!g2699) & (!g2700)) + ((!g1346) & (!g1376) & (!g2098) & (g2129) & (!g2699) & (g2700)) + ((!g1346) & (!g1376) & (!g2098) & (g2129) & (g2699) & (!g2700)) + ((!g1346) & (!g1376) & (!g2098) & (g2129) & (g2699) & (g2700)) + ((!g1346) & (!g1376) & (g2098) & (!g2129) & (!g2699) & (!g2700)) + ((!g1346) & (!g1376) & (g2098) & (!g2129) & (!g2699) & (g2700)) + ((!g1346) & (!g1376) & (g2098) & (!g2129) & (g2699) & (!g2700)) + ((!g1346) & (!g1376) & (g2098) & (!g2129) & (g2699) & (g2700)) + ((!g1346) & (!g1376) & (g2098) & (g2129) & (!g2699) & (!g2700)) + ((!g1346) & (g1376) & (!g2098) & (!g2129) & (!g2699) & (!g2700)) + ((!g1346) & (g1376) & (!g2098) & (!g2129) & (!g2699) & (g2700)) + ((!g1346) & (g1376) & (!g2098) & (!g2129) & (g2699) & (!g2700)) + ((!g1346) & (g1376) & (!g2098) & (!g2129) & (g2699) & (g2700)) + ((!g1346) & (g1376) & (g2098) & (!g2129) & (!g2699) & (!g2700)) + ((g1346) & (!g1376) & (!g2098) & (!g2129) & (!g2699) & (!g2700)) + ((g1346) & (!g1376) & (!g2098) & (!g2129) & (!g2699) & (g2700)) + ((g1346) & (!g1376) & (!g2098) & (!g2129) & (g2699) & (!g2700)) + ((g1346) & (!g1376) & (!g2098) & (!g2129) & (g2699) & (g2700)) + ((g1346) & (!g1376) & (!g2098) & (g2129) & (!g2699) & (!g2700)) + ((g1346) & (!g1376) & (g2098) & (!g2129) & (!g2699) & (!g2700)) + ((g1346) & (!g1376) & (g2098) & (!g2129) & (!g2699) & (g2700)) + ((g1346) & (!g1376) & (g2098) & (!g2129) & (g2699) & (!g2700)) + ((g1346) & (!g1376) & (g2098) & (!g2129) & (g2699) & (g2700)) + ((g1346) & (g1376) & (!g2098) & (!g2129) & (!g2699) & (!g2700)));
	assign g2803 = (((!g827) & (!g1415) & (g2177) & (!g2802)) + ((!g827) & (!g1415) & (g2177) & (g2802)) + ((!g827) & (g1415) & (g2177) & (!g2802)) + ((!g827) & (g1415) & (g2177) & (g2802)) + ((g827) & (!g1415) & (!g2177) & (!g2802)) + ((g827) & (!g1415) & (g2177) & (g2802)) + ((g827) & (g1415) & (!g2177) & (g2802)) + ((g827) & (g1415) & (g2177) & (!g2802)));
	assign g8123 = (((!g2017) & (g6193) & (!g2804)) + ((!g2017) & (g6193) & (g2804)) + ((g2017) & (!g6193) & (g2804)) + ((g2017) & (g6193) & (g2804)));
	assign g2805 = (((!g1348) & (!g1384) & (!g2703) & (!g2768) & (!g2704) & (!g2705)) + ((!g1348) & (!g1384) & (!g2703) & (!g2768) & (!g2704) & (g2705)) + ((!g1348) & (!g1384) & (!g2703) & (!g2768) & (g2704) & (!g2705)) + ((!g1348) & (!g1384) & (!g2703) & (!g2768) & (g2704) & (g2705)) + ((!g1348) & (!g1384) & (!g2703) & (g2768) & (!g2704) & (!g2705)) + ((!g1348) & (!g1384) & (!g2703) & (g2768) & (!g2704) & (g2705)) + ((!g1348) & (!g1384) & (!g2703) & (g2768) & (g2704) & (!g2705)) + ((!g1348) & (!g1384) & (!g2703) & (g2768) & (g2704) & (g2705)) + ((!g1348) & (!g1384) & (g2703) & (!g2768) & (!g2704) & (!g2705)) + ((!g1348) & (!g1384) & (g2703) & (!g2768) & (!g2704) & (g2705)) + ((!g1348) & (!g1384) & (g2703) & (!g2768) & (g2704) & (!g2705)) + ((!g1348) & (!g1384) & (g2703) & (!g2768) & (g2704) & (g2705)) + ((!g1348) & (!g1384) & (g2703) & (g2768) & (!g2704) & (!g2705)) + ((!g1348) & (g1384) & (!g2703) & (!g2768) & (!g2704) & (!g2705)) + ((!g1348) & (g1384) & (!g2703) & (!g2768) & (!g2704) & (g2705)) + ((!g1348) & (g1384) & (!g2703) & (!g2768) & (g2704) & (!g2705)) + ((!g1348) & (g1384) & (!g2703) & (!g2768) & (g2704) & (g2705)) + ((!g1348) & (g1384) & (g2703) & (!g2768) & (!g2704) & (!g2705)) + ((g1348) & (!g1384) & (!g2703) & (!g2768) & (!g2704) & (!g2705)) + ((g1348) & (!g1384) & (!g2703) & (!g2768) & (!g2704) & (g2705)) + ((g1348) & (!g1384) & (!g2703) & (!g2768) & (g2704) & (!g2705)) + ((g1348) & (!g1384) & (!g2703) & (!g2768) & (g2704) & (g2705)) + ((g1348) & (!g1384) & (!g2703) & (g2768) & (!g2704) & (!g2705)) + ((g1348) & (!g1384) & (g2703) & (!g2768) & (!g2704) & (!g2705)) + ((g1348) & (!g1384) & (g2703) & (!g2768) & (!g2704) & (g2705)) + ((g1348) & (!g1384) & (g2703) & (!g2768) & (g2704) & (!g2705)) + ((g1348) & (!g1384) & (g2703) & (!g2768) & (g2704) & (g2705)) + ((g1348) & (g1384) & (!g2703) & (!g2768) & (!g2704) & (!g2705)));
	assign g2806 = (((!g827) & (!g1417) & (g2804) & (!g2805)) + ((!g827) & (!g1417) & (g2804) & (g2805)) + ((!g827) & (g1417) & (g2804) & (!g2805)) + ((!g827) & (g1417) & (g2804) & (g2805)) + ((g827) & (!g1417) & (!g2804) & (!g2805)) + ((g827) & (!g1417) & (g2804) & (g2805)) + ((g827) & (g1417) & (!g2804) & (g2805)) + ((g827) & (g1417) & (g2804) & (!g2805)));
	assign g8124 = (((!g3499) & (g5045) & (!g2807)) + ((!g3499) & (g5045) & (g2807)) + ((g3499) & (!g5045) & (g2807)) + ((g3499) & (g5045) & (g2807)));
	assign g2808 = (((!g1350) & (!g1392) & (!g2708) & (!g2776) & (!g2709) & (!g2710)) + ((!g1350) & (!g1392) & (!g2708) & (!g2776) & (!g2709) & (g2710)) + ((!g1350) & (!g1392) & (!g2708) & (!g2776) & (g2709) & (!g2710)) + ((!g1350) & (!g1392) & (!g2708) & (!g2776) & (g2709) & (g2710)) + ((!g1350) & (!g1392) & (!g2708) & (g2776) & (!g2709) & (!g2710)) + ((!g1350) & (!g1392) & (!g2708) & (g2776) & (!g2709) & (g2710)) + ((!g1350) & (!g1392) & (!g2708) & (g2776) & (g2709) & (!g2710)) + ((!g1350) & (!g1392) & (!g2708) & (g2776) & (g2709) & (g2710)) + ((!g1350) & (!g1392) & (g2708) & (!g2776) & (!g2709) & (!g2710)) + ((!g1350) & (!g1392) & (g2708) & (!g2776) & (!g2709) & (g2710)) + ((!g1350) & (!g1392) & (g2708) & (!g2776) & (g2709) & (!g2710)) + ((!g1350) & (!g1392) & (g2708) & (!g2776) & (g2709) & (g2710)) + ((!g1350) & (!g1392) & (g2708) & (g2776) & (!g2709) & (!g2710)) + ((!g1350) & (g1392) & (!g2708) & (!g2776) & (!g2709) & (!g2710)) + ((!g1350) & (g1392) & (!g2708) & (!g2776) & (!g2709) & (g2710)) + ((!g1350) & (g1392) & (!g2708) & (!g2776) & (g2709) & (!g2710)) + ((!g1350) & (g1392) & (!g2708) & (!g2776) & (g2709) & (g2710)) + ((!g1350) & (g1392) & (g2708) & (!g2776) & (!g2709) & (!g2710)) + ((g1350) & (!g1392) & (!g2708) & (!g2776) & (!g2709) & (!g2710)) + ((g1350) & (!g1392) & (!g2708) & (!g2776) & (!g2709) & (g2710)) + ((g1350) & (!g1392) & (!g2708) & (!g2776) & (g2709) & (!g2710)) + ((g1350) & (!g1392) & (!g2708) & (!g2776) & (g2709) & (g2710)) + ((g1350) & (!g1392) & (!g2708) & (g2776) & (!g2709) & (!g2710)) + ((g1350) & (!g1392) & (g2708) & (!g2776) & (!g2709) & (!g2710)) + ((g1350) & (!g1392) & (g2708) & (!g2776) & (!g2709) & (g2710)) + ((g1350) & (!g1392) & (g2708) & (!g2776) & (g2709) & (!g2710)) + ((g1350) & (!g1392) & (g2708) & (!g2776) & (g2709) & (g2710)) + ((g1350) & (g1392) & (!g2708) & (!g2776) & (!g2709) & (!g2710)));
	assign g2809 = (((!g827) & (!g1419) & (g2807) & (!g2808)) + ((!g827) & (!g1419) & (g2807) & (g2808)) + ((!g827) & (g1419) & (g2807) & (!g2808)) + ((!g827) & (g1419) & (g2807) & (g2808)) + ((g827) & (!g1419) & (!g2807) & (!g2808)) + ((g827) & (!g1419) & (g2807) & (g2808)) + ((g827) & (g1419) & (!g2807) & (g2808)) + ((g827) & (g1419) & (g2807) & (!g2808)));
	assign g8125 = (((!g3464) & (g5049) & (!g2810)) + ((!g3464) & (g5049) & (g2810)) + ((g3464) & (!g5049) & (g2810)) + ((g3464) & (g5049) & (g2810)));
	assign g2811 = (((!g1352) & (!g1400) & (!g2713) & (!g2783) & (!g2714) & (!g2715)) + ((!g1352) & (!g1400) & (!g2713) & (!g2783) & (!g2714) & (g2715)) + ((!g1352) & (!g1400) & (!g2713) & (!g2783) & (g2714) & (!g2715)) + ((!g1352) & (!g1400) & (!g2713) & (!g2783) & (g2714) & (g2715)) + ((!g1352) & (!g1400) & (!g2713) & (g2783) & (!g2714) & (!g2715)) + ((!g1352) & (!g1400) & (!g2713) & (g2783) & (!g2714) & (g2715)) + ((!g1352) & (!g1400) & (!g2713) & (g2783) & (g2714) & (!g2715)) + ((!g1352) & (!g1400) & (!g2713) & (g2783) & (g2714) & (g2715)) + ((!g1352) & (!g1400) & (g2713) & (!g2783) & (!g2714) & (!g2715)) + ((!g1352) & (!g1400) & (g2713) & (!g2783) & (!g2714) & (g2715)) + ((!g1352) & (!g1400) & (g2713) & (!g2783) & (g2714) & (!g2715)) + ((!g1352) & (!g1400) & (g2713) & (!g2783) & (g2714) & (g2715)) + ((!g1352) & (!g1400) & (g2713) & (g2783) & (!g2714) & (!g2715)) + ((!g1352) & (g1400) & (!g2713) & (!g2783) & (!g2714) & (!g2715)) + ((!g1352) & (g1400) & (!g2713) & (!g2783) & (!g2714) & (g2715)) + ((!g1352) & (g1400) & (!g2713) & (!g2783) & (g2714) & (!g2715)) + ((!g1352) & (g1400) & (!g2713) & (!g2783) & (g2714) & (g2715)) + ((!g1352) & (g1400) & (g2713) & (!g2783) & (!g2714) & (!g2715)) + ((g1352) & (!g1400) & (!g2713) & (!g2783) & (!g2714) & (!g2715)) + ((g1352) & (!g1400) & (!g2713) & (!g2783) & (!g2714) & (g2715)) + ((g1352) & (!g1400) & (!g2713) & (!g2783) & (g2714) & (!g2715)) + ((g1352) & (!g1400) & (!g2713) & (!g2783) & (g2714) & (g2715)) + ((g1352) & (!g1400) & (!g2713) & (g2783) & (!g2714) & (!g2715)) + ((g1352) & (!g1400) & (g2713) & (!g2783) & (!g2714) & (!g2715)) + ((g1352) & (!g1400) & (g2713) & (!g2783) & (!g2714) & (g2715)) + ((g1352) & (!g1400) & (g2713) & (!g2783) & (g2714) & (!g2715)) + ((g1352) & (!g1400) & (g2713) & (!g2783) & (g2714) & (g2715)) + ((g1352) & (g1400) & (!g2713) & (!g2783) & (!g2714) & (!g2715)));
	assign g2812 = (((!g827) & (!g1421) & (g2810) & (!g2811)) + ((!g827) & (!g1421) & (g2810) & (g2811)) + ((!g827) & (g1421) & (g2810) & (!g2811)) + ((!g827) & (g1421) & (g2810) & (g2811)) + ((g827) & (!g1421) & (!g2810) & (!g2811)) + ((g827) & (!g1421) & (g2810) & (g2811)) + ((g827) & (g1421) & (!g2810) & (g2811)) + ((g827) & (g1421) & (g2810) & (!g2811)));
	assign g8126 = (((!g3499) & (g5053) & (!g2813)) + ((!g3499) & (g5053) & (g2813)) + ((g3499) & (!g5053) & (g2813)) + ((g3499) & (g5053) & (g2813)));
	assign g2814 = (((!g1354) & (!g1378) & (!g2718) & (!g2764) & (!g2719) & (!g2720)) + ((!g1354) & (!g1378) & (!g2718) & (!g2764) & (!g2719) & (g2720)) + ((!g1354) & (!g1378) & (!g2718) & (!g2764) & (g2719) & (!g2720)) + ((!g1354) & (!g1378) & (!g2718) & (!g2764) & (g2719) & (g2720)) + ((!g1354) & (!g1378) & (!g2718) & (g2764) & (!g2719) & (!g2720)) + ((!g1354) & (!g1378) & (!g2718) & (g2764) & (!g2719) & (g2720)) + ((!g1354) & (!g1378) & (!g2718) & (g2764) & (g2719) & (!g2720)) + ((!g1354) & (!g1378) & (!g2718) & (g2764) & (g2719) & (g2720)) + ((!g1354) & (!g1378) & (g2718) & (!g2764) & (!g2719) & (!g2720)) + ((!g1354) & (!g1378) & (g2718) & (!g2764) & (!g2719) & (g2720)) + ((!g1354) & (!g1378) & (g2718) & (!g2764) & (g2719) & (!g2720)) + ((!g1354) & (!g1378) & (g2718) & (!g2764) & (g2719) & (g2720)) + ((!g1354) & (!g1378) & (g2718) & (g2764) & (!g2719) & (!g2720)) + ((!g1354) & (g1378) & (!g2718) & (!g2764) & (!g2719) & (!g2720)) + ((!g1354) & (g1378) & (!g2718) & (!g2764) & (!g2719) & (g2720)) + ((!g1354) & (g1378) & (!g2718) & (!g2764) & (g2719) & (!g2720)) + ((!g1354) & (g1378) & (!g2718) & (!g2764) & (g2719) & (g2720)) + ((!g1354) & (g1378) & (g2718) & (!g2764) & (!g2719) & (!g2720)) + ((g1354) & (!g1378) & (!g2718) & (!g2764) & (!g2719) & (!g2720)) + ((g1354) & (!g1378) & (!g2718) & (!g2764) & (!g2719) & (g2720)) + ((g1354) & (!g1378) & (!g2718) & (!g2764) & (g2719) & (!g2720)) + ((g1354) & (!g1378) & (!g2718) & (!g2764) & (g2719) & (g2720)) + ((g1354) & (!g1378) & (!g2718) & (g2764) & (!g2719) & (!g2720)) + ((g1354) & (!g1378) & (g2718) & (!g2764) & (!g2719) & (!g2720)) + ((g1354) & (!g1378) & (g2718) & (!g2764) & (!g2719) & (g2720)) + ((g1354) & (!g1378) & (g2718) & (!g2764) & (g2719) & (!g2720)) + ((g1354) & (!g1378) & (g2718) & (!g2764) & (g2719) & (g2720)) + ((g1354) & (g1378) & (!g2718) & (!g2764) & (!g2719) & (!g2720)));
	assign g2815 = (((!g827) & (!g1423) & (g2813) & (!g2814)) + ((!g827) & (!g1423) & (g2813) & (g2814)) + ((!g827) & (g1423) & (g2813) & (!g2814)) + ((!g827) & (g1423) & (g2813) & (g2814)) + ((g827) & (!g1423) & (!g2813) & (!g2814)) + ((g827) & (!g1423) & (g2813) & (g2814)) + ((g827) & (g1423) & (!g2813) & (g2814)) + ((g827) & (g1423) & (g2813) & (!g2814)));
	assign g8127 = (((!g3464) & (g5058) & (!g2816)) + ((!g3464) & (g5058) & (g2816)) + ((g3464) & (!g5058) & (g2816)) + ((g3464) & (g5058) & (g2816)));
	assign g2817 = (((!g1356) & (!g1386) & (!g2723) & (!g2770) & (!g2724) & (!g2725)) + ((!g1356) & (!g1386) & (!g2723) & (!g2770) & (!g2724) & (g2725)) + ((!g1356) & (!g1386) & (!g2723) & (!g2770) & (g2724) & (!g2725)) + ((!g1356) & (!g1386) & (!g2723) & (!g2770) & (g2724) & (g2725)) + ((!g1356) & (!g1386) & (!g2723) & (g2770) & (!g2724) & (!g2725)) + ((!g1356) & (!g1386) & (!g2723) & (g2770) & (!g2724) & (g2725)) + ((!g1356) & (!g1386) & (!g2723) & (g2770) & (g2724) & (!g2725)) + ((!g1356) & (!g1386) & (!g2723) & (g2770) & (g2724) & (g2725)) + ((!g1356) & (!g1386) & (g2723) & (!g2770) & (!g2724) & (!g2725)) + ((!g1356) & (!g1386) & (g2723) & (!g2770) & (!g2724) & (g2725)) + ((!g1356) & (!g1386) & (g2723) & (!g2770) & (g2724) & (!g2725)) + ((!g1356) & (!g1386) & (g2723) & (!g2770) & (g2724) & (g2725)) + ((!g1356) & (!g1386) & (g2723) & (g2770) & (!g2724) & (!g2725)) + ((!g1356) & (g1386) & (!g2723) & (!g2770) & (!g2724) & (!g2725)) + ((!g1356) & (g1386) & (!g2723) & (!g2770) & (!g2724) & (g2725)) + ((!g1356) & (g1386) & (!g2723) & (!g2770) & (g2724) & (!g2725)) + ((!g1356) & (g1386) & (!g2723) & (!g2770) & (g2724) & (g2725)) + ((!g1356) & (g1386) & (g2723) & (!g2770) & (!g2724) & (!g2725)) + ((g1356) & (!g1386) & (!g2723) & (!g2770) & (!g2724) & (!g2725)) + ((g1356) & (!g1386) & (!g2723) & (!g2770) & (!g2724) & (g2725)) + ((g1356) & (!g1386) & (!g2723) & (!g2770) & (g2724) & (!g2725)) + ((g1356) & (!g1386) & (!g2723) & (!g2770) & (g2724) & (g2725)) + ((g1356) & (!g1386) & (!g2723) & (g2770) & (!g2724) & (!g2725)) + ((g1356) & (!g1386) & (g2723) & (!g2770) & (!g2724) & (!g2725)) + ((g1356) & (!g1386) & (g2723) & (!g2770) & (!g2724) & (g2725)) + ((g1356) & (!g1386) & (g2723) & (!g2770) & (g2724) & (!g2725)) + ((g1356) & (!g1386) & (g2723) & (!g2770) & (g2724) & (g2725)) + ((g1356) & (g1386) & (!g2723) & (!g2770) & (!g2724) & (!g2725)));
	assign g2818 = (((!g827) & (!g1425) & (g2816) & (!g2817)) + ((!g827) & (!g1425) & (g2816) & (g2817)) + ((!g827) & (g1425) & (g2816) & (!g2817)) + ((!g827) & (g1425) & (g2816) & (g2817)) + ((g827) & (!g1425) & (!g2816) & (!g2817)) + ((g827) & (!g1425) & (g2816) & (g2817)) + ((g827) & (g1425) & (!g2816) & (g2817)) + ((g827) & (g1425) & (g2816) & (!g2817)));
	assign g8128 = (((!g2017) & (g6187) & (!g2819)) + ((!g2017) & (g6187) & (g2819)) + ((g2017) & (!g6187) & (g2819)) + ((g2017) & (g6187) & (g2819)));
	assign g2820 = (((!g1358) & (!g1394) & (!g2728) & (!g2778) & (!g2729) & (!g2730)) + ((!g1358) & (!g1394) & (!g2728) & (!g2778) & (!g2729) & (g2730)) + ((!g1358) & (!g1394) & (!g2728) & (!g2778) & (g2729) & (!g2730)) + ((!g1358) & (!g1394) & (!g2728) & (!g2778) & (g2729) & (g2730)) + ((!g1358) & (!g1394) & (!g2728) & (g2778) & (!g2729) & (!g2730)) + ((!g1358) & (!g1394) & (!g2728) & (g2778) & (!g2729) & (g2730)) + ((!g1358) & (!g1394) & (!g2728) & (g2778) & (g2729) & (!g2730)) + ((!g1358) & (!g1394) & (!g2728) & (g2778) & (g2729) & (g2730)) + ((!g1358) & (!g1394) & (g2728) & (!g2778) & (!g2729) & (!g2730)) + ((!g1358) & (!g1394) & (g2728) & (!g2778) & (!g2729) & (g2730)) + ((!g1358) & (!g1394) & (g2728) & (!g2778) & (g2729) & (!g2730)) + ((!g1358) & (!g1394) & (g2728) & (!g2778) & (g2729) & (g2730)) + ((!g1358) & (!g1394) & (g2728) & (g2778) & (!g2729) & (!g2730)) + ((!g1358) & (g1394) & (!g2728) & (!g2778) & (!g2729) & (!g2730)) + ((!g1358) & (g1394) & (!g2728) & (!g2778) & (!g2729) & (g2730)) + ((!g1358) & (g1394) & (!g2728) & (!g2778) & (g2729) & (!g2730)) + ((!g1358) & (g1394) & (!g2728) & (!g2778) & (g2729) & (g2730)) + ((!g1358) & (g1394) & (g2728) & (!g2778) & (!g2729) & (!g2730)) + ((g1358) & (!g1394) & (!g2728) & (!g2778) & (!g2729) & (!g2730)) + ((g1358) & (!g1394) & (!g2728) & (!g2778) & (!g2729) & (g2730)) + ((g1358) & (!g1394) & (!g2728) & (!g2778) & (g2729) & (!g2730)) + ((g1358) & (!g1394) & (!g2728) & (!g2778) & (g2729) & (g2730)) + ((g1358) & (!g1394) & (!g2728) & (g2778) & (!g2729) & (!g2730)) + ((g1358) & (!g1394) & (g2728) & (!g2778) & (!g2729) & (!g2730)) + ((g1358) & (!g1394) & (g2728) & (!g2778) & (!g2729) & (g2730)) + ((g1358) & (!g1394) & (g2728) & (!g2778) & (g2729) & (!g2730)) + ((g1358) & (!g1394) & (g2728) & (!g2778) & (g2729) & (g2730)) + ((g1358) & (g1394) & (!g2728) & (!g2778) & (!g2729) & (!g2730)));
	assign g2821 = (((!g827) & (!g1427) & (g2819) & (!g2820)) + ((!g827) & (!g1427) & (g2819) & (g2820)) + ((!g827) & (g1427) & (g2819) & (!g2820)) + ((!g827) & (g1427) & (g2819) & (g2820)) + ((g827) & (!g1427) & (!g2819) & (!g2820)) + ((g827) & (!g1427) & (g2819) & (g2820)) + ((g827) & (g1427) & (!g2819) & (g2820)) + ((g827) & (g1427) & (g2819) & (!g2820)));
	assign g8129 = (((!g3429) & (g5063) & (!g2822)) + ((!g3429) & (g5063) & (g2822)) + ((g3429) & (!g5063) & (g2822)) + ((g3429) & (g5063) & (g2822)));
	assign g2823 = (((!g1360) & (!g1402) & (!g2733) & (!g2785) & (!g2734) & (!g2735)) + ((!g1360) & (!g1402) & (!g2733) & (!g2785) & (!g2734) & (g2735)) + ((!g1360) & (!g1402) & (!g2733) & (!g2785) & (g2734) & (!g2735)) + ((!g1360) & (!g1402) & (!g2733) & (!g2785) & (g2734) & (g2735)) + ((!g1360) & (!g1402) & (!g2733) & (g2785) & (!g2734) & (!g2735)) + ((!g1360) & (!g1402) & (!g2733) & (g2785) & (!g2734) & (g2735)) + ((!g1360) & (!g1402) & (!g2733) & (g2785) & (g2734) & (!g2735)) + ((!g1360) & (!g1402) & (!g2733) & (g2785) & (g2734) & (g2735)) + ((!g1360) & (!g1402) & (g2733) & (!g2785) & (!g2734) & (!g2735)) + ((!g1360) & (!g1402) & (g2733) & (!g2785) & (!g2734) & (g2735)) + ((!g1360) & (!g1402) & (g2733) & (!g2785) & (g2734) & (!g2735)) + ((!g1360) & (!g1402) & (g2733) & (!g2785) & (g2734) & (g2735)) + ((!g1360) & (!g1402) & (g2733) & (g2785) & (!g2734) & (!g2735)) + ((!g1360) & (g1402) & (!g2733) & (!g2785) & (!g2734) & (!g2735)) + ((!g1360) & (g1402) & (!g2733) & (!g2785) & (!g2734) & (g2735)) + ((!g1360) & (g1402) & (!g2733) & (!g2785) & (g2734) & (!g2735)) + ((!g1360) & (g1402) & (!g2733) & (!g2785) & (g2734) & (g2735)) + ((!g1360) & (g1402) & (g2733) & (!g2785) & (!g2734) & (!g2735)) + ((g1360) & (!g1402) & (!g2733) & (!g2785) & (!g2734) & (!g2735)) + ((g1360) & (!g1402) & (!g2733) & (!g2785) & (!g2734) & (g2735)) + ((g1360) & (!g1402) & (!g2733) & (!g2785) & (g2734) & (!g2735)) + ((g1360) & (!g1402) & (!g2733) & (!g2785) & (g2734) & (g2735)) + ((g1360) & (!g1402) & (!g2733) & (g2785) & (!g2734) & (!g2735)) + ((g1360) & (!g1402) & (g2733) & (!g2785) & (!g2734) & (!g2735)) + ((g1360) & (!g1402) & (g2733) & (!g2785) & (!g2734) & (g2735)) + ((g1360) & (!g1402) & (g2733) & (!g2785) & (g2734) & (!g2735)) + ((g1360) & (!g1402) & (g2733) & (!g2785) & (g2734) & (g2735)) + ((g1360) & (g1402) & (!g2733) & (!g2785) & (!g2734) & (!g2735)));
	assign g2824 = (((!g827) & (!g1429) & (g2822) & (!g2823)) + ((!g827) & (!g1429) & (g2822) & (g2823)) + ((!g827) & (g1429) & (g2822) & (!g2823)) + ((!g827) & (g1429) & (g2822) & (g2823)) + ((g827) & (!g1429) & (!g2822) & (!g2823)) + ((g827) & (!g1429) & (g2822) & (g2823)) + ((g827) & (g1429) & (!g2822) & (g2823)) + ((g827) & (g1429) & (g2822) & (!g2823)));
	assign g2825 = (((!g1362) & (!g1380) & (!g2099) & (!g2130) & (!g2738) & (!g2739)) + ((!g1362) & (!g1380) & (!g2099) & (!g2130) & (!g2738) & (g2739)) + ((!g1362) & (!g1380) & (!g2099) & (!g2130) & (g2738) & (!g2739)) + ((!g1362) & (!g1380) & (!g2099) & (!g2130) & (g2738) & (g2739)) + ((!g1362) & (!g1380) & (!g2099) & (g2130) & (!g2738) & (!g2739)) + ((!g1362) & (!g1380) & (!g2099) & (g2130) & (!g2738) & (g2739)) + ((!g1362) & (!g1380) & (!g2099) & (g2130) & (g2738) & (!g2739)) + ((!g1362) & (!g1380) & (!g2099) & (g2130) & (g2738) & (g2739)) + ((!g1362) & (!g1380) & (g2099) & (!g2130) & (!g2738) & (!g2739)) + ((!g1362) & (!g1380) & (g2099) & (!g2130) & (!g2738) & (g2739)) + ((!g1362) & (!g1380) & (g2099) & (!g2130) & (g2738) & (!g2739)) + ((!g1362) & (!g1380) & (g2099) & (!g2130) & (g2738) & (g2739)) + ((!g1362) & (!g1380) & (g2099) & (g2130) & (!g2738) & (!g2739)) + ((!g1362) & (g1380) & (!g2099) & (!g2130) & (!g2738) & (!g2739)) + ((!g1362) & (g1380) & (!g2099) & (!g2130) & (!g2738) & (g2739)) + ((!g1362) & (g1380) & (!g2099) & (!g2130) & (g2738) & (!g2739)) + ((!g1362) & (g1380) & (!g2099) & (!g2130) & (g2738) & (g2739)) + ((!g1362) & (g1380) & (g2099) & (!g2130) & (!g2738) & (!g2739)) + ((g1362) & (!g1380) & (!g2099) & (!g2130) & (!g2738) & (!g2739)) + ((g1362) & (!g1380) & (!g2099) & (!g2130) & (!g2738) & (g2739)) + ((g1362) & (!g1380) & (!g2099) & (!g2130) & (g2738) & (!g2739)) + ((g1362) & (!g1380) & (!g2099) & (!g2130) & (g2738) & (g2739)) + ((g1362) & (!g1380) & (!g2099) & (g2130) & (!g2738) & (!g2739)) + ((g1362) & (!g1380) & (g2099) & (!g2130) & (!g2738) & (!g2739)) + ((g1362) & (!g1380) & (g2099) & (!g2130) & (!g2738) & (g2739)) + ((g1362) & (!g1380) & (g2099) & (!g2130) & (g2738) & (!g2739)) + ((g1362) & (!g1380) & (g2099) & (!g2130) & (g2738) & (g2739)) + ((g1362) & (g1380) & (!g2099) & (!g2130) & (!g2738) & (!g2739)));
	assign g2826 = (((!g827) & (!g1431) & (g2178) & (!g2825)) + ((!g827) & (!g1431) & (g2178) & (g2825)) + ((!g827) & (g1431) & (g2178) & (!g2825)) + ((!g827) & (g1431) & (g2178) & (g2825)) + ((g827) & (!g1431) & (!g2178) & (!g2825)) + ((g827) & (!g1431) & (g2178) & (g2825)) + ((g827) & (g1431) & (!g2178) & (g2825)) + ((g827) & (g1431) & (g2178) & (!g2825)));
	assign g8130 = (((!g3499) & (g5067) & (!g2827)) + ((!g3499) & (g5067) & (g2827)) + ((g3499) & (!g5067) & (g2827)) + ((g3499) & (g5067) & (g2827)));
	assign g2828 = (((!g1364) & (!g1388) & (!g2742) & (!g2772) & (!g2743) & (!g2744)) + ((!g1364) & (!g1388) & (!g2742) & (!g2772) & (!g2743) & (g2744)) + ((!g1364) & (!g1388) & (!g2742) & (!g2772) & (g2743) & (!g2744)) + ((!g1364) & (!g1388) & (!g2742) & (!g2772) & (g2743) & (g2744)) + ((!g1364) & (!g1388) & (!g2742) & (g2772) & (!g2743) & (!g2744)) + ((!g1364) & (!g1388) & (!g2742) & (g2772) & (!g2743) & (g2744)) + ((!g1364) & (!g1388) & (!g2742) & (g2772) & (g2743) & (!g2744)) + ((!g1364) & (!g1388) & (!g2742) & (g2772) & (g2743) & (g2744)) + ((!g1364) & (!g1388) & (g2742) & (!g2772) & (!g2743) & (!g2744)) + ((!g1364) & (!g1388) & (g2742) & (!g2772) & (!g2743) & (g2744)) + ((!g1364) & (!g1388) & (g2742) & (!g2772) & (g2743) & (!g2744)) + ((!g1364) & (!g1388) & (g2742) & (!g2772) & (g2743) & (g2744)) + ((!g1364) & (!g1388) & (g2742) & (g2772) & (!g2743) & (!g2744)) + ((!g1364) & (g1388) & (!g2742) & (!g2772) & (!g2743) & (!g2744)) + ((!g1364) & (g1388) & (!g2742) & (!g2772) & (!g2743) & (g2744)) + ((!g1364) & (g1388) & (!g2742) & (!g2772) & (g2743) & (!g2744)) + ((!g1364) & (g1388) & (!g2742) & (!g2772) & (g2743) & (g2744)) + ((!g1364) & (g1388) & (g2742) & (!g2772) & (!g2743) & (!g2744)) + ((g1364) & (!g1388) & (!g2742) & (!g2772) & (!g2743) & (!g2744)) + ((g1364) & (!g1388) & (!g2742) & (!g2772) & (!g2743) & (g2744)) + ((g1364) & (!g1388) & (!g2742) & (!g2772) & (g2743) & (!g2744)) + ((g1364) & (!g1388) & (!g2742) & (!g2772) & (g2743) & (g2744)) + ((g1364) & (!g1388) & (!g2742) & (g2772) & (!g2743) & (!g2744)) + ((g1364) & (!g1388) & (g2742) & (!g2772) & (!g2743) & (!g2744)) + ((g1364) & (!g1388) & (g2742) & (!g2772) & (!g2743) & (g2744)) + ((g1364) & (!g1388) & (g2742) & (!g2772) & (g2743) & (!g2744)) + ((g1364) & (!g1388) & (g2742) & (!g2772) & (g2743) & (g2744)) + ((g1364) & (g1388) & (!g2742) & (!g2772) & (!g2743) & (!g2744)));
	assign g2829 = (((!g827) & (!g1433) & (g2827) & (!g2828)) + ((!g827) & (!g1433) & (g2827) & (g2828)) + ((!g827) & (g1433) & (g2827) & (!g2828)) + ((!g827) & (g1433) & (g2827) & (g2828)) + ((g827) & (!g1433) & (!g2827) & (!g2828)) + ((g827) & (!g1433) & (g2827) & (g2828)) + ((g827) & (g1433) & (!g2827) & (g2828)) + ((g827) & (g1433) & (g2827) & (!g2828)));
	assign g8131 = (((!g3429) & (g5072) & (!g2830)) + ((!g3429) & (g5072) & (g2830)) + ((g3429) & (!g5072) & (g2830)) + ((g3429) & (g5072) & (g2830)));
	assign g2831 = (((!g1366) & (!g1396) & (!g2747) & (!g2780) & (!g2748) & (!g2749)) + ((!g1366) & (!g1396) & (!g2747) & (!g2780) & (!g2748) & (g2749)) + ((!g1366) & (!g1396) & (!g2747) & (!g2780) & (g2748) & (!g2749)) + ((!g1366) & (!g1396) & (!g2747) & (!g2780) & (g2748) & (g2749)) + ((!g1366) & (!g1396) & (!g2747) & (g2780) & (!g2748) & (!g2749)) + ((!g1366) & (!g1396) & (!g2747) & (g2780) & (!g2748) & (g2749)) + ((!g1366) & (!g1396) & (!g2747) & (g2780) & (g2748) & (!g2749)) + ((!g1366) & (!g1396) & (!g2747) & (g2780) & (g2748) & (g2749)) + ((!g1366) & (!g1396) & (g2747) & (!g2780) & (!g2748) & (!g2749)) + ((!g1366) & (!g1396) & (g2747) & (!g2780) & (!g2748) & (g2749)) + ((!g1366) & (!g1396) & (g2747) & (!g2780) & (g2748) & (!g2749)) + ((!g1366) & (!g1396) & (g2747) & (!g2780) & (g2748) & (g2749)) + ((!g1366) & (!g1396) & (g2747) & (g2780) & (!g2748) & (!g2749)) + ((!g1366) & (g1396) & (!g2747) & (!g2780) & (!g2748) & (!g2749)) + ((!g1366) & (g1396) & (!g2747) & (!g2780) & (!g2748) & (g2749)) + ((!g1366) & (g1396) & (!g2747) & (!g2780) & (g2748) & (!g2749)) + ((!g1366) & (g1396) & (!g2747) & (!g2780) & (g2748) & (g2749)) + ((!g1366) & (g1396) & (g2747) & (!g2780) & (!g2748) & (!g2749)) + ((g1366) & (!g1396) & (!g2747) & (!g2780) & (!g2748) & (!g2749)) + ((g1366) & (!g1396) & (!g2747) & (!g2780) & (!g2748) & (g2749)) + ((g1366) & (!g1396) & (!g2747) & (!g2780) & (g2748) & (!g2749)) + ((g1366) & (!g1396) & (!g2747) & (!g2780) & (g2748) & (g2749)) + ((g1366) & (!g1396) & (!g2747) & (g2780) & (!g2748) & (!g2749)) + ((g1366) & (!g1396) & (g2747) & (!g2780) & (!g2748) & (!g2749)) + ((g1366) & (!g1396) & (g2747) & (!g2780) & (!g2748) & (g2749)) + ((g1366) & (!g1396) & (g2747) & (!g2780) & (g2748) & (!g2749)) + ((g1366) & (!g1396) & (g2747) & (!g2780) & (g2748) & (g2749)) + ((g1366) & (g1396) & (!g2747) & (!g2780) & (!g2748) & (!g2749)));
	assign g2832 = (((!g827) & (!g1435) & (g2830) & (!g2831)) + ((!g827) & (!g1435) & (g2830) & (g2831)) + ((!g827) & (g1435) & (g2830) & (!g2831)) + ((!g827) & (g1435) & (g2830) & (g2831)) + ((g827) & (!g1435) & (!g2830) & (!g2831)) + ((g827) & (!g1435) & (g2830) & (g2831)) + ((g827) & (g1435) & (!g2830) & (g2831)) + ((g827) & (g1435) & (g2830) & (!g2831)));
	assign g8132 = (((!g2017) & (g6181) & (!g2833)) + ((!g2017) & (g6181) & (g2833)) + ((g2017) & (!g6181) & (g2833)) + ((g2017) & (g6181) & (g2833)));
	assign g2834 = (((!g1368) & (!g1404) & (!g2752) & (!g2787) & (!g2753) & (!g2754)) + ((!g1368) & (!g1404) & (!g2752) & (!g2787) & (!g2753) & (g2754)) + ((!g1368) & (!g1404) & (!g2752) & (!g2787) & (g2753) & (!g2754)) + ((!g1368) & (!g1404) & (!g2752) & (!g2787) & (g2753) & (g2754)) + ((!g1368) & (!g1404) & (!g2752) & (g2787) & (!g2753) & (!g2754)) + ((!g1368) & (!g1404) & (!g2752) & (g2787) & (!g2753) & (g2754)) + ((!g1368) & (!g1404) & (!g2752) & (g2787) & (g2753) & (!g2754)) + ((!g1368) & (!g1404) & (!g2752) & (g2787) & (g2753) & (g2754)) + ((!g1368) & (!g1404) & (g2752) & (!g2787) & (!g2753) & (!g2754)) + ((!g1368) & (!g1404) & (g2752) & (!g2787) & (!g2753) & (g2754)) + ((!g1368) & (!g1404) & (g2752) & (!g2787) & (g2753) & (!g2754)) + ((!g1368) & (!g1404) & (g2752) & (!g2787) & (g2753) & (g2754)) + ((!g1368) & (!g1404) & (g2752) & (g2787) & (!g2753) & (!g2754)) + ((!g1368) & (g1404) & (!g2752) & (!g2787) & (!g2753) & (!g2754)) + ((!g1368) & (g1404) & (!g2752) & (!g2787) & (!g2753) & (g2754)) + ((!g1368) & (g1404) & (!g2752) & (!g2787) & (g2753) & (!g2754)) + ((!g1368) & (g1404) & (!g2752) & (!g2787) & (g2753) & (g2754)) + ((!g1368) & (g1404) & (g2752) & (!g2787) & (!g2753) & (!g2754)) + ((g1368) & (!g1404) & (!g2752) & (!g2787) & (!g2753) & (!g2754)) + ((g1368) & (!g1404) & (!g2752) & (!g2787) & (!g2753) & (g2754)) + ((g1368) & (!g1404) & (!g2752) & (!g2787) & (g2753) & (!g2754)) + ((g1368) & (!g1404) & (!g2752) & (!g2787) & (g2753) & (g2754)) + ((g1368) & (!g1404) & (!g2752) & (g2787) & (!g2753) & (!g2754)) + ((g1368) & (!g1404) & (g2752) & (!g2787) & (!g2753) & (!g2754)) + ((g1368) & (!g1404) & (g2752) & (!g2787) & (!g2753) & (g2754)) + ((g1368) & (!g1404) & (g2752) & (!g2787) & (g2753) & (!g2754)) + ((g1368) & (!g1404) & (g2752) & (!g2787) & (g2753) & (g2754)) + ((g1368) & (g1404) & (!g2752) & (!g2787) & (!g2753) & (!g2754)));
	assign g2835 = (((!g827) & (!g1437) & (g2833) & (!g2834)) + ((!g827) & (!g1437) & (g2833) & (g2834)) + ((!g827) & (g1437) & (g2833) & (!g2834)) + ((!g827) & (g1437) & (g2833) & (g2834)) + ((g827) & (!g1437) & (!g2833) & (!g2834)) + ((g827) & (!g1437) & (g2833) & (g2834)) + ((g827) & (g1437) & (!g2833) & (g2834)) + ((g827) & (g1437) & (g2833) & (!g2834)));
	assign g2836 = (((!g1415) & (g2177) & (!g2802)) + ((g1415) & (!g2177) & (!g2802)) + ((g1415) & (g2177) & (!g2802)) + ((g1415) & (g2177) & (g2802)));
	assign g2837 = (((!g827) & (!g1443) & (g2210) & (!g2836)) + ((!g827) & (!g1443) & (g2210) & (g2836)) + ((!g827) & (g1443) & (g2210) & (!g2836)) + ((!g827) & (g1443) & (g2210) & (g2836)) + ((g827) & (!g1443) & (!g2210) & (g2836)) + ((g827) & (!g1443) & (g2210) & (!g2836)) + ((g827) & (g1443) & (!g2210) & (!g2836)) + ((g827) & (g1443) & (g2210) & (g2836)));
	assign g8133 = (((!g3499) & (g5076) & (!g2838)) + ((!g3499) & (g5076) & (g2838)) + ((g3499) & (!g5076) & (g2838)) + ((g3499) & (g5076) & (g2838)));
	assign g2839 = (((!g1423) & (g2813) & (!g2814)) + ((g1423) & (!g2813) & (!g2814)) + ((g1423) & (g2813) & (!g2814)) + ((g1423) & (g2813) & (g2814)));
	assign g2840 = (((!g827) & (!g1445) & (g2838) & (!g2839)) + ((!g827) & (!g1445) & (g2838) & (g2839)) + ((!g827) & (g1445) & (g2838) & (!g2839)) + ((!g827) & (g1445) & (g2838) & (g2839)) + ((g827) & (!g1445) & (!g2838) & (g2839)) + ((g827) & (!g1445) & (g2838) & (!g2839)) + ((g827) & (g1445) & (!g2838) & (!g2839)) + ((g827) & (g1445) & (g2838) & (g2839)));
	assign g2841 = (((!g1431) & (g2178) & (!g2825)) + ((g1431) & (!g2178) & (!g2825)) + ((g1431) & (g2178) & (!g2825)) + ((g1431) & (g2178) & (g2825)));
	assign g2842 = (((!g827) & (!g1447) & (g2211) & (!g2841)) + ((!g827) & (!g1447) & (g2211) & (g2841)) + ((!g827) & (g1447) & (g2211) & (!g2841)) + ((!g827) & (g1447) & (g2211) & (g2841)) + ((g827) & (!g1447) & (!g2211) & (g2841)) + ((g827) & (!g1447) & (g2211) & (!g2841)) + ((g827) & (g1447) & (!g2211) & (!g2841)) + ((g827) & (g1447) & (g2211) & (g2841)));
	assign g2843 = (((!g1409) & (g2180) & (!g2795)) + ((g1409) & (!g2180) & (!g2795)) + ((g1409) & (g2180) & (!g2795)) + ((g1409) & (g2180) & (g2795)));
	assign g2844 = (((!g827) & (!g1449) & (g2212) & (!g2843)) + ((!g827) & (!g1449) & (g2212) & (g2843)) + ((!g827) & (g1449) & (g2212) & (!g2843)) + ((!g827) & (g1449) & (g2212) & (g2843)) + ((g827) & (!g1449) & (!g2212) & (g2843)) + ((g827) & (!g1449) & (g2212) & (!g2843)) + ((g827) & (g1449) & (!g2212) & (!g2843)) + ((g827) & (g1449) & (g2212) & (g2843)));
	assign g8134 = (((!g2017) & (g5079) & (!g2845)) + ((!g2017) & (g5079) & (g2845)) + ((g2017) & (!g5079) & (g2845)) + ((g2017) & (g5079) & (g2845)));
	assign g2846 = (((!g1417) & (g2804) & (!g2805)) + ((g1417) & (!g2804) & (!g2805)) + ((g1417) & (g2804) & (!g2805)) + ((g1417) & (g2804) & (g2805)));
	assign g2847 = (((!g827) & (!g1451) & (g2845) & (!g2846)) + ((!g827) & (!g1451) & (g2845) & (g2846)) + ((!g827) & (g1451) & (g2845) & (!g2846)) + ((!g827) & (g1451) & (g2845) & (g2846)) + ((g827) & (!g1451) & (!g2845) & (g2846)) + ((g827) & (!g1451) & (g2845) & (!g2846)) + ((g827) & (g1451) & (!g2845) & (!g2846)) + ((g827) & (g1451) & (g2845) & (g2846)));
	assign g8135 = (((!g3464) & (g5084) & (!g2848)) + ((!g3464) & (g5084) & (g2848)) + ((g3464) & (!g5084) & (g2848)) + ((g3464) & (g5084) & (g2848)));
	assign g2849 = (((!g1425) & (g2816) & (!g2817)) + ((g1425) & (!g2816) & (!g2817)) + ((g1425) & (g2816) & (!g2817)) + ((g1425) & (g2816) & (g2817)));
	assign g2850 = (((!g827) & (!g1453) & (g2848) & (!g2849)) + ((!g827) & (!g1453) & (g2848) & (g2849)) + ((!g827) & (g1453) & (g2848) & (!g2849)) + ((!g827) & (g1453) & (g2848) & (g2849)) + ((g827) & (!g1453) & (!g2848) & (g2849)) + ((g827) & (!g1453) & (g2848) & (!g2849)) + ((g827) & (g1453) & (!g2848) & (!g2849)) + ((g827) & (g1453) & (g2848) & (g2849)));
	assign g8136 = (((!g3499) & (g5088) & (!g2851)) + ((!g3499) & (g5088) & (g2851)) + ((g3499) & (!g5088) & (g2851)) + ((g3499) & (g5088) & (g2851)));
	assign g2852 = (((!g1433) & (g2827) & (!g2828)) + ((g1433) & (!g2827) & (!g2828)) + ((g1433) & (g2827) & (!g2828)) + ((g1433) & (g2827) & (g2828)));
	assign g2853 = (((!g827) & (!g1455) & (g2851) & (!g2852)) + ((!g827) & (!g1455) & (g2851) & (g2852)) + ((!g827) & (g1455) & (g2851) & (!g2852)) + ((!g827) & (g1455) & (g2851) & (g2852)) + ((g827) & (!g1455) & (!g2851) & (g2852)) + ((g827) & (!g1455) & (g2851) & (!g2852)) + ((g827) & (g1455) & (!g2851) & (!g2852)) + ((g827) & (g1455) & (g2851) & (g2852)));
	assign g8137 = (((!g3464) & (g5092) & (!g2854)) + ((!g3464) & (g5092) & (g2854)) + ((g3464) & (!g5092) & (g2854)) + ((g3464) & (g5092) & (g2854)));
	assign g2855 = (((!g1411) & (g2797) & (!g2798)) + ((g1411) & (!g2797) & (!g2798)) + ((g1411) & (g2797) & (!g2798)) + ((g1411) & (g2797) & (g2798)));
	assign g2856 = (((!g827) & (!g1457) & (g2854) & (!g2855)) + ((!g827) & (!g1457) & (g2854) & (g2855)) + ((!g827) & (g1457) & (g2854) & (!g2855)) + ((!g827) & (g1457) & (g2854) & (g2855)) + ((g827) & (!g1457) & (!g2854) & (g2855)) + ((g827) & (!g1457) & (g2854) & (!g2855)) + ((g827) & (g1457) & (!g2854) & (!g2855)) + ((g827) & (g1457) & (g2854) & (g2855)));
	assign g8138 = (((!g3499) & (g5096) & (!g2857)) + ((!g3499) & (g5096) & (g2857)) + ((g3499) & (!g5096) & (g2857)) + ((g3499) & (g5096) & (g2857)));
	assign g2858 = (((!g1419) & (g2807) & (!g2808)) + ((g1419) & (!g2807) & (!g2808)) + ((g1419) & (g2807) & (!g2808)) + ((g1419) & (g2807) & (g2808)));
	assign g2859 = (((!g827) & (!g1459) & (g2857) & (!g2858)) + ((!g827) & (!g1459) & (g2857) & (g2858)) + ((!g827) & (g1459) & (g2857) & (!g2858)) + ((!g827) & (g1459) & (g2857) & (g2858)) + ((g827) & (!g1459) & (!g2857) & (g2858)) + ((g827) & (!g1459) & (g2857) & (!g2858)) + ((g827) & (g1459) & (!g2857) & (!g2858)) + ((g827) & (g1459) & (g2857) & (g2858)));
	assign g8139 = (((!g2017) & (g5099) & (!g2860)) + ((!g2017) & (g5099) & (g2860)) + ((g2017) & (!g5099) & (g2860)) + ((g2017) & (g5099) & (g2860)));
	assign g2861 = (((!g1427) & (g2819) & (!g2820)) + ((g1427) & (!g2819) & (!g2820)) + ((g1427) & (g2819) & (!g2820)) + ((g1427) & (g2819) & (g2820)));
	assign g2862 = (((!g827) & (!g1461) & (g2860) & (!g2861)) + ((!g827) & (!g1461) & (g2860) & (g2861)) + ((!g827) & (g1461) & (g2860) & (!g2861)) + ((!g827) & (g1461) & (g2860) & (g2861)) + ((g827) & (!g1461) & (!g2860) & (g2861)) + ((g827) & (!g1461) & (g2860) & (!g2861)) + ((g827) & (g1461) & (!g2860) & (!g2861)) + ((g827) & (g1461) & (g2860) & (g2861)));
	assign g8140 = (((!g3429) & (g5102) & (!g2863)) + ((!g3429) & (g5102) & (g2863)) + ((g3429) & (!g5102) & (g2863)) + ((g3429) & (g5102) & (g2863)));
	assign g2864 = (((!g1435) & (g2830) & (!g2831)) + ((g1435) & (!g2830) & (!g2831)) + ((g1435) & (g2830) & (!g2831)) + ((g1435) & (g2830) & (g2831)));
	assign g2865 = (((!g827) & (!g1463) & (g2863) & (!g2864)) + ((!g827) & (!g1463) & (g2863) & (g2864)) + ((!g827) & (g1463) & (g2863) & (!g2864)) + ((!g827) & (g1463) & (g2863) & (g2864)) + ((g827) & (!g1463) & (!g2863) & (g2864)) + ((g827) & (!g1463) & (g2863) & (!g2864)) + ((g827) & (g1463) & (!g2863) & (!g2864)) + ((g827) & (g1463) & (g2863) & (g2864)));
	assign g2866 = (((!g1413) & (g2181) & (!g2800)) + ((g1413) & (!g2181) & (!g2800)) + ((g1413) & (g2181) & (!g2800)) + ((g1413) & (g2181) & (g2800)));
	assign g2867 = (((!g827) & (!g1465) & (g2213) & (!g2866)) + ((!g827) & (!g1465) & (g2213) & (g2866)) + ((!g827) & (g1465) & (g2213) & (!g2866)) + ((!g827) & (g1465) & (g2213) & (g2866)) + ((g827) & (!g1465) & (!g2213) & (g2866)) + ((g827) & (!g1465) & (g2213) & (!g2866)) + ((g827) & (g1465) & (!g2213) & (!g2866)) + ((g827) & (g1465) & (g2213) & (g2866)));
	assign g8141 = (((!g3464) & (g5106) & (!g2868)) + ((!g3464) & (g5106) & (g2868)) + ((g3464) & (!g5106) & (g2868)) + ((g3464) & (g5106) & (g2868)));
	assign g2869 = (((!g1421) & (g2810) & (!g2811)) + ((g1421) & (!g2810) & (!g2811)) + ((g1421) & (g2810) & (!g2811)) + ((g1421) & (g2810) & (g2811)));
	assign g2870 = (((!g827) & (!g1467) & (g2868) & (!g2869)) + ((!g827) & (!g1467) & (g2868) & (g2869)) + ((!g827) & (g1467) & (g2868) & (!g2869)) + ((!g827) & (g1467) & (g2868) & (g2869)) + ((g827) & (!g1467) & (!g2868) & (g2869)) + ((g827) & (!g1467) & (g2868) & (!g2869)) + ((g827) & (g1467) & (!g2868) & (!g2869)) + ((g827) & (g1467) & (g2868) & (g2869)));
	assign g8142 = (((!g3429) & (g5109) & (!g2871)) + ((!g3429) & (g5109) & (g2871)) + ((g3429) & (!g5109) & (g2871)) + ((g3429) & (g5109) & (g2871)));
	assign g2872 = (((!g1429) & (g2822) & (!g2823)) + ((g1429) & (!g2822) & (!g2823)) + ((g1429) & (g2822) & (!g2823)) + ((g1429) & (g2822) & (g2823)));
	assign g2873 = (((!g827) & (!g1469) & (g2871) & (!g2872)) + ((!g827) & (!g1469) & (g2871) & (g2872)) + ((!g827) & (g1469) & (g2871) & (!g2872)) + ((!g827) & (g1469) & (g2871) & (g2872)) + ((g827) & (!g1469) & (!g2871) & (g2872)) + ((g827) & (!g1469) & (g2871) & (!g2872)) + ((g827) & (g1469) & (!g2871) & (!g2872)) + ((g827) & (g1469) & (g2871) & (g2872)));
	assign g8143 = (((!g2017) & (g5112) & (!g2874)) + ((!g2017) & (g5112) & (g2874)) + ((g2017) & (!g5112) & (g2874)) + ((g2017) & (g5112) & (g2874)));
	assign g2875 = (((!g1437) & (g2833) & (!g2834)) + ((g1437) & (!g2833) & (!g2834)) + ((g1437) & (g2833) & (!g2834)) + ((g1437) & (g2833) & (g2834)));
	assign g2876 = (((!g827) & (!g1471) & (g2874) & (!g2875)) + ((!g827) & (!g1471) & (g2874) & (g2875)) + ((!g827) & (g1471) & (g2874) & (!g2875)) + ((!g827) & (g1471) & (g2874) & (g2875)) + ((g827) & (!g1471) & (!g2874) & (g2875)) + ((g827) & (!g1471) & (g2874) & (!g2875)) + ((g827) & (g1471) & (!g2874) & (!g2875)) + ((g827) & (g1471) & (g2874) & (g2875)));
	assign g2877 = (((!g1890) & (!g1906) & (!g1939) & (g1940)) + ((!g1890) & (!g1906) & (g1939) & (!g1940)) + ((!g1890) & (g1906) & (!g1939) & (g1940)) + ((!g1890) & (g1906) & (g1939) & (!g1940)) + ((g1890) & (!g1906) & (!g1939) & (g1940)) + ((g1890) & (!g1906) & (g1939) & (!g1940)) + ((g1890) & (g1906) & (!g1939) & (!g1940)) + ((g1890) & (g1906) & (g1939) & (g1940)));
	assign g2878 = (((!g1884) & (!g1888) & (!g1977) & (g1978)) + ((!g1884) & (!g1888) & (g1977) & (!g1978)) + ((!g1884) & (g1888) & (!g1977) & (g1978)) + ((!g1884) & (g1888) & (g1977) & (!g1978)) + ((g1884) & (!g1888) & (!g1977) & (g1978)) + ((g1884) & (!g1888) & (g1977) & (!g1978)) + ((g1884) & (g1888) & (!g1977) & (!g1978)) + ((g1884) & (g1888) & (g1977) & (g1978)));
	assign g2879 = (((g830) & (!g1914) & (!g2877) & (!g2878) & (g1473)) + ((g830) & (!g1914) & (!g2877) & (g2878) & (!g1473)) + ((g830) & (!g1914) & (g2877) & (!g2878) & (g1473)) + ((g830) & (!g1914) & (g2877) & (g2878) & (!g1473)) + ((g830) & (g1914) & (!g2877) & (!g2878) & (g1473)) + ((g830) & (g1914) & (!g2877) & (g2878) & (g1473)) + ((g830) & (g1914) & (g2877) & (!g2878) & (!g1473)) + ((g830) & (g1914) & (g2877) & (g2878) & (!g1473)));
	assign g2880 = (((!g827) & (!g1449) & (!g1477) & (!g2212) & (g2262) & (!g2843)) + ((!g827) & (!g1449) & (!g1477) & (!g2212) & (g2262) & (g2843)) + ((!g827) & (!g1449) & (!g1477) & (g2212) & (g2262) & (!g2843)) + ((!g827) & (!g1449) & (!g1477) & (g2212) & (g2262) & (g2843)) + ((!g827) & (!g1449) & (g1477) & (!g2212) & (g2262) & (!g2843)) + ((!g827) & (!g1449) & (g1477) & (!g2212) & (g2262) & (g2843)) + ((!g827) & (!g1449) & (g1477) & (g2212) & (g2262) & (!g2843)) + ((!g827) & (!g1449) & (g1477) & (g2212) & (g2262) & (g2843)) + ((!g827) & (g1449) & (!g1477) & (!g2212) & (g2262) & (!g2843)) + ((!g827) & (g1449) & (!g1477) & (!g2212) & (g2262) & (g2843)) + ((!g827) & (g1449) & (!g1477) & (g2212) & (g2262) & (!g2843)) + ((!g827) & (g1449) & (!g1477) & (g2212) & (g2262) & (g2843)) + ((!g827) & (g1449) & (g1477) & (!g2212) & (g2262) & (!g2843)) + ((!g827) & (g1449) & (g1477) & (!g2212) & (g2262) & (g2843)) + ((!g827) & (g1449) & (g1477) & (g2212) & (g2262) & (!g2843)) + ((!g827) & (g1449) & (g1477) & (g2212) & (g2262) & (g2843)) + ((g827) & (!g1449) & (!g1477) & (!g2212) & (g2262) & (!g2843)) + ((g827) & (!g1449) & (!g1477) & (!g2212) & (g2262) & (g2843)) + ((g827) & (!g1449) & (!g1477) & (g2212) & (!g2262) & (g2843)) + ((g827) & (!g1449) & (!g1477) & (g2212) & (g2262) & (!g2843)) + ((g827) & (!g1449) & (g1477) & (!g2212) & (!g2262) & (!g2843)) + ((g827) & (!g1449) & (g1477) & (!g2212) & (!g2262) & (g2843)) + ((g827) & (!g1449) & (g1477) & (g2212) & (!g2262) & (!g2843)) + ((g827) & (!g1449) & (g1477) & (g2212) & (g2262) & (g2843)) + ((g827) & (g1449) & (!g1477) & (!g2212) & (!g2262) & (g2843)) + ((g827) & (g1449) & (!g1477) & (!g2212) & (g2262) & (!g2843)) + ((g827) & (g1449) & (!g1477) & (g2212) & (!g2262) & (!g2843)) + ((g827) & (g1449) & (!g1477) & (g2212) & (!g2262) & (g2843)) + ((g827) & (g1449) & (g1477) & (!g2212) & (!g2262) & (!g2843)) + ((g827) & (g1449) & (g1477) & (!g2212) & (g2262) & (g2843)) + ((g827) & (g1449) & (g1477) & (g2212) & (g2262) & (!g2843)) + ((g827) & (g1449) & (g1477) & (g2212) & (g2262) & (g2843)));
	assign g8144 = (((!g3464) & (g5115) & (!g2881)) + ((!g3464) & (g5115) & (g2881)) + ((g3464) & (!g5115) & (g2881)) + ((g3464) & (g5115) & (g2881)));
	assign g2882 = (((!g827) & (!g1457) & (!g1479) & (!g2854) & (g2881) & (!g2855)) + ((!g827) & (!g1457) & (!g1479) & (!g2854) & (g2881) & (g2855)) + ((!g827) & (!g1457) & (!g1479) & (g2854) & (g2881) & (!g2855)) + ((!g827) & (!g1457) & (!g1479) & (g2854) & (g2881) & (g2855)) + ((!g827) & (!g1457) & (g1479) & (!g2854) & (g2881) & (!g2855)) + ((!g827) & (!g1457) & (g1479) & (!g2854) & (g2881) & (g2855)) + ((!g827) & (!g1457) & (g1479) & (g2854) & (g2881) & (!g2855)) + ((!g827) & (!g1457) & (g1479) & (g2854) & (g2881) & (g2855)) + ((!g827) & (g1457) & (!g1479) & (!g2854) & (g2881) & (!g2855)) + ((!g827) & (g1457) & (!g1479) & (!g2854) & (g2881) & (g2855)) + ((!g827) & (g1457) & (!g1479) & (g2854) & (g2881) & (!g2855)) + ((!g827) & (g1457) & (!g1479) & (g2854) & (g2881) & (g2855)) + ((!g827) & (g1457) & (g1479) & (!g2854) & (g2881) & (!g2855)) + ((!g827) & (g1457) & (g1479) & (!g2854) & (g2881) & (g2855)) + ((!g827) & (g1457) & (g1479) & (g2854) & (g2881) & (!g2855)) + ((!g827) & (g1457) & (g1479) & (g2854) & (g2881) & (g2855)) + ((g827) & (!g1457) & (!g1479) & (!g2854) & (g2881) & (!g2855)) + ((g827) & (!g1457) & (!g1479) & (!g2854) & (g2881) & (g2855)) + ((g827) & (!g1457) & (!g1479) & (g2854) & (!g2881) & (g2855)) + ((g827) & (!g1457) & (!g1479) & (g2854) & (g2881) & (!g2855)) + ((g827) & (!g1457) & (g1479) & (!g2854) & (!g2881) & (!g2855)) + ((g827) & (!g1457) & (g1479) & (!g2854) & (!g2881) & (g2855)) + ((g827) & (!g1457) & (g1479) & (g2854) & (!g2881) & (!g2855)) + ((g827) & (!g1457) & (g1479) & (g2854) & (g2881) & (g2855)) + ((g827) & (g1457) & (!g1479) & (!g2854) & (!g2881) & (g2855)) + ((g827) & (g1457) & (!g1479) & (!g2854) & (g2881) & (!g2855)) + ((g827) & (g1457) & (!g1479) & (g2854) & (!g2881) & (!g2855)) + ((g827) & (g1457) & (!g1479) & (g2854) & (!g2881) & (g2855)) + ((g827) & (g1457) & (g1479) & (!g2854) & (!g2881) & (!g2855)) + ((g827) & (g1457) & (g1479) & (!g2854) & (g2881) & (g2855)) + ((g827) & (g1457) & (g1479) & (g2854) & (g2881) & (!g2855)) + ((g827) & (g1457) & (g1479) & (g2854) & (g2881) & (g2855)));
	assign g2883 = (((!g827) & (!g1465) & (!g1481) & (!g2213) & (g2263) & (!g2866)) + ((!g827) & (!g1465) & (!g1481) & (!g2213) & (g2263) & (g2866)) + ((!g827) & (!g1465) & (!g1481) & (g2213) & (g2263) & (!g2866)) + ((!g827) & (!g1465) & (!g1481) & (g2213) & (g2263) & (g2866)) + ((!g827) & (!g1465) & (g1481) & (!g2213) & (g2263) & (!g2866)) + ((!g827) & (!g1465) & (g1481) & (!g2213) & (g2263) & (g2866)) + ((!g827) & (!g1465) & (g1481) & (g2213) & (g2263) & (!g2866)) + ((!g827) & (!g1465) & (g1481) & (g2213) & (g2263) & (g2866)) + ((!g827) & (g1465) & (!g1481) & (!g2213) & (g2263) & (!g2866)) + ((!g827) & (g1465) & (!g1481) & (!g2213) & (g2263) & (g2866)) + ((!g827) & (g1465) & (!g1481) & (g2213) & (g2263) & (!g2866)) + ((!g827) & (g1465) & (!g1481) & (g2213) & (g2263) & (g2866)) + ((!g827) & (g1465) & (g1481) & (!g2213) & (g2263) & (!g2866)) + ((!g827) & (g1465) & (g1481) & (!g2213) & (g2263) & (g2866)) + ((!g827) & (g1465) & (g1481) & (g2213) & (g2263) & (!g2866)) + ((!g827) & (g1465) & (g1481) & (g2213) & (g2263) & (g2866)) + ((g827) & (!g1465) & (!g1481) & (!g2213) & (g2263) & (!g2866)) + ((g827) & (!g1465) & (!g1481) & (!g2213) & (g2263) & (g2866)) + ((g827) & (!g1465) & (!g1481) & (g2213) & (!g2263) & (g2866)) + ((g827) & (!g1465) & (!g1481) & (g2213) & (g2263) & (!g2866)) + ((g827) & (!g1465) & (g1481) & (!g2213) & (!g2263) & (!g2866)) + ((g827) & (!g1465) & (g1481) & (!g2213) & (!g2263) & (g2866)) + ((g827) & (!g1465) & (g1481) & (g2213) & (!g2263) & (!g2866)) + ((g827) & (!g1465) & (g1481) & (g2213) & (g2263) & (g2866)) + ((g827) & (g1465) & (!g1481) & (!g2213) & (!g2263) & (g2866)) + ((g827) & (g1465) & (!g1481) & (!g2213) & (g2263) & (!g2866)) + ((g827) & (g1465) & (!g1481) & (g2213) & (!g2263) & (!g2866)) + ((g827) & (g1465) & (!g1481) & (g2213) & (!g2263) & (g2866)) + ((g827) & (g1465) & (g1481) & (!g2213) & (!g2263) & (!g2866)) + ((g827) & (g1465) & (g1481) & (!g2213) & (g2263) & (g2866)) + ((g827) & (g1465) & (g1481) & (g2213) & (g2263) & (!g2866)) + ((g827) & (g1465) & (g1481) & (g2213) & (g2263) & (g2866)));
	assign g2884 = (((!g827) & (!g1443) & (!g1483) & (!g2210) & (g2256) & (!g2836)) + ((!g827) & (!g1443) & (!g1483) & (!g2210) & (g2256) & (g2836)) + ((!g827) & (!g1443) & (!g1483) & (g2210) & (g2256) & (!g2836)) + ((!g827) & (!g1443) & (!g1483) & (g2210) & (g2256) & (g2836)) + ((!g827) & (!g1443) & (g1483) & (!g2210) & (g2256) & (!g2836)) + ((!g827) & (!g1443) & (g1483) & (!g2210) & (g2256) & (g2836)) + ((!g827) & (!g1443) & (g1483) & (g2210) & (g2256) & (!g2836)) + ((!g827) & (!g1443) & (g1483) & (g2210) & (g2256) & (g2836)) + ((!g827) & (g1443) & (!g1483) & (!g2210) & (g2256) & (!g2836)) + ((!g827) & (g1443) & (!g1483) & (!g2210) & (g2256) & (g2836)) + ((!g827) & (g1443) & (!g1483) & (g2210) & (g2256) & (!g2836)) + ((!g827) & (g1443) & (!g1483) & (g2210) & (g2256) & (g2836)) + ((!g827) & (g1443) & (g1483) & (!g2210) & (g2256) & (!g2836)) + ((!g827) & (g1443) & (g1483) & (!g2210) & (g2256) & (g2836)) + ((!g827) & (g1443) & (g1483) & (g2210) & (g2256) & (!g2836)) + ((!g827) & (g1443) & (g1483) & (g2210) & (g2256) & (g2836)) + ((g827) & (!g1443) & (!g1483) & (!g2210) & (g2256) & (!g2836)) + ((g827) & (!g1443) & (!g1483) & (!g2210) & (g2256) & (g2836)) + ((g827) & (!g1443) & (!g1483) & (g2210) & (!g2256) & (g2836)) + ((g827) & (!g1443) & (!g1483) & (g2210) & (g2256) & (!g2836)) + ((g827) & (!g1443) & (g1483) & (!g2210) & (!g2256) & (!g2836)) + ((g827) & (!g1443) & (g1483) & (!g2210) & (!g2256) & (g2836)) + ((g827) & (!g1443) & (g1483) & (g2210) & (!g2256) & (!g2836)) + ((g827) & (!g1443) & (g1483) & (g2210) & (g2256) & (g2836)) + ((g827) & (g1443) & (!g1483) & (!g2210) & (!g2256) & (g2836)) + ((g827) & (g1443) & (!g1483) & (!g2210) & (g2256) & (!g2836)) + ((g827) & (g1443) & (!g1483) & (g2210) & (!g2256) & (!g2836)) + ((g827) & (g1443) & (!g1483) & (g2210) & (!g2256) & (g2836)) + ((g827) & (g1443) & (g1483) & (!g2210) & (!g2256) & (!g2836)) + ((g827) & (g1443) & (g1483) & (!g2210) & (g2256) & (g2836)) + ((g827) & (g1443) & (g1483) & (g2210) & (g2256) & (!g2836)) + ((g827) & (g1443) & (g1483) & (g2210) & (g2256) & (g2836)));
	assign g8145 = (((!g2017) & (g5120) & (!g2885)) + ((!g2017) & (g5120) & (g2885)) + ((g2017) & (!g5120) & (g2885)) + ((g2017) & (g5120) & (g2885)));
	assign g2886 = (((!g827) & (!g1451) & (!g1485) & (!g2845) & (g2885) & (!g2846)) + ((!g827) & (!g1451) & (!g1485) & (!g2845) & (g2885) & (g2846)) + ((!g827) & (!g1451) & (!g1485) & (g2845) & (g2885) & (!g2846)) + ((!g827) & (!g1451) & (!g1485) & (g2845) & (g2885) & (g2846)) + ((!g827) & (!g1451) & (g1485) & (!g2845) & (g2885) & (!g2846)) + ((!g827) & (!g1451) & (g1485) & (!g2845) & (g2885) & (g2846)) + ((!g827) & (!g1451) & (g1485) & (g2845) & (g2885) & (!g2846)) + ((!g827) & (!g1451) & (g1485) & (g2845) & (g2885) & (g2846)) + ((!g827) & (g1451) & (!g1485) & (!g2845) & (g2885) & (!g2846)) + ((!g827) & (g1451) & (!g1485) & (!g2845) & (g2885) & (g2846)) + ((!g827) & (g1451) & (!g1485) & (g2845) & (g2885) & (!g2846)) + ((!g827) & (g1451) & (!g1485) & (g2845) & (g2885) & (g2846)) + ((!g827) & (g1451) & (g1485) & (!g2845) & (g2885) & (!g2846)) + ((!g827) & (g1451) & (g1485) & (!g2845) & (g2885) & (g2846)) + ((!g827) & (g1451) & (g1485) & (g2845) & (g2885) & (!g2846)) + ((!g827) & (g1451) & (g1485) & (g2845) & (g2885) & (g2846)) + ((g827) & (!g1451) & (!g1485) & (!g2845) & (g2885) & (!g2846)) + ((g827) & (!g1451) & (!g1485) & (!g2845) & (g2885) & (g2846)) + ((g827) & (!g1451) & (!g1485) & (g2845) & (!g2885) & (g2846)) + ((g827) & (!g1451) & (!g1485) & (g2845) & (g2885) & (!g2846)) + ((g827) & (!g1451) & (g1485) & (!g2845) & (!g2885) & (!g2846)) + ((g827) & (!g1451) & (g1485) & (!g2845) & (!g2885) & (g2846)) + ((g827) & (!g1451) & (g1485) & (g2845) & (!g2885) & (!g2846)) + ((g827) & (!g1451) & (g1485) & (g2845) & (g2885) & (g2846)) + ((g827) & (g1451) & (!g1485) & (!g2845) & (!g2885) & (g2846)) + ((g827) & (g1451) & (!g1485) & (!g2845) & (g2885) & (!g2846)) + ((g827) & (g1451) & (!g1485) & (g2845) & (!g2885) & (!g2846)) + ((g827) & (g1451) & (!g1485) & (g2845) & (!g2885) & (g2846)) + ((g827) & (g1451) & (g1485) & (!g2845) & (!g2885) & (!g2846)) + ((g827) & (g1451) & (g1485) & (!g2845) & (g2885) & (g2846)) + ((g827) & (g1451) & (g1485) & (g2845) & (g2885) & (!g2846)) + ((g827) & (g1451) & (g1485) & (g2845) & (g2885) & (g2846)));
	assign g8146 = (((!g3499) & (g5123) & (!g2887)) + ((!g3499) & (g5123) & (g2887)) + ((g3499) & (!g5123) & (g2887)) + ((g3499) & (g5123) & (g2887)));
	assign g2888 = (((!g827) & (!g1459) & (!g1487) & (!g2857) & (g2887) & (!g2858)) + ((!g827) & (!g1459) & (!g1487) & (!g2857) & (g2887) & (g2858)) + ((!g827) & (!g1459) & (!g1487) & (g2857) & (g2887) & (!g2858)) + ((!g827) & (!g1459) & (!g1487) & (g2857) & (g2887) & (g2858)) + ((!g827) & (!g1459) & (g1487) & (!g2857) & (g2887) & (!g2858)) + ((!g827) & (!g1459) & (g1487) & (!g2857) & (g2887) & (g2858)) + ((!g827) & (!g1459) & (g1487) & (g2857) & (g2887) & (!g2858)) + ((!g827) & (!g1459) & (g1487) & (g2857) & (g2887) & (g2858)) + ((!g827) & (g1459) & (!g1487) & (!g2857) & (g2887) & (!g2858)) + ((!g827) & (g1459) & (!g1487) & (!g2857) & (g2887) & (g2858)) + ((!g827) & (g1459) & (!g1487) & (g2857) & (g2887) & (!g2858)) + ((!g827) & (g1459) & (!g1487) & (g2857) & (g2887) & (g2858)) + ((!g827) & (g1459) & (g1487) & (!g2857) & (g2887) & (!g2858)) + ((!g827) & (g1459) & (g1487) & (!g2857) & (g2887) & (g2858)) + ((!g827) & (g1459) & (g1487) & (g2857) & (g2887) & (!g2858)) + ((!g827) & (g1459) & (g1487) & (g2857) & (g2887) & (g2858)) + ((g827) & (!g1459) & (!g1487) & (!g2857) & (g2887) & (!g2858)) + ((g827) & (!g1459) & (!g1487) & (!g2857) & (g2887) & (g2858)) + ((g827) & (!g1459) & (!g1487) & (g2857) & (!g2887) & (g2858)) + ((g827) & (!g1459) & (!g1487) & (g2857) & (g2887) & (!g2858)) + ((g827) & (!g1459) & (g1487) & (!g2857) & (!g2887) & (!g2858)) + ((g827) & (!g1459) & (g1487) & (!g2857) & (!g2887) & (g2858)) + ((g827) & (!g1459) & (g1487) & (g2857) & (!g2887) & (!g2858)) + ((g827) & (!g1459) & (g1487) & (g2857) & (g2887) & (g2858)) + ((g827) & (g1459) & (!g1487) & (!g2857) & (!g2887) & (g2858)) + ((g827) & (g1459) & (!g1487) & (!g2857) & (g2887) & (!g2858)) + ((g827) & (g1459) & (!g1487) & (g2857) & (!g2887) & (!g2858)) + ((g827) & (g1459) & (!g1487) & (g2857) & (!g2887) & (g2858)) + ((g827) & (g1459) & (g1487) & (!g2857) & (!g2887) & (!g2858)) + ((g827) & (g1459) & (g1487) & (!g2857) & (g2887) & (g2858)) + ((g827) & (g1459) & (g1487) & (g2857) & (g2887) & (!g2858)) + ((g827) & (g1459) & (g1487) & (g2857) & (g2887) & (g2858)));
	assign g8147 = (((!g3464) & (g5126) & (!g2889)) + ((!g3464) & (g5126) & (g2889)) + ((g3464) & (!g5126) & (g2889)) + ((g3464) & (g5126) & (g2889)));
	assign g2890 = (((!g827) & (!g1467) & (!g1489) & (!g2868) & (g2889) & (!g2869)) + ((!g827) & (!g1467) & (!g1489) & (!g2868) & (g2889) & (g2869)) + ((!g827) & (!g1467) & (!g1489) & (g2868) & (g2889) & (!g2869)) + ((!g827) & (!g1467) & (!g1489) & (g2868) & (g2889) & (g2869)) + ((!g827) & (!g1467) & (g1489) & (!g2868) & (g2889) & (!g2869)) + ((!g827) & (!g1467) & (g1489) & (!g2868) & (g2889) & (g2869)) + ((!g827) & (!g1467) & (g1489) & (g2868) & (g2889) & (!g2869)) + ((!g827) & (!g1467) & (g1489) & (g2868) & (g2889) & (g2869)) + ((!g827) & (g1467) & (!g1489) & (!g2868) & (g2889) & (!g2869)) + ((!g827) & (g1467) & (!g1489) & (!g2868) & (g2889) & (g2869)) + ((!g827) & (g1467) & (!g1489) & (g2868) & (g2889) & (!g2869)) + ((!g827) & (g1467) & (!g1489) & (g2868) & (g2889) & (g2869)) + ((!g827) & (g1467) & (g1489) & (!g2868) & (g2889) & (!g2869)) + ((!g827) & (g1467) & (g1489) & (!g2868) & (g2889) & (g2869)) + ((!g827) & (g1467) & (g1489) & (g2868) & (g2889) & (!g2869)) + ((!g827) & (g1467) & (g1489) & (g2868) & (g2889) & (g2869)) + ((g827) & (!g1467) & (!g1489) & (!g2868) & (g2889) & (!g2869)) + ((g827) & (!g1467) & (!g1489) & (!g2868) & (g2889) & (g2869)) + ((g827) & (!g1467) & (!g1489) & (g2868) & (!g2889) & (g2869)) + ((g827) & (!g1467) & (!g1489) & (g2868) & (g2889) & (!g2869)) + ((g827) & (!g1467) & (g1489) & (!g2868) & (!g2889) & (!g2869)) + ((g827) & (!g1467) & (g1489) & (!g2868) & (!g2889) & (g2869)) + ((g827) & (!g1467) & (g1489) & (g2868) & (!g2889) & (!g2869)) + ((g827) & (!g1467) & (g1489) & (g2868) & (g2889) & (g2869)) + ((g827) & (g1467) & (!g1489) & (!g2868) & (!g2889) & (g2869)) + ((g827) & (g1467) & (!g1489) & (!g2868) & (g2889) & (!g2869)) + ((g827) & (g1467) & (!g1489) & (g2868) & (!g2889) & (!g2869)) + ((g827) & (g1467) & (!g1489) & (g2868) & (!g2889) & (g2869)) + ((g827) & (g1467) & (g1489) & (!g2868) & (!g2889) & (!g2869)) + ((g827) & (g1467) & (g1489) & (!g2868) & (g2889) & (g2869)) + ((g827) & (g1467) & (g1489) & (g2868) & (g2889) & (!g2869)) + ((g827) & (g1467) & (g1489) & (g2868) & (g2889) & (g2869)));
	assign g8148 = (((!g3499) & (g5129) & (!g2891)) + ((!g3499) & (g5129) & (g2891)) + ((g3499) & (!g5129) & (g2891)) + ((g3499) & (g5129) & (g2891)));
	assign g2892 = (((!g827) & (!g1445) & (!g1491) & (!g2838) & (g2891) & (!g2839)) + ((!g827) & (!g1445) & (!g1491) & (!g2838) & (g2891) & (g2839)) + ((!g827) & (!g1445) & (!g1491) & (g2838) & (g2891) & (!g2839)) + ((!g827) & (!g1445) & (!g1491) & (g2838) & (g2891) & (g2839)) + ((!g827) & (!g1445) & (g1491) & (!g2838) & (g2891) & (!g2839)) + ((!g827) & (!g1445) & (g1491) & (!g2838) & (g2891) & (g2839)) + ((!g827) & (!g1445) & (g1491) & (g2838) & (g2891) & (!g2839)) + ((!g827) & (!g1445) & (g1491) & (g2838) & (g2891) & (g2839)) + ((!g827) & (g1445) & (!g1491) & (!g2838) & (g2891) & (!g2839)) + ((!g827) & (g1445) & (!g1491) & (!g2838) & (g2891) & (g2839)) + ((!g827) & (g1445) & (!g1491) & (g2838) & (g2891) & (!g2839)) + ((!g827) & (g1445) & (!g1491) & (g2838) & (g2891) & (g2839)) + ((!g827) & (g1445) & (g1491) & (!g2838) & (g2891) & (!g2839)) + ((!g827) & (g1445) & (g1491) & (!g2838) & (g2891) & (g2839)) + ((!g827) & (g1445) & (g1491) & (g2838) & (g2891) & (!g2839)) + ((!g827) & (g1445) & (g1491) & (g2838) & (g2891) & (g2839)) + ((g827) & (!g1445) & (!g1491) & (!g2838) & (g2891) & (!g2839)) + ((g827) & (!g1445) & (!g1491) & (!g2838) & (g2891) & (g2839)) + ((g827) & (!g1445) & (!g1491) & (g2838) & (!g2891) & (g2839)) + ((g827) & (!g1445) & (!g1491) & (g2838) & (g2891) & (!g2839)) + ((g827) & (!g1445) & (g1491) & (!g2838) & (!g2891) & (!g2839)) + ((g827) & (!g1445) & (g1491) & (!g2838) & (!g2891) & (g2839)) + ((g827) & (!g1445) & (g1491) & (g2838) & (!g2891) & (!g2839)) + ((g827) & (!g1445) & (g1491) & (g2838) & (g2891) & (g2839)) + ((g827) & (g1445) & (!g1491) & (!g2838) & (!g2891) & (g2839)) + ((g827) & (g1445) & (!g1491) & (!g2838) & (g2891) & (!g2839)) + ((g827) & (g1445) & (!g1491) & (g2838) & (!g2891) & (!g2839)) + ((g827) & (g1445) & (!g1491) & (g2838) & (!g2891) & (g2839)) + ((g827) & (g1445) & (g1491) & (!g2838) & (!g2891) & (!g2839)) + ((g827) & (g1445) & (g1491) & (!g2838) & (g2891) & (g2839)) + ((g827) & (g1445) & (g1491) & (g2838) & (g2891) & (!g2839)) + ((g827) & (g1445) & (g1491) & (g2838) & (g2891) & (g2839)));
	assign g8149 = (((!g3464) & (g5133) & (!g2893)) + ((!g3464) & (g5133) & (g2893)) + ((g3464) & (!g5133) & (g2893)) + ((g3464) & (g5133) & (g2893)));
	assign g2894 = (((!g827) & (!g1453) & (!g1493) & (!g2848) & (g2893) & (!g2849)) + ((!g827) & (!g1453) & (!g1493) & (!g2848) & (g2893) & (g2849)) + ((!g827) & (!g1453) & (!g1493) & (g2848) & (g2893) & (!g2849)) + ((!g827) & (!g1453) & (!g1493) & (g2848) & (g2893) & (g2849)) + ((!g827) & (!g1453) & (g1493) & (!g2848) & (g2893) & (!g2849)) + ((!g827) & (!g1453) & (g1493) & (!g2848) & (g2893) & (g2849)) + ((!g827) & (!g1453) & (g1493) & (g2848) & (g2893) & (!g2849)) + ((!g827) & (!g1453) & (g1493) & (g2848) & (g2893) & (g2849)) + ((!g827) & (g1453) & (!g1493) & (!g2848) & (g2893) & (!g2849)) + ((!g827) & (g1453) & (!g1493) & (!g2848) & (g2893) & (g2849)) + ((!g827) & (g1453) & (!g1493) & (g2848) & (g2893) & (!g2849)) + ((!g827) & (g1453) & (!g1493) & (g2848) & (g2893) & (g2849)) + ((!g827) & (g1453) & (g1493) & (!g2848) & (g2893) & (!g2849)) + ((!g827) & (g1453) & (g1493) & (!g2848) & (g2893) & (g2849)) + ((!g827) & (g1453) & (g1493) & (g2848) & (g2893) & (!g2849)) + ((!g827) & (g1453) & (g1493) & (g2848) & (g2893) & (g2849)) + ((g827) & (!g1453) & (!g1493) & (!g2848) & (g2893) & (!g2849)) + ((g827) & (!g1453) & (!g1493) & (!g2848) & (g2893) & (g2849)) + ((g827) & (!g1453) & (!g1493) & (g2848) & (!g2893) & (g2849)) + ((g827) & (!g1453) & (!g1493) & (g2848) & (g2893) & (!g2849)) + ((g827) & (!g1453) & (g1493) & (!g2848) & (!g2893) & (!g2849)) + ((g827) & (!g1453) & (g1493) & (!g2848) & (!g2893) & (g2849)) + ((g827) & (!g1453) & (g1493) & (g2848) & (!g2893) & (!g2849)) + ((g827) & (!g1453) & (g1493) & (g2848) & (g2893) & (g2849)) + ((g827) & (g1453) & (!g1493) & (!g2848) & (!g2893) & (g2849)) + ((g827) & (g1453) & (!g1493) & (!g2848) & (g2893) & (!g2849)) + ((g827) & (g1453) & (!g1493) & (g2848) & (!g2893) & (!g2849)) + ((g827) & (g1453) & (!g1493) & (g2848) & (!g2893) & (g2849)) + ((g827) & (g1453) & (g1493) & (!g2848) & (!g2893) & (!g2849)) + ((g827) & (g1453) & (g1493) & (!g2848) & (g2893) & (g2849)) + ((g827) & (g1453) & (g1493) & (g2848) & (g2893) & (!g2849)) + ((g827) & (g1453) & (g1493) & (g2848) & (g2893) & (g2849)));
	assign g8150 = (((!g2017) & (g5138) & (!g2895)) + ((!g2017) & (g5138) & (g2895)) + ((g2017) & (!g5138) & (g2895)) + ((g2017) & (g5138) & (g2895)));
	assign g2896 = (((!g827) & (!g1461) & (!g1495) & (!g2860) & (g2895) & (!g2861)) + ((!g827) & (!g1461) & (!g1495) & (!g2860) & (g2895) & (g2861)) + ((!g827) & (!g1461) & (!g1495) & (g2860) & (g2895) & (!g2861)) + ((!g827) & (!g1461) & (!g1495) & (g2860) & (g2895) & (g2861)) + ((!g827) & (!g1461) & (g1495) & (!g2860) & (g2895) & (!g2861)) + ((!g827) & (!g1461) & (g1495) & (!g2860) & (g2895) & (g2861)) + ((!g827) & (!g1461) & (g1495) & (g2860) & (g2895) & (!g2861)) + ((!g827) & (!g1461) & (g1495) & (g2860) & (g2895) & (g2861)) + ((!g827) & (g1461) & (!g1495) & (!g2860) & (g2895) & (!g2861)) + ((!g827) & (g1461) & (!g1495) & (!g2860) & (g2895) & (g2861)) + ((!g827) & (g1461) & (!g1495) & (g2860) & (g2895) & (!g2861)) + ((!g827) & (g1461) & (!g1495) & (g2860) & (g2895) & (g2861)) + ((!g827) & (g1461) & (g1495) & (!g2860) & (g2895) & (!g2861)) + ((!g827) & (g1461) & (g1495) & (!g2860) & (g2895) & (g2861)) + ((!g827) & (g1461) & (g1495) & (g2860) & (g2895) & (!g2861)) + ((!g827) & (g1461) & (g1495) & (g2860) & (g2895) & (g2861)) + ((g827) & (!g1461) & (!g1495) & (!g2860) & (g2895) & (!g2861)) + ((g827) & (!g1461) & (!g1495) & (!g2860) & (g2895) & (g2861)) + ((g827) & (!g1461) & (!g1495) & (g2860) & (!g2895) & (g2861)) + ((g827) & (!g1461) & (!g1495) & (g2860) & (g2895) & (!g2861)) + ((g827) & (!g1461) & (g1495) & (!g2860) & (!g2895) & (!g2861)) + ((g827) & (!g1461) & (g1495) & (!g2860) & (!g2895) & (g2861)) + ((g827) & (!g1461) & (g1495) & (g2860) & (!g2895) & (!g2861)) + ((g827) & (!g1461) & (g1495) & (g2860) & (g2895) & (g2861)) + ((g827) & (g1461) & (!g1495) & (!g2860) & (!g2895) & (g2861)) + ((g827) & (g1461) & (!g1495) & (!g2860) & (g2895) & (!g2861)) + ((g827) & (g1461) & (!g1495) & (g2860) & (!g2895) & (!g2861)) + ((g827) & (g1461) & (!g1495) & (g2860) & (!g2895) & (g2861)) + ((g827) & (g1461) & (g1495) & (!g2860) & (!g2895) & (!g2861)) + ((g827) & (g1461) & (g1495) & (!g2860) & (g2895) & (g2861)) + ((g827) & (g1461) & (g1495) & (g2860) & (g2895) & (!g2861)) + ((g827) & (g1461) & (g1495) & (g2860) & (g2895) & (g2861)));
	assign g8151 = (((!g3429) & (g5143) & (!g2897)) + ((!g3429) & (g5143) & (g2897)) + ((g3429) & (!g5143) & (g2897)) + ((g3429) & (g5143) & (g2897)));
	assign g2898 = (((!g827) & (!g1469) & (!g1497) & (!g2871) & (g2897) & (!g2872)) + ((!g827) & (!g1469) & (!g1497) & (!g2871) & (g2897) & (g2872)) + ((!g827) & (!g1469) & (!g1497) & (g2871) & (g2897) & (!g2872)) + ((!g827) & (!g1469) & (!g1497) & (g2871) & (g2897) & (g2872)) + ((!g827) & (!g1469) & (g1497) & (!g2871) & (g2897) & (!g2872)) + ((!g827) & (!g1469) & (g1497) & (!g2871) & (g2897) & (g2872)) + ((!g827) & (!g1469) & (g1497) & (g2871) & (g2897) & (!g2872)) + ((!g827) & (!g1469) & (g1497) & (g2871) & (g2897) & (g2872)) + ((!g827) & (g1469) & (!g1497) & (!g2871) & (g2897) & (!g2872)) + ((!g827) & (g1469) & (!g1497) & (!g2871) & (g2897) & (g2872)) + ((!g827) & (g1469) & (!g1497) & (g2871) & (g2897) & (!g2872)) + ((!g827) & (g1469) & (!g1497) & (g2871) & (g2897) & (g2872)) + ((!g827) & (g1469) & (g1497) & (!g2871) & (g2897) & (!g2872)) + ((!g827) & (g1469) & (g1497) & (!g2871) & (g2897) & (g2872)) + ((!g827) & (g1469) & (g1497) & (g2871) & (g2897) & (!g2872)) + ((!g827) & (g1469) & (g1497) & (g2871) & (g2897) & (g2872)) + ((g827) & (!g1469) & (!g1497) & (!g2871) & (g2897) & (!g2872)) + ((g827) & (!g1469) & (!g1497) & (!g2871) & (g2897) & (g2872)) + ((g827) & (!g1469) & (!g1497) & (g2871) & (!g2897) & (g2872)) + ((g827) & (!g1469) & (!g1497) & (g2871) & (g2897) & (!g2872)) + ((g827) & (!g1469) & (g1497) & (!g2871) & (!g2897) & (!g2872)) + ((g827) & (!g1469) & (g1497) & (!g2871) & (!g2897) & (g2872)) + ((g827) & (!g1469) & (g1497) & (g2871) & (!g2897) & (!g2872)) + ((g827) & (!g1469) & (g1497) & (g2871) & (g2897) & (g2872)) + ((g827) & (g1469) & (!g1497) & (!g2871) & (!g2897) & (g2872)) + ((g827) & (g1469) & (!g1497) & (!g2871) & (g2897) & (!g2872)) + ((g827) & (g1469) & (!g1497) & (g2871) & (!g2897) & (!g2872)) + ((g827) & (g1469) & (!g1497) & (g2871) & (!g2897) & (g2872)) + ((g827) & (g1469) & (g1497) & (!g2871) & (!g2897) & (!g2872)) + ((g827) & (g1469) & (g1497) & (!g2871) & (g2897) & (g2872)) + ((g827) & (g1469) & (g1497) & (g2871) & (g2897) & (!g2872)) + ((g827) & (g1469) & (g1497) & (g2871) & (g2897) & (g2872)));
	assign g2899 = (((!g827) & (!g1447) & (!g1499) & (!g2211) & (g2257) & (!g2841)) + ((!g827) & (!g1447) & (!g1499) & (!g2211) & (g2257) & (g2841)) + ((!g827) & (!g1447) & (!g1499) & (g2211) & (g2257) & (!g2841)) + ((!g827) & (!g1447) & (!g1499) & (g2211) & (g2257) & (g2841)) + ((!g827) & (!g1447) & (g1499) & (!g2211) & (g2257) & (!g2841)) + ((!g827) & (!g1447) & (g1499) & (!g2211) & (g2257) & (g2841)) + ((!g827) & (!g1447) & (g1499) & (g2211) & (g2257) & (!g2841)) + ((!g827) & (!g1447) & (g1499) & (g2211) & (g2257) & (g2841)) + ((!g827) & (g1447) & (!g1499) & (!g2211) & (g2257) & (!g2841)) + ((!g827) & (g1447) & (!g1499) & (!g2211) & (g2257) & (g2841)) + ((!g827) & (g1447) & (!g1499) & (g2211) & (g2257) & (!g2841)) + ((!g827) & (g1447) & (!g1499) & (g2211) & (g2257) & (g2841)) + ((!g827) & (g1447) & (g1499) & (!g2211) & (g2257) & (!g2841)) + ((!g827) & (g1447) & (g1499) & (!g2211) & (g2257) & (g2841)) + ((!g827) & (g1447) & (g1499) & (g2211) & (g2257) & (!g2841)) + ((!g827) & (g1447) & (g1499) & (g2211) & (g2257) & (g2841)) + ((g827) & (!g1447) & (!g1499) & (!g2211) & (g2257) & (!g2841)) + ((g827) & (!g1447) & (!g1499) & (!g2211) & (g2257) & (g2841)) + ((g827) & (!g1447) & (!g1499) & (g2211) & (!g2257) & (g2841)) + ((g827) & (!g1447) & (!g1499) & (g2211) & (g2257) & (!g2841)) + ((g827) & (!g1447) & (g1499) & (!g2211) & (!g2257) & (!g2841)) + ((g827) & (!g1447) & (g1499) & (!g2211) & (!g2257) & (g2841)) + ((g827) & (!g1447) & (g1499) & (g2211) & (!g2257) & (!g2841)) + ((g827) & (!g1447) & (g1499) & (g2211) & (g2257) & (g2841)) + ((g827) & (g1447) & (!g1499) & (!g2211) & (!g2257) & (g2841)) + ((g827) & (g1447) & (!g1499) & (!g2211) & (g2257) & (!g2841)) + ((g827) & (g1447) & (!g1499) & (g2211) & (!g2257) & (!g2841)) + ((g827) & (g1447) & (!g1499) & (g2211) & (!g2257) & (g2841)) + ((g827) & (g1447) & (g1499) & (!g2211) & (!g2257) & (!g2841)) + ((g827) & (g1447) & (g1499) & (!g2211) & (g2257) & (g2841)) + ((g827) & (g1447) & (g1499) & (g2211) & (g2257) & (!g2841)) + ((g827) & (g1447) & (g1499) & (g2211) & (g2257) & (g2841)));
	assign g8152 = (((!g3499) & (g5146) & (!g2900)) + ((!g3499) & (g5146) & (g2900)) + ((g3499) & (!g5146) & (g2900)) + ((g3499) & (g5146) & (g2900)));
	assign g2901 = (((!g827) & (!g1455) & (!g1501) & (!g2851) & (g2900) & (!g2852)) + ((!g827) & (!g1455) & (!g1501) & (!g2851) & (g2900) & (g2852)) + ((!g827) & (!g1455) & (!g1501) & (g2851) & (g2900) & (!g2852)) + ((!g827) & (!g1455) & (!g1501) & (g2851) & (g2900) & (g2852)) + ((!g827) & (!g1455) & (g1501) & (!g2851) & (g2900) & (!g2852)) + ((!g827) & (!g1455) & (g1501) & (!g2851) & (g2900) & (g2852)) + ((!g827) & (!g1455) & (g1501) & (g2851) & (g2900) & (!g2852)) + ((!g827) & (!g1455) & (g1501) & (g2851) & (g2900) & (g2852)) + ((!g827) & (g1455) & (!g1501) & (!g2851) & (g2900) & (!g2852)) + ((!g827) & (g1455) & (!g1501) & (!g2851) & (g2900) & (g2852)) + ((!g827) & (g1455) & (!g1501) & (g2851) & (g2900) & (!g2852)) + ((!g827) & (g1455) & (!g1501) & (g2851) & (g2900) & (g2852)) + ((!g827) & (g1455) & (g1501) & (!g2851) & (g2900) & (!g2852)) + ((!g827) & (g1455) & (g1501) & (!g2851) & (g2900) & (g2852)) + ((!g827) & (g1455) & (g1501) & (g2851) & (g2900) & (!g2852)) + ((!g827) & (g1455) & (g1501) & (g2851) & (g2900) & (g2852)) + ((g827) & (!g1455) & (!g1501) & (!g2851) & (g2900) & (!g2852)) + ((g827) & (!g1455) & (!g1501) & (!g2851) & (g2900) & (g2852)) + ((g827) & (!g1455) & (!g1501) & (g2851) & (!g2900) & (g2852)) + ((g827) & (!g1455) & (!g1501) & (g2851) & (g2900) & (!g2852)) + ((g827) & (!g1455) & (g1501) & (!g2851) & (!g2900) & (!g2852)) + ((g827) & (!g1455) & (g1501) & (!g2851) & (!g2900) & (g2852)) + ((g827) & (!g1455) & (g1501) & (g2851) & (!g2900) & (!g2852)) + ((g827) & (!g1455) & (g1501) & (g2851) & (g2900) & (g2852)) + ((g827) & (g1455) & (!g1501) & (!g2851) & (!g2900) & (g2852)) + ((g827) & (g1455) & (!g1501) & (!g2851) & (g2900) & (!g2852)) + ((g827) & (g1455) & (!g1501) & (g2851) & (!g2900) & (!g2852)) + ((g827) & (g1455) & (!g1501) & (g2851) & (!g2900) & (g2852)) + ((g827) & (g1455) & (g1501) & (!g2851) & (!g2900) & (!g2852)) + ((g827) & (g1455) & (g1501) & (!g2851) & (g2900) & (g2852)) + ((g827) & (g1455) & (g1501) & (g2851) & (g2900) & (!g2852)) + ((g827) & (g1455) & (g1501) & (g2851) & (g2900) & (g2852)));
	assign g8153 = (((!g3429) & (g5151) & (!g2902)) + ((!g3429) & (g5151) & (g2902)) + ((g3429) & (!g5151) & (g2902)) + ((g3429) & (g5151) & (g2902)));
	assign g2903 = (((!g827) & (!g1463) & (!g1503) & (!g2863) & (g2902) & (!g2864)) + ((!g827) & (!g1463) & (!g1503) & (!g2863) & (g2902) & (g2864)) + ((!g827) & (!g1463) & (!g1503) & (g2863) & (g2902) & (!g2864)) + ((!g827) & (!g1463) & (!g1503) & (g2863) & (g2902) & (g2864)) + ((!g827) & (!g1463) & (g1503) & (!g2863) & (g2902) & (!g2864)) + ((!g827) & (!g1463) & (g1503) & (!g2863) & (g2902) & (g2864)) + ((!g827) & (!g1463) & (g1503) & (g2863) & (g2902) & (!g2864)) + ((!g827) & (!g1463) & (g1503) & (g2863) & (g2902) & (g2864)) + ((!g827) & (g1463) & (!g1503) & (!g2863) & (g2902) & (!g2864)) + ((!g827) & (g1463) & (!g1503) & (!g2863) & (g2902) & (g2864)) + ((!g827) & (g1463) & (!g1503) & (g2863) & (g2902) & (!g2864)) + ((!g827) & (g1463) & (!g1503) & (g2863) & (g2902) & (g2864)) + ((!g827) & (g1463) & (g1503) & (!g2863) & (g2902) & (!g2864)) + ((!g827) & (g1463) & (g1503) & (!g2863) & (g2902) & (g2864)) + ((!g827) & (g1463) & (g1503) & (g2863) & (g2902) & (!g2864)) + ((!g827) & (g1463) & (g1503) & (g2863) & (g2902) & (g2864)) + ((g827) & (!g1463) & (!g1503) & (!g2863) & (g2902) & (!g2864)) + ((g827) & (!g1463) & (!g1503) & (!g2863) & (g2902) & (g2864)) + ((g827) & (!g1463) & (!g1503) & (g2863) & (!g2902) & (g2864)) + ((g827) & (!g1463) & (!g1503) & (g2863) & (g2902) & (!g2864)) + ((g827) & (!g1463) & (g1503) & (!g2863) & (!g2902) & (!g2864)) + ((g827) & (!g1463) & (g1503) & (!g2863) & (!g2902) & (g2864)) + ((g827) & (!g1463) & (g1503) & (g2863) & (!g2902) & (!g2864)) + ((g827) & (!g1463) & (g1503) & (g2863) & (g2902) & (g2864)) + ((g827) & (g1463) & (!g1503) & (!g2863) & (!g2902) & (g2864)) + ((g827) & (g1463) & (!g1503) & (!g2863) & (g2902) & (!g2864)) + ((g827) & (g1463) & (!g1503) & (g2863) & (!g2902) & (!g2864)) + ((g827) & (g1463) & (!g1503) & (g2863) & (!g2902) & (g2864)) + ((g827) & (g1463) & (g1503) & (!g2863) & (!g2902) & (!g2864)) + ((g827) & (g1463) & (g1503) & (!g2863) & (g2902) & (g2864)) + ((g827) & (g1463) & (g1503) & (g2863) & (g2902) & (!g2864)) + ((g827) & (g1463) & (g1503) & (g2863) & (g2902) & (g2864)));
	assign g8154 = (((!g2017) & (g5156) & (!g2904)) + ((!g2017) & (g5156) & (g2904)) + ((g2017) & (!g5156) & (g2904)) + ((g2017) & (g5156) & (g2904)));
	assign g2905 = (((!g827) & (!g1471) & (!g1505) & (!g2874) & (g2904) & (!g2875)) + ((!g827) & (!g1471) & (!g1505) & (!g2874) & (g2904) & (g2875)) + ((!g827) & (!g1471) & (!g1505) & (g2874) & (g2904) & (!g2875)) + ((!g827) & (!g1471) & (!g1505) & (g2874) & (g2904) & (g2875)) + ((!g827) & (!g1471) & (g1505) & (!g2874) & (g2904) & (!g2875)) + ((!g827) & (!g1471) & (g1505) & (!g2874) & (g2904) & (g2875)) + ((!g827) & (!g1471) & (g1505) & (g2874) & (g2904) & (!g2875)) + ((!g827) & (!g1471) & (g1505) & (g2874) & (g2904) & (g2875)) + ((!g827) & (g1471) & (!g1505) & (!g2874) & (g2904) & (!g2875)) + ((!g827) & (g1471) & (!g1505) & (!g2874) & (g2904) & (g2875)) + ((!g827) & (g1471) & (!g1505) & (g2874) & (g2904) & (!g2875)) + ((!g827) & (g1471) & (!g1505) & (g2874) & (g2904) & (g2875)) + ((!g827) & (g1471) & (g1505) & (!g2874) & (g2904) & (!g2875)) + ((!g827) & (g1471) & (g1505) & (!g2874) & (g2904) & (g2875)) + ((!g827) & (g1471) & (g1505) & (g2874) & (g2904) & (!g2875)) + ((!g827) & (g1471) & (g1505) & (g2874) & (g2904) & (g2875)) + ((g827) & (!g1471) & (!g1505) & (!g2874) & (g2904) & (!g2875)) + ((g827) & (!g1471) & (!g1505) & (!g2874) & (g2904) & (g2875)) + ((g827) & (!g1471) & (!g1505) & (g2874) & (!g2904) & (g2875)) + ((g827) & (!g1471) & (!g1505) & (g2874) & (g2904) & (!g2875)) + ((g827) & (!g1471) & (g1505) & (!g2874) & (!g2904) & (!g2875)) + ((g827) & (!g1471) & (g1505) & (!g2874) & (!g2904) & (g2875)) + ((g827) & (!g1471) & (g1505) & (g2874) & (!g2904) & (!g2875)) + ((g827) & (!g1471) & (g1505) & (g2874) & (g2904) & (g2875)) + ((g827) & (g1471) & (!g1505) & (!g2874) & (!g2904) & (g2875)) + ((g827) & (g1471) & (!g1505) & (!g2874) & (g2904) & (!g2875)) + ((g827) & (g1471) & (!g1505) & (g2874) & (!g2904) & (!g2875)) + ((g827) & (g1471) & (!g1505) & (g2874) & (!g2904) & (g2875)) + ((g827) & (g1471) & (g1505) & (!g2874) & (!g2904) & (!g2875)) + ((g827) & (g1471) & (g1505) & (!g2874) & (g2904) & (g2875)) + ((g827) & (g1471) & (g1505) & (g2874) & (g2904) & (!g2875)) + ((g827) & (g1471) & (g1505) & (g2874) & (g2904) & (g2875)));
	assign g2906 = (((!g1890) & (!g1906) & (g1939) & (g1940)) + ((!g1890) & (g1906) & (g1939) & (g1940)) + ((g1890) & (!g1906) & (g1939) & (g1940)) + ((g1890) & (g1906) & (!g1939) & (g1940)) + ((g1890) & (g1906) & (g1939) & (!g1940)) + ((g1890) & (g1906) & (g1939) & (g1940)));
	assign g2907 = (((g1914) & (!g2906) & (!g1941) & (g1942)) + ((g1914) & (!g2906) & (g1941) & (!g1942)) + ((g1914) & (g2906) & (!g1941) & (!g1942)) + ((g1914) & (g2906) & (g1941) & (g1942)));
	assign g2908 = (((!g1884) & (!g1888) & (g1977) & (g1978)) + ((!g1884) & (g1888) & (g1977) & (g1978)) + ((g1884) & (!g1888) & (g1977) & (g1978)) + ((g1884) & (g1888) & (!g1977) & (g1978)) + ((g1884) & (g1888) & (g1977) & (!g1978)) + ((g1884) & (g1888) & (g1977) & (g1978)));
	assign g2909 = (((!g1914) & (!g2908) & (!g1979) & (g1980)) + ((!g1914) & (!g2908) & (g1979) & (!g1980)) + ((!g1914) & (g2908) & (!g1979) & (!g1980)) + ((!g1914) & (g2908) & (g1979) & (g1980)));
	assign g2910 = (((!g830) & (!g2907) & (!g2909) & (!g1507)) + ((!g830) & (!g2907) & (!g2909) & (g1507)) + ((!g830) & (!g2907) & (g2909) & (!g1507)) + ((!g830) & (!g2907) & (g2909) & (g1507)) + ((!g830) & (g2907) & (!g2909) & (!g1507)) + ((!g830) & (g2907) & (!g2909) & (g1507)) + ((!g830) & (g2907) & (g2909) & (!g1507)) + ((!g830) & (g2907) & (g2909) & (g1507)) + ((g830) & (!g2907) & (!g2909) & (g1507)) + ((g830) & (!g2907) & (g2909) & (!g1507)) + ((g830) & (g2907) & (!g2909) & (!g1507)) + ((g830) & (g2907) & (g2909) & (!g1507)));
	assign g2911 = (((!g1483) & (g2256)) + ((g1483) & (!g2256)));
	assign g2912 = (((!g1415) & (!g1443) & (g2177) & (g2210) & (!g2802) & (g2911)) + ((!g1415) & (g1443) & (!g2177) & (g2210) & (!g2802) & (g2911)) + ((!g1415) & (g1443) & (!g2177) & (g2210) & (g2802) & (g2911)) + ((!g1415) & (g1443) & (g2177) & (!g2210) & (!g2802) & (g2911)) + ((!g1415) & (g1443) & (g2177) & (g2210) & (!g2802) & (g2911)) + ((!g1415) & (g1443) & (g2177) & (g2210) & (g2802) & (g2911)) + ((g1415) & (!g1443) & (!g2177) & (g2210) & (!g2802) & (g2911)) + ((g1415) & (!g1443) & (g2177) & (g2210) & (!g2802) & (g2911)) + ((g1415) & (!g1443) & (g2177) & (g2210) & (g2802) & (g2911)) + ((g1415) & (g1443) & (!g2177) & (!g2210) & (!g2802) & (g2911)) + ((g1415) & (g1443) & (!g2177) & (g2210) & (!g2802) & (g2911)) + ((g1415) & (g1443) & (!g2177) & (g2210) & (g2802) & (g2911)) + ((g1415) & (g1443) & (g2177) & (!g2210) & (!g2802) & (g2911)) + ((g1415) & (g1443) & (g2177) & (!g2210) & (g2802) & (g2911)) + ((g1415) & (g1443) & (g2177) & (g2210) & (!g2802) & (g2911)) + ((g1415) & (g1443) & (g2177) & (g2210) & (g2802) & (g2911)));
	assign g2913 = (((g1483) & (g2256)));
	assign g2914 = (((!g2912) & (!g2913)));
	assign g2915 = (((!g827) & (!g1510) & (g2295) & (!g2914)) + ((!g827) & (!g1510) & (g2295) & (g2914)) + ((!g827) & (g1510) & (g2295) & (!g2914)) + ((!g827) & (g1510) & (g2295) & (g2914)) + ((g827) & (!g1510) & (!g2295) & (!g2914)) + ((g827) & (!g1510) & (g2295) & (g2914)) + ((g827) & (g1510) & (!g2295) & (g2914)) + ((g827) & (g1510) & (g2295) & (!g2914)));
	assign g8155 = (((!g3499) & (g5160) & (!g2916)) + ((!g3499) & (g5160) & (g2916)) + ((g3499) & (!g5160) & (g2916)) + ((g3499) & (g5160) & (g2916)));
	assign g2917 = (((!g1491) & (g2891)) + ((g1491) & (!g2891)));
	assign g2918 = (((!g1423) & (!g1445) & (g2813) & (g2838) & (!g2814) & (g2917)) + ((!g1423) & (g1445) & (!g2813) & (g2838) & (!g2814) & (g2917)) + ((!g1423) & (g1445) & (!g2813) & (g2838) & (g2814) & (g2917)) + ((!g1423) & (g1445) & (g2813) & (!g2838) & (!g2814) & (g2917)) + ((!g1423) & (g1445) & (g2813) & (g2838) & (!g2814) & (g2917)) + ((!g1423) & (g1445) & (g2813) & (g2838) & (g2814) & (g2917)) + ((g1423) & (!g1445) & (!g2813) & (g2838) & (!g2814) & (g2917)) + ((g1423) & (!g1445) & (g2813) & (g2838) & (!g2814) & (g2917)) + ((g1423) & (!g1445) & (g2813) & (g2838) & (g2814) & (g2917)) + ((g1423) & (g1445) & (!g2813) & (!g2838) & (!g2814) & (g2917)) + ((g1423) & (g1445) & (!g2813) & (g2838) & (!g2814) & (g2917)) + ((g1423) & (g1445) & (!g2813) & (g2838) & (g2814) & (g2917)) + ((g1423) & (g1445) & (g2813) & (!g2838) & (!g2814) & (g2917)) + ((g1423) & (g1445) & (g2813) & (!g2838) & (g2814) & (g2917)) + ((g1423) & (g1445) & (g2813) & (g2838) & (!g2814) & (g2917)) + ((g1423) & (g1445) & (g2813) & (g2838) & (g2814) & (g2917)));
	assign g2919 = (((g1491) & (g2891)));
	assign g2920 = (((!g2918) & (!g2919)));
	assign g2921 = (((!g827) & (!g1512) & (g2916) & (!g2920)) + ((!g827) & (!g1512) & (g2916) & (g2920)) + ((!g827) & (g1512) & (g2916) & (!g2920)) + ((!g827) & (g1512) & (g2916) & (g2920)) + ((g827) & (!g1512) & (!g2916) & (!g2920)) + ((g827) & (!g1512) & (g2916) & (g2920)) + ((g827) & (g1512) & (!g2916) & (g2920)) + ((g827) & (g1512) & (g2916) & (!g2920)));
	assign g2922 = (((!g1499) & (g2257)) + ((g1499) & (!g2257)));
	assign g2923 = (((!g1431) & (!g1447) & (g2178) & (g2211) & (!g2825) & (g2922)) + ((!g1431) & (g1447) & (!g2178) & (g2211) & (!g2825) & (g2922)) + ((!g1431) & (g1447) & (!g2178) & (g2211) & (g2825) & (g2922)) + ((!g1431) & (g1447) & (g2178) & (!g2211) & (!g2825) & (g2922)) + ((!g1431) & (g1447) & (g2178) & (g2211) & (!g2825) & (g2922)) + ((!g1431) & (g1447) & (g2178) & (g2211) & (g2825) & (g2922)) + ((g1431) & (!g1447) & (!g2178) & (g2211) & (!g2825) & (g2922)) + ((g1431) & (!g1447) & (g2178) & (g2211) & (!g2825) & (g2922)) + ((g1431) & (!g1447) & (g2178) & (g2211) & (g2825) & (g2922)) + ((g1431) & (g1447) & (!g2178) & (!g2211) & (!g2825) & (g2922)) + ((g1431) & (g1447) & (!g2178) & (g2211) & (!g2825) & (g2922)) + ((g1431) & (g1447) & (!g2178) & (g2211) & (g2825) & (g2922)) + ((g1431) & (g1447) & (g2178) & (!g2211) & (!g2825) & (g2922)) + ((g1431) & (g1447) & (g2178) & (!g2211) & (g2825) & (g2922)) + ((g1431) & (g1447) & (g2178) & (g2211) & (!g2825) & (g2922)) + ((g1431) & (g1447) & (g2178) & (g2211) & (g2825) & (g2922)));
	assign g2924 = (((g1499) & (g2257)));
	assign g2925 = (((!g2923) & (!g2924)));
	assign g2926 = (((!g827) & (!g1514) & (g2296) & (!g2925)) + ((!g827) & (!g1514) & (g2296) & (g2925)) + ((!g827) & (g1514) & (g2296) & (!g2925)) + ((!g827) & (g1514) & (g2296) & (g2925)) + ((g827) & (!g1514) & (!g2296) & (!g2925)) + ((g827) & (!g1514) & (g2296) & (g2925)) + ((g827) & (g1514) & (!g2296) & (g2925)) + ((g827) & (g1514) & (g2296) & (!g2925)));
	assign g2927 = (((!g1477) & (g2262)) + ((g1477) & (!g2262)));
	assign g2928 = (((!g1409) & (!g1449) & (g2180) & (g2212) & (!g2795) & (g2927)) + ((!g1409) & (g1449) & (!g2180) & (g2212) & (!g2795) & (g2927)) + ((!g1409) & (g1449) & (!g2180) & (g2212) & (g2795) & (g2927)) + ((!g1409) & (g1449) & (g2180) & (!g2212) & (!g2795) & (g2927)) + ((!g1409) & (g1449) & (g2180) & (g2212) & (!g2795) & (g2927)) + ((!g1409) & (g1449) & (g2180) & (g2212) & (g2795) & (g2927)) + ((g1409) & (!g1449) & (!g2180) & (g2212) & (!g2795) & (g2927)) + ((g1409) & (!g1449) & (g2180) & (g2212) & (!g2795) & (g2927)) + ((g1409) & (!g1449) & (g2180) & (g2212) & (g2795) & (g2927)) + ((g1409) & (g1449) & (!g2180) & (!g2212) & (!g2795) & (g2927)) + ((g1409) & (g1449) & (!g2180) & (g2212) & (!g2795) & (g2927)) + ((g1409) & (g1449) & (!g2180) & (g2212) & (g2795) & (g2927)) + ((g1409) & (g1449) & (g2180) & (!g2212) & (!g2795) & (g2927)) + ((g1409) & (g1449) & (g2180) & (!g2212) & (g2795) & (g2927)) + ((g1409) & (g1449) & (g2180) & (g2212) & (!g2795) & (g2927)) + ((g1409) & (g1449) & (g2180) & (g2212) & (g2795) & (g2927)));
	assign g2929 = (((g1477) & (g2262)));
	assign g2930 = (((!g2928) & (!g2929)));
	assign g2931 = (((!g827) & (!g1516) & (g2298) & (!g2930)) + ((!g827) & (!g1516) & (g2298) & (g2930)) + ((!g827) & (g1516) & (g2298) & (!g2930)) + ((!g827) & (g1516) & (g2298) & (g2930)) + ((g827) & (!g1516) & (!g2298) & (!g2930)) + ((g827) & (!g1516) & (g2298) & (g2930)) + ((g827) & (g1516) & (!g2298) & (g2930)) + ((g827) & (g1516) & (g2298) & (!g2930)));
	assign g8156 = (((!g2017) & (g6174) & (!g2932)) + ((!g2017) & (g6174) & (g2932)) + ((g2017) & (!g6174) & (g2932)) + ((g2017) & (g6174) & (g2932)));
	assign g2933 = (((!g1485) & (g2885)) + ((g1485) & (!g2885)));
	assign g2934 = (((!g1417) & (!g1451) & (g2804) & (g2845) & (!g2805) & (g2933)) + ((!g1417) & (g1451) & (!g2804) & (g2845) & (!g2805) & (g2933)) + ((!g1417) & (g1451) & (!g2804) & (g2845) & (g2805) & (g2933)) + ((!g1417) & (g1451) & (g2804) & (!g2845) & (!g2805) & (g2933)) + ((!g1417) & (g1451) & (g2804) & (g2845) & (!g2805) & (g2933)) + ((!g1417) & (g1451) & (g2804) & (g2845) & (g2805) & (g2933)) + ((g1417) & (!g1451) & (!g2804) & (g2845) & (!g2805) & (g2933)) + ((g1417) & (!g1451) & (g2804) & (g2845) & (!g2805) & (g2933)) + ((g1417) & (!g1451) & (g2804) & (g2845) & (g2805) & (g2933)) + ((g1417) & (g1451) & (!g2804) & (!g2845) & (!g2805) & (g2933)) + ((g1417) & (g1451) & (!g2804) & (g2845) & (!g2805) & (g2933)) + ((g1417) & (g1451) & (!g2804) & (g2845) & (g2805) & (g2933)) + ((g1417) & (g1451) & (g2804) & (!g2845) & (!g2805) & (g2933)) + ((g1417) & (g1451) & (g2804) & (!g2845) & (g2805) & (g2933)) + ((g1417) & (g1451) & (g2804) & (g2845) & (!g2805) & (g2933)) + ((g1417) & (g1451) & (g2804) & (g2845) & (g2805) & (g2933)));
	assign g2935 = (((g1485) & (g2885)));
	assign g2936 = (((!g2934) & (!g2935)));
	assign g2937 = (((!g827) & (!g1518) & (g2932) & (!g2936)) + ((!g827) & (!g1518) & (g2932) & (g2936)) + ((!g827) & (g1518) & (g2932) & (!g2936)) + ((!g827) & (g1518) & (g2932) & (g2936)) + ((g827) & (!g1518) & (!g2932) & (!g2936)) + ((g827) & (!g1518) & (g2932) & (g2936)) + ((g827) & (g1518) & (!g2932) & (g2936)) + ((g827) & (g1518) & (g2932) & (!g2936)));
	assign g8157 = (((!g3464) & (g5166) & (!g2938)) + ((!g3464) & (g5166) & (g2938)) + ((g3464) & (!g5166) & (g2938)) + ((g3464) & (g5166) & (g2938)));
	assign g2939 = (((!g1493) & (g2893)) + ((g1493) & (!g2893)));
	assign g2940 = (((!g1425) & (!g1453) & (g2816) & (g2848) & (!g2817) & (g2939)) + ((!g1425) & (g1453) & (!g2816) & (g2848) & (!g2817) & (g2939)) + ((!g1425) & (g1453) & (!g2816) & (g2848) & (g2817) & (g2939)) + ((!g1425) & (g1453) & (g2816) & (!g2848) & (!g2817) & (g2939)) + ((!g1425) & (g1453) & (g2816) & (g2848) & (!g2817) & (g2939)) + ((!g1425) & (g1453) & (g2816) & (g2848) & (g2817) & (g2939)) + ((g1425) & (!g1453) & (!g2816) & (g2848) & (!g2817) & (g2939)) + ((g1425) & (!g1453) & (g2816) & (g2848) & (!g2817) & (g2939)) + ((g1425) & (!g1453) & (g2816) & (g2848) & (g2817) & (g2939)) + ((g1425) & (g1453) & (!g2816) & (!g2848) & (!g2817) & (g2939)) + ((g1425) & (g1453) & (!g2816) & (g2848) & (!g2817) & (g2939)) + ((g1425) & (g1453) & (!g2816) & (g2848) & (g2817) & (g2939)) + ((g1425) & (g1453) & (g2816) & (!g2848) & (!g2817) & (g2939)) + ((g1425) & (g1453) & (g2816) & (!g2848) & (g2817) & (g2939)) + ((g1425) & (g1453) & (g2816) & (g2848) & (!g2817) & (g2939)) + ((g1425) & (g1453) & (g2816) & (g2848) & (g2817) & (g2939)));
	assign g2941 = (((g1493) & (g2893)));
	assign g2942 = (((!g2940) & (!g2941)));
	assign g2943 = (((!g827) & (!g1520) & (g2938) & (!g2942)) + ((!g827) & (!g1520) & (g2938) & (g2942)) + ((!g827) & (g1520) & (g2938) & (!g2942)) + ((!g827) & (g1520) & (g2938) & (g2942)) + ((g827) & (!g1520) & (!g2938) & (!g2942)) + ((g827) & (!g1520) & (g2938) & (g2942)) + ((g827) & (g1520) & (!g2938) & (g2942)) + ((g827) & (g1520) & (g2938) & (!g2942)));
	assign g8158 = (((!g3499) & (g5170) & (!g2944)) + ((!g3499) & (g5170) & (g2944)) + ((g3499) & (!g5170) & (g2944)) + ((g3499) & (g5170) & (g2944)));
	assign g2945 = (((!g1501) & (g2900)) + ((g1501) & (!g2900)));
	assign g2946 = (((!g1433) & (!g1455) & (g2827) & (g2851) & (!g2828) & (g2945)) + ((!g1433) & (g1455) & (!g2827) & (g2851) & (!g2828) & (g2945)) + ((!g1433) & (g1455) & (!g2827) & (g2851) & (g2828) & (g2945)) + ((!g1433) & (g1455) & (g2827) & (!g2851) & (!g2828) & (g2945)) + ((!g1433) & (g1455) & (g2827) & (g2851) & (!g2828) & (g2945)) + ((!g1433) & (g1455) & (g2827) & (g2851) & (g2828) & (g2945)) + ((g1433) & (!g1455) & (!g2827) & (g2851) & (!g2828) & (g2945)) + ((g1433) & (!g1455) & (g2827) & (g2851) & (!g2828) & (g2945)) + ((g1433) & (!g1455) & (g2827) & (g2851) & (g2828) & (g2945)) + ((g1433) & (g1455) & (!g2827) & (!g2851) & (!g2828) & (g2945)) + ((g1433) & (g1455) & (!g2827) & (g2851) & (!g2828) & (g2945)) + ((g1433) & (g1455) & (!g2827) & (g2851) & (g2828) & (g2945)) + ((g1433) & (g1455) & (g2827) & (!g2851) & (!g2828) & (g2945)) + ((g1433) & (g1455) & (g2827) & (!g2851) & (g2828) & (g2945)) + ((g1433) & (g1455) & (g2827) & (g2851) & (!g2828) & (g2945)) + ((g1433) & (g1455) & (g2827) & (g2851) & (g2828) & (g2945)));
	assign g2947 = (((g1501) & (g2900)));
	assign g2948 = (((!g2946) & (!g2947)));
	assign g2949 = (((!g827) & (!g1522) & (g2944) & (!g2948)) + ((!g827) & (!g1522) & (g2944) & (g2948)) + ((!g827) & (g1522) & (g2944) & (!g2948)) + ((!g827) & (g1522) & (g2944) & (g2948)) + ((g827) & (!g1522) & (!g2944) & (!g2948)) + ((g827) & (!g1522) & (g2944) & (g2948)) + ((g827) & (g1522) & (!g2944) & (g2948)) + ((g827) & (g1522) & (g2944) & (!g2948)));
	assign g8159 = (((!g3464) & (g5174) & (!g2950)) + ((!g3464) & (g5174) & (g2950)) + ((g3464) & (!g5174) & (g2950)) + ((g3464) & (g5174) & (g2950)));
	assign g2951 = (((!g1479) & (g2881)) + ((g1479) & (!g2881)));
	assign g2952 = (((!g1411) & (!g1457) & (g2797) & (g2854) & (!g2798) & (g2951)) + ((!g1411) & (g1457) & (!g2797) & (g2854) & (!g2798) & (g2951)) + ((!g1411) & (g1457) & (!g2797) & (g2854) & (g2798) & (g2951)) + ((!g1411) & (g1457) & (g2797) & (!g2854) & (!g2798) & (g2951)) + ((!g1411) & (g1457) & (g2797) & (g2854) & (!g2798) & (g2951)) + ((!g1411) & (g1457) & (g2797) & (g2854) & (g2798) & (g2951)) + ((g1411) & (!g1457) & (!g2797) & (g2854) & (!g2798) & (g2951)) + ((g1411) & (!g1457) & (g2797) & (g2854) & (!g2798) & (g2951)) + ((g1411) & (!g1457) & (g2797) & (g2854) & (g2798) & (g2951)) + ((g1411) & (g1457) & (!g2797) & (!g2854) & (!g2798) & (g2951)) + ((g1411) & (g1457) & (!g2797) & (g2854) & (!g2798) & (g2951)) + ((g1411) & (g1457) & (!g2797) & (g2854) & (g2798) & (g2951)) + ((g1411) & (g1457) & (g2797) & (!g2854) & (!g2798) & (g2951)) + ((g1411) & (g1457) & (g2797) & (!g2854) & (g2798) & (g2951)) + ((g1411) & (g1457) & (g2797) & (g2854) & (!g2798) & (g2951)) + ((g1411) & (g1457) & (g2797) & (g2854) & (g2798) & (g2951)));
	assign g2953 = (((g1479) & (g2881)));
	assign g2954 = (((!g2952) & (!g2953)));
	assign g2955 = (((!g827) & (!g1524) & (g2950) & (!g2954)) + ((!g827) & (!g1524) & (g2950) & (g2954)) + ((!g827) & (g1524) & (g2950) & (!g2954)) + ((!g827) & (g1524) & (g2950) & (g2954)) + ((g827) & (!g1524) & (!g2950) & (!g2954)) + ((g827) & (!g1524) & (g2950) & (g2954)) + ((g827) & (g1524) & (!g2950) & (g2954)) + ((g827) & (g1524) & (g2950) & (!g2954)));
	assign g8160 = (((!g3499) & (g5178) & (!g2956)) + ((!g3499) & (g5178) & (g2956)) + ((g3499) & (!g5178) & (g2956)) + ((g3499) & (g5178) & (g2956)));
	assign g2957 = (((!g1487) & (g2887)) + ((g1487) & (!g2887)));
	assign g2958 = (((!g1419) & (!g1459) & (g2807) & (g2857) & (!g2808) & (g2957)) + ((!g1419) & (g1459) & (!g2807) & (g2857) & (!g2808) & (g2957)) + ((!g1419) & (g1459) & (!g2807) & (g2857) & (g2808) & (g2957)) + ((!g1419) & (g1459) & (g2807) & (!g2857) & (!g2808) & (g2957)) + ((!g1419) & (g1459) & (g2807) & (g2857) & (!g2808) & (g2957)) + ((!g1419) & (g1459) & (g2807) & (g2857) & (g2808) & (g2957)) + ((g1419) & (!g1459) & (!g2807) & (g2857) & (!g2808) & (g2957)) + ((g1419) & (!g1459) & (g2807) & (g2857) & (!g2808) & (g2957)) + ((g1419) & (!g1459) & (g2807) & (g2857) & (g2808) & (g2957)) + ((g1419) & (g1459) & (!g2807) & (!g2857) & (!g2808) & (g2957)) + ((g1419) & (g1459) & (!g2807) & (g2857) & (!g2808) & (g2957)) + ((g1419) & (g1459) & (!g2807) & (g2857) & (g2808) & (g2957)) + ((g1419) & (g1459) & (g2807) & (!g2857) & (!g2808) & (g2957)) + ((g1419) & (g1459) & (g2807) & (!g2857) & (g2808) & (g2957)) + ((g1419) & (g1459) & (g2807) & (g2857) & (!g2808) & (g2957)) + ((g1419) & (g1459) & (g2807) & (g2857) & (g2808) & (g2957)));
	assign g2959 = (((g1487) & (g2887)));
	assign g2960 = (((!g2958) & (!g2959)));
	assign g2961 = (((!g827) & (!g1526) & (g2956) & (!g2960)) + ((!g827) & (!g1526) & (g2956) & (g2960)) + ((!g827) & (g1526) & (g2956) & (!g2960)) + ((!g827) & (g1526) & (g2956) & (g2960)) + ((g827) & (!g1526) & (!g2956) & (!g2960)) + ((g827) & (!g1526) & (g2956) & (g2960)) + ((g827) & (g1526) & (!g2956) & (g2960)) + ((g827) & (g1526) & (g2956) & (!g2960)));
	assign g8161 = (((!g2017) & (g6167) & (!g2962)) + ((!g2017) & (g6167) & (g2962)) + ((g2017) & (!g6167) & (g2962)) + ((g2017) & (g6167) & (g2962)));
	assign g2963 = (((!g1495) & (g2895)) + ((g1495) & (!g2895)));
	assign g2964 = (((!g1427) & (!g1461) & (g2819) & (g2860) & (!g2820) & (g2963)) + ((!g1427) & (g1461) & (!g2819) & (g2860) & (!g2820) & (g2963)) + ((!g1427) & (g1461) & (!g2819) & (g2860) & (g2820) & (g2963)) + ((!g1427) & (g1461) & (g2819) & (!g2860) & (!g2820) & (g2963)) + ((!g1427) & (g1461) & (g2819) & (g2860) & (!g2820) & (g2963)) + ((!g1427) & (g1461) & (g2819) & (g2860) & (g2820) & (g2963)) + ((g1427) & (!g1461) & (!g2819) & (g2860) & (!g2820) & (g2963)) + ((g1427) & (!g1461) & (g2819) & (g2860) & (!g2820) & (g2963)) + ((g1427) & (!g1461) & (g2819) & (g2860) & (g2820) & (g2963)) + ((g1427) & (g1461) & (!g2819) & (!g2860) & (!g2820) & (g2963)) + ((g1427) & (g1461) & (!g2819) & (g2860) & (!g2820) & (g2963)) + ((g1427) & (g1461) & (!g2819) & (g2860) & (g2820) & (g2963)) + ((g1427) & (g1461) & (g2819) & (!g2860) & (!g2820) & (g2963)) + ((g1427) & (g1461) & (g2819) & (!g2860) & (g2820) & (g2963)) + ((g1427) & (g1461) & (g2819) & (g2860) & (!g2820) & (g2963)) + ((g1427) & (g1461) & (g2819) & (g2860) & (g2820) & (g2963)));
	assign g2965 = (((g1495) & (g2895)));
	assign g2966 = (((!g2964) & (!g2965)));
	assign g2967 = (((!g827) & (!g1528) & (g2962) & (!g2966)) + ((!g827) & (!g1528) & (g2962) & (g2966)) + ((!g827) & (g1528) & (g2962) & (!g2966)) + ((!g827) & (g1528) & (g2962) & (g2966)) + ((g827) & (!g1528) & (!g2962) & (!g2966)) + ((g827) & (!g1528) & (g2962) & (g2966)) + ((g827) & (g1528) & (!g2962) & (g2966)) + ((g827) & (g1528) & (g2962) & (!g2966)));
	assign g8162 = (((!g3429) & (g5182) & (!g2968)) + ((!g3429) & (g5182) & (g2968)) + ((g3429) & (!g5182) & (g2968)) + ((g3429) & (g5182) & (g2968)));
	assign g2969 = (((!g1503) & (g2902)) + ((g1503) & (!g2902)));
	assign g2970 = (((!g1435) & (!g1463) & (g2830) & (g2863) & (!g2831) & (g2969)) + ((!g1435) & (g1463) & (!g2830) & (g2863) & (!g2831) & (g2969)) + ((!g1435) & (g1463) & (!g2830) & (g2863) & (g2831) & (g2969)) + ((!g1435) & (g1463) & (g2830) & (!g2863) & (!g2831) & (g2969)) + ((!g1435) & (g1463) & (g2830) & (g2863) & (!g2831) & (g2969)) + ((!g1435) & (g1463) & (g2830) & (g2863) & (g2831) & (g2969)) + ((g1435) & (!g1463) & (!g2830) & (g2863) & (!g2831) & (g2969)) + ((g1435) & (!g1463) & (g2830) & (g2863) & (!g2831) & (g2969)) + ((g1435) & (!g1463) & (g2830) & (g2863) & (g2831) & (g2969)) + ((g1435) & (g1463) & (!g2830) & (!g2863) & (!g2831) & (g2969)) + ((g1435) & (g1463) & (!g2830) & (g2863) & (!g2831) & (g2969)) + ((g1435) & (g1463) & (!g2830) & (g2863) & (g2831) & (g2969)) + ((g1435) & (g1463) & (g2830) & (!g2863) & (!g2831) & (g2969)) + ((g1435) & (g1463) & (g2830) & (!g2863) & (g2831) & (g2969)) + ((g1435) & (g1463) & (g2830) & (g2863) & (!g2831) & (g2969)) + ((g1435) & (g1463) & (g2830) & (g2863) & (g2831) & (g2969)));
	assign g2971 = (((g1503) & (g2902)));
	assign g2972 = (((!g2970) & (!g2971)));
	assign g2973 = (((!g827) & (!g1530) & (g2968) & (!g2972)) + ((!g827) & (!g1530) & (g2968) & (g2972)) + ((!g827) & (g1530) & (g2968) & (!g2972)) + ((!g827) & (g1530) & (g2968) & (g2972)) + ((g827) & (!g1530) & (!g2968) & (!g2972)) + ((g827) & (!g1530) & (g2968) & (g2972)) + ((g827) & (g1530) & (!g2968) & (g2972)) + ((g827) & (g1530) & (g2968) & (!g2972)));
	assign g2974 = (((!g1481) & (g2263)) + ((g1481) & (!g2263)));
	assign g2975 = (((!g1413) & (!g1465) & (g2181) & (g2213) & (!g2800) & (g2974)) + ((!g1413) & (g1465) & (!g2181) & (g2213) & (!g2800) & (g2974)) + ((!g1413) & (g1465) & (!g2181) & (g2213) & (g2800) & (g2974)) + ((!g1413) & (g1465) & (g2181) & (!g2213) & (!g2800) & (g2974)) + ((!g1413) & (g1465) & (g2181) & (g2213) & (!g2800) & (g2974)) + ((!g1413) & (g1465) & (g2181) & (g2213) & (g2800) & (g2974)) + ((g1413) & (!g1465) & (!g2181) & (g2213) & (!g2800) & (g2974)) + ((g1413) & (!g1465) & (g2181) & (g2213) & (!g2800) & (g2974)) + ((g1413) & (!g1465) & (g2181) & (g2213) & (g2800) & (g2974)) + ((g1413) & (g1465) & (!g2181) & (!g2213) & (!g2800) & (g2974)) + ((g1413) & (g1465) & (!g2181) & (g2213) & (!g2800) & (g2974)) + ((g1413) & (g1465) & (!g2181) & (g2213) & (g2800) & (g2974)) + ((g1413) & (g1465) & (g2181) & (!g2213) & (!g2800) & (g2974)) + ((g1413) & (g1465) & (g2181) & (!g2213) & (g2800) & (g2974)) + ((g1413) & (g1465) & (g2181) & (g2213) & (!g2800) & (g2974)) + ((g1413) & (g1465) & (g2181) & (g2213) & (g2800) & (g2974)));
	assign g2976 = (((g1481) & (g2263)));
	assign g2977 = (((!g2975) & (!g2976)));
	assign g2978 = (((!g827) & (!g1532) & (g2299) & (!g2977)) + ((!g827) & (!g1532) & (g2299) & (g2977)) + ((!g827) & (g1532) & (g2299) & (!g2977)) + ((!g827) & (g1532) & (g2299) & (g2977)) + ((g827) & (!g1532) & (!g2299) & (!g2977)) + ((g827) & (!g1532) & (g2299) & (g2977)) + ((g827) & (g1532) & (!g2299) & (g2977)) + ((g827) & (g1532) & (g2299) & (!g2977)));
	assign g8163 = (((!g3464) & (g5186) & (!g2979)) + ((!g3464) & (g5186) & (g2979)) + ((g3464) & (!g5186) & (g2979)) + ((g3464) & (g5186) & (g2979)));
	assign g2980 = (((!g1489) & (g2889)) + ((g1489) & (!g2889)));
	assign g2981 = (((!g1421) & (!g1467) & (g2810) & (g2868) & (!g2811) & (g2980)) + ((!g1421) & (g1467) & (!g2810) & (g2868) & (!g2811) & (g2980)) + ((!g1421) & (g1467) & (!g2810) & (g2868) & (g2811) & (g2980)) + ((!g1421) & (g1467) & (g2810) & (!g2868) & (!g2811) & (g2980)) + ((!g1421) & (g1467) & (g2810) & (g2868) & (!g2811) & (g2980)) + ((!g1421) & (g1467) & (g2810) & (g2868) & (g2811) & (g2980)) + ((g1421) & (!g1467) & (!g2810) & (g2868) & (!g2811) & (g2980)) + ((g1421) & (!g1467) & (g2810) & (g2868) & (!g2811) & (g2980)) + ((g1421) & (!g1467) & (g2810) & (g2868) & (g2811) & (g2980)) + ((g1421) & (g1467) & (!g2810) & (!g2868) & (!g2811) & (g2980)) + ((g1421) & (g1467) & (!g2810) & (g2868) & (!g2811) & (g2980)) + ((g1421) & (g1467) & (!g2810) & (g2868) & (g2811) & (g2980)) + ((g1421) & (g1467) & (g2810) & (!g2868) & (!g2811) & (g2980)) + ((g1421) & (g1467) & (g2810) & (!g2868) & (g2811) & (g2980)) + ((g1421) & (g1467) & (g2810) & (g2868) & (!g2811) & (g2980)) + ((g1421) & (g1467) & (g2810) & (g2868) & (g2811) & (g2980)));
	assign g2982 = (((g1489) & (g2889)));
	assign g2983 = (((!g2981) & (!g2982)));
	assign g2984 = (((!g827) & (!g1534) & (g2979) & (!g2983)) + ((!g827) & (!g1534) & (g2979) & (g2983)) + ((!g827) & (g1534) & (g2979) & (!g2983)) + ((!g827) & (g1534) & (g2979) & (g2983)) + ((g827) & (!g1534) & (!g2979) & (!g2983)) + ((g827) & (!g1534) & (g2979) & (g2983)) + ((g827) & (g1534) & (!g2979) & (g2983)) + ((g827) & (g1534) & (g2979) & (!g2983)));
	assign g8164 = (((!g3429) & (g5189) & (!g2985)) + ((!g3429) & (g5189) & (g2985)) + ((g3429) & (!g5189) & (g2985)) + ((g3429) & (g5189) & (g2985)));
	assign g2986 = (((!g1497) & (g2897)) + ((g1497) & (!g2897)));
	assign g2987 = (((!g1429) & (!g1469) & (g2822) & (g2871) & (!g2823) & (g2986)) + ((!g1429) & (g1469) & (!g2822) & (g2871) & (!g2823) & (g2986)) + ((!g1429) & (g1469) & (!g2822) & (g2871) & (g2823) & (g2986)) + ((!g1429) & (g1469) & (g2822) & (!g2871) & (!g2823) & (g2986)) + ((!g1429) & (g1469) & (g2822) & (g2871) & (!g2823) & (g2986)) + ((!g1429) & (g1469) & (g2822) & (g2871) & (g2823) & (g2986)) + ((g1429) & (!g1469) & (!g2822) & (g2871) & (!g2823) & (g2986)) + ((g1429) & (!g1469) & (g2822) & (g2871) & (!g2823) & (g2986)) + ((g1429) & (!g1469) & (g2822) & (g2871) & (g2823) & (g2986)) + ((g1429) & (g1469) & (!g2822) & (!g2871) & (!g2823) & (g2986)) + ((g1429) & (g1469) & (!g2822) & (g2871) & (!g2823) & (g2986)) + ((g1429) & (g1469) & (!g2822) & (g2871) & (g2823) & (g2986)) + ((g1429) & (g1469) & (g2822) & (!g2871) & (!g2823) & (g2986)) + ((g1429) & (g1469) & (g2822) & (!g2871) & (g2823) & (g2986)) + ((g1429) & (g1469) & (g2822) & (g2871) & (!g2823) & (g2986)) + ((g1429) & (g1469) & (g2822) & (g2871) & (g2823) & (g2986)));
	assign g2988 = (((g1497) & (g2897)));
	assign g2989 = (((!g2987) & (!g2988)));
	assign g2990 = (((!g827) & (!g1536) & (g2985) & (!g2989)) + ((!g827) & (!g1536) & (g2985) & (g2989)) + ((!g827) & (g1536) & (g2985) & (!g2989)) + ((!g827) & (g1536) & (g2985) & (g2989)) + ((g827) & (!g1536) & (!g2985) & (!g2989)) + ((g827) & (!g1536) & (g2985) & (g2989)) + ((g827) & (g1536) & (!g2985) & (g2989)) + ((g827) & (g1536) & (g2985) & (!g2989)));
	assign g8165 = (((!g2017) & (g6160) & (!g2991)) + ((!g2017) & (g6160) & (g2991)) + ((g2017) & (!g6160) & (g2991)) + ((g2017) & (g6160) & (g2991)));
	assign g2992 = (((!g1505) & (g2904)) + ((g1505) & (!g2904)));
	assign g2993 = (((!g1437) & (!g1471) & (g2833) & (g2874) & (!g2834) & (g2992)) + ((!g1437) & (g1471) & (!g2833) & (g2874) & (!g2834) & (g2992)) + ((!g1437) & (g1471) & (!g2833) & (g2874) & (g2834) & (g2992)) + ((!g1437) & (g1471) & (g2833) & (!g2874) & (!g2834) & (g2992)) + ((!g1437) & (g1471) & (g2833) & (g2874) & (!g2834) & (g2992)) + ((!g1437) & (g1471) & (g2833) & (g2874) & (g2834) & (g2992)) + ((g1437) & (!g1471) & (!g2833) & (g2874) & (!g2834) & (g2992)) + ((g1437) & (!g1471) & (g2833) & (g2874) & (!g2834) & (g2992)) + ((g1437) & (!g1471) & (g2833) & (g2874) & (g2834) & (g2992)) + ((g1437) & (g1471) & (!g2833) & (!g2874) & (!g2834) & (g2992)) + ((g1437) & (g1471) & (!g2833) & (g2874) & (!g2834) & (g2992)) + ((g1437) & (g1471) & (!g2833) & (g2874) & (g2834) & (g2992)) + ((g1437) & (g1471) & (g2833) & (!g2874) & (!g2834) & (g2992)) + ((g1437) & (g1471) & (g2833) & (!g2874) & (g2834) & (g2992)) + ((g1437) & (g1471) & (g2833) & (g2874) & (!g2834) & (g2992)) + ((g1437) & (g1471) & (g2833) & (g2874) & (g2834) & (g2992)));
	assign g2994 = (((g1505) & (g2904)));
	assign g2995 = (((!g2993) & (!g2994)));
	assign g2996 = (((!g827) & (!g1538) & (g2991) & (!g2995)) + ((!g827) & (!g1538) & (g2991) & (g2995)) + ((!g827) & (g1538) & (g2991) & (!g2995)) + ((!g827) & (g1538) & (g2991) & (g2995)) + ((g827) & (!g1538) & (!g2991) & (!g2995)) + ((g827) & (!g1538) & (g2991) & (g2995)) + ((g827) & (g1538) & (!g2991) & (g2995)) + ((g827) & (g1538) & (g2991) & (!g2995)));
	assign g2997 = (((!g1981) & (!g1982) & (g1983)) + ((!g1981) & (g1982) & (!g1983)) + ((g1981) & (!g1982) & (!g1983)) + ((g1981) & (g1982) & (g1983)));
	assign g2998 = (((!g827) & (!g1516) & (!g1547) & (!g2298) & (g2347) & (!g2930)) + ((!g827) & (!g1516) & (!g1547) & (!g2298) & (g2347) & (g2930)) + ((!g827) & (!g1516) & (!g1547) & (g2298) & (g2347) & (!g2930)) + ((!g827) & (!g1516) & (!g1547) & (g2298) & (g2347) & (g2930)) + ((!g827) & (!g1516) & (g1547) & (!g2298) & (g2347) & (!g2930)) + ((!g827) & (!g1516) & (g1547) & (!g2298) & (g2347) & (g2930)) + ((!g827) & (!g1516) & (g1547) & (g2298) & (g2347) & (!g2930)) + ((!g827) & (!g1516) & (g1547) & (g2298) & (g2347) & (g2930)) + ((!g827) & (g1516) & (!g1547) & (!g2298) & (g2347) & (!g2930)) + ((!g827) & (g1516) & (!g1547) & (!g2298) & (g2347) & (g2930)) + ((!g827) & (g1516) & (!g1547) & (g2298) & (g2347) & (!g2930)) + ((!g827) & (g1516) & (!g1547) & (g2298) & (g2347) & (g2930)) + ((!g827) & (g1516) & (g1547) & (!g2298) & (g2347) & (!g2930)) + ((!g827) & (g1516) & (g1547) & (!g2298) & (g2347) & (g2930)) + ((!g827) & (g1516) & (g1547) & (g2298) & (g2347) & (!g2930)) + ((!g827) & (g1516) & (g1547) & (g2298) & (g2347) & (g2930)) + ((g827) & (!g1516) & (!g1547) & (!g2298) & (g2347) & (!g2930)) + ((g827) & (!g1516) & (!g1547) & (!g2298) & (g2347) & (g2930)) + ((g827) & (!g1516) & (!g1547) & (g2298) & (!g2347) & (!g2930)) + ((g827) & (!g1516) & (!g1547) & (g2298) & (g2347) & (g2930)) + ((g827) & (!g1516) & (g1547) & (!g2298) & (!g2347) & (!g2930)) + ((g827) & (!g1516) & (g1547) & (!g2298) & (!g2347) & (g2930)) + ((g827) & (!g1516) & (g1547) & (g2298) & (!g2347) & (g2930)) + ((g827) & (!g1516) & (g1547) & (g2298) & (g2347) & (!g2930)) + ((g827) & (g1516) & (!g1547) & (!g2298) & (!g2347) & (!g2930)) + ((g827) & (g1516) & (!g1547) & (!g2298) & (g2347) & (g2930)) + ((g827) & (g1516) & (!g1547) & (g2298) & (!g2347) & (!g2930)) + ((g827) & (g1516) & (!g1547) & (g2298) & (!g2347) & (g2930)) + ((g827) & (g1516) & (g1547) & (!g2298) & (!g2347) & (g2930)) + ((g827) & (g1516) & (g1547) & (!g2298) & (g2347) & (!g2930)) + ((g827) & (g1516) & (g1547) & (g2298) & (g2347) & (!g2930)) + ((g827) & (g1516) & (g1547) & (g2298) & (g2347) & (g2930)));
	assign g8166 = (((!g3464) & (g5193) & (!g2999)) + ((!g3464) & (g5193) & (g2999)) + ((g3464) & (!g5193) & (g2999)) + ((g3464) & (g5193) & (g2999)));
	assign g3000 = (((!g827) & (!g1524) & (!g1549) & (!g2950) & (g2999) & (!g2954)) + ((!g827) & (!g1524) & (!g1549) & (!g2950) & (g2999) & (g2954)) + ((!g827) & (!g1524) & (!g1549) & (g2950) & (g2999) & (!g2954)) + ((!g827) & (!g1524) & (!g1549) & (g2950) & (g2999) & (g2954)) + ((!g827) & (!g1524) & (g1549) & (!g2950) & (g2999) & (!g2954)) + ((!g827) & (!g1524) & (g1549) & (!g2950) & (g2999) & (g2954)) + ((!g827) & (!g1524) & (g1549) & (g2950) & (g2999) & (!g2954)) + ((!g827) & (!g1524) & (g1549) & (g2950) & (g2999) & (g2954)) + ((!g827) & (g1524) & (!g1549) & (!g2950) & (g2999) & (!g2954)) + ((!g827) & (g1524) & (!g1549) & (!g2950) & (g2999) & (g2954)) + ((!g827) & (g1524) & (!g1549) & (g2950) & (g2999) & (!g2954)) + ((!g827) & (g1524) & (!g1549) & (g2950) & (g2999) & (g2954)) + ((!g827) & (g1524) & (g1549) & (!g2950) & (g2999) & (!g2954)) + ((!g827) & (g1524) & (g1549) & (!g2950) & (g2999) & (g2954)) + ((!g827) & (g1524) & (g1549) & (g2950) & (g2999) & (!g2954)) + ((!g827) & (g1524) & (g1549) & (g2950) & (g2999) & (g2954)) + ((g827) & (!g1524) & (!g1549) & (!g2950) & (g2999) & (!g2954)) + ((g827) & (!g1524) & (!g1549) & (!g2950) & (g2999) & (g2954)) + ((g827) & (!g1524) & (!g1549) & (g2950) & (!g2999) & (!g2954)) + ((g827) & (!g1524) & (!g1549) & (g2950) & (g2999) & (g2954)) + ((g827) & (!g1524) & (g1549) & (!g2950) & (!g2999) & (!g2954)) + ((g827) & (!g1524) & (g1549) & (!g2950) & (!g2999) & (g2954)) + ((g827) & (!g1524) & (g1549) & (g2950) & (!g2999) & (g2954)) + ((g827) & (!g1524) & (g1549) & (g2950) & (g2999) & (!g2954)) + ((g827) & (g1524) & (!g1549) & (!g2950) & (!g2999) & (!g2954)) + ((g827) & (g1524) & (!g1549) & (!g2950) & (g2999) & (g2954)) + ((g827) & (g1524) & (!g1549) & (g2950) & (!g2999) & (!g2954)) + ((g827) & (g1524) & (!g1549) & (g2950) & (!g2999) & (g2954)) + ((g827) & (g1524) & (g1549) & (!g2950) & (!g2999) & (g2954)) + ((g827) & (g1524) & (g1549) & (!g2950) & (g2999) & (!g2954)) + ((g827) & (g1524) & (g1549) & (g2950) & (g2999) & (!g2954)) + ((g827) & (g1524) & (g1549) & (g2950) & (g2999) & (g2954)));
	assign g3001 = (((!g827) & (!g1532) & (!g1551) & (!g2299) & (g2348) & (!g2977)) + ((!g827) & (!g1532) & (!g1551) & (!g2299) & (g2348) & (g2977)) + ((!g827) & (!g1532) & (!g1551) & (g2299) & (g2348) & (!g2977)) + ((!g827) & (!g1532) & (!g1551) & (g2299) & (g2348) & (g2977)) + ((!g827) & (!g1532) & (g1551) & (!g2299) & (g2348) & (!g2977)) + ((!g827) & (!g1532) & (g1551) & (!g2299) & (g2348) & (g2977)) + ((!g827) & (!g1532) & (g1551) & (g2299) & (g2348) & (!g2977)) + ((!g827) & (!g1532) & (g1551) & (g2299) & (g2348) & (g2977)) + ((!g827) & (g1532) & (!g1551) & (!g2299) & (g2348) & (!g2977)) + ((!g827) & (g1532) & (!g1551) & (!g2299) & (g2348) & (g2977)) + ((!g827) & (g1532) & (!g1551) & (g2299) & (g2348) & (!g2977)) + ((!g827) & (g1532) & (!g1551) & (g2299) & (g2348) & (g2977)) + ((!g827) & (g1532) & (g1551) & (!g2299) & (g2348) & (!g2977)) + ((!g827) & (g1532) & (g1551) & (!g2299) & (g2348) & (g2977)) + ((!g827) & (g1532) & (g1551) & (g2299) & (g2348) & (!g2977)) + ((!g827) & (g1532) & (g1551) & (g2299) & (g2348) & (g2977)) + ((g827) & (!g1532) & (!g1551) & (!g2299) & (g2348) & (!g2977)) + ((g827) & (!g1532) & (!g1551) & (!g2299) & (g2348) & (g2977)) + ((g827) & (!g1532) & (!g1551) & (g2299) & (!g2348) & (!g2977)) + ((g827) & (!g1532) & (!g1551) & (g2299) & (g2348) & (g2977)) + ((g827) & (!g1532) & (g1551) & (!g2299) & (!g2348) & (!g2977)) + ((g827) & (!g1532) & (g1551) & (!g2299) & (!g2348) & (g2977)) + ((g827) & (!g1532) & (g1551) & (g2299) & (!g2348) & (g2977)) + ((g827) & (!g1532) & (g1551) & (g2299) & (g2348) & (!g2977)) + ((g827) & (g1532) & (!g1551) & (!g2299) & (!g2348) & (!g2977)) + ((g827) & (g1532) & (!g1551) & (!g2299) & (g2348) & (g2977)) + ((g827) & (g1532) & (!g1551) & (g2299) & (!g2348) & (!g2977)) + ((g827) & (g1532) & (!g1551) & (g2299) & (!g2348) & (g2977)) + ((g827) & (g1532) & (g1551) & (!g2299) & (!g2348) & (g2977)) + ((g827) & (g1532) & (g1551) & (!g2299) & (g2348) & (!g2977)) + ((g827) & (g1532) & (g1551) & (g2299) & (g2348) & (!g2977)) + ((g827) & (g1532) & (g1551) & (g2299) & (g2348) & (g2977)));
	assign g3002 = (((!g827) & (!g1510) & (!g1553) & (!g2295) & (g2343) & (!g2914)) + ((!g827) & (!g1510) & (!g1553) & (!g2295) & (g2343) & (g2914)) + ((!g827) & (!g1510) & (!g1553) & (g2295) & (g2343) & (!g2914)) + ((!g827) & (!g1510) & (!g1553) & (g2295) & (g2343) & (g2914)) + ((!g827) & (!g1510) & (g1553) & (!g2295) & (g2343) & (!g2914)) + ((!g827) & (!g1510) & (g1553) & (!g2295) & (g2343) & (g2914)) + ((!g827) & (!g1510) & (g1553) & (g2295) & (g2343) & (!g2914)) + ((!g827) & (!g1510) & (g1553) & (g2295) & (g2343) & (g2914)) + ((!g827) & (g1510) & (!g1553) & (!g2295) & (g2343) & (!g2914)) + ((!g827) & (g1510) & (!g1553) & (!g2295) & (g2343) & (g2914)) + ((!g827) & (g1510) & (!g1553) & (g2295) & (g2343) & (!g2914)) + ((!g827) & (g1510) & (!g1553) & (g2295) & (g2343) & (g2914)) + ((!g827) & (g1510) & (g1553) & (!g2295) & (g2343) & (!g2914)) + ((!g827) & (g1510) & (g1553) & (!g2295) & (g2343) & (g2914)) + ((!g827) & (g1510) & (g1553) & (g2295) & (g2343) & (!g2914)) + ((!g827) & (g1510) & (g1553) & (g2295) & (g2343) & (g2914)) + ((g827) & (!g1510) & (!g1553) & (!g2295) & (g2343) & (!g2914)) + ((g827) & (!g1510) & (!g1553) & (!g2295) & (g2343) & (g2914)) + ((g827) & (!g1510) & (!g1553) & (g2295) & (!g2343) & (!g2914)) + ((g827) & (!g1510) & (!g1553) & (g2295) & (g2343) & (g2914)) + ((g827) & (!g1510) & (g1553) & (!g2295) & (!g2343) & (!g2914)) + ((g827) & (!g1510) & (g1553) & (!g2295) & (!g2343) & (g2914)) + ((g827) & (!g1510) & (g1553) & (g2295) & (!g2343) & (g2914)) + ((g827) & (!g1510) & (g1553) & (g2295) & (g2343) & (!g2914)) + ((g827) & (g1510) & (!g1553) & (!g2295) & (!g2343) & (!g2914)) + ((g827) & (g1510) & (!g1553) & (!g2295) & (g2343) & (g2914)) + ((g827) & (g1510) & (!g1553) & (g2295) & (!g2343) & (!g2914)) + ((g827) & (g1510) & (!g1553) & (g2295) & (!g2343) & (g2914)) + ((g827) & (g1510) & (g1553) & (!g2295) & (!g2343) & (g2914)) + ((g827) & (g1510) & (g1553) & (!g2295) & (g2343) & (!g2914)) + ((g827) & (g1510) & (g1553) & (g2295) & (g2343) & (!g2914)) + ((g827) & (g1510) & (g1553) & (g2295) & (g2343) & (g2914)));
	assign g8167 = (((!g2017) & (g5198) & (!g3003)) + ((!g2017) & (g5198) & (g3003)) + ((g2017) & (!g5198) & (g3003)) + ((g2017) & (g5198) & (g3003)));
	assign g3004 = (((!g827) & (!g1518) & (!g1555) & (!g2932) & (g3003) & (!g2936)) + ((!g827) & (!g1518) & (!g1555) & (!g2932) & (g3003) & (g2936)) + ((!g827) & (!g1518) & (!g1555) & (g2932) & (g3003) & (!g2936)) + ((!g827) & (!g1518) & (!g1555) & (g2932) & (g3003) & (g2936)) + ((!g827) & (!g1518) & (g1555) & (!g2932) & (g3003) & (!g2936)) + ((!g827) & (!g1518) & (g1555) & (!g2932) & (g3003) & (g2936)) + ((!g827) & (!g1518) & (g1555) & (g2932) & (g3003) & (!g2936)) + ((!g827) & (!g1518) & (g1555) & (g2932) & (g3003) & (g2936)) + ((!g827) & (g1518) & (!g1555) & (!g2932) & (g3003) & (!g2936)) + ((!g827) & (g1518) & (!g1555) & (!g2932) & (g3003) & (g2936)) + ((!g827) & (g1518) & (!g1555) & (g2932) & (g3003) & (!g2936)) + ((!g827) & (g1518) & (!g1555) & (g2932) & (g3003) & (g2936)) + ((!g827) & (g1518) & (g1555) & (!g2932) & (g3003) & (!g2936)) + ((!g827) & (g1518) & (g1555) & (!g2932) & (g3003) & (g2936)) + ((!g827) & (g1518) & (g1555) & (g2932) & (g3003) & (!g2936)) + ((!g827) & (g1518) & (g1555) & (g2932) & (g3003) & (g2936)) + ((g827) & (!g1518) & (!g1555) & (!g2932) & (g3003) & (!g2936)) + ((g827) & (!g1518) & (!g1555) & (!g2932) & (g3003) & (g2936)) + ((g827) & (!g1518) & (!g1555) & (g2932) & (!g3003) & (!g2936)) + ((g827) & (!g1518) & (!g1555) & (g2932) & (g3003) & (g2936)) + ((g827) & (!g1518) & (g1555) & (!g2932) & (!g3003) & (!g2936)) + ((g827) & (!g1518) & (g1555) & (!g2932) & (!g3003) & (g2936)) + ((g827) & (!g1518) & (g1555) & (g2932) & (!g3003) & (g2936)) + ((g827) & (!g1518) & (g1555) & (g2932) & (g3003) & (!g2936)) + ((g827) & (g1518) & (!g1555) & (!g2932) & (!g3003) & (!g2936)) + ((g827) & (g1518) & (!g1555) & (!g2932) & (g3003) & (g2936)) + ((g827) & (g1518) & (!g1555) & (g2932) & (!g3003) & (!g2936)) + ((g827) & (g1518) & (!g1555) & (g2932) & (!g3003) & (g2936)) + ((g827) & (g1518) & (g1555) & (!g2932) & (!g3003) & (g2936)) + ((g827) & (g1518) & (g1555) & (!g2932) & (g3003) & (!g2936)) + ((g827) & (g1518) & (g1555) & (g2932) & (g3003) & (!g2936)) + ((g827) & (g1518) & (g1555) & (g2932) & (g3003) & (g2936)));
	assign g8168 = (((!g3499) & (g5201) & (!g3005)) + ((!g3499) & (g5201) & (g3005)) + ((g3499) & (!g5201) & (g3005)) + ((g3499) & (g5201) & (g3005)));
	assign g3006 = (((!g827) & (!g1526) & (!g1557) & (!g2956) & (g3005) & (!g2960)) + ((!g827) & (!g1526) & (!g1557) & (!g2956) & (g3005) & (g2960)) + ((!g827) & (!g1526) & (!g1557) & (g2956) & (g3005) & (!g2960)) + ((!g827) & (!g1526) & (!g1557) & (g2956) & (g3005) & (g2960)) + ((!g827) & (!g1526) & (g1557) & (!g2956) & (g3005) & (!g2960)) + ((!g827) & (!g1526) & (g1557) & (!g2956) & (g3005) & (g2960)) + ((!g827) & (!g1526) & (g1557) & (g2956) & (g3005) & (!g2960)) + ((!g827) & (!g1526) & (g1557) & (g2956) & (g3005) & (g2960)) + ((!g827) & (g1526) & (!g1557) & (!g2956) & (g3005) & (!g2960)) + ((!g827) & (g1526) & (!g1557) & (!g2956) & (g3005) & (g2960)) + ((!g827) & (g1526) & (!g1557) & (g2956) & (g3005) & (!g2960)) + ((!g827) & (g1526) & (!g1557) & (g2956) & (g3005) & (g2960)) + ((!g827) & (g1526) & (g1557) & (!g2956) & (g3005) & (!g2960)) + ((!g827) & (g1526) & (g1557) & (!g2956) & (g3005) & (g2960)) + ((!g827) & (g1526) & (g1557) & (g2956) & (g3005) & (!g2960)) + ((!g827) & (g1526) & (g1557) & (g2956) & (g3005) & (g2960)) + ((g827) & (!g1526) & (!g1557) & (!g2956) & (g3005) & (!g2960)) + ((g827) & (!g1526) & (!g1557) & (!g2956) & (g3005) & (g2960)) + ((g827) & (!g1526) & (!g1557) & (g2956) & (!g3005) & (!g2960)) + ((g827) & (!g1526) & (!g1557) & (g2956) & (g3005) & (g2960)) + ((g827) & (!g1526) & (g1557) & (!g2956) & (!g3005) & (!g2960)) + ((g827) & (!g1526) & (g1557) & (!g2956) & (!g3005) & (g2960)) + ((g827) & (!g1526) & (g1557) & (g2956) & (!g3005) & (g2960)) + ((g827) & (!g1526) & (g1557) & (g2956) & (g3005) & (!g2960)) + ((g827) & (g1526) & (!g1557) & (!g2956) & (!g3005) & (!g2960)) + ((g827) & (g1526) & (!g1557) & (!g2956) & (g3005) & (g2960)) + ((g827) & (g1526) & (!g1557) & (g2956) & (!g3005) & (!g2960)) + ((g827) & (g1526) & (!g1557) & (g2956) & (!g3005) & (g2960)) + ((g827) & (g1526) & (g1557) & (!g2956) & (!g3005) & (g2960)) + ((g827) & (g1526) & (g1557) & (!g2956) & (g3005) & (!g2960)) + ((g827) & (g1526) & (g1557) & (g2956) & (g3005) & (!g2960)) + ((g827) & (g1526) & (g1557) & (g2956) & (g3005) & (g2960)));
	assign g8169 = (((!g3464) & (g5204) & (!g3007)) + ((!g3464) & (g5204) & (g3007)) + ((g3464) & (!g5204) & (g3007)) + ((g3464) & (g5204) & (g3007)));
	assign g3008 = (((!g827) & (!g1534) & (!g1559) & (!g2979) & (g3007) & (!g2983)) + ((!g827) & (!g1534) & (!g1559) & (!g2979) & (g3007) & (g2983)) + ((!g827) & (!g1534) & (!g1559) & (g2979) & (g3007) & (!g2983)) + ((!g827) & (!g1534) & (!g1559) & (g2979) & (g3007) & (g2983)) + ((!g827) & (!g1534) & (g1559) & (!g2979) & (g3007) & (!g2983)) + ((!g827) & (!g1534) & (g1559) & (!g2979) & (g3007) & (g2983)) + ((!g827) & (!g1534) & (g1559) & (g2979) & (g3007) & (!g2983)) + ((!g827) & (!g1534) & (g1559) & (g2979) & (g3007) & (g2983)) + ((!g827) & (g1534) & (!g1559) & (!g2979) & (g3007) & (!g2983)) + ((!g827) & (g1534) & (!g1559) & (!g2979) & (g3007) & (g2983)) + ((!g827) & (g1534) & (!g1559) & (g2979) & (g3007) & (!g2983)) + ((!g827) & (g1534) & (!g1559) & (g2979) & (g3007) & (g2983)) + ((!g827) & (g1534) & (g1559) & (!g2979) & (g3007) & (!g2983)) + ((!g827) & (g1534) & (g1559) & (!g2979) & (g3007) & (g2983)) + ((!g827) & (g1534) & (g1559) & (g2979) & (g3007) & (!g2983)) + ((!g827) & (g1534) & (g1559) & (g2979) & (g3007) & (g2983)) + ((g827) & (!g1534) & (!g1559) & (!g2979) & (g3007) & (!g2983)) + ((g827) & (!g1534) & (!g1559) & (!g2979) & (g3007) & (g2983)) + ((g827) & (!g1534) & (!g1559) & (g2979) & (!g3007) & (!g2983)) + ((g827) & (!g1534) & (!g1559) & (g2979) & (g3007) & (g2983)) + ((g827) & (!g1534) & (g1559) & (!g2979) & (!g3007) & (!g2983)) + ((g827) & (!g1534) & (g1559) & (!g2979) & (!g3007) & (g2983)) + ((g827) & (!g1534) & (g1559) & (g2979) & (!g3007) & (g2983)) + ((g827) & (!g1534) & (g1559) & (g2979) & (g3007) & (!g2983)) + ((g827) & (g1534) & (!g1559) & (!g2979) & (!g3007) & (!g2983)) + ((g827) & (g1534) & (!g1559) & (!g2979) & (g3007) & (g2983)) + ((g827) & (g1534) & (!g1559) & (g2979) & (!g3007) & (!g2983)) + ((g827) & (g1534) & (!g1559) & (g2979) & (!g3007) & (g2983)) + ((g827) & (g1534) & (g1559) & (!g2979) & (!g3007) & (g2983)) + ((g827) & (g1534) & (g1559) & (!g2979) & (g3007) & (!g2983)) + ((g827) & (g1534) & (g1559) & (g2979) & (g3007) & (!g2983)) + ((g827) & (g1534) & (g1559) & (g2979) & (g3007) & (g2983)));
	assign g8170 = (((!g3499) & (g5207) & (!g3009)) + ((!g3499) & (g5207) & (g3009)) + ((g3499) & (!g5207) & (g3009)) + ((g3499) & (g5207) & (g3009)));
	assign g3010 = (((!g827) & (!g1512) & (!g1561) & (!g2916) & (g3009) & (!g2920)) + ((!g827) & (!g1512) & (!g1561) & (!g2916) & (g3009) & (g2920)) + ((!g827) & (!g1512) & (!g1561) & (g2916) & (g3009) & (!g2920)) + ((!g827) & (!g1512) & (!g1561) & (g2916) & (g3009) & (g2920)) + ((!g827) & (!g1512) & (g1561) & (!g2916) & (g3009) & (!g2920)) + ((!g827) & (!g1512) & (g1561) & (!g2916) & (g3009) & (g2920)) + ((!g827) & (!g1512) & (g1561) & (g2916) & (g3009) & (!g2920)) + ((!g827) & (!g1512) & (g1561) & (g2916) & (g3009) & (g2920)) + ((!g827) & (g1512) & (!g1561) & (!g2916) & (g3009) & (!g2920)) + ((!g827) & (g1512) & (!g1561) & (!g2916) & (g3009) & (g2920)) + ((!g827) & (g1512) & (!g1561) & (g2916) & (g3009) & (!g2920)) + ((!g827) & (g1512) & (!g1561) & (g2916) & (g3009) & (g2920)) + ((!g827) & (g1512) & (g1561) & (!g2916) & (g3009) & (!g2920)) + ((!g827) & (g1512) & (g1561) & (!g2916) & (g3009) & (g2920)) + ((!g827) & (g1512) & (g1561) & (g2916) & (g3009) & (!g2920)) + ((!g827) & (g1512) & (g1561) & (g2916) & (g3009) & (g2920)) + ((g827) & (!g1512) & (!g1561) & (!g2916) & (g3009) & (!g2920)) + ((g827) & (!g1512) & (!g1561) & (!g2916) & (g3009) & (g2920)) + ((g827) & (!g1512) & (!g1561) & (g2916) & (!g3009) & (!g2920)) + ((g827) & (!g1512) & (!g1561) & (g2916) & (g3009) & (g2920)) + ((g827) & (!g1512) & (g1561) & (!g2916) & (!g3009) & (!g2920)) + ((g827) & (!g1512) & (g1561) & (!g2916) & (!g3009) & (g2920)) + ((g827) & (!g1512) & (g1561) & (g2916) & (!g3009) & (g2920)) + ((g827) & (!g1512) & (g1561) & (g2916) & (g3009) & (!g2920)) + ((g827) & (g1512) & (!g1561) & (!g2916) & (!g3009) & (!g2920)) + ((g827) & (g1512) & (!g1561) & (!g2916) & (g3009) & (g2920)) + ((g827) & (g1512) & (!g1561) & (g2916) & (!g3009) & (!g2920)) + ((g827) & (g1512) & (!g1561) & (g2916) & (!g3009) & (g2920)) + ((g827) & (g1512) & (g1561) & (!g2916) & (!g3009) & (g2920)) + ((g827) & (g1512) & (g1561) & (!g2916) & (g3009) & (!g2920)) + ((g827) & (g1512) & (g1561) & (g2916) & (g3009) & (!g2920)) + ((g827) & (g1512) & (g1561) & (g2916) & (g3009) & (g2920)));
	assign g8171 = (((!g3464) & (g5211) & (!g3011)) + ((!g3464) & (g5211) & (g3011)) + ((g3464) & (!g5211) & (g3011)) + ((g3464) & (g5211) & (g3011)));
	assign g3012 = (((!g827) & (!g1520) & (!g1563) & (!g2938) & (g3011) & (!g2942)) + ((!g827) & (!g1520) & (!g1563) & (!g2938) & (g3011) & (g2942)) + ((!g827) & (!g1520) & (!g1563) & (g2938) & (g3011) & (!g2942)) + ((!g827) & (!g1520) & (!g1563) & (g2938) & (g3011) & (g2942)) + ((!g827) & (!g1520) & (g1563) & (!g2938) & (g3011) & (!g2942)) + ((!g827) & (!g1520) & (g1563) & (!g2938) & (g3011) & (g2942)) + ((!g827) & (!g1520) & (g1563) & (g2938) & (g3011) & (!g2942)) + ((!g827) & (!g1520) & (g1563) & (g2938) & (g3011) & (g2942)) + ((!g827) & (g1520) & (!g1563) & (!g2938) & (g3011) & (!g2942)) + ((!g827) & (g1520) & (!g1563) & (!g2938) & (g3011) & (g2942)) + ((!g827) & (g1520) & (!g1563) & (g2938) & (g3011) & (!g2942)) + ((!g827) & (g1520) & (!g1563) & (g2938) & (g3011) & (g2942)) + ((!g827) & (g1520) & (g1563) & (!g2938) & (g3011) & (!g2942)) + ((!g827) & (g1520) & (g1563) & (!g2938) & (g3011) & (g2942)) + ((!g827) & (g1520) & (g1563) & (g2938) & (g3011) & (!g2942)) + ((!g827) & (g1520) & (g1563) & (g2938) & (g3011) & (g2942)) + ((g827) & (!g1520) & (!g1563) & (!g2938) & (g3011) & (!g2942)) + ((g827) & (!g1520) & (!g1563) & (!g2938) & (g3011) & (g2942)) + ((g827) & (!g1520) & (!g1563) & (g2938) & (!g3011) & (!g2942)) + ((g827) & (!g1520) & (!g1563) & (g2938) & (g3011) & (g2942)) + ((g827) & (!g1520) & (g1563) & (!g2938) & (!g3011) & (!g2942)) + ((g827) & (!g1520) & (g1563) & (!g2938) & (!g3011) & (g2942)) + ((g827) & (!g1520) & (g1563) & (g2938) & (!g3011) & (g2942)) + ((g827) & (!g1520) & (g1563) & (g2938) & (g3011) & (!g2942)) + ((g827) & (g1520) & (!g1563) & (!g2938) & (!g3011) & (!g2942)) + ((g827) & (g1520) & (!g1563) & (!g2938) & (g3011) & (g2942)) + ((g827) & (g1520) & (!g1563) & (g2938) & (!g3011) & (!g2942)) + ((g827) & (g1520) & (!g1563) & (g2938) & (!g3011) & (g2942)) + ((g827) & (g1520) & (g1563) & (!g2938) & (!g3011) & (g2942)) + ((g827) & (g1520) & (g1563) & (!g2938) & (g3011) & (!g2942)) + ((g827) & (g1520) & (g1563) & (g2938) & (g3011) & (!g2942)) + ((g827) & (g1520) & (g1563) & (g2938) & (g3011) & (g2942)));
	assign g8172 = (((!g2017) & (g5216) & (!g3013)) + ((!g2017) & (g5216) & (g3013)) + ((g2017) & (!g5216) & (g3013)) + ((g2017) & (g5216) & (g3013)));
	assign g3014 = (((!g827) & (!g1528) & (!g1565) & (!g2962) & (g3013) & (!g2966)) + ((!g827) & (!g1528) & (!g1565) & (!g2962) & (g3013) & (g2966)) + ((!g827) & (!g1528) & (!g1565) & (g2962) & (g3013) & (!g2966)) + ((!g827) & (!g1528) & (!g1565) & (g2962) & (g3013) & (g2966)) + ((!g827) & (!g1528) & (g1565) & (!g2962) & (g3013) & (!g2966)) + ((!g827) & (!g1528) & (g1565) & (!g2962) & (g3013) & (g2966)) + ((!g827) & (!g1528) & (g1565) & (g2962) & (g3013) & (!g2966)) + ((!g827) & (!g1528) & (g1565) & (g2962) & (g3013) & (g2966)) + ((!g827) & (g1528) & (!g1565) & (!g2962) & (g3013) & (!g2966)) + ((!g827) & (g1528) & (!g1565) & (!g2962) & (g3013) & (g2966)) + ((!g827) & (g1528) & (!g1565) & (g2962) & (g3013) & (!g2966)) + ((!g827) & (g1528) & (!g1565) & (g2962) & (g3013) & (g2966)) + ((!g827) & (g1528) & (g1565) & (!g2962) & (g3013) & (!g2966)) + ((!g827) & (g1528) & (g1565) & (!g2962) & (g3013) & (g2966)) + ((!g827) & (g1528) & (g1565) & (g2962) & (g3013) & (!g2966)) + ((!g827) & (g1528) & (g1565) & (g2962) & (g3013) & (g2966)) + ((g827) & (!g1528) & (!g1565) & (!g2962) & (g3013) & (!g2966)) + ((g827) & (!g1528) & (!g1565) & (!g2962) & (g3013) & (g2966)) + ((g827) & (!g1528) & (!g1565) & (g2962) & (!g3013) & (!g2966)) + ((g827) & (!g1528) & (!g1565) & (g2962) & (g3013) & (g2966)) + ((g827) & (!g1528) & (g1565) & (!g2962) & (!g3013) & (!g2966)) + ((g827) & (!g1528) & (g1565) & (!g2962) & (!g3013) & (g2966)) + ((g827) & (!g1528) & (g1565) & (g2962) & (!g3013) & (g2966)) + ((g827) & (!g1528) & (g1565) & (g2962) & (g3013) & (!g2966)) + ((g827) & (g1528) & (!g1565) & (!g2962) & (!g3013) & (!g2966)) + ((g827) & (g1528) & (!g1565) & (!g2962) & (g3013) & (g2966)) + ((g827) & (g1528) & (!g1565) & (g2962) & (!g3013) & (!g2966)) + ((g827) & (g1528) & (!g1565) & (g2962) & (!g3013) & (g2966)) + ((g827) & (g1528) & (g1565) & (!g2962) & (!g3013) & (g2966)) + ((g827) & (g1528) & (g1565) & (!g2962) & (g3013) & (!g2966)) + ((g827) & (g1528) & (g1565) & (g2962) & (g3013) & (!g2966)) + ((g827) & (g1528) & (g1565) & (g2962) & (g3013) & (g2966)));
	assign g8173 = (((!g3429) & (g5219) & (!g3015)) + ((!g3429) & (g5219) & (g3015)) + ((g3429) & (!g5219) & (g3015)) + ((g3429) & (g5219) & (g3015)));
	assign g3016 = (((!g827) & (!g1536) & (!g1567) & (!g2985) & (g3015) & (!g2989)) + ((!g827) & (!g1536) & (!g1567) & (!g2985) & (g3015) & (g2989)) + ((!g827) & (!g1536) & (!g1567) & (g2985) & (g3015) & (!g2989)) + ((!g827) & (!g1536) & (!g1567) & (g2985) & (g3015) & (g2989)) + ((!g827) & (!g1536) & (g1567) & (!g2985) & (g3015) & (!g2989)) + ((!g827) & (!g1536) & (g1567) & (!g2985) & (g3015) & (g2989)) + ((!g827) & (!g1536) & (g1567) & (g2985) & (g3015) & (!g2989)) + ((!g827) & (!g1536) & (g1567) & (g2985) & (g3015) & (g2989)) + ((!g827) & (g1536) & (!g1567) & (!g2985) & (g3015) & (!g2989)) + ((!g827) & (g1536) & (!g1567) & (!g2985) & (g3015) & (g2989)) + ((!g827) & (g1536) & (!g1567) & (g2985) & (g3015) & (!g2989)) + ((!g827) & (g1536) & (!g1567) & (g2985) & (g3015) & (g2989)) + ((!g827) & (g1536) & (g1567) & (!g2985) & (g3015) & (!g2989)) + ((!g827) & (g1536) & (g1567) & (!g2985) & (g3015) & (g2989)) + ((!g827) & (g1536) & (g1567) & (g2985) & (g3015) & (!g2989)) + ((!g827) & (g1536) & (g1567) & (g2985) & (g3015) & (g2989)) + ((g827) & (!g1536) & (!g1567) & (!g2985) & (g3015) & (!g2989)) + ((g827) & (!g1536) & (!g1567) & (!g2985) & (g3015) & (g2989)) + ((g827) & (!g1536) & (!g1567) & (g2985) & (!g3015) & (!g2989)) + ((g827) & (!g1536) & (!g1567) & (g2985) & (g3015) & (g2989)) + ((g827) & (!g1536) & (g1567) & (!g2985) & (!g3015) & (!g2989)) + ((g827) & (!g1536) & (g1567) & (!g2985) & (!g3015) & (g2989)) + ((g827) & (!g1536) & (g1567) & (g2985) & (!g3015) & (g2989)) + ((g827) & (!g1536) & (g1567) & (g2985) & (g3015) & (!g2989)) + ((g827) & (g1536) & (!g1567) & (!g2985) & (!g3015) & (!g2989)) + ((g827) & (g1536) & (!g1567) & (!g2985) & (g3015) & (g2989)) + ((g827) & (g1536) & (!g1567) & (g2985) & (!g3015) & (!g2989)) + ((g827) & (g1536) & (!g1567) & (g2985) & (!g3015) & (g2989)) + ((g827) & (g1536) & (g1567) & (!g2985) & (!g3015) & (g2989)) + ((g827) & (g1536) & (g1567) & (!g2985) & (g3015) & (!g2989)) + ((g827) & (g1536) & (g1567) & (g2985) & (g3015) & (!g2989)) + ((g827) & (g1536) & (g1567) & (g2985) & (g3015) & (g2989)));
	assign g3017 = (((!g827) & (!g1514) & (!g1569) & (!g2296) & (g2344) & (!g2925)) + ((!g827) & (!g1514) & (!g1569) & (!g2296) & (g2344) & (g2925)) + ((!g827) & (!g1514) & (!g1569) & (g2296) & (g2344) & (!g2925)) + ((!g827) & (!g1514) & (!g1569) & (g2296) & (g2344) & (g2925)) + ((!g827) & (!g1514) & (g1569) & (!g2296) & (g2344) & (!g2925)) + ((!g827) & (!g1514) & (g1569) & (!g2296) & (g2344) & (g2925)) + ((!g827) & (!g1514) & (g1569) & (g2296) & (g2344) & (!g2925)) + ((!g827) & (!g1514) & (g1569) & (g2296) & (g2344) & (g2925)) + ((!g827) & (g1514) & (!g1569) & (!g2296) & (g2344) & (!g2925)) + ((!g827) & (g1514) & (!g1569) & (!g2296) & (g2344) & (g2925)) + ((!g827) & (g1514) & (!g1569) & (g2296) & (g2344) & (!g2925)) + ((!g827) & (g1514) & (!g1569) & (g2296) & (g2344) & (g2925)) + ((!g827) & (g1514) & (g1569) & (!g2296) & (g2344) & (!g2925)) + ((!g827) & (g1514) & (g1569) & (!g2296) & (g2344) & (g2925)) + ((!g827) & (g1514) & (g1569) & (g2296) & (g2344) & (!g2925)) + ((!g827) & (g1514) & (g1569) & (g2296) & (g2344) & (g2925)) + ((g827) & (!g1514) & (!g1569) & (!g2296) & (g2344) & (!g2925)) + ((g827) & (!g1514) & (!g1569) & (!g2296) & (g2344) & (g2925)) + ((g827) & (!g1514) & (!g1569) & (g2296) & (!g2344) & (!g2925)) + ((g827) & (!g1514) & (!g1569) & (g2296) & (g2344) & (g2925)) + ((g827) & (!g1514) & (g1569) & (!g2296) & (!g2344) & (!g2925)) + ((g827) & (!g1514) & (g1569) & (!g2296) & (!g2344) & (g2925)) + ((g827) & (!g1514) & (g1569) & (g2296) & (!g2344) & (g2925)) + ((g827) & (!g1514) & (g1569) & (g2296) & (g2344) & (!g2925)) + ((g827) & (g1514) & (!g1569) & (!g2296) & (!g2344) & (!g2925)) + ((g827) & (g1514) & (!g1569) & (!g2296) & (g2344) & (g2925)) + ((g827) & (g1514) & (!g1569) & (g2296) & (!g2344) & (!g2925)) + ((g827) & (g1514) & (!g1569) & (g2296) & (!g2344) & (g2925)) + ((g827) & (g1514) & (g1569) & (!g2296) & (!g2344) & (g2925)) + ((g827) & (g1514) & (g1569) & (!g2296) & (g2344) & (!g2925)) + ((g827) & (g1514) & (g1569) & (g2296) & (g2344) & (!g2925)) + ((g827) & (g1514) & (g1569) & (g2296) & (g2344) & (g2925)));
	assign g8174 = (((!g3499) & (g5222) & (!g3018)) + ((!g3499) & (g5222) & (g3018)) + ((g3499) & (!g5222) & (g3018)) + ((g3499) & (g5222) & (g3018)));
	assign g3019 = (((!g827) & (!g1522) & (!g1571) & (!g2944) & (g3018) & (!g2948)) + ((!g827) & (!g1522) & (!g1571) & (!g2944) & (g3018) & (g2948)) + ((!g827) & (!g1522) & (!g1571) & (g2944) & (g3018) & (!g2948)) + ((!g827) & (!g1522) & (!g1571) & (g2944) & (g3018) & (g2948)) + ((!g827) & (!g1522) & (g1571) & (!g2944) & (g3018) & (!g2948)) + ((!g827) & (!g1522) & (g1571) & (!g2944) & (g3018) & (g2948)) + ((!g827) & (!g1522) & (g1571) & (g2944) & (g3018) & (!g2948)) + ((!g827) & (!g1522) & (g1571) & (g2944) & (g3018) & (g2948)) + ((!g827) & (g1522) & (!g1571) & (!g2944) & (g3018) & (!g2948)) + ((!g827) & (g1522) & (!g1571) & (!g2944) & (g3018) & (g2948)) + ((!g827) & (g1522) & (!g1571) & (g2944) & (g3018) & (!g2948)) + ((!g827) & (g1522) & (!g1571) & (g2944) & (g3018) & (g2948)) + ((!g827) & (g1522) & (g1571) & (!g2944) & (g3018) & (!g2948)) + ((!g827) & (g1522) & (g1571) & (!g2944) & (g3018) & (g2948)) + ((!g827) & (g1522) & (g1571) & (g2944) & (g3018) & (!g2948)) + ((!g827) & (g1522) & (g1571) & (g2944) & (g3018) & (g2948)) + ((g827) & (!g1522) & (!g1571) & (!g2944) & (g3018) & (!g2948)) + ((g827) & (!g1522) & (!g1571) & (!g2944) & (g3018) & (g2948)) + ((g827) & (!g1522) & (!g1571) & (g2944) & (!g3018) & (!g2948)) + ((g827) & (!g1522) & (!g1571) & (g2944) & (g3018) & (g2948)) + ((g827) & (!g1522) & (g1571) & (!g2944) & (!g3018) & (!g2948)) + ((g827) & (!g1522) & (g1571) & (!g2944) & (!g3018) & (g2948)) + ((g827) & (!g1522) & (g1571) & (g2944) & (!g3018) & (g2948)) + ((g827) & (!g1522) & (g1571) & (g2944) & (g3018) & (!g2948)) + ((g827) & (g1522) & (!g1571) & (!g2944) & (!g3018) & (!g2948)) + ((g827) & (g1522) & (!g1571) & (!g2944) & (g3018) & (g2948)) + ((g827) & (g1522) & (!g1571) & (g2944) & (!g3018) & (!g2948)) + ((g827) & (g1522) & (!g1571) & (g2944) & (!g3018) & (g2948)) + ((g827) & (g1522) & (g1571) & (!g2944) & (!g3018) & (g2948)) + ((g827) & (g1522) & (g1571) & (!g2944) & (g3018) & (!g2948)) + ((g827) & (g1522) & (g1571) & (g2944) & (g3018) & (!g2948)) + ((g827) & (g1522) & (g1571) & (g2944) & (g3018) & (g2948)));
	assign g8175 = (((!g3429) & (g5225) & (!g3020)) + ((!g3429) & (g5225) & (g3020)) + ((g3429) & (!g5225) & (g3020)) + ((g3429) & (g5225) & (g3020)));
	assign g3021 = (((!g827) & (!g1530) & (!g1573) & (!g2968) & (g3020) & (!g2972)) + ((!g827) & (!g1530) & (!g1573) & (!g2968) & (g3020) & (g2972)) + ((!g827) & (!g1530) & (!g1573) & (g2968) & (g3020) & (!g2972)) + ((!g827) & (!g1530) & (!g1573) & (g2968) & (g3020) & (g2972)) + ((!g827) & (!g1530) & (g1573) & (!g2968) & (g3020) & (!g2972)) + ((!g827) & (!g1530) & (g1573) & (!g2968) & (g3020) & (g2972)) + ((!g827) & (!g1530) & (g1573) & (g2968) & (g3020) & (!g2972)) + ((!g827) & (!g1530) & (g1573) & (g2968) & (g3020) & (g2972)) + ((!g827) & (g1530) & (!g1573) & (!g2968) & (g3020) & (!g2972)) + ((!g827) & (g1530) & (!g1573) & (!g2968) & (g3020) & (g2972)) + ((!g827) & (g1530) & (!g1573) & (g2968) & (g3020) & (!g2972)) + ((!g827) & (g1530) & (!g1573) & (g2968) & (g3020) & (g2972)) + ((!g827) & (g1530) & (g1573) & (!g2968) & (g3020) & (!g2972)) + ((!g827) & (g1530) & (g1573) & (!g2968) & (g3020) & (g2972)) + ((!g827) & (g1530) & (g1573) & (g2968) & (g3020) & (!g2972)) + ((!g827) & (g1530) & (g1573) & (g2968) & (g3020) & (g2972)) + ((g827) & (!g1530) & (!g1573) & (!g2968) & (g3020) & (!g2972)) + ((g827) & (!g1530) & (!g1573) & (!g2968) & (g3020) & (g2972)) + ((g827) & (!g1530) & (!g1573) & (g2968) & (!g3020) & (!g2972)) + ((g827) & (!g1530) & (!g1573) & (g2968) & (g3020) & (g2972)) + ((g827) & (!g1530) & (g1573) & (!g2968) & (!g3020) & (!g2972)) + ((g827) & (!g1530) & (g1573) & (!g2968) & (!g3020) & (g2972)) + ((g827) & (!g1530) & (g1573) & (g2968) & (!g3020) & (g2972)) + ((g827) & (!g1530) & (g1573) & (g2968) & (g3020) & (!g2972)) + ((g827) & (g1530) & (!g1573) & (!g2968) & (!g3020) & (!g2972)) + ((g827) & (g1530) & (!g1573) & (!g2968) & (g3020) & (g2972)) + ((g827) & (g1530) & (!g1573) & (g2968) & (!g3020) & (!g2972)) + ((g827) & (g1530) & (!g1573) & (g2968) & (!g3020) & (g2972)) + ((g827) & (g1530) & (g1573) & (!g2968) & (!g3020) & (g2972)) + ((g827) & (g1530) & (g1573) & (!g2968) & (g3020) & (!g2972)) + ((g827) & (g1530) & (g1573) & (g2968) & (g3020) & (!g2972)) + ((g827) & (g1530) & (g1573) & (g2968) & (g3020) & (g2972)));
	assign g8176 = (((!g2017) & (g5230) & (!g3022)) + ((!g2017) & (g5230) & (g3022)) + ((g2017) & (!g5230) & (g3022)) + ((g2017) & (g5230) & (g3022)));
	assign g3023 = (((!g827) & (!g1538) & (!g1575) & (!g2991) & (g3022) & (!g2995)) + ((!g827) & (!g1538) & (!g1575) & (!g2991) & (g3022) & (g2995)) + ((!g827) & (!g1538) & (!g1575) & (g2991) & (g3022) & (!g2995)) + ((!g827) & (!g1538) & (!g1575) & (g2991) & (g3022) & (g2995)) + ((!g827) & (!g1538) & (g1575) & (!g2991) & (g3022) & (!g2995)) + ((!g827) & (!g1538) & (g1575) & (!g2991) & (g3022) & (g2995)) + ((!g827) & (!g1538) & (g1575) & (g2991) & (g3022) & (!g2995)) + ((!g827) & (!g1538) & (g1575) & (g2991) & (g3022) & (g2995)) + ((!g827) & (g1538) & (!g1575) & (!g2991) & (g3022) & (!g2995)) + ((!g827) & (g1538) & (!g1575) & (!g2991) & (g3022) & (g2995)) + ((!g827) & (g1538) & (!g1575) & (g2991) & (g3022) & (!g2995)) + ((!g827) & (g1538) & (!g1575) & (g2991) & (g3022) & (g2995)) + ((!g827) & (g1538) & (g1575) & (!g2991) & (g3022) & (!g2995)) + ((!g827) & (g1538) & (g1575) & (!g2991) & (g3022) & (g2995)) + ((!g827) & (g1538) & (g1575) & (g2991) & (g3022) & (!g2995)) + ((!g827) & (g1538) & (g1575) & (g2991) & (g3022) & (g2995)) + ((g827) & (!g1538) & (!g1575) & (!g2991) & (g3022) & (!g2995)) + ((g827) & (!g1538) & (!g1575) & (!g2991) & (g3022) & (g2995)) + ((g827) & (!g1538) & (!g1575) & (g2991) & (!g3022) & (!g2995)) + ((g827) & (!g1538) & (!g1575) & (g2991) & (g3022) & (g2995)) + ((g827) & (!g1538) & (g1575) & (!g2991) & (!g3022) & (!g2995)) + ((g827) & (!g1538) & (g1575) & (!g2991) & (!g3022) & (g2995)) + ((g827) & (!g1538) & (g1575) & (g2991) & (!g3022) & (g2995)) + ((g827) & (!g1538) & (g1575) & (g2991) & (g3022) & (!g2995)) + ((g827) & (g1538) & (!g1575) & (!g2991) & (!g3022) & (!g2995)) + ((g827) & (g1538) & (!g1575) & (!g2991) & (g3022) & (g2995)) + ((g827) & (g1538) & (!g1575) & (g2991) & (!g3022) & (!g2995)) + ((g827) & (g1538) & (!g1575) & (g2991) & (!g3022) & (g2995)) + ((g827) & (g1538) & (g1575) & (!g2991) & (!g3022) & (g2995)) + ((g827) & (g1538) & (g1575) & (!g2991) & (g3022) & (!g2995)) + ((g827) & (g1538) & (g1575) & (g2991) & (g3022) & (!g2995)) + ((g827) & (g1538) & (g1575) & (g2991) & (g3022) & (g2995)));
	assign g3024 = (((!g1943) & (g1944) & (g1945)) + ((g1943) & (!g1944) & (g1945)) + ((g1943) & (g1944) & (!g1945)) + ((g1943) & (g1944) & (g1945)));
	assign g3025 = (((g1914) & (!g3024) & (!g1946) & (g1947)) + ((g1914) & (!g3024) & (g1946) & (!g1947)) + ((g1914) & (g3024) & (!g1946) & (!g1947)) + ((g1914) & (g3024) & (g1946) & (g1947)));
	assign g3026 = (((!g1981) & (g1982) & (g1983)) + ((g1981) & (!g1982) & (g1983)) + ((g1981) & (g1982) & (!g1983)) + ((g1981) & (g1982) & (g1983)));
	assign g3027 = (((!g1914) & (!g3026) & (!g1984) & (g1985)) + ((!g1914) & (!g3026) & (g1984) & (!g1985)) + ((!g1914) & (g3026) & (!g1984) & (!g1985)) + ((!g1914) & (g3026) & (g1984) & (g1985)));
	assign g3028 = (((!g830) & (!g3025) & (!g3027) & (!g1577)) + ((!g830) & (!g3025) & (!g3027) & (g1577)) + ((!g830) & (!g3025) & (g3027) & (!g1577)) + ((!g830) & (!g3025) & (g3027) & (g1577)) + ((!g830) & (g3025) & (!g3027) & (!g1577)) + ((!g830) & (g3025) & (!g3027) & (g1577)) + ((!g830) & (g3025) & (g3027) & (!g1577)) + ((!g830) & (g3025) & (g3027) & (g1577)) + ((g830) & (!g3025) & (!g3027) & (g1577)) + ((g830) & (!g3025) & (g3027) & (!g1577)) + ((g830) & (g3025) & (!g3027) & (!g1577)) + ((g830) & (g3025) & (g3027) & (!g1577)));
	assign g3029 = (((!g1510) & (!g1553) & (!g2295) & (!g2343) & (!g2912) & (!g2913)) + ((!g1510) & (!g1553) & (!g2295) & (!g2343) & (!g2912) & (g2913)) + ((!g1510) & (!g1553) & (!g2295) & (!g2343) & (g2912) & (!g2913)) + ((!g1510) & (!g1553) & (!g2295) & (!g2343) & (g2912) & (g2913)) + ((!g1510) & (!g1553) & (!g2295) & (g2343) & (!g2912) & (!g2913)) + ((!g1510) & (!g1553) & (!g2295) & (g2343) & (!g2912) & (g2913)) + ((!g1510) & (!g1553) & (!g2295) & (g2343) & (g2912) & (!g2913)) + ((!g1510) & (!g1553) & (!g2295) & (g2343) & (g2912) & (g2913)) + ((!g1510) & (!g1553) & (g2295) & (!g2343) & (!g2912) & (!g2913)) + ((!g1510) & (!g1553) & (g2295) & (!g2343) & (!g2912) & (g2913)) + ((!g1510) & (!g1553) & (g2295) & (!g2343) & (g2912) & (!g2913)) + ((!g1510) & (!g1553) & (g2295) & (!g2343) & (g2912) & (g2913)) + ((!g1510) & (!g1553) & (g2295) & (g2343) & (!g2912) & (!g2913)) + ((!g1510) & (g1553) & (!g2295) & (!g2343) & (!g2912) & (!g2913)) + ((!g1510) & (g1553) & (!g2295) & (!g2343) & (!g2912) & (g2913)) + ((!g1510) & (g1553) & (!g2295) & (!g2343) & (g2912) & (!g2913)) + ((!g1510) & (g1553) & (!g2295) & (!g2343) & (g2912) & (g2913)) + ((!g1510) & (g1553) & (g2295) & (!g2343) & (!g2912) & (!g2913)) + ((g1510) & (!g1553) & (!g2295) & (!g2343) & (!g2912) & (!g2913)) + ((g1510) & (!g1553) & (!g2295) & (!g2343) & (!g2912) & (g2913)) + ((g1510) & (!g1553) & (!g2295) & (!g2343) & (g2912) & (!g2913)) + ((g1510) & (!g1553) & (!g2295) & (!g2343) & (g2912) & (g2913)) + ((g1510) & (!g1553) & (!g2295) & (g2343) & (!g2912) & (!g2913)) + ((g1510) & (!g1553) & (g2295) & (!g2343) & (!g2912) & (!g2913)) + ((g1510) & (!g1553) & (g2295) & (!g2343) & (!g2912) & (g2913)) + ((g1510) & (!g1553) & (g2295) & (!g2343) & (g2912) & (!g2913)) + ((g1510) & (!g1553) & (g2295) & (!g2343) & (g2912) & (g2913)) + ((g1510) & (g1553) & (!g2295) & (!g2343) & (!g2912) & (!g2913)));
	assign g3030 = (((!g827) & (!g1580) & (g2376) & (!g3029)) + ((!g827) & (!g1580) & (g2376) & (g3029)) + ((!g827) & (g1580) & (g2376) & (!g3029)) + ((!g827) & (g1580) & (g2376) & (g3029)) + ((g827) & (!g1580) & (!g2376) & (!g3029)) + ((g827) & (!g1580) & (g2376) & (g3029)) + ((g827) & (g1580) & (!g2376) & (g3029)) + ((g827) & (g1580) & (g2376) & (!g3029)));
	assign g8177 = (((!g3499) & (g5234) & (!g3031)) + ((!g3499) & (g5234) & (g3031)) + ((g3499) & (!g5234) & (g3031)) + ((g3499) & (g5234) & (g3031)));
	assign g3032 = (((!g1512) & (!g1561) & (!g2916) & (!g3009) & (!g2918) & (!g2919)) + ((!g1512) & (!g1561) & (!g2916) & (!g3009) & (!g2918) & (g2919)) + ((!g1512) & (!g1561) & (!g2916) & (!g3009) & (g2918) & (!g2919)) + ((!g1512) & (!g1561) & (!g2916) & (!g3009) & (g2918) & (g2919)) + ((!g1512) & (!g1561) & (!g2916) & (g3009) & (!g2918) & (!g2919)) + ((!g1512) & (!g1561) & (!g2916) & (g3009) & (!g2918) & (g2919)) + ((!g1512) & (!g1561) & (!g2916) & (g3009) & (g2918) & (!g2919)) + ((!g1512) & (!g1561) & (!g2916) & (g3009) & (g2918) & (g2919)) + ((!g1512) & (!g1561) & (g2916) & (!g3009) & (!g2918) & (!g2919)) + ((!g1512) & (!g1561) & (g2916) & (!g3009) & (!g2918) & (g2919)) + ((!g1512) & (!g1561) & (g2916) & (!g3009) & (g2918) & (!g2919)) + ((!g1512) & (!g1561) & (g2916) & (!g3009) & (g2918) & (g2919)) + ((!g1512) & (!g1561) & (g2916) & (g3009) & (!g2918) & (!g2919)) + ((!g1512) & (g1561) & (!g2916) & (!g3009) & (!g2918) & (!g2919)) + ((!g1512) & (g1561) & (!g2916) & (!g3009) & (!g2918) & (g2919)) + ((!g1512) & (g1561) & (!g2916) & (!g3009) & (g2918) & (!g2919)) + ((!g1512) & (g1561) & (!g2916) & (!g3009) & (g2918) & (g2919)) + ((!g1512) & (g1561) & (g2916) & (!g3009) & (!g2918) & (!g2919)) + ((g1512) & (!g1561) & (!g2916) & (!g3009) & (!g2918) & (!g2919)) + ((g1512) & (!g1561) & (!g2916) & (!g3009) & (!g2918) & (g2919)) + ((g1512) & (!g1561) & (!g2916) & (!g3009) & (g2918) & (!g2919)) + ((g1512) & (!g1561) & (!g2916) & (!g3009) & (g2918) & (g2919)) + ((g1512) & (!g1561) & (!g2916) & (g3009) & (!g2918) & (!g2919)) + ((g1512) & (!g1561) & (g2916) & (!g3009) & (!g2918) & (!g2919)) + ((g1512) & (!g1561) & (g2916) & (!g3009) & (!g2918) & (g2919)) + ((g1512) & (!g1561) & (g2916) & (!g3009) & (g2918) & (!g2919)) + ((g1512) & (!g1561) & (g2916) & (!g3009) & (g2918) & (g2919)) + ((g1512) & (g1561) & (!g2916) & (!g3009) & (!g2918) & (!g2919)));
	assign g3033 = (((!g827) & (!g1582) & (g3031) & (!g3032)) + ((!g827) & (!g1582) & (g3031) & (g3032)) + ((!g827) & (g1582) & (g3031) & (!g3032)) + ((!g827) & (g1582) & (g3031) & (g3032)) + ((g827) & (!g1582) & (!g3031) & (!g3032)) + ((g827) & (!g1582) & (g3031) & (g3032)) + ((g827) & (g1582) & (!g3031) & (g3032)) + ((g827) & (g1582) & (g3031) & (!g3032)));
	assign g3034 = (((!g1514) & (!g1569) & (!g2296) & (!g2344) & (!g2923) & (!g2924)) + ((!g1514) & (!g1569) & (!g2296) & (!g2344) & (!g2923) & (g2924)) + ((!g1514) & (!g1569) & (!g2296) & (!g2344) & (g2923) & (!g2924)) + ((!g1514) & (!g1569) & (!g2296) & (!g2344) & (g2923) & (g2924)) + ((!g1514) & (!g1569) & (!g2296) & (g2344) & (!g2923) & (!g2924)) + ((!g1514) & (!g1569) & (!g2296) & (g2344) & (!g2923) & (g2924)) + ((!g1514) & (!g1569) & (!g2296) & (g2344) & (g2923) & (!g2924)) + ((!g1514) & (!g1569) & (!g2296) & (g2344) & (g2923) & (g2924)) + ((!g1514) & (!g1569) & (g2296) & (!g2344) & (!g2923) & (!g2924)) + ((!g1514) & (!g1569) & (g2296) & (!g2344) & (!g2923) & (g2924)) + ((!g1514) & (!g1569) & (g2296) & (!g2344) & (g2923) & (!g2924)) + ((!g1514) & (!g1569) & (g2296) & (!g2344) & (g2923) & (g2924)) + ((!g1514) & (!g1569) & (g2296) & (g2344) & (!g2923) & (!g2924)) + ((!g1514) & (g1569) & (!g2296) & (!g2344) & (!g2923) & (!g2924)) + ((!g1514) & (g1569) & (!g2296) & (!g2344) & (!g2923) & (g2924)) + ((!g1514) & (g1569) & (!g2296) & (!g2344) & (g2923) & (!g2924)) + ((!g1514) & (g1569) & (!g2296) & (!g2344) & (g2923) & (g2924)) + ((!g1514) & (g1569) & (g2296) & (!g2344) & (!g2923) & (!g2924)) + ((g1514) & (!g1569) & (!g2296) & (!g2344) & (!g2923) & (!g2924)) + ((g1514) & (!g1569) & (!g2296) & (!g2344) & (!g2923) & (g2924)) + ((g1514) & (!g1569) & (!g2296) & (!g2344) & (g2923) & (!g2924)) + ((g1514) & (!g1569) & (!g2296) & (!g2344) & (g2923) & (g2924)) + ((g1514) & (!g1569) & (!g2296) & (g2344) & (!g2923) & (!g2924)) + ((g1514) & (!g1569) & (g2296) & (!g2344) & (!g2923) & (!g2924)) + ((g1514) & (!g1569) & (g2296) & (!g2344) & (!g2923) & (g2924)) + ((g1514) & (!g1569) & (g2296) & (!g2344) & (g2923) & (!g2924)) + ((g1514) & (!g1569) & (g2296) & (!g2344) & (g2923) & (g2924)) + ((g1514) & (g1569) & (!g2296) & (!g2344) & (!g2923) & (!g2924)));
	assign g3035 = (((!g827) & (!g1584) & (g2377) & (!g3034)) + ((!g827) & (!g1584) & (g2377) & (g3034)) + ((!g827) & (g1584) & (g2377) & (!g3034)) + ((!g827) & (g1584) & (g2377) & (g3034)) + ((g827) & (!g1584) & (!g2377) & (!g3034)) + ((g827) & (!g1584) & (g2377) & (g3034)) + ((g827) & (g1584) & (!g2377) & (g3034)) + ((g827) & (g1584) & (g2377) & (!g3034)));
	assign g3036 = (((!g1516) & (!g1547) & (!g2298) & (!g2347) & (!g2928) & (!g2929)) + ((!g1516) & (!g1547) & (!g2298) & (!g2347) & (!g2928) & (g2929)) + ((!g1516) & (!g1547) & (!g2298) & (!g2347) & (g2928) & (!g2929)) + ((!g1516) & (!g1547) & (!g2298) & (!g2347) & (g2928) & (g2929)) + ((!g1516) & (!g1547) & (!g2298) & (g2347) & (!g2928) & (!g2929)) + ((!g1516) & (!g1547) & (!g2298) & (g2347) & (!g2928) & (g2929)) + ((!g1516) & (!g1547) & (!g2298) & (g2347) & (g2928) & (!g2929)) + ((!g1516) & (!g1547) & (!g2298) & (g2347) & (g2928) & (g2929)) + ((!g1516) & (!g1547) & (g2298) & (!g2347) & (!g2928) & (!g2929)) + ((!g1516) & (!g1547) & (g2298) & (!g2347) & (!g2928) & (g2929)) + ((!g1516) & (!g1547) & (g2298) & (!g2347) & (g2928) & (!g2929)) + ((!g1516) & (!g1547) & (g2298) & (!g2347) & (g2928) & (g2929)) + ((!g1516) & (!g1547) & (g2298) & (g2347) & (!g2928) & (!g2929)) + ((!g1516) & (g1547) & (!g2298) & (!g2347) & (!g2928) & (!g2929)) + ((!g1516) & (g1547) & (!g2298) & (!g2347) & (!g2928) & (g2929)) + ((!g1516) & (g1547) & (!g2298) & (!g2347) & (g2928) & (!g2929)) + ((!g1516) & (g1547) & (!g2298) & (!g2347) & (g2928) & (g2929)) + ((!g1516) & (g1547) & (g2298) & (!g2347) & (!g2928) & (!g2929)) + ((g1516) & (!g1547) & (!g2298) & (!g2347) & (!g2928) & (!g2929)) + ((g1516) & (!g1547) & (!g2298) & (!g2347) & (!g2928) & (g2929)) + ((g1516) & (!g1547) & (!g2298) & (!g2347) & (g2928) & (!g2929)) + ((g1516) & (!g1547) & (!g2298) & (!g2347) & (g2928) & (g2929)) + ((g1516) & (!g1547) & (!g2298) & (g2347) & (!g2928) & (!g2929)) + ((g1516) & (!g1547) & (g2298) & (!g2347) & (!g2928) & (!g2929)) + ((g1516) & (!g1547) & (g2298) & (!g2347) & (!g2928) & (g2929)) + ((g1516) & (!g1547) & (g2298) & (!g2347) & (g2928) & (!g2929)) + ((g1516) & (!g1547) & (g2298) & (!g2347) & (g2928) & (g2929)) + ((g1516) & (g1547) & (!g2298) & (!g2347) & (!g2928) & (!g2929)));
	assign g3037 = (((!g827) & (!g1586) & (g2378) & (!g3036)) + ((!g827) & (!g1586) & (g2378) & (g3036)) + ((!g827) & (g1586) & (g2378) & (!g3036)) + ((!g827) & (g1586) & (g2378) & (g3036)) + ((g827) & (!g1586) & (!g2378) & (!g3036)) + ((g827) & (!g1586) & (g2378) & (g3036)) + ((g827) & (g1586) & (!g2378) & (g3036)) + ((g827) & (g1586) & (g2378) & (!g3036)));
	assign g8178 = (((!g2017) & (g5237) & (!g3038)) + ((!g2017) & (g5237) & (g3038)) + ((g2017) & (!g5237) & (g3038)) + ((g2017) & (g5237) & (g3038)));
	assign g3039 = (((!g1518) & (!g1555) & (!g2932) & (!g3003) & (!g2934) & (!g2935)) + ((!g1518) & (!g1555) & (!g2932) & (!g3003) & (!g2934) & (g2935)) + ((!g1518) & (!g1555) & (!g2932) & (!g3003) & (g2934) & (!g2935)) + ((!g1518) & (!g1555) & (!g2932) & (!g3003) & (g2934) & (g2935)) + ((!g1518) & (!g1555) & (!g2932) & (g3003) & (!g2934) & (!g2935)) + ((!g1518) & (!g1555) & (!g2932) & (g3003) & (!g2934) & (g2935)) + ((!g1518) & (!g1555) & (!g2932) & (g3003) & (g2934) & (!g2935)) + ((!g1518) & (!g1555) & (!g2932) & (g3003) & (g2934) & (g2935)) + ((!g1518) & (!g1555) & (g2932) & (!g3003) & (!g2934) & (!g2935)) + ((!g1518) & (!g1555) & (g2932) & (!g3003) & (!g2934) & (g2935)) + ((!g1518) & (!g1555) & (g2932) & (!g3003) & (g2934) & (!g2935)) + ((!g1518) & (!g1555) & (g2932) & (!g3003) & (g2934) & (g2935)) + ((!g1518) & (!g1555) & (g2932) & (g3003) & (!g2934) & (!g2935)) + ((!g1518) & (g1555) & (!g2932) & (!g3003) & (!g2934) & (!g2935)) + ((!g1518) & (g1555) & (!g2932) & (!g3003) & (!g2934) & (g2935)) + ((!g1518) & (g1555) & (!g2932) & (!g3003) & (g2934) & (!g2935)) + ((!g1518) & (g1555) & (!g2932) & (!g3003) & (g2934) & (g2935)) + ((!g1518) & (g1555) & (g2932) & (!g3003) & (!g2934) & (!g2935)) + ((g1518) & (!g1555) & (!g2932) & (!g3003) & (!g2934) & (!g2935)) + ((g1518) & (!g1555) & (!g2932) & (!g3003) & (!g2934) & (g2935)) + ((g1518) & (!g1555) & (!g2932) & (!g3003) & (g2934) & (!g2935)) + ((g1518) & (!g1555) & (!g2932) & (!g3003) & (g2934) & (g2935)) + ((g1518) & (!g1555) & (!g2932) & (g3003) & (!g2934) & (!g2935)) + ((g1518) & (!g1555) & (g2932) & (!g3003) & (!g2934) & (!g2935)) + ((g1518) & (!g1555) & (g2932) & (!g3003) & (!g2934) & (g2935)) + ((g1518) & (!g1555) & (g2932) & (!g3003) & (g2934) & (!g2935)) + ((g1518) & (!g1555) & (g2932) & (!g3003) & (g2934) & (g2935)) + ((g1518) & (g1555) & (!g2932) & (!g3003) & (!g2934) & (!g2935)));
	assign g3040 = (((!g827) & (!g1588) & (g3038) & (!g3039)) + ((!g827) & (!g1588) & (g3038) & (g3039)) + ((!g827) & (g1588) & (g3038) & (!g3039)) + ((!g827) & (g1588) & (g3038) & (g3039)) + ((g827) & (!g1588) & (!g3038) & (!g3039)) + ((g827) & (!g1588) & (g3038) & (g3039)) + ((g827) & (g1588) & (!g3038) & (g3039)) + ((g827) & (g1588) & (g3038) & (!g3039)));
	assign g8179 = (((!g3464) & (g5242) & (!g3041)) + ((!g3464) & (g5242) & (g3041)) + ((g3464) & (!g5242) & (g3041)) + ((g3464) & (g5242) & (g3041)));
	assign g3042 = (((!g1520) & (!g1563) & (!g2938) & (!g3011) & (!g2940) & (!g2941)) + ((!g1520) & (!g1563) & (!g2938) & (!g3011) & (!g2940) & (g2941)) + ((!g1520) & (!g1563) & (!g2938) & (!g3011) & (g2940) & (!g2941)) + ((!g1520) & (!g1563) & (!g2938) & (!g3011) & (g2940) & (g2941)) + ((!g1520) & (!g1563) & (!g2938) & (g3011) & (!g2940) & (!g2941)) + ((!g1520) & (!g1563) & (!g2938) & (g3011) & (!g2940) & (g2941)) + ((!g1520) & (!g1563) & (!g2938) & (g3011) & (g2940) & (!g2941)) + ((!g1520) & (!g1563) & (!g2938) & (g3011) & (g2940) & (g2941)) + ((!g1520) & (!g1563) & (g2938) & (!g3011) & (!g2940) & (!g2941)) + ((!g1520) & (!g1563) & (g2938) & (!g3011) & (!g2940) & (g2941)) + ((!g1520) & (!g1563) & (g2938) & (!g3011) & (g2940) & (!g2941)) + ((!g1520) & (!g1563) & (g2938) & (!g3011) & (g2940) & (g2941)) + ((!g1520) & (!g1563) & (g2938) & (g3011) & (!g2940) & (!g2941)) + ((!g1520) & (g1563) & (!g2938) & (!g3011) & (!g2940) & (!g2941)) + ((!g1520) & (g1563) & (!g2938) & (!g3011) & (!g2940) & (g2941)) + ((!g1520) & (g1563) & (!g2938) & (!g3011) & (g2940) & (!g2941)) + ((!g1520) & (g1563) & (!g2938) & (!g3011) & (g2940) & (g2941)) + ((!g1520) & (g1563) & (g2938) & (!g3011) & (!g2940) & (!g2941)) + ((g1520) & (!g1563) & (!g2938) & (!g3011) & (!g2940) & (!g2941)) + ((g1520) & (!g1563) & (!g2938) & (!g3011) & (!g2940) & (g2941)) + ((g1520) & (!g1563) & (!g2938) & (!g3011) & (g2940) & (!g2941)) + ((g1520) & (!g1563) & (!g2938) & (!g3011) & (g2940) & (g2941)) + ((g1520) & (!g1563) & (!g2938) & (g3011) & (!g2940) & (!g2941)) + ((g1520) & (!g1563) & (g2938) & (!g3011) & (!g2940) & (!g2941)) + ((g1520) & (!g1563) & (g2938) & (!g3011) & (!g2940) & (g2941)) + ((g1520) & (!g1563) & (g2938) & (!g3011) & (g2940) & (!g2941)) + ((g1520) & (!g1563) & (g2938) & (!g3011) & (g2940) & (g2941)) + ((g1520) & (g1563) & (!g2938) & (!g3011) & (!g2940) & (!g2941)));
	assign g3043 = (((!g827) & (!g1590) & (g3041) & (!g3042)) + ((!g827) & (!g1590) & (g3041) & (g3042)) + ((!g827) & (g1590) & (g3041) & (!g3042)) + ((!g827) & (g1590) & (g3041) & (g3042)) + ((g827) & (!g1590) & (!g3041) & (!g3042)) + ((g827) & (!g1590) & (g3041) & (g3042)) + ((g827) & (g1590) & (!g3041) & (g3042)) + ((g827) & (g1590) & (g3041) & (!g3042)));
	assign g8180 = (((!g3499) & (g5246) & (!g3044)) + ((!g3499) & (g5246) & (g3044)) + ((g3499) & (!g5246) & (g3044)) + ((g3499) & (g5246) & (g3044)));
	assign g3045 = (((!g1522) & (!g1571) & (!g2944) & (!g3018) & (!g2946) & (!g2947)) + ((!g1522) & (!g1571) & (!g2944) & (!g3018) & (!g2946) & (g2947)) + ((!g1522) & (!g1571) & (!g2944) & (!g3018) & (g2946) & (!g2947)) + ((!g1522) & (!g1571) & (!g2944) & (!g3018) & (g2946) & (g2947)) + ((!g1522) & (!g1571) & (!g2944) & (g3018) & (!g2946) & (!g2947)) + ((!g1522) & (!g1571) & (!g2944) & (g3018) & (!g2946) & (g2947)) + ((!g1522) & (!g1571) & (!g2944) & (g3018) & (g2946) & (!g2947)) + ((!g1522) & (!g1571) & (!g2944) & (g3018) & (g2946) & (g2947)) + ((!g1522) & (!g1571) & (g2944) & (!g3018) & (!g2946) & (!g2947)) + ((!g1522) & (!g1571) & (g2944) & (!g3018) & (!g2946) & (g2947)) + ((!g1522) & (!g1571) & (g2944) & (!g3018) & (g2946) & (!g2947)) + ((!g1522) & (!g1571) & (g2944) & (!g3018) & (g2946) & (g2947)) + ((!g1522) & (!g1571) & (g2944) & (g3018) & (!g2946) & (!g2947)) + ((!g1522) & (g1571) & (!g2944) & (!g3018) & (!g2946) & (!g2947)) + ((!g1522) & (g1571) & (!g2944) & (!g3018) & (!g2946) & (g2947)) + ((!g1522) & (g1571) & (!g2944) & (!g3018) & (g2946) & (!g2947)) + ((!g1522) & (g1571) & (!g2944) & (!g3018) & (g2946) & (g2947)) + ((!g1522) & (g1571) & (g2944) & (!g3018) & (!g2946) & (!g2947)) + ((g1522) & (!g1571) & (!g2944) & (!g3018) & (!g2946) & (!g2947)) + ((g1522) & (!g1571) & (!g2944) & (!g3018) & (!g2946) & (g2947)) + ((g1522) & (!g1571) & (!g2944) & (!g3018) & (g2946) & (!g2947)) + ((g1522) & (!g1571) & (!g2944) & (!g3018) & (g2946) & (g2947)) + ((g1522) & (!g1571) & (!g2944) & (g3018) & (!g2946) & (!g2947)) + ((g1522) & (!g1571) & (g2944) & (!g3018) & (!g2946) & (!g2947)) + ((g1522) & (!g1571) & (g2944) & (!g3018) & (!g2946) & (g2947)) + ((g1522) & (!g1571) & (g2944) & (!g3018) & (g2946) & (!g2947)) + ((g1522) & (!g1571) & (g2944) & (!g3018) & (g2946) & (g2947)) + ((g1522) & (g1571) & (!g2944) & (!g3018) & (!g2946) & (!g2947)));
	assign g3046 = (((!g827) & (!g1592) & (g3044) & (!g3045)) + ((!g827) & (!g1592) & (g3044) & (g3045)) + ((!g827) & (g1592) & (g3044) & (!g3045)) + ((!g827) & (g1592) & (g3044) & (g3045)) + ((g827) & (!g1592) & (!g3044) & (!g3045)) + ((g827) & (!g1592) & (g3044) & (g3045)) + ((g827) & (g1592) & (!g3044) & (g3045)) + ((g827) & (g1592) & (g3044) & (!g3045)));
	assign g8181 = (((!g3464) & (g5250) & (!g3047)) + ((!g3464) & (g5250) & (g3047)) + ((g3464) & (!g5250) & (g3047)) + ((g3464) & (g5250) & (g3047)));
	assign g3048 = (((!g1524) & (!g1549) & (!g2950) & (!g2999) & (!g2952) & (!g2953)) + ((!g1524) & (!g1549) & (!g2950) & (!g2999) & (!g2952) & (g2953)) + ((!g1524) & (!g1549) & (!g2950) & (!g2999) & (g2952) & (!g2953)) + ((!g1524) & (!g1549) & (!g2950) & (!g2999) & (g2952) & (g2953)) + ((!g1524) & (!g1549) & (!g2950) & (g2999) & (!g2952) & (!g2953)) + ((!g1524) & (!g1549) & (!g2950) & (g2999) & (!g2952) & (g2953)) + ((!g1524) & (!g1549) & (!g2950) & (g2999) & (g2952) & (!g2953)) + ((!g1524) & (!g1549) & (!g2950) & (g2999) & (g2952) & (g2953)) + ((!g1524) & (!g1549) & (g2950) & (!g2999) & (!g2952) & (!g2953)) + ((!g1524) & (!g1549) & (g2950) & (!g2999) & (!g2952) & (g2953)) + ((!g1524) & (!g1549) & (g2950) & (!g2999) & (g2952) & (!g2953)) + ((!g1524) & (!g1549) & (g2950) & (!g2999) & (g2952) & (g2953)) + ((!g1524) & (!g1549) & (g2950) & (g2999) & (!g2952) & (!g2953)) + ((!g1524) & (g1549) & (!g2950) & (!g2999) & (!g2952) & (!g2953)) + ((!g1524) & (g1549) & (!g2950) & (!g2999) & (!g2952) & (g2953)) + ((!g1524) & (g1549) & (!g2950) & (!g2999) & (g2952) & (!g2953)) + ((!g1524) & (g1549) & (!g2950) & (!g2999) & (g2952) & (g2953)) + ((!g1524) & (g1549) & (g2950) & (!g2999) & (!g2952) & (!g2953)) + ((g1524) & (!g1549) & (!g2950) & (!g2999) & (!g2952) & (!g2953)) + ((g1524) & (!g1549) & (!g2950) & (!g2999) & (!g2952) & (g2953)) + ((g1524) & (!g1549) & (!g2950) & (!g2999) & (g2952) & (!g2953)) + ((g1524) & (!g1549) & (!g2950) & (!g2999) & (g2952) & (g2953)) + ((g1524) & (!g1549) & (!g2950) & (g2999) & (!g2952) & (!g2953)) + ((g1524) & (!g1549) & (g2950) & (!g2999) & (!g2952) & (!g2953)) + ((g1524) & (!g1549) & (g2950) & (!g2999) & (!g2952) & (g2953)) + ((g1524) & (!g1549) & (g2950) & (!g2999) & (g2952) & (!g2953)) + ((g1524) & (!g1549) & (g2950) & (!g2999) & (g2952) & (g2953)) + ((g1524) & (g1549) & (!g2950) & (!g2999) & (!g2952) & (!g2953)));
	assign g3049 = (((!g827) & (!g1594) & (g3047) & (!g3048)) + ((!g827) & (!g1594) & (g3047) & (g3048)) + ((!g827) & (g1594) & (g3047) & (!g3048)) + ((!g827) & (g1594) & (g3047) & (g3048)) + ((g827) & (!g1594) & (!g3047) & (!g3048)) + ((g827) & (!g1594) & (g3047) & (g3048)) + ((g827) & (g1594) & (!g3047) & (g3048)) + ((g827) & (g1594) & (g3047) & (!g3048)));
	assign g8182 = (((!g3499) & (g5254) & (!g3050)) + ((!g3499) & (g5254) & (g3050)) + ((g3499) & (!g5254) & (g3050)) + ((g3499) & (g5254) & (g3050)));
	assign g3051 = (((!g1526) & (!g1557) & (!g2956) & (!g3005) & (!g2958) & (!g2959)) + ((!g1526) & (!g1557) & (!g2956) & (!g3005) & (!g2958) & (g2959)) + ((!g1526) & (!g1557) & (!g2956) & (!g3005) & (g2958) & (!g2959)) + ((!g1526) & (!g1557) & (!g2956) & (!g3005) & (g2958) & (g2959)) + ((!g1526) & (!g1557) & (!g2956) & (g3005) & (!g2958) & (!g2959)) + ((!g1526) & (!g1557) & (!g2956) & (g3005) & (!g2958) & (g2959)) + ((!g1526) & (!g1557) & (!g2956) & (g3005) & (g2958) & (!g2959)) + ((!g1526) & (!g1557) & (!g2956) & (g3005) & (g2958) & (g2959)) + ((!g1526) & (!g1557) & (g2956) & (!g3005) & (!g2958) & (!g2959)) + ((!g1526) & (!g1557) & (g2956) & (!g3005) & (!g2958) & (g2959)) + ((!g1526) & (!g1557) & (g2956) & (!g3005) & (g2958) & (!g2959)) + ((!g1526) & (!g1557) & (g2956) & (!g3005) & (g2958) & (g2959)) + ((!g1526) & (!g1557) & (g2956) & (g3005) & (!g2958) & (!g2959)) + ((!g1526) & (g1557) & (!g2956) & (!g3005) & (!g2958) & (!g2959)) + ((!g1526) & (g1557) & (!g2956) & (!g3005) & (!g2958) & (g2959)) + ((!g1526) & (g1557) & (!g2956) & (!g3005) & (g2958) & (!g2959)) + ((!g1526) & (g1557) & (!g2956) & (!g3005) & (g2958) & (g2959)) + ((!g1526) & (g1557) & (g2956) & (!g3005) & (!g2958) & (!g2959)) + ((g1526) & (!g1557) & (!g2956) & (!g3005) & (!g2958) & (!g2959)) + ((g1526) & (!g1557) & (!g2956) & (!g3005) & (!g2958) & (g2959)) + ((g1526) & (!g1557) & (!g2956) & (!g3005) & (g2958) & (!g2959)) + ((g1526) & (!g1557) & (!g2956) & (!g3005) & (g2958) & (g2959)) + ((g1526) & (!g1557) & (!g2956) & (g3005) & (!g2958) & (!g2959)) + ((g1526) & (!g1557) & (g2956) & (!g3005) & (!g2958) & (!g2959)) + ((g1526) & (!g1557) & (g2956) & (!g3005) & (!g2958) & (g2959)) + ((g1526) & (!g1557) & (g2956) & (!g3005) & (g2958) & (!g2959)) + ((g1526) & (!g1557) & (g2956) & (!g3005) & (g2958) & (g2959)) + ((g1526) & (g1557) & (!g2956) & (!g3005) & (!g2958) & (!g2959)));
	assign g3052 = (((!g827) & (!g1596) & (g3050) & (!g3051)) + ((!g827) & (!g1596) & (g3050) & (g3051)) + ((!g827) & (g1596) & (g3050) & (!g3051)) + ((!g827) & (g1596) & (g3050) & (g3051)) + ((g827) & (!g1596) & (!g3050) & (!g3051)) + ((g827) & (!g1596) & (g3050) & (g3051)) + ((g827) & (g1596) & (!g3050) & (g3051)) + ((g827) & (g1596) & (g3050) & (!g3051)));
	assign g8183 = (((!g2017) & (g5257) & (!g3053)) + ((!g2017) & (g5257) & (g3053)) + ((g2017) & (!g5257) & (g3053)) + ((g2017) & (g5257) & (g3053)));
	assign g3054 = (((!g1528) & (!g1565) & (!g2962) & (!g3013) & (!g2964) & (!g2965)) + ((!g1528) & (!g1565) & (!g2962) & (!g3013) & (!g2964) & (g2965)) + ((!g1528) & (!g1565) & (!g2962) & (!g3013) & (g2964) & (!g2965)) + ((!g1528) & (!g1565) & (!g2962) & (!g3013) & (g2964) & (g2965)) + ((!g1528) & (!g1565) & (!g2962) & (g3013) & (!g2964) & (!g2965)) + ((!g1528) & (!g1565) & (!g2962) & (g3013) & (!g2964) & (g2965)) + ((!g1528) & (!g1565) & (!g2962) & (g3013) & (g2964) & (!g2965)) + ((!g1528) & (!g1565) & (!g2962) & (g3013) & (g2964) & (g2965)) + ((!g1528) & (!g1565) & (g2962) & (!g3013) & (!g2964) & (!g2965)) + ((!g1528) & (!g1565) & (g2962) & (!g3013) & (!g2964) & (g2965)) + ((!g1528) & (!g1565) & (g2962) & (!g3013) & (g2964) & (!g2965)) + ((!g1528) & (!g1565) & (g2962) & (!g3013) & (g2964) & (g2965)) + ((!g1528) & (!g1565) & (g2962) & (g3013) & (!g2964) & (!g2965)) + ((!g1528) & (g1565) & (!g2962) & (!g3013) & (!g2964) & (!g2965)) + ((!g1528) & (g1565) & (!g2962) & (!g3013) & (!g2964) & (g2965)) + ((!g1528) & (g1565) & (!g2962) & (!g3013) & (g2964) & (!g2965)) + ((!g1528) & (g1565) & (!g2962) & (!g3013) & (g2964) & (g2965)) + ((!g1528) & (g1565) & (g2962) & (!g3013) & (!g2964) & (!g2965)) + ((g1528) & (!g1565) & (!g2962) & (!g3013) & (!g2964) & (!g2965)) + ((g1528) & (!g1565) & (!g2962) & (!g3013) & (!g2964) & (g2965)) + ((g1528) & (!g1565) & (!g2962) & (!g3013) & (g2964) & (!g2965)) + ((g1528) & (!g1565) & (!g2962) & (!g3013) & (g2964) & (g2965)) + ((g1528) & (!g1565) & (!g2962) & (g3013) & (!g2964) & (!g2965)) + ((g1528) & (!g1565) & (g2962) & (!g3013) & (!g2964) & (!g2965)) + ((g1528) & (!g1565) & (g2962) & (!g3013) & (!g2964) & (g2965)) + ((g1528) & (!g1565) & (g2962) & (!g3013) & (g2964) & (!g2965)) + ((g1528) & (!g1565) & (g2962) & (!g3013) & (g2964) & (g2965)) + ((g1528) & (g1565) & (!g2962) & (!g3013) & (!g2964) & (!g2965)));
	assign g3055 = (((!g827) & (!g1598) & (g3053) & (!g3054)) + ((!g827) & (!g1598) & (g3053) & (g3054)) + ((!g827) & (g1598) & (g3053) & (!g3054)) + ((!g827) & (g1598) & (g3053) & (g3054)) + ((g827) & (!g1598) & (!g3053) & (!g3054)) + ((g827) & (!g1598) & (g3053) & (g3054)) + ((g827) & (g1598) & (!g3053) & (g3054)) + ((g827) & (g1598) & (g3053) & (!g3054)));
	assign g8184 = (((!g3429) & (g5262) & (!g3056)) + ((!g3429) & (g5262) & (g3056)) + ((g3429) & (!g5262) & (g3056)) + ((g3429) & (g5262) & (g3056)));
	assign g3057 = (((!g1530) & (!g1573) & (!g2968) & (!g3020) & (!g2970) & (!g2971)) + ((!g1530) & (!g1573) & (!g2968) & (!g3020) & (!g2970) & (g2971)) + ((!g1530) & (!g1573) & (!g2968) & (!g3020) & (g2970) & (!g2971)) + ((!g1530) & (!g1573) & (!g2968) & (!g3020) & (g2970) & (g2971)) + ((!g1530) & (!g1573) & (!g2968) & (g3020) & (!g2970) & (!g2971)) + ((!g1530) & (!g1573) & (!g2968) & (g3020) & (!g2970) & (g2971)) + ((!g1530) & (!g1573) & (!g2968) & (g3020) & (g2970) & (!g2971)) + ((!g1530) & (!g1573) & (!g2968) & (g3020) & (g2970) & (g2971)) + ((!g1530) & (!g1573) & (g2968) & (!g3020) & (!g2970) & (!g2971)) + ((!g1530) & (!g1573) & (g2968) & (!g3020) & (!g2970) & (g2971)) + ((!g1530) & (!g1573) & (g2968) & (!g3020) & (g2970) & (!g2971)) + ((!g1530) & (!g1573) & (g2968) & (!g3020) & (g2970) & (g2971)) + ((!g1530) & (!g1573) & (g2968) & (g3020) & (!g2970) & (!g2971)) + ((!g1530) & (g1573) & (!g2968) & (!g3020) & (!g2970) & (!g2971)) + ((!g1530) & (g1573) & (!g2968) & (!g3020) & (!g2970) & (g2971)) + ((!g1530) & (g1573) & (!g2968) & (!g3020) & (g2970) & (!g2971)) + ((!g1530) & (g1573) & (!g2968) & (!g3020) & (g2970) & (g2971)) + ((!g1530) & (g1573) & (g2968) & (!g3020) & (!g2970) & (!g2971)) + ((g1530) & (!g1573) & (!g2968) & (!g3020) & (!g2970) & (!g2971)) + ((g1530) & (!g1573) & (!g2968) & (!g3020) & (!g2970) & (g2971)) + ((g1530) & (!g1573) & (!g2968) & (!g3020) & (g2970) & (!g2971)) + ((g1530) & (!g1573) & (!g2968) & (!g3020) & (g2970) & (g2971)) + ((g1530) & (!g1573) & (!g2968) & (g3020) & (!g2970) & (!g2971)) + ((g1530) & (!g1573) & (g2968) & (!g3020) & (!g2970) & (!g2971)) + ((g1530) & (!g1573) & (g2968) & (!g3020) & (!g2970) & (g2971)) + ((g1530) & (!g1573) & (g2968) & (!g3020) & (g2970) & (!g2971)) + ((g1530) & (!g1573) & (g2968) & (!g3020) & (g2970) & (g2971)) + ((g1530) & (g1573) & (!g2968) & (!g3020) & (!g2970) & (!g2971)));
	assign g3058 = (((!g827) & (!g1600) & (g3056) & (!g3057)) + ((!g827) & (!g1600) & (g3056) & (g3057)) + ((!g827) & (g1600) & (g3056) & (!g3057)) + ((!g827) & (g1600) & (g3056) & (g3057)) + ((g827) & (!g1600) & (!g3056) & (!g3057)) + ((g827) & (!g1600) & (g3056) & (g3057)) + ((g827) & (g1600) & (!g3056) & (g3057)) + ((g827) & (g1600) & (g3056) & (!g3057)));
	assign g3059 = (((!g1532) & (!g1551) & (!g2299) & (!g2348) & (!g2975) & (!g2976)) + ((!g1532) & (!g1551) & (!g2299) & (!g2348) & (!g2975) & (g2976)) + ((!g1532) & (!g1551) & (!g2299) & (!g2348) & (g2975) & (!g2976)) + ((!g1532) & (!g1551) & (!g2299) & (!g2348) & (g2975) & (g2976)) + ((!g1532) & (!g1551) & (!g2299) & (g2348) & (!g2975) & (!g2976)) + ((!g1532) & (!g1551) & (!g2299) & (g2348) & (!g2975) & (g2976)) + ((!g1532) & (!g1551) & (!g2299) & (g2348) & (g2975) & (!g2976)) + ((!g1532) & (!g1551) & (!g2299) & (g2348) & (g2975) & (g2976)) + ((!g1532) & (!g1551) & (g2299) & (!g2348) & (!g2975) & (!g2976)) + ((!g1532) & (!g1551) & (g2299) & (!g2348) & (!g2975) & (g2976)) + ((!g1532) & (!g1551) & (g2299) & (!g2348) & (g2975) & (!g2976)) + ((!g1532) & (!g1551) & (g2299) & (!g2348) & (g2975) & (g2976)) + ((!g1532) & (!g1551) & (g2299) & (g2348) & (!g2975) & (!g2976)) + ((!g1532) & (g1551) & (!g2299) & (!g2348) & (!g2975) & (!g2976)) + ((!g1532) & (g1551) & (!g2299) & (!g2348) & (!g2975) & (g2976)) + ((!g1532) & (g1551) & (!g2299) & (!g2348) & (g2975) & (!g2976)) + ((!g1532) & (g1551) & (!g2299) & (!g2348) & (g2975) & (g2976)) + ((!g1532) & (g1551) & (g2299) & (!g2348) & (!g2975) & (!g2976)) + ((g1532) & (!g1551) & (!g2299) & (!g2348) & (!g2975) & (!g2976)) + ((g1532) & (!g1551) & (!g2299) & (!g2348) & (!g2975) & (g2976)) + ((g1532) & (!g1551) & (!g2299) & (!g2348) & (g2975) & (!g2976)) + ((g1532) & (!g1551) & (!g2299) & (!g2348) & (g2975) & (g2976)) + ((g1532) & (!g1551) & (!g2299) & (g2348) & (!g2975) & (!g2976)) + ((g1532) & (!g1551) & (g2299) & (!g2348) & (!g2975) & (!g2976)) + ((g1532) & (!g1551) & (g2299) & (!g2348) & (!g2975) & (g2976)) + ((g1532) & (!g1551) & (g2299) & (!g2348) & (g2975) & (!g2976)) + ((g1532) & (!g1551) & (g2299) & (!g2348) & (g2975) & (g2976)) + ((g1532) & (g1551) & (!g2299) & (!g2348) & (!g2975) & (!g2976)));
	assign g3060 = (((!g827) & (!g1602) & (g2379) & (!g3059)) + ((!g827) & (!g1602) & (g2379) & (g3059)) + ((!g827) & (g1602) & (g2379) & (!g3059)) + ((!g827) & (g1602) & (g2379) & (g3059)) + ((g827) & (!g1602) & (!g2379) & (!g3059)) + ((g827) & (!g1602) & (g2379) & (g3059)) + ((g827) & (g1602) & (!g2379) & (g3059)) + ((g827) & (g1602) & (g2379) & (!g3059)));
	assign g8185 = (((!g3464) & (g5266) & (!g3061)) + ((!g3464) & (g5266) & (g3061)) + ((g3464) & (!g5266) & (g3061)) + ((g3464) & (g5266) & (g3061)));
	assign g3062 = (((!g1534) & (!g1559) & (!g2979) & (!g3007) & (!g2981) & (!g2982)) + ((!g1534) & (!g1559) & (!g2979) & (!g3007) & (!g2981) & (g2982)) + ((!g1534) & (!g1559) & (!g2979) & (!g3007) & (g2981) & (!g2982)) + ((!g1534) & (!g1559) & (!g2979) & (!g3007) & (g2981) & (g2982)) + ((!g1534) & (!g1559) & (!g2979) & (g3007) & (!g2981) & (!g2982)) + ((!g1534) & (!g1559) & (!g2979) & (g3007) & (!g2981) & (g2982)) + ((!g1534) & (!g1559) & (!g2979) & (g3007) & (g2981) & (!g2982)) + ((!g1534) & (!g1559) & (!g2979) & (g3007) & (g2981) & (g2982)) + ((!g1534) & (!g1559) & (g2979) & (!g3007) & (!g2981) & (!g2982)) + ((!g1534) & (!g1559) & (g2979) & (!g3007) & (!g2981) & (g2982)) + ((!g1534) & (!g1559) & (g2979) & (!g3007) & (g2981) & (!g2982)) + ((!g1534) & (!g1559) & (g2979) & (!g3007) & (g2981) & (g2982)) + ((!g1534) & (!g1559) & (g2979) & (g3007) & (!g2981) & (!g2982)) + ((!g1534) & (g1559) & (!g2979) & (!g3007) & (!g2981) & (!g2982)) + ((!g1534) & (g1559) & (!g2979) & (!g3007) & (!g2981) & (g2982)) + ((!g1534) & (g1559) & (!g2979) & (!g3007) & (g2981) & (!g2982)) + ((!g1534) & (g1559) & (!g2979) & (!g3007) & (g2981) & (g2982)) + ((!g1534) & (g1559) & (g2979) & (!g3007) & (!g2981) & (!g2982)) + ((g1534) & (!g1559) & (!g2979) & (!g3007) & (!g2981) & (!g2982)) + ((g1534) & (!g1559) & (!g2979) & (!g3007) & (!g2981) & (g2982)) + ((g1534) & (!g1559) & (!g2979) & (!g3007) & (g2981) & (!g2982)) + ((g1534) & (!g1559) & (!g2979) & (!g3007) & (g2981) & (g2982)) + ((g1534) & (!g1559) & (!g2979) & (g3007) & (!g2981) & (!g2982)) + ((g1534) & (!g1559) & (g2979) & (!g3007) & (!g2981) & (!g2982)) + ((g1534) & (!g1559) & (g2979) & (!g3007) & (!g2981) & (g2982)) + ((g1534) & (!g1559) & (g2979) & (!g3007) & (g2981) & (!g2982)) + ((g1534) & (!g1559) & (g2979) & (!g3007) & (g2981) & (g2982)) + ((g1534) & (g1559) & (!g2979) & (!g3007) & (!g2981) & (!g2982)));
	assign g3063 = (((!g827) & (!g1604) & (g3061) & (!g3062)) + ((!g827) & (!g1604) & (g3061) & (g3062)) + ((!g827) & (g1604) & (g3061) & (!g3062)) + ((!g827) & (g1604) & (g3061) & (g3062)) + ((g827) & (!g1604) & (!g3061) & (!g3062)) + ((g827) & (!g1604) & (g3061) & (g3062)) + ((g827) & (g1604) & (!g3061) & (g3062)) + ((g827) & (g1604) & (g3061) & (!g3062)));
	assign g8186 = (((!g3429) & (g5271) & (!g3064)) + ((!g3429) & (g5271) & (g3064)) + ((g3429) & (!g5271) & (g3064)) + ((g3429) & (g5271) & (g3064)));
	assign g3065 = (((!g1536) & (!g1567) & (!g2985) & (!g3015) & (!g2987) & (!g2988)) + ((!g1536) & (!g1567) & (!g2985) & (!g3015) & (!g2987) & (g2988)) + ((!g1536) & (!g1567) & (!g2985) & (!g3015) & (g2987) & (!g2988)) + ((!g1536) & (!g1567) & (!g2985) & (!g3015) & (g2987) & (g2988)) + ((!g1536) & (!g1567) & (!g2985) & (g3015) & (!g2987) & (!g2988)) + ((!g1536) & (!g1567) & (!g2985) & (g3015) & (!g2987) & (g2988)) + ((!g1536) & (!g1567) & (!g2985) & (g3015) & (g2987) & (!g2988)) + ((!g1536) & (!g1567) & (!g2985) & (g3015) & (g2987) & (g2988)) + ((!g1536) & (!g1567) & (g2985) & (!g3015) & (!g2987) & (!g2988)) + ((!g1536) & (!g1567) & (g2985) & (!g3015) & (!g2987) & (g2988)) + ((!g1536) & (!g1567) & (g2985) & (!g3015) & (g2987) & (!g2988)) + ((!g1536) & (!g1567) & (g2985) & (!g3015) & (g2987) & (g2988)) + ((!g1536) & (!g1567) & (g2985) & (g3015) & (!g2987) & (!g2988)) + ((!g1536) & (g1567) & (!g2985) & (!g3015) & (!g2987) & (!g2988)) + ((!g1536) & (g1567) & (!g2985) & (!g3015) & (!g2987) & (g2988)) + ((!g1536) & (g1567) & (!g2985) & (!g3015) & (g2987) & (!g2988)) + ((!g1536) & (g1567) & (!g2985) & (!g3015) & (g2987) & (g2988)) + ((!g1536) & (g1567) & (g2985) & (!g3015) & (!g2987) & (!g2988)) + ((g1536) & (!g1567) & (!g2985) & (!g3015) & (!g2987) & (!g2988)) + ((g1536) & (!g1567) & (!g2985) & (!g3015) & (!g2987) & (g2988)) + ((g1536) & (!g1567) & (!g2985) & (!g3015) & (g2987) & (!g2988)) + ((g1536) & (!g1567) & (!g2985) & (!g3015) & (g2987) & (g2988)) + ((g1536) & (!g1567) & (!g2985) & (g3015) & (!g2987) & (!g2988)) + ((g1536) & (!g1567) & (g2985) & (!g3015) & (!g2987) & (!g2988)) + ((g1536) & (!g1567) & (g2985) & (!g3015) & (!g2987) & (g2988)) + ((g1536) & (!g1567) & (g2985) & (!g3015) & (g2987) & (!g2988)) + ((g1536) & (!g1567) & (g2985) & (!g3015) & (g2987) & (g2988)) + ((g1536) & (g1567) & (!g2985) & (!g3015) & (!g2987) & (!g2988)));
	assign g3066 = (((!g827) & (!g1606) & (g3064) & (!g3065)) + ((!g827) & (!g1606) & (g3064) & (g3065)) + ((!g827) & (g1606) & (g3064) & (!g3065)) + ((!g827) & (g1606) & (g3064) & (g3065)) + ((g827) & (!g1606) & (!g3064) & (!g3065)) + ((g827) & (!g1606) & (g3064) & (g3065)) + ((g827) & (g1606) & (!g3064) & (g3065)) + ((g827) & (g1606) & (g3064) & (!g3065)));
	assign g8187 = (((!g2017) & (g5274) & (!g3067)) + ((!g2017) & (g5274) & (g3067)) + ((g2017) & (!g5274) & (g3067)) + ((g2017) & (g5274) & (g3067)));
	assign g3068 = (((!g1538) & (!g1575) & (!g2991) & (!g3022) & (!g2993) & (!g2994)) + ((!g1538) & (!g1575) & (!g2991) & (!g3022) & (!g2993) & (g2994)) + ((!g1538) & (!g1575) & (!g2991) & (!g3022) & (g2993) & (!g2994)) + ((!g1538) & (!g1575) & (!g2991) & (!g3022) & (g2993) & (g2994)) + ((!g1538) & (!g1575) & (!g2991) & (g3022) & (!g2993) & (!g2994)) + ((!g1538) & (!g1575) & (!g2991) & (g3022) & (!g2993) & (g2994)) + ((!g1538) & (!g1575) & (!g2991) & (g3022) & (g2993) & (!g2994)) + ((!g1538) & (!g1575) & (!g2991) & (g3022) & (g2993) & (g2994)) + ((!g1538) & (!g1575) & (g2991) & (!g3022) & (!g2993) & (!g2994)) + ((!g1538) & (!g1575) & (g2991) & (!g3022) & (!g2993) & (g2994)) + ((!g1538) & (!g1575) & (g2991) & (!g3022) & (g2993) & (!g2994)) + ((!g1538) & (!g1575) & (g2991) & (!g3022) & (g2993) & (g2994)) + ((!g1538) & (!g1575) & (g2991) & (g3022) & (!g2993) & (!g2994)) + ((!g1538) & (g1575) & (!g2991) & (!g3022) & (!g2993) & (!g2994)) + ((!g1538) & (g1575) & (!g2991) & (!g3022) & (!g2993) & (g2994)) + ((!g1538) & (g1575) & (!g2991) & (!g3022) & (g2993) & (!g2994)) + ((!g1538) & (g1575) & (!g2991) & (!g3022) & (g2993) & (g2994)) + ((!g1538) & (g1575) & (g2991) & (!g3022) & (!g2993) & (!g2994)) + ((g1538) & (!g1575) & (!g2991) & (!g3022) & (!g2993) & (!g2994)) + ((g1538) & (!g1575) & (!g2991) & (!g3022) & (!g2993) & (g2994)) + ((g1538) & (!g1575) & (!g2991) & (!g3022) & (g2993) & (!g2994)) + ((g1538) & (!g1575) & (!g2991) & (!g3022) & (g2993) & (g2994)) + ((g1538) & (!g1575) & (!g2991) & (g3022) & (!g2993) & (!g2994)) + ((g1538) & (!g1575) & (g2991) & (!g3022) & (!g2993) & (!g2994)) + ((g1538) & (!g1575) & (g2991) & (!g3022) & (!g2993) & (g2994)) + ((g1538) & (!g1575) & (g2991) & (!g3022) & (g2993) & (!g2994)) + ((g1538) & (!g1575) & (g2991) & (!g3022) & (g2993) & (g2994)) + ((g1538) & (g1575) & (!g2991) & (!g3022) & (!g2993) & (!g2994)));
	assign g3069 = (((!g827) & (!g1608) & (g3067) & (!g3068)) + ((!g827) & (!g1608) & (g3067) & (g3068)) + ((!g827) & (g1608) & (g3067) & (!g3068)) + ((!g827) & (g1608) & (g3067) & (g3068)) + ((g827) & (!g1608) & (!g3067) & (!g3068)) + ((g827) & (!g1608) & (g3067) & (g3068)) + ((g827) & (g1608) & (!g3067) & (g3068)) + ((g827) & (g1608) & (g3067) & (!g3068)));
	assign g3070 = (((!g3024) & (!g1946) & (!g1947) & (!g1948) & (g1949)) + ((!g3024) & (!g1946) & (!g1947) & (g1948) & (!g1949)) + ((!g3024) & (!g1946) & (g1947) & (!g1948) & (g1949)) + ((!g3024) & (!g1946) & (g1947) & (g1948) & (!g1949)) + ((!g3024) & (g1946) & (!g1947) & (!g1948) & (g1949)) + ((!g3024) & (g1946) & (!g1947) & (g1948) & (!g1949)) + ((!g3024) & (g1946) & (g1947) & (!g1948) & (!g1949)) + ((!g3024) & (g1946) & (g1947) & (g1948) & (g1949)) + ((g3024) & (!g1946) & (!g1947) & (!g1948) & (g1949)) + ((g3024) & (!g1946) & (!g1947) & (g1948) & (!g1949)) + ((g3024) & (!g1946) & (g1947) & (!g1948) & (!g1949)) + ((g3024) & (!g1946) & (g1947) & (g1948) & (g1949)) + ((g3024) & (g1946) & (!g1947) & (!g1948) & (!g1949)) + ((g3024) & (g1946) & (!g1947) & (g1948) & (g1949)) + ((g3024) & (g1946) & (g1947) & (!g1948) & (!g1949)) + ((g3024) & (g1946) & (g1947) & (g1948) & (g1949)));
	assign g3071 = (((!g3026) & (!g1984) & (!g1985) & (!g1986) & (g1987)) + ((!g3026) & (!g1984) & (!g1985) & (g1986) & (!g1987)) + ((!g3026) & (!g1984) & (g1985) & (!g1986) & (g1987)) + ((!g3026) & (!g1984) & (g1985) & (g1986) & (!g1987)) + ((!g3026) & (g1984) & (!g1985) & (!g1986) & (g1987)) + ((!g3026) & (g1984) & (!g1985) & (g1986) & (!g1987)) + ((!g3026) & (g1984) & (g1985) & (!g1986) & (!g1987)) + ((!g3026) & (g1984) & (g1985) & (g1986) & (g1987)) + ((g3026) & (!g1984) & (!g1985) & (!g1986) & (g1987)) + ((g3026) & (!g1984) & (!g1985) & (g1986) & (!g1987)) + ((g3026) & (!g1984) & (g1985) & (!g1986) & (!g1987)) + ((g3026) & (!g1984) & (g1985) & (g1986) & (g1987)) + ((g3026) & (g1984) & (!g1985) & (!g1986) & (!g1987)) + ((g3026) & (g1984) & (!g1985) & (g1986) & (g1987)) + ((g3026) & (g1984) & (g1985) & (!g1986) & (!g1987)) + ((g3026) & (g1984) & (g1985) & (g1986) & (g1987)));
	assign g3072 = (((g830) & (!g1914) & (!g3070) & (!g3071) & (g1610)) + ((g830) & (!g1914) & (!g3070) & (g3071) & (!g1610)) + ((g830) & (!g1914) & (g3070) & (!g3071) & (g1610)) + ((g830) & (!g1914) & (g3070) & (g3071) & (!g1610)) + ((g830) & (g1914) & (!g3070) & (!g3071) & (g1610)) + ((g830) & (g1914) & (!g3070) & (g3071) & (g1610)) + ((g830) & (g1914) & (g3070) & (!g3071) & (!g1610)) + ((g830) & (g1914) & (g3070) & (g3071) & (!g1610)));
	assign g3073 = (((!g827) & (!g1586) & (!g1614) & (!g2378) & (g2426) & (!g3036)) + ((!g827) & (!g1586) & (!g1614) & (!g2378) & (g2426) & (g3036)) + ((!g827) & (!g1586) & (!g1614) & (g2378) & (g2426) & (!g3036)) + ((!g827) & (!g1586) & (!g1614) & (g2378) & (g2426) & (g3036)) + ((!g827) & (!g1586) & (g1614) & (!g2378) & (g2426) & (!g3036)) + ((!g827) & (!g1586) & (g1614) & (!g2378) & (g2426) & (g3036)) + ((!g827) & (!g1586) & (g1614) & (g2378) & (g2426) & (!g3036)) + ((!g827) & (!g1586) & (g1614) & (g2378) & (g2426) & (g3036)) + ((!g827) & (g1586) & (!g1614) & (!g2378) & (g2426) & (!g3036)) + ((!g827) & (g1586) & (!g1614) & (!g2378) & (g2426) & (g3036)) + ((!g827) & (g1586) & (!g1614) & (g2378) & (g2426) & (!g3036)) + ((!g827) & (g1586) & (!g1614) & (g2378) & (g2426) & (g3036)) + ((!g827) & (g1586) & (g1614) & (!g2378) & (g2426) & (!g3036)) + ((!g827) & (g1586) & (g1614) & (!g2378) & (g2426) & (g3036)) + ((!g827) & (g1586) & (g1614) & (g2378) & (g2426) & (!g3036)) + ((!g827) & (g1586) & (g1614) & (g2378) & (g2426) & (g3036)) + ((g827) & (!g1586) & (!g1614) & (!g2378) & (g2426) & (!g3036)) + ((g827) & (!g1586) & (!g1614) & (!g2378) & (g2426) & (g3036)) + ((g827) & (!g1586) & (!g1614) & (g2378) & (!g2426) & (!g3036)) + ((g827) & (!g1586) & (!g1614) & (g2378) & (g2426) & (g3036)) + ((g827) & (!g1586) & (g1614) & (!g2378) & (!g2426) & (!g3036)) + ((g827) & (!g1586) & (g1614) & (!g2378) & (!g2426) & (g3036)) + ((g827) & (!g1586) & (g1614) & (g2378) & (!g2426) & (g3036)) + ((g827) & (!g1586) & (g1614) & (g2378) & (g2426) & (!g3036)) + ((g827) & (g1586) & (!g1614) & (!g2378) & (!g2426) & (!g3036)) + ((g827) & (g1586) & (!g1614) & (!g2378) & (g2426) & (g3036)) + ((g827) & (g1586) & (!g1614) & (g2378) & (!g2426) & (!g3036)) + ((g827) & (g1586) & (!g1614) & (g2378) & (!g2426) & (g3036)) + ((g827) & (g1586) & (g1614) & (!g2378) & (!g2426) & (g3036)) + ((g827) & (g1586) & (g1614) & (!g2378) & (g2426) & (!g3036)) + ((g827) & (g1586) & (g1614) & (g2378) & (g2426) & (!g3036)) + ((g827) & (g1586) & (g1614) & (g2378) & (g2426) & (g3036)));
	assign g8188 = (((!g3464) & (g5277) & (!g3074)) + ((!g3464) & (g5277) & (g3074)) + ((g3464) & (!g5277) & (g3074)) + ((g3464) & (g5277) & (g3074)));
	assign g3075 = (((!g827) & (!g1594) & (!g1616) & (!g3047) & (g3074) & (!g3048)) + ((!g827) & (!g1594) & (!g1616) & (!g3047) & (g3074) & (g3048)) + ((!g827) & (!g1594) & (!g1616) & (g3047) & (g3074) & (!g3048)) + ((!g827) & (!g1594) & (!g1616) & (g3047) & (g3074) & (g3048)) + ((!g827) & (!g1594) & (g1616) & (!g3047) & (g3074) & (!g3048)) + ((!g827) & (!g1594) & (g1616) & (!g3047) & (g3074) & (g3048)) + ((!g827) & (!g1594) & (g1616) & (g3047) & (g3074) & (!g3048)) + ((!g827) & (!g1594) & (g1616) & (g3047) & (g3074) & (g3048)) + ((!g827) & (g1594) & (!g1616) & (!g3047) & (g3074) & (!g3048)) + ((!g827) & (g1594) & (!g1616) & (!g3047) & (g3074) & (g3048)) + ((!g827) & (g1594) & (!g1616) & (g3047) & (g3074) & (!g3048)) + ((!g827) & (g1594) & (!g1616) & (g3047) & (g3074) & (g3048)) + ((!g827) & (g1594) & (g1616) & (!g3047) & (g3074) & (!g3048)) + ((!g827) & (g1594) & (g1616) & (!g3047) & (g3074) & (g3048)) + ((!g827) & (g1594) & (g1616) & (g3047) & (g3074) & (!g3048)) + ((!g827) & (g1594) & (g1616) & (g3047) & (g3074) & (g3048)) + ((g827) & (!g1594) & (!g1616) & (!g3047) & (g3074) & (!g3048)) + ((g827) & (!g1594) & (!g1616) & (!g3047) & (g3074) & (g3048)) + ((g827) & (!g1594) & (!g1616) & (g3047) & (!g3074) & (!g3048)) + ((g827) & (!g1594) & (!g1616) & (g3047) & (g3074) & (g3048)) + ((g827) & (!g1594) & (g1616) & (!g3047) & (!g3074) & (!g3048)) + ((g827) & (!g1594) & (g1616) & (!g3047) & (!g3074) & (g3048)) + ((g827) & (!g1594) & (g1616) & (g3047) & (!g3074) & (g3048)) + ((g827) & (!g1594) & (g1616) & (g3047) & (g3074) & (!g3048)) + ((g827) & (g1594) & (!g1616) & (!g3047) & (!g3074) & (!g3048)) + ((g827) & (g1594) & (!g1616) & (!g3047) & (g3074) & (g3048)) + ((g827) & (g1594) & (!g1616) & (g3047) & (!g3074) & (!g3048)) + ((g827) & (g1594) & (!g1616) & (g3047) & (!g3074) & (g3048)) + ((g827) & (g1594) & (g1616) & (!g3047) & (!g3074) & (g3048)) + ((g827) & (g1594) & (g1616) & (!g3047) & (g3074) & (!g3048)) + ((g827) & (g1594) & (g1616) & (g3047) & (g3074) & (!g3048)) + ((g827) & (g1594) & (g1616) & (g3047) & (g3074) & (g3048)));
	assign g3076 = (((!g827) & (!g1602) & (!g1618) & (!g2379) & (g2427) & (!g3059)) + ((!g827) & (!g1602) & (!g1618) & (!g2379) & (g2427) & (g3059)) + ((!g827) & (!g1602) & (!g1618) & (g2379) & (g2427) & (!g3059)) + ((!g827) & (!g1602) & (!g1618) & (g2379) & (g2427) & (g3059)) + ((!g827) & (!g1602) & (g1618) & (!g2379) & (g2427) & (!g3059)) + ((!g827) & (!g1602) & (g1618) & (!g2379) & (g2427) & (g3059)) + ((!g827) & (!g1602) & (g1618) & (g2379) & (g2427) & (!g3059)) + ((!g827) & (!g1602) & (g1618) & (g2379) & (g2427) & (g3059)) + ((!g827) & (g1602) & (!g1618) & (!g2379) & (g2427) & (!g3059)) + ((!g827) & (g1602) & (!g1618) & (!g2379) & (g2427) & (g3059)) + ((!g827) & (g1602) & (!g1618) & (g2379) & (g2427) & (!g3059)) + ((!g827) & (g1602) & (!g1618) & (g2379) & (g2427) & (g3059)) + ((!g827) & (g1602) & (g1618) & (!g2379) & (g2427) & (!g3059)) + ((!g827) & (g1602) & (g1618) & (!g2379) & (g2427) & (g3059)) + ((!g827) & (g1602) & (g1618) & (g2379) & (g2427) & (!g3059)) + ((!g827) & (g1602) & (g1618) & (g2379) & (g2427) & (g3059)) + ((g827) & (!g1602) & (!g1618) & (!g2379) & (g2427) & (!g3059)) + ((g827) & (!g1602) & (!g1618) & (!g2379) & (g2427) & (g3059)) + ((g827) & (!g1602) & (!g1618) & (g2379) & (!g2427) & (!g3059)) + ((g827) & (!g1602) & (!g1618) & (g2379) & (g2427) & (g3059)) + ((g827) & (!g1602) & (g1618) & (!g2379) & (!g2427) & (!g3059)) + ((g827) & (!g1602) & (g1618) & (!g2379) & (!g2427) & (g3059)) + ((g827) & (!g1602) & (g1618) & (g2379) & (!g2427) & (g3059)) + ((g827) & (!g1602) & (g1618) & (g2379) & (g2427) & (!g3059)) + ((g827) & (g1602) & (!g1618) & (!g2379) & (!g2427) & (!g3059)) + ((g827) & (g1602) & (!g1618) & (!g2379) & (g2427) & (g3059)) + ((g827) & (g1602) & (!g1618) & (g2379) & (!g2427) & (!g3059)) + ((g827) & (g1602) & (!g1618) & (g2379) & (!g2427) & (g3059)) + ((g827) & (g1602) & (g1618) & (!g2379) & (!g2427) & (g3059)) + ((g827) & (g1602) & (g1618) & (!g2379) & (g2427) & (!g3059)) + ((g827) & (g1602) & (g1618) & (g2379) & (g2427) & (!g3059)) + ((g827) & (g1602) & (g1618) & (g2379) & (g2427) & (g3059)));
	assign g3077 = (((!g827) & (!g1580) & (!g1620) & (!g2376) & (g2423) & (!g3029)) + ((!g827) & (!g1580) & (!g1620) & (!g2376) & (g2423) & (g3029)) + ((!g827) & (!g1580) & (!g1620) & (g2376) & (g2423) & (!g3029)) + ((!g827) & (!g1580) & (!g1620) & (g2376) & (g2423) & (g3029)) + ((!g827) & (!g1580) & (g1620) & (!g2376) & (g2423) & (!g3029)) + ((!g827) & (!g1580) & (g1620) & (!g2376) & (g2423) & (g3029)) + ((!g827) & (!g1580) & (g1620) & (g2376) & (g2423) & (!g3029)) + ((!g827) & (!g1580) & (g1620) & (g2376) & (g2423) & (g3029)) + ((!g827) & (g1580) & (!g1620) & (!g2376) & (g2423) & (!g3029)) + ((!g827) & (g1580) & (!g1620) & (!g2376) & (g2423) & (g3029)) + ((!g827) & (g1580) & (!g1620) & (g2376) & (g2423) & (!g3029)) + ((!g827) & (g1580) & (!g1620) & (g2376) & (g2423) & (g3029)) + ((!g827) & (g1580) & (g1620) & (!g2376) & (g2423) & (!g3029)) + ((!g827) & (g1580) & (g1620) & (!g2376) & (g2423) & (g3029)) + ((!g827) & (g1580) & (g1620) & (g2376) & (g2423) & (!g3029)) + ((!g827) & (g1580) & (g1620) & (g2376) & (g2423) & (g3029)) + ((g827) & (!g1580) & (!g1620) & (!g2376) & (g2423) & (!g3029)) + ((g827) & (!g1580) & (!g1620) & (!g2376) & (g2423) & (g3029)) + ((g827) & (!g1580) & (!g1620) & (g2376) & (!g2423) & (!g3029)) + ((g827) & (!g1580) & (!g1620) & (g2376) & (g2423) & (g3029)) + ((g827) & (!g1580) & (g1620) & (!g2376) & (!g2423) & (!g3029)) + ((g827) & (!g1580) & (g1620) & (!g2376) & (!g2423) & (g3029)) + ((g827) & (!g1580) & (g1620) & (g2376) & (!g2423) & (g3029)) + ((g827) & (!g1580) & (g1620) & (g2376) & (g2423) & (!g3029)) + ((g827) & (g1580) & (!g1620) & (!g2376) & (!g2423) & (!g3029)) + ((g827) & (g1580) & (!g1620) & (!g2376) & (g2423) & (g3029)) + ((g827) & (g1580) & (!g1620) & (g2376) & (!g2423) & (!g3029)) + ((g827) & (g1580) & (!g1620) & (g2376) & (!g2423) & (g3029)) + ((g827) & (g1580) & (g1620) & (!g2376) & (!g2423) & (g3029)) + ((g827) & (g1580) & (g1620) & (!g2376) & (g2423) & (!g3029)) + ((g827) & (g1580) & (g1620) & (g2376) & (g2423) & (!g3029)) + ((g827) & (g1580) & (g1620) & (g2376) & (g2423) & (g3029)));
	assign g8189 = (((!g2017) & (g5282) & (!g3078)) + ((!g2017) & (g5282) & (g3078)) + ((g2017) & (!g5282) & (g3078)) + ((g2017) & (g5282) & (g3078)));
	assign g3079 = (((!g827) & (!g1588) & (!g1622) & (!g3038) & (g3078) & (!g3039)) + ((!g827) & (!g1588) & (!g1622) & (!g3038) & (g3078) & (g3039)) + ((!g827) & (!g1588) & (!g1622) & (g3038) & (g3078) & (!g3039)) + ((!g827) & (!g1588) & (!g1622) & (g3038) & (g3078) & (g3039)) + ((!g827) & (!g1588) & (g1622) & (!g3038) & (g3078) & (!g3039)) + ((!g827) & (!g1588) & (g1622) & (!g3038) & (g3078) & (g3039)) + ((!g827) & (!g1588) & (g1622) & (g3038) & (g3078) & (!g3039)) + ((!g827) & (!g1588) & (g1622) & (g3038) & (g3078) & (g3039)) + ((!g827) & (g1588) & (!g1622) & (!g3038) & (g3078) & (!g3039)) + ((!g827) & (g1588) & (!g1622) & (!g3038) & (g3078) & (g3039)) + ((!g827) & (g1588) & (!g1622) & (g3038) & (g3078) & (!g3039)) + ((!g827) & (g1588) & (!g1622) & (g3038) & (g3078) & (g3039)) + ((!g827) & (g1588) & (g1622) & (!g3038) & (g3078) & (!g3039)) + ((!g827) & (g1588) & (g1622) & (!g3038) & (g3078) & (g3039)) + ((!g827) & (g1588) & (g1622) & (g3038) & (g3078) & (!g3039)) + ((!g827) & (g1588) & (g1622) & (g3038) & (g3078) & (g3039)) + ((g827) & (!g1588) & (!g1622) & (!g3038) & (g3078) & (!g3039)) + ((g827) & (!g1588) & (!g1622) & (!g3038) & (g3078) & (g3039)) + ((g827) & (!g1588) & (!g1622) & (g3038) & (!g3078) & (!g3039)) + ((g827) & (!g1588) & (!g1622) & (g3038) & (g3078) & (g3039)) + ((g827) & (!g1588) & (g1622) & (!g3038) & (!g3078) & (!g3039)) + ((g827) & (!g1588) & (g1622) & (!g3038) & (!g3078) & (g3039)) + ((g827) & (!g1588) & (g1622) & (g3038) & (!g3078) & (g3039)) + ((g827) & (!g1588) & (g1622) & (g3038) & (g3078) & (!g3039)) + ((g827) & (g1588) & (!g1622) & (!g3038) & (!g3078) & (!g3039)) + ((g827) & (g1588) & (!g1622) & (!g3038) & (g3078) & (g3039)) + ((g827) & (g1588) & (!g1622) & (g3038) & (!g3078) & (!g3039)) + ((g827) & (g1588) & (!g1622) & (g3038) & (!g3078) & (g3039)) + ((g827) & (g1588) & (g1622) & (!g3038) & (!g3078) & (g3039)) + ((g827) & (g1588) & (g1622) & (!g3038) & (g3078) & (!g3039)) + ((g827) & (g1588) & (g1622) & (g3038) & (g3078) & (!g3039)) + ((g827) & (g1588) & (g1622) & (g3038) & (g3078) & (g3039)));
	assign g8190 = (((!g3499) & (g5285) & (!g3080)) + ((!g3499) & (g5285) & (g3080)) + ((g3499) & (!g5285) & (g3080)) + ((g3499) & (g5285) & (g3080)));
	assign g3081 = (((!g827) & (!g1596) & (!g1624) & (!g3050) & (g3080) & (!g3051)) + ((!g827) & (!g1596) & (!g1624) & (!g3050) & (g3080) & (g3051)) + ((!g827) & (!g1596) & (!g1624) & (g3050) & (g3080) & (!g3051)) + ((!g827) & (!g1596) & (!g1624) & (g3050) & (g3080) & (g3051)) + ((!g827) & (!g1596) & (g1624) & (!g3050) & (g3080) & (!g3051)) + ((!g827) & (!g1596) & (g1624) & (!g3050) & (g3080) & (g3051)) + ((!g827) & (!g1596) & (g1624) & (g3050) & (g3080) & (!g3051)) + ((!g827) & (!g1596) & (g1624) & (g3050) & (g3080) & (g3051)) + ((!g827) & (g1596) & (!g1624) & (!g3050) & (g3080) & (!g3051)) + ((!g827) & (g1596) & (!g1624) & (!g3050) & (g3080) & (g3051)) + ((!g827) & (g1596) & (!g1624) & (g3050) & (g3080) & (!g3051)) + ((!g827) & (g1596) & (!g1624) & (g3050) & (g3080) & (g3051)) + ((!g827) & (g1596) & (g1624) & (!g3050) & (g3080) & (!g3051)) + ((!g827) & (g1596) & (g1624) & (!g3050) & (g3080) & (g3051)) + ((!g827) & (g1596) & (g1624) & (g3050) & (g3080) & (!g3051)) + ((!g827) & (g1596) & (g1624) & (g3050) & (g3080) & (g3051)) + ((g827) & (!g1596) & (!g1624) & (!g3050) & (g3080) & (!g3051)) + ((g827) & (!g1596) & (!g1624) & (!g3050) & (g3080) & (g3051)) + ((g827) & (!g1596) & (!g1624) & (g3050) & (!g3080) & (!g3051)) + ((g827) & (!g1596) & (!g1624) & (g3050) & (g3080) & (g3051)) + ((g827) & (!g1596) & (g1624) & (!g3050) & (!g3080) & (!g3051)) + ((g827) & (!g1596) & (g1624) & (!g3050) & (!g3080) & (g3051)) + ((g827) & (!g1596) & (g1624) & (g3050) & (!g3080) & (g3051)) + ((g827) & (!g1596) & (g1624) & (g3050) & (g3080) & (!g3051)) + ((g827) & (g1596) & (!g1624) & (!g3050) & (!g3080) & (!g3051)) + ((g827) & (g1596) & (!g1624) & (!g3050) & (g3080) & (g3051)) + ((g827) & (g1596) & (!g1624) & (g3050) & (!g3080) & (!g3051)) + ((g827) & (g1596) & (!g1624) & (g3050) & (!g3080) & (g3051)) + ((g827) & (g1596) & (g1624) & (!g3050) & (!g3080) & (g3051)) + ((g827) & (g1596) & (g1624) & (!g3050) & (g3080) & (!g3051)) + ((g827) & (g1596) & (g1624) & (g3050) & (g3080) & (!g3051)) + ((g827) & (g1596) & (g1624) & (g3050) & (g3080) & (g3051)));
	assign g8191 = (((!g3464) & (g5288) & (!g3082)) + ((!g3464) & (g5288) & (g3082)) + ((g3464) & (!g5288) & (g3082)) + ((g3464) & (g5288) & (g3082)));
	assign g3083 = (((!g827) & (!g1604) & (!g1626) & (!g3061) & (g3082) & (!g3062)) + ((!g827) & (!g1604) & (!g1626) & (!g3061) & (g3082) & (g3062)) + ((!g827) & (!g1604) & (!g1626) & (g3061) & (g3082) & (!g3062)) + ((!g827) & (!g1604) & (!g1626) & (g3061) & (g3082) & (g3062)) + ((!g827) & (!g1604) & (g1626) & (!g3061) & (g3082) & (!g3062)) + ((!g827) & (!g1604) & (g1626) & (!g3061) & (g3082) & (g3062)) + ((!g827) & (!g1604) & (g1626) & (g3061) & (g3082) & (!g3062)) + ((!g827) & (!g1604) & (g1626) & (g3061) & (g3082) & (g3062)) + ((!g827) & (g1604) & (!g1626) & (!g3061) & (g3082) & (!g3062)) + ((!g827) & (g1604) & (!g1626) & (!g3061) & (g3082) & (g3062)) + ((!g827) & (g1604) & (!g1626) & (g3061) & (g3082) & (!g3062)) + ((!g827) & (g1604) & (!g1626) & (g3061) & (g3082) & (g3062)) + ((!g827) & (g1604) & (g1626) & (!g3061) & (g3082) & (!g3062)) + ((!g827) & (g1604) & (g1626) & (!g3061) & (g3082) & (g3062)) + ((!g827) & (g1604) & (g1626) & (g3061) & (g3082) & (!g3062)) + ((!g827) & (g1604) & (g1626) & (g3061) & (g3082) & (g3062)) + ((g827) & (!g1604) & (!g1626) & (!g3061) & (g3082) & (!g3062)) + ((g827) & (!g1604) & (!g1626) & (!g3061) & (g3082) & (g3062)) + ((g827) & (!g1604) & (!g1626) & (g3061) & (!g3082) & (!g3062)) + ((g827) & (!g1604) & (!g1626) & (g3061) & (g3082) & (g3062)) + ((g827) & (!g1604) & (g1626) & (!g3061) & (!g3082) & (!g3062)) + ((g827) & (!g1604) & (g1626) & (!g3061) & (!g3082) & (g3062)) + ((g827) & (!g1604) & (g1626) & (g3061) & (!g3082) & (g3062)) + ((g827) & (!g1604) & (g1626) & (g3061) & (g3082) & (!g3062)) + ((g827) & (g1604) & (!g1626) & (!g3061) & (!g3082) & (!g3062)) + ((g827) & (g1604) & (!g1626) & (!g3061) & (g3082) & (g3062)) + ((g827) & (g1604) & (!g1626) & (g3061) & (!g3082) & (!g3062)) + ((g827) & (g1604) & (!g1626) & (g3061) & (!g3082) & (g3062)) + ((g827) & (g1604) & (g1626) & (!g3061) & (!g3082) & (g3062)) + ((g827) & (g1604) & (g1626) & (!g3061) & (g3082) & (!g3062)) + ((g827) & (g1604) & (g1626) & (g3061) & (g3082) & (!g3062)) + ((g827) & (g1604) & (g1626) & (g3061) & (g3082) & (g3062)));
	assign g8192 = (((!g3499) & (g5291) & (!g3084)) + ((!g3499) & (g5291) & (g3084)) + ((g3499) & (!g5291) & (g3084)) + ((g3499) & (g5291) & (g3084)));
	assign g3085 = (((!g827) & (!g1582) & (!g1628) & (!g3031) & (g3084) & (!g3032)) + ((!g827) & (!g1582) & (!g1628) & (!g3031) & (g3084) & (g3032)) + ((!g827) & (!g1582) & (!g1628) & (g3031) & (g3084) & (!g3032)) + ((!g827) & (!g1582) & (!g1628) & (g3031) & (g3084) & (g3032)) + ((!g827) & (!g1582) & (g1628) & (!g3031) & (g3084) & (!g3032)) + ((!g827) & (!g1582) & (g1628) & (!g3031) & (g3084) & (g3032)) + ((!g827) & (!g1582) & (g1628) & (g3031) & (g3084) & (!g3032)) + ((!g827) & (!g1582) & (g1628) & (g3031) & (g3084) & (g3032)) + ((!g827) & (g1582) & (!g1628) & (!g3031) & (g3084) & (!g3032)) + ((!g827) & (g1582) & (!g1628) & (!g3031) & (g3084) & (g3032)) + ((!g827) & (g1582) & (!g1628) & (g3031) & (g3084) & (!g3032)) + ((!g827) & (g1582) & (!g1628) & (g3031) & (g3084) & (g3032)) + ((!g827) & (g1582) & (g1628) & (!g3031) & (g3084) & (!g3032)) + ((!g827) & (g1582) & (g1628) & (!g3031) & (g3084) & (g3032)) + ((!g827) & (g1582) & (g1628) & (g3031) & (g3084) & (!g3032)) + ((!g827) & (g1582) & (g1628) & (g3031) & (g3084) & (g3032)) + ((g827) & (!g1582) & (!g1628) & (!g3031) & (g3084) & (!g3032)) + ((g827) & (!g1582) & (!g1628) & (!g3031) & (g3084) & (g3032)) + ((g827) & (!g1582) & (!g1628) & (g3031) & (!g3084) & (!g3032)) + ((g827) & (!g1582) & (!g1628) & (g3031) & (g3084) & (g3032)) + ((g827) & (!g1582) & (g1628) & (!g3031) & (!g3084) & (!g3032)) + ((g827) & (!g1582) & (g1628) & (!g3031) & (!g3084) & (g3032)) + ((g827) & (!g1582) & (g1628) & (g3031) & (!g3084) & (g3032)) + ((g827) & (!g1582) & (g1628) & (g3031) & (g3084) & (!g3032)) + ((g827) & (g1582) & (!g1628) & (!g3031) & (!g3084) & (!g3032)) + ((g827) & (g1582) & (!g1628) & (!g3031) & (g3084) & (g3032)) + ((g827) & (g1582) & (!g1628) & (g3031) & (!g3084) & (!g3032)) + ((g827) & (g1582) & (!g1628) & (g3031) & (!g3084) & (g3032)) + ((g827) & (g1582) & (g1628) & (!g3031) & (!g3084) & (g3032)) + ((g827) & (g1582) & (g1628) & (!g3031) & (g3084) & (!g3032)) + ((g827) & (g1582) & (g1628) & (g3031) & (g3084) & (!g3032)) + ((g827) & (g1582) & (g1628) & (g3031) & (g3084) & (g3032)));
	assign g8193 = (((!g3464) & (g5295) & (!g3086)) + ((!g3464) & (g5295) & (g3086)) + ((g3464) & (!g5295) & (g3086)) + ((g3464) & (g5295) & (g3086)));
	assign g3087 = (((!g827) & (!g1590) & (!g1630) & (!g3041) & (g3086) & (!g3042)) + ((!g827) & (!g1590) & (!g1630) & (!g3041) & (g3086) & (g3042)) + ((!g827) & (!g1590) & (!g1630) & (g3041) & (g3086) & (!g3042)) + ((!g827) & (!g1590) & (!g1630) & (g3041) & (g3086) & (g3042)) + ((!g827) & (!g1590) & (g1630) & (!g3041) & (g3086) & (!g3042)) + ((!g827) & (!g1590) & (g1630) & (!g3041) & (g3086) & (g3042)) + ((!g827) & (!g1590) & (g1630) & (g3041) & (g3086) & (!g3042)) + ((!g827) & (!g1590) & (g1630) & (g3041) & (g3086) & (g3042)) + ((!g827) & (g1590) & (!g1630) & (!g3041) & (g3086) & (!g3042)) + ((!g827) & (g1590) & (!g1630) & (!g3041) & (g3086) & (g3042)) + ((!g827) & (g1590) & (!g1630) & (g3041) & (g3086) & (!g3042)) + ((!g827) & (g1590) & (!g1630) & (g3041) & (g3086) & (g3042)) + ((!g827) & (g1590) & (g1630) & (!g3041) & (g3086) & (!g3042)) + ((!g827) & (g1590) & (g1630) & (!g3041) & (g3086) & (g3042)) + ((!g827) & (g1590) & (g1630) & (g3041) & (g3086) & (!g3042)) + ((!g827) & (g1590) & (g1630) & (g3041) & (g3086) & (g3042)) + ((g827) & (!g1590) & (!g1630) & (!g3041) & (g3086) & (!g3042)) + ((g827) & (!g1590) & (!g1630) & (!g3041) & (g3086) & (g3042)) + ((g827) & (!g1590) & (!g1630) & (g3041) & (!g3086) & (!g3042)) + ((g827) & (!g1590) & (!g1630) & (g3041) & (g3086) & (g3042)) + ((g827) & (!g1590) & (g1630) & (!g3041) & (!g3086) & (!g3042)) + ((g827) & (!g1590) & (g1630) & (!g3041) & (!g3086) & (g3042)) + ((g827) & (!g1590) & (g1630) & (g3041) & (!g3086) & (g3042)) + ((g827) & (!g1590) & (g1630) & (g3041) & (g3086) & (!g3042)) + ((g827) & (g1590) & (!g1630) & (!g3041) & (!g3086) & (!g3042)) + ((g827) & (g1590) & (!g1630) & (!g3041) & (g3086) & (g3042)) + ((g827) & (g1590) & (!g1630) & (g3041) & (!g3086) & (!g3042)) + ((g827) & (g1590) & (!g1630) & (g3041) & (!g3086) & (g3042)) + ((g827) & (g1590) & (g1630) & (!g3041) & (!g3086) & (g3042)) + ((g827) & (g1590) & (g1630) & (!g3041) & (g3086) & (!g3042)) + ((g827) & (g1590) & (g1630) & (g3041) & (g3086) & (!g3042)) + ((g827) & (g1590) & (g1630) & (g3041) & (g3086) & (g3042)));
	assign g8194 = (((!g2017) & (g5300) & (!g3088)) + ((!g2017) & (g5300) & (g3088)) + ((g2017) & (!g5300) & (g3088)) + ((g2017) & (g5300) & (g3088)));
	assign g3089 = (((!g827) & (!g1598) & (!g1632) & (!g3053) & (g3088) & (!g3054)) + ((!g827) & (!g1598) & (!g1632) & (!g3053) & (g3088) & (g3054)) + ((!g827) & (!g1598) & (!g1632) & (g3053) & (g3088) & (!g3054)) + ((!g827) & (!g1598) & (!g1632) & (g3053) & (g3088) & (g3054)) + ((!g827) & (!g1598) & (g1632) & (!g3053) & (g3088) & (!g3054)) + ((!g827) & (!g1598) & (g1632) & (!g3053) & (g3088) & (g3054)) + ((!g827) & (!g1598) & (g1632) & (g3053) & (g3088) & (!g3054)) + ((!g827) & (!g1598) & (g1632) & (g3053) & (g3088) & (g3054)) + ((!g827) & (g1598) & (!g1632) & (!g3053) & (g3088) & (!g3054)) + ((!g827) & (g1598) & (!g1632) & (!g3053) & (g3088) & (g3054)) + ((!g827) & (g1598) & (!g1632) & (g3053) & (g3088) & (!g3054)) + ((!g827) & (g1598) & (!g1632) & (g3053) & (g3088) & (g3054)) + ((!g827) & (g1598) & (g1632) & (!g3053) & (g3088) & (!g3054)) + ((!g827) & (g1598) & (g1632) & (!g3053) & (g3088) & (g3054)) + ((!g827) & (g1598) & (g1632) & (g3053) & (g3088) & (!g3054)) + ((!g827) & (g1598) & (g1632) & (g3053) & (g3088) & (g3054)) + ((g827) & (!g1598) & (!g1632) & (!g3053) & (g3088) & (!g3054)) + ((g827) & (!g1598) & (!g1632) & (!g3053) & (g3088) & (g3054)) + ((g827) & (!g1598) & (!g1632) & (g3053) & (!g3088) & (!g3054)) + ((g827) & (!g1598) & (!g1632) & (g3053) & (g3088) & (g3054)) + ((g827) & (!g1598) & (g1632) & (!g3053) & (!g3088) & (!g3054)) + ((g827) & (!g1598) & (g1632) & (!g3053) & (!g3088) & (g3054)) + ((g827) & (!g1598) & (g1632) & (g3053) & (!g3088) & (g3054)) + ((g827) & (!g1598) & (g1632) & (g3053) & (g3088) & (!g3054)) + ((g827) & (g1598) & (!g1632) & (!g3053) & (!g3088) & (!g3054)) + ((g827) & (g1598) & (!g1632) & (!g3053) & (g3088) & (g3054)) + ((g827) & (g1598) & (!g1632) & (g3053) & (!g3088) & (!g3054)) + ((g827) & (g1598) & (!g1632) & (g3053) & (!g3088) & (g3054)) + ((g827) & (g1598) & (g1632) & (!g3053) & (!g3088) & (g3054)) + ((g827) & (g1598) & (g1632) & (!g3053) & (g3088) & (!g3054)) + ((g827) & (g1598) & (g1632) & (g3053) & (g3088) & (!g3054)) + ((g827) & (g1598) & (g1632) & (g3053) & (g3088) & (g3054)));
	assign g8195 = (((!g3429) & (g5303) & (!g3090)) + ((!g3429) & (g5303) & (g3090)) + ((g3429) & (!g5303) & (g3090)) + ((g3429) & (g5303) & (g3090)));
	assign g3091 = (((!g827) & (!g1606) & (!g1634) & (!g3064) & (g3090) & (!g3065)) + ((!g827) & (!g1606) & (!g1634) & (!g3064) & (g3090) & (g3065)) + ((!g827) & (!g1606) & (!g1634) & (g3064) & (g3090) & (!g3065)) + ((!g827) & (!g1606) & (!g1634) & (g3064) & (g3090) & (g3065)) + ((!g827) & (!g1606) & (g1634) & (!g3064) & (g3090) & (!g3065)) + ((!g827) & (!g1606) & (g1634) & (!g3064) & (g3090) & (g3065)) + ((!g827) & (!g1606) & (g1634) & (g3064) & (g3090) & (!g3065)) + ((!g827) & (!g1606) & (g1634) & (g3064) & (g3090) & (g3065)) + ((!g827) & (g1606) & (!g1634) & (!g3064) & (g3090) & (!g3065)) + ((!g827) & (g1606) & (!g1634) & (!g3064) & (g3090) & (g3065)) + ((!g827) & (g1606) & (!g1634) & (g3064) & (g3090) & (!g3065)) + ((!g827) & (g1606) & (!g1634) & (g3064) & (g3090) & (g3065)) + ((!g827) & (g1606) & (g1634) & (!g3064) & (g3090) & (!g3065)) + ((!g827) & (g1606) & (g1634) & (!g3064) & (g3090) & (g3065)) + ((!g827) & (g1606) & (g1634) & (g3064) & (g3090) & (!g3065)) + ((!g827) & (g1606) & (g1634) & (g3064) & (g3090) & (g3065)) + ((g827) & (!g1606) & (!g1634) & (!g3064) & (g3090) & (!g3065)) + ((g827) & (!g1606) & (!g1634) & (!g3064) & (g3090) & (g3065)) + ((g827) & (!g1606) & (!g1634) & (g3064) & (!g3090) & (!g3065)) + ((g827) & (!g1606) & (!g1634) & (g3064) & (g3090) & (g3065)) + ((g827) & (!g1606) & (g1634) & (!g3064) & (!g3090) & (!g3065)) + ((g827) & (!g1606) & (g1634) & (!g3064) & (!g3090) & (g3065)) + ((g827) & (!g1606) & (g1634) & (g3064) & (!g3090) & (g3065)) + ((g827) & (!g1606) & (g1634) & (g3064) & (g3090) & (!g3065)) + ((g827) & (g1606) & (!g1634) & (!g3064) & (!g3090) & (!g3065)) + ((g827) & (g1606) & (!g1634) & (!g3064) & (g3090) & (g3065)) + ((g827) & (g1606) & (!g1634) & (g3064) & (!g3090) & (!g3065)) + ((g827) & (g1606) & (!g1634) & (g3064) & (!g3090) & (g3065)) + ((g827) & (g1606) & (g1634) & (!g3064) & (!g3090) & (g3065)) + ((g827) & (g1606) & (g1634) & (!g3064) & (g3090) & (!g3065)) + ((g827) & (g1606) & (g1634) & (g3064) & (g3090) & (!g3065)) + ((g827) & (g1606) & (g1634) & (g3064) & (g3090) & (g3065)));
	assign g3092 = (((!g827) & (!g1584) & (!g1636) & (!g2377) & (g2424) & (!g3034)) + ((!g827) & (!g1584) & (!g1636) & (!g2377) & (g2424) & (g3034)) + ((!g827) & (!g1584) & (!g1636) & (g2377) & (g2424) & (!g3034)) + ((!g827) & (!g1584) & (!g1636) & (g2377) & (g2424) & (g3034)) + ((!g827) & (!g1584) & (g1636) & (!g2377) & (g2424) & (!g3034)) + ((!g827) & (!g1584) & (g1636) & (!g2377) & (g2424) & (g3034)) + ((!g827) & (!g1584) & (g1636) & (g2377) & (g2424) & (!g3034)) + ((!g827) & (!g1584) & (g1636) & (g2377) & (g2424) & (g3034)) + ((!g827) & (g1584) & (!g1636) & (!g2377) & (g2424) & (!g3034)) + ((!g827) & (g1584) & (!g1636) & (!g2377) & (g2424) & (g3034)) + ((!g827) & (g1584) & (!g1636) & (g2377) & (g2424) & (!g3034)) + ((!g827) & (g1584) & (!g1636) & (g2377) & (g2424) & (g3034)) + ((!g827) & (g1584) & (g1636) & (!g2377) & (g2424) & (!g3034)) + ((!g827) & (g1584) & (g1636) & (!g2377) & (g2424) & (g3034)) + ((!g827) & (g1584) & (g1636) & (g2377) & (g2424) & (!g3034)) + ((!g827) & (g1584) & (g1636) & (g2377) & (g2424) & (g3034)) + ((g827) & (!g1584) & (!g1636) & (!g2377) & (g2424) & (!g3034)) + ((g827) & (!g1584) & (!g1636) & (!g2377) & (g2424) & (g3034)) + ((g827) & (!g1584) & (!g1636) & (g2377) & (!g2424) & (!g3034)) + ((g827) & (!g1584) & (!g1636) & (g2377) & (g2424) & (g3034)) + ((g827) & (!g1584) & (g1636) & (!g2377) & (!g2424) & (!g3034)) + ((g827) & (!g1584) & (g1636) & (!g2377) & (!g2424) & (g3034)) + ((g827) & (!g1584) & (g1636) & (g2377) & (!g2424) & (g3034)) + ((g827) & (!g1584) & (g1636) & (g2377) & (g2424) & (!g3034)) + ((g827) & (g1584) & (!g1636) & (!g2377) & (!g2424) & (!g3034)) + ((g827) & (g1584) & (!g1636) & (!g2377) & (g2424) & (g3034)) + ((g827) & (g1584) & (!g1636) & (g2377) & (!g2424) & (!g3034)) + ((g827) & (g1584) & (!g1636) & (g2377) & (!g2424) & (g3034)) + ((g827) & (g1584) & (g1636) & (!g2377) & (!g2424) & (g3034)) + ((g827) & (g1584) & (g1636) & (!g2377) & (g2424) & (!g3034)) + ((g827) & (g1584) & (g1636) & (g2377) & (g2424) & (!g3034)) + ((g827) & (g1584) & (g1636) & (g2377) & (g2424) & (g3034)));
	assign g8196 = (((!g3499) & (g5306) & (!g3093)) + ((!g3499) & (g5306) & (g3093)) + ((g3499) & (!g5306) & (g3093)) + ((g3499) & (g5306) & (g3093)));
	assign g3094 = (((!g827) & (!g1592) & (!g1638) & (!g3044) & (g3093) & (!g3045)) + ((!g827) & (!g1592) & (!g1638) & (!g3044) & (g3093) & (g3045)) + ((!g827) & (!g1592) & (!g1638) & (g3044) & (g3093) & (!g3045)) + ((!g827) & (!g1592) & (!g1638) & (g3044) & (g3093) & (g3045)) + ((!g827) & (!g1592) & (g1638) & (!g3044) & (g3093) & (!g3045)) + ((!g827) & (!g1592) & (g1638) & (!g3044) & (g3093) & (g3045)) + ((!g827) & (!g1592) & (g1638) & (g3044) & (g3093) & (!g3045)) + ((!g827) & (!g1592) & (g1638) & (g3044) & (g3093) & (g3045)) + ((!g827) & (g1592) & (!g1638) & (!g3044) & (g3093) & (!g3045)) + ((!g827) & (g1592) & (!g1638) & (!g3044) & (g3093) & (g3045)) + ((!g827) & (g1592) & (!g1638) & (g3044) & (g3093) & (!g3045)) + ((!g827) & (g1592) & (!g1638) & (g3044) & (g3093) & (g3045)) + ((!g827) & (g1592) & (g1638) & (!g3044) & (g3093) & (!g3045)) + ((!g827) & (g1592) & (g1638) & (!g3044) & (g3093) & (g3045)) + ((!g827) & (g1592) & (g1638) & (g3044) & (g3093) & (!g3045)) + ((!g827) & (g1592) & (g1638) & (g3044) & (g3093) & (g3045)) + ((g827) & (!g1592) & (!g1638) & (!g3044) & (g3093) & (!g3045)) + ((g827) & (!g1592) & (!g1638) & (!g3044) & (g3093) & (g3045)) + ((g827) & (!g1592) & (!g1638) & (g3044) & (!g3093) & (!g3045)) + ((g827) & (!g1592) & (!g1638) & (g3044) & (g3093) & (g3045)) + ((g827) & (!g1592) & (g1638) & (!g3044) & (!g3093) & (!g3045)) + ((g827) & (!g1592) & (g1638) & (!g3044) & (!g3093) & (g3045)) + ((g827) & (!g1592) & (g1638) & (g3044) & (!g3093) & (g3045)) + ((g827) & (!g1592) & (g1638) & (g3044) & (g3093) & (!g3045)) + ((g827) & (g1592) & (!g1638) & (!g3044) & (!g3093) & (!g3045)) + ((g827) & (g1592) & (!g1638) & (!g3044) & (g3093) & (g3045)) + ((g827) & (g1592) & (!g1638) & (g3044) & (!g3093) & (!g3045)) + ((g827) & (g1592) & (!g1638) & (g3044) & (!g3093) & (g3045)) + ((g827) & (g1592) & (g1638) & (!g3044) & (!g3093) & (g3045)) + ((g827) & (g1592) & (g1638) & (!g3044) & (g3093) & (!g3045)) + ((g827) & (g1592) & (g1638) & (g3044) & (g3093) & (!g3045)) + ((g827) & (g1592) & (g1638) & (g3044) & (g3093) & (g3045)));
	assign g8197 = (((!g3429) & (g5309) & (!g3095)) + ((!g3429) & (g5309) & (g3095)) + ((g3429) & (!g5309) & (g3095)) + ((g3429) & (g5309) & (g3095)));
	assign g3096 = (((!g827) & (!g1600) & (!g1640) & (!g3056) & (g3095) & (!g3057)) + ((!g827) & (!g1600) & (!g1640) & (!g3056) & (g3095) & (g3057)) + ((!g827) & (!g1600) & (!g1640) & (g3056) & (g3095) & (!g3057)) + ((!g827) & (!g1600) & (!g1640) & (g3056) & (g3095) & (g3057)) + ((!g827) & (!g1600) & (g1640) & (!g3056) & (g3095) & (!g3057)) + ((!g827) & (!g1600) & (g1640) & (!g3056) & (g3095) & (g3057)) + ((!g827) & (!g1600) & (g1640) & (g3056) & (g3095) & (!g3057)) + ((!g827) & (!g1600) & (g1640) & (g3056) & (g3095) & (g3057)) + ((!g827) & (g1600) & (!g1640) & (!g3056) & (g3095) & (!g3057)) + ((!g827) & (g1600) & (!g1640) & (!g3056) & (g3095) & (g3057)) + ((!g827) & (g1600) & (!g1640) & (g3056) & (g3095) & (!g3057)) + ((!g827) & (g1600) & (!g1640) & (g3056) & (g3095) & (g3057)) + ((!g827) & (g1600) & (g1640) & (!g3056) & (g3095) & (!g3057)) + ((!g827) & (g1600) & (g1640) & (!g3056) & (g3095) & (g3057)) + ((!g827) & (g1600) & (g1640) & (g3056) & (g3095) & (!g3057)) + ((!g827) & (g1600) & (g1640) & (g3056) & (g3095) & (g3057)) + ((g827) & (!g1600) & (!g1640) & (!g3056) & (g3095) & (!g3057)) + ((g827) & (!g1600) & (!g1640) & (!g3056) & (g3095) & (g3057)) + ((g827) & (!g1600) & (!g1640) & (g3056) & (!g3095) & (!g3057)) + ((g827) & (!g1600) & (!g1640) & (g3056) & (g3095) & (g3057)) + ((g827) & (!g1600) & (g1640) & (!g3056) & (!g3095) & (!g3057)) + ((g827) & (!g1600) & (g1640) & (!g3056) & (!g3095) & (g3057)) + ((g827) & (!g1600) & (g1640) & (g3056) & (!g3095) & (g3057)) + ((g827) & (!g1600) & (g1640) & (g3056) & (g3095) & (!g3057)) + ((g827) & (g1600) & (!g1640) & (!g3056) & (!g3095) & (!g3057)) + ((g827) & (g1600) & (!g1640) & (!g3056) & (g3095) & (g3057)) + ((g827) & (g1600) & (!g1640) & (g3056) & (!g3095) & (!g3057)) + ((g827) & (g1600) & (!g1640) & (g3056) & (!g3095) & (g3057)) + ((g827) & (g1600) & (g1640) & (!g3056) & (!g3095) & (g3057)) + ((g827) & (g1600) & (g1640) & (!g3056) & (g3095) & (!g3057)) + ((g827) & (g1600) & (g1640) & (g3056) & (g3095) & (!g3057)) + ((g827) & (g1600) & (g1640) & (g3056) & (g3095) & (g3057)));
	assign g8198 = (((!g2017) & (g5314) & (!g3097)) + ((!g2017) & (g5314) & (g3097)) + ((g2017) & (!g5314) & (g3097)) + ((g2017) & (g5314) & (g3097)));
	assign g3098 = (((!g827) & (!g1608) & (!g1642) & (!g3067) & (g3097) & (!g3068)) + ((!g827) & (!g1608) & (!g1642) & (!g3067) & (g3097) & (g3068)) + ((!g827) & (!g1608) & (!g1642) & (g3067) & (g3097) & (!g3068)) + ((!g827) & (!g1608) & (!g1642) & (g3067) & (g3097) & (g3068)) + ((!g827) & (!g1608) & (g1642) & (!g3067) & (g3097) & (!g3068)) + ((!g827) & (!g1608) & (g1642) & (!g3067) & (g3097) & (g3068)) + ((!g827) & (!g1608) & (g1642) & (g3067) & (g3097) & (!g3068)) + ((!g827) & (!g1608) & (g1642) & (g3067) & (g3097) & (g3068)) + ((!g827) & (g1608) & (!g1642) & (!g3067) & (g3097) & (!g3068)) + ((!g827) & (g1608) & (!g1642) & (!g3067) & (g3097) & (g3068)) + ((!g827) & (g1608) & (!g1642) & (g3067) & (g3097) & (!g3068)) + ((!g827) & (g1608) & (!g1642) & (g3067) & (g3097) & (g3068)) + ((!g827) & (g1608) & (g1642) & (!g3067) & (g3097) & (!g3068)) + ((!g827) & (g1608) & (g1642) & (!g3067) & (g3097) & (g3068)) + ((!g827) & (g1608) & (g1642) & (g3067) & (g3097) & (!g3068)) + ((!g827) & (g1608) & (g1642) & (g3067) & (g3097) & (g3068)) + ((g827) & (!g1608) & (!g1642) & (!g3067) & (g3097) & (!g3068)) + ((g827) & (!g1608) & (!g1642) & (!g3067) & (g3097) & (g3068)) + ((g827) & (!g1608) & (!g1642) & (g3067) & (!g3097) & (!g3068)) + ((g827) & (!g1608) & (!g1642) & (g3067) & (g3097) & (g3068)) + ((g827) & (!g1608) & (g1642) & (!g3067) & (!g3097) & (!g3068)) + ((g827) & (!g1608) & (g1642) & (!g3067) & (!g3097) & (g3068)) + ((g827) & (!g1608) & (g1642) & (g3067) & (!g3097) & (g3068)) + ((g827) & (!g1608) & (g1642) & (g3067) & (g3097) & (!g3068)) + ((g827) & (g1608) & (!g1642) & (!g3067) & (!g3097) & (!g3068)) + ((g827) & (g1608) & (!g1642) & (!g3067) & (g3097) & (g3068)) + ((g827) & (g1608) & (!g1642) & (g3067) & (!g3097) & (!g3068)) + ((g827) & (g1608) & (!g1642) & (g3067) & (!g3097) & (g3068)) + ((g827) & (g1608) & (g1642) & (!g3067) & (!g3097) & (g3068)) + ((g827) & (g1608) & (g1642) & (!g3067) & (g3097) & (!g3068)) + ((g827) & (g1608) & (g1642) & (g3067) & (g3097) & (!g3068)) + ((g827) & (g1608) & (g1642) & (g3067) & (g3097) & (g3068)));
	assign g3099 = (((!g1951) & (!g1952)));
	assign g3100 = (((g1914) & (!g3099) & (!g1953) & (!g1954)) + ((g1914) & (!g3099) & (g1953) & (g1954)) + ((g1914) & (g3099) & (!g1953) & (g1954)) + ((g1914) & (g3099) & (g1953) & (!g1954)));
	assign g3101 = (((!g1989) & (!g1990)));
	assign g3102 = (((!g1914) & (!g3101) & (!g1991) & (!g1992)) + ((!g1914) & (!g3101) & (g1991) & (g1992)) + ((!g1914) & (g3101) & (!g1991) & (g1992)) + ((!g1914) & (g3101) & (g1991) & (!g1992)));
	assign g3103 = (((!g830) & (!g3100) & (!g3102) & (!g1644)) + ((!g830) & (!g3100) & (!g3102) & (g1644)) + ((!g830) & (!g3100) & (g3102) & (!g1644)) + ((!g830) & (!g3100) & (g3102) & (g1644)) + ((!g830) & (g3100) & (!g3102) & (!g1644)) + ((!g830) & (g3100) & (!g3102) & (g1644)) + ((!g830) & (g3100) & (g3102) & (!g1644)) + ((!g830) & (g3100) & (g3102) & (g1644)) + ((g830) & (!g3100) & (!g3102) & (g1644)) + ((g830) & (!g3100) & (g3102) & (!g1644)) + ((g830) & (g3100) & (!g3102) & (!g1644)) + ((g830) & (g3100) & (g3102) & (!g1644)));
	assign g3104 = (((!g1580) & (!g1620) & (g2376) & (g2423) & (!g3029)) + ((!g1580) & (g1620) & (!g2376) & (g2423) & (!g3029)) + ((!g1580) & (g1620) & (!g2376) & (g2423) & (g3029)) + ((!g1580) & (g1620) & (g2376) & (!g2423) & (!g3029)) + ((!g1580) & (g1620) & (g2376) & (g2423) & (!g3029)) + ((!g1580) & (g1620) & (g2376) & (g2423) & (g3029)) + ((g1580) & (!g1620) & (!g2376) & (g2423) & (!g3029)) + ((g1580) & (!g1620) & (g2376) & (g2423) & (!g3029)) + ((g1580) & (!g1620) & (g2376) & (g2423) & (g3029)) + ((g1580) & (g1620) & (!g2376) & (!g2423) & (!g3029)) + ((g1580) & (g1620) & (!g2376) & (g2423) & (!g3029)) + ((g1580) & (g1620) & (!g2376) & (g2423) & (g3029)) + ((g1580) & (g1620) & (g2376) & (!g2423) & (!g3029)) + ((g1580) & (g1620) & (g2376) & (!g2423) & (g3029)) + ((g1580) & (g1620) & (g2376) & (g2423) & (!g3029)) + ((g1580) & (g1620) & (g2376) & (g2423) & (g3029)));
	assign g3105 = (((!g827) & (!g1647) & (g2515) & (!g3104)) + ((!g827) & (!g1647) & (g2515) & (g3104)) + ((!g827) & (g1647) & (g2515) & (!g3104)) + ((!g827) & (g1647) & (g2515) & (g3104)) + ((g827) & (!g1647) & (!g2515) & (g3104)) + ((g827) & (!g1647) & (g2515) & (!g3104)) + ((g827) & (g1647) & (!g2515) & (!g3104)) + ((g827) & (g1647) & (g2515) & (g3104)));
	assign g8199 = (((!g3499) & (g5317) & (!g3106)) + ((!g3499) & (g5317) & (g3106)) + ((g3499) & (!g5317) & (g3106)) + ((g3499) & (g5317) & (g3106)));
	assign g3107 = (((!g1582) & (!g1628) & (g3031) & (g3084) & (!g3032)) + ((!g1582) & (g1628) & (!g3031) & (g3084) & (!g3032)) + ((!g1582) & (g1628) & (!g3031) & (g3084) & (g3032)) + ((!g1582) & (g1628) & (g3031) & (!g3084) & (!g3032)) + ((!g1582) & (g1628) & (g3031) & (g3084) & (!g3032)) + ((!g1582) & (g1628) & (g3031) & (g3084) & (g3032)) + ((g1582) & (!g1628) & (!g3031) & (g3084) & (!g3032)) + ((g1582) & (!g1628) & (g3031) & (g3084) & (!g3032)) + ((g1582) & (!g1628) & (g3031) & (g3084) & (g3032)) + ((g1582) & (g1628) & (!g3031) & (!g3084) & (!g3032)) + ((g1582) & (g1628) & (!g3031) & (g3084) & (!g3032)) + ((g1582) & (g1628) & (!g3031) & (g3084) & (g3032)) + ((g1582) & (g1628) & (g3031) & (!g3084) & (!g3032)) + ((g1582) & (g1628) & (g3031) & (!g3084) & (g3032)) + ((g1582) & (g1628) & (g3031) & (g3084) & (!g3032)) + ((g1582) & (g1628) & (g3031) & (g3084) & (g3032)));
	assign g3108 = (((!g827) & (!g1649) & (g3106) & (!g3107)) + ((!g827) & (!g1649) & (g3106) & (g3107)) + ((!g827) & (g1649) & (g3106) & (!g3107)) + ((!g827) & (g1649) & (g3106) & (g3107)) + ((g827) & (!g1649) & (!g3106) & (g3107)) + ((g827) & (!g1649) & (g3106) & (!g3107)) + ((g827) & (g1649) & (!g3106) & (!g3107)) + ((g827) & (g1649) & (g3106) & (g3107)));
	assign g3109 = (((!g1584) & (!g1636) & (g2377) & (g2424) & (!g3034)) + ((!g1584) & (g1636) & (!g2377) & (g2424) & (!g3034)) + ((!g1584) & (g1636) & (!g2377) & (g2424) & (g3034)) + ((!g1584) & (g1636) & (g2377) & (!g2424) & (!g3034)) + ((!g1584) & (g1636) & (g2377) & (g2424) & (!g3034)) + ((!g1584) & (g1636) & (g2377) & (g2424) & (g3034)) + ((g1584) & (!g1636) & (!g2377) & (g2424) & (!g3034)) + ((g1584) & (!g1636) & (g2377) & (g2424) & (!g3034)) + ((g1584) & (!g1636) & (g2377) & (g2424) & (g3034)) + ((g1584) & (g1636) & (!g2377) & (!g2424) & (!g3034)) + ((g1584) & (g1636) & (!g2377) & (g2424) & (!g3034)) + ((g1584) & (g1636) & (!g2377) & (g2424) & (g3034)) + ((g1584) & (g1636) & (g2377) & (!g2424) & (!g3034)) + ((g1584) & (g1636) & (g2377) & (!g2424) & (g3034)) + ((g1584) & (g1636) & (g2377) & (g2424) & (!g3034)) + ((g1584) & (g1636) & (g2377) & (g2424) & (g3034)));
	assign g3110 = (((!g827) & (!g1651) & (g2516) & (!g3109)) + ((!g827) & (!g1651) & (g2516) & (g3109)) + ((!g827) & (g1651) & (g2516) & (!g3109)) + ((!g827) & (g1651) & (g2516) & (g3109)) + ((g827) & (!g1651) & (!g2516) & (g3109)) + ((g827) & (!g1651) & (g2516) & (!g3109)) + ((g827) & (g1651) & (!g2516) & (!g3109)) + ((g827) & (g1651) & (g2516) & (g3109)));
	assign g3111 = (((!g1586) & (!g1614) & (g2378) & (g2426) & (!g3036)) + ((!g1586) & (g1614) & (!g2378) & (g2426) & (!g3036)) + ((!g1586) & (g1614) & (!g2378) & (g2426) & (g3036)) + ((!g1586) & (g1614) & (g2378) & (!g2426) & (!g3036)) + ((!g1586) & (g1614) & (g2378) & (g2426) & (!g3036)) + ((!g1586) & (g1614) & (g2378) & (g2426) & (g3036)) + ((g1586) & (!g1614) & (!g2378) & (g2426) & (!g3036)) + ((g1586) & (!g1614) & (g2378) & (g2426) & (!g3036)) + ((g1586) & (!g1614) & (g2378) & (g2426) & (g3036)) + ((g1586) & (g1614) & (!g2378) & (!g2426) & (!g3036)) + ((g1586) & (g1614) & (!g2378) & (g2426) & (!g3036)) + ((g1586) & (g1614) & (!g2378) & (g2426) & (g3036)) + ((g1586) & (g1614) & (g2378) & (!g2426) & (!g3036)) + ((g1586) & (g1614) & (g2378) & (!g2426) & (g3036)) + ((g1586) & (g1614) & (g2378) & (g2426) & (!g3036)) + ((g1586) & (g1614) & (g2378) & (g2426) & (g3036)));
	assign g3112 = (((!g827) & (!g1653) & (g2518) & (!g3111)) + ((!g827) & (!g1653) & (g2518) & (g3111)) + ((!g827) & (g1653) & (g2518) & (!g3111)) + ((!g827) & (g1653) & (g2518) & (g3111)) + ((g827) & (!g1653) & (!g2518) & (g3111)) + ((g827) & (!g1653) & (g2518) & (!g3111)) + ((g827) & (g1653) & (!g2518) & (!g3111)) + ((g827) & (g1653) & (g2518) & (g3111)));
	assign g8200 = (((!g2017) & (g5320) & (!g3113)) + ((!g2017) & (g5320) & (g3113)) + ((g2017) & (!g5320) & (g3113)) + ((g2017) & (g5320) & (g3113)));
	assign g3114 = (((!g1588) & (!g1622) & (g3038) & (g3078) & (!g3039)) + ((!g1588) & (g1622) & (!g3038) & (g3078) & (!g3039)) + ((!g1588) & (g1622) & (!g3038) & (g3078) & (g3039)) + ((!g1588) & (g1622) & (g3038) & (!g3078) & (!g3039)) + ((!g1588) & (g1622) & (g3038) & (g3078) & (!g3039)) + ((!g1588) & (g1622) & (g3038) & (g3078) & (g3039)) + ((g1588) & (!g1622) & (!g3038) & (g3078) & (!g3039)) + ((g1588) & (!g1622) & (g3038) & (g3078) & (!g3039)) + ((g1588) & (!g1622) & (g3038) & (g3078) & (g3039)) + ((g1588) & (g1622) & (!g3038) & (!g3078) & (!g3039)) + ((g1588) & (g1622) & (!g3038) & (g3078) & (!g3039)) + ((g1588) & (g1622) & (!g3038) & (g3078) & (g3039)) + ((g1588) & (g1622) & (g3038) & (!g3078) & (!g3039)) + ((g1588) & (g1622) & (g3038) & (!g3078) & (g3039)) + ((g1588) & (g1622) & (g3038) & (g3078) & (!g3039)) + ((g1588) & (g1622) & (g3038) & (g3078) & (g3039)));
	assign g3115 = (((!g827) & (!g1655) & (g3113) & (!g3114)) + ((!g827) & (!g1655) & (g3113) & (g3114)) + ((!g827) & (g1655) & (g3113) & (!g3114)) + ((!g827) & (g1655) & (g3113) & (g3114)) + ((g827) & (!g1655) & (!g3113) & (g3114)) + ((g827) & (!g1655) & (g3113) & (!g3114)) + ((g827) & (g1655) & (!g3113) & (!g3114)) + ((g827) & (g1655) & (g3113) & (g3114)));
	assign g8201 = (((!g3464) & (g5324) & (!g3116)) + ((!g3464) & (g5324) & (g3116)) + ((g3464) & (!g5324) & (g3116)) + ((g3464) & (g5324) & (g3116)));
	assign g3117 = (((!g1590) & (!g1630) & (g3041) & (g3086) & (!g3042)) + ((!g1590) & (g1630) & (!g3041) & (g3086) & (!g3042)) + ((!g1590) & (g1630) & (!g3041) & (g3086) & (g3042)) + ((!g1590) & (g1630) & (g3041) & (!g3086) & (!g3042)) + ((!g1590) & (g1630) & (g3041) & (g3086) & (!g3042)) + ((!g1590) & (g1630) & (g3041) & (g3086) & (g3042)) + ((g1590) & (!g1630) & (!g3041) & (g3086) & (!g3042)) + ((g1590) & (!g1630) & (g3041) & (g3086) & (!g3042)) + ((g1590) & (!g1630) & (g3041) & (g3086) & (g3042)) + ((g1590) & (g1630) & (!g3041) & (!g3086) & (!g3042)) + ((g1590) & (g1630) & (!g3041) & (g3086) & (!g3042)) + ((g1590) & (g1630) & (!g3041) & (g3086) & (g3042)) + ((g1590) & (g1630) & (g3041) & (!g3086) & (!g3042)) + ((g1590) & (g1630) & (g3041) & (!g3086) & (g3042)) + ((g1590) & (g1630) & (g3041) & (g3086) & (!g3042)) + ((g1590) & (g1630) & (g3041) & (g3086) & (g3042)));
	assign g3118 = (((!g827) & (!g1657) & (g3116) & (!g3117)) + ((!g827) & (!g1657) & (g3116) & (g3117)) + ((!g827) & (g1657) & (g3116) & (!g3117)) + ((!g827) & (g1657) & (g3116) & (g3117)) + ((g827) & (!g1657) & (!g3116) & (g3117)) + ((g827) & (!g1657) & (g3116) & (!g3117)) + ((g827) & (g1657) & (!g3116) & (!g3117)) + ((g827) & (g1657) & (g3116) & (g3117)));
	assign g8202 = (((!g3499) & (g5327) & (!g3119)) + ((!g3499) & (g5327) & (g3119)) + ((g3499) & (!g5327) & (g3119)) + ((g3499) & (g5327) & (g3119)));
	assign g3120 = (((!g1592) & (!g1638) & (g3044) & (g3093) & (!g3045)) + ((!g1592) & (g1638) & (!g3044) & (g3093) & (!g3045)) + ((!g1592) & (g1638) & (!g3044) & (g3093) & (g3045)) + ((!g1592) & (g1638) & (g3044) & (!g3093) & (!g3045)) + ((!g1592) & (g1638) & (g3044) & (g3093) & (!g3045)) + ((!g1592) & (g1638) & (g3044) & (g3093) & (g3045)) + ((g1592) & (!g1638) & (!g3044) & (g3093) & (!g3045)) + ((g1592) & (!g1638) & (g3044) & (g3093) & (!g3045)) + ((g1592) & (!g1638) & (g3044) & (g3093) & (g3045)) + ((g1592) & (g1638) & (!g3044) & (!g3093) & (!g3045)) + ((g1592) & (g1638) & (!g3044) & (g3093) & (!g3045)) + ((g1592) & (g1638) & (!g3044) & (g3093) & (g3045)) + ((g1592) & (g1638) & (g3044) & (!g3093) & (!g3045)) + ((g1592) & (g1638) & (g3044) & (!g3093) & (g3045)) + ((g1592) & (g1638) & (g3044) & (g3093) & (!g3045)) + ((g1592) & (g1638) & (g3044) & (g3093) & (g3045)));
	assign g3121 = (((!g827) & (!g1659) & (g3119) & (!g3120)) + ((!g827) & (!g1659) & (g3119) & (g3120)) + ((!g827) & (g1659) & (g3119) & (!g3120)) + ((!g827) & (g1659) & (g3119) & (g3120)) + ((g827) & (!g1659) & (!g3119) & (g3120)) + ((g827) & (!g1659) & (g3119) & (!g3120)) + ((g827) & (g1659) & (!g3119) & (!g3120)) + ((g827) & (g1659) & (g3119) & (g3120)));
	assign g8203 = (((!g3464) & (g5330) & (!g3122)) + ((!g3464) & (g5330) & (g3122)) + ((g3464) & (!g5330) & (g3122)) + ((g3464) & (g5330) & (g3122)));
	assign g3123 = (((!g1594) & (!g1616) & (g3047) & (g3074) & (!g3048)) + ((!g1594) & (g1616) & (!g3047) & (g3074) & (!g3048)) + ((!g1594) & (g1616) & (!g3047) & (g3074) & (g3048)) + ((!g1594) & (g1616) & (g3047) & (!g3074) & (!g3048)) + ((!g1594) & (g1616) & (g3047) & (g3074) & (!g3048)) + ((!g1594) & (g1616) & (g3047) & (g3074) & (g3048)) + ((g1594) & (!g1616) & (!g3047) & (g3074) & (!g3048)) + ((g1594) & (!g1616) & (g3047) & (g3074) & (!g3048)) + ((g1594) & (!g1616) & (g3047) & (g3074) & (g3048)) + ((g1594) & (g1616) & (!g3047) & (!g3074) & (!g3048)) + ((g1594) & (g1616) & (!g3047) & (g3074) & (!g3048)) + ((g1594) & (g1616) & (!g3047) & (g3074) & (g3048)) + ((g1594) & (g1616) & (g3047) & (!g3074) & (!g3048)) + ((g1594) & (g1616) & (g3047) & (!g3074) & (g3048)) + ((g1594) & (g1616) & (g3047) & (g3074) & (!g3048)) + ((g1594) & (g1616) & (g3047) & (g3074) & (g3048)));
	assign g3124 = (((!g827) & (!g1661) & (g3122) & (!g3123)) + ((!g827) & (!g1661) & (g3122) & (g3123)) + ((!g827) & (g1661) & (g3122) & (!g3123)) + ((!g827) & (g1661) & (g3122) & (g3123)) + ((g827) & (!g1661) & (!g3122) & (g3123)) + ((g827) & (!g1661) & (g3122) & (!g3123)) + ((g827) & (g1661) & (!g3122) & (!g3123)) + ((g827) & (g1661) & (g3122) & (g3123)));
	assign g8204 = (((!g3499) & (g5333) & (!g3125)) + ((!g3499) & (g5333) & (g3125)) + ((g3499) & (!g5333) & (g3125)) + ((g3499) & (g5333) & (g3125)));
	assign g3126 = (((!g1596) & (!g1624) & (g3050) & (g3080) & (!g3051)) + ((!g1596) & (g1624) & (!g3050) & (g3080) & (!g3051)) + ((!g1596) & (g1624) & (!g3050) & (g3080) & (g3051)) + ((!g1596) & (g1624) & (g3050) & (!g3080) & (!g3051)) + ((!g1596) & (g1624) & (g3050) & (g3080) & (!g3051)) + ((!g1596) & (g1624) & (g3050) & (g3080) & (g3051)) + ((g1596) & (!g1624) & (!g3050) & (g3080) & (!g3051)) + ((g1596) & (!g1624) & (g3050) & (g3080) & (!g3051)) + ((g1596) & (!g1624) & (g3050) & (g3080) & (g3051)) + ((g1596) & (g1624) & (!g3050) & (!g3080) & (!g3051)) + ((g1596) & (g1624) & (!g3050) & (g3080) & (!g3051)) + ((g1596) & (g1624) & (!g3050) & (g3080) & (g3051)) + ((g1596) & (g1624) & (g3050) & (!g3080) & (!g3051)) + ((g1596) & (g1624) & (g3050) & (!g3080) & (g3051)) + ((g1596) & (g1624) & (g3050) & (g3080) & (!g3051)) + ((g1596) & (g1624) & (g3050) & (g3080) & (g3051)));
	assign g3127 = (((!g827) & (!g1663) & (g3125) & (!g3126)) + ((!g827) & (!g1663) & (g3125) & (g3126)) + ((!g827) & (g1663) & (g3125) & (!g3126)) + ((!g827) & (g1663) & (g3125) & (g3126)) + ((g827) & (!g1663) & (!g3125) & (g3126)) + ((g827) & (!g1663) & (g3125) & (!g3126)) + ((g827) & (g1663) & (!g3125) & (!g3126)) + ((g827) & (g1663) & (g3125) & (g3126)));
	assign g8205 = (((!g2017) & (g5336) & (!g3128)) + ((!g2017) & (g5336) & (g3128)) + ((g2017) & (!g5336) & (g3128)) + ((g2017) & (g5336) & (g3128)));
	assign g3129 = (((!g1598) & (!g1632) & (g3053) & (g3088) & (!g3054)) + ((!g1598) & (g1632) & (!g3053) & (g3088) & (!g3054)) + ((!g1598) & (g1632) & (!g3053) & (g3088) & (g3054)) + ((!g1598) & (g1632) & (g3053) & (!g3088) & (!g3054)) + ((!g1598) & (g1632) & (g3053) & (g3088) & (!g3054)) + ((!g1598) & (g1632) & (g3053) & (g3088) & (g3054)) + ((g1598) & (!g1632) & (!g3053) & (g3088) & (!g3054)) + ((g1598) & (!g1632) & (g3053) & (g3088) & (!g3054)) + ((g1598) & (!g1632) & (g3053) & (g3088) & (g3054)) + ((g1598) & (g1632) & (!g3053) & (!g3088) & (!g3054)) + ((g1598) & (g1632) & (!g3053) & (g3088) & (!g3054)) + ((g1598) & (g1632) & (!g3053) & (g3088) & (g3054)) + ((g1598) & (g1632) & (g3053) & (!g3088) & (!g3054)) + ((g1598) & (g1632) & (g3053) & (!g3088) & (g3054)) + ((g1598) & (g1632) & (g3053) & (g3088) & (!g3054)) + ((g1598) & (g1632) & (g3053) & (g3088) & (g3054)));
	assign g3130 = (((!g827) & (!g1665) & (g3128) & (!g3129)) + ((!g827) & (!g1665) & (g3128) & (g3129)) + ((!g827) & (g1665) & (g3128) & (!g3129)) + ((!g827) & (g1665) & (g3128) & (g3129)) + ((g827) & (!g1665) & (!g3128) & (g3129)) + ((g827) & (!g1665) & (g3128) & (!g3129)) + ((g827) & (g1665) & (!g3128) & (!g3129)) + ((g827) & (g1665) & (g3128) & (g3129)));
	assign g8206 = (((!g3429) & (g5341) & (!g3131)) + ((!g3429) & (g5341) & (g3131)) + ((g3429) & (!g5341) & (g3131)) + ((g3429) & (g5341) & (g3131)));
	assign g3132 = (((!g1600) & (!g1640) & (g3056) & (g3095) & (!g3057)) + ((!g1600) & (g1640) & (!g3056) & (g3095) & (!g3057)) + ((!g1600) & (g1640) & (!g3056) & (g3095) & (g3057)) + ((!g1600) & (g1640) & (g3056) & (!g3095) & (!g3057)) + ((!g1600) & (g1640) & (g3056) & (g3095) & (!g3057)) + ((!g1600) & (g1640) & (g3056) & (g3095) & (g3057)) + ((g1600) & (!g1640) & (!g3056) & (g3095) & (!g3057)) + ((g1600) & (!g1640) & (g3056) & (g3095) & (!g3057)) + ((g1600) & (!g1640) & (g3056) & (g3095) & (g3057)) + ((g1600) & (g1640) & (!g3056) & (!g3095) & (!g3057)) + ((g1600) & (g1640) & (!g3056) & (g3095) & (!g3057)) + ((g1600) & (g1640) & (!g3056) & (g3095) & (g3057)) + ((g1600) & (g1640) & (g3056) & (!g3095) & (!g3057)) + ((g1600) & (g1640) & (g3056) & (!g3095) & (g3057)) + ((g1600) & (g1640) & (g3056) & (g3095) & (!g3057)) + ((g1600) & (g1640) & (g3056) & (g3095) & (g3057)));
	assign g3133 = (((!g827) & (!g1667) & (g3131) & (!g3132)) + ((!g827) & (!g1667) & (g3131) & (g3132)) + ((!g827) & (g1667) & (g3131) & (!g3132)) + ((!g827) & (g1667) & (g3131) & (g3132)) + ((g827) & (!g1667) & (!g3131) & (g3132)) + ((g827) & (!g1667) & (g3131) & (!g3132)) + ((g827) & (g1667) & (!g3131) & (!g3132)) + ((g827) & (g1667) & (g3131) & (g3132)));
	assign g3134 = (((!g1602) & (!g1618) & (g2379) & (g2427) & (!g3059)) + ((!g1602) & (g1618) & (!g2379) & (g2427) & (!g3059)) + ((!g1602) & (g1618) & (!g2379) & (g2427) & (g3059)) + ((!g1602) & (g1618) & (g2379) & (!g2427) & (!g3059)) + ((!g1602) & (g1618) & (g2379) & (g2427) & (!g3059)) + ((!g1602) & (g1618) & (g2379) & (g2427) & (g3059)) + ((g1602) & (!g1618) & (!g2379) & (g2427) & (!g3059)) + ((g1602) & (!g1618) & (g2379) & (g2427) & (!g3059)) + ((g1602) & (!g1618) & (g2379) & (g2427) & (g3059)) + ((g1602) & (g1618) & (!g2379) & (!g2427) & (!g3059)) + ((g1602) & (g1618) & (!g2379) & (g2427) & (!g3059)) + ((g1602) & (g1618) & (!g2379) & (g2427) & (g3059)) + ((g1602) & (g1618) & (g2379) & (!g2427) & (!g3059)) + ((g1602) & (g1618) & (g2379) & (!g2427) & (g3059)) + ((g1602) & (g1618) & (g2379) & (g2427) & (!g3059)) + ((g1602) & (g1618) & (g2379) & (g2427) & (g3059)));
	assign g3135 = (((!g827) & (!g1669) & (g2519) & (!g3134)) + ((!g827) & (!g1669) & (g2519) & (g3134)) + ((!g827) & (g1669) & (g2519) & (!g3134)) + ((!g827) & (g1669) & (g2519) & (g3134)) + ((g827) & (!g1669) & (!g2519) & (g3134)) + ((g827) & (!g1669) & (g2519) & (!g3134)) + ((g827) & (g1669) & (!g2519) & (!g3134)) + ((g827) & (g1669) & (g2519) & (g3134)));
	assign g8207 = (((!g3464) & (g5344) & (!g3136)) + ((!g3464) & (g5344) & (g3136)) + ((g3464) & (!g5344) & (g3136)) + ((g3464) & (g5344) & (g3136)));
	assign g3137 = (((!g1604) & (!g1626) & (g3061) & (g3082) & (!g3062)) + ((!g1604) & (g1626) & (!g3061) & (g3082) & (!g3062)) + ((!g1604) & (g1626) & (!g3061) & (g3082) & (g3062)) + ((!g1604) & (g1626) & (g3061) & (!g3082) & (!g3062)) + ((!g1604) & (g1626) & (g3061) & (g3082) & (!g3062)) + ((!g1604) & (g1626) & (g3061) & (g3082) & (g3062)) + ((g1604) & (!g1626) & (!g3061) & (g3082) & (!g3062)) + ((g1604) & (!g1626) & (g3061) & (g3082) & (!g3062)) + ((g1604) & (!g1626) & (g3061) & (g3082) & (g3062)) + ((g1604) & (g1626) & (!g3061) & (!g3082) & (!g3062)) + ((g1604) & (g1626) & (!g3061) & (g3082) & (!g3062)) + ((g1604) & (g1626) & (!g3061) & (g3082) & (g3062)) + ((g1604) & (g1626) & (g3061) & (!g3082) & (!g3062)) + ((g1604) & (g1626) & (g3061) & (!g3082) & (g3062)) + ((g1604) & (g1626) & (g3061) & (g3082) & (!g3062)) + ((g1604) & (g1626) & (g3061) & (g3082) & (g3062)));
	assign g3138 = (((!g827) & (!g1671) & (g3136) & (!g3137)) + ((!g827) & (!g1671) & (g3136) & (g3137)) + ((!g827) & (g1671) & (g3136) & (!g3137)) + ((!g827) & (g1671) & (g3136) & (g3137)) + ((g827) & (!g1671) & (!g3136) & (g3137)) + ((g827) & (!g1671) & (g3136) & (!g3137)) + ((g827) & (g1671) & (!g3136) & (!g3137)) + ((g827) & (g1671) & (g3136) & (g3137)));
	assign g8208 = (((!g3429) & (g5349) & (!g3139)) + ((!g3429) & (g5349) & (g3139)) + ((g3429) & (!g5349) & (g3139)) + ((g3429) & (g5349) & (g3139)));
	assign g3140 = (((!g1606) & (!g1634) & (g3064) & (g3090) & (!g3065)) + ((!g1606) & (g1634) & (!g3064) & (g3090) & (!g3065)) + ((!g1606) & (g1634) & (!g3064) & (g3090) & (g3065)) + ((!g1606) & (g1634) & (g3064) & (!g3090) & (!g3065)) + ((!g1606) & (g1634) & (g3064) & (g3090) & (!g3065)) + ((!g1606) & (g1634) & (g3064) & (g3090) & (g3065)) + ((g1606) & (!g1634) & (!g3064) & (g3090) & (!g3065)) + ((g1606) & (!g1634) & (g3064) & (g3090) & (!g3065)) + ((g1606) & (!g1634) & (g3064) & (g3090) & (g3065)) + ((g1606) & (g1634) & (!g3064) & (!g3090) & (!g3065)) + ((g1606) & (g1634) & (!g3064) & (g3090) & (!g3065)) + ((g1606) & (g1634) & (!g3064) & (g3090) & (g3065)) + ((g1606) & (g1634) & (g3064) & (!g3090) & (!g3065)) + ((g1606) & (g1634) & (g3064) & (!g3090) & (g3065)) + ((g1606) & (g1634) & (g3064) & (g3090) & (!g3065)) + ((g1606) & (g1634) & (g3064) & (g3090) & (g3065)));
	assign g3141 = (((!g827) & (!g1673) & (g3139) & (!g3140)) + ((!g827) & (!g1673) & (g3139) & (g3140)) + ((!g827) & (g1673) & (g3139) & (!g3140)) + ((!g827) & (g1673) & (g3139) & (g3140)) + ((g827) & (!g1673) & (!g3139) & (g3140)) + ((g827) & (!g1673) & (g3139) & (!g3140)) + ((g827) & (g1673) & (!g3139) & (!g3140)) + ((g827) & (g1673) & (g3139) & (g3140)));
	assign g8209 = (((!g2017) & (g5352) & (!g3142)) + ((!g2017) & (g5352) & (g3142)) + ((g2017) & (!g5352) & (g3142)) + ((g2017) & (g5352) & (g3142)));
	assign g3143 = (((!g1608) & (!g1642) & (g3067) & (g3097) & (!g3068)) + ((!g1608) & (g1642) & (!g3067) & (g3097) & (!g3068)) + ((!g1608) & (g1642) & (!g3067) & (g3097) & (g3068)) + ((!g1608) & (g1642) & (g3067) & (!g3097) & (!g3068)) + ((!g1608) & (g1642) & (g3067) & (g3097) & (!g3068)) + ((!g1608) & (g1642) & (g3067) & (g3097) & (g3068)) + ((g1608) & (!g1642) & (!g3067) & (g3097) & (!g3068)) + ((g1608) & (!g1642) & (g3067) & (g3097) & (!g3068)) + ((g1608) & (!g1642) & (g3067) & (g3097) & (g3068)) + ((g1608) & (g1642) & (!g3067) & (!g3097) & (!g3068)) + ((g1608) & (g1642) & (!g3067) & (g3097) & (!g3068)) + ((g1608) & (g1642) & (!g3067) & (g3097) & (g3068)) + ((g1608) & (g1642) & (g3067) & (!g3097) & (!g3068)) + ((g1608) & (g1642) & (g3067) & (!g3097) & (g3068)) + ((g1608) & (g1642) & (g3067) & (g3097) & (!g3068)) + ((g1608) & (g1642) & (g3067) & (g3097) & (g3068)));
	assign g3144 = (((!g827) & (!g1675) & (g3142) & (!g3143)) + ((!g827) & (!g1675) & (g3142) & (g3143)) + ((!g827) & (g1675) & (g3142) & (!g3143)) + ((!g827) & (g1675) & (g3142) & (g3143)) + ((g827) & (!g1675) & (!g3142) & (g3143)) + ((g827) & (!g1675) & (g3142) & (!g3143)) + ((g827) & (g1675) & (!g3142) & (!g3143)) + ((g827) & (g1675) & (g3142) & (g3143)));
	assign g3145 = (((!g3099) & (!g1953) & (!g1954) & (!g1955) & (g1956)) + ((!g3099) & (!g1953) & (!g1954) & (g1955) & (!g1956)) + ((!g3099) & (!g1953) & (g1954) & (!g1955) & (!g1956)) + ((!g3099) & (!g1953) & (g1954) & (g1955) & (g1956)) + ((!g3099) & (g1953) & (!g1954) & (!g1955) & (!g1956)) + ((!g3099) & (g1953) & (!g1954) & (g1955) & (g1956)) + ((!g3099) & (g1953) & (g1954) & (!g1955) & (!g1956)) + ((!g3099) & (g1953) & (g1954) & (g1955) & (g1956)) + ((g3099) & (!g1953) & (!g1954) & (!g1955) & (g1956)) + ((g3099) & (!g1953) & (!g1954) & (g1955) & (!g1956)) + ((g3099) & (!g1953) & (g1954) & (!g1955) & (g1956)) + ((g3099) & (!g1953) & (g1954) & (g1955) & (!g1956)) + ((g3099) & (g1953) & (!g1954) & (!g1955) & (g1956)) + ((g3099) & (g1953) & (!g1954) & (g1955) & (!g1956)) + ((g3099) & (g1953) & (g1954) & (!g1955) & (!g1956)) + ((g3099) & (g1953) & (g1954) & (g1955) & (g1956)));
	assign g3146 = (((!g3101) & (!g1991) & (!g1992) & (!g1993) & (g1994)) + ((!g3101) & (!g1991) & (!g1992) & (g1993) & (!g1994)) + ((!g3101) & (!g1991) & (g1992) & (!g1993) & (!g1994)) + ((!g3101) & (!g1991) & (g1992) & (g1993) & (g1994)) + ((!g3101) & (g1991) & (!g1992) & (!g1993) & (!g1994)) + ((!g3101) & (g1991) & (!g1992) & (g1993) & (g1994)) + ((!g3101) & (g1991) & (g1992) & (!g1993) & (!g1994)) + ((!g3101) & (g1991) & (g1992) & (g1993) & (g1994)) + ((g3101) & (!g1991) & (!g1992) & (!g1993) & (g1994)) + ((g3101) & (!g1991) & (!g1992) & (g1993) & (!g1994)) + ((g3101) & (!g1991) & (g1992) & (!g1993) & (g1994)) + ((g3101) & (!g1991) & (g1992) & (g1993) & (!g1994)) + ((g3101) & (g1991) & (!g1992) & (!g1993) & (g1994)) + ((g3101) & (g1991) & (!g1992) & (g1993) & (!g1994)) + ((g3101) & (g1991) & (g1992) & (!g1993) & (!g1994)) + ((g3101) & (g1991) & (g1992) & (g1993) & (g1994)));
	assign g3147 = (((g830) & (!g1914) & (!g3145) & (!g3146) & (g1677)) + ((g830) & (!g1914) & (!g3145) & (g3146) & (!g1677)) + ((g830) & (!g1914) & (g3145) & (!g3146) & (g1677)) + ((g830) & (!g1914) & (g3145) & (g3146) & (!g1677)) + ((g830) & (g1914) & (!g3145) & (!g3146) & (g1677)) + ((g830) & (g1914) & (!g3145) & (g3146) & (g1677)) + ((g830) & (g1914) & (g3145) & (!g3146) & (!g1677)) + ((g830) & (g1914) & (g3145) & (g3146) & (!g1677)));
	assign g3148 = (((!g827) & (!g1653) & (!g1681) & (!g2518) & (g2555) & (!g3111)) + ((!g827) & (!g1653) & (!g1681) & (!g2518) & (g2555) & (g3111)) + ((!g827) & (!g1653) & (!g1681) & (g2518) & (g2555) & (!g3111)) + ((!g827) & (!g1653) & (!g1681) & (g2518) & (g2555) & (g3111)) + ((!g827) & (!g1653) & (g1681) & (!g2518) & (g2555) & (!g3111)) + ((!g827) & (!g1653) & (g1681) & (!g2518) & (g2555) & (g3111)) + ((!g827) & (!g1653) & (g1681) & (g2518) & (g2555) & (!g3111)) + ((!g827) & (!g1653) & (g1681) & (g2518) & (g2555) & (g3111)) + ((!g827) & (g1653) & (!g1681) & (!g2518) & (g2555) & (!g3111)) + ((!g827) & (g1653) & (!g1681) & (!g2518) & (g2555) & (g3111)) + ((!g827) & (g1653) & (!g1681) & (g2518) & (g2555) & (!g3111)) + ((!g827) & (g1653) & (!g1681) & (g2518) & (g2555) & (g3111)) + ((!g827) & (g1653) & (g1681) & (!g2518) & (g2555) & (!g3111)) + ((!g827) & (g1653) & (g1681) & (!g2518) & (g2555) & (g3111)) + ((!g827) & (g1653) & (g1681) & (g2518) & (g2555) & (!g3111)) + ((!g827) & (g1653) & (g1681) & (g2518) & (g2555) & (g3111)) + ((g827) & (!g1653) & (!g1681) & (!g2518) & (g2555) & (!g3111)) + ((g827) & (!g1653) & (!g1681) & (!g2518) & (g2555) & (g3111)) + ((g827) & (!g1653) & (!g1681) & (g2518) & (!g2555) & (g3111)) + ((g827) & (!g1653) & (!g1681) & (g2518) & (g2555) & (!g3111)) + ((g827) & (!g1653) & (g1681) & (!g2518) & (!g2555) & (!g3111)) + ((g827) & (!g1653) & (g1681) & (!g2518) & (!g2555) & (g3111)) + ((g827) & (!g1653) & (g1681) & (g2518) & (!g2555) & (!g3111)) + ((g827) & (!g1653) & (g1681) & (g2518) & (g2555) & (g3111)) + ((g827) & (g1653) & (!g1681) & (!g2518) & (!g2555) & (g3111)) + ((g827) & (g1653) & (!g1681) & (!g2518) & (g2555) & (!g3111)) + ((g827) & (g1653) & (!g1681) & (g2518) & (!g2555) & (!g3111)) + ((g827) & (g1653) & (!g1681) & (g2518) & (!g2555) & (g3111)) + ((g827) & (g1653) & (g1681) & (!g2518) & (!g2555) & (!g3111)) + ((g827) & (g1653) & (g1681) & (!g2518) & (g2555) & (g3111)) + ((g827) & (g1653) & (g1681) & (g2518) & (g2555) & (!g3111)) + ((g827) & (g1653) & (g1681) & (g2518) & (g2555) & (g3111)));
	assign g8210 = (((!g3464) & (g5356) & (!g3149)) + ((!g3464) & (g5356) & (g3149)) + ((g3464) & (!g5356) & (g3149)) + ((g3464) & (g5356) & (g3149)));
	assign g3150 = (((!g827) & (!g1661) & (!g1683) & (!g3122) & (g3149) & (!g3123)) + ((!g827) & (!g1661) & (!g1683) & (!g3122) & (g3149) & (g3123)) + ((!g827) & (!g1661) & (!g1683) & (g3122) & (g3149) & (!g3123)) + ((!g827) & (!g1661) & (!g1683) & (g3122) & (g3149) & (g3123)) + ((!g827) & (!g1661) & (g1683) & (!g3122) & (g3149) & (!g3123)) + ((!g827) & (!g1661) & (g1683) & (!g3122) & (g3149) & (g3123)) + ((!g827) & (!g1661) & (g1683) & (g3122) & (g3149) & (!g3123)) + ((!g827) & (!g1661) & (g1683) & (g3122) & (g3149) & (g3123)) + ((!g827) & (g1661) & (!g1683) & (!g3122) & (g3149) & (!g3123)) + ((!g827) & (g1661) & (!g1683) & (!g3122) & (g3149) & (g3123)) + ((!g827) & (g1661) & (!g1683) & (g3122) & (g3149) & (!g3123)) + ((!g827) & (g1661) & (!g1683) & (g3122) & (g3149) & (g3123)) + ((!g827) & (g1661) & (g1683) & (!g3122) & (g3149) & (!g3123)) + ((!g827) & (g1661) & (g1683) & (!g3122) & (g3149) & (g3123)) + ((!g827) & (g1661) & (g1683) & (g3122) & (g3149) & (!g3123)) + ((!g827) & (g1661) & (g1683) & (g3122) & (g3149) & (g3123)) + ((g827) & (!g1661) & (!g1683) & (!g3122) & (g3149) & (!g3123)) + ((g827) & (!g1661) & (!g1683) & (!g3122) & (g3149) & (g3123)) + ((g827) & (!g1661) & (!g1683) & (g3122) & (!g3149) & (g3123)) + ((g827) & (!g1661) & (!g1683) & (g3122) & (g3149) & (!g3123)) + ((g827) & (!g1661) & (g1683) & (!g3122) & (!g3149) & (!g3123)) + ((g827) & (!g1661) & (g1683) & (!g3122) & (!g3149) & (g3123)) + ((g827) & (!g1661) & (g1683) & (g3122) & (!g3149) & (!g3123)) + ((g827) & (!g1661) & (g1683) & (g3122) & (g3149) & (g3123)) + ((g827) & (g1661) & (!g1683) & (!g3122) & (!g3149) & (g3123)) + ((g827) & (g1661) & (!g1683) & (!g3122) & (g3149) & (!g3123)) + ((g827) & (g1661) & (!g1683) & (g3122) & (!g3149) & (!g3123)) + ((g827) & (g1661) & (!g1683) & (g3122) & (!g3149) & (g3123)) + ((g827) & (g1661) & (g1683) & (!g3122) & (!g3149) & (!g3123)) + ((g827) & (g1661) & (g1683) & (!g3122) & (g3149) & (g3123)) + ((g827) & (g1661) & (g1683) & (g3122) & (g3149) & (!g3123)) + ((g827) & (g1661) & (g1683) & (g3122) & (g3149) & (g3123)));
	assign g3151 = (((!g827) & (!g1669) & (!g1685) & (!g2519) & (g2556) & (!g3134)) + ((!g827) & (!g1669) & (!g1685) & (!g2519) & (g2556) & (g3134)) + ((!g827) & (!g1669) & (!g1685) & (g2519) & (g2556) & (!g3134)) + ((!g827) & (!g1669) & (!g1685) & (g2519) & (g2556) & (g3134)) + ((!g827) & (!g1669) & (g1685) & (!g2519) & (g2556) & (!g3134)) + ((!g827) & (!g1669) & (g1685) & (!g2519) & (g2556) & (g3134)) + ((!g827) & (!g1669) & (g1685) & (g2519) & (g2556) & (!g3134)) + ((!g827) & (!g1669) & (g1685) & (g2519) & (g2556) & (g3134)) + ((!g827) & (g1669) & (!g1685) & (!g2519) & (g2556) & (!g3134)) + ((!g827) & (g1669) & (!g1685) & (!g2519) & (g2556) & (g3134)) + ((!g827) & (g1669) & (!g1685) & (g2519) & (g2556) & (!g3134)) + ((!g827) & (g1669) & (!g1685) & (g2519) & (g2556) & (g3134)) + ((!g827) & (g1669) & (g1685) & (!g2519) & (g2556) & (!g3134)) + ((!g827) & (g1669) & (g1685) & (!g2519) & (g2556) & (g3134)) + ((!g827) & (g1669) & (g1685) & (g2519) & (g2556) & (!g3134)) + ((!g827) & (g1669) & (g1685) & (g2519) & (g2556) & (g3134)) + ((g827) & (!g1669) & (!g1685) & (!g2519) & (g2556) & (!g3134)) + ((g827) & (!g1669) & (!g1685) & (!g2519) & (g2556) & (g3134)) + ((g827) & (!g1669) & (!g1685) & (g2519) & (!g2556) & (g3134)) + ((g827) & (!g1669) & (!g1685) & (g2519) & (g2556) & (!g3134)) + ((g827) & (!g1669) & (g1685) & (!g2519) & (!g2556) & (!g3134)) + ((g827) & (!g1669) & (g1685) & (!g2519) & (!g2556) & (g3134)) + ((g827) & (!g1669) & (g1685) & (g2519) & (!g2556) & (!g3134)) + ((g827) & (!g1669) & (g1685) & (g2519) & (g2556) & (g3134)) + ((g827) & (g1669) & (!g1685) & (!g2519) & (!g2556) & (g3134)) + ((g827) & (g1669) & (!g1685) & (!g2519) & (g2556) & (!g3134)) + ((g827) & (g1669) & (!g1685) & (g2519) & (!g2556) & (!g3134)) + ((g827) & (g1669) & (!g1685) & (g2519) & (!g2556) & (g3134)) + ((g827) & (g1669) & (g1685) & (!g2519) & (!g2556) & (!g3134)) + ((g827) & (g1669) & (g1685) & (!g2519) & (g2556) & (g3134)) + ((g827) & (g1669) & (g1685) & (g2519) & (g2556) & (!g3134)) + ((g827) & (g1669) & (g1685) & (g2519) & (g2556) & (g3134)));
	assign g3152 = (((!g827) & (!g1647) & (!g1687) & (!g2515) & (g2551) & (!g3104)) + ((!g827) & (!g1647) & (!g1687) & (!g2515) & (g2551) & (g3104)) + ((!g827) & (!g1647) & (!g1687) & (g2515) & (g2551) & (!g3104)) + ((!g827) & (!g1647) & (!g1687) & (g2515) & (g2551) & (g3104)) + ((!g827) & (!g1647) & (g1687) & (!g2515) & (g2551) & (!g3104)) + ((!g827) & (!g1647) & (g1687) & (!g2515) & (g2551) & (g3104)) + ((!g827) & (!g1647) & (g1687) & (g2515) & (g2551) & (!g3104)) + ((!g827) & (!g1647) & (g1687) & (g2515) & (g2551) & (g3104)) + ((!g827) & (g1647) & (!g1687) & (!g2515) & (g2551) & (!g3104)) + ((!g827) & (g1647) & (!g1687) & (!g2515) & (g2551) & (g3104)) + ((!g827) & (g1647) & (!g1687) & (g2515) & (g2551) & (!g3104)) + ((!g827) & (g1647) & (!g1687) & (g2515) & (g2551) & (g3104)) + ((!g827) & (g1647) & (g1687) & (!g2515) & (g2551) & (!g3104)) + ((!g827) & (g1647) & (g1687) & (!g2515) & (g2551) & (g3104)) + ((!g827) & (g1647) & (g1687) & (g2515) & (g2551) & (!g3104)) + ((!g827) & (g1647) & (g1687) & (g2515) & (g2551) & (g3104)) + ((g827) & (!g1647) & (!g1687) & (!g2515) & (g2551) & (!g3104)) + ((g827) & (!g1647) & (!g1687) & (!g2515) & (g2551) & (g3104)) + ((g827) & (!g1647) & (!g1687) & (g2515) & (!g2551) & (g3104)) + ((g827) & (!g1647) & (!g1687) & (g2515) & (g2551) & (!g3104)) + ((g827) & (!g1647) & (g1687) & (!g2515) & (!g2551) & (!g3104)) + ((g827) & (!g1647) & (g1687) & (!g2515) & (!g2551) & (g3104)) + ((g827) & (!g1647) & (g1687) & (g2515) & (!g2551) & (!g3104)) + ((g827) & (!g1647) & (g1687) & (g2515) & (g2551) & (g3104)) + ((g827) & (g1647) & (!g1687) & (!g2515) & (!g2551) & (g3104)) + ((g827) & (g1647) & (!g1687) & (!g2515) & (g2551) & (!g3104)) + ((g827) & (g1647) & (!g1687) & (g2515) & (!g2551) & (!g3104)) + ((g827) & (g1647) & (!g1687) & (g2515) & (!g2551) & (g3104)) + ((g827) & (g1647) & (g1687) & (!g2515) & (!g2551) & (!g3104)) + ((g827) & (g1647) & (g1687) & (!g2515) & (g2551) & (g3104)) + ((g827) & (g1647) & (g1687) & (g2515) & (g2551) & (!g3104)) + ((g827) & (g1647) & (g1687) & (g2515) & (g2551) & (g3104)));
	assign g8211 = (((!g2017) & (g6022) & (!g3153)) + ((!g2017) & (g6022) & (g3153)) + ((g2017) & (!g6022) & (g3153)) + ((g2017) & (g6022) & (g3153)));
	assign g3154 = (((!g827) & (!g1655) & (!g1689) & (!g3113) & (g3153) & (!g3114)) + ((!g827) & (!g1655) & (!g1689) & (!g3113) & (g3153) & (g3114)) + ((!g827) & (!g1655) & (!g1689) & (g3113) & (g3153) & (!g3114)) + ((!g827) & (!g1655) & (!g1689) & (g3113) & (g3153) & (g3114)) + ((!g827) & (!g1655) & (g1689) & (!g3113) & (g3153) & (!g3114)) + ((!g827) & (!g1655) & (g1689) & (!g3113) & (g3153) & (g3114)) + ((!g827) & (!g1655) & (g1689) & (g3113) & (g3153) & (!g3114)) + ((!g827) & (!g1655) & (g1689) & (g3113) & (g3153) & (g3114)) + ((!g827) & (g1655) & (!g1689) & (!g3113) & (g3153) & (!g3114)) + ((!g827) & (g1655) & (!g1689) & (!g3113) & (g3153) & (g3114)) + ((!g827) & (g1655) & (!g1689) & (g3113) & (g3153) & (!g3114)) + ((!g827) & (g1655) & (!g1689) & (g3113) & (g3153) & (g3114)) + ((!g827) & (g1655) & (g1689) & (!g3113) & (g3153) & (!g3114)) + ((!g827) & (g1655) & (g1689) & (!g3113) & (g3153) & (g3114)) + ((!g827) & (g1655) & (g1689) & (g3113) & (g3153) & (!g3114)) + ((!g827) & (g1655) & (g1689) & (g3113) & (g3153) & (g3114)) + ((g827) & (!g1655) & (!g1689) & (!g3113) & (g3153) & (!g3114)) + ((g827) & (!g1655) & (!g1689) & (!g3113) & (g3153) & (g3114)) + ((g827) & (!g1655) & (!g1689) & (g3113) & (!g3153) & (g3114)) + ((g827) & (!g1655) & (!g1689) & (g3113) & (g3153) & (!g3114)) + ((g827) & (!g1655) & (g1689) & (!g3113) & (!g3153) & (!g3114)) + ((g827) & (!g1655) & (g1689) & (!g3113) & (!g3153) & (g3114)) + ((g827) & (!g1655) & (g1689) & (g3113) & (!g3153) & (!g3114)) + ((g827) & (!g1655) & (g1689) & (g3113) & (g3153) & (g3114)) + ((g827) & (g1655) & (!g1689) & (!g3113) & (!g3153) & (g3114)) + ((g827) & (g1655) & (!g1689) & (!g3113) & (g3153) & (!g3114)) + ((g827) & (g1655) & (!g1689) & (g3113) & (!g3153) & (!g3114)) + ((g827) & (g1655) & (!g1689) & (g3113) & (!g3153) & (g3114)) + ((g827) & (g1655) & (g1689) & (!g3113) & (!g3153) & (!g3114)) + ((g827) & (g1655) & (g1689) & (!g3113) & (g3153) & (g3114)) + ((g827) & (g1655) & (g1689) & (g3113) & (g3153) & (!g3114)) + ((g827) & (g1655) & (g1689) & (g3113) & (g3153) & (g3114)));
	assign g8212 = (((!g3499) & (g5361) & (!g3155)) + ((!g3499) & (g5361) & (g3155)) + ((g3499) & (!g5361) & (g3155)) + ((g3499) & (g5361) & (g3155)));
	assign g3156 = (((!g827) & (!g1663) & (!g1691) & (!g3125) & (g3155) & (!g3126)) + ((!g827) & (!g1663) & (!g1691) & (!g3125) & (g3155) & (g3126)) + ((!g827) & (!g1663) & (!g1691) & (g3125) & (g3155) & (!g3126)) + ((!g827) & (!g1663) & (!g1691) & (g3125) & (g3155) & (g3126)) + ((!g827) & (!g1663) & (g1691) & (!g3125) & (g3155) & (!g3126)) + ((!g827) & (!g1663) & (g1691) & (!g3125) & (g3155) & (g3126)) + ((!g827) & (!g1663) & (g1691) & (g3125) & (g3155) & (!g3126)) + ((!g827) & (!g1663) & (g1691) & (g3125) & (g3155) & (g3126)) + ((!g827) & (g1663) & (!g1691) & (!g3125) & (g3155) & (!g3126)) + ((!g827) & (g1663) & (!g1691) & (!g3125) & (g3155) & (g3126)) + ((!g827) & (g1663) & (!g1691) & (g3125) & (g3155) & (!g3126)) + ((!g827) & (g1663) & (!g1691) & (g3125) & (g3155) & (g3126)) + ((!g827) & (g1663) & (g1691) & (!g3125) & (g3155) & (!g3126)) + ((!g827) & (g1663) & (g1691) & (!g3125) & (g3155) & (g3126)) + ((!g827) & (g1663) & (g1691) & (g3125) & (g3155) & (!g3126)) + ((!g827) & (g1663) & (g1691) & (g3125) & (g3155) & (g3126)) + ((g827) & (!g1663) & (!g1691) & (!g3125) & (g3155) & (!g3126)) + ((g827) & (!g1663) & (!g1691) & (!g3125) & (g3155) & (g3126)) + ((g827) & (!g1663) & (!g1691) & (g3125) & (!g3155) & (g3126)) + ((g827) & (!g1663) & (!g1691) & (g3125) & (g3155) & (!g3126)) + ((g827) & (!g1663) & (g1691) & (!g3125) & (!g3155) & (!g3126)) + ((g827) & (!g1663) & (g1691) & (!g3125) & (!g3155) & (g3126)) + ((g827) & (!g1663) & (g1691) & (g3125) & (!g3155) & (!g3126)) + ((g827) & (!g1663) & (g1691) & (g3125) & (g3155) & (g3126)) + ((g827) & (g1663) & (!g1691) & (!g3125) & (!g3155) & (g3126)) + ((g827) & (g1663) & (!g1691) & (!g3125) & (g3155) & (!g3126)) + ((g827) & (g1663) & (!g1691) & (g3125) & (!g3155) & (!g3126)) + ((g827) & (g1663) & (!g1691) & (g3125) & (!g3155) & (g3126)) + ((g827) & (g1663) & (g1691) & (!g3125) & (!g3155) & (!g3126)) + ((g827) & (g1663) & (g1691) & (!g3125) & (g3155) & (g3126)) + ((g827) & (g1663) & (g1691) & (g3125) & (g3155) & (!g3126)) + ((g827) & (g1663) & (g1691) & (g3125) & (g3155) & (g3126)));
	assign g8213 = (((!g3464) & (g5365) & (!g3157)) + ((!g3464) & (g5365) & (g3157)) + ((g3464) & (!g5365) & (g3157)) + ((g3464) & (g5365) & (g3157)));
	assign g3158 = (((!g827) & (!g1671) & (!g1693) & (!g3136) & (g3157) & (!g3137)) + ((!g827) & (!g1671) & (!g1693) & (!g3136) & (g3157) & (g3137)) + ((!g827) & (!g1671) & (!g1693) & (g3136) & (g3157) & (!g3137)) + ((!g827) & (!g1671) & (!g1693) & (g3136) & (g3157) & (g3137)) + ((!g827) & (!g1671) & (g1693) & (!g3136) & (g3157) & (!g3137)) + ((!g827) & (!g1671) & (g1693) & (!g3136) & (g3157) & (g3137)) + ((!g827) & (!g1671) & (g1693) & (g3136) & (g3157) & (!g3137)) + ((!g827) & (!g1671) & (g1693) & (g3136) & (g3157) & (g3137)) + ((!g827) & (g1671) & (!g1693) & (!g3136) & (g3157) & (!g3137)) + ((!g827) & (g1671) & (!g1693) & (!g3136) & (g3157) & (g3137)) + ((!g827) & (g1671) & (!g1693) & (g3136) & (g3157) & (!g3137)) + ((!g827) & (g1671) & (!g1693) & (g3136) & (g3157) & (g3137)) + ((!g827) & (g1671) & (g1693) & (!g3136) & (g3157) & (!g3137)) + ((!g827) & (g1671) & (g1693) & (!g3136) & (g3157) & (g3137)) + ((!g827) & (g1671) & (g1693) & (g3136) & (g3157) & (!g3137)) + ((!g827) & (g1671) & (g1693) & (g3136) & (g3157) & (g3137)) + ((g827) & (!g1671) & (!g1693) & (!g3136) & (g3157) & (!g3137)) + ((g827) & (!g1671) & (!g1693) & (!g3136) & (g3157) & (g3137)) + ((g827) & (!g1671) & (!g1693) & (g3136) & (!g3157) & (g3137)) + ((g827) & (!g1671) & (!g1693) & (g3136) & (g3157) & (!g3137)) + ((g827) & (!g1671) & (g1693) & (!g3136) & (!g3157) & (!g3137)) + ((g827) & (!g1671) & (g1693) & (!g3136) & (!g3157) & (g3137)) + ((g827) & (!g1671) & (g1693) & (g3136) & (!g3157) & (!g3137)) + ((g827) & (!g1671) & (g1693) & (g3136) & (g3157) & (g3137)) + ((g827) & (g1671) & (!g1693) & (!g3136) & (!g3157) & (g3137)) + ((g827) & (g1671) & (!g1693) & (!g3136) & (g3157) & (!g3137)) + ((g827) & (g1671) & (!g1693) & (g3136) & (!g3157) & (!g3137)) + ((g827) & (g1671) & (!g1693) & (g3136) & (!g3157) & (g3137)) + ((g827) & (g1671) & (g1693) & (!g3136) & (!g3157) & (!g3137)) + ((g827) & (g1671) & (g1693) & (!g3136) & (g3157) & (g3137)) + ((g827) & (g1671) & (g1693) & (g3136) & (g3157) & (!g3137)) + ((g827) & (g1671) & (g1693) & (g3136) & (g3157) & (g3137)));
	assign g8214 = (((!g3499) & (g5369) & (!g3159)) + ((!g3499) & (g5369) & (g3159)) + ((g3499) & (!g5369) & (g3159)) + ((g3499) & (g5369) & (g3159)));
	assign g3160 = (((!g827) & (!g1649) & (!g1695) & (!g3106) & (g3159) & (!g3107)) + ((!g827) & (!g1649) & (!g1695) & (!g3106) & (g3159) & (g3107)) + ((!g827) & (!g1649) & (!g1695) & (g3106) & (g3159) & (!g3107)) + ((!g827) & (!g1649) & (!g1695) & (g3106) & (g3159) & (g3107)) + ((!g827) & (!g1649) & (g1695) & (!g3106) & (g3159) & (!g3107)) + ((!g827) & (!g1649) & (g1695) & (!g3106) & (g3159) & (g3107)) + ((!g827) & (!g1649) & (g1695) & (g3106) & (g3159) & (!g3107)) + ((!g827) & (!g1649) & (g1695) & (g3106) & (g3159) & (g3107)) + ((!g827) & (g1649) & (!g1695) & (!g3106) & (g3159) & (!g3107)) + ((!g827) & (g1649) & (!g1695) & (!g3106) & (g3159) & (g3107)) + ((!g827) & (g1649) & (!g1695) & (g3106) & (g3159) & (!g3107)) + ((!g827) & (g1649) & (!g1695) & (g3106) & (g3159) & (g3107)) + ((!g827) & (g1649) & (g1695) & (!g3106) & (g3159) & (!g3107)) + ((!g827) & (g1649) & (g1695) & (!g3106) & (g3159) & (g3107)) + ((!g827) & (g1649) & (g1695) & (g3106) & (g3159) & (!g3107)) + ((!g827) & (g1649) & (g1695) & (g3106) & (g3159) & (g3107)) + ((g827) & (!g1649) & (!g1695) & (!g3106) & (g3159) & (!g3107)) + ((g827) & (!g1649) & (!g1695) & (!g3106) & (g3159) & (g3107)) + ((g827) & (!g1649) & (!g1695) & (g3106) & (!g3159) & (g3107)) + ((g827) & (!g1649) & (!g1695) & (g3106) & (g3159) & (!g3107)) + ((g827) & (!g1649) & (g1695) & (!g3106) & (!g3159) & (!g3107)) + ((g827) & (!g1649) & (g1695) & (!g3106) & (!g3159) & (g3107)) + ((g827) & (!g1649) & (g1695) & (g3106) & (!g3159) & (!g3107)) + ((g827) & (!g1649) & (g1695) & (g3106) & (g3159) & (g3107)) + ((g827) & (g1649) & (!g1695) & (!g3106) & (!g3159) & (g3107)) + ((g827) & (g1649) & (!g1695) & (!g3106) & (g3159) & (!g3107)) + ((g827) & (g1649) & (!g1695) & (g3106) & (!g3159) & (!g3107)) + ((g827) & (g1649) & (!g1695) & (g3106) & (!g3159) & (g3107)) + ((g827) & (g1649) & (g1695) & (!g3106) & (!g3159) & (!g3107)) + ((g827) & (g1649) & (g1695) & (!g3106) & (g3159) & (g3107)) + ((g827) & (g1649) & (g1695) & (g3106) & (g3159) & (!g3107)) + ((g827) & (g1649) & (g1695) & (g3106) & (g3159) & (g3107)));
	assign g8215 = (((!g3464) & (g5374) & (!g3161)) + ((!g3464) & (g5374) & (g3161)) + ((g3464) & (!g5374) & (g3161)) + ((g3464) & (g5374) & (g3161)));
	assign g3162 = (((!g827) & (!g1657) & (!g1697) & (!g3116) & (g3161) & (!g3117)) + ((!g827) & (!g1657) & (!g1697) & (!g3116) & (g3161) & (g3117)) + ((!g827) & (!g1657) & (!g1697) & (g3116) & (g3161) & (!g3117)) + ((!g827) & (!g1657) & (!g1697) & (g3116) & (g3161) & (g3117)) + ((!g827) & (!g1657) & (g1697) & (!g3116) & (g3161) & (!g3117)) + ((!g827) & (!g1657) & (g1697) & (!g3116) & (g3161) & (g3117)) + ((!g827) & (!g1657) & (g1697) & (g3116) & (g3161) & (!g3117)) + ((!g827) & (!g1657) & (g1697) & (g3116) & (g3161) & (g3117)) + ((!g827) & (g1657) & (!g1697) & (!g3116) & (g3161) & (!g3117)) + ((!g827) & (g1657) & (!g1697) & (!g3116) & (g3161) & (g3117)) + ((!g827) & (g1657) & (!g1697) & (g3116) & (g3161) & (!g3117)) + ((!g827) & (g1657) & (!g1697) & (g3116) & (g3161) & (g3117)) + ((!g827) & (g1657) & (g1697) & (!g3116) & (g3161) & (!g3117)) + ((!g827) & (g1657) & (g1697) & (!g3116) & (g3161) & (g3117)) + ((!g827) & (g1657) & (g1697) & (g3116) & (g3161) & (!g3117)) + ((!g827) & (g1657) & (g1697) & (g3116) & (g3161) & (g3117)) + ((g827) & (!g1657) & (!g1697) & (!g3116) & (g3161) & (!g3117)) + ((g827) & (!g1657) & (!g1697) & (!g3116) & (g3161) & (g3117)) + ((g827) & (!g1657) & (!g1697) & (g3116) & (!g3161) & (g3117)) + ((g827) & (!g1657) & (!g1697) & (g3116) & (g3161) & (!g3117)) + ((g827) & (!g1657) & (g1697) & (!g3116) & (!g3161) & (!g3117)) + ((g827) & (!g1657) & (g1697) & (!g3116) & (!g3161) & (g3117)) + ((g827) & (!g1657) & (g1697) & (g3116) & (!g3161) & (!g3117)) + ((g827) & (!g1657) & (g1697) & (g3116) & (g3161) & (g3117)) + ((g827) & (g1657) & (!g1697) & (!g3116) & (!g3161) & (g3117)) + ((g827) & (g1657) & (!g1697) & (!g3116) & (g3161) & (!g3117)) + ((g827) & (g1657) & (!g1697) & (g3116) & (!g3161) & (!g3117)) + ((g827) & (g1657) & (!g1697) & (g3116) & (!g3161) & (g3117)) + ((g827) & (g1657) & (g1697) & (!g3116) & (!g3161) & (!g3117)) + ((g827) & (g1657) & (g1697) & (!g3116) & (g3161) & (g3117)) + ((g827) & (g1657) & (g1697) & (g3116) & (g3161) & (!g3117)) + ((g827) & (g1657) & (g1697) & (g3116) & (g3161) & (g3117)));
	assign g8216 = (((!g2017) & (g6016) & (!g3163)) + ((!g2017) & (g6016) & (g3163)) + ((g2017) & (!g6016) & (g3163)) + ((g2017) & (g6016) & (g3163)));
	assign g3164 = (((!g827) & (!g1665) & (!g1699) & (!g3128) & (g3163) & (!g3129)) + ((!g827) & (!g1665) & (!g1699) & (!g3128) & (g3163) & (g3129)) + ((!g827) & (!g1665) & (!g1699) & (g3128) & (g3163) & (!g3129)) + ((!g827) & (!g1665) & (!g1699) & (g3128) & (g3163) & (g3129)) + ((!g827) & (!g1665) & (g1699) & (!g3128) & (g3163) & (!g3129)) + ((!g827) & (!g1665) & (g1699) & (!g3128) & (g3163) & (g3129)) + ((!g827) & (!g1665) & (g1699) & (g3128) & (g3163) & (!g3129)) + ((!g827) & (!g1665) & (g1699) & (g3128) & (g3163) & (g3129)) + ((!g827) & (g1665) & (!g1699) & (!g3128) & (g3163) & (!g3129)) + ((!g827) & (g1665) & (!g1699) & (!g3128) & (g3163) & (g3129)) + ((!g827) & (g1665) & (!g1699) & (g3128) & (g3163) & (!g3129)) + ((!g827) & (g1665) & (!g1699) & (g3128) & (g3163) & (g3129)) + ((!g827) & (g1665) & (g1699) & (!g3128) & (g3163) & (!g3129)) + ((!g827) & (g1665) & (g1699) & (!g3128) & (g3163) & (g3129)) + ((!g827) & (g1665) & (g1699) & (g3128) & (g3163) & (!g3129)) + ((!g827) & (g1665) & (g1699) & (g3128) & (g3163) & (g3129)) + ((g827) & (!g1665) & (!g1699) & (!g3128) & (g3163) & (!g3129)) + ((g827) & (!g1665) & (!g1699) & (!g3128) & (g3163) & (g3129)) + ((g827) & (!g1665) & (!g1699) & (g3128) & (!g3163) & (g3129)) + ((g827) & (!g1665) & (!g1699) & (g3128) & (g3163) & (!g3129)) + ((g827) & (!g1665) & (g1699) & (!g3128) & (!g3163) & (!g3129)) + ((g827) & (!g1665) & (g1699) & (!g3128) & (!g3163) & (g3129)) + ((g827) & (!g1665) & (g1699) & (g3128) & (!g3163) & (!g3129)) + ((g827) & (!g1665) & (g1699) & (g3128) & (g3163) & (g3129)) + ((g827) & (g1665) & (!g1699) & (!g3128) & (!g3163) & (g3129)) + ((g827) & (g1665) & (!g1699) & (!g3128) & (g3163) & (!g3129)) + ((g827) & (g1665) & (!g1699) & (g3128) & (!g3163) & (!g3129)) + ((g827) & (g1665) & (!g1699) & (g3128) & (!g3163) & (g3129)) + ((g827) & (g1665) & (g1699) & (!g3128) & (!g3163) & (!g3129)) + ((g827) & (g1665) & (g1699) & (!g3128) & (g3163) & (g3129)) + ((g827) & (g1665) & (g1699) & (g3128) & (g3163) & (!g3129)) + ((g827) & (g1665) & (g1699) & (g3128) & (g3163) & (g3129)));
	assign g8217 = (((!g3429) & (g5378) & (!g3165)) + ((!g3429) & (g5378) & (g3165)) + ((g3429) & (!g5378) & (g3165)) + ((g3429) & (g5378) & (g3165)));
	assign g3166 = (((!g827) & (!g1673) & (!g1701) & (!g3139) & (g3165) & (!g3140)) + ((!g827) & (!g1673) & (!g1701) & (!g3139) & (g3165) & (g3140)) + ((!g827) & (!g1673) & (!g1701) & (g3139) & (g3165) & (!g3140)) + ((!g827) & (!g1673) & (!g1701) & (g3139) & (g3165) & (g3140)) + ((!g827) & (!g1673) & (g1701) & (!g3139) & (g3165) & (!g3140)) + ((!g827) & (!g1673) & (g1701) & (!g3139) & (g3165) & (g3140)) + ((!g827) & (!g1673) & (g1701) & (g3139) & (g3165) & (!g3140)) + ((!g827) & (!g1673) & (g1701) & (g3139) & (g3165) & (g3140)) + ((!g827) & (g1673) & (!g1701) & (!g3139) & (g3165) & (!g3140)) + ((!g827) & (g1673) & (!g1701) & (!g3139) & (g3165) & (g3140)) + ((!g827) & (g1673) & (!g1701) & (g3139) & (g3165) & (!g3140)) + ((!g827) & (g1673) & (!g1701) & (g3139) & (g3165) & (g3140)) + ((!g827) & (g1673) & (g1701) & (!g3139) & (g3165) & (!g3140)) + ((!g827) & (g1673) & (g1701) & (!g3139) & (g3165) & (g3140)) + ((!g827) & (g1673) & (g1701) & (g3139) & (g3165) & (!g3140)) + ((!g827) & (g1673) & (g1701) & (g3139) & (g3165) & (g3140)) + ((g827) & (!g1673) & (!g1701) & (!g3139) & (g3165) & (!g3140)) + ((g827) & (!g1673) & (!g1701) & (!g3139) & (g3165) & (g3140)) + ((g827) & (!g1673) & (!g1701) & (g3139) & (!g3165) & (g3140)) + ((g827) & (!g1673) & (!g1701) & (g3139) & (g3165) & (!g3140)) + ((g827) & (!g1673) & (g1701) & (!g3139) & (!g3165) & (!g3140)) + ((g827) & (!g1673) & (g1701) & (!g3139) & (!g3165) & (g3140)) + ((g827) & (!g1673) & (g1701) & (g3139) & (!g3165) & (!g3140)) + ((g827) & (!g1673) & (g1701) & (g3139) & (g3165) & (g3140)) + ((g827) & (g1673) & (!g1701) & (!g3139) & (!g3165) & (g3140)) + ((g827) & (g1673) & (!g1701) & (!g3139) & (g3165) & (!g3140)) + ((g827) & (g1673) & (!g1701) & (g3139) & (!g3165) & (!g3140)) + ((g827) & (g1673) & (!g1701) & (g3139) & (!g3165) & (g3140)) + ((g827) & (g1673) & (g1701) & (!g3139) & (!g3165) & (!g3140)) + ((g827) & (g1673) & (g1701) & (!g3139) & (g3165) & (g3140)) + ((g827) & (g1673) & (g1701) & (g3139) & (g3165) & (!g3140)) + ((g827) & (g1673) & (g1701) & (g3139) & (g3165) & (g3140)));
	assign g3167 = (((!g827) & (!g1651) & (!g1703) & (!g2516) & (g2552) & (!g3109)) + ((!g827) & (!g1651) & (!g1703) & (!g2516) & (g2552) & (g3109)) + ((!g827) & (!g1651) & (!g1703) & (g2516) & (g2552) & (!g3109)) + ((!g827) & (!g1651) & (!g1703) & (g2516) & (g2552) & (g3109)) + ((!g827) & (!g1651) & (g1703) & (!g2516) & (g2552) & (!g3109)) + ((!g827) & (!g1651) & (g1703) & (!g2516) & (g2552) & (g3109)) + ((!g827) & (!g1651) & (g1703) & (g2516) & (g2552) & (!g3109)) + ((!g827) & (!g1651) & (g1703) & (g2516) & (g2552) & (g3109)) + ((!g827) & (g1651) & (!g1703) & (!g2516) & (g2552) & (!g3109)) + ((!g827) & (g1651) & (!g1703) & (!g2516) & (g2552) & (g3109)) + ((!g827) & (g1651) & (!g1703) & (g2516) & (g2552) & (!g3109)) + ((!g827) & (g1651) & (!g1703) & (g2516) & (g2552) & (g3109)) + ((!g827) & (g1651) & (g1703) & (!g2516) & (g2552) & (!g3109)) + ((!g827) & (g1651) & (g1703) & (!g2516) & (g2552) & (g3109)) + ((!g827) & (g1651) & (g1703) & (g2516) & (g2552) & (!g3109)) + ((!g827) & (g1651) & (g1703) & (g2516) & (g2552) & (g3109)) + ((g827) & (!g1651) & (!g1703) & (!g2516) & (g2552) & (!g3109)) + ((g827) & (!g1651) & (!g1703) & (!g2516) & (g2552) & (g3109)) + ((g827) & (!g1651) & (!g1703) & (g2516) & (!g2552) & (g3109)) + ((g827) & (!g1651) & (!g1703) & (g2516) & (g2552) & (!g3109)) + ((g827) & (!g1651) & (g1703) & (!g2516) & (!g2552) & (!g3109)) + ((g827) & (!g1651) & (g1703) & (!g2516) & (!g2552) & (g3109)) + ((g827) & (!g1651) & (g1703) & (g2516) & (!g2552) & (!g3109)) + ((g827) & (!g1651) & (g1703) & (g2516) & (g2552) & (g3109)) + ((g827) & (g1651) & (!g1703) & (!g2516) & (!g2552) & (g3109)) + ((g827) & (g1651) & (!g1703) & (!g2516) & (g2552) & (!g3109)) + ((g827) & (g1651) & (!g1703) & (g2516) & (!g2552) & (!g3109)) + ((g827) & (g1651) & (!g1703) & (g2516) & (!g2552) & (g3109)) + ((g827) & (g1651) & (g1703) & (!g2516) & (!g2552) & (!g3109)) + ((g827) & (g1651) & (g1703) & (!g2516) & (g2552) & (g3109)) + ((g827) & (g1651) & (g1703) & (g2516) & (g2552) & (!g3109)) + ((g827) & (g1651) & (g1703) & (g2516) & (g2552) & (g3109)));
	assign g8218 = (((!g3499) & (g5382) & (!g3168)) + ((!g3499) & (g5382) & (g3168)) + ((g3499) & (!g5382) & (g3168)) + ((g3499) & (g5382) & (g3168)));
	assign g3169 = (((!g827) & (!g1659) & (!g1705) & (!g3119) & (g3168) & (!g3120)) + ((!g827) & (!g1659) & (!g1705) & (!g3119) & (g3168) & (g3120)) + ((!g827) & (!g1659) & (!g1705) & (g3119) & (g3168) & (!g3120)) + ((!g827) & (!g1659) & (!g1705) & (g3119) & (g3168) & (g3120)) + ((!g827) & (!g1659) & (g1705) & (!g3119) & (g3168) & (!g3120)) + ((!g827) & (!g1659) & (g1705) & (!g3119) & (g3168) & (g3120)) + ((!g827) & (!g1659) & (g1705) & (g3119) & (g3168) & (!g3120)) + ((!g827) & (!g1659) & (g1705) & (g3119) & (g3168) & (g3120)) + ((!g827) & (g1659) & (!g1705) & (!g3119) & (g3168) & (!g3120)) + ((!g827) & (g1659) & (!g1705) & (!g3119) & (g3168) & (g3120)) + ((!g827) & (g1659) & (!g1705) & (g3119) & (g3168) & (!g3120)) + ((!g827) & (g1659) & (!g1705) & (g3119) & (g3168) & (g3120)) + ((!g827) & (g1659) & (g1705) & (!g3119) & (g3168) & (!g3120)) + ((!g827) & (g1659) & (g1705) & (!g3119) & (g3168) & (g3120)) + ((!g827) & (g1659) & (g1705) & (g3119) & (g3168) & (!g3120)) + ((!g827) & (g1659) & (g1705) & (g3119) & (g3168) & (g3120)) + ((g827) & (!g1659) & (!g1705) & (!g3119) & (g3168) & (!g3120)) + ((g827) & (!g1659) & (!g1705) & (!g3119) & (g3168) & (g3120)) + ((g827) & (!g1659) & (!g1705) & (g3119) & (!g3168) & (g3120)) + ((g827) & (!g1659) & (!g1705) & (g3119) & (g3168) & (!g3120)) + ((g827) & (!g1659) & (g1705) & (!g3119) & (!g3168) & (!g3120)) + ((g827) & (!g1659) & (g1705) & (!g3119) & (!g3168) & (g3120)) + ((g827) & (!g1659) & (g1705) & (g3119) & (!g3168) & (!g3120)) + ((g827) & (!g1659) & (g1705) & (g3119) & (g3168) & (g3120)) + ((g827) & (g1659) & (!g1705) & (!g3119) & (!g3168) & (g3120)) + ((g827) & (g1659) & (!g1705) & (!g3119) & (g3168) & (!g3120)) + ((g827) & (g1659) & (!g1705) & (g3119) & (!g3168) & (!g3120)) + ((g827) & (g1659) & (!g1705) & (g3119) & (!g3168) & (g3120)) + ((g827) & (g1659) & (g1705) & (!g3119) & (!g3168) & (!g3120)) + ((g827) & (g1659) & (g1705) & (!g3119) & (g3168) & (g3120)) + ((g827) & (g1659) & (g1705) & (g3119) & (g3168) & (!g3120)) + ((g827) & (g1659) & (g1705) & (g3119) & (g3168) & (g3120)));
	assign g8219 = (((!g3429) & (g5385) & (!g3170)) + ((!g3429) & (g5385) & (g3170)) + ((g3429) & (!g5385) & (g3170)) + ((g3429) & (g5385) & (g3170)));
	assign g3171 = (((!g827) & (!g1667) & (!g1707) & (!g3131) & (g3170) & (!g3132)) + ((!g827) & (!g1667) & (!g1707) & (!g3131) & (g3170) & (g3132)) + ((!g827) & (!g1667) & (!g1707) & (g3131) & (g3170) & (!g3132)) + ((!g827) & (!g1667) & (!g1707) & (g3131) & (g3170) & (g3132)) + ((!g827) & (!g1667) & (g1707) & (!g3131) & (g3170) & (!g3132)) + ((!g827) & (!g1667) & (g1707) & (!g3131) & (g3170) & (g3132)) + ((!g827) & (!g1667) & (g1707) & (g3131) & (g3170) & (!g3132)) + ((!g827) & (!g1667) & (g1707) & (g3131) & (g3170) & (g3132)) + ((!g827) & (g1667) & (!g1707) & (!g3131) & (g3170) & (!g3132)) + ((!g827) & (g1667) & (!g1707) & (!g3131) & (g3170) & (g3132)) + ((!g827) & (g1667) & (!g1707) & (g3131) & (g3170) & (!g3132)) + ((!g827) & (g1667) & (!g1707) & (g3131) & (g3170) & (g3132)) + ((!g827) & (g1667) & (g1707) & (!g3131) & (g3170) & (!g3132)) + ((!g827) & (g1667) & (g1707) & (!g3131) & (g3170) & (g3132)) + ((!g827) & (g1667) & (g1707) & (g3131) & (g3170) & (!g3132)) + ((!g827) & (g1667) & (g1707) & (g3131) & (g3170) & (g3132)) + ((g827) & (!g1667) & (!g1707) & (!g3131) & (g3170) & (!g3132)) + ((g827) & (!g1667) & (!g1707) & (!g3131) & (g3170) & (g3132)) + ((g827) & (!g1667) & (!g1707) & (g3131) & (!g3170) & (g3132)) + ((g827) & (!g1667) & (!g1707) & (g3131) & (g3170) & (!g3132)) + ((g827) & (!g1667) & (g1707) & (!g3131) & (!g3170) & (!g3132)) + ((g827) & (!g1667) & (g1707) & (!g3131) & (!g3170) & (g3132)) + ((g827) & (!g1667) & (g1707) & (g3131) & (!g3170) & (!g3132)) + ((g827) & (!g1667) & (g1707) & (g3131) & (g3170) & (g3132)) + ((g827) & (g1667) & (!g1707) & (!g3131) & (!g3170) & (g3132)) + ((g827) & (g1667) & (!g1707) & (!g3131) & (g3170) & (!g3132)) + ((g827) & (g1667) & (!g1707) & (g3131) & (!g3170) & (!g3132)) + ((g827) & (g1667) & (!g1707) & (g3131) & (!g3170) & (g3132)) + ((g827) & (g1667) & (g1707) & (!g3131) & (!g3170) & (!g3132)) + ((g827) & (g1667) & (g1707) & (!g3131) & (g3170) & (g3132)) + ((g827) & (g1667) & (g1707) & (g3131) & (g3170) & (!g3132)) + ((g827) & (g1667) & (g1707) & (g3131) & (g3170) & (g3132)));
	assign g8220 = (((!g2017) & (g6010) & (!g3172)) + ((!g2017) & (g6010) & (g3172)) + ((g2017) & (!g6010) & (g3172)) + ((g2017) & (g6010) & (g3172)));
	assign g3173 = (((!g827) & (!g1675) & (!g1709) & (!g3142) & (g3172) & (!g3143)) + ((!g827) & (!g1675) & (!g1709) & (!g3142) & (g3172) & (g3143)) + ((!g827) & (!g1675) & (!g1709) & (g3142) & (g3172) & (!g3143)) + ((!g827) & (!g1675) & (!g1709) & (g3142) & (g3172) & (g3143)) + ((!g827) & (!g1675) & (g1709) & (!g3142) & (g3172) & (!g3143)) + ((!g827) & (!g1675) & (g1709) & (!g3142) & (g3172) & (g3143)) + ((!g827) & (!g1675) & (g1709) & (g3142) & (g3172) & (!g3143)) + ((!g827) & (!g1675) & (g1709) & (g3142) & (g3172) & (g3143)) + ((!g827) & (g1675) & (!g1709) & (!g3142) & (g3172) & (!g3143)) + ((!g827) & (g1675) & (!g1709) & (!g3142) & (g3172) & (g3143)) + ((!g827) & (g1675) & (!g1709) & (g3142) & (g3172) & (!g3143)) + ((!g827) & (g1675) & (!g1709) & (g3142) & (g3172) & (g3143)) + ((!g827) & (g1675) & (g1709) & (!g3142) & (g3172) & (!g3143)) + ((!g827) & (g1675) & (g1709) & (!g3142) & (g3172) & (g3143)) + ((!g827) & (g1675) & (g1709) & (g3142) & (g3172) & (!g3143)) + ((!g827) & (g1675) & (g1709) & (g3142) & (g3172) & (g3143)) + ((g827) & (!g1675) & (!g1709) & (!g3142) & (g3172) & (!g3143)) + ((g827) & (!g1675) & (!g1709) & (!g3142) & (g3172) & (g3143)) + ((g827) & (!g1675) & (!g1709) & (g3142) & (!g3172) & (g3143)) + ((g827) & (!g1675) & (!g1709) & (g3142) & (g3172) & (!g3143)) + ((g827) & (!g1675) & (g1709) & (!g3142) & (!g3172) & (!g3143)) + ((g827) & (!g1675) & (g1709) & (!g3142) & (!g3172) & (g3143)) + ((g827) & (!g1675) & (g1709) & (g3142) & (!g3172) & (!g3143)) + ((g827) & (!g1675) & (g1709) & (g3142) & (g3172) & (g3143)) + ((g827) & (g1675) & (!g1709) & (!g3142) & (!g3172) & (g3143)) + ((g827) & (g1675) & (!g1709) & (!g3142) & (g3172) & (!g3143)) + ((g827) & (g1675) & (!g1709) & (g3142) & (!g3172) & (!g3143)) + ((g827) & (g1675) & (!g1709) & (g3142) & (!g3172) & (g3143)) + ((g827) & (g1675) & (g1709) & (!g3142) & (!g3172) & (!g3143)) + ((g827) & (g1675) & (g1709) & (!g3142) & (g3172) & (g3143)) + ((g827) & (g1675) & (g1709) & (g3142) & (g3172) & (!g3143)) + ((g827) & (g1675) & (g1709) & (g3142) & (g3172) & (g3143)));
	assign g3174 = (((!g1995) & (!g1996) & (!g1997)) + ((!g1995) & (g1996) & (g1997)) + ((g1995) & (!g1996) & (g1997)) + ((g1995) & (g1996) & (!g1997)));
	assign g3175 = (((!g1647) & (!g1687) & (g2515) & (g2551) & (g3104)) + ((!g1647) & (g1687) & (!g2515) & (g2551) & (!g3104)) + ((!g1647) & (g1687) & (!g2515) & (g2551) & (g3104)) + ((!g1647) & (g1687) & (g2515) & (!g2551) & (g3104)) + ((!g1647) & (g1687) & (g2515) & (g2551) & (!g3104)) + ((!g1647) & (g1687) & (g2515) & (g2551) & (g3104)) + ((g1647) & (!g1687) & (!g2515) & (g2551) & (g3104)) + ((g1647) & (!g1687) & (g2515) & (g2551) & (!g3104)) + ((g1647) & (!g1687) & (g2515) & (g2551) & (g3104)) + ((g1647) & (g1687) & (!g2515) & (!g2551) & (g3104)) + ((g1647) & (g1687) & (!g2515) & (g2551) & (!g3104)) + ((g1647) & (g1687) & (!g2515) & (g2551) & (g3104)) + ((g1647) & (g1687) & (g2515) & (!g2551) & (!g3104)) + ((g1647) & (g1687) & (g2515) & (!g2551) & (g3104)) + ((g1647) & (g1687) & (g2515) & (g2551) & (!g3104)) + ((g1647) & (g1687) & (g2515) & (g2551) & (g3104)));
	assign g3176 = (((!g827) & (!g1714) & (g2598) & (!g3175)) + ((!g827) & (!g1714) & (g2598) & (g3175)) + ((!g827) & (g1714) & (g2598) & (!g3175)) + ((!g827) & (g1714) & (g2598) & (g3175)) + ((g827) & (!g1714) & (!g2598) & (g3175)) + ((g827) & (!g1714) & (g2598) & (!g3175)) + ((g827) & (g1714) & (!g2598) & (!g3175)) + ((g827) & (g1714) & (g2598) & (g3175)));
	assign g8221 = (((!g3499) & (g5388) & (!g3177)) + ((!g3499) & (g5388) & (g3177)) + ((g3499) & (!g5388) & (g3177)) + ((g3499) & (g5388) & (g3177)));
	assign g3178 = (((!g1649) & (!g1695) & (g3106) & (g3159) & (g3107)) + ((!g1649) & (g1695) & (!g3106) & (g3159) & (!g3107)) + ((!g1649) & (g1695) & (!g3106) & (g3159) & (g3107)) + ((!g1649) & (g1695) & (g3106) & (!g3159) & (g3107)) + ((!g1649) & (g1695) & (g3106) & (g3159) & (!g3107)) + ((!g1649) & (g1695) & (g3106) & (g3159) & (g3107)) + ((g1649) & (!g1695) & (!g3106) & (g3159) & (g3107)) + ((g1649) & (!g1695) & (g3106) & (g3159) & (!g3107)) + ((g1649) & (!g1695) & (g3106) & (g3159) & (g3107)) + ((g1649) & (g1695) & (!g3106) & (!g3159) & (g3107)) + ((g1649) & (g1695) & (!g3106) & (g3159) & (!g3107)) + ((g1649) & (g1695) & (!g3106) & (g3159) & (g3107)) + ((g1649) & (g1695) & (g3106) & (!g3159) & (!g3107)) + ((g1649) & (g1695) & (g3106) & (!g3159) & (g3107)) + ((g1649) & (g1695) & (g3106) & (g3159) & (!g3107)) + ((g1649) & (g1695) & (g3106) & (g3159) & (g3107)));
	assign g3179 = (((!g827) & (!g1716) & (g3177) & (!g3178)) + ((!g827) & (!g1716) & (g3177) & (g3178)) + ((!g827) & (g1716) & (g3177) & (!g3178)) + ((!g827) & (g1716) & (g3177) & (g3178)) + ((g827) & (!g1716) & (!g3177) & (g3178)) + ((g827) & (!g1716) & (g3177) & (!g3178)) + ((g827) & (g1716) & (!g3177) & (!g3178)) + ((g827) & (g1716) & (g3177) & (g3178)));
	assign g3180 = (((!g1651) & (!g1703) & (g2516) & (g2552) & (g3109)) + ((!g1651) & (g1703) & (!g2516) & (g2552) & (!g3109)) + ((!g1651) & (g1703) & (!g2516) & (g2552) & (g3109)) + ((!g1651) & (g1703) & (g2516) & (!g2552) & (g3109)) + ((!g1651) & (g1703) & (g2516) & (g2552) & (!g3109)) + ((!g1651) & (g1703) & (g2516) & (g2552) & (g3109)) + ((g1651) & (!g1703) & (!g2516) & (g2552) & (g3109)) + ((g1651) & (!g1703) & (g2516) & (g2552) & (!g3109)) + ((g1651) & (!g1703) & (g2516) & (g2552) & (g3109)) + ((g1651) & (g1703) & (!g2516) & (!g2552) & (g3109)) + ((g1651) & (g1703) & (!g2516) & (g2552) & (!g3109)) + ((g1651) & (g1703) & (!g2516) & (g2552) & (g3109)) + ((g1651) & (g1703) & (g2516) & (!g2552) & (!g3109)) + ((g1651) & (g1703) & (g2516) & (!g2552) & (g3109)) + ((g1651) & (g1703) & (g2516) & (g2552) & (!g3109)) + ((g1651) & (g1703) & (g2516) & (g2552) & (g3109)));
	assign g3181 = (((!g827) & (!g1718) & (g2599) & (!g3180)) + ((!g827) & (!g1718) & (g2599) & (g3180)) + ((!g827) & (g1718) & (g2599) & (!g3180)) + ((!g827) & (g1718) & (g2599) & (g3180)) + ((g827) & (!g1718) & (!g2599) & (g3180)) + ((g827) & (!g1718) & (g2599) & (!g3180)) + ((g827) & (g1718) & (!g2599) & (!g3180)) + ((g827) & (g1718) & (g2599) & (g3180)));
	assign g3182 = (((!g1653) & (!g1681) & (g2518) & (g2555) & (g3111)) + ((!g1653) & (g1681) & (!g2518) & (g2555) & (!g3111)) + ((!g1653) & (g1681) & (!g2518) & (g2555) & (g3111)) + ((!g1653) & (g1681) & (g2518) & (!g2555) & (g3111)) + ((!g1653) & (g1681) & (g2518) & (g2555) & (!g3111)) + ((!g1653) & (g1681) & (g2518) & (g2555) & (g3111)) + ((g1653) & (!g1681) & (!g2518) & (g2555) & (g3111)) + ((g1653) & (!g1681) & (g2518) & (g2555) & (!g3111)) + ((g1653) & (!g1681) & (g2518) & (g2555) & (g3111)) + ((g1653) & (g1681) & (!g2518) & (!g2555) & (g3111)) + ((g1653) & (g1681) & (!g2518) & (g2555) & (!g3111)) + ((g1653) & (g1681) & (!g2518) & (g2555) & (g3111)) + ((g1653) & (g1681) & (g2518) & (!g2555) & (!g3111)) + ((g1653) & (g1681) & (g2518) & (!g2555) & (g3111)) + ((g1653) & (g1681) & (g2518) & (g2555) & (!g3111)) + ((g1653) & (g1681) & (g2518) & (g2555) & (g3111)));
	assign g3183 = (((!g827) & (!g1720) & (g2601) & (!g3182)) + ((!g827) & (!g1720) & (g2601) & (g3182)) + ((!g827) & (g1720) & (g2601) & (!g3182)) + ((!g827) & (g1720) & (g2601) & (g3182)) + ((g827) & (!g1720) & (!g2601) & (g3182)) + ((g827) & (!g1720) & (g2601) & (!g3182)) + ((g827) & (g1720) & (!g2601) & (!g3182)) + ((g827) & (g1720) & (g2601) & (g3182)));
	assign g8222 = (((!g2017) & (g5992) & (!g3184)) + ((!g2017) & (g5992) & (g3184)) + ((g2017) & (!g5992) & (g3184)) + ((g2017) & (g5992) & (g3184)));
	assign g3185 = (((!g1655) & (!g1689) & (g3113) & (g3153) & (g3114)) + ((!g1655) & (g1689) & (!g3113) & (g3153) & (!g3114)) + ((!g1655) & (g1689) & (!g3113) & (g3153) & (g3114)) + ((!g1655) & (g1689) & (g3113) & (!g3153) & (g3114)) + ((!g1655) & (g1689) & (g3113) & (g3153) & (!g3114)) + ((!g1655) & (g1689) & (g3113) & (g3153) & (g3114)) + ((g1655) & (!g1689) & (!g3113) & (g3153) & (g3114)) + ((g1655) & (!g1689) & (g3113) & (g3153) & (!g3114)) + ((g1655) & (!g1689) & (g3113) & (g3153) & (g3114)) + ((g1655) & (g1689) & (!g3113) & (!g3153) & (g3114)) + ((g1655) & (g1689) & (!g3113) & (g3153) & (!g3114)) + ((g1655) & (g1689) & (!g3113) & (g3153) & (g3114)) + ((g1655) & (g1689) & (g3113) & (!g3153) & (!g3114)) + ((g1655) & (g1689) & (g3113) & (!g3153) & (g3114)) + ((g1655) & (g1689) & (g3113) & (g3153) & (!g3114)) + ((g1655) & (g1689) & (g3113) & (g3153) & (g3114)));
	assign g3186 = (((!g827) & (!g1722) & (g3184) & (!g3185)) + ((!g827) & (!g1722) & (g3184) & (g3185)) + ((!g827) & (g1722) & (g3184) & (!g3185)) + ((!g827) & (g1722) & (g3184) & (g3185)) + ((g827) & (!g1722) & (!g3184) & (g3185)) + ((g827) & (!g1722) & (g3184) & (!g3185)) + ((g827) & (g1722) & (!g3184) & (!g3185)) + ((g827) & (g1722) & (g3184) & (g3185)));
	assign g8223 = (((!g3464) & (g5394) & (!g3187)) + ((!g3464) & (g5394) & (g3187)) + ((g3464) & (!g5394) & (g3187)) + ((g3464) & (g5394) & (g3187)));
	assign g3188 = (((!g1657) & (!g1697) & (g3116) & (g3161) & (g3117)) + ((!g1657) & (g1697) & (!g3116) & (g3161) & (!g3117)) + ((!g1657) & (g1697) & (!g3116) & (g3161) & (g3117)) + ((!g1657) & (g1697) & (g3116) & (!g3161) & (g3117)) + ((!g1657) & (g1697) & (g3116) & (g3161) & (!g3117)) + ((!g1657) & (g1697) & (g3116) & (g3161) & (g3117)) + ((g1657) & (!g1697) & (!g3116) & (g3161) & (g3117)) + ((g1657) & (!g1697) & (g3116) & (g3161) & (!g3117)) + ((g1657) & (!g1697) & (g3116) & (g3161) & (g3117)) + ((g1657) & (g1697) & (!g3116) & (!g3161) & (g3117)) + ((g1657) & (g1697) & (!g3116) & (g3161) & (!g3117)) + ((g1657) & (g1697) & (!g3116) & (g3161) & (g3117)) + ((g1657) & (g1697) & (g3116) & (!g3161) & (!g3117)) + ((g1657) & (g1697) & (g3116) & (!g3161) & (g3117)) + ((g1657) & (g1697) & (g3116) & (g3161) & (!g3117)) + ((g1657) & (g1697) & (g3116) & (g3161) & (g3117)));
	assign g3189 = (((!g827) & (!g1724) & (g3187) & (!g3188)) + ((!g827) & (!g1724) & (g3187) & (g3188)) + ((!g827) & (g1724) & (g3187) & (!g3188)) + ((!g827) & (g1724) & (g3187) & (g3188)) + ((g827) & (!g1724) & (!g3187) & (g3188)) + ((g827) & (!g1724) & (g3187) & (!g3188)) + ((g827) & (g1724) & (!g3187) & (!g3188)) + ((g827) & (g1724) & (g3187) & (g3188)));
	assign g8224 = (((!g3499) & (g5396) & (!g3190)) + ((!g3499) & (g5396) & (g3190)) + ((g3499) & (!g5396) & (g3190)) + ((g3499) & (g5396) & (g3190)));
	assign g3191 = (((!g1659) & (!g1705) & (g3119) & (g3168) & (g3120)) + ((!g1659) & (g1705) & (!g3119) & (g3168) & (!g3120)) + ((!g1659) & (g1705) & (!g3119) & (g3168) & (g3120)) + ((!g1659) & (g1705) & (g3119) & (!g3168) & (g3120)) + ((!g1659) & (g1705) & (g3119) & (g3168) & (!g3120)) + ((!g1659) & (g1705) & (g3119) & (g3168) & (g3120)) + ((g1659) & (!g1705) & (!g3119) & (g3168) & (g3120)) + ((g1659) & (!g1705) & (g3119) & (g3168) & (!g3120)) + ((g1659) & (!g1705) & (g3119) & (g3168) & (g3120)) + ((g1659) & (g1705) & (!g3119) & (!g3168) & (g3120)) + ((g1659) & (g1705) & (!g3119) & (g3168) & (!g3120)) + ((g1659) & (g1705) & (!g3119) & (g3168) & (g3120)) + ((g1659) & (g1705) & (g3119) & (!g3168) & (!g3120)) + ((g1659) & (g1705) & (g3119) & (!g3168) & (g3120)) + ((g1659) & (g1705) & (g3119) & (g3168) & (!g3120)) + ((g1659) & (g1705) & (g3119) & (g3168) & (g3120)));
	assign g3192 = (((!g827) & (!g1726) & (g3190) & (!g3191)) + ((!g827) & (!g1726) & (g3190) & (g3191)) + ((!g827) & (g1726) & (g3190) & (!g3191)) + ((!g827) & (g1726) & (g3190) & (g3191)) + ((g827) & (!g1726) & (!g3190) & (g3191)) + ((g827) & (!g1726) & (g3190) & (!g3191)) + ((g827) & (g1726) & (!g3190) & (!g3191)) + ((g827) & (g1726) & (g3190) & (g3191)));
	assign g8225 = (((!g3464) & (g5398) & (!g3193)) + ((!g3464) & (g5398) & (g3193)) + ((g3464) & (!g5398) & (g3193)) + ((g3464) & (g5398) & (g3193)));
	assign g3194 = (((!g1661) & (!g1683) & (g3122) & (g3149) & (g3123)) + ((!g1661) & (g1683) & (!g3122) & (g3149) & (!g3123)) + ((!g1661) & (g1683) & (!g3122) & (g3149) & (g3123)) + ((!g1661) & (g1683) & (g3122) & (!g3149) & (g3123)) + ((!g1661) & (g1683) & (g3122) & (g3149) & (!g3123)) + ((!g1661) & (g1683) & (g3122) & (g3149) & (g3123)) + ((g1661) & (!g1683) & (!g3122) & (g3149) & (g3123)) + ((g1661) & (!g1683) & (g3122) & (g3149) & (!g3123)) + ((g1661) & (!g1683) & (g3122) & (g3149) & (g3123)) + ((g1661) & (g1683) & (!g3122) & (!g3149) & (g3123)) + ((g1661) & (g1683) & (!g3122) & (g3149) & (!g3123)) + ((g1661) & (g1683) & (!g3122) & (g3149) & (g3123)) + ((g1661) & (g1683) & (g3122) & (!g3149) & (!g3123)) + ((g1661) & (g1683) & (g3122) & (!g3149) & (g3123)) + ((g1661) & (g1683) & (g3122) & (g3149) & (!g3123)) + ((g1661) & (g1683) & (g3122) & (g3149) & (g3123)));
	assign g3195 = (((!g827) & (!g1728) & (g3193) & (!g3194)) + ((!g827) & (!g1728) & (g3193) & (g3194)) + ((!g827) & (g1728) & (g3193) & (!g3194)) + ((!g827) & (g1728) & (g3193) & (g3194)) + ((g827) & (!g1728) & (!g3193) & (g3194)) + ((g827) & (!g1728) & (g3193) & (!g3194)) + ((g827) & (g1728) & (!g3193) & (!g3194)) + ((g827) & (g1728) & (g3193) & (g3194)));
	assign g8226 = (((!g3499) & (g5400) & (!g3196)) + ((!g3499) & (g5400) & (g3196)) + ((g3499) & (!g5400) & (g3196)) + ((g3499) & (g5400) & (g3196)));
	assign g3197 = (((!g1663) & (!g1691) & (g3125) & (g3155) & (g3126)) + ((!g1663) & (g1691) & (!g3125) & (g3155) & (!g3126)) + ((!g1663) & (g1691) & (!g3125) & (g3155) & (g3126)) + ((!g1663) & (g1691) & (g3125) & (!g3155) & (g3126)) + ((!g1663) & (g1691) & (g3125) & (g3155) & (!g3126)) + ((!g1663) & (g1691) & (g3125) & (g3155) & (g3126)) + ((g1663) & (!g1691) & (!g3125) & (g3155) & (g3126)) + ((g1663) & (!g1691) & (g3125) & (g3155) & (!g3126)) + ((g1663) & (!g1691) & (g3125) & (g3155) & (g3126)) + ((g1663) & (g1691) & (!g3125) & (!g3155) & (g3126)) + ((g1663) & (g1691) & (!g3125) & (g3155) & (!g3126)) + ((g1663) & (g1691) & (!g3125) & (g3155) & (g3126)) + ((g1663) & (g1691) & (g3125) & (!g3155) & (!g3126)) + ((g1663) & (g1691) & (g3125) & (!g3155) & (g3126)) + ((g1663) & (g1691) & (g3125) & (g3155) & (!g3126)) + ((g1663) & (g1691) & (g3125) & (g3155) & (g3126)));
	assign g3198 = (((!g827) & (!g1730) & (g3196) & (!g3197)) + ((!g827) & (!g1730) & (g3196) & (g3197)) + ((!g827) & (g1730) & (g3196) & (!g3197)) + ((!g827) & (g1730) & (g3196) & (g3197)) + ((g827) & (!g1730) & (!g3196) & (g3197)) + ((g827) & (!g1730) & (g3196) & (!g3197)) + ((g827) & (g1730) & (!g3196) & (!g3197)) + ((g827) & (g1730) & (g3196) & (g3197)));
	assign g8227 = (((!g2017) & (g5953) & (!g3199)) + ((!g2017) & (g5953) & (g3199)) + ((g2017) & (!g5953) & (g3199)) + ((g2017) & (g5953) & (g3199)));
	assign g3200 = (((!g1665) & (!g1699) & (g3128) & (g3163) & (g3129)) + ((!g1665) & (g1699) & (!g3128) & (g3163) & (!g3129)) + ((!g1665) & (g1699) & (!g3128) & (g3163) & (g3129)) + ((!g1665) & (g1699) & (g3128) & (!g3163) & (g3129)) + ((!g1665) & (g1699) & (g3128) & (g3163) & (!g3129)) + ((!g1665) & (g1699) & (g3128) & (g3163) & (g3129)) + ((g1665) & (!g1699) & (!g3128) & (g3163) & (g3129)) + ((g1665) & (!g1699) & (g3128) & (g3163) & (!g3129)) + ((g1665) & (!g1699) & (g3128) & (g3163) & (g3129)) + ((g1665) & (g1699) & (!g3128) & (!g3163) & (g3129)) + ((g1665) & (g1699) & (!g3128) & (g3163) & (!g3129)) + ((g1665) & (g1699) & (!g3128) & (g3163) & (g3129)) + ((g1665) & (g1699) & (g3128) & (!g3163) & (!g3129)) + ((g1665) & (g1699) & (g3128) & (!g3163) & (g3129)) + ((g1665) & (g1699) & (g3128) & (g3163) & (!g3129)) + ((g1665) & (g1699) & (g3128) & (g3163) & (g3129)));
	assign g3201 = (((!g827) & (!g1732) & (g3199) & (!g3200)) + ((!g827) & (!g1732) & (g3199) & (g3200)) + ((!g827) & (g1732) & (g3199) & (!g3200)) + ((!g827) & (g1732) & (g3199) & (g3200)) + ((g827) & (!g1732) & (!g3199) & (g3200)) + ((g827) & (!g1732) & (g3199) & (!g3200)) + ((g827) & (g1732) & (!g3199) & (!g3200)) + ((g827) & (g1732) & (g3199) & (g3200)));
	assign g8228 = (((!g3429) & (g5405) & (!g3202)) + ((!g3429) & (g5405) & (g3202)) + ((g3429) & (!g5405) & (g3202)) + ((g3429) & (g5405) & (g3202)));
	assign g3203 = (((!g1667) & (!g1707) & (g3131) & (g3170) & (g3132)) + ((!g1667) & (g1707) & (!g3131) & (g3170) & (!g3132)) + ((!g1667) & (g1707) & (!g3131) & (g3170) & (g3132)) + ((!g1667) & (g1707) & (g3131) & (!g3170) & (g3132)) + ((!g1667) & (g1707) & (g3131) & (g3170) & (!g3132)) + ((!g1667) & (g1707) & (g3131) & (g3170) & (g3132)) + ((g1667) & (!g1707) & (!g3131) & (g3170) & (g3132)) + ((g1667) & (!g1707) & (g3131) & (g3170) & (!g3132)) + ((g1667) & (!g1707) & (g3131) & (g3170) & (g3132)) + ((g1667) & (g1707) & (!g3131) & (!g3170) & (g3132)) + ((g1667) & (g1707) & (!g3131) & (g3170) & (!g3132)) + ((g1667) & (g1707) & (!g3131) & (g3170) & (g3132)) + ((g1667) & (g1707) & (g3131) & (!g3170) & (!g3132)) + ((g1667) & (g1707) & (g3131) & (!g3170) & (g3132)) + ((g1667) & (g1707) & (g3131) & (g3170) & (!g3132)) + ((g1667) & (g1707) & (g3131) & (g3170) & (g3132)));
	assign g3204 = (((!g827) & (!g1734) & (g3202) & (!g3203)) + ((!g827) & (!g1734) & (g3202) & (g3203)) + ((!g827) & (g1734) & (g3202) & (!g3203)) + ((!g827) & (g1734) & (g3202) & (g3203)) + ((g827) & (!g1734) & (!g3202) & (g3203)) + ((g827) & (!g1734) & (g3202) & (!g3203)) + ((g827) & (g1734) & (!g3202) & (!g3203)) + ((g827) & (g1734) & (g3202) & (g3203)));
	assign g3205 = (((!g1669) & (!g1685) & (g2519) & (g2556) & (g3134)) + ((!g1669) & (g1685) & (!g2519) & (g2556) & (!g3134)) + ((!g1669) & (g1685) & (!g2519) & (g2556) & (g3134)) + ((!g1669) & (g1685) & (g2519) & (!g2556) & (g3134)) + ((!g1669) & (g1685) & (g2519) & (g2556) & (!g3134)) + ((!g1669) & (g1685) & (g2519) & (g2556) & (g3134)) + ((g1669) & (!g1685) & (!g2519) & (g2556) & (g3134)) + ((g1669) & (!g1685) & (g2519) & (g2556) & (!g3134)) + ((g1669) & (!g1685) & (g2519) & (g2556) & (g3134)) + ((g1669) & (g1685) & (!g2519) & (!g2556) & (g3134)) + ((g1669) & (g1685) & (!g2519) & (g2556) & (!g3134)) + ((g1669) & (g1685) & (!g2519) & (g2556) & (g3134)) + ((g1669) & (g1685) & (g2519) & (!g2556) & (!g3134)) + ((g1669) & (g1685) & (g2519) & (!g2556) & (g3134)) + ((g1669) & (g1685) & (g2519) & (g2556) & (!g3134)) + ((g1669) & (g1685) & (g2519) & (g2556) & (g3134)));
	assign g3206 = (((!g827) & (!g1736) & (g2602) & (!g3205)) + ((!g827) & (!g1736) & (g2602) & (g3205)) + ((!g827) & (g1736) & (g2602) & (!g3205)) + ((!g827) & (g1736) & (g2602) & (g3205)) + ((g827) & (!g1736) & (!g2602) & (g3205)) + ((g827) & (!g1736) & (g2602) & (!g3205)) + ((g827) & (g1736) & (!g2602) & (!g3205)) + ((g827) & (g1736) & (g2602) & (g3205)));
	assign g8229 = (((!g3464) & (g5407) & (!g3207)) + ((!g3464) & (g5407) & (g3207)) + ((g3464) & (!g5407) & (g3207)) + ((g3464) & (g5407) & (g3207)));
	assign g3208 = (((!g1671) & (!g1693) & (g3136) & (g3157) & (g3137)) + ((!g1671) & (g1693) & (!g3136) & (g3157) & (!g3137)) + ((!g1671) & (g1693) & (!g3136) & (g3157) & (g3137)) + ((!g1671) & (g1693) & (g3136) & (!g3157) & (g3137)) + ((!g1671) & (g1693) & (g3136) & (g3157) & (!g3137)) + ((!g1671) & (g1693) & (g3136) & (g3157) & (g3137)) + ((g1671) & (!g1693) & (!g3136) & (g3157) & (g3137)) + ((g1671) & (!g1693) & (g3136) & (g3157) & (!g3137)) + ((g1671) & (!g1693) & (g3136) & (g3157) & (g3137)) + ((g1671) & (g1693) & (!g3136) & (!g3157) & (g3137)) + ((g1671) & (g1693) & (!g3136) & (g3157) & (!g3137)) + ((g1671) & (g1693) & (!g3136) & (g3157) & (g3137)) + ((g1671) & (g1693) & (g3136) & (!g3157) & (!g3137)) + ((g1671) & (g1693) & (g3136) & (!g3157) & (g3137)) + ((g1671) & (g1693) & (g3136) & (g3157) & (!g3137)) + ((g1671) & (g1693) & (g3136) & (g3157) & (g3137)));
	assign g3209 = (((!g827) & (!g1738) & (g3207) & (!g3208)) + ((!g827) & (!g1738) & (g3207) & (g3208)) + ((!g827) & (g1738) & (g3207) & (!g3208)) + ((!g827) & (g1738) & (g3207) & (g3208)) + ((g827) & (!g1738) & (!g3207) & (g3208)) + ((g827) & (!g1738) & (g3207) & (!g3208)) + ((g827) & (g1738) & (!g3207) & (!g3208)) + ((g827) & (g1738) & (g3207) & (g3208)));
	assign g8230 = (((!g3429) & (g5410) & (!g3210)) + ((!g3429) & (g5410) & (g3210)) + ((g3429) & (!g5410) & (g3210)) + ((g3429) & (g5410) & (g3210)));
	assign g3211 = (((!g1673) & (!g1701) & (g3139) & (g3165) & (g3140)) + ((!g1673) & (g1701) & (!g3139) & (g3165) & (!g3140)) + ((!g1673) & (g1701) & (!g3139) & (g3165) & (g3140)) + ((!g1673) & (g1701) & (g3139) & (!g3165) & (g3140)) + ((!g1673) & (g1701) & (g3139) & (g3165) & (!g3140)) + ((!g1673) & (g1701) & (g3139) & (g3165) & (g3140)) + ((g1673) & (!g1701) & (!g3139) & (g3165) & (g3140)) + ((g1673) & (!g1701) & (g3139) & (g3165) & (!g3140)) + ((g1673) & (!g1701) & (g3139) & (g3165) & (g3140)) + ((g1673) & (g1701) & (!g3139) & (!g3165) & (g3140)) + ((g1673) & (g1701) & (!g3139) & (g3165) & (!g3140)) + ((g1673) & (g1701) & (!g3139) & (g3165) & (g3140)) + ((g1673) & (g1701) & (g3139) & (!g3165) & (!g3140)) + ((g1673) & (g1701) & (g3139) & (!g3165) & (g3140)) + ((g1673) & (g1701) & (g3139) & (g3165) & (!g3140)) + ((g1673) & (g1701) & (g3139) & (g3165) & (g3140)));
	assign g3212 = (((!g827) & (!g1740) & (g3210) & (!g3211)) + ((!g827) & (!g1740) & (g3210) & (g3211)) + ((!g827) & (g1740) & (g3210) & (!g3211)) + ((!g827) & (g1740) & (g3210) & (g3211)) + ((g827) & (!g1740) & (!g3210) & (g3211)) + ((g827) & (!g1740) & (g3210) & (!g3211)) + ((g827) & (g1740) & (!g3210) & (!g3211)) + ((g827) & (g1740) & (g3210) & (g3211)));
	assign g8231 = (((!g2017) & (g5935) & (!g3213)) + ((!g2017) & (g5935) & (g3213)) + ((g2017) & (!g5935) & (g3213)) + ((g2017) & (g5935) & (g3213)));
	assign g3214 = (((!g1675) & (!g1709) & (g3142) & (g3172) & (g3143)) + ((!g1675) & (g1709) & (!g3142) & (g3172) & (!g3143)) + ((!g1675) & (g1709) & (!g3142) & (g3172) & (g3143)) + ((!g1675) & (g1709) & (g3142) & (!g3172) & (g3143)) + ((!g1675) & (g1709) & (g3142) & (g3172) & (!g3143)) + ((!g1675) & (g1709) & (g3142) & (g3172) & (g3143)) + ((g1675) & (!g1709) & (!g3142) & (g3172) & (g3143)) + ((g1675) & (!g1709) & (g3142) & (g3172) & (!g3143)) + ((g1675) & (!g1709) & (g3142) & (g3172) & (g3143)) + ((g1675) & (g1709) & (!g3142) & (!g3172) & (g3143)) + ((g1675) & (g1709) & (!g3142) & (g3172) & (!g3143)) + ((g1675) & (g1709) & (!g3142) & (g3172) & (g3143)) + ((g1675) & (g1709) & (g3142) & (!g3172) & (!g3143)) + ((g1675) & (g1709) & (g3142) & (!g3172) & (g3143)) + ((g1675) & (g1709) & (g3142) & (g3172) & (!g3143)) + ((g1675) & (g1709) & (g3142) & (g3172) & (g3143)));
	assign g3215 = (((!g827) & (!g1742) & (g3213) & (!g3214)) + ((!g827) & (!g1742) & (g3213) & (g3214)) + ((!g827) & (g1742) & (g3213) & (!g3214)) + ((!g827) & (g1742) & (g3213) & (g3214)) + ((g827) & (!g1742) & (!g3213) & (g3214)) + ((g827) & (!g1742) & (g3213) & (!g3214)) + ((g827) & (g1742) & (!g3213) & (!g3214)) + ((g827) & (g1742) & (g3213) & (g3214)));
	assign g3216 = (((!g1957) & (g1958) & (g1959)) + ((g1957) & (!g1958) & (g1959)) + ((g1957) & (g1958) & (!g1959)) + ((g1957) & (g1958) & (g1959)));
	assign g3217 = (((!g1995) & (!g1996) & (!g1997) & (!g1998) & (g1999)) + ((!g1995) & (!g1996) & (!g1997) & (g1998) & (!g1999)) + ((!g1995) & (!g1996) & (g1997) & (!g1998) & (!g1999)) + ((!g1995) & (!g1996) & (g1997) & (g1998) & (g1999)) + ((!g1995) & (g1996) & (!g1997) & (!g1998) & (!g1999)) + ((!g1995) & (g1996) & (!g1997) & (g1998) & (g1999)) + ((!g1995) & (g1996) & (g1997) & (!g1998) & (!g1999)) + ((!g1995) & (g1996) & (g1997) & (g1998) & (g1999)) + ((g1995) & (!g1996) & (!g1997) & (!g1998) & (g1999)) + ((g1995) & (!g1996) & (!g1997) & (g1998) & (!g1999)) + ((g1995) & (!g1996) & (g1997) & (!g1998) & (g1999)) + ((g1995) & (!g1996) & (g1997) & (g1998) & (!g1999)) + ((g1995) & (g1996) & (!g1997) & (!g1998) & (g1999)) + ((g1995) & (g1996) & (!g1997) & (g1998) & (!g1999)) + ((g1995) & (g1996) & (g1997) & (!g1998) & (!g1999)) + ((g1995) & (g1996) & (g1997) & (g1998) & (g1999)));
	assign g3218 = (((!g1720) & (g2601)) + ((g1720) & (!g2601)));
	assign g3219 = (((!g1653) & (!g1681) & (g2518) & (g2555) & (g3111) & (g3218)) + ((!g1653) & (g1681) & (!g2518) & (g2555) & (!g3111) & (g3218)) + ((!g1653) & (g1681) & (!g2518) & (g2555) & (g3111) & (g3218)) + ((!g1653) & (g1681) & (g2518) & (!g2555) & (g3111) & (g3218)) + ((!g1653) & (g1681) & (g2518) & (g2555) & (!g3111) & (g3218)) + ((!g1653) & (g1681) & (g2518) & (g2555) & (g3111) & (g3218)) + ((g1653) & (!g1681) & (!g2518) & (g2555) & (g3111) & (g3218)) + ((g1653) & (!g1681) & (g2518) & (g2555) & (!g3111) & (g3218)) + ((g1653) & (!g1681) & (g2518) & (g2555) & (g3111) & (g3218)) + ((g1653) & (g1681) & (!g2518) & (!g2555) & (g3111) & (g3218)) + ((g1653) & (g1681) & (!g2518) & (g2555) & (!g3111) & (g3218)) + ((g1653) & (g1681) & (!g2518) & (g2555) & (g3111) & (g3218)) + ((g1653) & (g1681) & (g2518) & (!g2555) & (!g3111) & (g3218)) + ((g1653) & (g1681) & (g2518) & (!g2555) & (g3111) & (g3218)) + ((g1653) & (g1681) & (g2518) & (g2555) & (!g3111) & (g3218)) + ((g1653) & (g1681) & (g2518) & (g2555) & (g3111) & (g3218)));
	assign g3220 = (((g1720) & (g2601)));
	assign g3221 = (((!g827) & (!g1748) & (g2649) & (!g3219) & (!g3220)) + ((!g827) & (!g1748) & (g2649) & (!g3219) & (g3220)) + ((!g827) & (!g1748) & (g2649) & (g3219) & (!g3220)) + ((!g827) & (!g1748) & (g2649) & (g3219) & (g3220)) + ((!g827) & (g1748) & (g2649) & (!g3219) & (!g3220)) + ((!g827) & (g1748) & (g2649) & (!g3219) & (g3220)) + ((!g827) & (g1748) & (g2649) & (g3219) & (!g3220)) + ((!g827) & (g1748) & (g2649) & (g3219) & (g3220)) + ((g827) & (!g1748) & (!g2649) & (!g3219) & (g3220)) + ((g827) & (!g1748) & (!g2649) & (g3219) & (!g3220)) + ((g827) & (!g1748) & (!g2649) & (g3219) & (g3220)) + ((g827) & (!g1748) & (g2649) & (!g3219) & (!g3220)) + ((g827) & (g1748) & (!g2649) & (!g3219) & (!g3220)) + ((g827) & (g1748) & (g2649) & (!g3219) & (g3220)) + ((g827) & (g1748) & (g2649) & (g3219) & (!g3220)) + ((g827) & (g1748) & (g2649) & (g3219) & (g3220)));
	assign g8232 = (((!g3464) & (g5416) & (!g3222)) + ((!g3464) & (g5416) & (g3222)) + ((g3464) & (!g5416) & (g3222)) + ((g3464) & (g5416) & (g3222)));
	assign g3223 = (((!g1728) & (g3193)) + ((g1728) & (!g3193)));
	assign g3224 = (((!g1661) & (!g1683) & (g3122) & (g3149) & (g3123) & (g3223)) + ((!g1661) & (g1683) & (!g3122) & (g3149) & (!g3123) & (g3223)) + ((!g1661) & (g1683) & (!g3122) & (g3149) & (g3123) & (g3223)) + ((!g1661) & (g1683) & (g3122) & (!g3149) & (g3123) & (g3223)) + ((!g1661) & (g1683) & (g3122) & (g3149) & (!g3123) & (g3223)) + ((!g1661) & (g1683) & (g3122) & (g3149) & (g3123) & (g3223)) + ((g1661) & (!g1683) & (!g3122) & (g3149) & (g3123) & (g3223)) + ((g1661) & (!g1683) & (g3122) & (g3149) & (!g3123) & (g3223)) + ((g1661) & (!g1683) & (g3122) & (g3149) & (g3123) & (g3223)) + ((g1661) & (g1683) & (!g3122) & (!g3149) & (g3123) & (g3223)) + ((g1661) & (g1683) & (!g3122) & (g3149) & (!g3123) & (g3223)) + ((g1661) & (g1683) & (!g3122) & (g3149) & (g3123) & (g3223)) + ((g1661) & (g1683) & (g3122) & (!g3149) & (!g3123) & (g3223)) + ((g1661) & (g1683) & (g3122) & (!g3149) & (g3123) & (g3223)) + ((g1661) & (g1683) & (g3122) & (g3149) & (!g3123) & (g3223)) + ((g1661) & (g1683) & (g3122) & (g3149) & (g3123) & (g3223)));
	assign g3225 = (((g1728) & (g3193)));
	assign g3226 = (((!g827) & (!g1750) & (g3222) & (!g3224) & (!g3225)) + ((!g827) & (!g1750) & (g3222) & (!g3224) & (g3225)) + ((!g827) & (!g1750) & (g3222) & (g3224) & (!g3225)) + ((!g827) & (!g1750) & (g3222) & (g3224) & (g3225)) + ((!g827) & (g1750) & (g3222) & (!g3224) & (!g3225)) + ((!g827) & (g1750) & (g3222) & (!g3224) & (g3225)) + ((!g827) & (g1750) & (g3222) & (g3224) & (!g3225)) + ((!g827) & (g1750) & (g3222) & (g3224) & (g3225)) + ((g827) & (!g1750) & (!g3222) & (!g3224) & (g3225)) + ((g827) & (!g1750) & (!g3222) & (g3224) & (!g3225)) + ((g827) & (!g1750) & (!g3222) & (g3224) & (g3225)) + ((g827) & (!g1750) & (g3222) & (!g3224) & (!g3225)) + ((g827) & (g1750) & (!g3222) & (!g3224) & (!g3225)) + ((g827) & (g1750) & (g3222) & (!g3224) & (g3225)) + ((g827) & (g1750) & (g3222) & (g3224) & (!g3225)) + ((g827) & (g1750) & (g3222) & (g3224) & (g3225)));
	assign g3227 = (((!g1736) & (g2602)) + ((g1736) & (!g2602)));
	assign g3228 = (((!g1669) & (!g1685) & (g2519) & (g2556) & (g3134) & (g3227)) + ((!g1669) & (g1685) & (!g2519) & (g2556) & (!g3134) & (g3227)) + ((!g1669) & (g1685) & (!g2519) & (g2556) & (g3134) & (g3227)) + ((!g1669) & (g1685) & (g2519) & (!g2556) & (g3134) & (g3227)) + ((!g1669) & (g1685) & (g2519) & (g2556) & (!g3134) & (g3227)) + ((!g1669) & (g1685) & (g2519) & (g2556) & (g3134) & (g3227)) + ((g1669) & (!g1685) & (!g2519) & (g2556) & (g3134) & (g3227)) + ((g1669) & (!g1685) & (g2519) & (g2556) & (!g3134) & (g3227)) + ((g1669) & (!g1685) & (g2519) & (g2556) & (g3134) & (g3227)) + ((g1669) & (g1685) & (!g2519) & (!g2556) & (g3134) & (g3227)) + ((g1669) & (g1685) & (!g2519) & (g2556) & (!g3134) & (g3227)) + ((g1669) & (g1685) & (!g2519) & (g2556) & (g3134) & (g3227)) + ((g1669) & (g1685) & (g2519) & (!g2556) & (!g3134) & (g3227)) + ((g1669) & (g1685) & (g2519) & (!g2556) & (g3134) & (g3227)) + ((g1669) & (g1685) & (g2519) & (g2556) & (!g3134) & (g3227)) + ((g1669) & (g1685) & (g2519) & (g2556) & (g3134) & (g3227)));
	assign g3229 = (((g1736) & (g2602)));
	assign g3230 = (((!g827) & (!g1752) & (g2650) & (!g3228) & (!g3229)) + ((!g827) & (!g1752) & (g2650) & (!g3228) & (g3229)) + ((!g827) & (!g1752) & (g2650) & (g3228) & (!g3229)) + ((!g827) & (!g1752) & (g2650) & (g3228) & (g3229)) + ((!g827) & (g1752) & (g2650) & (!g3228) & (!g3229)) + ((!g827) & (g1752) & (g2650) & (!g3228) & (g3229)) + ((!g827) & (g1752) & (g2650) & (g3228) & (!g3229)) + ((!g827) & (g1752) & (g2650) & (g3228) & (g3229)) + ((g827) & (!g1752) & (!g2650) & (!g3228) & (g3229)) + ((g827) & (!g1752) & (!g2650) & (g3228) & (!g3229)) + ((g827) & (!g1752) & (!g2650) & (g3228) & (g3229)) + ((g827) & (!g1752) & (g2650) & (!g3228) & (!g3229)) + ((g827) & (g1752) & (!g2650) & (!g3228) & (!g3229)) + ((g827) & (g1752) & (g2650) & (!g3228) & (g3229)) + ((g827) & (g1752) & (g2650) & (g3228) & (!g3229)) + ((g827) & (g1752) & (g2650) & (g3228) & (g3229)));
	assign g3231 = (((!g1714) & (g2598)) + ((g1714) & (!g2598)));
	assign g3232 = (((!g1647) & (!g1687) & (g2515) & (g2551) & (g3104) & (g3231)) + ((!g1647) & (g1687) & (!g2515) & (g2551) & (!g3104) & (g3231)) + ((!g1647) & (g1687) & (!g2515) & (g2551) & (g3104) & (g3231)) + ((!g1647) & (g1687) & (g2515) & (!g2551) & (g3104) & (g3231)) + ((!g1647) & (g1687) & (g2515) & (g2551) & (!g3104) & (g3231)) + ((!g1647) & (g1687) & (g2515) & (g2551) & (g3104) & (g3231)) + ((g1647) & (!g1687) & (!g2515) & (g2551) & (g3104) & (g3231)) + ((g1647) & (!g1687) & (g2515) & (g2551) & (!g3104) & (g3231)) + ((g1647) & (!g1687) & (g2515) & (g2551) & (g3104) & (g3231)) + ((g1647) & (g1687) & (!g2515) & (!g2551) & (g3104) & (g3231)) + ((g1647) & (g1687) & (!g2515) & (g2551) & (!g3104) & (g3231)) + ((g1647) & (g1687) & (!g2515) & (g2551) & (g3104) & (g3231)) + ((g1647) & (g1687) & (g2515) & (!g2551) & (!g3104) & (g3231)) + ((g1647) & (g1687) & (g2515) & (!g2551) & (g3104) & (g3231)) + ((g1647) & (g1687) & (g2515) & (g2551) & (!g3104) & (g3231)) + ((g1647) & (g1687) & (g2515) & (g2551) & (g3104) & (g3231)));
	assign g3233 = (((g1714) & (g2598)));
	assign g3234 = (((!g827) & (!g1754) & (g2647) & (!g3232) & (!g3233)) + ((!g827) & (!g1754) & (g2647) & (!g3232) & (g3233)) + ((!g827) & (!g1754) & (g2647) & (g3232) & (!g3233)) + ((!g827) & (!g1754) & (g2647) & (g3232) & (g3233)) + ((!g827) & (g1754) & (g2647) & (!g3232) & (!g3233)) + ((!g827) & (g1754) & (g2647) & (!g3232) & (g3233)) + ((!g827) & (g1754) & (g2647) & (g3232) & (!g3233)) + ((!g827) & (g1754) & (g2647) & (g3232) & (g3233)) + ((g827) & (!g1754) & (!g2647) & (!g3232) & (g3233)) + ((g827) & (!g1754) & (!g2647) & (g3232) & (!g3233)) + ((g827) & (!g1754) & (!g2647) & (g3232) & (g3233)) + ((g827) & (!g1754) & (g2647) & (!g3232) & (!g3233)) + ((g827) & (g1754) & (!g2647) & (!g3232) & (!g3233)) + ((g827) & (g1754) & (g2647) & (!g3232) & (g3233)) + ((g827) & (g1754) & (g2647) & (g3232) & (!g3233)) + ((g827) & (g1754) & (g2647) & (g3232) & (g3233)));
	assign g8233 = (((!g2017) & (g5928) & (!g3235)) + ((!g2017) & (g5928) & (g3235)) + ((g2017) & (!g5928) & (g3235)) + ((g2017) & (g5928) & (g3235)));
	assign g3236 = (((!g1722) & (g3184)) + ((g1722) & (!g3184)));
	assign g3237 = (((!g1655) & (!g1689) & (g3113) & (g3153) & (g3114) & (g3236)) + ((!g1655) & (g1689) & (!g3113) & (g3153) & (!g3114) & (g3236)) + ((!g1655) & (g1689) & (!g3113) & (g3153) & (g3114) & (g3236)) + ((!g1655) & (g1689) & (g3113) & (!g3153) & (g3114) & (g3236)) + ((!g1655) & (g1689) & (g3113) & (g3153) & (!g3114) & (g3236)) + ((!g1655) & (g1689) & (g3113) & (g3153) & (g3114) & (g3236)) + ((g1655) & (!g1689) & (!g3113) & (g3153) & (g3114) & (g3236)) + ((g1655) & (!g1689) & (g3113) & (g3153) & (!g3114) & (g3236)) + ((g1655) & (!g1689) & (g3113) & (g3153) & (g3114) & (g3236)) + ((g1655) & (g1689) & (!g3113) & (!g3153) & (g3114) & (g3236)) + ((g1655) & (g1689) & (!g3113) & (g3153) & (!g3114) & (g3236)) + ((g1655) & (g1689) & (!g3113) & (g3153) & (g3114) & (g3236)) + ((g1655) & (g1689) & (g3113) & (!g3153) & (!g3114) & (g3236)) + ((g1655) & (g1689) & (g3113) & (!g3153) & (g3114) & (g3236)) + ((g1655) & (g1689) & (g3113) & (g3153) & (!g3114) & (g3236)) + ((g1655) & (g1689) & (g3113) & (g3153) & (g3114) & (g3236)));
	assign g3238 = (((g1722) & (g3184)));
	assign g3239 = (((!g827) & (!g1756) & (g3235) & (!g3237) & (!g3238)) + ((!g827) & (!g1756) & (g3235) & (!g3237) & (g3238)) + ((!g827) & (!g1756) & (g3235) & (g3237) & (!g3238)) + ((!g827) & (!g1756) & (g3235) & (g3237) & (g3238)) + ((!g827) & (g1756) & (g3235) & (!g3237) & (!g3238)) + ((!g827) & (g1756) & (g3235) & (!g3237) & (g3238)) + ((!g827) & (g1756) & (g3235) & (g3237) & (!g3238)) + ((!g827) & (g1756) & (g3235) & (g3237) & (g3238)) + ((g827) & (!g1756) & (!g3235) & (!g3237) & (g3238)) + ((g827) & (!g1756) & (!g3235) & (g3237) & (!g3238)) + ((g827) & (!g1756) & (!g3235) & (g3237) & (g3238)) + ((g827) & (!g1756) & (g3235) & (!g3237) & (!g3238)) + ((g827) & (g1756) & (!g3235) & (!g3237) & (!g3238)) + ((g827) & (g1756) & (g3235) & (!g3237) & (g3238)) + ((g827) & (g1756) & (g3235) & (g3237) & (!g3238)) + ((g827) & (g1756) & (g3235) & (g3237) & (g3238)));
	assign g8234 = (((!g3499) & (g5421) & (!g3240)) + ((!g3499) & (g5421) & (g3240)) + ((g3499) & (!g5421) & (g3240)) + ((g3499) & (g5421) & (g3240)));
	assign g3241 = (((!g1730) & (g3196)) + ((g1730) & (!g3196)));
	assign g3242 = (((!g1663) & (!g1691) & (g3125) & (g3155) & (g3126) & (g3241)) + ((!g1663) & (g1691) & (!g3125) & (g3155) & (!g3126) & (g3241)) + ((!g1663) & (g1691) & (!g3125) & (g3155) & (g3126) & (g3241)) + ((!g1663) & (g1691) & (g3125) & (!g3155) & (g3126) & (g3241)) + ((!g1663) & (g1691) & (g3125) & (g3155) & (!g3126) & (g3241)) + ((!g1663) & (g1691) & (g3125) & (g3155) & (g3126) & (g3241)) + ((g1663) & (!g1691) & (!g3125) & (g3155) & (g3126) & (g3241)) + ((g1663) & (!g1691) & (g3125) & (g3155) & (!g3126) & (g3241)) + ((g1663) & (!g1691) & (g3125) & (g3155) & (g3126) & (g3241)) + ((g1663) & (g1691) & (!g3125) & (!g3155) & (g3126) & (g3241)) + ((g1663) & (g1691) & (!g3125) & (g3155) & (!g3126) & (g3241)) + ((g1663) & (g1691) & (!g3125) & (g3155) & (g3126) & (g3241)) + ((g1663) & (g1691) & (g3125) & (!g3155) & (!g3126) & (g3241)) + ((g1663) & (g1691) & (g3125) & (!g3155) & (g3126) & (g3241)) + ((g1663) & (g1691) & (g3125) & (g3155) & (!g3126) & (g3241)) + ((g1663) & (g1691) & (g3125) & (g3155) & (g3126) & (g3241)));
	assign g3243 = (((g1730) & (g3196)));
	assign g3244 = (((!g827) & (!g1758) & (g3240) & (!g3242) & (!g3243)) + ((!g827) & (!g1758) & (g3240) & (!g3242) & (g3243)) + ((!g827) & (!g1758) & (g3240) & (g3242) & (!g3243)) + ((!g827) & (!g1758) & (g3240) & (g3242) & (g3243)) + ((!g827) & (g1758) & (g3240) & (!g3242) & (!g3243)) + ((!g827) & (g1758) & (g3240) & (!g3242) & (g3243)) + ((!g827) & (g1758) & (g3240) & (g3242) & (!g3243)) + ((!g827) & (g1758) & (g3240) & (g3242) & (g3243)) + ((g827) & (!g1758) & (!g3240) & (!g3242) & (g3243)) + ((g827) & (!g1758) & (!g3240) & (g3242) & (!g3243)) + ((g827) & (!g1758) & (!g3240) & (g3242) & (g3243)) + ((g827) & (!g1758) & (g3240) & (!g3242) & (!g3243)) + ((g827) & (g1758) & (!g3240) & (!g3242) & (!g3243)) + ((g827) & (g1758) & (g3240) & (!g3242) & (g3243)) + ((g827) & (g1758) & (g3240) & (g3242) & (!g3243)) + ((g827) & (g1758) & (g3240) & (g3242) & (g3243)));
	assign g8235 = (((!g3464) & (g5425) & (!g3245)) + ((!g3464) & (g5425) & (g3245)) + ((g3464) & (!g5425) & (g3245)) + ((g3464) & (g5425) & (g3245)));
	assign g3246 = (((!g1738) & (g3207)) + ((g1738) & (!g3207)));
	assign g3247 = (((!g1671) & (!g1693) & (g3136) & (g3157) & (g3137) & (g3246)) + ((!g1671) & (g1693) & (!g3136) & (g3157) & (!g3137) & (g3246)) + ((!g1671) & (g1693) & (!g3136) & (g3157) & (g3137) & (g3246)) + ((!g1671) & (g1693) & (g3136) & (!g3157) & (g3137) & (g3246)) + ((!g1671) & (g1693) & (g3136) & (g3157) & (!g3137) & (g3246)) + ((!g1671) & (g1693) & (g3136) & (g3157) & (g3137) & (g3246)) + ((g1671) & (!g1693) & (!g3136) & (g3157) & (g3137) & (g3246)) + ((g1671) & (!g1693) & (g3136) & (g3157) & (!g3137) & (g3246)) + ((g1671) & (!g1693) & (g3136) & (g3157) & (g3137) & (g3246)) + ((g1671) & (g1693) & (!g3136) & (!g3157) & (g3137) & (g3246)) + ((g1671) & (g1693) & (!g3136) & (g3157) & (!g3137) & (g3246)) + ((g1671) & (g1693) & (!g3136) & (g3157) & (g3137) & (g3246)) + ((g1671) & (g1693) & (g3136) & (!g3157) & (!g3137) & (g3246)) + ((g1671) & (g1693) & (g3136) & (!g3157) & (g3137) & (g3246)) + ((g1671) & (g1693) & (g3136) & (g3157) & (!g3137) & (g3246)) + ((g1671) & (g1693) & (g3136) & (g3157) & (g3137) & (g3246)));
	assign g3248 = (((g1738) & (g3207)));
	assign g3249 = (((!g827) & (!g1760) & (g3245) & (!g3247) & (!g3248)) + ((!g827) & (!g1760) & (g3245) & (!g3247) & (g3248)) + ((!g827) & (!g1760) & (g3245) & (g3247) & (!g3248)) + ((!g827) & (!g1760) & (g3245) & (g3247) & (g3248)) + ((!g827) & (g1760) & (g3245) & (!g3247) & (!g3248)) + ((!g827) & (g1760) & (g3245) & (!g3247) & (g3248)) + ((!g827) & (g1760) & (g3245) & (g3247) & (!g3248)) + ((!g827) & (g1760) & (g3245) & (g3247) & (g3248)) + ((g827) & (!g1760) & (!g3245) & (!g3247) & (g3248)) + ((g827) & (!g1760) & (!g3245) & (g3247) & (!g3248)) + ((g827) & (!g1760) & (!g3245) & (g3247) & (g3248)) + ((g827) & (!g1760) & (g3245) & (!g3247) & (!g3248)) + ((g827) & (g1760) & (!g3245) & (!g3247) & (!g3248)) + ((g827) & (g1760) & (g3245) & (!g3247) & (g3248)) + ((g827) & (g1760) & (g3245) & (g3247) & (!g3248)) + ((g827) & (g1760) & (g3245) & (g3247) & (g3248)));
	assign g8236 = (((!g3499) & (g5429) & (!g3250)) + ((!g3499) & (g5429) & (g3250)) + ((g3499) & (!g5429) & (g3250)) + ((g3499) & (g5429) & (g3250)));
	assign g3251 = (((!g1716) & (g3177)) + ((g1716) & (!g3177)));
	assign g3252 = (((!g1649) & (!g1695) & (g3106) & (g3159) & (g3107) & (g3251)) + ((!g1649) & (g1695) & (!g3106) & (g3159) & (!g3107) & (g3251)) + ((!g1649) & (g1695) & (!g3106) & (g3159) & (g3107) & (g3251)) + ((!g1649) & (g1695) & (g3106) & (!g3159) & (g3107) & (g3251)) + ((!g1649) & (g1695) & (g3106) & (g3159) & (!g3107) & (g3251)) + ((!g1649) & (g1695) & (g3106) & (g3159) & (g3107) & (g3251)) + ((g1649) & (!g1695) & (!g3106) & (g3159) & (g3107) & (g3251)) + ((g1649) & (!g1695) & (g3106) & (g3159) & (!g3107) & (g3251)) + ((g1649) & (!g1695) & (g3106) & (g3159) & (g3107) & (g3251)) + ((g1649) & (g1695) & (!g3106) & (!g3159) & (g3107) & (g3251)) + ((g1649) & (g1695) & (!g3106) & (g3159) & (!g3107) & (g3251)) + ((g1649) & (g1695) & (!g3106) & (g3159) & (g3107) & (g3251)) + ((g1649) & (g1695) & (g3106) & (!g3159) & (!g3107) & (g3251)) + ((g1649) & (g1695) & (g3106) & (!g3159) & (g3107) & (g3251)) + ((g1649) & (g1695) & (g3106) & (g3159) & (!g3107) & (g3251)) + ((g1649) & (g1695) & (g3106) & (g3159) & (g3107) & (g3251)));
	assign g3253 = (((g1716) & (g3177)));
	assign g3254 = (((!g827) & (!g1762) & (g3250) & (!g3252) & (!g3253)) + ((!g827) & (!g1762) & (g3250) & (!g3252) & (g3253)) + ((!g827) & (!g1762) & (g3250) & (g3252) & (!g3253)) + ((!g827) & (!g1762) & (g3250) & (g3252) & (g3253)) + ((!g827) & (g1762) & (g3250) & (!g3252) & (!g3253)) + ((!g827) & (g1762) & (g3250) & (!g3252) & (g3253)) + ((!g827) & (g1762) & (g3250) & (g3252) & (!g3253)) + ((!g827) & (g1762) & (g3250) & (g3252) & (g3253)) + ((g827) & (!g1762) & (!g3250) & (!g3252) & (g3253)) + ((g827) & (!g1762) & (!g3250) & (g3252) & (!g3253)) + ((g827) & (!g1762) & (!g3250) & (g3252) & (g3253)) + ((g827) & (!g1762) & (g3250) & (!g3252) & (!g3253)) + ((g827) & (g1762) & (!g3250) & (!g3252) & (!g3253)) + ((g827) & (g1762) & (g3250) & (!g3252) & (g3253)) + ((g827) & (g1762) & (g3250) & (g3252) & (!g3253)) + ((g827) & (g1762) & (g3250) & (g3252) & (g3253)));
	assign g8237 = (((!g3464) & (g5435) & (!g3255)) + ((!g3464) & (g5435) & (g3255)) + ((g3464) & (!g5435) & (g3255)) + ((g3464) & (g5435) & (g3255)));
	assign g3256 = (((!g1724) & (g3187)) + ((g1724) & (!g3187)));
	assign g3257 = (((!g1657) & (!g1697) & (g3116) & (g3161) & (g3117) & (g3256)) + ((!g1657) & (g1697) & (!g3116) & (g3161) & (!g3117) & (g3256)) + ((!g1657) & (g1697) & (!g3116) & (g3161) & (g3117) & (g3256)) + ((!g1657) & (g1697) & (g3116) & (!g3161) & (g3117) & (g3256)) + ((!g1657) & (g1697) & (g3116) & (g3161) & (!g3117) & (g3256)) + ((!g1657) & (g1697) & (g3116) & (g3161) & (g3117) & (g3256)) + ((g1657) & (!g1697) & (!g3116) & (g3161) & (g3117) & (g3256)) + ((g1657) & (!g1697) & (g3116) & (g3161) & (!g3117) & (g3256)) + ((g1657) & (!g1697) & (g3116) & (g3161) & (g3117) & (g3256)) + ((g1657) & (g1697) & (!g3116) & (!g3161) & (g3117) & (g3256)) + ((g1657) & (g1697) & (!g3116) & (g3161) & (!g3117) & (g3256)) + ((g1657) & (g1697) & (!g3116) & (g3161) & (g3117) & (g3256)) + ((g1657) & (g1697) & (g3116) & (!g3161) & (!g3117) & (g3256)) + ((g1657) & (g1697) & (g3116) & (!g3161) & (g3117) & (g3256)) + ((g1657) & (g1697) & (g3116) & (g3161) & (!g3117) & (g3256)) + ((g1657) & (g1697) & (g3116) & (g3161) & (g3117) & (g3256)));
	assign g3258 = (((g1724) & (g3187)));
	assign g3259 = (((!g827) & (!g1764) & (g3255) & (!g3257) & (!g3258)) + ((!g827) & (!g1764) & (g3255) & (!g3257) & (g3258)) + ((!g827) & (!g1764) & (g3255) & (g3257) & (!g3258)) + ((!g827) & (!g1764) & (g3255) & (g3257) & (g3258)) + ((!g827) & (g1764) & (g3255) & (!g3257) & (!g3258)) + ((!g827) & (g1764) & (g3255) & (!g3257) & (g3258)) + ((!g827) & (g1764) & (g3255) & (g3257) & (!g3258)) + ((!g827) & (g1764) & (g3255) & (g3257) & (g3258)) + ((g827) & (!g1764) & (!g3255) & (!g3257) & (g3258)) + ((g827) & (!g1764) & (!g3255) & (g3257) & (!g3258)) + ((g827) & (!g1764) & (!g3255) & (g3257) & (g3258)) + ((g827) & (!g1764) & (g3255) & (!g3257) & (!g3258)) + ((g827) & (g1764) & (!g3255) & (!g3257) & (!g3258)) + ((g827) & (g1764) & (g3255) & (!g3257) & (g3258)) + ((g827) & (g1764) & (g3255) & (g3257) & (!g3258)) + ((g827) & (g1764) & (g3255) & (g3257) & (g3258)));
	assign g8238 = (((!g2017) & (g5921) & (!g3260)) + ((!g2017) & (g5921) & (g3260)) + ((g2017) & (!g5921) & (g3260)) + ((g2017) & (g5921) & (g3260)));
	assign g3261 = (((!g1732) & (g3199)) + ((g1732) & (!g3199)));
	assign g3262 = (((!g1665) & (!g1699) & (g3128) & (g3163) & (g3129) & (g3261)) + ((!g1665) & (g1699) & (!g3128) & (g3163) & (!g3129) & (g3261)) + ((!g1665) & (g1699) & (!g3128) & (g3163) & (g3129) & (g3261)) + ((!g1665) & (g1699) & (g3128) & (!g3163) & (g3129) & (g3261)) + ((!g1665) & (g1699) & (g3128) & (g3163) & (!g3129) & (g3261)) + ((!g1665) & (g1699) & (g3128) & (g3163) & (g3129) & (g3261)) + ((g1665) & (!g1699) & (!g3128) & (g3163) & (g3129) & (g3261)) + ((g1665) & (!g1699) & (g3128) & (g3163) & (!g3129) & (g3261)) + ((g1665) & (!g1699) & (g3128) & (g3163) & (g3129) & (g3261)) + ((g1665) & (g1699) & (!g3128) & (!g3163) & (g3129) & (g3261)) + ((g1665) & (g1699) & (!g3128) & (g3163) & (!g3129) & (g3261)) + ((g1665) & (g1699) & (!g3128) & (g3163) & (g3129) & (g3261)) + ((g1665) & (g1699) & (g3128) & (!g3163) & (!g3129) & (g3261)) + ((g1665) & (g1699) & (g3128) & (!g3163) & (g3129) & (g3261)) + ((g1665) & (g1699) & (g3128) & (g3163) & (!g3129) & (g3261)) + ((g1665) & (g1699) & (g3128) & (g3163) & (g3129) & (g3261)));
	assign g3263 = (((g1732) & (g3199)));
	assign g3264 = (((!g827) & (!g1766) & (g3260) & (!g3262) & (!g3263)) + ((!g827) & (!g1766) & (g3260) & (!g3262) & (g3263)) + ((!g827) & (!g1766) & (g3260) & (g3262) & (!g3263)) + ((!g827) & (!g1766) & (g3260) & (g3262) & (g3263)) + ((!g827) & (g1766) & (g3260) & (!g3262) & (!g3263)) + ((!g827) & (g1766) & (g3260) & (!g3262) & (g3263)) + ((!g827) & (g1766) & (g3260) & (g3262) & (!g3263)) + ((!g827) & (g1766) & (g3260) & (g3262) & (g3263)) + ((g827) & (!g1766) & (!g3260) & (!g3262) & (g3263)) + ((g827) & (!g1766) & (!g3260) & (g3262) & (!g3263)) + ((g827) & (!g1766) & (!g3260) & (g3262) & (g3263)) + ((g827) & (!g1766) & (g3260) & (!g3262) & (!g3263)) + ((g827) & (g1766) & (!g3260) & (!g3262) & (!g3263)) + ((g827) & (g1766) & (g3260) & (!g3262) & (g3263)) + ((g827) & (g1766) & (g3260) & (g3262) & (!g3263)) + ((g827) & (g1766) & (g3260) & (g3262) & (g3263)));
	assign g8239 = (((!g3429) & (g5441) & (!g3265)) + ((!g3429) & (g5441) & (g3265)) + ((g3429) & (!g5441) & (g3265)) + ((g3429) & (g5441) & (g3265)));
	assign g3266 = (((!g1740) & (g3210)) + ((g1740) & (!g3210)));
	assign g3267 = (((!g1673) & (!g1701) & (g3139) & (g3165) & (g3140) & (g3266)) + ((!g1673) & (g1701) & (!g3139) & (g3165) & (!g3140) & (g3266)) + ((!g1673) & (g1701) & (!g3139) & (g3165) & (g3140) & (g3266)) + ((!g1673) & (g1701) & (g3139) & (!g3165) & (g3140) & (g3266)) + ((!g1673) & (g1701) & (g3139) & (g3165) & (!g3140) & (g3266)) + ((!g1673) & (g1701) & (g3139) & (g3165) & (g3140) & (g3266)) + ((g1673) & (!g1701) & (!g3139) & (g3165) & (g3140) & (g3266)) + ((g1673) & (!g1701) & (g3139) & (g3165) & (!g3140) & (g3266)) + ((g1673) & (!g1701) & (g3139) & (g3165) & (g3140) & (g3266)) + ((g1673) & (g1701) & (!g3139) & (!g3165) & (g3140) & (g3266)) + ((g1673) & (g1701) & (!g3139) & (g3165) & (!g3140) & (g3266)) + ((g1673) & (g1701) & (!g3139) & (g3165) & (g3140) & (g3266)) + ((g1673) & (g1701) & (g3139) & (!g3165) & (!g3140) & (g3266)) + ((g1673) & (g1701) & (g3139) & (!g3165) & (g3140) & (g3266)) + ((g1673) & (g1701) & (g3139) & (g3165) & (!g3140) & (g3266)) + ((g1673) & (g1701) & (g3139) & (g3165) & (g3140) & (g3266)));
	assign g3268 = (((g1740) & (g3210)));
	assign g3269 = (((!g827) & (!g1768) & (g3265) & (!g3267) & (!g3268)) + ((!g827) & (!g1768) & (g3265) & (!g3267) & (g3268)) + ((!g827) & (!g1768) & (g3265) & (g3267) & (!g3268)) + ((!g827) & (!g1768) & (g3265) & (g3267) & (g3268)) + ((!g827) & (g1768) & (g3265) & (!g3267) & (!g3268)) + ((!g827) & (g1768) & (g3265) & (!g3267) & (g3268)) + ((!g827) & (g1768) & (g3265) & (g3267) & (!g3268)) + ((!g827) & (g1768) & (g3265) & (g3267) & (g3268)) + ((g827) & (!g1768) & (!g3265) & (!g3267) & (g3268)) + ((g827) & (!g1768) & (!g3265) & (g3267) & (!g3268)) + ((g827) & (!g1768) & (!g3265) & (g3267) & (g3268)) + ((g827) & (!g1768) & (g3265) & (!g3267) & (!g3268)) + ((g827) & (g1768) & (!g3265) & (!g3267) & (!g3268)) + ((g827) & (g1768) & (g3265) & (!g3267) & (g3268)) + ((g827) & (g1768) & (g3265) & (g3267) & (!g3268)) + ((g827) & (g1768) & (g3265) & (g3267) & (g3268)));
	assign g3270 = (((!g1718) & (g2599)) + ((g1718) & (!g2599)));
	assign g3271 = (((!g1651) & (!g1703) & (g2516) & (g2552) & (g3109) & (g3270)) + ((!g1651) & (g1703) & (!g2516) & (g2552) & (!g3109) & (g3270)) + ((!g1651) & (g1703) & (!g2516) & (g2552) & (g3109) & (g3270)) + ((!g1651) & (g1703) & (g2516) & (!g2552) & (g3109) & (g3270)) + ((!g1651) & (g1703) & (g2516) & (g2552) & (!g3109) & (g3270)) + ((!g1651) & (g1703) & (g2516) & (g2552) & (g3109) & (g3270)) + ((g1651) & (!g1703) & (!g2516) & (g2552) & (g3109) & (g3270)) + ((g1651) & (!g1703) & (g2516) & (g2552) & (!g3109) & (g3270)) + ((g1651) & (!g1703) & (g2516) & (g2552) & (g3109) & (g3270)) + ((g1651) & (g1703) & (!g2516) & (!g2552) & (g3109) & (g3270)) + ((g1651) & (g1703) & (!g2516) & (g2552) & (!g3109) & (g3270)) + ((g1651) & (g1703) & (!g2516) & (g2552) & (g3109) & (g3270)) + ((g1651) & (g1703) & (g2516) & (!g2552) & (!g3109) & (g3270)) + ((g1651) & (g1703) & (g2516) & (!g2552) & (g3109) & (g3270)) + ((g1651) & (g1703) & (g2516) & (g2552) & (!g3109) & (g3270)) + ((g1651) & (g1703) & (g2516) & (g2552) & (g3109) & (g3270)));
	assign g3272 = (((g1718) & (g2599)));
	assign g3273 = (((!g827) & (!g1770) & (g2648) & (!g3271) & (!g3272)) + ((!g827) & (!g1770) & (g2648) & (!g3271) & (g3272)) + ((!g827) & (!g1770) & (g2648) & (g3271) & (!g3272)) + ((!g827) & (!g1770) & (g2648) & (g3271) & (g3272)) + ((!g827) & (g1770) & (g2648) & (!g3271) & (!g3272)) + ((!g827) & (g1770) & (g2648) & (!g3271) & (g3272)) + ((!g827) & (g1770) & (g2648) & (g3271) & (!g3272)) + ((!g827) & (g1770) & (g2648) & (g3271) & (g3272)) + ((g827) & (!g1770) & (!g2648) & (!g3271) & (g3272)) + ((g827) & (!g1770) & (!g2648) & (g3271) & (!g3272)) + ((g827) & (!g1770) & (!g2648) & (g3271) & (g3272)) + ((g827) & (!g1770) & (g2648) & (!g3271) & (!g3272)) + ((g827) & (g1770) & (!g2648) & (!g3271) & (!g3272)) + ((g827) & (g1770) & (g2648) & (!g3271) & (g3272)) + ((g827) & (g1770) & (g2648) & (g3271) & (!g3272)) + ((g827) & (g1770) & (g2648) & (g3271) & (g3272)));
	assign g8240 = (((!g3499) & (g5445) & (!g3274)) + ((!g3499) & (g5445) & (g3274)) + ((g3499) & (!g5445) & (g3274)) + ((g3499) & (g5445) & (g3274)));
	assign g3275 = (((!g1726) & (g3190)) + ((g1726) & (!g3190)));
	assign g3276 = (((!g1659) & (!g1705) & (g3119) & (g3168) & (g3120) & (g3275)) + ((!g1659) & (g1705) & (!g3119) & (g3168) & (!g3120) & (g3275)) + ((!g1659) & (g1705) & (!g3119) & (g3168) & (g3120) & (g3275)) + ((!g1659) & (g1705) & (g3119) & (!g3168) & (g3120) & (g3275)) + ((!g1659) & (g1705) & (g3119) & (g3168) & (!g3120) & (g3275)) + ((!g1659) & (g1705) & (g3119) & (g3168) & (g3120) & (g3275)) + ((g1659) & (!g1705) & (!g3119) & (g3168) & (g3120) & (g3275)) + ((g1659) & (!g1705) & (g3119) & (g3168) & (!g3120) & (g3275)) + ((g1659) & (!g1705) & (g3119) & (g3168) & (g3120) & (g3275)) + ((g1659) & (g1705) & (!g3119) & (!g3168) & (g3120) & (g3275)) + ((g1659) & (g1705) & (!g3119) & (g3168) & (!g3120) & (g3275)) + ((g1659) & (g1705) & (!g3119) & (g3168) & (g3120) & (g3275)) + ((g1659) & (g1705) & (g3119) & (!g3168) & (!g3120) & (g3275)) + ((g1659) & (g1705) & (g3119) & (!g3168) & (g3120) & (g3275)) + ((g1659) & (g1705) & (g3119) & (g3168) & (!g3120) & (g3275)) + ((g1659) & (g1705) & (g3119) & (g3168) & (g3120) & (g3275)));
	assign g3277 = (((g1726) & (g3190)));
	assign g3278 = (((!g827) & (!g1772) & (g3274) & (!g3276) & (!g3277)) + ((!g827) & (!g1772) & (g3274) & (!g3276) & (g3277)) + ((!g827) & (!g1772) & (g3274) & (g3276) & (!g3277)) + ((!g827) & (!g1772) & (g3274) & (g3276) & (g3277)) + ((!g827) & (g1772) & (g3274) & (!g3276) & (!g3277)) + ((!g827) & (g1772) & (g3274) & (!g3276) & (g3277)) + ((!g827) & (g1772) & (g3274) & (g3276) & (!g3277)) + ((!g827) & (g1772) & (g3274) & (g3276) & (g3277)) + ((g827) & (!g1772) & (!g3274) & (!g3276) & (g3277)) + ((g827) & (!g1772) & (!g3274) & (g3276) & (!g3277)) + ((g827) & (!g1772) & (!g3274) & (g3276) & (g3277)) + ((g827) & (!g1772) & (g3274) & (!g3276) & (!g3277)) + ((g827) & (g1772) & (!g3274) & (!g3276) & (!g3277)) + ((g827) & (g1772) & (g3274) & (!g3276) & (g3277)) + ((g827) & (g1772) & (g3274) & (g3276) & (!g3277)) + ((g827) & (g1772) & (g3274) & (g3276) & (g3277)));
	assign g8241 = (((!g3429) & (g5450) & (!g3279)) + ((!g3429) & (g5450) & (g3279)) + ((g3429) & (!g5450) & (g3279)) + ((g3429) & (g5450) & (g3279)));
	assign g3280 = (((!g1734) & (g3202)) + ((g1734) & (!g3202)));
	assign g3281 = (((!g1667) & (!g1707) & (g3131) & (g3170) & (g3132) & (g3280)) + ((!g1667) & (g1707) & (!g3131) & (g3170) & (!g3132) & (g3280)) + ((!g1667) & (g1707) & (!g3131) & (g3170) & (g3132) & (g3280)) + ((!g1667) & (g1707) & (g3131) & (!g3170) & (g3132) & (g3280)) + ((!g1667) & (g1707) & (g3131) & (g3170) & (!g3132) & (g3280)) + ((!g1667) & (g1707) & (g3131) & (g3170) & (g3132) & (g3280)) + ((g1667) & (!g1707) & (!g3131) & (g3170) & (g3132) & (g3280)) + ((g1667) & (!g1707) & (g3131) & (g3170) & (!g3132) & (g3280)) + ((g1667) & (!g1707) & (g3131) & (g3170) & (g3132) & (g3280)) + ((g1667) & (g1707) & (!g3131) & (!g3170) & (g3132) & (g3280)) + ((g1667) & (g1707) & (!g3131) & (g3170) & (!g3132) & (g3280)) + ((g1667) & (g1707) & (!g3131) & (g3170) & (g3132) & (g3280)) + ((g1667) & (g1707) & (g3131) & (!g3170) & (!g3132) & (g3280)) + ((g1667) & (g1707) & (g3131) & (!g3170) & (g3132) & (g3280)) + ((g1667) & (g1707) & (g3131) & (g3170) & (!g3132) & (g3280)) + ((g1667) & (g1707) & (g3131) & (g3170) & (g3132) & (g3280)));
	assign g3282 = (((g1734) & (g3202)));
	assign g3283 = (((!g827) & (!g1774) & (g3279) & (!g3281) & (!g3282)) + ((!g827) & (!g1774) & (g3279) & (!g3281) & (g3282)) + ((!g827) & (!g1774) & (g3279) & (g3281) & (!g3282)) + ((!g827) & (!g1774) & (g3279) & (g3281) & (g3282)) + ((!g827) & (g1774) & (g3279) & (!g3281) & (!g3282)) + ((!g827) & (g1774) & (g3279) & (!g3281) & (g3282)) + ((!g827) & (g1774) & (g3279) & (g3281) & (!g3282)) + ((!g827) & (g1774) & (g3279) & (g3281) & (g3282)) + ((g827) & (!g1774) & (!g3279) & (!g3281) & (g3282)) + ((g827) & (!g1774) & (!g3279) & (g3281) & (!g3282)) + ((g827) & (!g1774) & (!g3279) & (g3281) & (g3282)) + ((g827) & (!g1774) & (g3279) & (!g3281) & (!g3282)) + ((g827) & (g1774) & (!g3279) & (!g3281) & (!g3282)) + ((g827) & (g1774) & (g3279) & (!g3281) & (g3282)) + ((g827) & (g1774) & (g3279) & (g3281) & (!g3282)) + ((g827) & (g1774) & (g3279) & (g3281) & (g3282)));
	assign g8242 = (((!g2017) & (g5915) & (!g3284)) + ((!g2017) & (g5915) & (g3284)) + ((g2017) & (!g5915) & (g3284)) + ((g2017) & (g5915) & (g3284)));
	assign g3285 = (((!g1742) & (g3213)) + ((g1742) & (!g3213)));
	assign g3286 = (((!g1675) & (!g1709) & (g3142) & (g3172) & (g3143) & (g3285)) + ((!g1675) & (g1709) & (!g3142) & (g3172) & (!g3143) & (g3285)) + ((!g1675) & (g1709) & (!g3142) & (g3172) & (g3143) & (g3285)) + ((!g1675) & (g1709) & (g3142) & (!g3172) & (g3143) & (g3285)) + ((!g1675) & (g1709) & (g3142) & (g3172) & (!g3143) & (g3285)) + ((!g1675) & (g1709) & (g3142) & (g3172) & (g3143) & (g3285)) + ((g1675) & (!g1709) & (!g3142) & (g3172) & (g3143) & (g3285)) + ((g1675) & (!g1709) & (g3142) & (g3172) & (!g3143) & (g3285)) + ((g1675) & (!g1709) & (g3142) & (g3172) & (g3143) & (g3285)) + ((g1675) & (g1709) & (!g3142) & (!g3172) & (g3143) & (g3285)) + ((g1675) & (g1709) & (!g3142) & (g3172) & (!g3143) & (g3285)) + ((g1675) & (g1709) & (!g3142) & (g3172) & (g3143) & (g3285)) + ((g1675) & (g1709) & (g3142) & (!g3172) & (!g3143) & (g3285)) + ((g1675) & (g1709) & (g3142) & (!g3172) & (g3143) & (g3285)) + ((g1675) & (g1709) & (g3142) & (g3172) & (!g3143) & (g3285)) + ((g1675) & (g1709) & (g3142) & (g3172) & (g3143) & (g3285)));
	assign g3287 = (((g1742) & (g3213)));
	assign g3288 = (((!g827) & (!g1776) & (g3284) & (!g3286) & (!g3287)) + ((!g827) & (!g1776) & (g3284) & (!g3286) & (g3287)) + ((!g827) & (!g1776) & (g3284) & (g3286) & (!g3287)) + ((!g827) & (!g1776) & (g3284) & (g3286) & (g3287)) + ((!g827) & (g1776) & (g3284) & (!g3286) & (!g3287)) + ((!g827) & (g1776) & (g3284) & (!g3286) & (g3287)) + ((!g827) & (g1776) & (g3284) & (g3286) & (!g3287)) + ((!g827) & (g1776) & (g3284) & (g3286) & (g3287)) + ((g827) & (!g1776) & (!g3284) & (!g3286) & (g3287)) + ((g827) & (!g1776) & (!g3284) & (g3286) & (!g3287)) + ((g827) & (!g1776) & (!g3284) & (g3286) & (g3287)) + ((g827) & (!g1776) & (g3284) & (!g3286) & (!g3287)) + ((g827) & (g1776) & (!g3284) & (!g3286) & (!g3287)) + ((g827) & (g1776) & (g3284) & (!g3286) & (g3287)) + ((g827) & (g1776) & (g3284) & (g3286) & (!g3287)) + ((g827) & (g1776) & (g3284) & (g3286) & (g3287)));
	assign g3289 = (((!g3216) & (!g1960) & (!g1961) & (!g1962) & (g1963)) + ((!g3216) & (!g1960) & (!g1961) & (g1962) & (!g1963)) + ((!g3216) & (!g1960) & (g1961) & (!g1962) & (g1963)) + ((!g3216) & (!g1960) & (g1961) & (g1962) & (!g1963)) + ((!g3216) & (g1960) & (!g1961) & (!g1962) & (g1963)) + ((!g3216) & (g1960) & (!g1961) & (g1962) & (!g1963)) + ((!g3216) & (g1960) & (g1961) & (!g1962) & (!g1963)) + ((!g3216) & (g1960) & (g1961) & (g1962) & (g1963)) + ((g3216) & (!g1960) & (!g1961) & (!g1962) & (g1963)) + ((g3216) & (!g1960) & (!g1961) & (g1962) & (!g1963)) + ((g3216) & (!g1960) & (g1961) & (!g1962) & (!g1963)) + ((g3216) & (!g1960) & (g1961) & (g1962) & (g1963)) + ((g3216) & (g1960) & (!g1961) & (!g1962) & (!g1963)) + ((g3216) & (g1960) & (!g1961) & (g1962) & (g1963)) + ((g3216) & (g1960) & (g1961) & (!g1962) & (!g1963)) + ((g3216) & (g1960) & (g1961) & (g1962) & (g1963)));
	assign g3290 = (((!g827) & (!g1754) & (!g2647) & (!g3232) & (!g3233) & (g5649)) + ((!g827) & (!g1754) & (!g2647) & (!g3232) & (g3233) & (g5649)) + ((!g827) & (!g1754) & (!g2647) & (g3232) & (!g3233) & (g5649)) + ((!g827) & (!g1754) & (!g2647) & (g3232) & (g3233) & (g5649)) + ((!g827) & (!g1754) & (g2647) & (!g3232) & (!g3233) & (g5649)) + ((!g827) & (!g1754) & (g2647) & (!g3232) & (g3233) & (g5649)) + ((!g827) & (!g1754) & (g2647) & (g3232) & (!g3233) & (g5649)) + ((!g827) & (!g1754) & (g2647) & (g3232) & (g3233) & (g5649)) + ((!g827) & (g1754) & (!g2647) & (!g3232) & (!g3233) & (g5649)) + ((!g827) & (g1754) & (!g2647) & (!g3232) & (g3233) & (g5649)) + ((!g827) & (g1754) & (!g2647) & (g3232) & (!g3233) & (g5649)) + ((!g827) & (g1754) & (!g2647) & (g3232) & (g3233) & (g5649)) + ((!g827) & (g1754) & (g2647) & (!g3232) & (!g3233) & (g5649)) + ((!g827) & (g1754) & (g2647) & (!g3232) & (g3233) & (g5649)) + ((!g827) & (g1754) & (g2647) & (g3232) & (!g3233) & (g5649)) + ((!g827) & (g1754) & (g2647) & (g3232) & (g3233) & (g5649)) + ((g827) & (!g1754) & (!g2647) & (!g3232) & (!g3233) & (!g5649)) + ((g827) & (!g1754) & (!g2647) & (!g3232) & (g3233) & (!g5649)) + ((g827) & (!g1754) & (!g2647) & (g3232) & (!g3233) & (!g5649)) + ((g827) & (!g1754) & (!g2647) & (g3232) & (g3233) & (!g5649)) + ((g827) & (!g1754) & (g2647) & (!g3232) & (!g3233) & (!g5649)) + ((g827) & (!g1754) & (g2647) & (!g3232) & (g3233) & (g5649)) + ((g827) & (!g1754) & (g2647) & (g3232) & (!g3233) & (g5649)) + ((g827) & (!g1754) & (g2647) & (g3232) & (g3233) & (g5649)) + ((g827) & (g1754) & (!g2647) & (!g3232) & (!g3233) & (!g5649)) + ((g827) & (g1754) & (!g2647) & (!g3232) & (g3233) & (g5649)) + ((g827) & (g1754) & (!g2647) & (g3232) & (!g3233) & (g5649)) + ((g827) & (g1754) & (!g2647) & (g3232) & (g3233) & (g5649)) + ((g827) & (g1754) & (g2647) & (!g3232) & (!g3233) & (g5649)) + ((g827) & (g1754) & (g2647) & (!g3232) & (g3233) & (g5649)) + ((g827) & (g1754) & (g2647) & (g3232) & (!g3233) & (g5649)) + ((g827) & (g1754) & (g2647) & (g3232) & (g3233) & (g5649)));
	assign g8243 = (((!g3499) & (g5454) & (!g3291)) + ((!g3499) & (g5454) & (g3291)) + ((g3499) & (!g5454) & (g3291)) + ((g3499) & (g5454) & (g3291)));
	assign g3292 = (((!g827) & (!g1762) & (!g3250) & (!g3252) & (!g3253) & (g5650)) + ((!g827) & (!g1762) & (!g3250) & (!g3252) & (g3253) & (g5650)) + ((!g827) & (!g1762) & (!g3250) & (g3252) & (!g3253) & (g5650)) + ((!g827) & (!g1762) & (!g3250) & (g3252) & (g3253) & (g5650)) + ((!g827) & (!g1762) & (g3250) & (!g3252) & (!g3253) & (g5650)) + ((!g827) & (!g1762) & (g3250) & (!g3252) & (g3253) & (g5650)) + ((!g827) & (!g1762) & (g3250) & (g3252) & (!g3253) & (g5650)) + ((!g827) & (!g1762) & (g3250) & (g3252) & (g3253) & (g5650)) + ((!g827) & (g1762) & (!g3250) & (!g3252) & (!g3253) & (g5650)) + ((!g827) & (g1762) & (!g3250) & (!g3252) & (g3253) & (g5650)) + ((!g827) & (g1762) & (!g3250) & (g3252) & (!g3253) & (g5650)) + ((!g827) & (g1762) & (!g3250) & (g3252) & (g3253) & (g5650)) + ((!g827) & (g1762) & (g3250) & (!g3252) & (!g3253) & (g5650)) + ((!g827) & (g1762) & (g3250) & (!g3252) & (g3253) & (g5650)) + ((!g827) & (g1762) & (g3250) & (g3252) & (!g3253) & (g5650)) + ((!g827) & (g1762) & (g3250) & (g3252) & (g3253) & (g5650)) + ((g827) & (!g1762) & (!g3250) & (!g3252) & (!g3253) & (!g5650)) + ((g827) & (!g1762) & (!g3250) & (!g3252) & (g3253) & (!g5650)) + ((g827) & (!g1762) & (!g3250) & (g3252) & (!g3253) & (!g5650)) + ((g827) & (!g1762) & (!g3250) & (g3252) & (g3253) & (!g5650)) + ((g827) & (!g1762) & (g3250) & (!g3252) & (!g3253) & (!g5650)) + ((g827) & (!g1762) & (g3250) & (!g3252) & (g3253) & (g5650)) + ((g827) & (!g1762) & (g3250) & (g3252) & (!g3253) & (g5650)) + ((g827) & (!g1762) & (g3250) & (g3252) & (g3253) & (g5650)) + ((g827) & (g1762) & (!g3250) & (!g3252) & (!g3253) & (!g5650)) + ((g827) & (g1762) & (!g3250) & (!g3252) & (g3253) & (g5650)) + ((g827) & (g1762) & (!g3250) & (g3252) & (!g3253) & (g5650)) + ((g827) & (g1762) & (!g3250) & (g3252) & (g3253) & (g5650)) + ((g827) & (g1762) & (g3250) & (!g3252) & (!g3253) & (g5650)) + ((g827) & (g1762) & (g3250) & (!g3252) & (g3253) & (g5650)) + ((g827) & (g1762) & (g3250) & (g3252) & (!g3253) & (g5650)) + ((g827) & (g1762) & (g3250) & (g3252) & (g3253) & (g5650)));
	assign g3293 = (((!g827) & (!g1770) & (!g2648) & (!g3271) & (!g3272) & (g5651)) + ((!g827) & (!g1770) & (!g2648) & (!g3271) & (g3272) & (g5651)) + ((!g827) & (!g1770) & (!g2648) & (g3271) & (!g3272) & (g5651)) + ((!g827) & (!g1770) & (!g2648) & (g3271) & (g3272) & (g5651)) + ((!g827) & (!g1770) & (g2648) & (!g3271) & (!g3272) & (g5651)) + ((!g827) & (!g1770) & (g2648) & (!g3271) & (g3272) & (g5651)) + ((!g827) & (!g1770) & (g2648) & (g3271) & (!g3272) & (g5651)) + ((!g827) & (!g1770) & (g2648) & (g3271) & (g3272) & (g5651)) + ((!g827) & (g1770) & (!g2648) & (!g3271) & (!g3272) & (g5651)) + ((!g827) & (g1770) & (!g2648) & (!g3271) & (g3272) & (g5651)) + ((!g827) & (g1770) & (!g2648) & (g3271) & (!g3272) & (g5651)) + ((!g827) & (g1770) & (!g2648) & (g3271) & (g3272) & (g5651)) + ((!g827) & (g1770) & (g2648) & (!g3271) & (!g3272) & (g5651)) + ((!g827) & (g1770) & (g2648) & (!g3271) & (g3272) & (g5651)) + ((!g827) & (g1770) & (g2648) & (g3271) & (!g3272) & (g5651)) + ((!g827) & (g1770) & (g2648) & (g3271) & (g3272) & (g5651)) + ((g827) & (!g1770) & (!g2648) & (!g3271) & (!g3272) & (!g5651)) + ((g827) & (!g1770) & (!g2648) & (!g3271) & (g3272) & (!g5651)) + ((g827) & (!g1770) & (!g2648) & (g3271) & (!g3272) & (!g5651)) + ((g827) & (!g1770) & (!g2648) & (g3271) & (g3272) & (!g5651)) + ((g827) & (!g1770) & (g2648) & (!g3271) & (!g3272) & (!g5651)) + ((g827) & (!g1770) & (g2648) & (!g3271) & (g3272) & (g5651)) + ((g827) & (!g1770) & (g2648) & (g3271) & (!g3272) & (g5651)) + ((g827) & (!g1770) & (g2648) & (g3271) & (g3272) & (g5651)) + ((g827) & (g1770) & (!g2648) & (!g3271) & (!g3272) & (!g5651)) + ((g827) & (g1770) & (!g2648) & (!g3271) & (g3272) & (g5651)) + ((g827) & (g1770) & (!g2648) & (g3271) & (!g3272) & (g5651)) + ((g827) & (g1770) & (!g2648) & (g3271) & (g3272) & (g5651)) + ((g827) & (g1770) & (g2648) & (!g3271) & (!g3272) & (g5651)) + ((g827) & (g1770) & (g2648) & (!g3271) & (g3272) & (g5651)) + ((g827) & (g1770) & (g2648) & (g3271) & (!g3272) & (g5651)) + ((g827) & (g1770) & (g2648) & (g3271) & (g3272) & (g5651)));
	assign g3294 = (((!g827) & (!g1748) & (!g2649) & (!g3219) & (!g3220) & (g5652)) + ((!g827) & (!g1748) & (!g2649) & (!g3219) & (g3220) & (g5652)) + ((!g827) & (!g1748) & (!g2649) & (g3219) & (!g3220) & (g5652)) + ((!g827) & (!g1748) & (!g2649) & (g3219) & (g3220) & (g5652)) + ((!g827) & (!g1748) & (g2649) & (!g3219) & (!g3220) & (g5652)) + ((!g827) & (!g1748) & (g2649) & (!g3219) & (g3220) & (g5652)) + ((!g827) & (!g1748) & (g2649) & (g3219) & (!g3220) & (g5652)) + ((!g827) & (!g1748) & (g2649) & (g3219) & (g3220) & (g5652)) + ((!g827) & (g1748) & (!g2649) & (!g3219) & (!g3220) & (g5652)) + ((!g827) & (g1748) & (!g2649) & (!g3219) & (g3220) & (g5652)) + ((!g827) & (g1748) & (!g2649) & (g3219) & (!g3220) & (g5652)) + ((!g827) & (g1748) & (!g2649) & (g3219) & (g3220) & (g5652)) + ((!g827) & (g1748) & (g2649) & (!g3219) & (!g3220) & (g5652)) + ((!g827) & (g1748) & (g2649) & (!g3219) & (g3220) & (g5652)) + ((!g827) & (g1748) & (g2649) & (g3219) & (!g3220) & (g5652)) + ((!g827) & (g1748) & (g2649) & (g3219) & (g3220) & (g5652)) + ((g827) & (!g1748) & (!g2649) & (!g3219) & (!g3220) & (!g5652)) + ((g827) & (!g1748) & (!g2649) & (!g3219) & (g3220) & (!g5652)) + ((g827) & (!g1748) & (!g2649) & (g3219) & (!g3220) & (!g5652)) + ((g827) & (!g1748) & (!g2649) & (g3219) & (g3220) & (!g5652)) + ((g827) & (!g1748) & (g2649) & (!g3219) & (!g3220) & (!g5652)) + ((g827) & (!g1748) & (g2649) & (!g3219) & (g3220) & (g5652)) + ((g827) & (!g1748) & (g2649) & (g3219) & (!g3220) & (g5652)) + ((g827) & (!g1748) & (g2649) & (g3219) & (g3220) & (g5652)) + ((g827) & (g1748) & (!g2649) & (!g3219) & (!g3220) & (!g5652)) + ((g827) & (g1748) & (!g2649) & (!g3219) & (g3220) & (g5652)) + ((g827) & (g1748) & (!g2649) & (g3219) & (!g3220) & (g5652)) + ((g827) & (g1748) & (!g2649) & (g3219) & (g3220) & (g5652)) + ((g827) & (g1748) & (g2649) & (!g3219) & (!g3220) & (g5652)) + ((g827) & (g1748) & (g2649) & (!g3219) & (g3220) & (g5652)) + ((g827) & (g1748) & (g2649) & (g3219) & (!g3220) & (g5652)) + ((g827) & (g1748) & (g2649) & (g3219) & (g3220) & (g5652)));
	assign g8244 = (((!g2017) & (g5459) & (!g3295)) + ((!g2017) & (g5459) & (g3295)) + ((g2017) & (!g5459) & (g3295)) + ((g2017) & (g5459) & (g3295)));
	assign g3296 = (((!g827) & (!g1756) & (!g3235) & (!g3237) & (!g3238) & (g5653)) + ((!g827) & (!g1756) & (!g3235) & (!g3237) & (g3238) & (g5653)) + ((!g827) & (!g1756) & (!g3235) & (g3237) & (!g3238) & (g5653)) + ((!g827) & (!g1756) & (!g3235) & (g3237) & (g3238) & (g5653)) + ((!g827) & (!g1756) & (g3235) & (!g3237) & (!g3238) & (g5653)) + ((!g827) & (!g1756) & (g3235) & (!g3237) & (g3238) & (g5653)) + ((!g827) & (!g1756) & (g3235) & (g3237) & (!g3238) & (g5653)) + ((!g827) & (!g1756) & (g3235) & (g3237) & (g3238) & (g5653)) + ((!g827) & (g1756) & (!g3235) & (!g3237) & (!g3238) & (g5653)) + ((!g827) & (g1756) & (!g3235) & (!g3237) & (g3238) & (g5653)) + ((!g827) & (g1756) & (!g3235) & (g3237) & (!g3238) & (g5653)) + ((!g827) & (g1756) & (!g3235) & (g3237) & (g3238) & (g5653)) + ((!g827) & (g1756) & (g3235) & (!g3237) & (!g3238) & (g5653)) + ((!g827) & (g1756) & (g3235) & (!g3237) & (g3238) & (g5653)) + ((!g827) & (g1756) & (g3235) & (g3237) & (!g3238) & (g5653)) + ((!g827) & (g1756) & (g3235) & (g3237) & (g3238) & (g5653)) + ((g827) & (!g1756) & (!g3235) & (!g3237) & (!g3238) & (!g5653)) + ((g827) & (!g1756) & (!g3235) & (!g3237) & (g3238) & (!g5653)) + ((g827) & (!g1756) & (!g3235) & (g3237) & (!g3238) & (!g5653)) + ((g827) & (!g1756) & (!g3235) & (g3237) & (g3238) & (!g5653)) + ((g827) & (!g1756) & (g3235) & (!g3237) & (!g3238) & (!g5653)) + ((g827) & (!g1756) & (g3235) & (!g3237) & (g3238) & (g5653)) + ((g827) & (!g1756) & (g3235) & (g3237) & (!g3238) & (g5653)) + ((g827) & (!g1756) & (g3235) & (g3237) & (g3238) & (g5653)) + ((g827) & (g1756) & (!g3235) & (!g3237) & (!g3238) & (!g5653)) + ((g827) & (g1756) & (!g3235) & (!g3237) & (g3238) & (g5653)) + ((g827) & (g1756) & (!g3235) & (g3237) & (!g3238) & (g5653)) + ((g827) & (g1756) & (!g3235) & (g3237) & (g3238) & (g5653)) + ((g827) & (g1756) & (g3235) & (!g3237) & (!g3238) & (g5653)) + ((g827) & (g1756) & (g3235) & (!g3237) & (g3238) & (g5653)) + ((g827) & (g1756) & (g3235) & (g3237) & (!g3238) & (g5653)) + ((g827) & (g1756) & (g3235) & (g3237) & (g3238) & (g5653)));
	assign g8245 = (((!g3464) & (g5464) & (!g3297)) + ((!g3464) & (g5464) & (g3297)) + ((g3464) & (!g5464) & (g3297)) + ((g3464) & (g5464) & (g3297)));
	assign g3298 = (((!g827) & (!g1764) & (!g3255) & (!g3257) & (!g3258) & (g5654)) + ((!g827) & (!g1764) & (!g3255) & (!g3257) & (g3258) & (g5654)) + ((!g827) & (!g1764) & (!g3255) & (g3257) & (!g3258) & (g5654)) + ((!g827) & (!g1764) & (!g3255) & (g3257) & (g3258) & (g5654)) + ((!g827) & (!g1764) & (g3255) & (!g3257) & (!g3258) & (g5654)) + ((!g827) & (!g1764) & (g3255) & (!g3257) & (g3258) & (g5654)) + ((!g827) & (!g1764) & (g3255) & (g3257) & (!g3258) & (g5654)) + ((!g827) & (!g1764) & (g3255) & (g3257) & (g3258) & (g5654)) + ((!g827) & (g1764) & (!g3255) & (!g3257) & (!g3258) & (g5654)) + ((!g827) & (g1764) & (!g3255) & (!g3257) & (g3258) & (g5654)) + ((!g827) & (g1764) & (!g3255) & (g3257) & (!g3258) & (g5654)) + ((!g827) & (g1764) & (!g3255) & (g3257) & (g3258) & (g5654)) + ((!g827) & (g1764) & (g3255) & (!g3257) & (!g3258) & (g5654)) + ((!g827) & (g1764) & (g3255) & (!g3257) & (g3258) & (g5654)) + ((!g827) & (g1764) & (g3255) & (g3257) & (!g3258) & (g5654)) + ((!g827) & (g1764) & (g3255) & (g3257) & (g3258) & (g5654)) + ((g827) & (!g1764) & (!g3255) & (!g3257) & (!g3258) & (!g5654)) + ((g827) & (!g1764) & (!g3255) & (!g3257) & (g3258) & (!g5654)) + ((g827) & (!g1764) & (!g3255) & (g3257) & (!g3258) & (!g5654)) + ((g827) & (!g1764) & (!g3255) & (g3257) & (g3258) & (!g5654)) + ((g827) & (!g1764) & (g3255) & (!g3257) & (!g3258) & (!g5654)) + ((g827) & (!g1764) & (g3255) & (!g3257) & (g3258) & (g5654)) + ((g827) & (!g1764) & (g3255) & (g3257) & (!g3258) & (g5654)) + ((g827) & (!g1764) & (g3255) & (g3257) & (g3258) & (g5654)) + ((g827) & (g1764) & (!g3255) & (!g3257) & (!g3258) & (!g5654)) + ((g827) & (g1764) & (!g3255) & (!g3257) & (g3258) & (g5654)) + ((g827) & (g1764) & (!g3255) & (g3257) & (!g3258) & (g5654)) + ((g827) & (g1764) & (!g3255) & (g3257) & (g3258) & (g5654)) + ((g827) & (g1764) & (g3255) & (!g3257) & (!g3258) & (g5654)) + ((g827) & (g1764) & (g3255) & (!g3257) & (g3258) & (g5654)) + ((g827) & (g1764) & (g3255) & (g3257) & (!g3258) & (g5654)) + ((g827) & (g1764) & (g3255) & (g3257) & (g3258) & (g5654)));
	assign g8246 = (((!g3499) & (g5467) & (!g3299)) + ((!g3499) & (g5467) & (g3299)) + ((g3499) & (!g5467) & (g3299)) + ((g3499) & (g5467) & (g3299)));
	assign g3300 = (((!g827) & (!g1772) & (!g3274) & (!g3276) & (!g3277) & (g5655)) + ((!g827) & (!g1772) & (!g3274) & (!g3276) & (g3277) & (g5655)) + ((!g827) & (!g1772) & (!g3274) & (g3276) & (!g3277) & (g5655)) + ((!g827) & (!g1772) & (!g3274) & (g3276) & (g3277) & (g5655)) + ((!g827) & (!g1772) & (g3274) & (!g3276) & (!g3277) & (g5655)) + ((!g827) & (!g1772) & (g3274) & (!g3276) & (g3277) & (g5655)) + ((!g827) & (!g1772) & (g3274) & (g3276) & (!g3277) & (g5655)) + ((!g827) & (!g1772) & (g3274) & (g3276) & (g3277) & (g5655)) + ((!g827) & (g1772) & (!g3274) & (!g3276) & (!g3277) & (g5655)) + ((!g827) & (g1772) & (!g3274) & (!g3276) & (g3277) & (g5655)) + ((!g827) & (g1772) & (!g3274) & (g3276) & (!g3277) & (g5655)) + ((!g827) & (g1772) & (!g3274) & (g3276) & (g3277) & (g5655)) + ((!g827) & (g1772) & (g3274) & (!g3276) & (!g3277) & (g5655)) + ((!g827) & (g1772) & (g3274) & (!g3276) & (g3277) & (g5655)) + ((!g827) & (g1772) & (g3274) & (g3276) & (!g3277) & (g5655)) + ((!g827) & (g1772) & (g3274) & (g3276) & (g3277) & (g5655)) + ((g827) & (!g1772) & (!g3274) & (!g3276) & (!g3277) & (!g5655)) + ((g827) & (!g1772) & (!g3274) & (!g3276) & (g3277) & (!g5655)) + ((g827) & (!g1772) & (!g3274) & (g3276) & (!g3277) & (!g5655)) + ((g827) & (!g1772) & (!g3274) & (g3276) & (g3277) & (!g5655)) + ((g827) & (!g1772) & (g3274) & (!g3276) & (!g3277) & (!g5655)) + ((g827) & (!g1772) & (g3274) & (!g3276) & (g3277) & (g5655)) + ((g827) & (!g1772) & (g3274) & (g3276) & (!g3277) & (g5655)) + ((g827) & (!g1772) & (g3274) & (g3276) & (g3277) & (g5655)) + ((g827) & (g1772) & (!g3274) & (!g3276) & (!g3277) & (!g5655)) + ((g827) & (g1772) & (!g3274) & (!g3276) & (g3277) & (g5655)) + ((g827) & (g1772) & (!g3274) & (g3276) & (!g3277) & (g5655)) + ((g827) & (g1772) & (!g3274) & (g3276) & (g3277) & (g5655)) + ((g827) & (g1772) & (g3274) & (!g3276) & (!g3277) & (g5655)) + ((g827) & (g1772) & (g3274) & (!g3276) & (g3277) & (g5655)) + ((g827) & (g1772) & (g3274) & (g3276) & (!g3277) & (g5655)) + ((g827) & (g1772) & (g3274) & (g3276) & (g3277) & (g5655)));
	assign g8247 = (((!g3464) & (g5470) & (!g3301)) + ((!g3464) & (g5470) & (g3301)) + ((g3464) & (!g5470) & (g3301)) + ((g3464) & (g5470) & (g3301)));
	assign g3302 = (((!g827) & (!g1750) & (!g3222) & (!g3224) & (!g3225) & (g5656)) + ((!g827) & (!g1750) & (!g3222) & (!g3224) & (g3225) & (g5656)) + ((!g827) & (!g1750) & (!g3222) & (g3224) & (!g3225) & (g5656)) + ((!g827) & (!g1750) & (!g3222) & (g3224) & (g3225) & (g5656)) + ((!g827) & (!g1750) & (g3222) & (!g3224) & (!g3225) & (g5656)) + ((!g827) & (!g1750) & (g3222) & (!g3224) & (g3225) & (g5656)) + ((!g827) & (!g1750) & (g3222) & (g3224) & (!g3225) & (g5656)) + ((!g827) & (!g1750) & (g3222) & (g3224) & (g3225) & (g5656)) + ((!g827) & (g1750) & (!g3222) & (!g3224) & (!g3225) & (g5656)) + ((!g827) & (g1750) & (!g3222) & (!g3224) & (g3225) & (g5656)) + ((!g827) & (g1750) & (!g3222) & (g3224) & (!g3225) & (g5656)) + ((!g827) & (g1750) & (!g3222) & (g3224) & (g3225) & (g5656)) + ((!g827) & (g1750) & (g3222) & (!g3224) & (!g3225) & (g5656)) + ((!g827) & (g1750) & (g3222) & (!g3224) & (g3225) & (g5656)) + ((!g827) & (g1750) & (g3222) & (g3224) & (!g3225) & (g5656)) + ((!g827) & (g1750) & (g3222) & (g3224) & (g3225) & (g5656)) + ((g827) & (!g1750) & (!g3222) & (!g3224) & (!g3225) & (!g5656)) + ((g827) & (!g1750) & (!g3222) & (!g3224) & (g3225) & (!g5656)) + ((g827) & (!g1750) & (!g3222) & (g3224) & (!g3225) & (!g5656)) + ((g827) & (!g1750) & (!g3222) & (g3224) & (g3225) & (!g5656)) + ((g827) & (!g1750) & (g3222) & (!g3224) & (!g3225) & (!g5656)) + ((g827) & (!g1750) & (g3222) & (!g3224) & (g3225) & (g5656)) + ((g827) & (!g1750) & (g3222) & (g3224) & (!g3225) & (g5656)) + ((g827) & (!g1750) & (g3222) & (g3224) & (g3225) & (g5656)) + ((g827) & (g1750) & (!g3222) & (!g3224) & (!g3225) & (!g5656)) + ((g827) & (g1750) & (!g3222) & (!g3224) & (g3225) & (g5656)) + ((g827) & (g1750) & (!g3222) & (g3224) & (!g3225) & (g5656)) + ((g827) & (g1750) & (!g3222) & (g3224) & (g3225) & (g5656)) + ((g827) & (g1750) & (g3222) & (!g3224) & (!g3225) & (g5656)) + ((g827) & (g1750) & (g3222) & (!g3224) & (g3225) & (g5656)) + ((g827) & (g1750) & (g3222) & (g3224) & (!g3225) & (g5656)) + ((g827) & (g1750) & (g3222) & (g3224) & (g3225) & (g5656)));
	assign g8248 = (((!g3499) & (g5473) & (!g3303)) + ((!g3499) & (g5473) & (g3303)) + ((g3499) & (!g5473) & (g3303)) + ((g3499) & (g5473) & (g3303)));
	assign g3304 = (((!g827) & (!g1758) & (!g3240) & (!g3242) & (!g3243) & (g5657)) + ((!g827) & (!g1758) & (!g3240) & (!g3242) & (g3243) & (g5657)) + ((!g827) & (!g1758) & (!g3240) & (g3242) & (!g3243) & (g5657)) + ((!g827) & (!g1758) & (!g3240) & (g3242) & (g3243) & (g5657)) + ((!g827) & (!g1758) & (g3240) & (!g3242) & (!g3243) & (g5657)) + ((!g827) & (!g1758) & (g3240) & (!g3242) & (g3243) & (g5657)) + ((!g827) & (!g1758) & (g3240) & (g3242) & (!g3243) & (g5657)) + ((!g827) & (!g1758) & (g3240) & (g3242) & (g3243) & (g5657)) + ((!g827) & (g1758) & (!g3240) & (!g3242) & (!g3243) & (g5657)) + ((!g827) & (g1758) & (!g3240) & (!g3242) & (g3243) & (g5657)) + ((!g827) & (g1758) & (!g3240) & (g3242) & (!g3243) & (g5657)) + ((!g827) & (g1758) & (!g3240) & (g3242) & (g3243) & (g5657)) + ((!g827) & (g1758) & (g3240) & (!g3242) & (!g3243) & (g5657)) + ((!g827) & (g1758) & (g3240) & (!g3242) & (g3243) & (g5657)) + ((!g827) & (g1758) & (g3240) & (g3242) & (!g3243) & (g5657)) + ((!g827) & (g1758) & (g3240) & (g3242) & (g3243) & (g5657)) + ((g827) & (!g1758) & (!g3240) & (!g3242) & (!g3243) & (!g5657)) + ((g827) & (!g1758) & (!g3240) & (!g3242) & (g3243) & (!g5657)) + ((g827) & (!g1758) & (!g3240) & (g3242) & (!g3243) & (!g5657)) + ((g827) & (!g1758) & (!g3240) & (g3242) & (g3243) & (!g5657)) + ((g827) & (!g1758) & (g3240) & (!g3242) & (!g3243) & (!g5657)) + ((g827) & (!g1758) & (g3240) & (!g3242) & (g3243) & (g5657)) + ((g827) & (!g1758) & (g3240) & (g3242) & (!g3243) & (g5657)) + ((g827) & (!g1758) & (g3240) & (g3242) & (g3243) & (g5657)) + ((g827) & (g1758) & (!g3240) & (!g3242) & (!g3243) & (!g5657)) + ((g827) & (g1758) & (!g3240) & (!g3242) & (g3243) & (g5657)) + ((g827) & (g1758) & (!g3240) & (g3242) & (!g3243) & (g5657)) + ((g827) & (g1758) & (!g3240) & (g3242) & (g3243) & (g5657)) + ((g827) & (g1758) & (g3240) & (!g3242) & (!g3243) & (g5657)) + ((g827) & (g1758) & (g3240) & (!g3242) & (g3243) & (g5657)) + ((g827) & (g1758) & (g3240) & (g3242) & (!g3243) & (g5657)) + ((g827) & (g1758) & (g3240) & (g3242) & (g3243) & (g5657)));
	assign g8249 = (((!g2017) & (g5478) & (!g3305)) + ((!g2017) & (g5478) & (g3305)) + ((g2017) & (!g5478) & (g3305)) + ((g2017) & (g5478) & (g3305)));
	assign g3306 = (((!g827) & (!g1766) & (!g3260) & (!g3262) & (!g3263) & (g5658)) + ((!g827) & (!g1766) & (!g3260) & (!g3262) & (g3263) & (g5658)) + ((!g827) & (!g1766) & (!g3260) & (g3262) & (!g3263) & (g5658)) + ((!g827) & (!g1766) & (!g3260) & (g3262) & (g3263) & (g5658)) + ((!g827) & (!g1766) & (g3260) & (!g3262) & (!g3263) & (g5658)) + ((!g827) & (!g1766) & (g3260) & (!g3262) & (g3263) & (g5658)) + ((!g827) & (!g1766) & (g3260) & (g3262) & (!g3263) & (g5658)) + ((!g827) & (!g1766) & (g3260) & (g3262) & (g3263) & (g5658)) + ((!g827) & (g1766) & (!g3260) & (!g3262) & (!g3263) & (g5658)) + ((!g827) & (g1766) & (!g3260) & (!g3262) & (g3263) & (g5658)) + ((!g827) & (g1766) & (!g3260) & (g3262) & (!g3263) & (g5658)) + ((!g827) & (g1766) & (!g3260) & (g3262) & (g3263) & (g5658)) + ((!g827) & (g1766) & (g3260) & (!g3262) & (!g3263) & (g5658)) + ((!g827) & (g1766) & (g3260) & (!g3262) & (g3263) & (g5658)) + ((!g827) & (g1766) & (g3260) & (g3262) & (!g3263) & (g5658)) + ((!g827) & (g1766) & (g3260) & (g3262) & (g3263) & (g5658)) + ((g827) & (!g1766) & (!g3260) & (!g3262) & (!g3263) & (!g5658)) + ((g827) & (!g1766) & (!g3260) & (!g3262) & (g3263) & (!g5658)) + ((g827) & (!g1766) & (!g3260) & (g3262) & (!g3263) & (!g5658)) + ((g827) & (!g1766) & (!g3260) & (g3262) & (g3263) & (!g5658)) + ((g827) & (!g1766) & (g3260) & (!g3262) & (!g3263) & (!g5658)) + ((g827) & (!g1766) & (g3260) & (!g3262) & (g3263) & (g5658)) + ((g827) & (!g1766) & (g3260) & (g3262) & (!g3263) & (g5658)) + ((g827) & (!g1766) & (g3260) & (g3262) & (g3263) & (g5658)) + ((g827) & (g1766) & (!g3260) & (!g3262) & (!g3263) & (!g5658)) + ((g827) & (g1766) & (!g3260) & (!g3262) & (g3263) & (g5658)) + ((g827) & (g1766) & (!g3260) & (g3262) & (!g3263) & (g5658)) + ((g827) & (g1766) & (!g3260) & (g3262) & (g3263) & (g5658)) + ((g827) & (g1766) & (g3260) & (!g3262) & (!g3263) & (g5658)) + ((g827) & (g1766) & (g3260) & (!g3262) & (g3263) & (g5658)) + ((g827) & (g1766) & (g3260) & (g3262) & (!g3263) & (g5658)) + ((g827) & (g1766) & (g3260) & (g3262) & (g3263) & (g5658)));
	assign g8250 = (((!g3429) & (g5481) & (!g3307)) + ((!g3429) & (g5481) & (g3307)) + ((g3429) & (!g5481) & (g3307)) + ((g3429) & (g5481) & (g3307)));
	assign g3308 = (((!g827) & (!g1774) & (!g3279) & (!g3281) & (!g3282) & (g5659)) + ((!g827) & (!g1774) & (!g3279) & (!g3281) & (g3282) & (g5659)) + ((!g827) & (!g1774) & (!g3279) & (g3281) & (!g3282) & (g5659)) + ((!g827) & (!g1774) & (!g3279) & (g3281) & (g3282) & (g5659)) + ((!g827) & (!g1774) & (g3279) & (!g3281) & (!g3282) & (g5659)) + ((!g827) & (!g1774) & (g3279) & (!g3281) & (g3282) & (g5659)) + ((!g827) & (!g1774) & (g3279) & (g3281) & (!g3282) & (g5659)) + ((!g827) & (!g1774) & (g3279) & (g3281) & (g3282) & (g5659)) + ((!g827) & (g1774) & (!g3279) & (!g3281) & (!g3282) & (g5659)) + ((!g827) & (g1774) & (!g3279) & (!g3281) & (g3282) & (g5659)) + ((!g827) & (g1774) & (!g3279) & (g3281) & (!g3282) & (g5659)) + ((!g827) & (g1774) & (!g3279) & (g3281) & (g3282) & (g5659)) + ((!g827) & (g1774) & (g3279) & (!g3281) & (!g3282) & (g5659)) + ((!g827) & (g1774) & (g3279) & (!g3281) & (g3282) & (g5659)) + ((!g827) & (g1774) & (g3279) & (g3281) & (!g3282) & (g5659)) + ((!g827) & (g1774) & (g3279) & (g3281) & (g3282) & (g5659)) + ((g827) & (!g1774) & (!g3279) & (!g3281) & (!g3282) & (!g5659)) + ((g827) & (!g1774) & (!g3279) & (!g3281) & (g3282) & (!g5659)) + ((g827) & (!g1774) & (!g3279) & (g3281) & (!g3282) & (!g5659)) + ((g827) & (!g1774) & (!g3279) & (g3281) & (g3282) & (!g5659)) + ((g827) & (!g1774) & (g3279) & (!g3281) & (!g3282) & (!g5659)) + ((g827) & (!g1774) & (g3279) & (!g3281) & (g3282) & (g5659)) + ((g827) & (!g1774) & (g3279) & (g3281) & (!g3282) & (g5659)) + ((g827) & (!g1774) & (g3279) & (g3281) & (g3282) & (g5659)) + ((g827) & (g1774) & (!g3279) & (!g3281) & (!g3282) & (!g5659)) + ((g827) & (g1774) & (!g3279) & (!g3281) & (g3282) & (g5659)) + ((g827) & (g1774) & (!g3279) & (g3281) & (!g3282) & (g5659)) + ((g827) & (g1774) & (!g3279) & (g3281) & (g3282) & (g5659)) + ((g827) & (g1774) & (g3279) & (!g3281) & (!g3282) & (g5659)) + ((g827) & (g1774) & (g3279) & (!g3281) & (g3282) & (g5659)) + ((g827) & (g1774) & (g3279) & (g3281) & (!g3282) & (g5659)) + ((g827) & (g1774) & (g3279) & (g3281) & (g3282) & (g5659)));
	assign g3309 = (((!g827) & (!g1752) & (!g2650) & (!g3228) & (!g3229) & (g5660)) + ((!g827) & (!g1752) & (!g2650) & (!g3228) & (g3229) & (g5660)) + ((!g827) & (!g1752) & (!g2650) & (g3228) & (!g3229) & (g5660)) + ((!g827) & (!g1752) & (!g2650) & (g3228) & (g3229) & (g5660)) + ((!g827) & (!g1752) & (g2650) & (!g3228) & (!g3229) & (g5660)) + ((!g827) & (!g1752) & (g2650) & (!g3228) & (g3229) & (g5660)) + ((!g827) & (!g1752) & (g2650) & (g3228) & (!g3229) & (g5660)) + ((!g827) & (!g1752) & (g2650) & (g3228) & (g3229) & (g5660)) + ((!g827) & (g1752) & (!g2650) & (!g3228) & (!g3229) & (g5660)) + ((!g827) & (g1752) & (!g2650) & (!g3228) & (g3229) & (g5660)) + ((!g827) & (g1752) & (!g2650) & (g3228) & (!g3229) & (g5660)) + ((!g827) & (g1752) & (!g2650) & (g3228) & (g3229) & (g5660)) + ((!g827) & (g1752) & (g2650) & (!g3228) & (!g3229) & (g5660)) + ((!g827) & (g1752) & (g2650) & (!g3228) & (g3229) & (g5660)) + ((!g827) & (g1752) & (g2650) & (g3228) & (!g3229) & (g5660)) + ((!g827) & (g1752) & (g2650) & (g3228) & (g3229) & (g5660)) + ((g827) & (!g1752) & (!g2650) & (!g3228) & (!g3229) & (!g5660)) + ((g827) & (!g1752) & (!g2650) & (!g3228) & (g3229) & (!g5660)) + ((g827) & (!g1752) & (!g2650) & (g3228) & (!g3229) & (!g5660)) + ((g827) & (!g1752) & (!g2650) & (g3228) & (g3229) & (!g5660)) + ((g827) & (!g1752) & (g2650) & (!g3228) & (!g3229) & (!g5660)) + ((g827) & (!g1752) & (g2650) & (!g3228) & (g3229) & (g5660)) + ((g827) & (!g1752) & (g2650) & (g3228) & (!g3229) & (g5660)) + ((g827) & (!g1752) & (g2650) & (g3228) & (g3229) & (g5660)) + ((g827) & (g1752) & (!g2650) & (!g3228) & (!g3229) & (!g5660)) + ((g827) & (g1752) & (!g2650) & (!g3228) & (g3229) & (g5660)) + ((g827) & (g1752) & (!g2650) & (g3228) & (!g3229) & (g5660)) + ((g827) & (g1752) & (!g2650) & (g3228) & (g3229) & (g5660)) + ((g827) & (g1752) & (g2650) & (!g3228) & (!g3229) & (g5660)) + ((g827) & (g1752) & (g2650) & (!g3228) & (g3229) & (g5660)) + ((g827) & (g1752) & (g2650) & (g3228) & (!g3229) & (g5660)) + ((g827) & (g1752) & (g2650) & (g3228) & (g3229) & (g5660)));
	assign g8251 = (((!g3464) & (g5484) & (!g3310)) + ((!g3464) & (g5484) & (g3310)) + ((g3464) & (!g5484) & (g3310)) + ((g3464) & (g5484) & (g3310)));
	assign g3311 = (((!g827) & (!g1760) & (!g3245) & (!g3247) & (!g3248) & (g5661)) + ((!g827) & (!g1760) & (!g3245) & (!g3247) & (g3248) & (g5661)) + ((!g827) & (!g1760) & (!g3245) & (g3247) & (!g3248) & (g5661)) + ((!g827) & (!g1760) & (!g3245) & (g3247) & (g3248) & (g5661)) + ((!g827) & (!g1760) & (g3245) & (!g3247) & (!g3248) & (g5661)) + ((!g827) & (!g1760) & (g3245) & (!g3247) & (g3248) & (g5661)) + ((!g827) & (!g1760) & (g3245) & (g3247) & (!g3248) & (g5661)) + ((!g827) & (!g1760) & (g3245) & (g3247) & (g3248) & (g5661)) + ((!g827) & (g1760) & (!g3245) & (!g3247) & (!g3248) & (g5661)) + ((!g827) & (g1760) & (!g3245) & (!g3247) & (g3248) & (g5661)) + ((!g827) & (g1760) & (!g3245) & (g3247) & (!g3248) & (g5661)) + ((!g827) & (g1760) & (!g3245) & (g3247) & (g3248) & (g5661)) + ((!g827) & (g1760) & (g3245) & (!g3247) & (!g3248) & (g5661)) + ((!g827) & (g1760) & (g3245) & (!g3247) & (g3248) & (g5661)) + ((!g827) & (g1760) & (g3245) & (g3247) & (!g3248) & (g5661)) + ((!g827) & (g1760) & (g3245) & (g3247) & (g3248) & (g5661)) + ((g827) & (!g1760) & (!g3245) & (!g3247) & (!g3248) & (!g5661)) + ((g827) & (!g1760) & (!g3245) & (!g3247) & (g3248) & (!g5661)) + ((g827) & (!g1760) & (!g3245) & (g3247) & (!g3248) & (!g5661)) + ((g827) & (!g1760) & (!g3245) & (g3247) & (g3248) & (!g5661)) + ((g827) & (!g1760) & (g3245) & (!g3247) & (!g3248) & (!g5661)) + ((g827) & (!g1760) & (g3245) & (!g3247) & (g3248) & (g5661)) + ((g827) & (!g1760) & (g3245) & (g3247) & (!g3248) & (g5661)) + ((g827) & (!g1760) & (g3245) & (g3247) & (g3248) & (g5661)) + ((g827) & (g1760) & (!g3245) & (!g3247) & (!g3248) & (!g5661)) + ((g827) & (g1760) & (!g3245) & (!g3247) & (g3248) & (g5661)) + ((g827) & (g1760) & (!g3245) & (g3247) & (!g3248) & (g5661)) + ((g827) & (g1760) & (!g3245) & (g3247) & (g3248) & (g5661)) + ((g827) & (g1760) & (g3245) & (!g3247) & (!g3248) & (g5661)) + ((g827) & (g1760) & (g3245) & (!g3247) & (g3248) & (g5661)) + ((g827) & (g1760) & (g3245) & (g3247) & (!g3248) & (g5661)) + ((g827) & (g1760) & (g3245) & (g3247) & (g3248) & (g5661)));
	assign g8252 = (((!g3429) & (g5487) & (!g3312)) + ((!g3429) & (g5487) & (g3312)) + ((g3429) & (!g5487) & (g3312)) + ((g3429) & (g5487) & (g3312)));
	assign g3313 = (((!g827) & (!g1768) & (!g3265) & (!g3267) & (!g3268) & (g5662)) + ((!g827) & (!g1768) & (!g3265) & (!g3267) & (g3268) & (g5662)) + ((!g827) & (!g1768) & (!g3265) & (g3267) & (!g3268) & (g5662)) + ((!g827) & (!g1768) & (!g3265) & (g3267) & (g3268) & (g5662)) + ((!g827) & (!g1768) & (g3265) & (!g3267) & (!g3268) & (g5662)) + ((!g827) & (!g1768) & (g3265) & (!g3267) & (g3268) & (g5662)) + ((!g827) & (!g1768) & (g3265) & (g3267) & (!g3268) & (g5662)) + ((!g827) & (!g1768) & (g3265) & (g3267) & (g3268) & (g5662)) + ((!g827) & (g1768) & (!g3265) & (!g3267) & (!g3268) & (g5662)) + ((!g827) & (g1768) & (!g3265) & (!g3267) & (g3268) & (g5662)) + ((!g827) & (g1768) & (!g3265) & (g3267) & (!g3268) & (g5662)) + ((!g827) & (g1768) & (!g3265) & (g3267) & (g3268) & (g5662)) + ((!g827) & (g1768) & (g3265) & (!g3267) & (!g3268) & (g5662)) + ((!g827) & (g1768) & (g3265) & (!g3267) & (g3268) & (g5662)) + ((!g827) & (g1768) & (g3265) & (g3267) & (!g3268) & (g5662)) + ((!g827) & (g1768) & (g3265) & (g3267) & (g3268) & (g5662)) + ((g827) & (!g1768) & (!g3265) & (!g3267) & (!g3268) & (!g5662)) + ((g827) & (!g1768) & (!g3265) & (!g3267) & (g3268) & (!g5662)) + ((g827) & (!g1768) & (!g3265) & (g3267) & (!g3268) & (!g5662)) + ((g827) & (!g1768) & (!g3265) & (g3267) & (g3268) & (!g5662)) + ((g827) & (!g1768) & (g3265) & (!g3267) & (!g3268) & (!g5662)) + ((g827) & (!g1768) & (g3265) & (!g3267) & (g3268) & (g5662)) + ((g827) & (!g1768) & (g3265) & (g3267) & (!g3268) & (g5662)) + ((g827) & (!g1768) & (g3265) & (g3267) & (g3268) & (g5662)) + ((g827) & (g1768) & (!g3265) & (!g3267) & (!g3268) & (!g5662)) + ((g827) & (g1768) & (!g3265) & (!g3267) & (g3268) & (g5662)) + ((g827) & (g1768) & (!g3265) & (g3267) & (!g3268) & (g5662)) + ((g827) & (g1768) & (!g3265) & (g3267) & (g3268) & (g5662)) + ((g827) & (g1768) & (g3265) & (!g3267) & (!g3268) & (g5662)) + ((g827) & (g1768) & (g3265) & (!g3267) & (g3268) & (g5662)) + ((g827) & (g1768) & (g3265) & (g3267) & (!g3268) & (g5662)) + ((g827) & (g1768) & (g3265) & (g3267) & (g3268) & (g5662)));
	assign g8253 = (((!g2017) & (g5492) & (!g3314)) + ((!g2017) & (g5492) & (g3314)) + ((g2017) & (!g5492) & (g3314)) + ((g2017) & (g5492) & (g3314)));
	assign g3315 = (((!g827) & (!g1776) & (!g3284) & (!g3286) & (!g3287) & (g5663)) + ((!g827) & (!g1776) & (!g3284) & (!g3286) & (g3287) & (g5663)) + ((!g827) & (!g1776) & (!g3284) & (g3286) & (!g3287) & (g5663)) + ((!g827) & (!g1776) & (!g3284) & (g3286) & (g3287) & (g5663)) + ((!g827) & (!g1776) & (g3284) & (!g3286) & (!g3287) & (g5663)) + ((!g827) & (!g1776) & (g3284) & (!g3286) & (g3287) & (g5663)) + ((!g827) & (!g1776) & (g3284) & (g3286) & (!g3287) & (g5663)) + ((!g827) & (!g1776) & (g3284) & (g3286) & (g3287) & (g5663)) + ((!g827) & (g1776) & (!g3284) & (!g3286) & (!g3287) & (g5663)) + ((!g827) & (g1776) & (!g3284) & (!g3286) & (g3287) & (g5663)) + ((!g827) & (g1776) & (!g3284) & (g3286) & (!g3287) & (g5663)) + ((!g827) & (g1776) & (!g3284) & (g3286) & (g3287) & (g5663)) + ((!g827) & (g1776) & (g3284) & (!g3286) & (!g3287) & (g5663)) + ((!g827) & (g1776) & (g3284) & (!g3286) & (g3287) & (g5663)) + ((!g827) & (g1776) & (g3284) & (g3286) & (!g3287) & (g5663)) + ((!g827) & (g1776) & (g3284) & (g3286) & (g3287) & (g5663)) + ((g827) & (!g1776) & (!g3284) & (!g3286) & (!g3287) & (!g5663)) + ((g827) & (!g1776) & (!g3284) & (!g3286) & (g3287) & (!g5663)) + ((g827) & (!g1776) & (!g3284) & (g3286) & (!g3287) & (!g5663)) + ((g827) & (!g1776) & (!g3284) & (g3286) & (g3287) & (!g5663)) + ((g827) & (!g1776) & (g3284) & (!g3286) & (!g3287) & (!g5663)) + ((g827) & (!g1776) & (g3284) & (!g3286) & (g3287) & (g5663)) + ((g827) & (!g1776) & (g3284) & (g3286) & (!g3287) & (g5663)) + ((g827) & (!g1776) & (g3284) & (g3286) & (g3287) & (g5663)) + ((g827) & (g1776) & (!g3284) & (!g3286) & (!g3287) & (!g5663)) + ((g827) & (g1776) & (!g3284) & (!g3286) & (g3287) & (g5663)) + ((g827) & (g1776) & (!g3284) & (g3286) & (!g3287) & (g5663)) + ((g827) & (g1776) & (!g3284) & (g3286) & (g3287) & (g5663)) + ((g827) & (g1776) & (g3284) & (!g3286) & (!g3287) & (g5663)) + ((g827) & (g1776) & (g3284) & (!g3286) & (g3287) & (g5663)) + ((g827) & (g1776) & (g3284) & (g3286) & (!g3287) & (g5663)) + ((g827) & (g1776) & (g3284) & (g3286) & (g3287) & (g5663)));
	assign g3316 = (((!g1965) & (!g1966)));
	assign g3317 = (((g1914) & (!g3316) & (!g1967) & (!g1968)) + ((g1914) & (!g3316) & (g1967) & (g1968)) + ((g1914) & (g3316) & (!g1967) & (g1968)) + ((g1914) & (g3316) & (g1967) & (!g1968)));
	assign g3318 = (((!g2000) & (g2001) & (g2002)) + ((g2000) & (!g2001) & (g2002)) + ((g2000) & (g2001) & (!g2002)) + ((g2000) & (g2001) & (g2002)));
	assign g3319 = (((!g1914) & (!g3318) & (!g2003) & (g2004)) + ((!g1914) & (!g3318) & (g2003) & (!g2004)) + ((!g1914) & (g3318) & (!g2003) & (!g2004)) + ((!g1914) & (g3318) & (g2003) & (g2004)));
	assign g3320 = (((!g830) & (!g3317) & (!g3319) & (!g1814)) + ((!g830) & (!g3317) & (!g3319) & (g1814)) + ((!g830) & (!g3317) & (g3319) & (!g1814)) + ((!g830) & (!g3317) & (g3319) & (g1814)) + ((!g830) & (g3317) & (!g3319) & (!g1814)) + ((!g830) & (g3317) & (!g3319) & (g1814)) + ((!g830) & (g3317) & (g3319) & (!g1814)) + ((!g830) & (g3317) & (g3319) & (g1814)) + ((g830) & (!g3317) & (!g3319) & (g1814)) + ((g830) & (!g3317) & (g3319) & (!g1814)) + ((g830) & (g3317) & (!g3319) & (!g1814)) + ((g830) & (g3317) & (g3319) & (!g1814)));
	assign g3321 = (((!g1748) & (!g1790) & (!g2649) & (!g2683) & (!g3219) & (!g3220)) + ((!g1748) & (!g1790) & (!g2649) & (!g2683) & (!g3219) & (g3220)) + ((!g1748) & (!g1790) & (!g2649) & (!g2683) & (g3219) & (!g3220)) + ((!g1748) & (!g1790) & (!g2649) & (!g2683) & (g3219) & (g3220)) + ((!g1748) & (!g1790) & (!g2649) & (g2683) & (!g3219) & (!g3220)) + ((!g1748) & (!g1790) & (!g2649) & (g2683) & (!g3219) & (g3220)) + ((!g1748) & (!g1790) & (!g2649) & (g2683) & (g3219) & (!g3220)) + ((!g1748) & (!g1790) & (!g2649) & (g2683) & (g3219) & (g3220)) + ((!g1748) & (!g1790) & (g2649) & (!g2683) & (!g3219) & (!g3220)) + ((!g1748) & (!g1790) & (g2649) & (!g2683) & (!g3219) & (g3220)) + ((!g1748) & (!g1790) & (g2649) & (!g2683) & (g3219) & (!g3220)) + ((!g1748) & (!g1790) & (g2649) & (!g2683) & (g3219) & (g3220)) + ((!g1748) & (!g1790) & (g2649) & (g2683) & (!g3219) & (!g3220)) + ((!g1748) & (g1790) & (!g2649) & (!g2683) & (!g3219) & (!g3220)) + ((!g1748) & (g1790) & (!g2649) & (!g2683) & (!g3219) & (g3220)) + ((!g1748) & (g1790) & (!g2649) & (!g2683) & (g3219) & (!g3220)) + ((!g1748) & (g1790) & (!g2649) & (!g2683) & (g3219) & (g3220)) + ((!g1748) & (g1790) & (g2649) & (!g2683) & (!g3219) & (!g3220)) + ((g1748) & (!g1790) & (!g2649) & (!g2683) & (!g3219) & (!g3220)) + ((g1748) & (!g1790) & (!g2649) & (!g2683) & (!g3219) & (g3220)) + ((g1748) & (!g1790) & (!g2649) & (!g2683) & (g3219) & (!g3220)) + ((g1748) & (!g1790) & (!g2649) & (!g2683) & (g3219) & (g3220)) + ((g1748) & (!g1790) & (!g2649) & (g2683) & (!g3219) & (!g3220)) + ((g1748) & (!g1790) & (g2649) & (!g2683) & (!g3219) & (!g3220)) + ((g1748) & (!g1790) & (g2649) & (!g2683) & (!g3219) & (g3220)) + ((g1748) & (!g1790) & (g2649) & (!g2683) & (g3219) & (!g3220)) + ((g1748) & (!g1790) & (g2649) & (!g2683) & (g3219) & (g3220)) + ((g1748) & (g1790) & (!g2649) & (!g2683) & (!g3219) & (!g3220)));
	assign g3322 = (((!g827) & (!g1817) & (g2760) & (!g3321)) + ((!g827) & (!g1817) & (g2760) & (g3321)) + ((!g827) & (g1817) & (g2760) & (!g3321)) + ((!g827) & (g1817) & (g2760) & (g3321)) + ((g827) & (!g1817) & (!g2760) & (!g3321)) + ((g827) & (!g1817) & (g2760) & (g3321)) + ((g827) & (g1817) & (!g2760) & (g3321)) + ((g827) & (g1817) & (g2760) & (!g3321)));
	assign g8254 = (((!g3464) & (g5495) & (!g3323)) + ((!g3464) & (g5495) & (g3323)) + ((g3464) & (!g5495) & (g3323)) + ((g3464) & (g5495) & (g3323)));
	assign g3324 = (((!g1750) & (!g1798) & (!g3222) & (!g3301) & (!g3224) & (!g3225)) + ((!g1750) & (!g1798) & (!g3222) & (!g3301) & (!g3224) & (g3225)) + ((!g1750) & (!g1798) & (!g3222) & (!g3301) & (g3224) & (!g3225)) + ((!g1750) & (!g1798) & (!g3222) & (!g3301) & (g3224) & (g3225)) + ((!g1750) & (!g1798) & (!g3222) & (g3301) & (!g3224) & (!g3225)) + ((!g1750) & (!g1798) & (!g3222) & (g3301) & (!g3224) & (g3225)) + ((!g1750) & (!g1798) & (!g3222) & (g3301) & (g3224) & (!g3225)) + ((!g1750) & (!g1798) & (!g3222) & (g3301) & (g3224) & (g3225)) + ((!g1750) & (!g1798) & (g3222) & (!g3301) & (!g3224) & (!g3225)) + ((!g1750) & (!g1798) & (g3222) & (!g3301) & (!g3224) & (g3225)) + ((!g1750) & (!g1798) & (g3222) & (!g3301) & (g3224) & (!g3225)) + ((!g1750) & (!g1798) & (g3222) & (!g3301) & (g3224) & (g3225)) + ((!g1750) & (!g1798) & (g3222) & (g3301) & (!g3224) & (!g3225)) + ((!g1750) & (g1798) & (!g3222) & (!g3301) & (!g3224) & (!g3225)) + ((!g1750) & (g1798) & (!g3222) & (!g3301) & (!g3224) & (g3225)) + ((!g1750) & (g1798) & (!g3222) & (!g3301) & (g3224) & (!g3225)) + ((!g1750) & (g1798) & (!g3222) & (!g3301) & (g3224) & (g3225)) + ((!g1750) & (g1798) & (g3222) & (!g3301) & (!g3224) & (!g3225)) + ((g1750) & (!g1798) & (!g3222) & (!g3301) & (!g3224) & (!g3225)) + ((g1750) & (!g1798) & (!g3222) & (!g3301) & (!g3224) & (g3225)) + ((g1750) & (!g1798) & (!g3222) & (!g3301) & (g3224) & (!g3225)) + ((g1750) & (!g1798) & (!g3222) & (!g3301) & (g3224) & (g3225)) + ((g1750) & (!g1798) & (!g3222) & (g3301) & (!g3224) & (!g3225)) + ((g1750) & (!g1798) & (g3222) & (!g3301) & (!g3224) & (!g3225)) + ((g1750) & (!g1798) & (g3222) & (!g3301) & (!g3224) & (g3225)) + ((g1750) & (!g1798) & (g3222) & (!g3301) & (g3224) & (!g3225)) + ((g1750) & (!g1798) & (g3222) & (!g3301) & (g3224) & (g3225)) + ((g1750) & (g1798) & (!g3222) & (!g3301) & (!g3224) & (!g3225)));
	assign g3325 = (((!g827) & (!g1819) & (g3323) & (!g3324)) + ((!g827) & (!g1819) & (g3323) & (g3324)) + ((!g827) & (g1819) & (g3323) & (!g3324)) + ((!g827) & (g1819) & (g3323) & (g3324)) + ((g827) & (!g1819) & (!g3323) & (!g3324)) + ((g827) & (!g1819) & (g3323) & (g3324)) + ((g827) & (g1819) & (!g3323) & (g3324)) + ((g827) & (g1819) & (g3323) & (!g3324)));
	assign g3326 = (((!g1752) & (!g1806) & (!g2650) & (!g2684) & (!g3228) & (!g3229)) + ((!g1752) & (!g1806) & (!g2650) & (!g2684) & (!g3228) & (g3229)) + ((!g1752) & (!g1806) & (!g2650) & (!g2684) & (g3228) & (!g3229)) + ((!g1752) & (!g1806) & (!g2650) & (!g2684) & (g3228) & (g3229)) + ((!g1752) & (!g1806) & (!g2650) & (g2684) & (!g3228) & (!g3229)) + ((!g1752) & (!g1806) & (!g2650) & (g2684) & (!g3228) & (g3229)) + ((!g1752) & (!g1806) & (!g2650) & (g2684) & (g3228) & (!g3229)) + ((!g1752) & (!g1806) & (!g2650) & (g2684) & (g3228) & (g3229)) + ((!g1752) & (!g1806) & (g2650) & (!g2684) & (!g3228) & (!g3229)) + ((!g1752) & (!g1806) & (g2650) & (!g2684) & (!g3228) & (g3229)) + ((!g1752) & (!g1806) & (g2650) & (!g2684) & (g3228) & (!g3229)) + ((!g1752) & (!g1806) & (g2650) & (!g2684) & (g3228) & (g3229)) + ((!g1752) & (!g1806) & (g2650) & (g2684) & (!g3228) & (!g3229)) + ((!g1752) & (g1806) & (!g2650) & (!g2684) & (!g3228) & (!g3229)) + ((!g1752) & (g1806) & (!g2650) & (!g2684) & (!g3228) & (g3229)) + ((!g1752) & (g1806) & (!g2650) & (!g2684) & (g3228) & (!g3229)) + ((!g1752) & (g1806) & (!g2650) & (!g2684) & (g3228) & (g3229)) + ((!g1752) & (g1806) & (g2650) & (!g2684) & (!g3228) & (!g3229)) + ((g1752) & (!g1806) & (!g2650) & (!g2684) & (!g3228) & (!g3229)) + ((g1752) & (!g1806) & (!g2650) & (!g2684) & (!g3228) & (g3229)) + ((g1752) & (!g1806) & (!g2650) & (!g2684) & (g3228) & (!g3229)) + ((g1752) & (!g1806) & (!g2650) & (!g2684) & (g3228) & (g3229)) + ((g1752) & (!g1806) & (!g2650) & (g2684) & (!g3228) & (!g3229)) + ((g1752) & (!g1806) & (g2650) & (!g2684) & (!g3228) & (!g3229)) + ((g1752) & (!g1806) & (g2650) & (!g2684) & (!g3228) & (g3229)) + ((g1752) & (!g1806) & (g2650) & (!g2684) & (g3228) & (!g3229)) + ((g1752) & (!g1806) & (g2650) & (!g2684) & (g3228) & (g3229)) + ((g1752) & (g1806) & (!g2650) & (!g2684) & (!g3228) & (!g3229)));
	assign g3327 = (((!g827) & (!g1821) & (g2761) & (!g3326)) + ((!g827) & (!g1821) & (g2761) & (g3326)) + ((!g827) & (g1821) & (g2761) & (!g3326)) + ((!g827) & (g1821) & (g2761) & (g3326)) + ((g827) & (!g1821) & (!g2761) & (!g3326)) + ((g827) & (!g1821) & (g2761) & (g3326)) + ((g827) & (g1821) & (!g2761) & (g3326)) + ((g827) & (g1821) & (g2761) & (!g3326)));
	assign g3328 = (((!g1754) & (!g1784) & (!g2647) & (!g2678) & (!g3232) & (!g3233)) + ((!g1754) & (!g1784) & (!g2647) & (!g2678) & (!g3232) & (g3233)) + ((!g1754) & (!g1784) & (!g2647) & (!g2678) & (g3232) & (!g3233)) + ((!g1754) & (!g1784) & (!g2647) & (!g2678) & (g3232) & (g3233)) + ((!g1754) & (!g1784) & (!g2647) & (g2678) & (!g3232) & (!g3233)) + ((!g1754) & (!g1784) & (!g2647) & (g2678) & (!g3232) & (g3233)) + ((!g1754) & (!g1784) & (!g2647) & (g2678) & (g3232) & (!g3233)) + ((!g1754) & (!g1784) & (!g2647) & (g2678) & (g3232) & (g3233)) + ((!g1754) & (!g1784) & (g2647) & (!g2678) & (!g3232) & (!g3233)) + ((!g1754) & (!g1784) & (g2647) & (!g2678) & (!g3232) & (g3233)) + ((!g1754) & (!g1784) & (g2647) & (!g2678) & (g3232) & (!g3233)) + ((!g1754) & (!g1784) & (g2647) & (!g2678) & (g3232) & (g3233)) + ((!g1754) & (!g1784) & (g2647) & (g2678) & (!g3232) & (!g3233)) + ((!g1754) & (g1784) & (!g2647) & (!g2678) & (!g3232) & (!g3233)) + ((!g1754) & (g1784) & (!g2647) & (!g2678) & (!g3232) & (g3233)) + ((!g1754) & (g1784) & (!g2647) & (!g2678) & (g3232) & (!g3233)) + ((!g1754) & (g1784) & (!g2647) & (!g2678) & (g3232) & (g3233)) + ((!g1754) & (g1784) & (g2647) & (!g2678) & (!g3232) & (!g3233)) + ((g1754) & (!g1784) & (!g2647) & (!g2678) & (!g3232) & (!g3233)) + ((g1754) & (!g1784) & (!g2647) & (!g2678) & (!g3232) & (g3233)) + ((g1754) & (!g1784) & (!g2647) & (!g2678) & (g3232) & (!g3233)) + ((g1754) & (!g1784) & (!g2647) & (!g2678) & (g3232) & (g3233)) + ((g1754) & (!g1784) & (!g2647) & (g2678) & (!g3232) & (!g3233)) + ((g1754) & (!g1784) & (g2647) & (!g2678) & (!g3232) & (!g3233)) + ((g1754) & (!g1784) & (g2647) & (!g2678) & (!g3232) & (g3233)) + ((g1754) & (!g1784) & (g2647) & (!g2678) & (g3232) & (!g3233)) + ((g1754) & (!g1784) & (g2647) & (!g2678) & (g3232) & (g3233)) + ((g1754) & (g1784) & (!g2647) & (!g2678) & (!g3232) & (!g3233)));
	assign g3329 = (((!g827) & (!g1823) & (g2758) & (!g3328)) + ((!g827) & (!g1823) & (g2758) & (g3328)) + ((!g827) & (g1823) & (g2758) & (!g3328)) + ((!g827) & (g1823) & (g2758) & (g3328)) + ((g827) & (!g1823) & (!g2758) & (!g3328)) + ((g827) & (!g1823) & (g2758) & (g3328)) + ((g827) & (g1823) & (!g2758) & (g3328)) + ((g827) & (g1823) & (g2758) & (!g3328)));
	assign g8255 = (((!g2017) & (g5498) & (!g3330)) + ((!g2017) & (g5498) & (g3330)) + ((g2017) & (!g5498) & (g3330)) + ((g2017) & (g5498) & (g3330)));
	assign g3331 = (((!g1756) & (!g1792) & (!g3235) & (!g3295) & (!g3237) & (!g3238)) + ((!g1756) & (!g1792) & (!g3235) & (!g3295) & (!g3237) & (g3238)) + ((!g1756) & (!g1792) & (!g3235) & (!g3295) & (g3237) & (!g3238)) + ((!g1756) & (!g1792) & (!g3235) & (!g3295) & (g3237) & (g3238)) + ((!g1756) & (!g1792) & (!g3235) & (g3295) & (!g3237) & (!g3238)) + ((!g1756) & (!g1792) & (!g3235) & (g3295) & (!g3237) & (g3238)) + ((!g1756) & (!g1792) & (!g3235) & (g3295) & (g3237) & (!g3238)) + ((!g1756) & (!g1792) & (!g3235) & (g3295) & (g3237) & (g3238)) + ((!g1756) & (!g1792) & (g3235) & (!g3295) & (!g3237) & (!g3238)) + ((!g1756) & (!g1792) & (g3235) & (!g3295) & (!g3237) & (g3238)) + ((!g1756) & (!g1792) & (g3235) & (!g3295) & (g3237) & (!g3238)) + ((!g1756) & (!g1792) & (g3235) & (!g3295) & (g3237) & (g3238)) + ((!g1756) & (!g1792) & (g3235) & (g3295) & (!g3237) & (!g3238)) + ((!g1756) & (g1792) & (!g3235) & (!g3295) & (!g3237) & (!g3238)) + ((!g1756) & (g1792) & (!g3235) & (!g3295) & (!g3237) & (g3238)) + ((!g1756) & (g1792) & (!g3235) & (!g3295) & (g3237) & (!g3238)) + ((!g1756) & (g1792) & (!g3235) & (!g3295) & (g3237) & (g3238)) + ((!g1756) & (g1792) & (g3235) & (!g3295) & (!g3237) & (!g3238)) + ((g1756) & (!g1792) & (!g3235) & (!g3295) & (!g3237) & (!g3238)) + ((g1756) & (!g1792) & (!g3235) & (!g3295) & (!g3237) & (g3238)) + ((g1756) & (!g1792) & (!g3235) & (!g3295) & (g3237) & (!g3238)) + ((g1756) & (!g1792) & (!g3235) & (!g3295) & (g3237) & (g3238)) + ((g1756) & (!g1792) & (!g3235) & (g3295) & (!g3237) & (!g3238)) + ((g1756) & (!g1792) & (g3235) & (!g3295) & (!g3237) & (!g3238)) + ((g1756) & (!g1792) & (g3235) & (!g3295) & (!g3237) & (g3238)) + ((g1756) & (!g1792) & (g3235) & (!g3295) & (g3237) & (!g3238)) + ((g1756) & (!g1792) & (g3235) & (!g3295) & (g3237) & (g3238)) + ((g1756) & (g1792) & (!g3235) & (!g3295) & (!g3237) & (!g3238)));
	assign g3332 = (((!g827) & (!g1825) & (g3330) & (!g3331)) + ((!g827) & (!g1825) & (g3330) & (g3331)) + ((!g827) & (g1825) & (g3330) & (!g3331)) + ((!g827) & (g1825) & (g3330) & (g3331)) + ((g827) & (!g1825) & (!g3330) & (!g3331)) + ((g827) & (!g1825) & (g3330) & (g3331)) + ((g827) & (g1825) & (!g3330) & (g3331)) + ((g827) & (g1825) & (g3330) & (!g3331)));
	assign g8256 = (((!g3499) & (g5501) & (!g3333)) + ((!g3499) & (g5501) & (g3333)) + ((g3499) & (!g5501) & (g3333)) + ((g3499) & (g5501) & (g3333)));
	assign g3334 = (((!g1758) & (!g1800) & (!g3240) & (!g3303) & (!g3242) & (!g3243)) + ((!g1758) & (!g1800) & (!g3240) & (!g3303) & (!g3242) & (g3243)) + ((!g1758) & (!g1800) & (!g3240) & (!g3303) & (g3242) & (!g3243)) + ((!g1758) & (!g1800) & (!g3240) & (!g3303) & (g3242) & (g3243)) + ((!g1758) & (!g1800) & (!g3240) & (g3303) & (!g3242) & (!g3243)) + ((!g1758) & (!g1800) & (!g3240) & (g3303) & (!g3242) & (g3243)) + ((!g1758) & (!g1800) & (!g3240) & (g3303) & (g3242) & (!g3243)) + ((!g1758) & (!g1800) & (!g3240) & (g3303) & (g3242) & (g3243)) + ((!g1758) & (!g1800) & (g3240) & (!g3303) & (!g3242) & (!g3243)) + ((!g1758) & (!g1800) & (g3240) & (!g3303) & (!g3242) & (g3243)) + ((!g1758) & (!g1800) & (g3240) & (!g3303) & (g3242) & (!g3243)) + ((!g1758) & (!g1800) & (g3240) & (!g3303) & (g3242) & (g3243)) + ((!g1758) & (!g1800) & (g3240) & (g3303) & (!g3242) & (!g3243)) + ((!g1758) & (g1800) & (!g3240) & (!g3303) & (!g3242) & (!g3243)) + ((!g1758) & (g1800) & (!g3240) & (!g3303) & (!g3242) & (g3243)) + ((!g1758) & (g1800) & (!g3240) & (!g3303) & (g3242) & (!g3243)) + ((!g1758) & (g1800) & (!g3240) & (!g3303) & (g3242) & (g3243)) + ((!g1758) & (g1800) & (g3240) & (!g3303) & (!g3242) & (!g3243)) + ((g1758) & (!g1800) & (!g3240) & (!g3303) & (!g3242) & (!g3243)) + ((g1758) & (!g1800) & (!g3240) & (!g3303) & (!g3242) & (g3243)) + ((g1758) & (!g1800) & (!g3240) & (!g3303) & (g3242) & (!g3243)) + ((g1758) & (!g1800) & (!g3240) & (!g3303) & (g3242) & (g3243)) + ((g1758) & (!g1800) & (!g3240) & (g3303) & (!g3242) & (!g3243)) + ((g1758) & (!g1800) & (g3240) & (!g3303) & (!g3242) & (!g3243)) + ((g1758) & (!g1800) & (g3240) & (!g3303) & (!g3242) & (g3243)) + ((g1758) & (!g1800) & (g3240) & (!g3303) & (g3242) & (!g3243)) + ((g1758) & (!g1800) & (g3240) & (!g3303) & (g3242) & (g3243)) + ((g1758) & (g1800) & (!g3240) & (!g3303) & (!g3242) & (!g3243)));
	assign g3335 = (((!g827) & (!g1827) & (g3333) & (!g3334)) + ((!g827) & (!g1827) & (g3333) & (g3334)) + ((!g827) & (g1827) & (g3333) & (!g3334)) + ((!g827) & (g1827) & (g3333) & (g3334)) + ((g827) & (!g1827) & (!g3333) & (!g3334)) + ((g827) & (!g1827) & (g3333) & (g3334)) + ((g827) & (g1827) & (!g3333) & (g3334)) + ((g827) & (g1827) & (g3333) & (!g3334)));
	assign g8257 = (((!g3464) & (g5504) & (!g3336)) + ((!g3464) & (g5504) & (g3336)) + ((g3464) & (!g5504) & (g3336)) + ((g3464) & (g5504) & (g3336)));
	assign g3337 = (((!g1760) & (!g1808) & (!g3245) & (!g3310) & (!g3247) & (!g3248)) + ((!g1760) & (!g1808) & (!g3245) & (!g3310) & (!g3247) & (g3248)) + ((!g1760) & (!g1808) & (!g3245) & (!g3310) & (g3247) & (!g3248)) + ((!g1760) & (!g1808) & (!g3245) & (!g3310) & (g3247) & (g3248)) + ((!g1760) & (!g1808) & (!g3245) & (g3310) & (!g3247) & (!g3248)) + ((!g1760) & (!g1808) & (!g3245) & (g3310) & (!g3247) & (g3248)) + ((!g1760) & (!g1808) & (!g3245) & (g3310) & (g3247) & (!g3248)) + ((!g1760) & (!g1808) & (!g3245) & (g3310) & (g3247) & (g3248)) + ((!g1760) & (!g1808) & (g3245) & (!g3310) & (!g3247) & (!g3248)) + ((!g1760) & (!g1808) & (g3245) & (!g3310) & (!g3247) & (g3248)) + ((!g1760) & (!g1808) & (g3245) & (!g3310) & (g3247) & (!g3248)) + ((!g1760) & (!g1808) & (g3245) & (!g3310) & (g3247) & (g3248)) + ((!g1760) & (!g1808) & (g3245) & (g3310) & (!g3247) & (!g3248)) + ((!g1760) & (g1808) & (!g3245) & (!g3310) & (!g3247) & (!g3248)) + ((!g1760) & (g1808) & (!g3245) & (!g3310) & (!g3247) & (g3248)) + ((!g1760) & (g1808) & (!g3245) & (!g3310) & (g3247) & (!g3248)) + ((!g1760) & (g1808) & (!g3245) & (!g3310) & (g3247) & (g3248)) + ((!g1760) & (g1808) & (g3245) & (!g3310) & (!g3247) & (!g3248)) + ((g1760) & (!g1808) & (!g3245) & (!g3310) & (!g3247) & (!g3248)) + ((g1760) & (!g1808) & (!g3245) & (!g3310) & (!g3247) & (g3248)) + ((g1760) & (!g1808) & (!g3245) & (!g3310) & (g3247) & (!g3248)) + ((g1760) & (!g1808) & (!g3245) & (!g3310) & (g3247) & (g3248)) + ((g1760) & (!g1808) & (!g3245) & (g3310) & (!g3247) & (!g3248)) + ((g1760) & (!g1808) & (g3245) & (!g3310) & (!g3247) & (!g3248)) + ((g1760) & (!g1808) & (g3245) & (!g3310) & (!g3247) & (g3248)) + ((g1760) & (!g1808) & (g3245) & (!g3310) & (g3247) & (!g3248)) + ((g1760) & (!g1808) & (g3245) & (!g3310) & (g3247) & (g3248)) + ((g1760) & (g1808) & (!g3245) & (!g3310) & (!g3247) & (!g3248)));
	assign g3338 = (((!g827) & (!g1829) & (g3336) & (!g3337)) + ((!g827) & (!g1829) & (g3336) & (g3337)) + ((!g827) & (g1829) & (g3336) & (!g3337)) + ((!g827) & (g1829) & (g3336) & (g3337)) + ((g827) & (!g1829) & (!g3336) & (!g3337)) + ((g827) & (!g1829) & (g3336) & (g3337)) + ((g827) & (g1829) & (!g3336) & (g3337)) + ((g827) & (g1829) & (g3336) & (!g3337)));
	assign g8258 = (((!g3499) & (g5507) & (!g3339)) + ((!g3499) & (g5507) & (g3339)) + ((g3499) & (!g5507) & (g3339)) + ((g3499) & (g5507) & (g3339)));
	assign g3340 = (((!g1762) & (!g1786) & (!g3250) & (!g3291) & (!g3252) & (!g3253)) + ((!g1762) & (!g1786) & (!g3250) & (!g3291) & (!g3252) & (g3253)) + ((!g1762) & (!g1786) & (!g3250) & (!g3291) & (g3252) & (!g3253)) + ((!g1762) & (!g1786) & (!g3250) & (!g3291) & (g3252) & (g3253)) + ((!g1762) & (!g1786) & (!g3250) & (g3291) & (!g3252) & (!g3253)) + ((!g1762) & (!g1786) & (!g3250) & (g3291) & (!g3252) & (g3253)) + ((!g1762) & (!g1786) & (!g3250) & (g3291) & (g3252) & (!g3253)) + ((!g1762) & (!g1786) & (!g3250) & (g3291) & (g3252) & (g3253)) + ((!g1762) & (!g1786) & (g3250) & (!g3291) & (!g3252) & (!g3253)) + ((!g1762) & (!g1786) & (g3250) & (!g3291) & (!g3252) & (g3253)) + ((!g1762) & (!g1786) & (g3250) & (!g3291) & (g3252) & (!g3253)) + ((!g1762) & (!g1786) & (g3250) & (!g3291) & (g3252) & (g3253)) + ((!g1762) & (!g1786) & (g3250) & (g3291) & (!g3252) & (!g3253)) + ((!g1762) & (g1786) & (!g3250) & (!g3291) & (!g3252) & (!g3253)) + ((!g1762) & (g1786) & (!g3250) & (!g3291) & (!g3252) & (g3253)) + ((!g1762) & (g1786) & (!g3250) & (!g3291) & (g3252) & (!g3253)) + ((!g1762) & (g1786) & (!g3250) & (!g3291) & (g3252) & (g3253)) + ((!g1762) & (g1786) & (g3250) & (!g3291) & (!g3252) & (!g3253)) + ((g1762) & (!g1786) & (!g3250) & (!g3291) & (!g3252) & (!g3253)) + ((g1762) & (!g1786) & (!g3250) & (!g3291) & (!g3252) & (g3253)) + ((g1762) & (!g1786) & (!g3250) & (!g3291) & (g3252) & (!g3253)) + ((g1762) & (!g1786) & (!g3250) & (!g3291) & (g3252) & (g3253)) + ((g1762) & (!g1786) & (!g3250) & (g3291) & (!g3252) & (!g3253)) + ((g1762) & (!g1786) & (g3250) & (!g3291) & (!g3252) & (!g3253)) + ((g1762) & (!g1786) & (g3250) & (!g3291) & (!g3252) & (g3253)) + ((g1762) & (!g1786) & (g3250) & (!g3291) & (g3252) & (!g3253)) + ((g1762) & (!g1786) & (g3250) & (!g3291) & (g3252) & (g3253)) + ((g1762) & (g1786) & (!g3250) & (!g3291) & (!g3252) & (!g3253)));
	assign g3341 = (((!g827) & (!g1831) & (g3339) & (!g3340)) + ((!g827) & (!g1831) & (g3339) & (g3340)) + ((!g827) & (g1831) & (g3339) & (!g3340)) + ((!g827) & (g1831) & (g3339) & (g3340)) + ((g827) & (!g1831) & (!g3339) & (!g3340)) + ((g827) & (!g1831) & (g3339) & (g3340)) + ((g827) & (g1831) & (!g3339) & (g3340)) + ((g827) & (g1831) & (g3339) & (!g3340)));
	assign g8259 = (((!g3464) & (g5511) & (!g3342)) + ((!g3464) & (g5511) & (g3342)) + ((g3464) & (!g5511) & (g3342)) + ((g3464) & (g5511) & (g3342)));
	assign g3343 = (((!g1764) & (!g1794) & (!g3255) & (!g3297) & (!g3257) & (!g3258)) + ((!g1764) & (!g1794) & (!g3255) & (!g3297) & (!g3257) & (g3258)) + ((!g1764) & (!g1794) & (!g3255) & (!g3297) & (g3257) & (!g3258)) + ((!g1764) & (!g1794) & (!g3255) & (!g3297) & (g3257) & (g3258)) + ((!g1764) & (!g1794) & (!g3255) & (g3297) & (!g3257) & (!g3258)) + ((!g1764) & (!g1794) & (!g3255) & (g3297) & (!g3257) & (g3258)) + ((!g1764) & (!g1794) & (!g3255) & (g3297) & (g3257) & (!g3258)) + ((!g1764) & (!g1794) & (!g3255) & (g3297) & (g3257) & (g3258)) + ((!g1764) & (!g1794) & (g3255) & (!g3297) & (!g3257) & (!g3258)) + ((!g1764) & (!g1794) & (g3255) & (!g3297) & (!g3257) & (g3258)) + ((!g1764) & (!g1794) & (g3255) & (!g3297) & (g3257) & (!g3258)) + ((!g1764) & (!g1794) & (g3255) & (!g3297) & (g3257) & (g3258)) + ((!g1764) & (!g1794) & (g3255) & (g3297) & (!g3257) & (!g3258)) + ((!g1764) & (g1794) & (!g3255) & (!g3297) & (!g3257) & (!g3258)) + ((!g1764) & (g1794) & (!g3255) & (!g3297) & (!g3257) & (g3258)) + ((!g1764) & (g1794) & (!g3255) & (!g3297) & (g3257) & (!g3258)) + ((!g1764) & (g1794) & (!g3255) & (!g3297) & (g3257) & (g3258)) + ((!g1764) & (g1794) & (g3255) & (!g3297) & (!g3257) & (!g3258)) + ((g1764) & (!g1794) & (!g3255) & (!g3297) & (!g3257) & (!g3258)) + ((g1764) & (!g1794) & (!g3255) & (!g3297) & (!g3257) & (g3258)) + ((g1764) & (!g1794) & (!g3255) & (!g3297) & (g3257) & (!g3258)) + ((g1764) & (!g1794) & (!g3255) & (!g3297) & (g3257) & (g3258)) + ((g1764) & (!g1794) & (!g3255) & (g3297) & (!g3257) & (!g3258)) + ((g1764) & (!g1794) & (g3255) & (!g3297) & (!g3257) & (!g3258)) + ((g1764) & (!g1794) & (g3255) & (!g3297) & (!g3257) & (g3258)) + ((g1764) & (!g1794) & (g3255) & (!g3297) & (g3257) & (!g3258)) + ((g1764) & (!g1794) & (g3255) & (!g3297) & (g3257) & (g3258)) + ((g1764) & (g1794) & (!g3255) & (!g3297) & (!g3257) & (!g3258)));
	assign g3344 = (((!g827) & (!g1833) & (g3342) & (!g3343)) + ((!g827) & (!g1833) & (g3342) & (g3343)) + ((!g827) & (g1833) & (g3342) & (!g3343)) + ((!g827) & (g1833) & (g3342) & (g3343)) + ((g827) & (!g1833) & (!g3342) & (!g3343)) + ((g827) & (!g1833) & (g3342) & (g3343)) + ((g827) & (g1833) & (!g3342) & (g3343)) + ((g827) & (g1833) & (g3342) & (!g3343)));
	assign g8260 = (((!g2017) & (g5514) & (!g3345)) + ((!g2017) & (g5514) & (g3345)) + ((g2017) & (!g5514) & (g3345)) + ((g2017) & (g5514) & (g3345)));
	assign g3346 = (((!g1766) & (!g1802) & (!g3260) & (!g3305) & (!g3262) & (!g3263)) + ((!g1766) & (!g1802) & (!g3260) & (!g3305) & (!g3262) & (g3263)) + ((!g1766) & (!g1802) & (!g3260) & (!g3305) & (g3262) & (!g3263)) + ((!g1766) & (!g1802) & (!g3260) & (!g3305) & (g3262) & (g3263)) + ((!g1766) & (!g1802) & (!g3260) & (g3305) & (!g3262) & (!g3263)) + ((!g1766) & (!g1802) & (!g3260) & (g3305) & (!g3262) & (g3263)) + ((!g1766) & (!g1802) & (!g3260) & (g3305) & (g3262) & (!g3263)) + ((!g1766) & (!g1802) & (!g3260) & (g3305) & (g3262) & (g3263)) + ((!g1766) & (!g1802) & (g3260) & (!g3305) & (!g3262) & (!g3263)) + ((!g1766) & (!g1802) & (g3260) & (!g3305) & (!g3262) & (g3263)) + ((!g1766) & (!g1802) & (g3260) & (!g3305) & (g3262) & (!g3263)) + ((!g1766) & (!g1802) & (g3260) & (!g3305) & (g3262) & (g3263)) + ((!g1766) & (!g1802) & (g3260) & (g3305) & (!g3262) & (!g3263)) + ((!g1766) & (g1802) & (!g3260) & (!g3305) & (!g3262) & (!g3263)) + ((!g1766) & (g1802) & (!g3260) & (!g3305) & (!g3262) & (g3263)) + ((!g1766) & (g1802) & (!g3260) & (!g3305) & (g3262) & (!g3263)) + ((!g1766) & (g1802) & (!g3260) & (!g3305) & (g3262) & (g3263)) + ((!g1766) & (g1802) & (g3260) & (!g3305) & (!g3262) & (!g3263)) + ((g1766) & (!g1802) & (!g3260) & (!g3305) & (!g3262) & (!g3263)) + ((g1766) & (!g1802) & (!g3260) & (!g3305) & (!g3262) & (g3263)) + ((g1766) & (!g1802) & (!g3260) & (!g3305) & (g3262) & (!g3263)) + ((g1766) & (!g1802) & (!g3260) & (!g3305) & (g3262) & (g3263)) + ((g1766) & (!g1802) & (!g3260) & (g3305) & (!g3262) & (!g3263)) + ((g1766) & (!g1802) & (g3260) & (!g3305) & (!g3262) & (!g3263)) + ((g1766) & (!g1802) & (g3260) & (!g3305) & (!g3262) & (g3263)) + ((g1766) & (!g1802) & (g3260) & (!g3305) & (g3262) & (!g3263)) + ((g1766) & (!g1802) & (g3260) & (!g3305) & (g3262) & (g3263)) + ((g1766) & (g1802) & (!g3260) & (!g3305) & (!g3262) & (!g3263)));
	assign g3347 = (((!g827) & (!g1835) & (g3345) & (!g3346)) + ((!g827) & (!g1835) & (g3345) & (g3346)) + ((!g827) & (g1835) & (g3345) & (!g3346)) + ((!g827) & (g1835) & (g3345) & (g3346)) + ((g827) & (!g1835) & (!g3345) & (!g3346)) + ((g827) & (!g1835) & (g3345) & (g3346)) + ((g827) & (g1835) & (!g3345) & (g3346)) + ((g827) & (g1835) & (g3345) & (!g3346)));
	assign g8261 = (((!g3429) & (g5517) & (!g3348)) + ((!g3429) & (g5517) & (g3348)) + ((g3429) & (!g5517) & (g3348)) + ((g3429) & (g5517) & (g3348)));
	assign g3349 = (((!g1768) & (!g1810) & (!g3265) & (!g3312) & (!g3267) & (!g3268)) + ((!g1768) & (!g1810) & (!g3265) & (!g3312) & (!g3267) & (g3268)) + ((!g1768) & (!g1810) & (!g3265) & (!g3312) & (g3267) & (!g3268)) + ((!g1768) & (!g1810) & (!g3265) & (!g3312) & (g3267) & (g3268)) + ((!g1768) & (!g1810) & (!g3265) & (g3312) & (!g3267) & (!g3268)) + ((!g1768) & (!g1810) & (!g3265) & (g3312) & (!g3267) & (g3268)) + ((!g1768) & (!g1810) & (!g3265) & (g3312) & (g3267) & (!g3268)) + ((!g1768) & (!g1810) & (!g3265) & (g3312) & (g3267) & (g3268)) + ((!g1768) & (!g1810) & (g3265) & (!g3312) & (!g3267) & (!g3268)) + ((!g1768) & (!g1810) & (g3265) & (!g3312) & (!g3267) & (g3268)) + ((!g1768) & (!g1810) & (g3265) & (!g3312) & (g3267) & (!g3268)) + ((!g1768) & (!g1810) & (g3265) & (!g3312) & (g3267) & (g3268)) + ((!g1768) & (!g1810) & (g3265) & (g3312) & (!g3267) & (!g3268)) + ((!g1768) & (g1810) & (!g3265) & (!g3312) & (!g3267) & (!g3268)) + ((!g1768) & (g1810) & (!g3265) & (!g3312) & (!g3267) & (g3268)) + ((!g1768) & (g1810) & (!g3265) & (!g3312) & (g3267) & (!g3268)) + ((!g1768) & (g1810) & (!g3265) & (!g3312) & (g3267) & (g3268)) + ((!g1768) & (g1810) & (g3265) & (!g3312) & (!g3267) & (!g3268)) + ((g1768) & (!g1810) & (!g3265) & (!g3312) & (!g3267) & (!g3268)) + ((g1768) & (!g1810) & (!g3265) & (!g3312) & (!g3267) & (g3268)) + ((g1768) & (!g1810) & (!g3265) & (!g3312) & (g3267) & (!g3268)) + ((g1768) & (!g1810) & (!g3265) & (!g3312) & (g3267) & (g3268)) + ((g1768) & (!g1810) & (!g3265) & (g3312) & (!g3267) & (!g3268)) + ((g1768) & (!g1810) & (g3265) & (!g3312) & (!g3267) & (!g3268)) + ((g1768) & (!g1810) & (g3265) & (!g3312) & (!g3267) & (g3268)) + ((g1768) & (!g1810) & (g3265) & (!g3312) & (g3267) & (!g3268)) + ((g1768) & (!g1810) & (g3265) & (!g3312) & (g3267) & (g3268)) + ((g1768) & (g1810) & (!g3265) & (!g3312) & (!g3267) & (!g3268)));
	assign g3350 = (((!g827) & (!g1837) & (g3348) & (!g3349)) + ((!g827) & (!g1837) & (g3348) & (g3349)) + ((!g827) & (g1837) & (g3348) & (!g3349)) + ((!g827) & (g1837) & (g3348) & (g3349)) + ((g827) & (!g1837) & (!g3348) & (!g3349)) + ((g827) & (!g1837) & (g3348) & (g3349)) + ((g827) & (g1837) & (!g3348) & (g3349)) + ((g827) & (g1837) & (g3348) & (!g3349)));
	assign g3351 = (((!g1770) & (!g1788) & (!g2648) & (!g2679) & (!g3271) & (!g3272)) + ((!g1770) & (!g1788) & (!g2648) & (!g2679) & (!g3271) & (g3272)) + ((!g1770) & (!g1788) & (!g2648) & (!g2679) & (g3271) & (!g3272)) + ((!g1770) & (!g1788) & (!g2648) & (!g2679) & (g3271) & (g3272)) + ((!g1770) & (!g1788) & (!g2648) & (g2679) & (!g3271) & (!g3272)) + ((!g1770) & (!g1788) & (!g2648) & (g2679) & (!g3271) & (g3272)) + ((!g1770) & (!g1788) & (!g2648) & (g2679) & (g3271) & (!g3272)) + ((!g1770) & (!g1788) & (!g2648) & (g2679) & (g3271) & (g3272)) + ((!g1770) & (!g1788) & (g2648) & (!g2679) & (!g3271) & (!g3272)) + ((!g1770) & (!g1788) & (g2648) & (!g2679) & (!g3271) & (g3272)) + ((!g1770) & (!g1788) & (g2648) & (!g2679) & (g3271) & (!g3272)) + ((!g1770) & (!g1788) & (g2648) & (!g2679) & (g3271) & (g3272)) + ((!g1770) & (!g1788) & (g2648) & (g2679) & (!g3271) & (!g3272)) + ((!g1770) & (g1788) & (!g2648) & (!g2679) & (!g3271) & (!g3272)) + ((!g1770) & (g1788) & (!g2648) & (!g2679) & (!g3271) & (g3272)) + ((!g1770) & (g1788) & (!g2648) & (!g2679) & (g3271) & (!g3272)) + ((!g1770) & (g1788) & (!g2648) & (!g2679) & (g3271) & (g3272)) + ((!g1770) & (g1788) & (g2648) & (!g2679) & (!g3271) & (!g3272)) + ((g1770) & (!g1788) & (!g2648) & (!g2679) & (!g3271) & (!g3272)) + ((g1770) & (!g1788) & (!g2648) & (!g2679) & (!g3271) & (g3272)) + ((g1770) & (!g1788) & (!g2648) & (!g2679) & (g3271) & (!g3272)) + ((g1770) & (!g1788) & (!g2648) & (!g2679) & (g3271) & (g3272)) + ((g1770) & (!g1788) & (!g2648) & (g2679) & (!g3271) & (!g3272)) + ((g1770) & (!g1788) & (g2648) & (!g2679) & (!g3271) & (!g3272)) + ((g1770) & (!g1788) & (g2648) & (!g2679) & (!g3271) & (g3272)) + ((g1770) & (!g1788) & (g2648) & (!g2679) & (g3271) & (!g3272)) + ((g1770) & (!g1788) & (g2648) & (!g2679) & (g3271) & (g3272)) + ((g1770) & (g1788) & (!g2648) & (!g2679) & (!g3271) & (!g3272)));
	assign g3352 = (((!g827) & (!g1839) & (g2759) & (!g3351)) + ((!g827) & (!g1839) & (g2759) & (g3351)) + ((!g827) & (g1839) & (g2759) & (!g3351)) + ((!g827) & (g1839) & (g2759) & (g3351)) + ((g827) & (!g1839) & (!g2759) & (!g3351)) + ((g827) & (!g1839) & (g2759) & (g3351)) + ((g827) & (g1839) & (!g2759) & (g3351)) + ((g827) & (g1839) & (g2759) & (!g3351)));
	assign g8262 = (((!g3499) & (g5520) & (!g3353)) + ((!g3499) & (g5520) & (g3353)) + ((g3499) & (!g5520) & (g3353)) + ((g3499) & (g5520) & (g3353)));
	assign g3354 = (((!g1772) & (!g1796) & (!g3274) & (!g3299) & (!g3276) & (!g3277)) + ((!g1772) & (!g1796) & (!g3274) & (!g3299) & (!g3276) & (g3277)) + ((!g1772) & (!g1796) & (!g3274) & (!g3299) & (g3276) & (!g3277)) + ((!g1772) & (!g1796) & (!g3274) & (!g3299) & (g3276) & (g3277)) + ((!g1772) & (!g1796) & (!g3274) & (g3299) & (!g3276) & (!g3277)) + ((!g1772) & (!g1796) & (!g3274) & (g3299) & (!g3276) & (g3277)) + ((!g1772) & (!g1796) & (!g3274) & (g3299) & (g3276) & (!g3277)) + ((!g1772) & (!g1796) & (!g3274) & (g3299) & (g3276) & (g3277)) + ((!g1772) & (!g1796) & (g3274) & (!g3299) & (!g3276) & (!g3277)) + ((!g1772) & (!g1796) & (g3274) & (!g3299) & (!g3276) & (g3277)) + ((!g1772) & (!g1796) & (g3274) & (!g3299) & (g3276) & (!g3277)) + ((!g1772) & (!g1796) & (g3274) & (!g3299) & (g3276) & (g3277)) + ((!g1772) & (!g1796) & (g3274) & (g3299) & (!g3276) & (!g3277)) + ((!g1772) & (g1796) & (!g3274) & (!g3299) & (!g3276) & (!g3277)) + ((!g1772) & (g1796) & (!g3274) & (!g3299) & (!g3276) & (g3277)) + ((!g1772) & (g1796) & (!g3274) & (!g3299) & (g3276) & (!g3277)) + ((!g1772) & (g1796) & (!g3274) & (!g3299) & (g3276) & (g3277)) + ((!g1772) & (g1796) & (g3274) & (!g3299) & (!g3276) & (!g3277)) + ((g1772) & (!g1796) & (!g3274) & (!g3299) & (!g3276) & (!g3277)) + ((g1772) & (!g1796) & (!g3274) & (!g3299) & (!g3276) & (g3277)) + ((g1772) & (!g1796) & (!g3274) & (!g3299) & (g3276) & (!g3277)) + ((g1772) & (!g1796) & (!g3274) & (!g3299) & (g3276) & (g3277)) + ((g1772) & (!g1796) & (!g3274) & (g3299) & (!g3276) & (!g3277)) + ((g1772) & (!g1796) & (g3274) & (!g3299) & (!g3276) & (!g3277)) + ((g1772) & (!g1796) & (g3274) & (!g3299) & (!g3276) & (g3277)) + ((g1772) & (!g1796) & (g3274) & (!g3299) & (g3276) & (!g3277)) + ((g1772) & (!g1796) & (g3274) & (!g3299) & (g3276) & (g3277)) + ((g1772) & (g1796) & (!g3274) & (!g3299) & (!g3276) & (!g3277)));
	assign g3355 = (((!g827) & (!g1841) & (g3353) & (!g3354)) + ((!g827) & (!g1841) & (g3353) & (g3354)) + ((!g827) & (g1841) & (g3353) & (!g3354)) + ((!g827) & (g1841) & (g3353) & (g3354)) + ((g827) & (!g1841) & (!g3353) & (!g3354)) + ((g827) & (!g1841) & (g3353) & (g3354)) + ((g827) & (g1841) & (!g3353) & (g3354)) + ((g827) & (g1841) & (g3353) & (!g3354)));
	assign g8263 = (((!g3429) & (g5523) & (!g3356)) + ((!g3429) & (g5523) & (g3356)) + ((g3429) & (!g5523) & (g3356)) + ((g3429) & (g5523) & (g3356)));
	assign g3357 = (((!g1774) & (!g1804) & (!g3279) & (!g3307) & (!g3281) & (!g3282)) + ((!g1774) & (!g1804) & (!g3279) & (!g3307) & (!g3281) & (g3282)) + ((!g1774) & (!g1804) & (!g3279) & (!g3307) & (g3281) & (!g3282)) + ((!g1774) & (!g1804) & (!g3279) & (!g3307) & (g3281) & (g3282)) + ((!g1774) & (!g1804) & (!g3279) & (g3307) & (!g3281) & (!g3282)) + ((!g1774) & (!g1804) & (!g3279) & (g3307) & (!g3281) & (g3282)) + ((!g1774) & (!g1804) & (!g3279) & (g3307) & (g3281) & (!g3282)) + ((!g1774) & (!g1804) & (!g3279) & (g3307) & (g3281) & (g3282)) + ((!g1774) & (!g1804) & (g3279) & (!g3307) & (!g3281) & (!g3282)) + ((!g1774) & (!g1804) & (g3279) & (!g3307) & (!g3281) & (g3282)) + ((!g1774) & (!g1804) & (g3279) & (!g3307) & (g3281) & (!g3282)) + ((!g1774) & (!g1804) & (g3279) & (!g3307) & (g3281) & (g3282)) + ((!g1774) & (!g1804) & (g3279) & (g3307) & (!g3281) & (!g3282)) + ((!g1774) & (g1804) & (!g3279) & (!g3307) & (!g3281) & (!g3282)) + ((!g1774) & (g1804) & (!g3279) & (!g3307) & (!g3281) & (g3282)) + ((!g1774) & (g1804) & (!g3279) & (!g3307) & (g3281) & (!g3282)) + ((!g1774) & (g1804) & (!g3279) & (!g3307) & (g3281) & (g3282)) + ((!g1774) & (g1804) & (g3279) & (!g3307) & (!g3281) & (!g3282)) + ((g1774) & (!g1804) & (!g3279) & (!g3307) & (!g3281) & (!g3282)) + ((g1774) & (!g1804) & (!g3279) & (!g3307) & (!g3281) & (g3282)) + ((g1774) & (!g1804) & (!g3279) & (!g3307) & (g3281) & (!g3282)) + ((g1774) & (!g1804) & (!g3279) & (!g3307) & (g3281) & (g3282)) + ((g1774) & (!g1804) & (!g3279) & (g3307) & (!g3281) & (!g3282)) + ((g1774) & (!g1804) & (g3279) & (!g3307) & (!g3281) & (!g3282)) + ((g1774) & (!g1804) & (g3279) & (!g3307) & (!g3281) & (g3282)) + ((g1774) & (!g1804) & (g3279) & (!g3307) & (g3281) & (!g3282)) + ((g1774) & (!g1804) & (g3279) & (!g3307) & (g3281) & (g3282)) + ((g1774) & (g1804) & (!g3279) & (!g3307) & (!g3281) & (!g3282)));
	assign g3358 = (((!g827) & (!g1843) & (g3356) & (!g3357)) + ((!g827) & (!g1843) & (g3356) & (g3357)) + ((!g827) & (g1843) & (g3356) & (!g3357)) + ((!g827) & (g1843) & (g3356) & (g3357)) + ((g827) & (!g1843) & (!g3356) & (!g3357)) + ((g827) & (!g1843) & (g3356) & (g3357)) + ((g827) & (g1843) & (!g3356) & (g3357)) + ((g827) & (g1843) & (g3356) & (!g3357)));
	assign g8264 = (((!g2017) & (g5526) & (!g3359)) + ((!g2017) & (g5526) & (g3359)) + ((g2017) & (!g5526) & (g3359)) + ((g2017) & (g5526) & (g3359)));
	assign g3360 = (((!g1776) & (!g1812) & (!g3284) & (!g3314) & (!g3286) & (!g3287)) + ((!g1776) & (!g1812) & (!g3284) & (!g3314) & (!g3286) & (g3287)) + ((!g1776) & (!g1812) & (!g3284) & (!g3314) & (g3286) & (!g3287)) + ((!g1776) & (!g1812) & (!g3284) & (!g3314) & (g3286) & (g3287)) + ((!g1776) & (!g1812) & (!g3284) & (g3314) & (!g3286) & (!g3287)) + ((!g1776) & (!g1812) & (!g3284) & (g3314) & (!g3286) & (g3287)) + ((!g1776) & (!g1812) & (!g3284) & (g3314) & (g3286) & (!g3287)) + ((!g1776) & (!g1812) & (!g3284) & (g3314) & (g3286) & (g3287)) + ((!g1776) & (!g1812) & (g3284) & (!g3314) & (!g3286) & (!g3287)) + ((!g1776) & (!g1812) & (g3284) & (!g3314) & (!g3286) & (g3287)) + ((!g1776) & (!g1812) & (g3284) & (!g3314) & (g3286) & (!g3287)) + ((!g1776) & (!g1812) & (g3284) & (!g3314) & (g3286) & (g3287)) + ((!g1776) & (!g1812) & (g3284) & (g3314) & (!g3286) & (!g3287)) + ((!g1776) & (g1812) & (!g3284) & (!g3314) & (!g3286) & (!g3287)) + ((!g1776) & (g1812) & (!g3284) & (!g3314) & (!g3286) & (g3287)) + ((!g1776) & (g1812) & (!g3284) & (!g3314) & (g3286) & (!g3287)) + ((!g1776) & (g1812) & (!g3284) & (!g3314) & (g3286) & (g3287)) + ((!g1776) & (g1812) & (g3284) & (!g3314) & (!g3286) & (!g3287)) + ((g1776) & (!g1812) & (!g3284) & (!g3314) & (!g3286) & (!g3287)) + ((g1776) & (!g1812) & (!g3284) & (!g3314) & (!g3286) & (g3287)) + ((g1776) & (!g1812) & (!g3284) & (!g3314) & (g3286) & (!g3287)) + ((g1776) & (!g1812) & (!g3284) & (!g3314) & (g3286) & (g3287)) + ((g1776) & (!g1812) & (!g3284) & (g3314) & (!g3286) & (!g3287)) + ((g1776) & (!g1812) & (g3284) & (!g3314) & (!g3286) & (!g3287)) + ((g1776) & (!g1812) & (g3284) & (!g3314) & (!g3286) & (g3287)) + ((g1776) & (!g1812) & (g3284) & (!g3314) & (g3286) & (!g3287)) + ((g1776) & (!g1812) & (g3284) & (!g3314) & (g3286) & (g3287)) + ((g1776) & (g1812) & (!g3284) & (!g3314) & (!g3286) & (!g3287)));
	assign g3361 = (((!g827) & (!g1845) & (g3359) & (!g3360)) + ((!g827) & (!g1845) & (g3359) & (g3360)) + ((!g827) & (g1845) & (g3359) & (!g3360)) + ((!g827) & (g1845) & (g3359) & (g3360)) + ((g827) & (!g1845) & (!g3359) & (!g3360)) + ((g827) & (!g1845) & (g3359) & (g3360)) + ((g827) & (g1845) & (!g3359) & (g3360)) + ((g827) & (g1845) & (g3359) & (!g3360)));
	assign g3362 = (((!g3316) & (!g1967) & (!g1968) & (!g1969) & (g1970)) + ((!g3316) & (!g1967) & (!g1968) & (g1969) & (!g1970)) + ((!g3316) & (!g1967) & (g1968) & (!g1969) & (!g1970)) + ((!g3316) & (!g1967) & (g1968) & (g1969) & (g1970)) + ((!g3316) & (g1967) & (!g1968) & (!g1969) & (!g1970)) + ((!g3316) & (g1967) & (!g1968) & (g1969) & (g1970)) + ((!g3316) & (g1967) & (g1968) & (!g1969) & (!g1970)) + ((!g3316) & (g1967) & (g1968) & (g1969) & (g1970)) + ((g3316) & (!g1967) & (!g1968) & (!g1969) & (g1970)) + ((g3316) & (!g1967) & (!g1968) & (g1969) & (!g1970)) + ((g3316) & (!g1967) & (g1968) & (!g1969) & (g1970)) + ((g3316) & (!g1967) & (g1968) & (g1969) & (!g1970)) + ((g3316) & (g1967) & (!g1968) & (!g1969) & (g1970)) + ((g3316) & (g1967) & (!g1968) & (g1969) & (!g1970)) + ((g3316) & (g1967) & (g1968) & (!g1969) & (!g1970)) + ((g3316) & (g1967) & (g1968) & (g1969) & (g1970)));
	assign g3363 = (((!g3318) & (!g2003) & (!g2004) & (!g2005) & (g2006)) + ((!g3318) & (!g2003) & (!g2004) & (g2005) & (!g2006)) + ((!g3318) & (!g2003) & (g2004) & (!g2005) & (g2006)) + ((!g3318) & (!g2003) & (g2004) & (g2005) & (!g2006)) + ((!g3318) & (g2003) & (!g2004) & (!g2005) & (g2006)) + ((!g3318) & (g2003) & (!g2004) & (g2005) & (!g2006)) + ((!g3318) & (g2003) & (g2004) & (!g2005) & (!g2006)) + ((!g3318) & (g2003) & (g2004) & (g2005) & (g2006)) + ((g3318) & (!g2003) & (!g2004) & (!g2005) & (g2006)) + ((g3318) & (!g2003) & (!g2004) & (g2005) & (!g2006)) + ((g3318) & (!g2003) & (g2004) & (!g2005) & (!g2006)) + ((g3318) & (!g2003) & (g2004) & (g2005) & (g2006)) + ((g3318) & (g2003) & (!g2004) & (!g2005) & (!g2006)) + ((g3318) & (g2003) & (!g2004) & (g2005) & (g2006)) + ((g3318) & (g2003) & (g2004) & (!g2005) & (!g2006)) + ((g3318) & (g2003) & (g2004) & (g2005) & (g2006)));
	assign g3364 = (((!g830) & (!g1914) & (!g3362) & (!g3363) & (!g1847)) + ((!g830) & (!g1914) & (!g3362) & (!g3363) & (g1847)) + ((!g830) & (!g1914) & (!g3362) & (g3363) & (!g1847)) + ((!g830) & (!g1914) & (!g3362) & (g3363) & (g1847)) + ((!g830) & (!g1914) & (g3362) & (!g3363) & (!g1847)) + ((!g830) & (!g1914) & (g3362) & (!g3363) & (g1847)) + ((!g830) & (!g1914) & (g3362) & (g3363) & (!g1847)) + ((!g830) & (!g1914) & (g3362) & (g3363) & (g1847)) + ((!g830) & (g1914) & (!g3362) & (!g3363) & (!g1847)) + ((!g830) & (g1914) & (!g3362) & (!g3363) & (g1847)) + ((!g830) & (g1914) & (!g3362) & (g3363) & (!g1847)) + ((!g830) & (g1914) & (!g3362) & (g3363) & (g1847)) + ((!g830) & (g1914) & (g3362) & (!g3363) & (!g1847)) + ((!g830) & (g1914) & (g3362) & (!g3363) & (g1847)) + ((!g830) & (g1914) & (g3362) & (g3363) & (!g1847)) + ((!g830) & (g1914) & (g3362) & (g3363) & (g1847)) + ((g830) & (!g1914) & (!g3362) & (!g3363) & (g1847)) + ((g830) & (!g1914) & (!g3362) & (g3363) & (!g1847)) + ((g830) & (!g1914) & (g3362) & (!g3363) & (g1847)) + ((g830) & (!g1914) & (g3362) & (g3363) & (!g1847)) + ((g830) & (g1914) & (!g3362) & (!g3363) & (g1847)) + ((g830) & (g1914) & (!g3362) & (g3363) & (g1847)) + ((g830) & (g1914) & (g3362) & (!g3363) & (!g1847)) + ((g830) & (g1914) & (g3362) & (g3363) & (!g1847)));
	assign g3365 = (((!g827) & (!g1823) & (!g1851) & (!g2758) & (g2789) & (!g3328)) + ((!g827) & (!g1823) & (!g1851) & (!g2758) & (g2789) & (g3328)) + ((!g827) & (!g1823) & (!g1851) & (g2758) & (g2789) & (!g3328)) + ((!g827) & (!g1823) & (!g1851) & (g2758) & (g2789) & (g3328)) + ((!g827) & (!g1823) & (g1851) & (!g2758) & (g2789) & (!g3328)) + ((!g827) & (!g1823) & (g1851) & (!g2758) & (g2789) & (g3328)) + ((!g827) & (!g1823) & (g1851) & (g2758) & (g2789) & (!g3328)) + ((!g827) & (!g1823) & (g1851) & (g2758) & (g2789) & (g3328)) + ((!g827) & (g1823) & (!g1851) & (!g2758) & (g2789) & (!g3328)) + ((!g827) & (g1823) & (!g1851) & (!g2758) & (g2789) & (g3328)) + ((!g827) & (g1823) & (!g1851) & (g2758) & (g2789) & (!g3328)) + ((!g827) & (g1823) & (!g1851) & (g2758) & (g2789) & (g3328)) + ((!g827) & (g1823) & (g1851) & (!g2758) & (g2789) & (!g3328)) + ((!g827) & (g1823) & (g1851) & (!g2758) & (g2789) & (g3328)) + ((!g827) & (g1823) & (g1851) & (g2758) & (g2789) & (!g3328)) + ((!g827) & (g1823) & (g1851) & (g2758) & (g2789) & (g3328)) + ((g827) & (!g1823) & (!g1851) & (!g2758) & (g2789) & (!g3328)) + ((g827) & (!g1823) & (!g1851) & (!g2758) & (g2789) & (g3328)) + ((g827) & (!g1823) & (!g1851) & (g2758) & (!g2789) & (!g3328)) + ((g827) & (!g1823) & (!g1851) & (g2758) & (g2789) & (g3328)) + ((g827) & (!g1823) & (g1851) & (!g2758) & (!g2789) & (!g3328)) + ((g827) & (!g1823) & (g1851) & (!g2758) & (!g2789) & (g3328)) + ((g827) & (!g1823) & (g1851) & (g2758) & (!g2789) & (g3328)) + ((g827) & (!g1823) & (g1851) & (g2758) & (g2789) & (!g3328)) + ((g827) & (g1823) & (!g1851) & (!g2758) & (!g2789) & (!g3328)) + ((g827) & (g1823) & (!g1851) & (!g2758) & (g2789) & (g3328)) + ((g827) & (g1823) & (!g1851) & (g2758) & (!g2789) & (!g3328)) + ((g827) & (g1823) & (!g1851) & (g2758) & (!g2789) & (g3328)) + ((g827) & (g1823) & (g1851) & (!g2758) & (!g2789) & (g3328)) + ((g827) & (g1823) & (g1851) & (!g2758) & (g2789) & (!g3328)) + ((g827) & (g1823) & (g1851) & (g2758) & (g2789) & (!g3328)) + ((g827) & (g1823) & (g1851) & (g2758) & (g2789) & (g3328)));
	assign g8265 = (((!g3499) & (g5529) & (!g3366)) + ((!g3499) & (g5529) & (g3366)) + ((g3499) & (!g5529) & (g3366)) + ((g3499) & (g5529) & (g3366)));
	assign g3367 = (((!g827) & (!g1831) & (!g1853) & (!g3339) & (g3366) & (!g3340)) + ((!g827) & (!g1831) & (!g1853) & (!g3339) & (g3366) & (g3340)) + ((!g827) & (!g1831) & (!g1853) & (g3339) & (g3366) & (!g3340)) + ((!g827) & (!g1831) & (!g1853) & (g3339) & (g3366) & (g3340)) + ((!g827) & (!g1831) & (g1853) & (!g3339) & (g3366) & (!g3340)) + ((!g827) & (!g1831) & (g1853) & (!g3339) & (g3366) & (g3340)) + ((!g827) & (!g1831) & (g1853) & (g3339) & (g3366) & (!g3340)) + ((!g827) & (!g1831) & (g1853) & (g3339) & (g3366) & (g3340)) + ((!g827) & (g1831) & (!g1853) & (!g3339) & (g3366) & (!g3340)) + ((!g827) & (g1831) & (!g1853) & (!g3339) & (g3366) & (g3340)) + ((!g827) & (g1831) & (!g1853) & (g3339) & (g3366) & (!g3340)) + ((!g827) & (g1831) & (!g1853) & (g3339) & (g3366) & (g3340)) + ((!g827) & (g1831) & (g1853) & (!g3339) & (g3366) & (!g3340)) + ((!g827) & (g1831) & (g1853) & (!g3339) & (g3366) & (g3340)) + ((!g827) & (g1831) & (g1853) & (g3339) & (g3366) & (!g3340)) + ((!g827) & (g1831) & (g1853) & (g3339) & (g3366) & (g3340)) + ((g827) & (!g1831) & (!g1853) & (!g3339) & (g3366) & (!g3340)) + ((g827) & (!g1831) & (!g1853) & (!g3339) & (g3366) & (g3340)) + ((g827) & (!g1831) & (!g1853) & (g3339) & (!g3366) & (!g3340)) + ((g827) & (!g1831) & (!g1853) & (g3339) & (g3366) & (g3340)) + ((g827) & (!g1831) & (g1853) & (!g3339) & (!g3366) & (!g3340)) + ((g827) & (!g1831) & (g1853) & (!g3339) & (!g3366) & (g3340)) + ((g827) & (!g1831) & (g1853) & (g3339) & (!g3366) & (g3340)) + ((g827) & (!g1831) & (g1853) & (g3339) & (g3366) & (!g3340)) + ((g827) & (g1831) & (!g1853) & (!g3339) & (!g3366) & (!g3340)) + ((g827) & (g1831) & (!g1853) & (!g3339) & (g3366) & (g3340)) + ((g827) & (g1831) & (!g1853) & (g3339) & (!g3366) & (!g3340)) + ((g827) & (g1831) & (!g1853) & (g3339) & (!g3366) & (g3340)) + ((g827) & (g1831) & (g1853) & (!g3339) & (!g3366) & (g3340)) + ((g827) & (g1831) & (g1853) & (!g3339) & (g3366) & (!g3340)) + ((g827) & (g1831) & (g1853) & (g3339) & (g3366) & (!g3340)) + ((g827) & (g1831) & (g1853) & (g3339) & (g3366) & (g3340)));
	assign g3368 = (((!g827) & (!g1839) & (!g1855) & (!g2759) & (g2790) & (!g3351)) + ((!g827) & (!g1839) & (!g1855) & (!g2759) & (g2790) & (g3351)) + ((!g827) & (!g1839) & (!g1855) & (g2759) & (g2790) & (!g3351)) + ((!g827) & (!g1839) & (!g1855) & (g2759) & (g2790) & (g3351)) + ((!g827) & (!g1839) & (g1855) & (!g2759) & (g2790) & (!g3351)) + ((!g827) & (!g1839) & (g1855) & (!g2759) & (g2790) & (g3351)) + ((!g827) & (!g1839) & (g1855) & (g2759) & (g2790) & (!g3351)) + ((!g827) & (!g1839) & (g1855) & (g2759) & (g2790) & (g3351)) + ((!g827) & (g1839) & (!g1855) & (!g2759) & (g2790) & (!g3351)) + ((!g827) & (g1839) & (!g1855) & (!g2759) & (g2790) & (g3351)) + ((!g827) & (g1839) & (!g1855) & (g2759) & (g2790) & (!g3351)) + ((!g827) & (g1839) & (!g1855) & (g2759) & (g2790) & (g3351)) + ((!g827) & (g1839) & (g1855) & (!g2759) & (g2790) & (!g3351)) + ((!g827) & (g1839) & (g1855) & (!g2759) & (g2790) & (g3351)) + ((!g827) & (g1839) & (g1855) & (g2759) & (g2790) & (!g3351)) + ((!g827) & (g1839) & (g1855) & (g2759) & (g2790) & (g3351)) + ((g827) & (!g1839) & (!g1855) & (!g2759) & (g2790) & (!g3351)) + ((g827) & (!g1839) & (!g1855) & (!g2759) & (g2790) & (g3351)) + ((g827) & (!g1839) & (!g1855) & (g2759) & (!g2790) & (!g3351)) + ((g827) & (!g1839) & (!g1855) & (g2759) & (g2790) & (g3351)) + ((g827) & (!g1839) & (g1855) & (!g2759) & (!g2790) & (!g3351)) + ((g827) & (!g1839) & (g1855) & (!g2759) & (!g2790) & (g3351)) + ((g827) & (!g1839) & (g1855) & (g2759) & (!g2790) & (g3351)) + ((g827) & (!g1839) & (g1855) & (g2759) & (g2790) & (!g3351)) + ((g827) & (g1839) & (!g1855) & (!g2759) & (!g2790) & (!g3351)) + ((g827) & (g1839) & (!g1855) & (!g2759) & (g2790) & (g3351)) + ((g827) & (g1839) & (!g1855) & (g2759) & (!g2790) & (!g3351)) + ((g827) & (g1839) & (!g1855) & (g2759) & (!g2790) & (g3351)) + ((g827) & (g1839) & (g1855) & (!g2759) & (!g2790) & (g3351)) + ((g827) & (g1839) & (g1855) & (!g2759) & (g2790) & (!g3351)) + ((g827) & (g1839) & (g1855) & (g2759) & (g2790) & (!g3351)) + ((g827) & (g1839) & (g1855) & (g2759) & (g2790) & (g3351)));
	assign g3369 = (((!g827) & (!g1817) & (!g1857) & (!g2760) & (g2793) & (!g3321)) + ((!g827) & (!g1817) & (!g1857) & (!g2760) & (g2793) & (g3321)) + ((!g827) & (!g1817) & (!g1857) & (g2760) & (g2793) & (!g3321)) + ((!g827) & (!g1817) & (!g1857) & (g2760) & (g2793) & (g3321)) + ((!g827) & (!g1817) & (g1857) & (!g2760) & (g2793) & (!g3321)) + ((!g827) & (!g1817) & (g1857) & (!g2760) & (g2793) & (g3321)) + ((!g827) & (!g1817) & (g1857) & (g2760) & (g2793) & (!g3321)) + ((!g827) & (!g1817) & (g1857) & (g2760) & (g2793) & (g3321)) + ((!g827) & (g1817) & (!g1857) & (!g2760) & (g2793) & (!g3321)) + ((!g827) & (g1817) & (!g1857) & (!g2760) & (g2793) & (g3321)) + ((!g827) & (g1817) & (!g1857) & (g2760) & (g2793) & (!g3321)) + ((!g827) & (g1817) & (!g1857) & (g2760) & (g2793) & (g3321)) + ((!g827) & (g1817) & (g1857) & (!g2760) & (g2793) & (!g3321)) + ((!g827) & (g1817) & (g1857) & (!g2760) & (g2793) & (g3321)) + ((!g827) & (g1817) & (g1857) & (g2760) & (g2793) & (!g3321)) + ((!g827) & (g1817) & (g1857) & (g2760) & (g2793) & (g3321)) + ((g827) & (!g1817) & (!g1857) & (!g2760) & (g2793) & (!g3321)) + ((g827) & (!g1817) & (!g1857) & (!g2760) & (g2793) & (g3321)) + ((g827) & (!g1817) & (!g1857) & (g2760) & (!g2793) & (!g3321)) + ((g827) & (!g1817) & (!g1857) & (g2760) & (g2793) & (g3321)) + ((g827) & (!g1817) & (g1857) & (!g2760) & (!g2793) & (!g3321)) + ((g827) & (!g1817) & (g1857) & (!g2760) & (!g2793) & (g3321)) + ((g827) & (!g1817) & (g1857) & (g2760) & (!g2793) & (g3321)) + ((g827) & (!g1817) & (g1857) & (g2760) & (g2793) & (!g3321)) + ((g827) & (g1817) & (!g1857) & (!g2760) & (!g2793) & (!g3321)) + ((g827) & (g1817) & (!g1857) & (!g2760) & (g2793) & (g3321)) + ((g827) & (g1817) & (!g1857) & (g2760) & (!g2793) & (!g3321)) + ((g827) & (g1817) & (!g1857) & (g2760) & (!g2793) & (g3321)) + ((g827) & (g1817) & (g1857) & (!g2760) & (!g2793) & (g3321)) + ((g827) & (g1817) & (g1857) & (!g2760) & (g2793) & (!g3321)) + ((g827) & (g1817) & (g1857) & (g2760) & (g2793) & (!g3321)) + ((g827) & (g1817) & (g1857) & (g2760) & (g2793) & (g3321)));
	assign g8266 = (((!g2017) & (g5844) & (!g3370)) + ((!g2017) & (g5844) & (g3370)) + ((g2017) & (!g5844) & (g3370)) + ((g2017) & (g5844) & (g3370)));
	assign g3371 = (((!g827) & (!g1825) & (!g1859) & (!g3330) & (g3370) & (!g3331)) + ((!g827) & (!g1825) & (!g1859) & (!g3330) & (g3370) & (g3331)) + ((!g827) & (!g1825) & (!g1859) & (g3330) & (g3370) & (!g3331)) + ((!g827) & (!g1825) & (!g1859) & (g3330) & (g3370) & (g3331)) + ((!g827) & (!g1825) & (g1859) & (!g3330) & (g3370) & (!g3331)) + ((!g827) & (!g1825) & (g1859) & (!g3330) & (g3370) & (g3331)) + ((!g827) & (!g1825) & (g1859) & (g3330) & (g3370) & (!g3331)) + ((!g827) & (!g1825) & (g1859) & (g3330) & (g3370) & (g3331)) + ((!g827) & (g1825) & (!g1859) & (!g3330) & (g3370) & (!g3331)) + ((!g827) & (g1825) & (!g1859) & (!g3330) & (g3370) & (g3331)) + ((!g827) & (g1825) & (!g1859) & (g3330) & (g3370) & (!g3331)) + ((!g827) & (g1825) & (!g1859) & (g3330) & (g3370) & (g3331)) + ((!g827) & (g1825) & (g1859) & (!g3330) & (g3370) & (!g3331)) + ((!g827) & (g1825) & (g1859) & (!g3330) & (g3370) & (g3331)) + ((!g827) & (g1825) & (g1859) & (g3330) & (g3370) & (!g3331)) + ((!g827) & (g1825) & (g1859) & (g3330) & (g3370) & (g3331)) + ((g827) & (!g1825) & (!g1859) & (!g3330) & (g3370) & (!g3331)) + ((g827) & (!g1825) & (!g1859) & (!g3330) & (g3370) & (g3331)) + ((g827) & (!g1825) & (!g1859) & (g3330) & (!g3370) & (!g3331)) + ((g827) & (!g1825) & (!g1859) & (g3330) & (g3370) & (g3331)) + ((g827) & (!g1825) & (g1859) & (!g3330) & (!g3370) & (!g3331)) + ((g827) & (!g1825) & (g1859) & (!g3330) & (!g3370) & (g3331)) + ((g827) & (!g1825) & (g1859) & (g3330) & (!g3370) & (g3331)) + ((g827) & (!g1825) & (g1859) & (g3330) & (g3370) & (!g3331)) + ((g827) & (g1825) & (!g1859) & (!g3330) & (!g3370) & (!g3331)) + ((g827) & (g1825) & (!g1859) & (!g3330) & (g3370) & (g3331)) + ((g827) & (g1825) & (!g1859) & (g3330) & (!g3370) & (!g3331)) + ((g827) & (g1825) & (!g1859) & (g3330) & (!g3370) & (g3331)) + ((g827) & (g1825) & (g1859) & (!g3330) & (!g3370) & (g3331)) + ((g827) & (g1825) & (g1859) & (!g3330) & (g3370) & (!g3331)) + ((g827) & (g1825) & (g1859) & (g3330) & (g3370) & (!g3331)) + ((g827) & (g1825) & (g1859) & (g3330) & (g3370) & (g3331)));
	assign g8267 = (((!g3464) & (g5534) & (!g3372)) + ((!g3464) & (g5534) & (g3372)) + ((g3464) & (!g5534) & (g3372)) + ((g3464) & (g5534) & (g3372)));
	assign g3373 = (((!g827) & (!g1833) & (!g1861) & (!g3342) & (g3372) & (!g3343)) + ((!g827) & (!g1833) & (!g1861) & (!g3342) & (g3372) & (g3343)) + ((!g827) & (!g1833) & (!g1861) & (g3342) & (g3372) & (!g3343)) + ((!g827) & (!g1833) & (!g1861) & (g3342) & (g3372) & (g3343)) + ((!g827) & (!g1833) & (g1861) & (!g3342) & (g3372) & (!g3343)) + ((!g827) & (!g1833) & (g1861) & (!g3342) & (g3372) & (g3343)) + ((!g827) & (!g1833) & (g1861) & (g3342) & (g3372) & (!g3343)) + ((!g827) & (!g1833) & (g1861) & (g3342) & (g3372) & (g3343)) + ((!g827) & (g1833) & (!g1861) & (!g3342) & (g3372) & (!g3343)) + ((!g827) & (g1833) & (!g1861) & (!g3342) & (g3372) & (g3343)) + ((!g827) & (g1833) & (!g1861) & (g3342) & (g3372) & (!g3343)) + ((!g827) & (g1833) & (!g1861) & (g3342) & (g3372) & (g3343)) + ((!g827) & (g1833) & (g1861) & (!g3342) & (g3372) & (!g3343)) + ((!g827) & (g1833) & (g1861) & (!g3342) & (g3372) & (g3343)) + ((!g827) & (g1833) & (g1861) & (g3342) & (g3372) & (!g3343)) + ((!g827) & (g1833) & (g1861) & (g3342) & (g3372) & (g3343)) + ((g827) & (!g1833) & (!g1861) & (!g3342) & (g3372) & (!g3343)) + ((g827) & (!g1833) & (!g1861) & (!g3342) & (g3372) & (g3343)) + ((g827) & (!g1833) & (!g1861) & (g3342) & (!g3372) & (!g3343)) + ((g827) & (!g1833) & (!g1861) & (g3342) & (g3372) & (g3343)) + ((g827) & (!g1833) & (g1861) & (!g3342) & (!g3372) & (!g3343)) + ((g827) & (!g1833) & (g1861) & (!g3342) & (!g3372) & (g3343)) + ((g827) & (!g1833) & (g1861) & (g3342) & (!g3372) & (g3343)) + ((g827) & (!g1833) & (g1861) & (g3342) & (g3372) & (!g3343)) + ((g827) & (g1833) & (!g1861) & (!g3342) & (!g3372) & (!g3343)) + ((g827) & (g1833) & (!g1861) & (!g3342) & (g3372) & (g3343)) + ((g827) & (g1833) & (!g1861) & (g3342) & (!g3372) & (!g3343)) + ((g827) & (g1833) & (!g1861) & (g3342) & (!g3372) & (g3343)) + ((g827) & (g1833) & (g1861) & (!g3342) & (!g3372) & (g3343)) + ((g827) & (g1833) & (g1861) & (!g3342) & (g3372) & (!g3343)) + ((g827) & (g1833) & (g1861) & (g3342) & (g3372) & (!g3343)) + ((g827) & (g1833) & (g1861) & (g3342) & (g3372) & (g3343)));
	assign g8268 = (((!g3499) & (g5537) & (!g3374)) + ((!g3499) & (g5537) & (g3374)) + ((g3499) & (!g5537) & (g3374)) + ((g3499) & (g5537) & (g3374)));
	assign g3375 = (((!g827) & (!g1841) & (!g1863) & (!g3353) & (g3374) & (!g3354)) + ((!g827) & (!g1841) & (!g1863) & (!g3353) & (g3374) & (g3354)) + ((!g827) & (!g1841) & (!g1863) & (g3353) & (g3374) & (!g3354)) + ((!g827) & (!g1841) & (!g1863) & (g3353) & (g3374) & (g3354)) + ((!g827) & (!g1841) & (g1863) & (!g3353) & (g3374) & (!g3354)) + ((!g827) & (!g1841) & (g1863) & (!g3353) & (g3374) & (g3354)) + ((!g827) & (!g1841) & (g1863) & (g3353) & (g3374) & (!g3354)) + ((!g827) & (!g1841) & (g1863) & (g3353) & (g3374) & (g3354)) + ((!g827) & (g1841) & (!g1863) & (!g3353) & (g3374) & (!g3354)) + ((!g827) & (g1841) & (!g1863) & (!g3353) & (g3374) & (g3354)) + ((!g827) & (g1841) & (!g1863) & (g3353) & (g3374) & (!g3354)) + ((!g827) & (g1841) & (!g1863) & (g3353) & (g3374) & (g3354)) + ((!g827) & (g1841) & (g1863) & (!g3353) & (g3374) & (!g3354)) + ((!g827) & (g1841) & (g1863) & (!g3353) & (g3374) & (g3354)) + ((!g827) & (g1841) & (g1863) & (g3353) & (g3374) & (!g3354)) + ((!g827) & (g1841) & (g1863) & (g3353) & (g3374) & (g3354)) + ((g827) & (!g1841) & (!g1863) & (!g3353) & (g3374) & (!g3354)) + ((g827) & (!g1841) & (!g1863) & (!g3353) & (g3374) & (g3354)) + ((g827) & (!g1841) & (!g1863) & (g3353) & (!g3374) & (!g3354)) + ((g827) & (!g1841) & (!g1863) & (g3353) & (g3374) & (g3354)) + ((g827) & (!g1841) & (g1863) & (!g3353) & (!g3374) & (!g3354)) + ((g827) & (!g1841) & (g1863) & (!g3353) & (!g3374) & (g3354)) + ((g827) & (!g1841) & (g1863) & (g3353) & (!g3374) & (g3354)) + ((g827) & (!g1841) & (g1863) & (g3353) & (g3374) & (!g3354)) + ((g827) & (g1841) & (!g1863) & (!g3353) & (!g3374) & (!g3354)) + ((g827) & (g1841) & (!g1863) & (!g3353) & (g3374) & (g3354)) + ((g827) & (g1841) & (!g1863) & (g3353) & (!g3374) & (!g3354)) + ((g827) & (g1841) & (!g1863) & (g3353) & (!g3374) & (g3354)) + ((g827) & (g1841) & (g1863) & (!g3353) & (!g3374) & (g3354)) + ((g827) & (g1841) & (g1863) & (!g3353) & (g3374) & (!g3354)) + ((g827) & (g1841) & (g1863) & (g3353) & (g3374) & (!g3354)) + ((g827) & (g1841) & (g1863) & (g3353) & (g3374) & (g3354)));
	assign g8269 = (((!g3464) & (g5540) & (!g3376)) + ((!g3464) & (g5540) & (g3376)) + ((g3464) & (!g5540) & (g3376)) + ((g3464) & (g5540) & (g3376)));
	assign g3377 = (((!g827) & (!g1819) & (!g1865) & (!g3323) & (g3376) & (!g3324)) + ((!g827) & (!g1819) & (!g1865) & (!g3323) & (g3376) & (g3324)) + ((!g827) & (!g1819) & (!g1865) & (g3323) & (g3376) & (!g3324)) + ((!g827) & (!g1819) & (!g1865) & (g3323) & (g3376) & (g3324)) + ((!g827) & (!g1819) & (g1865) & (!g3323) & (g3376) & (!g3324)) + ((!g827) & (!g1819) & (g1865) & (!g3323) & (g3376) & (g3324)) + ((!g827) & (!g1819) & (g1865) & (g3323) & (g3376) & (!g3324)) + ((!g827) & (!g1819) & (g1865) & (g3323) & (g3376) & (g3324)) + ((!g827) & (g1819) & (!g1865) & (!g3323) & (g3376) & (!g3324)) + ((!g827) & (g1819) & (!g1865) & (!g3323) & (g3376) & (g3324)) + ((!g827) & (g1819) & (!g1865) & (g3323) & (g3376) & (!g3324)) + ((!g827) & (g1819) & (!g1865) & (g3323) & (g3376) & (g3324)) + ((!g827) & (g1819) & (g1865) & (!g3323) & (g3376) & (!g3324)) + ((!g827) & (g1819) & (g1865) & (!g3323) & (g3376) & (g3324)) + ((!g827) & (g1819) & (g1865) & (g3323) & (g3376) & (!g3324)) + ((!g827) & (g1819) & (g1865) & (g3323) & (g3376) & (g3324)) + ((g827) & (!g1819) & (!g1865) & (!g3323) & (g3376) & (!g3324)) + ((g827) & (!g1819) & (!g1865) & (!g3323) & (g3376) & (g3324)) + ((g827) & (!g1819) & (!g1865) & (g3323) & (!g3376) & (!g3324)) + ((g827) & (!g1819) & (!g1865) & (g3323) & (g3376) & (g3324)) + ((g827) & (!g1819) & (g1865) & (!g3323) & (!g3376) & (!g3324)) + ((g827) & (!g1819) & (g1865) & (!g3323) & (!g3376) & (g3324)) + ((g827) & (!g1819) & (g1865) & (g3323) & (!g3376) & (g3324)) + ((g827) & (!g1819) & (g1865) & (g3323) & (g3376) & (!g3324)) + ((g827) & (g1819) & (!g1865) & (!g3323) & (!g3376) & (!g3324)) + ((g827) & (g1819) & (!g1865) & (!g3323) & (g3376) & (g3324)) + ((g827) & (g1819) & (!g1865) & (g3323) & (!g3376) & (!g3324)) + ((g827) & (g1819) & (!g1865) & (g3323) & (!g3376) & (g3324)) + ((g827) & (g1819) & (g1865) & (!g3323) & (!g3376) & (g3324)) + ((g827) & (g1819) & (g1865) & (!g3323) & (g3376) & (!g3324)) + ((g827) & (g1819) & (g1865) & (g3323) & (g3376) & (!g3324)) + ((g827) & (g1819) & (g1865) & (g3323) & (g3376) & (g3324)));
	assign g8270 = (((!g3499) & (g5543) & (!g3378)) + ((!g3499) & (g5543) & (g3378)) + ((g3499) & (!g5543) & (g3378)) + ((g3499) & (g5543) & (g3378)));
	assign g3379 = (((!g827) & (!g1827) & (!g1867) & (!g3333) & (g3378) & (!g3334)) + ((!g827) & (!g1827) & (!g1867) & (!g3333) & (g3378) & (g3334)) + ((!g827) & (!g1827) & (!g1867) & (g3333) & (g3378) & (!g3334)) + ((!g827) & (!g1827) & (!g1867) & (g3333) & (g3378) & (g3334)) + ((!g827) & (!g1827) & (g1867) & (!g3333) & (g3378) & (!g3334)) + ((!g827) & (!g1827) & (g1867) & (!g3333) & (g3378) & (g3334)) + ((!g827) & (!g1827) & (g1867) & (g3333) & (g3378) & (!g3334)) + ((!g827) & (!g1827) & (g1867) & (g3333) & (g3378) & (g3334)) + ((!g827) & (g1827) & (!g1867) & (!g3333) & (g3378) & (!g3334)) + ((!g827) & (g1827) & (!g1867) & (!g3333) & (g3378) & (g3334)) + ((!g827) & (g1827) & (!g1867) & (g3333) & (g3378) & (!g3334)) + ((!g827) & (g1827) & (!g1867) & (g3333) & (g3378) & (g3334)) + ((!g827) & (g1827) & (g1867) & (!g3333) & (g3378) & (!g3334)) + ((!g827) & (g1827) & (g1867) & (!g3333) & (g3378) & (g3334)) + ((!g827) & (g1827) & (g1867) & (g3333) & (g3378) & (!g3334)) + ((!g827) & (g1827) & (g1867) & (g3333) & (g3378) & (g3334)) + ((g827) & (!g1827) & (!g1867) & (!g3333) & (g3378) & (!g3334)) + ((g827) & (!g1827) & (!g1867) & (!g3333) & (g3378) & (g3334)) + ((g827) & (!g1827) & (!g1867) & (g3333) & (!g3378) & (!g3334)) + ((g827) & (!g1827) & (!g1867) & (g3333) & (g3378) & (g3334)) + ((g827) & (!g1827) & (g1867) & (!g3333) & (!g3378) & (!g3334)) + ((g827) & (!g1827) & (g1867) & (!g3333) & (!g3378) & (g3334)) + ((g827) & (!g1827) & (g1867) & (g3333) & (!g3378) & (g3334)) + ((g827) & (!g1827) & (g1867) & (g3333) & (g3378) & (!g3334)) + ((g827) & (g1827) & (!g1867) & (!g3333) & (!g3378) & (!g3334)) + ((g827) & (g1827) & (!g1867) & (!g3333) & (g3378) & (g3334)) + ((g827) & (g1827) & (!g1867) & (g3333) & (!g3378) & (!g3334)) + ((g827) & (g1827) & (!g1867) & (g3333) & (!g3378) & (g3334)) + ((g827) & (g1827) & (g1867) & (!g3333) & (!g3378) & (g3334)) + ((g827) & (g1827) & (g1867) & (!g3333) & (g3378) & (!g3334)) + ((g827) & (g1827) & (g1867) & (g3333) & (g3378) & (!g3334)) + ((g827) & (g1827) & (g1867) & (g3333) & (g3378) & (g3334)));
	assign g8271 = (((!g2017) & (g5838) & (!g3380)) + ((!g2017) & (g5838) & (g3380)) + ((g2017) & (!g5838) & (g3380)) + ((g2017) & (g5838) & (g3380)));
	assign g3381 = (((!g827) & (!g1835) & (!g1869) & (!g3345) & (g3380) & (!g3346)) + ((!g827) & (!g1835) & (!g1869) & (!g3345) & (g3380) & (g3346)) + ((!g827) & (!g1835) & (!g1869) & (g3345) & (g3380) & (!g3346)) + ((!g827) & (!g1835) & (!g1869) & (g3345) & (g3380) & (g3346)) + ((!g827) & (!g1835) & (g1869) & (!g3345) & (g3380) & (!g3346)) + ((!g827) & (!g1835) & (g1869) & (!g3345) & (g3380) & (g3346)) + ((!g827) & (!g1835) & (g1869) & (g3345) & (g3380) & (!g3346)) + ((!g827) & (!g1835) & (g1869) & (g3345) & (g3380) & (g3346)) + ((!g827) & (g1835) & (!g1869) & (!g3345) & (g3380) & (!g3346)) + ((!g827) & (g1835) & (!g1869) & (!g3345) & (g3380) & (g3346)) + ((!g827) & (g1835) & (!g1869) & (g3345) & (g3380) & (!g3346)) + ((!g827) & (g1835) & (!g1869) & (g3345) & (g3380) & (g3346)) + ((!g827) & (g1835) & (g1869) & (!g3345) & (g3380) & (!g3346)) + ((!g827) & (g1835) & (g1869) & (!g3345) & (g3380) & (g3346)) + ((!g827) & (g1835) & (g1869) & (g3345) & (g3380) & (!g3346)) + ((!g827) & (g1835) & (g1869) & (g3345) & (g3380) & (g3346)) + ((g827) & (!g1835) & (!g1869) & (!g3345) & (g3380) & (!g3346)) + ((g827) & (!g1835) & (!g1869) & (!g3345) & (g3380) & (g3346)) + ((g827) & (!g1835) & (!g1869) & (g3345) & (!g3380) & (!g3346)) + ((g827) & (!g1835) & (!g1869) & (g3345) & (g3380) & (g3346)) + ((g827) & (!g1835) & (g1869) & (!g3345) & (!g3380) & (!g3346)) + ((g827) & (!g1835) & (g1869) & (!g3345) & (!g3380) & (g3346)) + ((g827) & (!g1835) & (g1869) & (g3345) & (!g3380) & (g3346)) + ((g827) & (!g1835) & (g1869) & (g3345) & (g3380) & (!g3346)) + ((g827) & (g1835) & (!g1869) & (!g3345) & (!g3380) & (!g3346)) + ((g827) & (g1835) & (!g1869) & (!g3345) & (g3380) & (g3346)) + ((g827) & (g1835) & (!g1869) & (g3345) & (!g3380) & (!g3346)) + ((g827) & (g1835) & (!g1869) & (g3345) & (!g3380) & (g3346)) + ((g827) & (g1835) & (g1869) & (!g3345) & (!g3380) & (g3346)) + ((g827) & (g1835) & (g1869) & (!g3345) & (g3380) & (!g3346)) + ((g827) & (g1835) & (g1869) & (g3345) & (g3380) & (!g3346)) + ((g827) & (g1835) & (g1869) & (g3345) & (g3380) & (g3346)));
	assign g8272 = (((!g3429) & (g5549) & (!g3382)) + ((!g3429) & (g5549) & (g3382)) + ((g3429) & (!g5549) & (g3382)) + ((g3429) & (g5549) & (g3382)));
	assign g3383 = (((!g827) & (!g1843) & (!g1871) & (!g3356) & (g3382) & (!g3357)) + ((!g827) & (!g1843) & (!g1871) & (!g3356) & (g3382) & (g3357)) + ((!g827) & (!g1843) & (!g1871) & (g3356) & (g3382) & (!g3357)) + ((!g827) & (!g1843) & (!g1871) & (g3356) & (g3382) & (g3357)) + ((!g827) & (!g1843) & (g1871) & (!g3356) & (g3382) & (!g3357)) + ((!g827) & (!g1843) & (g1871) & (!g3356) & (g3382) & (g3357)) + ((!g827) & (!g1843) & (g1871) & (g3356) & (g3382) & (!g3357)) + ((!g827) & (!g1843) & (g1871) & (g3356) & (g3382) & (g3357)) + ((!g827) & (g1843) & (!g1871) & (!g3356) & (g3382) & (!g3357)) + ((!g827) & (g1843) & (!g1871) & (!g3356) & (g3382) & (g3357)) + ((!g827) & (g1843) & (!g1871) & (g3356) & (g3382) & (!g3357)) + ((!g827) & (g1843) & (!g1871) & (g3356) & (g3382) & (g3357)) + ((!g827) & (g1843) & (g1871) & (!g3356) & (g3382) & (!g3357)) + ((!g827) & (g1843) & (g1871) & (!g3356) & (g3382) & (g3357)) + ((!g827) & (g1843) & (g1871) & (g3356) & (g3382) & (!g3357)) + ((!g827) & (g1843) & (g1871) & (g3356) & (g3382) & (g3357)) + ((g827) & (!g1843) & (!g1871) & (!g3356) & (g3382) & (!g3357)) + ((g827) & (!g1843) & (!g1871) & (!g3356) & (g3382) & (g3357)) + ((g827) & (!g1843) & (!g1871) & (g3356) & (!g3382) & (!g3357)) + ((g827) & (!g1843) & (!g1871) & (g3356) & (g3382) & (g3357)) + ((g827) & (!g1843) & (g1871) & (!g3356) & (!g3382) & (!g3357)) + ((g827) & (!g1843) & (g1871) & (!g3356) & (!g3382) & (g3357)) + ((g827) & (!g1843) & (g1871) & (g3356) & (!g3382) & (g3357)) + ((g827) & (!g1843) & (g1871) & (g3356) & (g3382) & (!g3357)) + ((g827) & (g1843) & (!g1871) & (!g3356) & (!g3382) & (!g3357)) + ((g827) & (g1843) & (!g1871) & (!g3356) & (g3382) & (g3357)) + ((g827) & (g1843) & (!g1871) & (g3356) & (!g3382) & (!g3357)) + ((g827) & (g1843) & (!g1871) & (g3356) & (!g3382) & (g3357)) + ((g827) & (g1843) & (g1871) & (!g3356) & (!g3382) & (g3357)) + ((g827) & (g1843) & (g1871) & (!g3356) & (g3382) & (!g3357)) + ((g827) & (g1843) & (g1871) & (g3356) & (g3382) & (!g3357)) + ((g827) & (g1843) & (g1871) & (g3356) & (g3382) & (g3357)));
	assign g3384 = (((!g827) & (!g1821) & (!g1873) & (!g2761) & (g2794) & (!g3326)) + ((!g827) & (!g1821) & (!g1873) & (!g2761) & (g2794) & (g3326)) + ((!g827) & (!g1821) & (!g1873) & (g2761) & (g2794) & (!g3326)) + ((!g827) & (!g1821) & (!g1873) & (g2761) & (g2794) & (g3326)) + ((!g827) & (!g1821) & (g1873) & (!g2761) & (g2794) & (!g3326)) + ((!g827) & (!g1821) & (g1873) & (!g2761) & (g2794) & (g3326)) + ((!g827) & (!g1821) & (g1873) & (g2761) & (g2794) & (!g3326)) + ((!g827) & (!g1821) & (g1873) & (g2761) & (g2794) & (g3326)) + ((!g827) & (g1821) & (!g1873) & (!g2761) & (g2794) & (!g3326)) + ((!g827) & (g1821) & (!g1873) & (!g2761) & (g2794) & (g3326)) + ((!g827) & (g1821) & (!g1873) & (g2761) & (g2794) & (!g3326)) + ((!g827) & (g1821) & (!g1873) & (g2761) & (g2794) & (g3326)) + ((!g827) & (g1821) & (g1873) & (!g2761) & (g2794) & (!g3326)) + ((!g827) & (g1821) & (g1873) & (!g2761) & (g2794) & (g3326)) + ((!g827) & (g1821) & (g1873) & (g2761) & (g2794) & (!g3326)) + ((!g827) & (g1821) & (g1873) & (g2761) & (g2794) & (g3326)) + ((g827) & (!g1821) & (!g1873) & (!g2761) & (g2794) & (!g3326)) + ((g827) & (!g1821) & (!g1873) & (!g2761) & (g2794) & (g3326)) + ((g827) & (!g1821) & (!g1873) & (g2761) & (!g2794) & (!g3326)) + ((g827) & (!g1821) & (!g1873) & (g2761) & (g2794) & (g3326)) + ((g827) & (!g1821) & (g1873) & (!g2761) & (!g2794) & (!g3326)) + ((g827) & (!g1821) & (g1873) & (!g2761) & (!g2794) & (g3326)) + ((g827) & (!g1821) & (g1873) & (g2761) & (!g2794) & (g3326)) + ((g827) & (!g1821) & (g1873) & (g2761) & (g2794) & (!g3326)) + ((g827) & (g1821) & (!g1873) & (!g2761) & (!g2794) & (!g3326)) + ((g827) & (g1821) & (!g1873) & (!g2761) & (g2794) & (g3326)) + ((g827) & (g1821) & (!g1873) & (g2761) & (!g2794) & (!g3326)) + ((g827) & (g1821) & (!g1873) & (g2761) & (!g2794) & (g3326)) + ((g827) & (g1821) & (g1873) & (!g2761) & (!g2794) & (g3326)) + ((g827) & (g1821) & (g1873) & (!g2761) & (g2794) & (!g3326)) + ((g827) & (g1821) & (g1873) & (g2761) & (g2794) & (!g3326)) + ((g827) & (g1821) & (g1873) & (g2761) & (g2794) & (g3326)));
	assign g8273 = (((!g3464) & (g5552) & (!g3385)) + ((!g3464) & (g5552) & (g3385)) + ((g3464) & (!g5552) & (g3385)) + ((g3464) & (g5552) & (g3385)));
	assign g3386 = (((!g827) & (!g1829) & (!g1875) & (!g3336) & (g3385) & (!g3337)) + ((!g827) & (!g1829) & (!g1875) & (!g3336) & (g3385) & (g3337)) + ((!g827) & (!g1829) & (!g1875) & (g3336) & (g3385) & (!g3337)) + ((!g827) & (!g1829) & (!g1875) & (g3336) & (g3385) & (g3337)) + ((!g827) & (!g1829) & (g1875) & (!g3336) & (g3385) & (!g3337)) + ((!g827) & (!g1829) & (g1875) & (!g3336) & (g3385) & (g3337)) + ((!g827) & (!g1829) & (g1875) & (g3336) & (g3385) & (!g3337)) + ((!g827) & (!g1829) & (g1875) & (g3336) & (g3385) & (g3337)) + ((!g827) & (g1829) & (!g1875) & (!g3336) & (g3385) & (!g3337)) + ((!g827) & (g1829) & (!g1875) & (!g3336) & (g3385) & (g3337)) + ((!g827) & (g1829) & (!g1875) & (g3336) & (g3385) & (!g3337)) + ((!g827) & (g1829) & (!g1875) & (g3336) & (g3385) & (g3337)) + ((!g827) & (g1829) & (g1875) & (!g3336) & (g3385) & (!g3337)) + ((!g827) & (g1829) & (g1875) & (!g3336) & (g3385) & (g3337)) + ((!g827) & (g1829) & (g1875) & (g3336) & (g3385) & (!g3337)) + ((!g827) & (g1829) & (g1875) & (g3336) & (g3385) & (g3337)) + ((g827) & (!g1829) & (!g1875) & (!g3336) & (g3385) & (!g3337)) + ((g827) & (!g1829) & (!g1875) & (!g3336) & (g3385) & (g3337)) + ((g827) & (!g1829) & (!g1875) & (g3336) & (!g3385) & (!g3337)) + ((g827) & (!g1829) & (!g1875) & (g3336) & (g3385) & (g3337)) + ((g827) & (!g1829) & (g1875) & (!g3336) & (!g3385) & (!g3337)) + ((g827) & (!g1829) & (g1875) & (!g3336) & (!g3385) & (g3337)) + ((g827) & (!g1829) & (g1875) & (g3336) & (!g3385) & (g3337)) + ((g827) & (!g1829) & (g1875) & (g3336) & (g3385) & (!g3337)) + ((g827) & (g1829) & (!g1875) & (!g3336) & (!g3385) & (!g3337)) + ((g827) & (g1829) & (!g1875) & (!g3336) & (g3385) & (g3337)) + ((g827) & (g1829) & (!g1875) & (g3336) & (!g3385) & (!g3337)) + ((g827) & (g1829) & (!g1875) & (g3336) & (!g3385) & (g3337)) + ((g827) & (g1829) & (g1875) & (!g3336) & (!g3385) & (g3337)) + ((g827) & (g1829) & (g1875) & (!g3336) & (g3385) & (!g3337)) + ((g827) & (g1829) & (g1875) & (g3336) & (g3385) & (!g3337)) + ((g827) & (g1829) & (g1875) & (g3336) & (g3385) & (g3337)));
	assign g8274 = (((!g3429) & (g5557) & (!g3387)) + ((!g3429) & (g5557) & (g3387)) + ((g3429) & (!g5557) & (g3387)) + ((g3429) & (g5557) & (g3387)));
	assign g3388 = (((!g827) & (!g1837) & (!g1877) & (!g3348) & (g3387) & (!g3349)) + ((!g827) & (!g1837) & (!g1877) & (!g3348) & (g3387) & (g3349)) + ((!g827) & (!g1837) & (!g1877) & (g3348) & (g3387) & (!g3349)) + ((!g827) & (!g1837) & (!g1877) & (g3348) & (g3387) & (g3349)) + ((!g827) & (!g1837) & (g1877) & (!g3348) & (g3387) & (!g3349)) + ((!g827) & (!g1837) & (g1877) & (!g3348) & (g3387) & (g3349)) + ((!g827) & (!g1837) & (g1877) & (g3348) & (g3387) & (!g3349)) + ((!g827) & (!g1837) & (g1877) & (g3348) & (g3387) & (g3349)) + ((!g827) & (g1837) & (!g1877) & (!g3348) & (g3387) & (!g3349)) + ((!g827) & (g1837) & (!g1877) & (!g3348) & (g3387) & (g3349)) + ((!g827) & (g1837) & (!g1877) & (g3348) & (g3387) & (!g3349)) + ((!g827) & (g1837) & (!g1877) & (g3348) & (g3387) & (g3349)) + ((!g827) & (g1837) & (g1877) & (!g3348) & (g3387) & (!g3349)) + ((!g827) & (g1837) & (g1877) & (!g3348) & (g3387) & (g3349)) + ((!g827) & (g1837) & (g1877) & (g3348) & (g3387) & (!g3349)) + ((!g827) & (g1837) & (g1877) & (g3348) & (g3387) & (g3349)) + ((g827) & (!g1837) & (!g1877) & (!g3348) & (g3387) & (!g3349)) + ((g827) & (!g1837) & (!g1877) & (!g3348) & (g3387) & (g3349)) + ((g827) & (!g1837) & (!g1877) & (g3348) & (!g3387) & (!g3349)) + ((g827) & (!g1837) & (!g1877) & (g3348) & (g3387) & (g3349)) + ((g827) & (!g1837) & (g1877) & (!g3348) & (!g3387) & (!g3349)) + ((g827) & (!g1837) & (g1877) & (!g3348) & (!g3387) & (g3349)) + ((g827) & (!g1837) & (g1877) & (g3348) & (!g3387) & (g3349)) + ((g827) & (!g1837) & (g1877) & (g3348) & (g3387) & (!g3349)) + ((g827) & (g1837) & (!g1877) & (!g3348) & (!g3387) & (!g3349)) + ((g827) & (g1837) & (!g1877) & (!g3348) & (g3387) & (g3349)) + ((g827) & (g1837) & (!g1877) & (g3348) & (!g3387) & (!g3349)) + ((g827) & (g1837) & (!g1877) & (g3348) & (!g3387) & (g3349)) + ((g827) & (g1837) & (g1877) & (!g3348) & (!g3387) & (g3349)) + ((g827) & (g1837) & (g1877) & (!g3348) & (g3387) & (!g3349)) + ((g827) & (g1837) & (g1877) & (g3348) & (g3387) & (!g3349)) + ((g827) & (g1837) & (g1877) & (g3348) & (g3387) & (g3349)));
	assign g8275 = (((!g2017) & (g5832) & (!g3389)) + ((!g2017) & (g5832) & (g3389)) + ((g2017) & (!g5832) & (g3389)) + ((g2017) & (g5832) & (g3389)));
	assign g3390 = (((!g827) & (!g1845) & (!g1879) & (!g3359) & (g3389) & (!g3360)) + ((!g827) & (!g1845) & (!g1879) & (!g3359) & (g3389) & (g3360)) + ((!g827) & (!g1845) & (!g1879) & (g3359) & (g3389) & (!g3360)) + ((!g827) & (!g1845) & (!g1879) & (g3359) & (g3389) & (g3360)) + ((!g827) & (!g1845) & (g1879) & (!g3359) & (g3389) & (!g3360)) + ((!g827) & (!g1845) & (g1879) & (!g3359) & (g3389) & (g3360)) + ((!g827) & (!g1845) & (g1879) & (g3359) & (g3389) & (!g3360)) + ((!g827) & (!g1845) & (g1879) & (g3359) & (g3389) & (g3360)) + ((!g827) & (g1845) & (!g1879) & (!g3359) & (g3389) & (!g3360)) + ((!g827) & (g1845) & (!g1879) & (!g3359) & (g3389) & (g3360)) + ((!g827) & (g1845) & (!g1879) & (g3359) & (g3389) & (!g3360)) + ((!g827) & (g1845) & (!g1879) & (g3359) & (g3389) & (g3360)) + ((!g827) & (g1845) & (g1879) & (!g3359) & (g3389) & (!g3360)) + ((!g827) & (g1845) & (g1879) & (!g3359) & (g3389) & (g3360)) + ((!g827) & (g1845) & (g1879) & (g3359) & (g3389) & (!g3360)) + ((!g827) & (g1845) & (g1879) & (g3359) & (g3389) & (g3360)) + ((g827) & (!g1845) & (!g1879) & (!g3359) & (g3389) & (!g3360)) + ((g827) & (!g1845) & (!g1879) & (!g3359) & (g3389) & (g3360)) + ((g827) & (!g1845) & (!g1879) & (g3359) & (!g3389) & (!g3360)) + ((g827) & (!g1845) & (!g1879) & (g3359) & (g3389) & (g3360)) + ((g827) & (!g1845) & (g1879) & (!g3359) & (!g3389) & (!g3360)) + ((g827) & (!g1845) & (g1879) & (!g3359) & (!g3389) & (g3360)) + ((g827) & (!g1845) & (g1879) & (g3359) & (!g3389) & (g3360)) + ((g827) & (!g1845) & (g1879) & (g3359) & (g3389) & (!g3360)) + ((g827) & (g1845) & (!g1879) & (!g3359) & (!g3389) & (!g3360)) + ((g827) & (g1845) & (!g1879) & (!g3359) & (g3389) & (g3360)) + ((g827) & (g1845) & (!g1879) & (g3359) & (!g3389) & (!g3360)) + ((g827) & (g1845) & (!g1879) & (g3359) & (!g3389) & (g3360)) + ((g827) & (g1845) & (g1879) & (!g3359) & (!g3389) & (g3360)) + ((g827) & (g1845) & (g1879) & (!g3359) & (g3389) & (!g3360)) + ((g827) & (g1845) & (g1879) & (g3359) & (g3389) & (!g3360)) + ((g827) & (g1845) & (g1879) & (g3359) & (g3389) & (g3360)));
	assign g3391 = (((!g2010) & (!g2011) & (!g2012)) + ((!g2010) & (g2011) & (g2012)) + ((g2010) & (!g2011) & (g2012)) + ((g2010) & (g2011) & (!g2012)));
	assign g3392 = (((!g1892) & (!g1908) & (!g2026) & (!g2030) & (g2062) & (g2085)) + ((!g1892) & (!g1908) & (!g2026) & (g2030) & (g2062) & (g2085)) + ((!g1892) & (!g1908) & (g2026) & (!g2030) & (g2062) & (g2085)) + ((!g1892) & (!g1908) & (g2026) & (g2030) & (!g2062) & (g2085)) + ((!g1892) & (!g1908) & (g2026) & (g2030) & (g2062) & (!g2085)) + ((!g1892) & (!g1908) & (g2026) & (g2030) & (g2062) & (g2085)) + ((!g1892) & (g1908) & (!g2026) & (!g2030) & (g2062) & (g2085)) + ((!g1892) & (g1908) & (!g2026) & (g2030) & (g2062) & (g2085)) + ((!g1892) & (g1908) & (g2026) & (!g2030) & (g2062) & (g2085)) + ((!g1892) & (g1908) & (g2026) & (g2030) & (!g2062) & (g2085)) + ((!g1892) & (g1908) & (g2026) & (g2030) & (g2062) & (!g2085)) + ((!g1892) & (g1908) & (g2026) & (g2030) & (g2062) & (g2085)) + ((g1892) & (!g1908) & (!g2026) & (!g2030) & (g2062) & (g2085)) + ((g1892) & (!g1908) & (!g2026) & (g2030) & (g2062) & (g2085)) + ((g1892) & (!g1908) & (g2026) & (!g2030) & (g2062) & (g2085)) + ((g1892) & (!g1908) & (g2026) & (g2030) & (!g2062) & (g2085)) + ((g1892) & (!g1908) & (g2026) & (g2030) & (g2062) & (!g2085)) + ((g1892) & (!g1908) & (g2026) & (g2030) & (g2062) & (g2085)) + ((g1892) & (g1908) & (!g2026) & (!g2030) & (g2062) & (g2085)) + ((g1892) & (g1908) & (!g2026) & (g2030) & (!g2062) & (g2085)) + ((g1892) & (g1908) & (!g2026) & (g2030) & (g2062) & (!g2085)) + ((g1892) & (g1908) & (!g2026) & (g2030) & (g2062) & (g2085)) + ((g1892) & (g1908) & (g2026) & (!g2030) & (!g2062) & (g2085)) + ((g1892) & (g1908) & (g2026) & (!g2030) & (g2062) & (!g2085)) + ((g1892) & (g1908) & (g2026) & (!g2030) & (g2062) & (g2085)) + ((g1892) & (g1908) & (g2026) & (g2030) & (!g2062) & (g2085)) + ((g1892) & (g1908) & (g2026) & (g2030) & (g2062) & (!g2085)) + ((g1892) & (g1908) & (g2026) & (g2030) & (g2062) & (g2085)));
	assign g3393 = (((!g2188) & (g2192)) + ((g2188) & (!g2192)));
	assign g3394 = (((!g3392) & (!g2108) & (!g2112) & (g2144) & (g2167) & (g3393)) + ((!g3392) & (!g2108) & (g2112) & (g2144) & (g2167) & (g3393)) + ((!g3392) & (g2108) & (!g2112) & (g2144) & (g2167) & (g3393)) + ((!g3392) & (g2108) & (g2112) & (!g2144) & (g2167) & (g3393)) + ((!g3392) & (g2108) & (g2112) & (g2144) & (!g2167) & (g3393)) + ((!g3392) & (g2108) & (g2112) & (g2144) & (g2167) & (g3393)) + ((g3392) & (!g2108) & (!g2112) & (g2144) & (g2167) & (g3393)) + ((g3392) & (!g2108) & (g2112) & (!g2144) & (g2167) & (g3393)) + ((g3392) & (!g2108) & (g2112) & (g2144) & (!g2167) & (g3393)) + ((g3392) & (!g2108) & (g2112) & (g2144) & (g2167) & (g3393)) + ((g3392) & (g2108) & (!g2112) & (!g2144) & (g2167) & (g3393)) + ((g3392) & (g2108) & (!g2112) & (g2144) & (!g2167) & (g3393)) + ((g3392) & (g2108) & (!g2112) & (g2144) & (g2167) & (g3393)) + ((g3392) & (g2108) & (g2112) & (!g2144) & (g2167) & (g3393)) + ((g3392) & (g2108) & (g2112) & (g2144) & (!g2167) & (g3393)) + ((g3392) & (g2108) & (g2112) & (g2144) & (g2167) & (g3393)));
	assign g3395 = (((g2188) & (g2192)));
	assign g3396 = (((!g3394) & (!g3395) & (!g2224) & (!g2247) & (!g2271) & (!g2275)) + ((!g3394) & (!g3395) & (!g2224) & (!g2247) & (!g2271) & (g2275)) + ((!g3394) & (!g3395) & (!g2224) & (!g2247) & (g2271) & (!g2275)) + ((!g3394) & (!g3395) & (!g2224) & (g2247) & (!g2271) & (!g2275)) + ((!g3394) & (!g3395) & (!g2224) & (g2247) & (!g2271) & (g2275)) + ((!g3394) & (!g3395) & (!g2224) & (g2247) & (g2271) & (!g2275)) + ((!g3394) & (!g3395) & (g2224) & (!g2247) & (!g2271) & (!g2275)) + ((!g3394) & (!g3395) & (g2224) & (!g2247) & (!g2271) & (g2275)) + ((!g3394) & (!g3395) & (g2224) & (!g2247) & (g2271) & (!g2275)) + ((!g3394) & (!g3395) & (g2224) & (g2247) & (!g2271) & (!g2275)) + ((!g3394) & (g3395) & (!g2224) & (!g2247) & (!g2271) & (!g2275)) + ((!g3394) & (g3395) & (!g2224) & (!g2247) & (!g2271) & (g2275)) + ((!g3394) & (g3395) & (!g2224) & (!g2247) & (g2271) & (!g2275)) + ((!g3394) & (g3395) & (!g2224) & (g2247) & (!g2271) & (!g2275)) + ((!g3394) & (g3395) & (g2224) & (!g2247) & (!g2271) & (!g2275)) + ((!g3394) & (g3395) & (g2224) & (g2247) & (!g2271) & (!g2275)) + ((g3394) & (!g3395) & (!g2224) & (!g2247) & (!g2271) & (!g2275)) + ((g3394) & (!g3395) & (!g2224) & (!g2247) & (!g2271) & (g2275)) + ((g3394) & (!g3395) & (!g2224) & (!g2247) & (g2271) & (!g2275)) + ((g3394) & (!g3395) & (!g2224) & (g2247) & (!g2271) & (!g2275)) + ((g3394) & (!g3395) & (g2224) & (!g2247) & (!g2271) & (!g2275)) + ((g3394) & (!g3395) & (g2224) & (g2247) & (!g2271) & (!g2275)) + ((g3394) & (g3395) & (!g2224) & (!g2247) & (!g2271) & (!g2275)) + ((g3394) & (g3395) & (!g2224) & (!g2247) & (!g2271) & (g2275)) + ((g3394) & (g3395) & (!g2224) & (!g2247) & (g2271) & (!g2275)) + ((g3394) & (g3395) & (!g2224) & (g2247) & (!g2271) & (!g2275)) + ((g3394) & (g3395) & (g2224) & (!g2247) & (!g2271) & (!g2275)) + ((g3394) & (g3395) & (g2224) & (g2247) & (!g2271) & (!g2275)));
	assign g3397 = (((!g2390) & (g2413)) + ((g2390) & (!g2413)));
	assign g3398 = (((!g3396) & (!g2311) & (!g2334) & (g2354) & (g2358) & (g3397)) + ((!g3396) & (!g2311) & (g2334) & (!g2354) & (g2358) & (g3397)) + ((!g3396) & (!g2311) & (g2334) & (g2354) & (!g2358) & (g3397)) + ((!g3396) & (!g2311) & (g2334) & (g2354) & (g2358) & (g3397)) + ((!g3396) & (g2311) & (!g2334) & (!g2354) & (g2358) & (g3397)) + ((!g3396) & (g2311) & (!g2334) & (g2354) & (!g2358) & (g3397)) + ((!g3396) & (g2311) & (!g2334) & (g2354) & (g2358) & (g3397)) + ((!g3396) & (g2311) & (g2334) & (!g2354) & (g2358) & (g3397)) + ((!g3396) & (g2311) & (g2334) & (g2354) & (!g2358) & (g3397)) + ((!g3396) & (g2311) & (g2334) & (g2354) & (g2358) & (g3397)) + ((g3396) & (!g2311) & (!g2334) & (g2354) & (g2358) & (g3397)) + ((g3396) & (!g2311) & (g2334) & (g2354) & (g2358) & (g3397)) + ((g3396) & (g2311) & (!g2334) & (g2354) & (g2358) & (g3397)) + ((g3396) & (g2311) & (g2334) & (!g2354) & (g2358) & (g3397)) + ((g3396) & (g2311) & (g2334) & (g2354) & (!g2358) & (g3397)) + ((g3396) & (g2311) & (g2334) & (g2354) & (g2358) & (g3397)));
	assign g3399 = (((g2390) & (g2413)));
	assign g3400 = (((!g3398) & (!g3399) & (!g2450) & (!g2462) & (!g2527) & (!g2542)) + ((!g3398) & (!g3399) & (!g2450) & (!g2462) & (!g2527) & (g2542)) + ((!g3398) & (!g3399) & (!g2450) & (!g2462) & (g2527) & (!g2542)) + ((!g3398) & (!g3399) & (!g2450) & (g2462) & (!g2527) & (!g2542)) + ((!g3398) & (!g3399) & (!g2450) & (g2462) & (!g2527) & (g2542)) + ((!g3398) & (!g3399) & (!g2450) & (g2462) & (g2527) & (!g2542)) + ((!g3398) & (!g3399) & (g2450) & (!g2462) & (!g2527) & (!g2542)) + ((!g3398) & (!g3399) & (g2450) & (!g2462) & (!g2527) & (g2542)) + ((!g3398) & (!g3399) & (g2450) & (!g2462) & (g2527) & (!g2542)) + ((!g3398) & (!g3399) & (g2450) & (g2462) & (!g2527) & (!g2542)) + ((!g3398) & (g3399) & (!g2450) & (!g2462) & (!g2527) & (!g2542)) + ((!g3398) & (g3399) & (!g2450) & (!g2462) & (!g2527) & (g2542)) + ((!g3398) & (g3399) & (!g2450) & (!g2462) & (g2527) & (!g2542)) + ((!g3398) & (g3399) & (!g2450) & (g2462) & (!g2527) & (!g2542)) + ((!g3398) & (g3399) & (g2450) & (!g2462) & (!g2527) & (!g2542)) + ((!g3398) & (g3399) & (g2450) & (g2462) & (!g2527) & (!g2542)) + ((g3398) & (!g3399) & (!g2450) & (!g2462) & (!g2527) & (!g2542)) + ((g3398) & (!g3399) & (!g2450) & (!g2462) & (!g2527) & (g2542)) + ((g3398) & (!g3399) & (!g2450) & (!g2462) & (g2527) & (!g2542)) + ((g3398) & (!g3399) & (!g2450) & (g2462) & (!g2527) & (!g2542)) + ((g3398) & (!g3399) & (g2450) & (!g2462) & (!g2527) & (!g2542)) + ((g3398) & (!g3399) & (g2450) & (g2462) & (!g2527) & (!g2542)) + ((g3398) & (g3399) & (!g2450) & (!g2462) & (!g2527) & (!g2542)) + ((g3398) & (g3399) & (!g2450) & (!g2462) & (!g2527) & (g2542)) + ((g3398) & (g3399) & (!g2450) & (!g2462) & (g2527) & (!g2542)) + ((g3398) & (g3399) & (!g2450) & (g2462) & (!g2527) & (!g2542)) + ((g3398) & (g3399) & (g2450) & (!g2462) & (!g2527) & (!g2542)) + ((g3398) & (g3399) & (g2450) & (g2462) & (!g2527) & (!g2542)));
	assign g3401 = (((!g2657) & (g2661)) + ((g2657) & (!g2661)));
	assign g3402 = (((!g3400) & (!g2566) & (!g2572) & (g2614) & (g2637) & (g3401)) + ((!g3400) & (!g2566) & (g2572) & (!g2614) & (g2637) & (g3401)) + ((!g3400) & (!g2566) & (g2572) & (g2614) & (!g2637) & (g3401)) + ((!g3400) & (!g2566) & (g2572) & (g2614) & (g2637) & (g3401)) + ((!g3400) & (g2566) & (!g2572) & (!g2614) & (g2637) & (g3401)) + ((!g3400) & (g2566) & (!g2572) & (g2614) & (!g2637) & (g3401)) + ((!g3400) & (g2566) & (!g2572) & (g2614) & (g2637) & (g3401)) + ((!g3400) & (g2566) & (g2572) & (!g2614) & (g2637) & (g3401)) + ((!g3400) & (g2566) & (g2572) & (g2614) & (!g2637) & (g3401)) + ((!g3400) & (g2566) & (g2572) & (g2614) & (g2637) & (g3401)) + ((g3400) & (!g2566) & (!g2572) & (g2614) & (g2637) & (g3401)) + ((g3400) & (!g2566) & (g2572) & (g2614) & (g2637) & (g3401)) + ((g3400) & (g2566) & (!g2572) & (g2614) & (g2637) & (g3401)) + ((g3400) & (g2566) & (g2572) & (!g2614) & (g2637) & (g3401)) + ((g3400) & (g2566) & (g2572) & (g2614) & (!g2637) & (g3401)) + ((g3400) & (g2566) & (g2572) & (g2614) & (g2637) & (g3401)));
	assign g3403 = (((g2657) & (g2661)));
	assign g3404 = (((!g3402) & (!g3403) & (!g2703) & (!g2742) & (!g2768) & (!g2772)) + ((!g3402) & (!g3403) & (!g2703) & (!g2742) & (!g2768) & (g2772)) + ((!g3402) & (!g3403) & (!g2703) & (!g2742) & (g2768) & (!g2772)) + ((!g3402) & (!g3403) & (!g2703) & (g2742) & (!g2768) & (!g2772)) + ((!g3402) & (!g3403) & (!g2703) & (g2742) & (!g2768) & (g2772)) + ((!g3402) & (!g3403) & (!g2703) & (g2742) & (g2768) & (!g2772)) + ((!g3402) & (!g3403) & (g2703) & (!g2742) & (!g2768) & (!g2772)) + ((!g3402) & (!g3403) & (g2703) & (!g2742) & (!g2768) & (g2772)) + ((!g3402) & (!g3403) & (g2703) & (!g2742) & (g2768) & (!g2772)) + ((!g3402) & (!g3403) & (g2703) & (g2742) & (!g2768) & (!g2772)) + ((!g3402) & (g3403) & (!g2703) & (!g2742) & (!g2768) & (!g2772)) + ((!g3402) & (g3403) & (!g2703) & (!g2742) & (!g2768) & (g2772)) + ((!g3402) & (g3403) & (!g2703) & (!g2742) & (g2768) & (!g2772)) + ((!g3402) & (g3403) & (!g2703) & (g2742) & (!g2768) & (!g2772)) + ((!g3402) & (g3403) & (g2703) & (!g2742) & (!g2768) & (!g2772)) + ((!g3402) & (g3403) & (g2703) & (g2742) & (!g2768) & (!g2772)) + ((g3402) & (!g3403) & (!g2703) & (!g2742) & (!g2768) & (!g2772)) + ((g3402) & (!g3403) & (!g2703) & (!g2742) & (!g2768) & (g2772)) + ((g3402) & (!g3403) & (!g2703) & (!g2742) & (g2768) & (!g2772)) + ((g3402) & (!g3403) & (!g2703) & (g2742) & (!g2768) & (!g2772)) + ((g3402) & (!g3403) & (g2703) & (!g2742) & (!g2768) & (!g2772)) + ((g3402) & (!g3403) & (g2703) & (g2742) & (!g2768) & (!g2772)) + ((g3402) & (g3403) & (!g2703) & (!g2742) & (!g2768) & (!g2772)) + ((g3402) & (g3403) & (!g2703) & (!g2742) & (!g2768) & (g2772)) + ((g3402) & (g3403) & (!g2703) & (!g2742) & (g2768) & (!g2772)) + ((g3402) & (g3403) & (!g2703) & (g2742) & (!g2768) & (!g2772)) + ((g3402) & (g3403) & (g2703) & (!g2742) & (!g2768) & (!g2772)) + ((g3402) & (g3403) & (g2703) & (g2742) & (!g2768) & (!g2772)));
	assign g3405 = (((!g2885) & (g2900)) + ((g2885) & (!g2900)));
	assign g3406 = (((!g3404) & (!g2804) & (!g2827) & (g2845) & (g2851) & (g3405)) + ((!g3404) & (!g2804) & (g2827) & (!g2845) & (g2851) & (g3405)) + ((!g3404) & (!g2804) & (g2827) & (g2845) & (!g2851) & (g3405)) + ((!g3404) & (!g2804) & (g2827) & (g2845) & (g2851) & (g3405)) + ((!g3404) & (g2804) & (!g2827) & (!g2845) & (g2851) & (g3405)) + ((!g3404) & (g2804) & (!g2827) & (g2845) & (!g2851) & (g3405)) + ((!g3404) & (g2804) & (!g2827) & (g2845) & (g2851) & (g3405)) + ((!g3404) & (g2804) & (g2827) & (!g2845) & (g2851) & (g3405)) + ((!g3404) & (g2804) & (g2827) & (g2845) & (!g2851) & (g3405)) + ((!g3404) & (g2804) & (g2827) & (g2845) & (g2851) & (g3405)) + ((g3404) & (!g2804) & (!g2827) & (g2845) & (g2851) & (g3405)) + ((g3404) & (!g2804) & (g2827) & (g2845) & (g2851) & (g3405)) + ((g3404) & (g2804) & (!g2827) & (g2845) & (g2851) & (g3405)) + ((g3404) & (g2804) & (g2827) & (!g2845) & (g2851) & (g3405)) + ((g3404) & (g2804) & (g2827) & (g2845) & (!g2851) & (g3405)) + ((g3404) & (g2804) & (g2827) & (g2845) & (g2851) & (g3405)));
	assign g3407 = (((g2885) & (g2900)));
	assign g3408 = (((!g3406) & (!g3407) & (!g2932) & (!g2944) & (!g3003) & (!g3018)) + ((!g3406) & (!g3407) & (!g2932) & (!g2944) & (!g3003) & (g3018)) + ((!g3406) & (!g3407) & (!g2932) & (!g2944) & (g3003) & (!g3018)) + ((!g3406) & (!g3407) & (!g2932) & (g2944) & (!g3003) & (!g3018)) + ((!g3406) & (!g3407) & (!g2932) & (g2944) & (!g3003) & (g3018)) + ((!g3406) & (!g3407) & (!g2932) & (g2944) & (g3003) & (!g3018)) + ((!g3406) & (!g3407) & (g2932) & (!g2944) & (!g3003) & (!g3018)) + ((!g3406) & (!g3407) & (g2932) & (!g2944) & (!g3003) & (g3018)) + ((!g3406) & (!g3407) & (g2932) & (!g2944) & (g3003) & (!g3018)) + ((!g3406) & (!g3407) & (g2932) & (g2944) & (!g3003) & (!g3018)) + ((!g3406) & (g3407) & (!g2932) & (!g2944) & (!g3003) & (!g3018)) + ((!g3406) & (g3407) & (!g2932) & (!g2944) & (!g3003) & (g3018)) + ((!g3406) & (g3407) & (!g2932) & (!g2944) & (g3003) & (!g3018)) + ((!g3406) & (g3407) & (!g2932) & (g2944) & (!g3003) & (!g3018)) + ((!g3406) & (g3407) & (g2932) & (!g2944) & (!g3003) & (!g3018)) + ((!g3406) & (g3407) & (g2932) & (g2944) & (!g3003) & (!g3018)) + ((g3406) & (!g3407) & (!g2932) & (!g2944) & (!g3003) & (!g3018)) + ((g3406) & (!g3407) & (!g2932) & (!g2944) & (!g3003) & (g3018)) + ((g3406) & (!g3407) & (!g2932) & (!g2944) & (g3003) & (!g3018)) + ((g3406) & (!g3407) & (!g2932) & (g2944) & (!g3003) & (!g3018)) + ((g3406) & (!g3407) & (g2932) & (!g2944) & (!g3003) & (!g3018)) + ((g3406) & (!g3407) & (g2932) & (g2944) & (!g3003) & (!g3018)) + ((g3406) & (g3407) & (!g2932) & (!g2944) & (!g3003) & (!g3018)) + ((g3406) & (g3407) & (!g2932) & (!g2944) & (!g3003) & (g3018)) + ((g3406) & (g3407) & (!g2932) & (!g2944) & (g3003) & (!g3018)) + ((g3406) & (g3407) & (!g2932) & (g2944) & (!g3003) & (!g3018)) + ((g3406) & (g3407) & (g2932) & (!g2944) & (!g3003) & (!g3018)) + ((g3406) & (g3407) & (g2932) & (g2944) & (!g3003) & (!g3018)));
	assign g3409 = (((!g3408) & (!g3038) & (!g3044)) + ((!g3408) & (g3038) & (g3044)) + ((g3408) & (!g3038) & (g3044)) + ((g3408) & (g3038) & (!g3044)));
	assign g3410 = (((!g828) & (!g864) & (g897) & (!g1886) & (!g2032) & (g2055)) + ((!g828) & (!g864) & (g897) & (!g1886) & (g2032) & (g2055)) + ((!g828) & (!g864) & (g897) & (g1886) & (!g2032) & (g2055)) + ((!g828) & (!g864) & (g897) & (g1886) & (g2032) & (g2055)) + ((!g828) & (g864) & (!g897) & (!g1886) & (g2032) & (g2055)) + ((!g828) & (g864) & (!g897) & (g1886) & (g2032) & (g2055)) + ((!g828) & (g864) & (g897) & (!g1886) & (!g2032) & (g2055)) + ((!g828) & (g864) & (g897) & (!g1886) & (g2032) & (!g2055)) + ((!g828) & (g864) & (g897) & (!g1886) & (g2032) & (g2055)) + ((!g828) & (g864) & (g897) & (g1886) & (!g2032) & (g2055)) + ((!g828) & (g864) & (g897) & (g1886) & (g2032) & (!g2055)) + ((!g828) & (g864) & (g897) & (g1886) & (g2032) & (g2055)) + ((g828) & (!g864) & (!g897) & (g1886) & (g2032) & (g2055)) + ((g828) & (!g864) & (g897) & (!g1886) & (!g2032) & (g2055)) + ((g828) & (!g864) & (g897) & (!g1886) & (g2032) & (g2055)) + ((g828) & (!g864) & (g897) & (g1886) & (!g2032) & (g2055)) + ((g828) & (!g864) & (g897) & (g1886) & (g2032) & (!g2055)) + ((g828) & (!g864) & (g897) & (g1886) & (g2032) & (g2055)) + ((g828) & (g864) & (!g897) & (!g1886) & (g2032) & (g2055)) + ((g828) & (g864) & (!g897) & (g1886) & (!g2032) & (g2055)) + ((g828) & (g864) & (!g897) & (g1886) & (g2032) & (g2055)) + ((g828) & (g864) & (g897) & (!g1886) & (!g2032) & (g2055)) + ((g828) & (g864) & (g897) & (!g1886) & (g2032) & (!g2055)) + ((g828) & (g864) & (g897) & (!g1886) & (g2032) & (g2055)) + ((g828) & (g864) & (g897) & (g1886) & (!g2032) & (!g2055)) + ((g828) & (g864) & (g897) & (g1886) & (!g2032) & (g2055)) + ((g828) & (g864) & (g897) & (g1886) & (g2032) & (!g2055)) + ((g828) & (g864) & (g897) & (g1886) & (g2032) & (g2055)));
	assign g3411 = (((!g998) & (g2194)) + ((g998) & (!g2194)));
	assign g3412 = (((!g931) & (!g964) & (g3410) & (g2114) & (g2137) & (g3411)) + ((!g931) & (g964) & (!g3410) & (!g2114) & (g2137) & (g3411)) + ((!g931) & (g964) & (!g3410) & (g2114) & (g2137) & (g3411)) + ((!g931) & (g964) & (g3410) & (!g2114) & (g2137) & (g3411)) + ((!g931) & (g964) & (g3410) & (g2114) & (!g2137) & (g3411)) + ((!g931) & (g964) & (g3410) & (g2114) & (g2137) & (g3411)) + ((g931) & (!g964) & (!g3410) & (g2114) & (g2137) & (g3411)) + ((g931) & (!g964) & (g3410) & (!g2114) & (g2137) & (g3411)) + ((g931) & (!g964) & (g3410) & (g2114) & (g2137) & (g3411)) + ((g931) & (g964) & (!g3410) & (!g2114) & (g2137) & (g3411)) + ((g931) & (g964) & (!g3410) & (g2114) & (!g2137) & (g3411)) + ((g931) & (g964) & (!g3410) & (g2114) & (g2137) & (g3411)) + ((g931) & (g964) & (g3410) & (!g2114) & (!g2137) & (g3411)) + ((g931) & (g964) & (g3410) & (!g2114) & (g2137) & (g3411)) + ((g931) & (g964) & (g3410) & (g2114) & (!g2137) & (g3411)) + ((g931) & (g964) & (g3410) & (g2114) & (g2137) & (g3411)));
	assign g3413 = (((g998) & (g2194)));
	assign g3414 = (((!g1031) & (!g1065) & (!g3412) & (!g3413) & (!g2217) & (!g2277)) + ((!g1031) & (!g1065) & (!g3412) & (!g3413) & (!g2217) & (g2277)) + ((!g1031) & (!g1065) & (!g3412) & (!g3413) & (g2217) & (!g2277)) + ((!g1031) & (!g1065) & (!g3412) & (!g3413) & (g2217) & (g2277)) + ((!g1031) & (!g1065) & (!g3412) & (g3413) & (!g2217) & (!g2277)) + ((!g1031) & (!g1065) & (!g3412) & (g3413) & (!g2217) & (g2277)) + ((!g1031) & (!g1065) & (!g3412) & (g3413) & (g2217) & (!g2277)) + ((!g1031) & (!g1065) & (g3412) & (!g3413) & (!g2217) & (!g2277)) + ((!g1031) & (!g1065) & (g3412) & (!g3413) & (!g2217) & (g2277)) + ((!g1031) & (!g1065) & (g3412) & (!g3413) & (g2217) & (!g2277)) + ((!g1031) & (!g1065) & (g3412) & (g3413) & (!g2217) & (!g2277)) + ((!g1031) & (!g1065) & (g3412) & (g3413) & (!g2217) & (g2277)) + ((!g1031) & (!g1065) & (g3412) & (g3413) & (g2217) & (!g2277)) + ((!g1031) & (g1065) & (!g3412) & (!g3413) & (!g2217) & (!g2277)) + ((!g1031) & (g1065) & (!g3412) & (!g3413) & (g2217) & (!g2277)) + ((!g1031) & (g1065) & (!g3412) & (g3413) & (!g2217) & (!g2277)) + ((!g1031) & (g1065) & (g3412) & (!g3413) & (!g2217) & (!g2277)) + ((!g1031) & (g1065) & (g3412) & (g3413) & (!g2217) & (!g2277)) + ((g1031) & (!g1065) & (!g3412) & (!g3413) & (!g2217) & (!g2277)) + ((g1031) & (!g1065) & (!g3412) & (!g3413) & (!g2217) & (g2277)) + ((g1031) & (!g1065) & (!g3412) & (!g3413) & (g2217) & (!g2277)) + ((g1031) & (!g1065) & (!g3412) & (g3413) & (!g2217) & (!g2277)) + ((g1031) & (!g1065) & (!g3412) & (g3413) & (g2217) & (!g2277)) + ((g1031) & (!g1065) & (g3412) & (!g3413) & (!g2217) & (!g2277)) + ((g1031) & (!g1065) & (g3412) & (!g3413) & (g2217) & (!g2277)) + ((g1031) & (!g1065) & (g3412) & (g3413) & (!g2217) & (!g2277)) + ((g1031) & (!g1065) & (g3412) & (g3413) & (g2217) & (!g2277)) + ((g1031) & (g1065) & (!g3412) & (!g3413) & (!g2217) & (!g2277)));
	assign g3415 = (((!g1031) & (!g3412) & (!g3413) & (!g2217) & (!g5794) & (g5795)) + ((!g1031) & (!g3412) & (!g3413) & (g2217) & (!g5794) & (g5795)) + ((!g1031) & (!g3412) & (g3413) & (!g2217) & (!g5794) & (g5795)) + ((!g1031) & (!g3412) & (g3413) & (g2217) & (!g5794) & (g5795)) + ((!g1031) & (!g3412) & (g3413) & (g2217) & (g5794) & (g5795)) + ((!g1031) & (g3412) & (!g3413) & (!g2217) & (!g5794) & (g5795)) + ((!g1031) & (g3412) & (!g3413) & (g2217) & (!g5794) & (g5795)) + ((!g1031) & (g3412) & (!g3413) & (g2217) & (g5794) & (g5795)) + ((!g1031) & (g3412) & (g3413) & (!g2217) & (!g5794) & (g5795)) + ((!g1031) & (g3412) & (g3413) & (g2217) & (!g5794) & (g5795)) + ((!g1031) & (g3412) & (g3413) & (g2217) & (g5794) & (g5795)) + ((g1031) & (!g3412) & (!g3413) & (!g2217) & (!g5794) & (g5795)) + ((g1031) & (!g3412) & (!g3413) & (g2217) & (!g5794) & (g5795)) + ((g1031) & (!g3412) & (!g3413) & (g2217) & (g5794) & (g5795)) + ((g1031) & (!g3412) & (g3413) & (!g2217) & (!g5794) & (g5795)) + ((g1031) & (!g3412) & (g3413) & (!g2217) & (g5794) & (g5795)) + ((g1031) & (!g3412) & (g3413) & (g2217) & (!g5794) & (g5795)) + ((g1031) & (!g3412) & (g3413) & (g2217) & (g5794) & (g5795)) + ((g1031) & (g3412) & (!g3413) & (!g2217) & (!g5794) & (g5795)) + ((g1031) & (g3412) & (!g3413) & (!g2217) & (g5794) & (g5795)) + ((g1031) & (g3412) & (!g3413) & (g2217) & (!g5794) & (g5795)) + ((g1031) & (g3412) & (!g3413) & (g2217) & (g5794) & (g5795)) + ((g1031) & (g3412) & (g3413) & (!g2217) & (!g5794) & (g5795)) + ((g1031) & (g3412) & (g3413) & (!g2217) & (g5794) & (g5795)) + ((g1031) & (g3412) & (g3413) & (g2217) & (!g5794) & (g5795)) + ((g1031) & (g3412) & (g3413) & (g2217) & (g5794) & (g5795)));
	assign g3416 = (((g1165) & (g2383)));
	assign g3417 = (((!g1199) & (!g1236) & (!g3415) & (!g3416) & (!g2468) & (!g2523)) + ((!g1199) & (!g1236) & (!g3415) & (!g3416) & (!g2468) & (g2523)) + ((!g1199) & (!g1236) & (!g3415) & (!g3416) & (g2468) & (!g2523)) + ((!g1199) & (!g1236) & (!g3415) & (!g3416) & (g2468) & (g2523)) + ((!g1199) & (!g1236) & (!g3415) & (g3416) & (!g2468) & (!g2523)) + ((!g1199) & (!g1236) & (!g3415) & (g3416) & (!g2468) & (g2523)) + ((!g1199) & (!g1236) & (!g3415) & (g3416) & (g2468) & (!g2523)) + ((!g1199) & (!g1236) & (g3415) & (!g3416) & (!g2468) & (!g2523)) + ((!g1199) & (!g1236) & (g3415) & (!g3416) & (!g2468) & (g2523)) + ((!g1199) & (!g1236) & (g3415) & (!g3416) & (g2468) & (!g2523)) + ((!g1199) & (!g1236) & (g3415) & (g3416) & (!g2468) & (!g2523)) + ((!g1199) & (!g1236) & (g3415) & (g3416) & (!g2468) & (g2523)) + ((!g1199) & (!g1236) & (g3415) & (g3416) & (g2468) & (!g2523)) + ((!g1199) & (g1236) & (!g3415) & (!g3416) & (!g2468) & (!g2523)) + ((!g1199) & (g1236) & (!g3415) & (!g3416) & (g2468) & (!g2523)) + ((!g1199) & (g1236) & (!g3415) & (g3416) & (!g2468) & (!g2523)) + ((!g1199) & (g1236) & (g3415) & (!g3416) & (!g2468) & (!g2523)) + ((!g1199) & (g1236) & (g3415) & (g3416) & (!g2468) & (!g2523)) + ((g1199) & (!g1236) & (!g3415) & (!g3416) & (!g2468) & (!g2523)) + ((g1199) & (!g1236) & (!g3415) & (!g3416) & (!g2468) & (g2523)) + ((g1199) & (!g1236) & (!g3415) & (!g3416) & (g2468) & (!g2523)) + ((g1199) & (!g1236) & (!g3415) & (g3416) & (!g2468) & (!g2523)) + ((g1199) & (!g1236) & (!g3415) & (g3416) & (g2468) & (!g2523)) + ((g1199) & (!g1236) & (g3415) & (!g3416) & (!g2468) & (!g2523)) + ((g1199) & (!g1236) & (g3415) & (!g3416) & (g2468) & (!g2523)) + ((g1199) & (!g1236) & (g3415) & (g3416) & (!g2468) & (!g2523)) + ((g1199) & (!g1236) & (g3415) & (g3416) & (g2468) & (!g2523)) + ((g1199) & (g1236) & (!g3415) & (!g3416) & (!g2468) & (!g2523)));
	assign g3418 = (((!g1337) & (g2663)) + ((g1337) & (!g2663)));
	assign g3419 = (((!g1269) & (!g1303) & (!g3417) & (g2575) & (g2607) & (g3418)) + ((!g1269) & (g1303) & (!g3417) & (!g2575) & (g2607) & (g3418)) + ((!g1269) & (g1303) & (!g3417) & (g2575) & (!g2607) & (g3418)) + ((!g1269) & (g1303) & (!g3417) & (g2575) & (g2607) & (g3418)) + ((!g1269) & (g1303) & (g3417) & (!g2575) & (g2607) & (g3418)) + ((!g1269) & (g1303) & (g3417) & (g2575) & (g2607) & (g3418)) + ((g1269) & (!g1303) & (!g3417) & (!g2575) & (g2607) & (g3418)) + ((g1269) & (!g1303) & (!g3417) & (g2575) & (g2607) & (g3418)) + ((g1269) & (!g1303) & (g3417) & (g2575) & (g2607) & (g3418)) + ((g1269) & (g1303) & (!g3417) & (!g2575) & (!g2607) & (g3418)) + ((g1269) & (g1303) & (!g3417) & (!g2575) & (g2607) & (g3418)) + ((g1269) & (g1303) & (!g3417) & (g2575) & (!g2607) & (g3418)) + ((g1269) & (g1303) & (!g3417) & (g2575) & (g2607) & (g3418)) + ((g1269) & (g1303) & (g3417) & (!g2575) & (g2607) & (g3418)) + ((g1269) & (g1303) & (g3417) & (g2575) & (!g2607) & (g3418)) + ((g1269) & (g1303) & (g3417) & (g2575) & (g2607) & (g3418)));
	assign g3420 = (((g1337) & (g2663)));
	assign g3421 = (((!g1370) & (!g1406) & (!g3419) & (!g3420) & (!g2690) & (!g2774)) + ((!g1370) & (!g1406) & (!g3419) & (!g3420) & (!g2690) & (g2774)) + ((!g1370) & (!g1406) & (!g3419) & (!g3420) & (g2690) & (!g2774)) + ((!g1370) & (!g1406) & (!g3419) & (!g3420) & (g2690) & (g2774)) + ((!g1370) & (!g1406) & (!g3419) & (g3420) & (!g2690) & (!g2774)) + ((!g1370) & (!g1406) & (!g3419) & (g3420) & (!g2690) & (g2774)) + ((!g1370) & (!g1406) & (!g3419) & (g3420) & (g2690) & (!g2774)) + ((!g1370) & (!g1406) & (g3419) & (!g3420) & (!g2690) & (!g2774)) + ((!g1370) & (!g1406) & (g3419) & (!g3420) & (!g2690) & (g2774)) + ((!g1370) & (!g1406) & (g3419) & (!g3420) & (g2690) & (!g2774)) + ((!g1370) & (!g1406) & (g3419) & (g3420) & (!g2690) & (!g2774)) + ((!g1370) & (!g1406) & (g3419) & (g3420) & (!g2690) & (g2774)) + ((!g1370) & (!g1406) & (g3419) & (g3420) & (g2690) & (!g2774)) + ((!g1370) & (g1406) & (!g3419) & (!g3420) & (!g2690) & (!g2774)) + ((!g1370) & (g1406) & (!g3419) & (!g3420) & (g2690) & (!g2774)) + ((!g1370) & (g1406) & (!g3419) & (g3420) & (!g2690) & (!g2774)) + ((!g1370) & (g1406) & (g3419) & (!g3420) & (!g2690) & (!g2774)) + ((!g1370) & (g1406) & (g3419) & (g3420) & (!g2690) & (!g2774)) + ((g1370) & (!g1406) & (!g3419) & (!g3420) & (!g2690) & (!g2774)) + ((g1370) & (!g1406) & (!g3419) & (!g3420) & (!g2690) & (g2774)) + ((g1370) & (!g1406) & (!g3419) & (!g3420) & (g2690) & (!g2774)) + ((g1370) & (!g1406) & (!g3419) & (g3420) & (!g2690) & (!g2774)) + ((g1370) & (!g1406) & (!g3419) & (g3420) & (g2690) & (!g2774)) + ((g1370) & (!g1406) & (g3419) & (!g3420) & (!g2690) & (!g2774)) + ((g1370) & (!g1406) & (g3419) & (!g3420) & (g2690) & (!g2774)) + ((g1370) & (!g1406) & (g3419) & (g3420) & (!g2690) & (!g2774)) + ((g1370) & (!g1406) & (g3419) & (g3420) & (g2690) & (!g2774)) + ((g1370) & (g1406) & (!g3419) & (!g3420) & (!g2690) & (!g2774)));
	assign g3422 = (((!g1507) & (g2881)) + ((g1507) & (!g2881)));
	assign g3423 = (((!g1439) & (!g1473) & (!g3421) & (g2797) & (g2854) & (g3422)) + ((!g1439) & (g1473) & (!g3421) & (!g2797) & (g2854) & (g3422)) + ((!g1439) & (g1473) & (!g3421) & (g2797) & (!g2854) & (g3422)) + ((!g1439) & (g1473) & (!g3421) & (g2797) & (g2854) & (g3422)) + ((!g1439) & (g1473) & (g3421) & (!g2797) & (g2854) & (g3422)) + ((!g1439) & (g1473) & (g3421) & (g2797) & (g2854) & (g3422)) + ((g1439) & (!g1473) & (!g3421) & (!g2797) & (g2854) & (g3422)) + ((g1439) & (!g1473) & (!g3421) & (g2797) & (g2854) & (g3422)) + ((g1439) & (!g1473) & (g3421) & (g2797) & (g2854) & (g3422)) + ((g1439) & (g1473) & (!g3421) & (!g2797) & (!g2854) & (g3422)) + ((g1439) & (g1473) & (!g3421) & (!g2797) & (g2854) & (g3422)) + ((g1439) & (g1473) & (!g3421) & (g2797) & (!g2854) & (g3422)) + ((g1439) & (g1473) & (!g3421) & (g2797) & (g2854) & (g3422)) + ((g1439) & (g1473) & (g3421) & (!g2797) & (g2854) & (g3422)) + ((g1439) & (g1473) & (g3421) & (g2797) & (!g2854) & (g3422)) + ((g1439) & (g1473) & (g3421) & (g2797) & (g2854) & (g3422)));
	assign g3424 = (((g1507) & (g2881)));
	assign g3425 = (((!g1540) & (!g1577) & (!g3423) & (!g3424) & (!g2950) & (!g2999)) + ((!g1540) & (!g1577) & (!g3423) & (!g3424) & (!g2950) & (g2999)) + ((!g1540) & (!g1577) & (!g3423) & (!g3424) & (g2950) & (!g2999)) + ((!g1540) & (!g1577) & (!g3423) & (!g3424) & (g2950) & (g2999)) + ((!g1540) & (!g1577) & (!g3423) & (g3424) & (!g2950) & (!g2999)) + ((!g1540) & (!g1577) & (!g3423) & (g3424) & (!g2950) & (g2999)) + ((!g1540) & (!g1577) & (!g3423) & (g3424) & (g2950) & (!g2999)) + ((!g1540) & (!g1577) & (g3423) & (!g3424) & (!g2950) & (!g2999)) + ((!g1540) & (!g1577) & (g3423) & (!g3424) & (!g2950) & (g2999)) + ((!g1540) & (!g1577) & (g3423) & (!g3424) & (g2950) & (!g2999)) + ((!g1540) & (!g1577) & (g3423) & (g3424) & (!g2950) & (!g2999)) + ((!g1540) & (!g1577) & (g3423) & (g3424) & (!g2950) & (g2999)) + ((!g1540) & (!g1577) & (g3423) & (g3424) & (g2950) & (!g2999)) + ((!g1540) & (g1577) & (!g3423) & (!g3424) & (!g2950) & (!g2999)) + ((!g1540) & (g1577) & (!g3423) & (!g3424) & (g2950) & (!g2999)) + ((!g1540) & (g1577) & (!g3423) & (g3424) & (!g2950) & (!g2999)) + ((!g1540) & (g1577) & (g3423) & (!g3424) & (!g2950) & (!g2999)) + ((!g1540) & (g1577) & (g3423) & (g3424) & (!g2950) & (!g2999)) + ((g1540) & (!g1577) & (!g3423) & (!g3424) & (!g2950) & (!g2999)) + ((g1540) & (!g1577) & (!g3423) & (!g3424) & (!g2950) & (g2999)) + ((g1540) & (!g1577) & (!g3423) & (!g3424) & (g2950) & (!g2999)) + ((g1540) & (!g1577) & (!g3423) & (g3424) & (!g2950) & (!g2999)) + ((g1540) & (!g1577) & (!g3423) & (g3424) & (g2950) & (!g2999)) + ((g1540) & (!g1577) & (g3423) & (!g3424) & (!g2950) & (!g2999)) + ((g1540) & (!g1577) & (g3423) & (!g3424) & (g2950) & (!g2999)) + ((g1540) & (!g1577) & (g3423) & (g3424) & (!g2950) & (!g2999)) + ((g1540) & (!g1577) & (g3423) & (g3424) & (g2950) & (!g2999)) + ((g1540) & (g1577) & (!g3423) & (!g3424) & (!g2950) & (!g2999)));
	assign g3426 = (((!g1610) & (!g3425) & (!g3047)) + ((!g1610) & (g3425) & (g3047)) + ((g1610) & (!g3425) & (g3047)) + ((g1610) & (g3425) & (!g3047)));
	assign g8276 = (((!g5560) & (g5559) & (!g3427)) + ((!g5560) & (g5559) & (g3427)) + ((g5560) & (!g5559) & (g3427)) + ((g5560) & (g5559) & (g3427)));
	assign g3428 = (((!g830) & (!g1914) & (!g1884) & (!g3409) & (!g3426) & (g3427)) + ((!g830) & (!g1914) & (!g1884) & (!g3409) & (g3426) & (g3427)) + ((!g830) & (!g1914) & (!g1884) & (g3409) & (!g3426) & (g3427)) + ((!g830) & (!g1914) & (!g1884) & (g3409) & (g3426) & (g3427)) + ((!g830) & (!g1914) & (g1884) & (!g3409) & (!g3426) & (g3427)) + ((!g830) & (!g1914) & (g1884) & (!g3409) & (g3426) & (g3427)) + ((!g830) & (!g1914) & (g1884) & (g3409) & (!g3426) & (g3427)) + ((!g830) & (!g1914) & (g1884) & (g3409) & (g3426) & (g3427)) + ((!g830) & (g1914) & (!g1884) & (!g3409) & (!g3426) & (g3427)) + ((!g830) & (g1914) & (!g1884) & (!g3409) & (g3426) & (g3427)) + ((!g830) & (g1914) & (!g1884) & (g3409) & (!g3426) & (g3427)) + ((!g830) & (g1914) & (!g1884) & (g3409) & (g3426) & (g3427)) + ((!g830) & (g1914) & (g1884) & (!g3409) & (!g3426) & (g3427)) + ((!g830) & (g1914) & (g1884) & (!g3409) & (g3426) & (g3427)) + ((!g830) & (g1914) & (g1884) & (g3409) & (!g3426) & (g3427)) + ((!g830) & (g1914) & (g1884) & (g3409) & (g3426) & (g3427)) + ((g830) & (!g1914) & (!g1884) & (!g3409) & (g3426) & (!g3427)) + ((g830) & (!g1914) & (!g1884) & (!g3409) & (g3426) & (g3427)) + ((g830) & (!g1914) & (!g1884) & (g3409) & (g3426) & (!g3427)) + ((g830) & (!g1914) & (!g1884) & (g3409) & (g3426) & (g3427)) + ((g830) & (!g1914) & (g1884) & (!g3409) & (!g3426) & (!g3427)) + ((g830) & (!g1914) & (g1884) & (!g3409) & (!g3426) & (g3427)) + ((g830) & (!g1914) & (g1884) & (g3409) & (!g3426) & (!g3427)) + ((g830) & (!g1914) & (g1884) & (g3409) & (!g3426) & (g3427)) + ((g830) & (g1914) & (!g1884) & (g3409) & (!g3426) & (!g3427)) + ((g830) & (g1914) & (!g1884) & (g3409) & (!g3426) & (g3427)) + ((g830) & (g1914) & (!g1884) & (g3409) & (g3426) & (!g3427)) + ((g830) & (g1914) & (!g1884) & (g3409) & (g3426) & (g3427)) + ((g830) & (g1914) & (g1884) & (!g3409) & (!g3426) & (!g3427)) + ((g830) & (g1914) & (g1884) & (!g3409) & (!g3426) & (g3427)) + ((g830) & (g1914) & (g1884) & (!g3409) & (g3426) & (!g3427)) + ((g830) & (g1914) & (g1884) & (!g3409) & (g3426) & (g3427)));
	assign g3429 = (((!reset) & (!g830) & (!g1921) & (!g1922) & (!g2016)) + ((!reset) & (!g830) & (!g1921) & (g1922) & (!g2016)) + ((!reset) & (!g830) & (g1921) & (!g1922) & (!g2016)) + ((!reset) & (!g830) & (g1921) & (g1922) & (!g2016)) + ((!reset) & (g830) & (!g1921) & (!g1922) & (!g2016)) + ((!reset) & (g830) & (!g1921) & (!g1922) & (g2016)) + ((!reset) & (g830) & (!g1921) & (g1922) & (!g2016)) + ((!reset) & (g830) & (!g1921) & (g1922) & (g2016)) + ((!reset) & (g830) & (g1921) & (!g1922) & (!g2016)) + ((!reset) & (g830) & (g1921) & (g1922) & (!g2016)) + ((!reset) & (g830) & (g1921) & (g1922) & (g2016)) + ((reset) & (!g830) & (!g1921) & (!g1922) & (!g2016)) + ((reset) & (!g830) & (!g1921) & (!g1922) & (g2016)) + ((reset) & (!g830) & (!g1921) & (g1922) & (!g2016)) + ((reset) & (!g830) & (!g1921) & (g1922) & (g2016)) + ((reset) & (!g830) & (g1921) & (!g1922) & (!g2016)) + ((reset) & (!g830) & (g1921) & (!g1922) & (g2016)) + ((reset) & (!g830) & (g1921) & (g1922) & (!g2016)) + ((reset) & (!g830) & (g1921) & (g1922) & (g2016)) + ((reset) & (g830) & (!g1921) & (!g1922) & (!g2016)) + ((reset) & (g830) & (!g1921) & (!g1922) & (g2016)) + ((reset) & (g830) & (!g1921) & (g1922) & (!g2016)) + ((reset) & (g830) & (!g1921) & (g1922) & (g2016)) + ((reset) & (g830) & (g1921) & (!g1922) & (!g2016)) + ((reset) & (g830) & (g1921) & (!g1922) & (g2016)) + ((reset) & (g830) & (g1921) & (g1922) & (!g2016)) + ((reset) & (g830) & (g1921) & (g1922) & (g2016)));
	assign g3430 = (((!g1894) & (!g1910) & (!g2034) & (!g2038) & (g2065) & (g2088)) + ((!g1894) & (!g1910) & (!g2034) & (g2038) & (g2065) & (g2088)) + ((!g1894) & (!g1910) & (g2034) & (!g2038) & (g2065) & (g2088)) + ((!g1894) & (!g1910) & (g2034) & (g2038) & (!g2065) & (g2088)) + ((!g1894) & (!g1910) & (g2034) & (g2038) & (g2065) & (!g2088)) + ((!g1894) & (!g1910) & (g2034) & (g2038) & (g2065) & (g2088)) + ((!g1894) & (g1910) & (!g2034) & (!g2038) & (g2065) & (g2088)) + ((!g1894) & (g1910) & (!g2034) & (g2038) & (g2065) & (g2088)) + ((!g1894) & (g1910) & (g2034) & (!g2038) & (g2065) & (g2088)) + ((!g1894) & (g1910) & (g2034) & (g2038) & (!g2065) & (g2088)) + ((!g1894) & (g1910) & (g2034) & (g2038) & (g2065) & (!g2088)) + ((!g1894) & (g1910) & (g2034) & (g2038) & (g2065) & (g2088)) + ((g1894) & (!g1910) & (!g2034) & (!g2038) & (g2065) & (g2088)) + ((g1894) & (!g1910) & (!g2034) & (g2038) & (g2065) & (g2088)) + ((g1894) & (!g1910) & (g2034) & (!g2038) & (g2065) & (g2088)) + ((g1894) & (!g1910) & (g2034) & (g2038) & (!g2065) & (g2088)) + ((g1894) & (!g1910) & (g2034) & (g2038) & (g2065) & (!g2088)) + ((g1894) & (!g1910) & (g2034) & (g2038) & (g2065) & (g2088)) + ((g1894) & (g1910) & (!g2034) & (!g2038) & (g2065) & (g2088)) + ((g1894) & (g1910) & (!g2034) & (g2038) & (!g2065) & (g2088)) + ((g1894) & (g1910) & (!g2034) & (g2038) & (g2065) & (!g2088)) + ((g1894) & (g1910) & (!g2034) & (g2038) & (g2065) & (g2088)) + ((g1894) & (g1910) & (g2034) & (!g2038) & (!g2065) & (g2088)) + ((g1894) & (g1910) & (g2034) & (!g2038) & (g2065) & (!g2088)) + ((g1894) & (g1910) & (g2034) & (!g2038) & (g2065) & (g2088)) + ((g1894) & (g1910) & (g2034) & (g2038) & (!g2065) & (g2088)) + ((g1894) & (g1910) & (g2034) & (g2038) & (g2065) & (!g2088)) + ((g1894) & (g1910) & (g2034) & (g2038) & (g2065) & (g2088)));
	assign g3431 = (((!g2196) & (g2200)) + ((g2196) & (!g2200)));
	assign g3432 = (((!g3430) & (!g2116) & (!g2120) & (g2147) & (g2170) & (g3431)) + ((!g3430) & (!g2116) & (g2120) & (g2147) & (g2170) & (g3431)) + ((!g3430) & (g2116) & (!g2120) & (g2147) & (g2170) & (g3431)) + ((!g3430) & (g2116) & (g2120) & (!g2147) & (g2170) & (g3431)) + ((!g3430) & (g2116) & (g2120) & (g2147) & (!g2170) & (g3431)) + ((!g3430) & (g2116) & (g2120) & (g2147) & (g2170) & (g3431)) + ((g3430) & (!g2116) & (!g2120) & (g2147) & (g2170) & (g3431)) + ((g3430) & (!g2116) & (g2120) & (!g2147) & (g2170) & (g3431)) + ((g3430) & (!g2116) & (g2120) & (g2147) & (!g2170) & (g3431)) + ((g3430) & (!g2116) & (g2120) & (g2147) & (g2170) & (g3431)) + ((g3430) & (g2116) & (!g2120) & (!g2147) & (g2170) & (g3431)) + ((g3430) & (g2116) & (!g2120) & (g2147) & (!g2170) & (g3431)) + ((g3430) & (g2116) & (!g2120) & (g2147) & (g2170) & (g3431)) + ((g3430) & (g2116) & (g2120) & (!g2147) & (g2170) & (g3431)) + ((g3430) & (g2116) & (g2120) & (g2147) & (!g2170) & (g3431)) + ((g3430) & (g2116) & (g2120) & (g2147) & (g2170) & (g3431)));
	assign g3433 = (((g2196) & (g2200)));
	assign g3434 = (((!g3432) & (!g3433) & (!g2227) & (!g2250) & (!g2279) & (!g2283)) + ((!g3432) & (!g3433) & (!g2227) & (!g2250) & (!g2279) & (g2283)) + ((!g3432) & (!g3433) & (!g2227) & (!g2250) & (g2279) & (!g2283)) + ((!g3432) & (!g3433) & (!g2227) & (g2250) & (!g2279) & (!g2283)) + ((!g3432) & (!g3433) & (!g2227) & (g2250) & (!g2279) & (g2283)) + ((!g3432) & (!g3433) & (!g2227) & (g2250) & (g2279) & (!g2283)) + ((!g3432) & (!g3433) & (g2227) & (!g2250) & (!g2279) & (!g2283)) + ((!g3432) & (!g3433) & (g2227) & (!g2250) & (!g2279) & (g2283)) + ((!g3432) & (!g3433) & (g2227) & (!g2250) & (g2279) & (!g2283)) + ((!g3432) & (!g3433) & (g2227) & (g2250) & (!g2279) & (!g2283)) + ((!g3432) & (g3433) & (!g2227) & (!g2250) & (!g2279) & (!g2283)) + ((!g3432) & (g3433) & (!g2227) & (!g2250) & (!g2279) & (g2283)) + ((!g3432) & (g3433) & (!g2227) & (!g2250) & (g2279) & (!g2283)) + ((!g3432) & (g3433) & (!g2227) & (g2250) & (!g2279) & (!g2283)) + ((!g3432) & (g3433) & (g2227) & (!g2250) & (!g2279) & (!g2283)) + ((!g3432) & (g3433) & (g2227) & (g2250) & (!g2279) & (!g2283)) + ((g3432) & (!g3433) & (!g2227) & (!g2250) & (!g2279) & (!g2283)) + ((g3432) & (!g3433) & (!g2227) & (!g2250) & (!g2279) & (g2283)) + ((g3432) & (!g3433) & (!g2227) & (!g2250) & (g2279) & (!g2283)) + ((g3432) & (!g3433) & (!g2227) & (g2250) & (!g2279) & (!g2283)) + ((g3432) & (!g3433) & (g2227) & (!g2250) & (!g2279) & (!g2283)) + ((g3432) & (!g3433) & (g2227) & (g2250) & (!g2279) & (!g2283)) + ((g3432) & (g3433) & (!g2227) & (!g2250) & (!g2279) & (!g2283)) + ((g3432) & (g3433) & (!g2227) & (!g2250) & (!g2279) & (g2283)) + ((g3432) & (g3433) & (!g2227) & (!g2250) & (g2279) & (!g2283)) + ((g3432) & (g3433) & (!g2227) & (g2250) & (!g2279) & (!g2283)) + ((g3432) & (g3433) & (g2227) & (!g2250) & (!g2279) & (!g2283)) + ((g3432) & (g3433) & (g2227) & (g2250) & (!g2279) & (!g2283)));
	assign g3435 = (((!g2393) & (g2416)) + ((g2393) & (!g2416)));
	assign g3436 = (((!g3434) & (!g2314) & (!g2337) & (g2362) & (g2366) & (g3435)) + ((!g3434) & (!g2314) & (g2337) & (!g2362) & (g2366) & (g3435)) + ((!g3434) & (!g2314) & (g2337) & (g2362) & (!g2366) & (g3435)) + ((!g3434) & (!g2314) & (g2337) & (g2362) & (g2366) & (g3435)) + ((!g3434) & (g2314) & (!g2337) & (!g2362) & (g2366) & (g3435)) + ((!g3434) & (g2314) & (!g2337) & (g2362) & (!g2366) & (g3435)) + ((!g3434) & (g2314) & (!g2337) & (g2362) & (g2366) & (g3435)) + ((!g3434) & (g2314) & (g2337) & (!g2362) & (g2366) & (g3435)) + ((!g3434) & (g2314) & (g2337) & (g2362) & (!g2366) & (g3435)) + ((!g3434) & (g2314) & (g2337) & (g2362) & (g2366) & (g3435)) + ((g3434) & (!g2314) & (!g2337) & (g2362) & (g2366) & (g3435)) + ((g3434) & (!g2314) & (g2337) & (g2362) & (g2366) & (g3435)) + ((g3434) & (g2314) & (!g2337) & (g2362) & (g2366) & (g3435)) + ((g3434) & (g2314) & (g2337) & (!g2362) & (g2366) & (g3435)) + ((g3434) & (g2314) & (g2337) & (g2362) & (!g2366) & (g3435)) + ((g3434) & (g2314) & (g2337) & (g2362) & (g2366) & (g3435)));
	assign g3437 = (((g2393) & (g2416)));
	assign g3438 = (((!g3436) & (!g3437) & (!g2474) & (!g2486) & (!g2529) & (!g2544)) + ((!g3436) & (!g3437) & (!g2474) & (!g2486) & (!g2529) & (g2544)) + ((!g3436) & (!g3437) & (!g2474) & (!g2486) & (g2529) & (!g2544)) + ((!g3436) & (!g3437) & (!g2474) & (g2486) & (!g2529) & (!g2544)) + ((!g3436) & (!g3437) & (!g2474) & (g2486) & (!g2529) & (g2544)) + ((!g3436) & (!g3437) & (!g2474) & (g2486) & (g2529) & (!g2544)) + ((!g3436) & (!g3437) & (g2474) & (!g2486) & (!g2529) & (!g2544)) + ((!g3436) & (!g3437) & (g2474) & (!g2486) & (!g2529) & (g2544)) + ((!g3436) & (!g3437) & (g2474) & (!g2486) & (g2529) & (!g2544)) + ((!g3436) & (!g3437) & (g2474) & (g2486) & (!g2529) & (!g2544)) + ((!g3436) & (g3437) & (!g2474) & (!g2486) & (!g2529) & (!g2544)) + ((!g3436) & (g3437) & (!g2474) & (!g2486) & (!g2529) & (g2544)) + ((!g3436) & (g3437) & (!g2474) & (!g2486) & (g2529) & (!g2544)) + ((!g3436) & (g3437) & (!g2474) & (g2486) & (!g2529) & (!g2544)) + ((!g3436) & (g3437) & (g2474) & (!g2486) & (!g2529) & (!g2544)) + ((!g3436) & (g3437) & (g2474) & (g2486) & (!g2529) & (!g2544)) + ((g3436) & (!g3437) & (!g2474) & (!g2486) & (!g2529) & (!g2544)) + ((g3436) & (!g3437) & (!g2474) & (!g2486) & (!g2529) & (g2544)) + ((g3436) & (!g3437) & (!g2474) & (!g2486) & (g2529) & (!g2544)) + ((g3436) & (!g3437) & (!g2474) & (g2486) & (!g2529) & (!g2544)) + ((g3436) & (!g3437) & (g2474) & (!g2486) & (!g2529) & (!g2544)) + ((g3436) & (!g3437) & (g2474) & (g2486) & (!g2529) & (!g2544)) + ((g3436) & (g3437) & (!g2474) & (!g2486) & (!g2529) & (!g2544)) + ((g3436) & (g3437) & (!g2474) & (!g2486) & (!g2529) & (g2544)) + ((g3436) & (g3437) & (!g2474) & (!g2486) & (g2529) & (!g2544)) + ((g3436) & (g3437) & (!g2474) & (g2486) & (!g2529) & (!g2544)) + ((g3436) & (g3437) & (g2474) & (!g2486) & (!g2529) & (!g2544)) + ((g3436) & (g3437) & (g2474) & (g2486) & (!g2529) & (!g2544)));
	assign g3439 = (((!g2665) & (g2669)) + ((g2665) & (!g2669)));
	assign g3440 = (((!g3438) & (!g2578) & (!g2584) & (g2617) & (g2640) & (g3439)) + ((!g3438) & (!g2578) & (g2584) & (!g2617) & (g2640) & (g3439)) + ((!g3438) & (!g2578) & (g2584) & (g2617) & (!g2640) & (g3439)) + ((!g3438) & (!g2578) & (g2584) & (g2617) & (g2640) & (g3439)) + ((!g3438) & (g2578) & (!g2584) & (!g2617) & (g2640) & (g3439)) + ((!g3438) & (g2578) & (!g2584) & (g2617) & (!g2640) & (g3439)) + ((!g3438) & (g2578) & (!g2584) & (g2617) & (g2640) & (g3439)) + ((!g3438) & (g2578) & (g2584) & (!g2617) & (g2640) & (g3439)) + ((!g3438) & (g2578) & (g2584) & (g2617) & (!g2640) & (g3439)) + ((!g3438) & (g2578) & (g2584) & (g2617) & (g2640) & (g3439)) + ((g3438) & (!g2578) & (!g2584) & (g2617) & (g2640) & (g3439)) + ((g3438) & (!g2578) & (g2584) & (g2617) & (g2640) & (g3439)) + ((g3438) & (g2578) & (!g2584) & (g2617) & (g2640) & (g3439)) + ((g3438) & (g2578) & (g2584) & (!g2617) & (g2640) & (g3439)) + ((g3438) & (g2578) & (g2584) & (g2617) & (!g2640) & (g3439)) + ((g3438) & (g2578) & (g2584) & (g2617) & (g2640) & (g3439)));
	assign g3441 = (((g2665) & (g2669)));
	assign g3442 = (((!g3440) & (!g3441) & (!g2708) & (!g2747) & (!g2776) & (!g2780)) + ((!g3440) & (!g3441) & (!g2708) & (!g2747) & (!g2776) & (g2780)) + ((!g3440) & (!g3441) & (!g2708) & (!g2747) & (g2776) & (!g2780)) + ((!g3440) & (!g3441) & (!g2708) & (g2747) & (!g2776) & (!g2780)) + ((!g3440) & (!g3441) & (!g2708) & (g2747) & (!g2776) & (g2780)) + ((!g3440) & (!g3441) & (!g2708) & (g2747) & (g2776) & (!g2780)) + ((!g3440) & (!g3441) & (g2708) & (!g2747) & (!g2776) & (!g2780)) + ((!g3440) & (!g3441) & (g2708) & (!g2747) & (!g2776) & (g2780)) + ((!g3440) & (!g3441) & (g2708) & (!g2747) & (g2776) & (!g2780)) + ((!g3440) & (!g3441) & (g2708) & (g2747) & (!g2776) & (!g2780)) + ((!g3440) & (g3441) & (!g2708) & (!g2747) & (!g2776) & (!g2780)) + ((!g3440) & (g3441) & (!g2708) & (!g2747) & (!g2776) & (g2780)) + ((!g3440) & (g3441) & (!g2708) & (!g2747) & (g2776) & (!g2780)) + ((!g3440) & (g3441) & (!g2708) & (g2747) & (!g2776) & (!g2780)) + ((!g3440) & (g3441) & (g2708) & (!g2747) & (!g2776) & (!g2780)) + ((!g3440) & (g3441) & (g2708) & (g2747) & (!g2776) & (!g2780)) + ((g3440) & (!g3441) & (!g2708) & (!g2747) & (!g2776) & (!g2780)) + ((g3440) & (!g3441) & (!g2708) & (!g2747) & (!g2776) & (g2780)) + ((g3440) & (!g3441) & (!g2708) & (!g2747) & (g2776) & (!g2780)) + ((g3440) & (!g3441) & (!g2708) & (g2747) & (!g2776) & (!g2780)) + ((g3440) & (!g3441) & (g2708) & (!g2747) & (!g2776) & (!g2780)) + ((g3440) & (!g3441) & (g2708) & (g2747) & (!g2776) & (!g2780)) + ((g3440) & (g3441) & (!g2708) & (!g2747) & (!g2776) & (!g2780)) + ((g3440) & (g3441) & (!g2708) & (!g2747) & (!g2776) & (g2780)) + ((g3440) & (g3441) & (!g2708) & (!g2747) & (g2776) & (!g2780)) + ((g3440) & (g3441) & (!g2708) & (g2747) & (!g2776) & (!g2780)) + ((g3440) & (g3441) & (g2708) & (!g2747) & (!g2776) & (!g2780)) + ((g3440) & (g3441) & (g2708) & (g2747) & (!g2776) & (!g2780)));
	assign g3443 = (((!g3442) & (!g2807) & (g2830)) + ((!g3442) & (g2807) & (!g2830)) + ((!g3442) & (g2807) & (g2830)) + ((g3442) & (g2807) & (g2830)));
	assign g3444 = (((!g1888) & (!g1978) & (g1980) & (!g828) & (!g864) & (g897)) + ((!g1888) & (!g1978) & (g1980) & (!g828) & (g864) & (g897)) + ((!g1888) & (!g1978) & (g1980) & (g828) & (!g864) & (g897)) + ((!g1888) & (!g1978) & (g1980) & (g828) & (g864) & (g897)) + ((!g1888) & (g1978) & (!g1980) & (!g828) & (g864) & (g897)) + ((!g1888) & (g1978) & (!g1980) & (g828) & (g864) & (g897)) + ((!g1888) & (g1978) & (g1980) & (!g828) & (!g864) & (g897)) + ((!g1888) & (g1978) & (g1980) & (!g828) & (g864) & (!g897)) + ((!g1888) & (g1978) & (g1980) & (!g828) & (g864) & (g897)) + ((!g1888) & (g1978) & (g1980) & (g828) & (!g864) & (g897)) + ((!g1888) & (g1978) & (g1980) & (g828) & (g864) & (!g897)) + ((!g1888) & (g1978) & (g1980) & (g828) & (g864) & (g897)) + ((g1888) & (!g1978) & (!g1980) & (g828) & (g864) & (g897)) + ((g1888) & (!g1978) & (g1980) & (!g828) & (!g864) & (g897)) + ((g1888) & (!g1978) & (g1980) & (!g828) & (g864) & (g897)) + ((g1888) & (!g1978) & (g1980) & (g828) & (!g864) & (g897)) + ((g1888) & (!g1978) & (g1980) & (g828) & (g864) & (!g897)) + ((g1888) & (!g1978) & (g1980) & (g828) & (g864) & (g897)) + ((g1888) & (g1978) & (!g1980) & (!g828) & (g864) & (g897)) + ((g1888) & (g1978) & (!g1980) & (g828) & (!g864) & (g897)) + ((g1888) & (g1978) & (!g1980) & (g828) & (g864) & (g897)) + ((g1888) & (g1978) & (g1980) & (!g828) & (!g864) & (g897)) + ((g1888) & (g1978) & (g1980) & (!g828) & (g864) & (!g897)) + ((g1888) & (g1978) & (g1980) & (!g828) & (g864) & (g897)) + ((g1888) & (g1978) & (g1980) & (g828) & (!g864) & (!g897)) + ((g1888) & (g1978) & (g1980) & (g828) & (!g864) & (g897)) + ((g1888) & (g1978) & (g1980) & (g828) & (g864) & (!g897)) + ((g1888) & (g1978) & (g1980) & (g828) & (g864) & (g897)));
	assign g3445 = (((!g1987) & (g998)) + ((g1987) & (!g998)));
	assign g3446 = (((!g1983) & (!g1985) & (g931) & (g964) & (g3444) & (g3445)) + ((!g1983) & (g1985) & (!g931) & (g964) & (!g3444) & (g3445)) + ((!g1983) & (g1985) & (!g931) & (g964) & (g3444) & (g3445)) + ((!g1983) & (g1985) & (g931) & (!g964) & (g3444) & (g3445)) + ((!g1983) & (g1985) & (g931) & (g964) & (!g3444) & (g3445)) + ((!g1983) & (g1985) & (g931) & (g964) & (g3444) & (g3445)) + ((g1983) & (!g1985) & (!g931) & (g964) & (g3444) & (g3445)) + ((g1983) & (!g1985) & (g931) & (g964) & (!g3444) & (g3445)) + ((g1983) & (!g1985) & (g931) & (g964) & (g3444) & (g3445)) + ((g1983) & (g1985) & (!g931) & (!g964) & (g3444) & (g3445)) + ((g1983) & (g1985) & (!g931) & (g964) & (!g3444) & (g3445)) + ((g1983) & (g1985) & (!g931) & (g964) & (g3444) & (g3445)) + ((g1983) & (g1985) & (g931) & (!g964) & (!g3444) & (g3445)) + ((g1983) & (g1985) & (g931) & (!g964) & (g3444) & (g3445)) + ((g1983) & (g1985) & (g931) & (g964) & (!g3444) & (g3445)) + ((g1983) & (g1985) & (g931) & (g964) & (g3444) & (g3445)));
	assign g3447 = (((g1987) & (g998)));
	assign g3448 = (((!g1992) & (!g1994) & (!g1031) & (!g1065) & (!g3446) & (!g3447)) + ((!g1992) & (!g1994) & (!g1031) & (!g1065) & (!g3446) & (g3447)) + ((!g1992) & (!g1994) & (!g1031) & (!g1065) & (g3446) & (!g3447)) + ((!g1992) & (!g1994) & (!g1031) & (!g1065) & (g3446) & (g3447)) + ((!g1992) & (!g1994) & (!g1031) & (g1065) & (!g3446) & (!g3447)) + ((!g1992) & (!g1994) & (!g1031) & (g1065) & (!g3446) & (g3447)) + ((!g1992) & (!g1994) & (!g1031) & (g1065) & (g3446) & (!g3447)) + ((!g1992) & (!g1994) & (!g1031) & (g1065) & (g3446) & (g3447)) + ((!g1992) & (!g1994) & (g1031) & (!g1065) & (!g3446) & (!g3447)) + ((!g1992) & (!g1994) & (g1031) & (!g1065) & (!g3446) & (g3447)) + ((!g1992) & (!g1994) & (g1031) & (!g1065) & (g3446) & (!g3447)) + ((!g1992) & (!g1994) & (g1031) & (!g1065) & (g3446) & (g3447)) + ((!g1992) & (!g1994) & (g1031) & (g1065) & (!g3446) & (!g3447)) + ((!g1992) & (g1994) & (!g1031) & (!g1065) & (!g3446) & (!g3447)) + ((!g1992) & (g1994) & (!g1031) & (!g1065) & (!g3446) & (g3447)) + ((!g1992) & (g1994) & (!g1031) & (!g1065) & (g3446) & (!g3447)) + ((!g1992) & (g1994) & (!g1031) & (!g1065) & (g3446) & (g3447)) + ((!g1992) & (g1994) & (g1031) & (!g1065) & (!g3446) & (!g3447)) + ((g1992) & (!g1994) & (!g1031) & (!g1065) & (!g3446) & (!g3447)) + ((g1992) & (!g1994) & (!g1031) & (!g1065) & (!g3446) & (g3447)) + ((g1992) & (!g1994) & (!g1031) & (!g1065) & (g3446) & (!g3447)) + ((g1992) & (!g1994) & (!g1031) & (!g1065) & (g3446) & (g3447)) + ((g1992) & (!g1994) & (!g1031) & (g1065) & (!g3446) & (!g3447)) + ((g1992) & (!g1994) & (g1031) & (!g1065) & (!g3446) & (!g3447)) + ((g1992) & (!g1994) & (g1031) & (!g1065) & (!g3446) & (g3447)) + ((g1992) & (!g1994) & (g1031) & (!g1065) & (g3446) & (!g3447)) + ((g1992) & (!g1994) & (g1031) & (!g1065) & (g3446) & (g3447)) + ((g1992) & (g1994) & (!g1031) & (!g1065) & (!g3446) & (!g3447)));
	assign g3449 = (((!g2002) & (g1165)) + ((g2002) & (!g1165)));
	assign g3450 = (((!g1997) & (!g1999) & (g1098) & (g1132) & (!g3448) & (g3449)) + ((!g1997) & (g1999) & (!g1098) & (g1132) & (!g3448) & (g3449)) + ((!g1997) & (g1999) & (!g1098) & (g1132) & (g3448) & (g3449)) + ((!g1997) & (g1999) & (g1098) & (!g1132) & (!g3448) & (g3449)) + ((!g1997) & (g1999) & (g1098) & (g1132) & (!g3448) & (g3449)) + ((!g1997) & (g1999) & (g1098) & (g1132) & (g3448) & (g3449)) + ((g1997) & (!g1999) & (!g1098) & (g1132) & (!g3448) & (g3449)) + ((g1997) & (!g1999) & (g1098) & (g1132) & (!g3448) & (g3449)) + ((g1997) & (!g1999) & (g1098) & (g1132) & (g3448) & (g3449)) + ((g1997) & (g1999) & (!g1098) & (!g1132) & (!g3448) & (g3449)) + ((g1997) & (g1999) & (!g1098) & (g1132) & (!g3448) & (g3449)) + ((g1997) & (g1999) & (!g1098) & (g1132) & (g3448) & (g3449)) + ((g1997) & (g1999) & (g1098) & (!g1132) & (!g3448) & (g3449)) + ((g1997) & (g1999) & (g1098) & (!g1132) & (g3448) & (g3449)) + ((g1997) & (g1999) & (g1098) & (g1132) & (!g3448) & (g3449)) + ((g1997) & (g1999) & (g1098) & (g1132) & (g3448) & (g3449)));
	assign g3451 = (((g2002) & (g1165)));
	assign g3452 = (((!g2004) & (!g2006) & (!g1199) & (!g1236) & (!g3450) & (!g3451)) + ((!g2004) & (!g2006) & (!g1199) & (!g1236) & (!g3450) & (g3451)) + ((!g2004) & (!g2006) & (!g1199) & (!g1236) & (g3450) & (!g3451)) + ((!g2004) & (!g2006) & (!g1199) & (!g1236) & (g3450) & (g3451)) + ((!g2004) & (!g2006) & (!g1199) & (g1236) & (!g3450) & (!g3451)) + ((!g2004) & (!g2006) & (!g1199) & (g1236) & (!g3450) & (g3451)) + ((!g2004) & (!g2006) & (!g1199) & (g1236) & (g3450) & (!g3451)) + ((!g2004) & (!g2006) & (!g1199) & (g1236) & (g3450) & (g3451)) + ((!g2004) & (!g2006) & (g1199) & (!g1236) & (!g3450) & (!g3451)) + ((!g2004) & (!g2006) & (g1199) & (!g1236) & (!g3450) & (g3451)) + ((!g2004) & (!g2006) & (g1199) & (!g1236) & (g3450) & (!g3451)) + ((!g2004) & (!g2006) & (g1199) & (!g1236) & (g3450) & (g3451)) + ((!g2004) & (!g2006) & (g1199) & (g1236) & (!g3450) & (!g3451)) + ((!g2004) & (g2006) & (!g1199) & (!g1236) & (!g3450) & (!g3451)) + ((!g2004) & (g2006) & (!g1199) & (!g1236) & (!g3450) & (g3451)) + ((!g2004) & (g2006) & (!g1199) & (!g1236) & (g3450) & (!g3451)) + ((!g2004) & (g2006) & (!g1199) & (!g1236) & (g3450) & (g3451)) + ((!g2004) & (g2006) & (g1199) & (!g1236) & (!g3450) & (!g3451)) + ((g2004) & (!g2006) & (!g1199) & (!g1236) & (!g3450) & (!g3451)) + ((g2004) & (!g2006) & (!g1199) & (!g1236) & (!g3450) & (g3451)) + ((g2004) & (!g2006) & (!g1199) & (!g1236) & (g3450) & (!g3451)) + ((g2004) & (!g2006) & (!g1199) & (!g1236) & (g3450) & (g3451)) + ((g2004) & (!g2006) & (!g1199) & (g1236) & (!g3450) & (!g3451)) + ((g2004) & (!g2006) & (g1199) & (!g1236) & (!g3450) & (!g3451)) + ((g2004) & (!g2006) & (g1199) & (!g1236) & (!g3450) & (g3451)) + ((g2004) & (!g2006) & (g1199) & (!g1236) & (g3450) & (!g3451)) + ((g2004) & (!g2006) & (g1199) & (!g1236) & (g3450) & (g3451)) + ((g2004) & (g2006) & (!g1199) & (!g1236) & (!g3450) & (!g3451)));
	assign g3453 = (((!g2004) & (!g1199) & (!g3450) & (!g3451) & (!g5797) & (g5798)) + ((!g2004) & (!g1199) & (!g3450) & (g3451) & (!g5797) & (g5798)) + ((!g2004) & (!g1199) & (g3450) & (!g3451) & (!g5797) & (g5798)) + ((!g2004) & (!g1199) & (g3450) & (g3451) & (!g5797) & (g5798)) + ((!g2004) & (g1199) & (!g3450) & (!g3451) & (!g5797) & (g5798)) + ((!g2004) & (g1199) & (!g3450) & (g3451) & (!g5797) & (g5798)) + ((!g2004) & (g1199) & (!g3450) & (g3451) & (g5797) & (g5798)) + ((!g2004) & (g1199) & (g3450) & (!g3451) & (!g5797) & (g5798)) + ((!g2004) & (g1199) & (g3450) & (!g3451) & (g5797) & (g5798)) + ((!g2004) & (g1199) & (g3450) & (g3451) & (!g5797) & (g5798)) + ((!g2004) & (g1199) & (g3450) & (g3451) & (g5797) & (g5798)) + ((g2004) & (!g1199) & (!g3450) & (!g3451) & (!g5797) & (g5798)) + ((g2004) & (!g1199) & (!g3450) & (g3451) & (!g5797) & (g5798)) + ((g2004) & (!g1199) & (!g3450) & (g3451) & (g5797) & (g5798)) + ((g2004) & (!g1199) & (g3450) & (!g3451) & (!g5797) & (g5798)) + ((g2004) & (!g1199) & (g3450) & (!g3451) & (g5797) & (g5798)) + ((g2004) & (!g1199) & (g3450) & (g3451) & (!g5797) & (g5798)) + ((g2004) & (!g1199) & (g3450) & (g3451) & (g5797) & (g5798)) + ((g2004) & (g1199) & (!g3450) & (!g3451) & (!g5797) & (g5798)) + ((g2004) & (g1199) & (!g3450) & (!g3451) & (g5797) & (g5798)) + ((g2004) & (g1199) & (!g3450) & (g3451) & (!g5797) & (g5798)) + ((g2004) & (g1199) & (!g3450) & (g3451) & (g5797) & (g5798)) + ((g2004) & (g1199) & (g3450) & (!g3451) & (!g5797) & (g5798)) + ((g2004) & (g1199) & (g3450) & (!g3451) & (g5797) & (g5798)) + ((g2004) & (g1199) & (g3450) & (g3451) & (!g5797) & (g5798)) + ((g2004) & (g1199) & (g3450) & (g3451) & (g5797) & (g5798)));
	assign g3454 = (((g2052) & (g1337)));
	assign g3455 = (((!g2101) & (!g2134) & (!g1370) & (!g1406) & (!g3453) & (!g3454)) + ((!g2101) & (!g2134) & (!g1370) & (!g1406) & (!g3453) & (g3454)) + ((!g2101) & (!g2134) & (!g1370) & (!g1406) & (g3453) & (!g3454)) + ((!g2101) & (!g2134) & (!g1370) & (!g1406) & (g3453) & (g3454)) + ((!g2101) & (!g2134) & (!g1370) & (g1406) & (!g3453) & (!g3454)) + ((!g2101) & (!g2134) & (!g1370) & (g1406) & (!g3453) & (g3454)) + ((!g2101) & (!g2134) & (!g1370) & (g1406) & (g3453) & (!g3454)) + ((!g2101) & (!g2134) & (!g1370) & (g1406) & (g3453) & (g3454)) + ((!g2101) & (!g2134) & (g1370) & (!g1406) & (!g3453) & (!g3454)) + ((!g2101) & (!g2134) & (g1370) & (!g1406) & (!g3453) & (g3454)) + ((!g2101) & (!g2134) & (g1370) & (!g1406) & (g3453) & (!g3454)) + ((!g2101) & (!g2134) & (g1370) & (!g1406) & (g3453) & (g3454)) + ((!g2101) & (!g2134) & (g1370) & (g1406) & (!g3453) & (!g3454)) + ((!g2101) & (g2134) & (!g1370) & (!g1406) & (!g3453) & (!g3454)) + ((!g2101) & (g2134) & (!g1370) & (!g1406) & (!g3453) & (g3454)) + ((!g2101) & (g2134) & (!g1370) & (!g1406) & (g3453) & (!g3454)) + ((!g2101) & (g2134) & (!g1370) & (!g1406) & (g3453) & (g3454)) + ((!g2101) & (g2134) & (g1370) & (!g1406) & (!g3453) & (!g3454)) + ((g2101) & (!g2134) & (!g1370) & (!g1406) & (!g3453) & (!g3454)) + ((g2101) & (!g2134) & (!g1370) & (!g1406) & (!g3453) & (g3454)) + ((g2101) & (!g2134) & (!g1370) & (!g1406) & (g3453) & (!g3454)) + ((g2101) & (!g2134) & (!g1370) & (!g1406) & (g3453) & (g3454)) + ((g2101) & (!g2134) & (!g1370) & (g1406) & (!g3453) & (!g3454)) + ((g2101) & (!g2134) & (g1370) & (!g1406) & (!g3453) & (!g3454)) + ((g2101) & (!g2134) & (g1370) & (!g1406) & (!g3453) & (g3454)) + ((g2101) & (!g2134) & (g1370) & (!g1406) & (g3453) & (!g3454)) + ((g2101) & (!g2134) & (g1370) & (!g1406) & (g3453) & (g3454)) + ((g2101) & (g2134) & (!g1370) & (!g1406) & (!g3453) & (!g3454)));
	assign g3456 = (((!g2263) & (g1507)) + ((g2263) & (!g1507)));
	assign g3457 = (((!g2181) & (!g2213) & (g1439) & (g1473) & (!g3455) & (g3456)) + ((!g2181) & (g2213) & (!g1439) & (g1473) & (!g3455) & (g3456)) + ((!g2181) & (g2213) & (!g1439) & (g1473) & (g3455) & (g3456)) + ((!g2181) & (g2213) & (g1439) & (!g1473) & (!g3455) & (g3456)) + ((!g2181) & (g2213) & (g1439) & (g1473) & (!g3455) & (g3456)) + ((!g2181) & (g2213) & (g1439) & (g1473) & (g3455) & (g3456)) + ((g2181) & (!g2213) & (!g1439) & (g1473) & (!g3455) & (g3456)) + ((g2181) & (!g2213) & (g1439) & (g1473) & (!g3455) & (g3456)) + ((g2181) & (!g2213) & (g1439) & (g1473) & (g3455) & (g3456)) + ((g2181) & (g2213) & (!g1439) & (!g1473) & (!g3455) & (g3456)) + ((g2181) & (g2213) & (!g1439) & (g1473) & (!g3455) & (g3456)) + ((g2181) & (g2213) & (!g1439) & (g1473) & (g3455) & (g3456)) + ((g2181) & (g2213) & (g1439) & (!g1473) & (!g3455) & (g3456)) + ((g2181) & (g2213) & (g1439) & (!g1473) & (g3455) & (g3456)) + ((g2181) & (g2213) & (g1439) & (g1473) & (!g3455) & (g3456)) + ((g2181) & (g2213) & (g1439) & (g1473) & (g3455) & (g3456)));
	assign g3458 = (((g2263) & (g1507)));
	assign g3459 = (((!g2299) & (!g2348) & (!g1540) & (!g1577) & (!g3457) & (!g3458)) + ((!g2299) & (!g2348) & (!g1540) & (!g1577) & (!g3457) & (g3458)) + ((!g2299) & (!g2348) & (!g1540) & (!g1577) & (g3457) & (!g3458)) + ((!g2299) & (!g2348) & (!g1540) & (!g1577) & (g3457) & (g3458)) + ((!g2299) & (!g2348) & (!g1540) & (g1577) & (!g3457) & (!g3458)) + ((!g2299) & (!g2348) & (!g1540) & (g1577) & (!g3457) & (g3458)) + ((!g2299) & (!g2348) & (!g1540) & (g1577) & (g3457) & (!g3458)) + ((!g2299) & (!g2348) & (!g1540) & (g1577) & (g3457) & (g3458)) + ((!g2299) & (!g2348) & (g1540) & (!g1577) & (!g3457) & (!g3458)) + ((!g2299) & (!g2348) & (g1540) & (!g1577) & (!g3457) & (g3458)) + ((!g2299) & (!g2348) & (g1540) & (!g1577) & (g3457) & (!g3458)) + ((!g2299) & (!g2348) & (g1540) & (!g1577) & (g3457) & (g3458)) + ((!g2299) & (!g2348) & (g1540) & (g1577) & (!g3457) & (!g3458)) + ((!g2299) & (g2348) & (!g1540) & (!g1577) & (!g3457) & (!g3458)) + ((!g2299) & (g2348) & (!g1540) & (!g1577) & (!g3457) & (g3458)) + ((!g2299) & (g2348) & (!g1540) & (!g1577) & (g3457) & (!g3458)) + ((!g2299) & (g2348) & (!g1540) & (!g1577) & (g3457) & (g3458)) + ((!g2299) & (g2348) & (g1540) & (!g1577) & (!g3457) & (!g3458)) + ((g2299) & (!g2348) & (!g1540) & (!g1577) & (!g3457) & (!g3458)) + ((g2299) & (!g2348) & (!g1540) & (!g1577) & (!g3457) & (g3458)) + ((g2299) & (!g2348) & (!g1540) & (!g1577) & (g3457) & (!g3458)) + ((g2299) & (!g2348) & (!g1540) & (!g1577) & (g3457) & (g3458)) + ((g2299) & (!g2348) & (!g1540) & (g1577) & (!g3457) & (!g3458)) + ((g2299) & (!g2348) & (g1540) & (!g1577) & (!g3457) & (!g3458)) + ((g2299) & (!g2348) & (g1540) & (!g1577) & (!g3457) & (g3458)) + ((g2299) & (!g2348) & (g1540) & (!g1577) & (g3457) & (!g3458)) + ((g2299) & (!g2348) & (g1540) & (!g1577) & (g3457) & (g3458)) + ((g2299) & (g2348) & (!g1540) & (!g1577) & (!g3457) & (!g3458)));
	assign g3460 = (((!g2379) & (g1610) & (!g3459)) + ((g2379) & (!g1610) & (!g3459)) + ((g2379) & (g1610) & (!g3459)) + ((g2379) & (g1610) & (g3459)));
	assign g3461 = (((!g2427) & (g1644) & (g3460)) + ((g2427) & (!g1644) & (g3460)) + ((g2427) & (g1644) & (!g3460)) + ((g2427) & (g1644) & (g3460)));
	assign g3462 = (((!g830) & (!g1886) & (!g7070) & (key[96])) + ((!g830) & (!g1886) & (g7070) & (key[96])) + ((!g830) & (g1886) & (!g7070) & (key[96])) + ((!g830) & (g1886) & (g7070) & (key[96])) + ((g830) & (!g1886) & (g7070) & (!key[96])) + ((g830) & (!g1886) & (g7070) & (key[96])) + ((g830) & (g1886) & (!g7070) & (!key[96])) + ((g830) & (g1886) & (!g7070) & (key[96])));
	assign g3463 = (((!g1915) & (!g1916) & (!g1917) & (!g1918) & (!g1919) & (!g1920)));
	assign g3464 = (((!reset) & (!g830) & (!g1914) & (!g1922) & (!g2016) & (!g3463)) + ((!reset) & (!g830) & (!g1914) & (!g1922) & (!g2016) & (g3463)) + ((!reset) & (!g830) & (!g1914) & (g1922) & (!g2016) & (!g3463)) + ((!reset) & (!g830) & (!g1914) & (g1922) & (!g2016) & (g3463)) + ((!reset) & (!g830) & (g1914) & (!g1922) & (!g2016) & (!g3463)) + ((!reset) & (!g830) & (g1914) & (!g1922) & (!g2016) & (g3463)) + ((!reset) & (!g830) & (g1914) & (g1922) & (!g2016) & (!g3463)) + ((!reset) & (!g830) & (g1914) & (g1922) & (!g2016) & (g3463)) + ((!reset) & (g830) & (!g1914) & (!g1922) & (!g2016) & (!g3463)) + ((!reset) & (g830) & (!g1914) & (!g1922) & (!g2016) & (g3463)) + ((!reset) & (g830) & (!g1914) & (!g1922) & (g2016) & (!g3463)) + ((!reset) & (g830) & (!g1914) & (g1922) & (!g2016) & (!g3463)) + ((!reset) & (g830) & (!g1914) & (g1922) & (!g2016) & (g3463)) + ((!reset) & (g830) & (!g1914) & (g1922) & (g2016) & (!g3463)) + ((!reset) & (g830) & (!g1914) & (g1922) & (g2016) & (g3463)) + ((!reset) & (g830) & (g1914) & (!g1922) & (!g2016) & (!g3463)) + ((!reset) & (g830) & (g1914) & (!g1922) & (!g2016) & (g3463)) + ((!reset) & (g830) & (g1914) & (!g1922) & (g2016) & (!g3463)) + ((!reset) & (g830) & (g1914) & (!g1922) & (g2016) & (g3463)) + ((!reset) & (g830) & (g1914) & (g1922) & (!g2016) & (!g3463)) + ((!reset) & (g830) & (g1914) & (g1922) & (!g2016) & (g3463)) + ((!reset) & (g830) & (g1914) & (g1922) & (g2016) & (!g3463)) + ((reset) & (!g830) & (!g1914) & (!g1922) & (!g2016) & (!g3463)) + ((reset) & (!g830) & (!g1914) & (!g1922) & (!g2016) & (g3463)) + ((reset) & (!g830) & (!g1914) & (!g1922) & (g2016) & (!g3463)) + ((reset) & (!g830) & (!g1914) & (!g1922) & (g2016) & (g3463)) + ((reset) & (!g830) & (!g1914) & (g1922) & (!g2016) & (!g3463)) + ((reset) & (!g830) & (!g1914) & (g1922) & (!g2016) & (g3463)) + ((reset) & (!g830) & (!g1914) & (g1922) & (g2016) & (!g3463)) + ((reset) & (!g830) & (!g1914) & (g1922) & (g2016) & (g3463)) + ((reset) & (!g830) & (g1914) & (!g1922) & (!g2016) & (!g3463)) + ((reset) & (!g830) & (g1914) & (!g1922) & (!g2016) & (g3463)) + ((reset) & (!g830) & (g1914) & (!g1922) & (g2016) & (!g3463)) + ((reset) & (!g830) & (g1914) & (!g1922) & (g2016) & (g3463)) + ((reset) & (!g830) & (g1914) & (g1922) & (!g2016) & (!g3463)) + ((reset) & (!g830) & (g1914) & (g1922) & (!g2016) & (g3463)) + ((reset) & (!g830) & (g1914) & (g1922) & (g2016) & (!g3463)) + ((reset) & (!g830) & (g1914) & (g1922) & (g2016) & (g3463)) + ((reset) & (g830) & (!g1914) & (!g1922) & (!g2016) & (!g3463)) + ((reset) & (g830) & (!g1914) & (!g1922) & (!g2016) & (g3463)) + ((reset) & (g830) & (!g1914) & (!g1922) & (g2016) & (!g3463)) + ((reset) & (g830) & (!g1914) & (!g1922) & (g2016) & (g3463)) + ((reset) & (g830) & (!g1914) & (g1922) & (!g2016) & (!g3463)) + ((reset) & (g830) & (!g1914) & (g1922) & (!g2016) & (g3463)) + ((reset) & (g830) & (!g1914) & (g1922) & (g2016) & (!g3463)) + ((reset) & (g830) & (!g1914) & (g1922) & (g2016) & (g3463)) + ((reset) & (g830) & (g1914) & (!g1922) & (!g2016) & (!g3463)) + ((reset) & (g830) & (g1914) & (!g1922) & (!g2016) & (g3463)) + ((reset) & (g830) & (g1914) & (!g1922) & (g2016) & (!g3463)) + ((reset) & (g830) & (g1914) & (!g1922) & (g2016) & (g3463)) + ((reset) & (g830) & (g1914) & (g1922) & (!g2016) & (!g3463)) + ((reset) & (g830) & (g1914) & (g1922) & (!g2016) & (g3463)) + ((reset) & (g830) & (g1914) & (g1922) & (g2016) & (!g3463)) + ((reset) & (g830) & (g1914) & (g1922) & (g2016) & (g3463)));
	assign g3465 = (((!g1896) & (!g1912) & (!g2041) & (!g2045) & (g2068) & (g2091)) + ((!g1896) & (!g1912) & (!g2041) & (g2045) & (g2068) & (g2091)) + ((!g1896) & (!g1912) & (g2041) & (!g2045) & (g2068) & (g2091)) + ((!g1896) & (!g1912) & (g2041) & (g2045) & (!g2068) & (g2091)) + ((!g1896) & (!g1912) & (g2041) & (g2045) & (g2068) & (!g2091)) + ((!g1896) & (!g1912) & (g2041) & (g2045) & (g2068) & (g2091)) + ((!g1896) & (g1912) & (!g2041) & (!g2045) & (g2068) & (g2091)) + ((!g1896) & (g1912) & (!g2041) & (g2045) & (g2068) & (g2091)) + ((!g1896) & (g1912) & (g2041) & (!g2045) & (g2068) & (g2091)) + ((!g1896) & (g1912) & (g2041) & (g2045) & (!g2068) & (g2091)) + ((!g1896) & (g1912) & (g2041) & (g2045) & (g2068) & (!g2091)) + ((!g1896) & (g1912) & (g2041) & (g2045) & (g2068) & (g2091)) + ((g1896) & (!g1912) & (!g2041) & (!g2045) & (g2068) & (g2091)) + ((g1896) & (!g1912) & (!g2041) & (g2045) & (g2068) & (g2091)) + ((g1896) & (!g1912) & (g2041) & (!g2045) & (g2068) & (g2091)) + ((g1896) & (!g1912) & (g2041) & (g2045) & (!g2068) & (g2091)) + ((g1896) & (!g1912) & (g2041) & (g2045) & (g2068) & (!g2091)) + ((g1896) & (!g1912) & (g2041) & (g2045) & (g2068) & (g2091)) + ((g1896) & (g1912) & (!g2041) & (!g2045) & (g2068) & (g2091)) + ((g1896) & (g1912) & (!g2041) & (g2045) & (!g2068) & (g2091)) + ((g1896) & (g1912) & (!g2041) & (g2045) & (g2068) & (!g2091)) + ((g1896) & (g1912) & (!g2041) & (g2045) & (g2068) & (g2091)) + ((g1896) & (g1912) & (g2041) & (!g2045) & (!g2068) & (g2091)) + ((g1896) & (g1912) & (g2041) & (!g2045) & (g2068) & (!g2091)) + ((g1896) & (g1912) & (g2041) & (!g2045) & (g2068) & (g2091)) + ((g1896) & (g1912) & (g2041) & (g2045) & (!g2068) & (g2091)) + ((g1896) & (g1912) & (g2041) & (g2045) & (g2068) & (!g2091)) + ((g1896) & (g1912) & (g2041) & (g2045) & (g2068) & (g2091)));
	assign g3466 = (((!g2203) & (g2207)) + ((g2203) & (!g2207)));
	assign g3467 = (((!g3465) & (!g2123) & (!g2127) & (g2150) & (g2173) & (g3466)) + ((!g3465) & (!g2123) & (g2127) & (g2150) & (g2173) & (g3466)) + ((!g3465) & (g2123) & (!g2127) & (g2150) & (g2173) & (g3466)) + ((!g3465) & (g2123) & (g2127) & (!g2150) & (g2173) & (g3466)) + ((!g3465) & (g2123) & (g2127) & (g2150) & (!g2173) & (g3466)) + ((!g3465) & (g2123) & (g2127) & (g2150) & (g2173) & (g3466)) + ((g3465) & (!g2123) & (!g2127) & (g2150) & (g2173) & (g3466)) + ((g3465) & (!g2123) & (g2127) & (!g2150) & (g2173) & (g3466)) + ((g3465) & (!g2123) & (g2127) & (g2150) & (!g2173) & (g3466)) + ((g3465) & (!g2123) & (g2127) & (g2150) & (g2173) & (g3466)) + ((g3465) & (g2123) & (!g2127) & (!g2150) & (g2173) & (g3466)) + ((g3465) & (g2123) & (!g2127) & (g2150) & (!g2173) & (g3466)) + ((g3465) & (g2123) & (!g2127) & (g2150) & (g2173) & (g3466)) + ((g3465) & (g2123) & (g2127) & (!g2150) & (g2173) & (g3466)) + ((g3465) & (g2123) & (g2127) & (g2150) & (!g2173) & (g3466)) + ((g3465) & (g2123) & (g2127) & (g2150) & (g2173) & (g3466)));
	assign g3468 = (((g2203) & (g2207)));
	assign g3469 = (((!g3467) & (!g3468) & (!g2230) & (!g2253) & (!g2286) & (!g2290)) + ((!g3467) & (!g3468) & (!g2230) & (!g2253) & (!g2286) & (g2290)) + ((!g3467) & (!g3468) & (!g2230) & (!g2253) & (g2286) & (!g2290)) + ((!g3467) & (!g3468) & (!g2230) & (g2253) & (!g2286) & (!g2290)) + ((!g3467) & (!g3468) & (!g2230) & (g2253) & (!g2286) & (g2290)) + ((!g3467) & (!g3468) & (!g2230) & (g2253) & (g2286) & (!g2290)) + ((!g3467) & (!g3468) & (g2230) & (!g2253) & (!g2286) & (!g2290)) + ((!g3467) & (!g3468) & (g2230) & (!g2253) & (!g2286) & (g2290)) + ((!g3467) & (!g3468) & (g2230) & (!g2253) & (g2286) & (!g2290)) + ((!g3467) & (!g3468) & (g2230) & (g2253) & (!g2286) & (!g2290)) + ((!g3467) & (g3468) & (!g2230) & (!g2253) & (!g2286) & (!g2290)) + ((!g3467) & (g3468) & (!g2230) & (!g2253) & (!g2286) & (g2290)) + ((!g3467) & (g3468) & (!g2230) & (!g2253) & (g2286) & (!g2290)) + ((!g3467) & (g3468) & (!g2230) & (g2253) & (!g2286) & (!g2290)) + ((!g3467) & (g3468) & (g2230) & (!g2253) & (!g2286) & (!g2290)) + ((!g3467) & (g3468) & (g2230) & (g2253) & (!g2286) & (!g2290)) + ((g3467) & (!g3468) & (!g2230) & (!g2253) & (!g2286) & (!g2290)) + ((g3467) & (!g3468) & (!g2230) & (!g2253) & (!g2286) & (g2290)) + ((g3467) & (!g3468) & (!g2230) & (!g2253) & (g2286) & (!g2290)) + ((g3467) & (!g3468) & (!g2230) & (g2253) & (!g2286) & (!g2290)) + ((g3467) & (!g3468) & (g2230) & (!g2253) & (!g2286) & (!g2290)) + ((g3467) & (!g3468) & (g2230) & (g2253) & (!g2286) & (!g2290)) + ((g3467) & (g3468) & (!g2230) & (!g2253) & (!g2286) & (!g2290)) + ((g3467) & (g3468) & (!g2230) & (!g2253) & (!g2286) & (g2290)) + ((g3467) & (g3468) & (!g2230) & (!g2253) & (g2286) & (!g2290)) + ((g3467) & (g3468) & (!g2230) & (g2253) & (!g2286) & (!g2290)) + ((g3467) & (g3468) & (g2230) & (!g2253) & (!g2286) & (!g2290)) + ((g3467) & (g3468) & (g2230) & (g2253) & (!g2286) & (!g2290)));
	assign g3470 = (((!g2396) & (g2419)) + ((g2396) & (!g2419)));
	assign g3471 = (((!g3469) & (!g2317) & (!g2340) & (g2369) & (g2373) & (g3470)) + ((!g3469) & (!g2317) & (g2340) & (!g2369) & (g2373) & (g3470)) + ((!g3469) & (!g2317) & (g2340) & (g2369) & (!g2373) & (g3470)) + ((!g3469) & (!g2317) & (g2340) & (g2369) & (g2373) & (g3470)) + ((!g3469) & (g2317) & (!g2340) & (!g2369) & (g2373) & (g3470)) + ((!g3469) & (g2317) & (!g2340) & (g2369) & (!g2373) & (g3470)) + ((!g3469) & (g2317) & (!g2340) & (g2369) & (g2373) & (g3470)) + ((!g3469) & (g2317) & (g2340) & (!g2369) & (g2373) & (g3470)) + ((!g3469) & (g2317) & (g2340) & (g2369) & (!g2373) & (g3470)) + ((!g3469) & (g2317) & (g2340) & (g2369) & (g2373) & (g3470)) + ((g3469) & (!g2317) & (!g2340) & (g2369) & (g2373) & (g3470)) + ((g3469) & (!g2317) & (g2340) & (g2369) & (g2373) & (g3470)) + ((g3469) & (g2317) & (!g2340) & (g2369) & (g2373) & (g3470)) + ((g3469) & (g2317) & (g2340) & (!g2369) & (g2373) & (g3470)) + ((g3469) & (g2317) & (g2340) & (g2369) & (!g2373) & (g3470)) + ((g3469) & (g2317) & (g2340) & (g2369) & (g2373) & (g3470)));
	assign g3472 = (((g2396) & (g2419)));
	assign g3473 = (((!g3471) & (!g3472) & (!g2497) & (!g2509) & (!g2531) & (!g2546)) + ((!g3471) & (!g3472) & (!g2497) & (!g2509) & (!g2531) & (g2546)) + ((!g3471) & (!g3472) & (!g2497) & (!g2509) & (g2531) & (!g2546)) + ((!g3471) & (!g3472) & (!g2497) & (g2509) & (!g2531) & (!g2546)) + ((!g3471) & (!g3472) & (!g2497) & (g2509) & (!g2531) & (g2546)) + ((!g3471) & (!g3472) & (!g2497) & (g2509) & (g2531) & (!g2546)) + ((!g3471) & (!g3472) & (g2497) & (!g2509) & (!g2531) & (!g2546)) + ((!g3471) & (!g3472) & (g2497) & (!g2509) & (!g2531) & (g2546)) + ((!g3471) & (!g3472) & (g2497) & (!g2509) & (g2531) & (!g2546)) + ((!g3471) & (!g3472) & (g2497) & (g2509) & (!g2531) & (!g2546)) + ((!g3471) & (g3472) & (!g2497) & (!g2509) & (!g2531) & (!g2546)) + ((!g3471) & (g3472) & (!g2497) & (!g2509) & (!g2531) & (g2546)) + ((!g3471) & (g3472) & (!g2497) & (!g2509) & (g2531) & (!g2546)) + ((!g3471) & (g3472) & (!g2497) & (g2509) & (!g2531) & (!g2546)) + ((!g3471) & (g3472) & (g2497) & (!g2509) & (!g2531) & (!g2546)) + ((!g3471) & (g3472) & (g2497) & (g2509) & (!g2531) & (!g2546)) + ((g3471) & (!g3472) & (!g2497) & (!g2509) & (!g2531) & (!g2546)) + ((g3471) & (!g3472) & (!g2497) & (!g2509) & (!g2531) & (g2546)) + ((g3471) & (!g3472) & (!g2497) & (!g2509) & (g2531) & (!g2546)) + ((g3471) & (!g3472) & (!g2497) & (g2509) & (!g2531) & (!g2546)) + ((g3471) & (!g3472) & (g2497) & (!g2509) & (!g2531) & (!g2546)) + ((g3471) & (!g3472) & (g2497) & (g2509) & (!g2531) & (!g2546)) + ((g3471) & (g3472) & (!g2497) & (!g2509) & (!g2531) & (!g2546)) + ((g3471) & (g3472) & (!g2497) & (!g2509) & (!g2531) & (g2546)) + ((g3471) & (g3472) & (!g2497) & (!g2509) & (g2531) & (!g2546)) + ((g3471) & (g3472) & (!g2497) & (g2509) & (!g2531) & (!g2546)) + ((g3471) & (g3472) & (g2497) & (!g2509) & (!g2531) & (!g2546)) + ((g3471) & (g3472) & (g2497) & (g2509) & (!g2531) & (!g2546)));
	assign g3474 = (((!g2672) & (g2676)) + ((g2672) & (!g2676)));
	assign g3475 = (((!g3473) & (!g2589) & (!g2595) & (g2620) & (g2643) & (g3474)) + ((!g3473) & (!g2589) & (g2595) & (!g2620) & (g2643) & (g3474)) + ((!g3473) & (!g2589) & (g2595) & (g2620) & (!g2643) & (g3474)) + ((!g3473) & (!g2589) & (g2595) & (g2620) & (g2643) & (g3474)) + ((!g3473) & (g2589) & (!g2595) & (!g2620) & (g2643) & (g3474)) + ((!g3473) & (g2589) & (!g2595) & (g2620) & (!g2643) & (g3474)) + ((!g3473) & (g2589) & (!g2595) & (g2620) & (g2643) & (g3474)) + ((!g3473) & (g2589) & (g2595) & (!g2620) & (g2643) & (g3474)) + ((!g3473) & (g2589) & (g2595) & (g2620) & (!g2643) & (g3474)) + ((!g3473) & (g2589) & (g2595) & (g2620) & (g2643) & (g3474)) + ((g3473) & (!g2589) & (!g2595) & (g2620) & (g2643) & (g3474)) + ((g3473) & (!g2589) & (g2595) & (g2620) & (g2643) & (g3474)) + ((g3473) & (g2589) & (!g2595) & (g2620) & (g2643) & (g3474)) + ((g3473) & (g2589) & (g2595) & (!g2620) & (g2643) & (g3474)) + ((g3473) & (g2589) & (g2595) & (g2620) & (!g2643) & (g3474)) + ((g3473) & (g2589) & (g2595) & (g2620) & (g2643) & (g3474)));
	assign g3476 = (((g2672) & (g2676)));
	assign g3477 = (((!g3475) & (!g3476) & (!g2713) & (!g2752) & (!g2783) & (!g2787)) + ((!g3475) & (!g3476) & (!g2713) & (!g2752) & (!g2783) & (g2787)) + ((!g3475) & (!g3476) & (!g2713) & (!g2752) & (g2783) & (!g2787)) + ((!g3475) & (!g3476) & (!g2713) & (g2752) & (!g2783) & (!g2787)) + ((!g3475) & (!g3476) & (!g2713) & (g2752) & (!g2783) & (g2787)) + ((!g3475) & (!g3476) & (!g2713) & (g2752) & (g2783) & (!g2787)) + ((!g3475) & (!g3476) & (g2713) & (!g2752) & (!g2783) & (!g2787)) + ((!g3475) & (!g3476) & (g2713) & (!g2752) & (!g2783) & (g2787)) + ((!g3475) & (!g3476) & (g2713) & (!g2752) & (g2783) & (!g2787)) + ((!g3475) & (!g3476) & (g2713) & (g2752) & (!g2783) & (!g2787)) + ((!g3475) & (g3476) & (!g2713) & (!g2752) & (!g2783) & (!g2787)) + ((!g3475) & (g3476) & (!g2713) & (!g2752) & (!g2783) & (g2787)) + ((!g3475) & (g3476) & (!g2713) & (!g2752) & (g2783) & (!g2787)) + ((!g3475) & (g3476) & (!g2713) & (g2752) & (!g2783) & (!g2787)) + ((!g3475) & (g3476) & (g2713) & (!g2752) & (!g2783) & (!g2787)) + ((!g3475) & (g3476) & (g2713) & (g2752) & (!g2783) & (!g2787)) + ((g3475) & (!g3476) & (!g2713) & (!g2752) & (!g2783) & (!g2787)) + ((g3475) & (!g3476) & (!g2713) & (!g2752) & (!g2783) & (g2787)) + ((g3475) & (!g3476) & (!g2713) & (!g2752) & (g2783) & (!g2787)) + ((g3475) & (!g3476) & (!g2713) & (g2752) & (!g2783) & (!g2787)) + ((g3475) & (!g3476) & (g2713) & (!g2752) & (!g2783) & (!g2787)) + ((g3475) & (!g3476) & (g2713) & (g2752) & (!g2783) & (!g2787)) + ((g3475) & (g3476) & (!g2713) & (!g2752) & (!g2783) & (!g2787)) + ((g3475) & (g3476) & (!g2713) & (!g2752) & (!g2783) & (g2787)) + ((g3475) & (g3476) & (!g2713) & (!g2752) & (g2783) & (!g2787)) + ((g3475) & (g3476) & (!g2713) & (g2752) & (!g2783) & (!g2787)) + ((g3475) & (g3476) & (g2713) & (!g2752) & (!g2783) & (!g2787)) + ((g3475) & (g3476) & (g2713) & (g2752) & (!g2783) & (!g2787)));
	assign g3478 = (((!g2889) & (g2904)) + ((g2889) & (!g2904)));
	assign g3479 = (((!g3477) & (!g2810) & (!g2833) & (g2868) & (g2874) & (g3478)) + ((!g3477) & (!g2810) & (g2833) & (!g2868) & (g2874) & (g3478)) + ((!g3477) & (!g2810) & (g2833) & (g2868) & (!g2874) & (g3478)) + ((!g3477) & (!g2810) & (g2833) & (g2868) & (g2874) & (g3478)) + ((!g3477) & (g2810) & (!g2833) & (!g2868) & (g2874) & (g3478)) + ((!g3477) & (g2810) & (!g2833) & (g2868) & (!g2874) & (g3478)) + ((!g3477) & (g2810) & (!g2833) & (g2868) & (g2874) & (g3478)) + ((!g3477) & (g2810) & (g2833) & (!g2868) & (g2874) & (g3478)) + ((!g3477) & (g2810) & (g2833) & (g2868) & (!g2874) & (g3478)) + ((!g3477) & (g2810) & (g2833) & (g2868) & (g2874) & (g3478)) + ((g3477) & (!g2810) & (!g2833) & (g2868) & (g2874) & (g3478)) + ((g3477) & (!g2810) & (g2833) & (g2868) & (g2874) & (g3478)) + ((g3477) & (g2810) & (!g2833) & (g2868) & (g2874) & (g3478)) + ((g3477) & (g2810) & (g2833) & (!g2868) & (g2874) & (g3478)) + ((g3477) & (g2810) & (g2833) & (g2868) & (!g2874) & (g3478)) + ((g3477) & (g2810) & (g2833) & (g2868) & (g2874) & (g3478)));
	assign g3480 = (((g2889) & (g2904)));
	assign g3481 = (((!g3479) & (!g3480) & (!g2979) & (!g2991) & (!g3007) & (!g3022)) + ((!g3479) & (!g3480) & (!g2979) & (!g2991) & (!g3007) & (g3022)) + ((!g3479) & (!g3480) & (!g2979) & (!g2991) & (g3007) & (!g3022)) + ((!g3479) & (!g3480) & (!g2979) & (g2991) & (!g3007) & (!g3022)) + ((!g3479) & (!g3480) & (!g2979) & (g2991) & (!g3007) & (g3022)) + ((!g3479) & (!g3480) & (!g2979) & (g2991) & (g3007) & (!g3022)) + ((!g3479) & (!g3480) & (g2979) & (!g2991) & (!g3007) & (!g3022)) + ((!g3479) & (!g3480) & (g2979) & (!g2991) & (!g3007) & (g3022)) + ((!g3479) & (!g3480) & (g2979) & (!g2991) & (g3007) & (!g3022)) + ((!g3479) & (!g3480) & (g2979) & (g2991) & (!g3007) & (!g3022)) + ((!g3479) & (g3480) & (!g2979) & (!g2991) & (!g3007) & (!g3022)) + ((!g3479) & (g3480) & (!g2979) & (!g2991) & (!g3007) & (g3022)) + ((!g3479) & (g3480) & (!g2979) & (!g2991) & (g3007) & (!g3022)) + ((!g3479) & (g3480) & (!g2979) & (g2991) & (!g3007) & (!g3022)) + ((!g3479) & (g3480) & (g2979) & (!g2991) & (!g3007) & (!g3022)) + ((!g3479) & (g3480) & (g2979) & (g2991) & (!g3007) & (!g3022)) + ((g3479) & (!g3480) & (!g2979) & (!g2991) & (!g3007) & (!g3022)) + ((g3479) & (!g3480) & (!g2979) & (!g2991) & (!g3007) & (g3022)) + ((g3479) & (!g3480) & (!g2979) & (!g2991) & (g3007) & (!g3022)) + ((g3479) & (!g3480) & (!g2979) & (g2991) & (!g3007) & (!g3022)) + ((g3479) & (!g3480) & (g2979) & (!g2991) & (!g3007) & (!g3022)) + ((g3479) & (!g3480) & (g2979) & (g2991) & (!g3007) & (!g3022)) + ((g3479) & (g3480) & (!g2979) & (!g2991) & (!g3007) & (!g3022)) + ((g3479) & (g3480) & (!g2979) & (!g2991) & (!g3007) & (g3022)) + ((g3479) & (g3480) & (!g2979) & (!g2991) & (g3007) & (!g3022)) + ((g3479) & (g3480) & (!g2979) & (g2991) & (!g3007) & (!g3022)) + ((g3479) & (g3480) & (g2979) & (!g2991) & (!g3007) & (!g3022)) + ((g3479) & (g3480) & (g2979) & (g2991) & (!g3007) & (!g3022)));
	assign g3482 = (((!g3481) & (!g3061) & (g3067)) + ((!g3481) & (g3061) & (!g3067)) + ((!g3481) & (g3061) & (g3067)) + ((g3481) & (g3061) & (g3067)));
	assign g3483 = (((!g1884) & (!g1977) & (g1979) & (!g1886) & (!g2032) & (g2055)) + ((!g1884) & (!g1977) & (g1979) & (!g1886) & (g2032) & (g2055)) + ((!g1884) & (!g1977) & (g1979) & (g1886) & (!g2032) & (g2055)) + ((!g1884) & (!g1977) & (g1979) & (g1886) & (g2032) & (g2055)) + ((!g1884) & (g1977) & (!g1979) & (!g1886) & (g2032) & (g2055)) + ((!g1884) & (g1977) & (!g1979) & (g1886) & (g2032) & (g2055)) + ((!g1884) & (g1977) & (g1979) & (!g1886) & (!g2032) & (g2055)) + ((!g1884) & (g1977) & (g1979) & (!g1886) & (g2032) & (!g2055)) + ((!g1884) & (g1977) & (g1979) & (!g1886) & (g2032) & (g2055)) + ((!g1884) & (g1977) & (g1979) & (g1886) & (!g2032) & (g2055)) + ((!g1884) & (g1977) & (g1979) & (g1886) & (g2032) & (!g2055)) + ((!g1884) & (g1977) & (g1979) & (g1886) & (g2032) & (g2055)) + ((g1884) & (!g1977) & (!g1979) & (g1886) & (g2032) & (g2055)) + ((g1884) & (!g1977) & (g1979) & (!g1886) & (!g2032) & (g2055)) + ((g1884) & (!g1977) & (g1979) & (!g1886) & (g2032) & (g2055)) + ((g1884) & (!g1977) & (g1979) & (g1886) & (!g2032) & (g2055)) + ((g1884) & (!g1977) & (g1979) & (g1886) & (g2032) & (!g2055)) + ((g1884) & (!g1977) & (g1979) & (g1886) & (g2032) & (g2055)) + ((g1884) & (g1977) & (!g1979) & (!g1886) & (g2032) & (g2055)) + ((g1884) & (g1977) & (!g1979) & (g1886) & (!g2032) & (g2055)) + ((g1884) & (g1977) & (!g1979) & (g1886) & (g2032) & (g2055)) + ((g1884) & (g1977) & (g1979) & (!g1886) & (!g2032) & (g2055)) + ((g1884) & (g1977) & (g1979) & (!g1886) & (g2032) & (!g2055)) + ((g1884) & (g1977) & (g1979) & (!g1886) & (g2032) & (g2055)) + ((g1884) & (g1977) & (g1979) & (g1886) & (!g2032) & (!g2055)) + ((g1884) & (g1977) & (g1979) & (g1886) & (!g2032) & (g2055)) + ((g1884) & (g1977) & (g1979) & (g1886) & (g2032) & (!g2055)) + ((g1884) & (g1977) & (g1979) & (g1886) & (g2032) & (g2055)));
	assign g3484 = (((!g1986) & (g2194)) + ((g1986) & (!g2194)));
	assign g3485 = (((!g1982) & (!g1984) & (g2114) & (g2137) & (g3483) & (g3484)) + ((!g1982) & (g1984) & (!g2114) & (g2137) & (!g3483) & (g3484)) + ((!g1982) & (g1984) & (!g2114) & (g2137) & (g3483) & (g3484)) + ((!g1982) & (g1984) & (g2114) & (!g2137) & (g3483) & (g3484)) + ((!g1982) & (g1984) & (g2114) & (g2137) & (!g3483) & (g3484)) + ((!g1982) & (g1984) & (g2114) & (g2137) & (g3483) & (g3484)) + ((g1982) & (!g1984) & (!g2114) & (g2137) & (g3483) & (g3484)) + ((g1982) & (!g1984) & (g2114) & (g2137) & (!g3483) & (g3484)) + ((g1982) & (!g1984) & (g2114) & (g2137) & (g3483) & (g3484)) + ((g1982) & (g1984) & (!g2114) & (!g2137) & (g3483) & (g3484)) + ((g1982) & (g1984) & (!g2114) & (g2137) & (!g3483) & (g3484)) + ((g1982) & (g1984) & (!g2114) & (g2137) & (g3483) & (g3484)) + ((g1982) & (g1984) & (g2114) & (!g2137) & (!g3483) & (g3484)) + ((g1982) & (g1984) & (g2114) & (!g2137) & (g3483) & (g3484)) + ((g1982) & (g1984) & (g2114) & (g2137) & (!g3483) & (g3484)) + ((g1982) & (g1984) & (g2114) & (g2137) & (g3483) & (g3484)));
	assign g3486 = (((g1986) & (g2194)));
	assign g3487 = (((!g1991) & (!g1993) & (!g2217) & (!g2277) & (!g3485) & (!g3486)) + ((!g1991) & (!g1993) & (!g2217) & (!g2277) & (!g3485) & (g3486)) + ((!g1991) & (!g1993) & (!g2217) & (!g2277) & (g3485) & (!g3486)) + ((!g1991) & (!g1993) & (!g2217) & (!g2277) & (g3485) & (g3486)) + ((!g1991) & (!g1993) & (!g2217) & (g2277) & (!g3485) & (!g3486)) + ((!g1991) & (!g1993) & (!g2217) & (g2277) & (!g3485) & (g3486)) + ((!g1991) & (!g1993) & (!g2217) & (g2277) & (g3485) & (!g3486)) + ((!g1991) & (!g1993) & (!g2217) & (g2277) & (g3485) & (g3486)) + ((!g1991) & (!g1993) & (g2217) & (!g2277) & (!g3485) & (!g3486)) + ((!g1991) & (!g1993) & (g2217) & (!g2277) & (!g3485) & (g3486)) + ((!g1991) & (!g1993) & (g2217) & (!g2277) & (g3485) & (!g3486)) + ((!g1991) & (!g1993) & (g2217) & (!g2277) & (g3485) & (g3486)) + ((!g1991) & (!g1993) & (g2217) & (g2277) & (!g3485) & (!g3486)) + ((!g1991) & (g1993) & (!g2217) & (!g2277) & (!g3485) & (!g3486)) + ((!g1991) & (g1993) & (!g2217) & (!g2277) & (!g3485) & (g3486)) + ((!g1991) & (g1993) & (!g2217) & (!g2277) & (g3485) & (!g3486)) + ((!g1991) & (g1993) & (!g2217) & (!g2277) & (g3485) & (g3486)) + ((!g1991) & (g1993) & (g2217) & (!g2277) & (!g3485) & (!g3486)) + ((g1991) & (!g1993) & (!g2217) & (!g2277) & (!g3485) & (!g3486)) + ((g1991) & (!g1993) & (!g2217) & (!g2277) & (!g3485) & (g3486)) + ((g1991) & (!g1993) & (!g2217) & (!g2277) & (g3485) & (!g3486)) + ((g1991) & (!g1993) & (!g2217) & (!g2277) & (g3485) & (g3486)) + ((g1991) & (!g1993) & (!g2217) & (g2277) & (!g3485) & (!g3486)) + ((g1991) & (!g1993) & (g2217) & (!g2277) & (!g3485) & (!g3486)) + ((g1991) & (!g1993) & (g2217) & (!g2277) & (!g3485) & (g3486)) + ((g1991) & (!g1993) & (g2217) & (!g2277) & (g3485) & (!g3486)) + ((g1991) & (!g1993) & (g2217) & (!g2277) & (g3485) & (g3486)) + ((g1991) & (g1993) & (!g2217) & (!g2277) & (!g3485) & (!g3486)));
	assign g3488 = (((!g2001) & (g2383)) + ((g2001) & (!g2383)));
	assign g3489 = (((!g1996) & (!g1998) & (g2304) & (g2360) & (!g3487) & (g3488)) + ((!g1996) & (g1998) & (!g2304) & (g2360) & (!g3487) & (g3488)) + ((!g1996) & (g1998) & (!g2304) & (g2360) & (g3487) & (g3488)) + ((!g1996) & (g1998) & (g2304) & (!g2360) & (!g3487) & (g3488)) + ((!g1996) & (g1998) & (g2304) & (g2360) & (!g3487) & (g3488)) + ((!g1996) & (g1998) & (g2304) & (g2360) & (g3487) & (g3488)) + ((g1996) & (!g1998) & (!g2304) & (g2360) & (!g3487) & (g3488)) + ((g1996) & (!g1998) & (g2304) & (g2360) & (!g3487) & (g3488)) + ((g1996) & (!g1998) & (g2304) & (g2360) & (g3487) & (g3488)) + ((g1996) & (g1998) & (!g2304) & (!g2360) & (!g3487) & (g3488)) + ((g1996) & (g1998) & (!g2304) & (g2360) & (!g3487) & (g3488)) + ((g1996) & (g1998) & (!g2304) & (g2360) & (g3487) & (g3488)) + ((g1996) & (g1998) & (g2304) & (!g2360) & (!g3487) & (g3488)) + ((g1996) & (g1998) & (g2304) & (!g2360) & (g3487) & (g3488)) + ((g1996) & (g1998) & (g2304) & (g2360) & (!g3487) & (g3488)) + ((g1996) & (g1998) & (g2304) & (g2360) & (g3487) & (g3488)));
	assign g3490 = (((g2001) & (g2383)));
	assign g3491 = (((!g2003) & (!g2005) & (!g2468) & (!g2523) & (!g3489) & (!g3490)) + ((!g2003) & (!g2005) & (!g2468) & (!g2523) & (!g3489) & (g3490)) + ((!g2003) & (!g2005) & (!g2468) & (!g2523) & (g3489) & (!g3490)) + ((!g2003) & (!g2005) & (!g2468) & (!g2523) & (g3489) & (g3490)) + ((!g2003) & (!g2005) & (!g2468) & (g2523) & (!g3489) & (!g3490)) + ((!g2003) & (!g2005) & (!g2468) & (g2523) & (!g3489) & (g3490)) + ((!g2003) & (!g2005) & (!g2468) & (g2523) & (g3489) & (!g3490)) + ((!g2003) & (!g2005) & (!g2468) & (g2523) & (g3489) & (g3490)) + ((!g2003) & (!g2005) & (g2468) & (!g2523) & (!g3489) & (!g3490)) + ((!g2003) & (!g2005) & (g2468) & (!g2523) & (!g3489) & (g3490)) + ((!g2003) & (!g2005) & (g2468) & (!g2523) & (g3489) & (!g3490)) + ((!g2003) & (!g2005) & (g2468) & (!g2523) & (g3489) & (g3490)) + ((!g2003) & (!g2005) & (g2468) & (g2523) & (!g3489) & (!g3490)) + ((!g2003) & (g2005) & (!g2468) & (!g2523) & (!g3489) & (!g3490)) + ((!g2003) & (g2005) & (!g2468) & (!g2523) & (!g3489) & (g3490)) + ((!g2003) & (g2005) & (!g2468) & (!g2523) & (g3489) & (!g3490)) + ((!g2003) & (g2005) & (!g2468) & (!g2523) & (g3489) & (g3490)) + ((!g2003) & (g2005) & (g2468) & (!g2523) & (!g3489) & (!g3490)) + ((g2003) & (!g2005) & (!g2468) & (!g2523) & (!g3489) & (!g3490)) + ((g2003) & (!g2005) & (!g2468) & (!g2523) & (!g3489) & (g3490)) + ((g2003) & (!g2005) & (!g2468) & (!g2523) & (g3489) & (!g3490)) + ((g2003) & (!g2005) & (!g2468) & (!g2523) & (g3489) & (g3490)) + ((g2003) & (!g2005) & (!g2468) & (g2523) & (!g3489) & (!g3490)) + ((g2003) & (!g2005) & (g2468) & (!g2523) & (!g3489) & (!g3490)) + ((g2003) & (!g2005) & (g2468) & (!g2523) & (!g3489) & (g3490)) + ((g2003) & (!g2005) & (g2468) & (!g2523) & (g3489) & (!g3490)) + ((g2003) & (!g2005) & (g2468) & (!g2523) & (g3489) & (g3490)) + ((g2003) & (g2005) & (!g2468) & (!g2523) & (!g3489) & (!g3490)));
	assign g3492 = (((!g2051) & (g2663)) + ((g2051) & (!g2663)));
	assign g3493 = (((!g2011) & (!g2013) & (g2575) & (g2607) & (!g3491) & (g3492)) + ((!g2011) & (g2013) & (!g2575) & (g2607) & (!g3491) & (g3492)) + ((!g2011) & (g2013) & (!g2575) & (g2607) & (g3491) & (g3492)) + ((!g2011) & (g2013) & (g2575) & (!g2607) & (!g3491) & (g3492)) + ((!g2011) & (g2013) & (g2575) & (g2607) & (!g3491) & (g3492)) + ((!g2011) & (g2013) & (g2575) & (g2607) & (g3491) & (g3492)) + ((g2011) & (!g2013) & (!g2575) & (g2607) & (!g3491) & (g3492)) + ((g2011) & (!g2013) & (g2575) & (g2607) & (!g3491) & (g3492)) + ((g2011) & (!g2013) & (g2575) & (g2607) & (g3491) & (g3492)) + ((g2011) & (g2013) & (!g2575) & (!g2607) & (!g3491) & (g3492)) + ((g2011) & (g2013) & (!g2575) & (g2607) & (!g3491) & (g3492)) + ((g2011) & (g2013) & (!g2575) & (g2607) & (g3491) & (g3492)) + ((g2011) & (g2013) & (g2575) & (!g2607) & (!g3491) & (g3492)) + ((g2011) & (g2013) & (g2575) & (!g2607) & (g3491) & (g3492)) + ((g2011) & (g2013) & (g2575) & (g2607) & (!g3491) & (g3492)) + ((g2011) & (g2013) & (g2575) & (g2607) & (g3491) & (g3492)));
	assign g3494 = (((g2051) & (g2663)));
	assign g3495 = (((!g2100) & (!g2133) & (!g2690) & (!g2774) & (!g3493) & (!g3494)) + ((!g2100) & (!g2133) & (!g2690) & (!g2774) & (!g3493) & (g3494)) + ((!g2100) & (!g2133) & (!g2690) & (!g2774) & (g3493) & (!g3494)) + ((!g2100) & (!g2133) & (!g2690) & (!g2774) & (g3493) & (g3494)) + ((!g2100) & (!g2133) & (!g2690) & (g2774) & (!g3493) & (!g3494)) + ((!g2100) & (!g2133) & (!g2690) & (g2774) & (!g3493) & (g3494)) + ((!g2100) & (!g2133) & (!g2690) & (g2774) & (g3493) & (!g3494)) + ((!g2100) & (!g2133) & (!g2690) & (g2774) & (g3493) & (g3494)) + ((!g2100) & (!g2133) & (g2690) & (!g2774) & (!g3493) & (!g3494)) + ((!g2100) & (!g2133) & (g2690) & (!g2774) & (!g3493) & (g3494)) + ((!g2100) & (!g2133) & (g2690) & (!g2774) & (g3493) & (!g3494)) + ((!g2100) & (!g2133) & (g2690) & (!g2774) & (g3493) & (g3494)) + ((!g2100) & (!g2133) & (g2690) & (g2774) & (!g3493) & (!g3494)) + ((!g2100) & (g2133) & (!g2690) & (!g2774) & (!g3493) & (!g3494)) + ((!g2100) & (g2133) & (!g2690) & (!g2774) & (!g3493) & (g3494)) + ((!g2100) & (g2133) & (!g2690) & (!g2774) & (g3493) & (!g3494)) + ((!g2100) & (g2133) & (!g2690) & (!g2774) & (g3493) & (g3494)) + ((!g2100) & (g2133) & (g2690) & (!g2774) & (!g3493) & (!g3494)) + ((g2100) & (!g2133) & (!g2690) & (!g2774) & (!g3493) & (!g3494)) + ((g2100) & (!g2133) & (!g2690) & (!g2774) & (!g3493) & (g3494)) + ((g2100) & (!g2133) & (!g2690) & (!g2774) & (g3493) & (!g3494)) + ((g2100) & (!g2133) & (!g2690) & (!g2774) & (g3493) & (g3494)) + ((g2100) & (!g2133) & (!g2690) & (g2774) & (!g3493) & (!g3494)) + ((g2100) & (!g2133) & (g2690) & (!g2774) & (!g3493) & (!g3494)) + ((g2100) & (!g2133) & (g2690) & (!g2774) & (!g3493) & (g3494)) + ((g2100) & (!g2133) & (g2690) & (!g2774) & (g3493) & (!g3494)) + ((g2100) & (!g2133) & (g2690) & (!g2774) & (g3493) & (g3494)) + ((g2100) & (g2133) & (!g2690) & (!g2774) & (!g3493) & (!g3494)));
	assign g3496 = (((!g2180) & (g2797) & (!g3495)) + ((g2180) & (!g2797) & (!g3495)) + ((g2180) & (g2797) & (!g3495)) + ((g2180) & (g2797) & (g3495)));
	assign g3497 = (((!g2212) & (!g2854) & (g3496)) + ((!g2212) & (g2854) & (!g3496)) + ((g2212) & (!g2854) & (!g3496)) + ((g2212) & (g2854) & (g3496)));
	assign g3498 = (((!g830) & (!g1888) & (!g7059) & (key[160])) + ((!g830) & (!g1888) & (g7059) & (key[160])) + ((!g830) & (g1888) & (!g7059) & (key[160])) + ((!g830) & (g1888) & (g7059) & (key[160])) + ((g830) & (!g1888) & (g7059) & (!key[160])) + ((g830) & (!g1888) & (g7059) & (key[160])) + ((g830) & (g1888) & (!g7059) & (!key[160])) + ((g830) & (g1888) & (!g7059) & (key[160])));
	assign g3499 = (((!reset) & (!g830) & (!g1914) & (!g1922) & (!g2016) & (!g3463)) + ((!reset) & (!g830) & (!g1914) & (!g1922) & (!g2016) & (g3463)) + ((!reset) & (!g830) & (!g1914) & (g1922) & (!g2016) & (!g3463)) + ((!reset) & (!g830) & (!g1914) & (g1922) & (!g2016) & (g3463)) + ((!reset) & (!g830) & (g1914) & (!g1922) & (!g2016) & (!g3463)) + ((!reset) & (!g830) & (g1914) & (!g1922) & (!g2016) & (g3463)) + ((!reset) & (!g830) & (g1914) & (g1922) & (!g2016) & (!g3463)) + ((!reset) & (!g830) & (g1914) & (g1922) & (!g2016) & (g3463)) + ((!reset) & (g830) & (!g1914) & (!g1922) & (!g2016) & (!g3463)) + ((!reset) & (g830) & (!g1914) & (!g1922) & (!g2016) & (g3463)) + ((!reset) & (g830) & (!g1914) & (!g1922) & (g2016) & (!g3463)) + ((!reset) & (g830) & (!g1914) & (!g1922) & (g2016) & (g3463)) + ((!reset) & (g830) & (!g1914) & (g1922) & (!g2016) & (!g3463)) + ((!reset) & (g830) & (!g1914) & (g1922) & (!g2016) & (g3463)) + ((!reset) & (g830) & (!g1914) & (g1922) & (g2016) & (!g3463)) + ((!reset) & (g830) & (g1914) & (!g1922) & (!g2016) & (!g3463)) + ((!reset) & (g830) & (g1914) & (!g1922) & (!g2016) & (g3463)) + ((!reset) & (g830) & (g1914) & (!g1922) & (g2016) & (!g3463)) + ((!reset) & (g830) & (g1914) & (g1922) & (!g2016) & (!g3463)) + ((!reset) & (g830) & (g1914) & (g1922) & (!g2016) & (g3463)) + ((!reset) & (g830) & (g1914) & (g1922) & (g2016) & (!g3463)) + ((!reset) & (g830) & (g1914) & (g1922) & (g2016) & (g3463)) + ((reset) & (!g830) & (!g1914) & (!g1922) & (!g2016) & (!g3463)) + ((reset) & (!g830) & (!g1914) & (!g1922) & (!g2016) & (g3463)) + ((reset) & (!g830) & (!g1914) & (!g1922) & (g2016) & (!g3463)) + ((reset) & (!g830) & (!g1914) & (!g1922) & (g2016) & (g3463)) + ((reset) & (!g830) & (!g1914) & (g1922) & (!g2016) & (!g3463)) + ((reset) & (!g830) & (!g1914) & (g1922) & (!g2016) & (g3463)) + ((reset) & (!g830) & (!g1914) & (g1922) & (g2016) & (!g3463)) + ((reset) & (!g830) & (!g1914) & (g1922) & (g2016) & (g3463)) + ((reset) & (!g830) & (g1914) & (!g1922) & (!g2016) & (!g3463)) + ((reset) & (!g830) & (g1914) & (!g1922) & (!g2016) & (g3463)) + ((reset) & (!g830) & (g1914) & (!g1922) & (g2016) & (!g3463)) + ((reset) & (!g830) & (g1914) & (!g1922) & (g2016) & (g3463)) + ((reset) & (!g830) & (g1914) & (g1922) & (!g2016) & (!g3463)) + ((reset) & (!g830) & (g1914) & (g1922) & (!g2016) & (g3463)) + ((reset) & (!g830) & (g1914) & (g1922) & (g2016) & (!g3463)) + ((reset) & (!g830) & (g1914) & (g1922) & (g2016) & (g3463)) + ((reset) & (g830) & (!g1914) & (!g1922) & (!g2016) & (!g3463)) + ((reset) & (g830) & (!g1914) & (!g1922) & (!g2016) & (g3463)) + ((reset) & (g830) & (!g1914) & (!g1922) & (g2016) & (!g3463)) + ((reset) & (g830) & (!g1914) & (!g1922) & (g2016) & (g3463)) + ((reset) & (g830) & (!g1914) & (g1922) & (!g2016) & (!g3463)) + ((reset) & (g830) & (!g1914) & (g1922) & (!g2016) & (g3463)) + ((reset) & (g830) & (!g1914) & (g1922) & (g2016) & (!g3463)) + ((reset) & (g830) & (!g1914) & (g1922) & (g2016) & (g3463)) + ((reset) & (g830) & (g1914) & (!g1922) & (!g2016) & (!g3463)) + ((reset) & (g830) & (g1914) & (!g1922) & (!g2016) & (g3463)) + ((reset) & (g830) & (g1914) & (!g1922) & (g2016) & (!g3463)) + ((reset) & (g830) & (g1914) & (!g1922) & (g2016) & (g3463)) + ((reset) & (g830) & (g1914) & (g1922) & (!g2016) & (!g3463)) + ((reset) & (g830) & (g1914) & (g1922) & (!g2016) & (g3463)) + ((reset) & (g830) & (g1914) & (g1922) & (g2016) & (!g3463)) + ((reset) & (g830) & (g1914) & (g1922) & (g2016) & (g3463)));
	assign g3500 = (((!g828) & (!g864) & (g897) & (!g1898) & (!g2022) & (g2071)) + ((!g828) & (!g864) & (g897) & (!g1898) & (g2022) & (g2071)) + ((!g828) & (!g864) & (g897) & (g1898) & (!g2022) & (g2071)) + ((!g828) & (!g864) & (g897) & (g1898) & (g2022) & (g2071)) + ((!g828) & (g864) & (!g897) & (!g1898) & (g2022) & (g2071)) + ((!g828) & (g864) & (!g897) & (g1898) & (g2022) & (g2071)) + ((!g828) & (g864) & (g897) & (!g1898) & (!g2022) & (g2071)) + ((!g828) & (g864) & (g897) & (!g1898) & (g2022) & (!g2071)) + ((!g828) & (g864) & (g897) & (!g1898) & (g2022) & (g2071)) + ((!g828) & (g864) & (g897) & (g1898) & (!g2022) & (g2071)) + ((!g828) & (g864) & (g897) & (g1898) & (g2022) & (!g2071)) + ((!g828) & (g864) & (g897) & (g1898) & (g2022) & (g2071)) + ((g828) & (!g864) & (!g897) & (g1898) & (g2022) & (g2071)) + ((g828) & (!g864) & (g897) & (!g1898) & (!g2022) & (g2071)) + ((g828) & (!g864) & (g897) & (!g1898) & (g2022) & (g2071)) + ((g828) & (!g864) & (g897) & (g1898) & (!g2022) & (g2071)) + ((g828) & (!g864) & (g897) & (g1898) & (g2022) & (!g2071)) + ((g828) & (!g864) & (g897) & (g1898) & (g2022) & (g2071)) + ((g828) & (g864) & (!g897) & (!g1898) & (g2022) & (g2071)) + ((g828) & (g864) & (!g897) & (g1898) & (!g2022) & (g2071)) + ((g828) & (g864) & (!g897) & (g1898) & (g2022) & (g2071)) + ((g828) & (g864) & (g897) & (!g1898) & (!g2022) & (g2071)) + ((g828) & (g864) & (g897) & (!g1898) & (g2022) & (!g2071)) + ((g828) & (g864) & (g897) & (!g1898) & (g2022) & (g2071)) + ((g828) & (g864) & (g897) & (g1898) & (!g2022) & (!g2071)) + ((g828) & (g864) & (g897) & (g1898) & (!g2022) & (g2071)) + ((g828) & (g864) & (g897) & (g1898) & (g2022) & (!g2071)) + ((g828) & (g864) & (g897) & (g1898) & (g2022) & (g2071)));
	assign g3501 = (((!g998) & (g2184)) + ((g998) & (!g2184)));
	assign g3502 = (((!g931) & (!g964) & (g3500) & (g2104) & (g2153) & (g3501)) + ((!g931) & (g964) & (!g3500) & (!g2104) & (g2153) & (g3501)) + ((!g931) & (g964) & (!g3500) & (g2104) & (g2153) & (g3501)) + ((!g931) & (g964) & (g3500) & (!g2104) & (g2153) & (g3501)) + ((!g931) & (g964) & (g3500) & (g2104) & (!g2153) & (g3501)) + ((!g931) & (g964) & (g3500) & (g2104) & (g2153) & (g3501)) + ((g931) & (!g964) & (!g3500) & (g2104) & (g2153) & (g3501)) + ((g931) & (!g964) & (g3500) & (!g2104) & (g2153) & (g3501)) + ((g931) & (!g964) & (g3500) & (g2104) & (g2153) & (g3501)) + ((g931) & (g964) & (!g3500) & (!g2104) & (g2153) & (g3501)) + ((g931) & (g964) & (!g3500) & (g2104) & (!g2153) & (g3501)) + ((g931) & (g964) & (!g3500) & (g2104) & (g2153) & (g3501)) + ((g931) & (g964) & (g3500) & (!g2104) & (!g2153) & (g3501)) + ((g931) & (g964) & (g3500) & (!g2104) & (g2153) & (g3501)) + ((g931) & (g964) & (g3500) & (g2104) & (!g2153) & (g3501)) + ((g931) & (g964) & (g3500) & (g2104) & (g2153) & (g3501)));
	assign g3503 = (((g998) & (g2184)));
	assign g3504 = (((!g1031) & (!g1065) & (!g3502) & (!g3503) & (!g2233) & (!g2267)) + ((!g1031) & (!g1065) & (!g3502) & (!g3503) & (!g2233) & (g2267)) + ((!g1031) & (!g1065) & (!g3502) & (!g3503) & (g2233) & (!g2267)) + ((!g1031) & (!g1065) & (!g3502) & (!g3503) & (g2233) & (g2267)) + ((!g1031) & (!g1065) & (!g3502) & (g3503) & (!g2233) & (!g2267)) + ((!g1031) & (!g1065) & (!g3502) & (g3503) & (!g2233) & (g2267)) + ((!g1031) & (!g1065) & (!g3502) & (g3503) & (g2233) & (!g2267)) + ((!g1031) & (!g1065) & (g3502) & (!g3503) & (!g2233) & (!g2267)) + ((!g1031) & (!g1065) & (g3502) & (!g3503) & (!g2233) & (g2267)) + ((!g1031) & (!g1065) & (g3502) & (!g3503) & (g2233) & (!g2267)) + ((!g1031) & (!g1065) & (g3502) & (g3503) & (!g2233) & (!g2267)) + ((!g1031) & (!g1065) & (g3502) & (g3503) & (!g2233) & (g2267)) + ((!g1031) & (!g1065) & (g3502) & (g3503) & (g2233) & (!g2267)) + ((!g1031) & (g1065) & (!g3502) & (!g3503) & (!g2233) & (!g2267)) + ((!g1031) & (g1065) & (!g3502) & (!g3503) & (g2233) & (!g2267)) + ((!g1031) & (g1065) & (!g3502) & (g3503) & (!g2233) & (!g2267)) + ((!g1031) & (g1065) & (g3502) & (!g3503) & (!g2233) & (!g2267)) + ((!g1031) & (g1065) & (g3502) & (g3503) & (!g2233) & (!g2267)) + ((g1031) & (!g1065) & (!g3502) & (!g3503) & (!g2233) & (!g2267)) + ((g1031) & (!g1065) & (!g3502) & (!g3503) & (!g2233) & (g2267)) + ((g1031) & (!g1065) & (!g3502) & (!g3503) & (g2233) & (!g2267)) + ((g1031) & (!g1065) & (!g3502) & (g3503) & (!g2233) & (!g2267)) + ((g1031) & (!g1065) & (!g3502) & (g3503) & (g2233) & (!g2267)) + ((g1031) & (!g1065) & (g3502) & (!g3503) & (!g2233) & (!g2267)) + ((g1031) & (!g1065) & (g3502) & (!g3503) & (g2233) & (!g2267)) + ((g1031) & (!g1065) & (g3502) & (g3503) & (!g2233) & (!g2267)) + ((g1031) & (!g1065) & (g3502) & (g3503) & (g2233) & (!g2267)) + ((g1031) & (g1065) & (!g3502) & (!g3503) & (!g2233) & (!g2267)));
	assign g3505 = (((!g1031) & (!g3502) & (!g3503) & (!g2233) & (!g5791) & (g5792)) + ((!g1031) & (!g3502) & (!g3503) & (g2233) & (!g5791) & (g5792)) + ((!g1031) & (!g3502) & (g3503) & (!g2233) & (!g5791) & (g5792)) + ((!g1031) & (!g3502) & (g3503) & (g2233) & (!g5791) & (g5792)) + ((!g1031) & (!g3502) & (g3503) & (g2233) & (g5791) & (g5792)) + ((!g1031) & (g3502) & (!g3503) & (!g2233) & (!g5791) & (g5792)) + ((!g1031) & (g3502) & (!g3503) & (g2233) & (!g5791) & (g5792)) + ((!g1031) & (g3502) & (!g3503) & (g2233) & (g5791) & (g5792)) + ((!g1031) & (g3502) & (g3503) & (!g2233) & (!g5791) & (g5792)) + ((!g1031) & (g3502) & (g3503) & (g2233) & (!g5791) & (g5792)) + ((!g1031) & (g3502) & (g3503) & (g2233) & (g5791) & (g5792)) + ((g1031) & (!g3502) & (!g3503) & (!g2233) & (!g5791) & (g5792)) + ((g1031) & (!g3502) & (!g3503) & (g2233) & (!g5791) & (g5792)) + ((g1031) & (!g3502) & (!g3503) & (g2233) & (g5791) & (g5792)) + ((g1031) & (!g3502) & (g3503) & (!g2233) & (!g5791) & (g5792)) + ((g1031) & (!g3502) & (g3503) & (!g2233) & (g5791) & (g5792)) + ((g1031) & (!g3502) & (g3503) & (g2233) & (!g5791) & (g5792)) + ((g1031) & (!g3502) & (g3503) & (g2233) & (g5791) & (g5792)) + ((g1031) & (g3502) & (!g3503) & (!g2233) & (!g5791) & (g5792)) + ((g1031) & (g3502) & (!g3503) & (!g2233) & (g5791) & (g5792)) + ((g1031) & (g3502) & (!g3503) & (g2233) & (!g5791) & (g5792)) + ((g1031) & (g3502) & (!g3503) & (g2233) & (g5791) & (g5792)) + ((g1031) & (g3502) & (g3503) & (!g2233) & (!g5791) & (g5792)) + ((g1031) & (g3502) & (g3503) & (!g2233) & (g5791) & (g5792)) + ((g1031) & (g3502) & (g3503) & (g2233) & (!g5791) & (g5792)) + ((g1031) & (g3502) & (g3503) & (g2233) & (g5791) & (g5792)));
	assign g3506 = (((g1165) & (g2399)));
	assign g3507 = (((!g1199) & (!g1236) & (!g3505) & (!g3506) & (!g2434) & (!g2533)) + ((!g1199) & (!g1236) & (!g3505) & (!g3506) & (!g2434) & (g2533)) + ((!g1199) & (!g1236) & (!g3505) & (!g3506) & (g2434) & (!g2533)) + ((!g1199) & (!g1236) & (!g3505) & (!g3506) & (g2434) & (g2533)) + ((!g1199) & (!g1236) & (!g3505) & (g3506) & (!g2434) & (!g2533)) + ((!g1199) & (!g1236) & (!g3505) & (g3506) & (!g2434) & (g2533)) + ((!g1199) & (!g1236) & (!g3505) & (g3506) & (g2434) & (!g2533)) + ((!g1199) & (!g1236) & (g3505) & (!g3506) & (!g2434) & (!g2533)) + ((!g1199) & (!g1236) & (g3505) & (!g3506) & (!g2434) & (g2533)) + ((!g1199) & (!g1236) & (g3505) & (!g3506) & (g2434) & (!g2533)) + ((!g1199) & (!g1236) & (g3505) & (g3506) & (!g2434) & (!g2533)) + ((!g1199) & (!g1236) & (g3505) & (g3506) & (!g2434) & (g2533)) + ((!g1199) & (!g1236) & (g3505) & (g3506) & (g2434) & (!g2533)) + ((!g1199) & (g1236) & (!g3505) & (!g3506) & (!g2434) & (!g2533)) + ((!g1199) & (g1236) & (!g3505) & (!g3506) & (g2434) & (!g2533)) + ((!g1199) & (g1236) & (!g3505) & (g3506) & (!g2434) & (!g2533)) + ((!g1199) & (g1236) & (g3505) & (!g3506) & (!g2434) & (!g2533)) + ((!g1199) & (g1236) & (g3505) & (g3506) & (!g2434) & (!g2533)) + ((g1199) & (!g1236) & (!g3505) & (!g3506) & (!g2434) & (!g2533)) + ((g1199) & (!g1236) & (!g3505) & (!g3506) & (!g2434) & (g2533)) + ((g1199) & (!g1236) & (!g3505) & (!g3506) & (g2434) & (!g2533)) + ((g1199) & (!g1236) & (!g3505) & (g3506) & (!g2434) & (!g2533)) + ((g1199) & (!g1236) & (!g3505) & (g3506) & (g2434) & (!g2533)) + ((g1199) & (!g1236) & (g3505) & (!g3506) & (!g2434) & (!g2533)) + ((g1199) & (!g1236) & (g3505) & (!g3506) & (g2434) & (!g2533)) + ((g1199) & (!g1236) & (g3505) & (g3506) & (!g2434) & (!g2533)) + ((g1199) & (!g1236) & (g3505) & (g3506) & (g2434) & (!g2533)) + ((g1199) & (g1236) & (!g3505) & (!g3506) & (!g2434) & (!g2533)));
	assign g3508 = (((!g1337) & (g2653)) + ((g1337) & (!g2653)));
	assign g3509 = (((!g1269) & (!g1303) & (!g3507) & (g2559) & (g2623) & (g3508)) + ((!g1269) & (g1303) & (!g3507) & (!g2559) & (g2623) & (g3508)) + ((!g1269) & (g1303) & (!g3507) & (g2559) & (!g2623) & (g3508)) + ((!g1269) & (g1303) & (!g3507) & (g2559) & (g2623) & (g3508)) + ((!g1269) & (g1303) & (g3507) & (!g2559) & (g2623) & (g3508)) + ((!g1269) & (g1303) & (g3507) & (g2559) & (g2623) & (g3508)) + ((g1269) & (!g1303) & (!g3507) & (!g2559) & (g2623) & (g3508)) + ((g1269) & (!g1303) & (!g3507) & (g2559) & (g2623) & (g3508)) + ((g1269) & (!g1303) & (g3507) & (g2559) & (g2623) & (g3508)) + ((g1269) & (g1303) & (!g3507) & (!g2559) & (!g2623) & (g3508)) + ((g1269) & (g1303) & (!g3507) & (!g2559) & (g2623) & (g3508)) + ((g1269) & (g1303) & (!g3507) & (g2559) & (!g2623) & (g3508)) + ((g1269) & (g1303) & (!g3507) & (g2559) & (g2623) & (g3508)) + ((g1269) & (g1303) & (g3507) & (!g2559) & (g2623) & (g3508)) + ((g1269) & (g1303) & (g3507) & (g2559) & (!g2623) & (g3508)) + ((g1269) & (g1303) & (g3507) & (g2559) & (g2623) & (g3508)));
	assign g3510 = (((g1337) & (g2653)));
	assign g3511 = (((!g1370) & (!g1406) & (!g3509) & (!g3510) & (!g2718) & (!g2764)) + ((!g1370) & (!g1406) & (!g3509) & (!g3510) & (!g2718) & (g2764)) + ((!g1370) & (!g1406) & (!g3509) & (!g3510) & (g2718) & (!g2764)) + ((!g1370) & (!g1406) & (!g3509) & (!g3510) & (g2718) & (g2764)) + ((!g1370) & (!g1406) & (!g3509) & (g3510) & (!g2718) & (!g2764)) + ((!g1370) & (!g1406) & (!g3509) & (g3510) & (!g2718) & (g2764)) + ((!g1370) & (!g1406) & (!g3509) & (g3510) & (g2718) & (!g2764)) + ((!g1370) & (!g1406) & (g3509) & (!g3510) & (!g2718) & (!g2764)) + ((!g1370) & (!g1406) & (g3509) & (!g3510) & (!g2718) & (g2764)) + ((!g1370) & (!g1406) & (g3509) & (!g3510) & (g2718) & (!g2764)) + ((!g1370) & (!g1406) & (g3509) & (g3510) & (!g2718) & (!g2764)) + ((!g1370) & (!g1406) & (g3509) & (g3510) & (!g2718) & (g2764)) + ((!g1370) & (!g1406) & (g3509) & (g3510) & (g2718) & (!g2764)) + ((!g1370) & (g1406) & (!g3509) & (!g3510) & (!g2718) & (!g2764)) + ((!g1370) & (g1406) & (!g3509) & (!g3510) & (g2718) & (!g2764)) + ((!g1370) & (g1406) & (!g3509) & (g3510) & (!g2718) & (!g2764)) + ((!g1370) & (g1406) & (g3509) & (!g3510) & (!g2718) & (!g2764)) + ((!g1370) & (g1406) & (g3509) & (g3510) & (!g2718) & (!g2764)) + ((g1370) & (!g1406) & (!g3509) & (!g3510) & (!g2718) & (!g2764)) + ((g1370) & (!g1406) & (!g3509) & (!g3510) & (!g2718) & (g2764)) + ((g1370) & (!g1406) & (!g3509) & (!g3510) & (g2718) & (!g2764)) + ((g1370) & (!g1406) & (!g3509) & (g3510) & (!g2718) & (!g2764)) + ((g1370) & (!g1406) & (!g3509) & (g3510) & (g2718) & (!g2764)) + ((g1370) & (!g1406) & (g3509) & (!g3510) & (!g2718) & (!g2764)) + ((g1370) & (!g1406) & (g3509) & (!g3510) & (g2718) & (!g2764)) + ((g1370) & (!g1406) & (g3509) & (g3510) & (!g2718) & (!g2764)) + ((g1370) & (!g1406) & (g3509) & (g3510) & (g2718) & (!g2764)) + ((g1370) & (g1406) & (!g3509) & (!g3510) & (!g2718) & (!g2764)));
	assign g3512 = (((!g1507) & (g2891)) + ((g1507) & (!g2891)));
	assign g3513 = (((!g1439) & (!g1473) & (!g3511) & (g2813) & (g2838) & (g3512)) + ((!g1439) & (g1473) & (!g3511) & (!g2813) & (g2838) & (g3512)) + ((!g1439) & (g1473) & (!g3511) & (g2813) & (!g2838) & (g3512)) + ((!g1439) & (g1473) & (!g3511) & (g2813) & (g2838) & (g3512)) + ((!g1439) & (g1473) & (g3511) & (!g2813) & (g2838) & (g3512)) + ((!g1439) & (g1473) & (g3511) & (g2813) & (g2838) & (g3512)) + ((g1439) & (!g1473) & (!g3511) & (!g2813) & (g2838) & (g3512)) + ((g1439) & (!g1473) & (!g3511) & (g2813) & (g2838) & (g3512)) + ((g1439) & (!g1473) & (g3511) & (g2813) & (g2838) & (g3512)) + ((g1439) & (g1473) & (!g3511) & (!g2813) & (!g2838) & (g3512)) + ((g1439) & (g1473) & (!g3511) & (!g2813) & (g2838) & (g3512)) + ((g1439) & (g1473) & (!g3511) & (g2813) & (!g2838) & (g3512)) + ((g1439) & (g1473) & (!g3511) & (g2813) & (g2838) & (g3512)) + ((g1439) & (g1473) & (g3511) & (!g2813) & (g2838) & (g3512)) + ((g1439) & (g1473) & (g3511) & (g2813) & (!g2838) & (g3512)) + ((g1439) & (g1473) & (g3511) & (g2813) & (g2838) & (g3512)));
	assign g3514 = (((g1507) & (g2891)));
	assign g3515 = (((!g1540) & (!g1577) & (!g3513) & (!g3514) & (!g2916) & (!g3009)) + ((!g1540) & (!g1577) & (!g3513) & (!g3514) & (!g2916) & (g3009)) + ((!g1540) & (!g1577) & (!g3513) & (!g3514) & (g2916) & (!g3009)) + ((!g1540) & (!g1577) & (!g3513) & (!g3514) & (g2916) & (g3009)) + ((!g1540) & (!g1577) & (!g3513) & (g3514) & (!g2916) & (!g3009)) + ((!g1540) & (!g1577) & (!g3513) & (g3514) & (!g2916) & (g3009)) + ((!g1540) & (!g1577) & (!g3513) & (g3514) & (g2916) & (!g3009)) + ((!g1540) & (!g1577) & (g3513) & (!g3514) & (!g2916) & (!g3009)) + ((!g1540) & (!g1577) & (g3513) & (!g3514) & (!g2916) & (g3009)) + ((!g1540) & (!g1577) & (g3513) & (!g3514) & (g2916) & (!g3009)) + ((!g1540) & (!g1577) & (g3513) & (g3514) & (!g2916) & (!g3009)) + ((!g1540) & (!g1577) & (g3513) & (g3514) & (!g2916) & (g3009)) + ((!g1540) & (!g1577) & (g3513) & (g3514) & (g2916) & (!g3009)) + ((!g1540) & (g1577) & (!g3513) & (!g3514) & (!g2916) & (!g3009)) + ((!g1540) & (g1577) & (!g3513) & (!g3514) & (g2916) & (!g3009)) + ((!g1540) & (g1577) & (!g3513) & (g3514) & (!g2916) & (!g3009)) + ((!g1540) & (g1577) & (g3513) & (!g3514) & (!g2916) & (!g3009)) + ((!g1540) & (g1577) & (g3513) & (g3514) & (!g2916) & (!g3009)) + ((g1540) & (!g1577) & (!g3513) & (!g3514) & (!g2916) & (!g3009)) + ((g1540) & (!g1577) & (!g3513) & (!g3514) & (!g2916) & (g3009)) + ((g1540) & (!g1577) & (!g3513) & (!g3514) & (g2916) & (!g3009)) + ((g1540) & (!g1577) & (!g3513) & (g3514) & (!g2916) & (!g3009)) + ((g1540) & (!g1577) & (!g3513) & (g3514) & (g2916) & (!g3009)) + ((g1540) & (!g1577) & (g3513) & (!g3514) & (!g2916) & (!g3009)) + ((g1540) & (!g1577) & (g3513) & (!g3514) & (g2916) & (!g3009)) + ((g1540) & (!g1577) & (g3513) & (g3514) & (!g2916) & (!g3009)) + ((g1540) & (!g1577) & (g3513) & (g3514) & (g2916) & (!g3009)) + ((g1540) & (g1577) & (!g3513) & (!g3514) & (!g2916) & (!g3009)));
	assign g3516 = (((g1914) & (!g1610) & (!g3515) & (!g3031)) + ((g1914) & (!g1610) & (g3515) & (g3031)) + ((g1914) & (g1610) & (!g3515) & (g3031)) + ((g1914) & (g1610) & (g3515) & (!g3031)));
	assign g3517 = (((!g1892) & (!g2026) & (g2062) & (!g1896) & (!g2041) & (g2068)) + ((!g1892) & (!g2026) & (g2062) & (!g1896) & (g2041) & (g2068)) + ((!g1892) & (!g2026) & (g2062) & (g1896) & (!g2041) & (g2068)) + ((!g1892) & (!g2026) & (g2062) & (g1896) & (g2041) & (g2068)) + ((!g1892) & (g2026) & (!g2062) & (!g1896) & (g2041) & (g2068)) + ((!g1892) & (g2026) & (!g2062) & (g1896) & (g2041) & (g2068)) + ((!g1892) & (g2026) & (g2062) & (!g1896) & (!g2041) & (g2068)) + ((!g1892) & (g2026) & (g2062) & (!g1896) & (g2041) & (!g2068)) + ((!g1892) & (g2026) & (g2062) & (!g1896) & (g2041) & (g2068)) + ((!g1892) & (g2026) & (g2062) & (g1896) & (!g2041) & (g2068)) + ((!g1892) & (g2026) & (g2062) & (g1896) & (g2041) & (!g2068)) + ((!g1892) & (g2026) & (g2062) & (g1896) & (g2041) & (g2068)) + ((g1892) & (!g2026) & (!g2062) & (g1896) & (g2041) & (g2068)) + ((g1892) & (!g2026) & (g2062) & (!g1896) & (!g2041) & (g2068)) + ((g1892) & (!g2026) & (g2062) & (!g1896) & (g2041) & (g2068)) + ((g1892) & (!g2026) & (g2062) & (g1896) & (!g2041) & (g2068)) + ((g1892) & (!g2026) & (g2062) & (g1896) & (g2041) & (!g2068)) + ((g1892) & (!g2026) & (g2062) & (g1896) & (g2041) & (g2068)) + ((g1892) & (g2026) & (!g2062) & (!g1896) & (g2041) & (g2068)) + ((g1892) & (g2026) & (!g2062) & (g1896) & (!g2041) & (g2068)) + ((g1892) & (g2026) & (!g2062) & (g1896) & (g2041) & (g2068)) + ((g1892) & (g2026) & (g2062) & (!g1896) & (!g2041) & (g2068)) + ((g1892) & (g2026) & (g2062) & (!g1896) & (g2041) & (!g2068)) + ((g1892) & (g2026) & (g2062) & (!g1896) & (g2041) & (g2068)) + ((g1892) & (g2026) & (g2062) & (g1896) & (!g2041) & (!g2068)) + ((g1892) & (g2026) & (g2062) & (g1896) & (!g2041) & (g2068)) + ((g1892) & (g2026) & (g2062) & (g1896) & (g2041) & (!g2068)) + ((g1892) & (g2026) & (g2062) & (g1896) & (g2041) & (g2068)));
	assign g3518 = (((!g2188) & (g2203)) + ((g2188) & (!g2203)));
	assign g3519 = (((!g2108) & (!g2144) & (g2123) & (g2150) & (g3517) & (g3518)) + ((!g2108) & (g2144) & (!g2123) & (g2150) & (!g3517) & (g3518)) + ((!g2108) & (g2144) & (!g2123) & (g2150) & (g3517) & (g3518)) + ((!g2108) & (g2144) & (g2123) & (!g2150) & (g3517) & (g3518)) + ((!g2108) & (g2144) & (g2123) & (g2150) & (!g3517) & (g3518)) + ((!g2108) & (g2144) & (g2123) & (g2150) & (g3517) & (g3518)) + ((g2108) & (!g2144) & (!g2123) & (g2150) & (g3517) & (g3518)) + ((g2108) & (!g2144) & (g2123) & (g2150) & (!g3517) & (g3518)) + ((g2108) & (!g2144) & (g2123) & (g2150) & (g3517) & (g3518)) + ((g2108) & (g2144) & (!g2123) & (!g2150) & (g3517) & (g3518)) + ((g2108) & (g2144) & (!g2123) & (g2150) & (!g3517) & (g3518)) + ((g2108) & (g2144) & (!g2123) & (g2150) & (g3517) & (g3518)) + ((g2108) & (g2144) & (g2123) & (!g2150) & (!g3517) & (g3518)) + ((g2108) & (g2144) & (g2123) & (!g2150) & (g3517) & (g3518)) + ((g2108) & (g2144) & (g2123) & (g2150) & (!g3517) & (g3518)) + ((g2108) & (g2144) & (g2123) & (g2150) & (g3517) & (g3518)));
	assign g3520 = (((g2188) & (g2203)));
	assign g3521 = (((!g2224) & (!g2271) & (!g2230) & (!g2286) & (!g3519) & (!g3520)) + ((!g2224) & (!g2271) & (!g2230) & (!g2286) & (!g3519) & (g3520)) + ((!g2224) & (!g2271) & (!g2230) & (!g2286) & (g3519) & (!g3520)) + ((!g2224) & (!g2271) & (!g2230) & (!g2286) & (g3519) & (g3520)) + ((!g2224) & (!g2271) & (!g2230) & (g2286) & (!g3519) & (!g3520)) + ((!g2224) & (!g2271) & (!g2230) & (g2286) & (!g3519) & (g3520)) + ((!g2224) & (!g2271) & (!g2230) & (g2286) & (g3519) & (!g3520)) + ((!g2224) & (!g2271) & (!g2230) & (g2286) & (g3519) & (g3520)) + ((!g2224) & (!g2271) & (g2230) & (!g2286) & (!g3519) & (!g3520)) + ((!g2224) & (!g2271) & (g2230) & (!g2286) & (!g3519) & (g3520)) + ((!g2224) & (!g2271) & (g2230) & (!g2286) & (g3519) & (!g3520)) + ((!g2224) & (!g2271) & (g2230) & (!g2286) & (g3519) & (g3520)) + ((!g2224) & (!g2271) & (g2230) & (g2286) & (!g3519) & (!g3520)) + ((!g2224) & (g2271) & (!g2230) & (!g2286) & (!g3519) & (!g3520)) + ((!g2224) & (g2271) & (!g2230) & (!g2286) & (!g3519) & (g3520)) + ((!g2224) & (g2271) & (!g2230) & (!g2286) & (g3519) & (!g3520)) + ((!g2224) & (g2271) & (!g2230) & (!g2286) & (g3519) & (g3520)) + ((!g2224) & (g2271) & (g2230) & (!g2286) & (!g3519) & (!g3520)) + ((g2224) & (!g2271) & (!g2230) & (!g2286) & (!g3519) & (!g3520)) + ((g2224) & (!g2271) & (!g2230) & (!g2286) & (!g3519) & (g3520)) + ((g2224) & (!g2271) & (!g2230) & (!g2286) & (g3519) & (!g3520)) + ((g2224) & (!g2271) & (!g2230) & (!g2286) & (g3519) & (g3520)) + ((g2224) & (!g2271) & (!g2230) & (g2286) & (!g3519) & (!g3520)) + ((g2224) & (!g2271) & (g2230) & (!g2286) & (!g3519) & (!g3520)) + ((g2224) & (!g2271) & (g2230) & (!g2286) & (!g3519) & (g3520)) + ((g2224) & (!g2271) & (g2230) & (!g2286) & (g3519) & (!g3520)) + ((g2224) & (!g2271) & (g2230) & (!g2286) & (g3519) & (g3520)) + ((g2224) & (g2271) & (!g2230) & (!g2286) & (!g3519) & (!g3520)));
	assign g3522 = (((!g2390) & (g2396)) + ((g2390) & (!g2396)));
	assign g3523 = (((!g2311) & (!g2354) & (g2317) & (g2369) & (!g3521) & (g3522)) + ((!g2311) & (g2354) & (!g2317) & (g2369) & (!g3521) & (g3522)) + ((!g2311) & (g2354) & (!g2317) & (g2369) & (g3521) & (g3522)) + ((!g2311) & (g2354) & (g2317) & (!g2369) & (!g3521) & (g3522)) + ((!g2311) & (g2354) & (g2317) & (g2369) & (!g3521) & (g3522)) + ((!g2311) & (g2354) & (g2317) & (g2369) & (g3521) & (g3522)) + ((g2311) & (!g2354) & (!g2317) & (g2369) & (!g3521) & (g3522)) + ((g2311) & (!g2354) & (g2317) & (g2369) & (!g3521) & (g3522)) + ((g2311) & (!g2354) & (g2317) & (g2369) & (g3521) & (g3522)) + ((g2311) & (g2354) & (!g2317) & (!g2369) & (!g3521) & (g3522)) + ((g2311) & (g2354) & (!g2317) & (g2369) & (!g3521) & (g3522)) + ((g2311) & (g2354) & (!g2317) & (g2369) & (g3521) & (g3522)) + ((g2311) & (g2354) & (g2317) & (!g2369) & (!g3521) & (g3522)) + ((g2311) & (g2354) & (g2317) & (!g2369) & (g3521) & (g3522)) + ((g2311) & (g2354) & (g2317) & (g2369) & (!g3521) & (g3522)) + ((g2311) & (g2354) & (g2317) & (g2369) & (g3521) & (g3522)));
	assign g3524 = (((g2390) & (g2396)));
	assign g3525 = (((!g2450) & (!g2527) & (!g2497) & (!g2531) & (!g3523) & (!g3524)) + ((!g2450) & (!g2527) & (!g2497) & (!g2531) & (!g3523) & (g3524)) + ((!g2450) & (!g2527) & (!g2497) & (!g2531) & (g3523) & (!g3524)) + ((!g2450) & (!g2527) & (!g2497) & (!g2531) & (g3523) & (g3524)) + ((!g2450) & (!g2527) & (!g2497) & (g2531) & (!g3523) & (!g3524)) + ((!g2450) & (!g2527) & (!g2497) & (g2531) & (!g3523) & (g3524)) + ((!g2450) & (!g2527) & (!g2497) & (g2531) & (g3523) & (!g3524)) + ((!g2450) & (!g2527) & (!g2497) & (g2531) & (g3523) & (g3524)) + ((!g2450) & (!g2527) & (g2497) & (!g2531) & (!g3523) & (!g3524)) + ((!g2450) & (!g2527) & (g2497) & (!g2531) & (!g3523) & (g3524)) + ((!g2450) & (!g2527) & (g2497) & (!g2531) & (g3523) & (!g3524)) + ((!g2450) & (!g2527) & (g2497) & (!g2531) & (g3523) & (g3524)) + ((!g2450) & (!g2527) & (g2497) & (g2531) & (!g3523) & (!g3524)) + ((!g2450) & (g2527) & (!g2497) & (!g2531) & (!g3523) & (!g3524)) + ((!g2450) & (g2527) & (!g2497) & (!g2531) & (!g3523) & (g3524)) + ((!g2450) & (g2527) & (!g2497) & (!g2531) & (g3523) & (!g3524)) + ((!g2450) & (g2527) & (!g2497) & (!g2531) & (g3523) & (g3524)) + ((!g2450) & (g2527) & (g2497) & (!g2531) & (!g3523) & (!g3524)) + ((g2450) & (!g2527) & (!g2497) & (!g2531) & (!g3523) & (!g3524)) + ((g2450) & (!g2527) & (!g2497) & (!g2531) & (!g3523) & (g3524)) + ((g2450) & (!g2527) & (!g2497) & (!g2531) & (g3523) & (!g3524)) + ((g2450) & (!g2527) & (!g2497) & (!g2531) & (g3523) & (g3524)) + ((g2450) & (!g2527) & (!g2497) & (g2531) & (!g3523) & (!g3524)) + ((g2450) & (!g2527) & (g2497) & (!g2531) & (!g3523) & (!g3524)) + ((g2450) & (!g2527) & (g2497) & (!g2531) & (!g3523) & (g3524)) + ((g2450) & (!g2527) & (g2497) & (!g2531) & (g3523) & (!g3524)) + ((g2450) & (!g2527) & (g2497) & (!g2531) & (g3523) & (g3524)) + ((g2450) & (g2527) & (!g2497) & (!g2531) & (!g3523) & (!g3524)));
	assign g3526 = (((!g2450) & (!g2497) & (!g3523) & (!g3524) & (!g5815) & (g5816)) + ((!g2450) & (!g2497) & (!g3523) & (g3524) & (!g5815) & (g5816)) + ((!g2450) & (!g2497) & (g3523) & (!g3524) & (!g5815) & (g5816)) + ((!g2450) & (!g2497) & (g3523) & (g3524) & (!g5815) & (g5816)) + ((!g2450) & (g2497) & (!g3523) & (!g3524) & (!g5815) & (g5816)) + ((!g2450) & (g2497) & (!g3523) & (g3524) & (!g5815) & (g5816)) + ((!g2450) & (g2497) & (!g3523) & (g3524) & (g5815) & (g5816)) + ((!g2450) & (g2497) & (g3523) & (!g3524) & (!g5815) & (g5816)) + ((!g2450) & (g2497) & (g3523) & (!g3524) & (g5815) & (g5816)) + ((!g2450) & (g2497) & (g3523) & (g3524) & (!g5815) & (g5816)) + ((!g2450) & (g2497) & (g3523) & (g3524) & (g5815) & (g5816)) + ((g2450) & (!g2497) & (!g3523) & (!g3524) & (!g5815) & (g5816)) + ((g2450) & (!g2497) & (!g3523) & (g3524) & (!g5815) & (g5816)) + ((g2450) & (!g2497) & (!g3523) & (g3524) & (g5815) & (g5816)) + ((g2450) & (!g2497) & (g3523) & (!g3524) & (!g5815) & (g5816)) + ((g2450) & (!g2497) & (g3523) & (!g3524) & (g5815) & (g5816)) + ((g2450) & (!g2497) & (g3523) & (g3524) & (!g5815) & (g5816)) + ((g2450) & (!g2497) & (g3523) & (g3524) & (g5815) & (g5816)) + ((g2450) & (g2497) & (!g3523) & (!g3524) & (!g5815) & (g5816)) + ((g2450) & (g2497) & (!g3523) & (!g3524) & (g5815) & (g5816)) + ((g2450) & (g2497) & (!g3523) & (g3524) & (!g5815) & (g5816)) + ((g2450) & (g2497) & (!g3523) & (g3524) & (g5815) & (g5816)) + ((g2450) & (g2497) & (g3523) & (!g3524) & (!g5815) & (g5816)) + ((g2450) & (g2497) & (g3523) & (!g3524) & (g5815) & (g5816)) + ((g2450) & (g2497) & (g3523) & (g3524) & (!g5815) & (g5816)) + ((g2450) & (g2497) & (g3523) & (g3524) & (g5815) & (g5816)));
	assign g3527 = (((g2657) & (g2672)));
	assign g3528 = (((!g2703) & (!g2768) & (!g2713) & (!g2783) & (!g3526) & (!g3527)) + ((!g2703) & (!g2768) & (!g2713) & (!g2783) & (!g3526) & (g3527)) + ((!g2703) & (!g2768) & (!g2713) & (!g2783) & (g3526) & (!g3527)) + ((!g2703) & (!g2768) & (!g2713) & (!g2783) & (g3526) & (g3527)) + ((!g2703) & (!g2768) & (!g2713) & (g2783) & (!g3526) & (!g3527)) + ((!g2703) & (!g2768) & (!g2713) & (g2783) & (!g3526) & (g3527)) + ((!g2703) & (!g2768) & (!g2713) & (g2783) & (g3526) & (!g3527)) + ((!g2703) & (!g2768) & (!g2713) & (g2783) & (g3526) & (g3527)) + ((!g2703) & (!g2768) & (g2713) & (!g2783) & (!g3526) & (!g3527)) + ((!g2703) & (!g2768) & (g2713) & (!g2783) & (!g3526) & (g3527)) + ((!g2703) & (!g2768) & (g2713) & (!g2783) & (g3526) & (!g3527)) + ((!g2703) & (!g2768) & (g2713) & (!g2783) & (g3526) & (g3527)) + ((!g2703) & (!g2768) & (g2713) & (g2783) & (!g3526) & (!g3527)) + ((!g2703) & (g2768) & (!g2713) & (!g2783) & (!g3526) & (!g3527)) + ((!g2703) & (g2768) & (!g2713) & (!g2783) & (!g3526) & (g3527)) + ((!g2703) & (g2768) & (!g2713) & (!g2783) & (g3526) & (!g3527)) + ((!g2703) & (g2768) & (!g2713) & (!g2783) & (g3526) & (g3527)) + ((!g2703) & (g2768) & (g2713) & (!g2783) & (!g3526) & (!g3527)) + ((g2703) & (!g2768) & (!g2713) & (!g2783) & (!g3526) & (!g3527)) + ((g2703) & (!g2768) & (!g2713) & (!g2783) & (!g3526) & (g3527)) + ((g2703) & (!g2768) & (!g2713) & (!g2783) & (g3526) & (!g3527)) + ((g2703) & (!g2768) & (!g2713) & (!g2783) & (g3526) & (g3527)) + ((g2703) & (!g2768) & (!g2713) & (g2783) & (!g3526) & (!g3527)) + ((g2703) & (!g2768) & (g2713) & (!g2783) & (!g3526) & (!g3527)) + ((g2703) & (!g2768) & (g2713) & (!g2783) & (!g3526) & (g3527)) + ((g2703) & (!g2768) & (g2713) & (!g2783) & (g3526) & (!g3527)) + ((g2703) & (!g2768) & (g2713) & (!g2783) & (g3526) & (g3527)) + ((g2703) & (g2768) & (!g2713) & (!g2783) & (!g3526) & (!g3527)));
	assign g3529 = (((!g2885) & (g2889)) + ((g2885) & (!g2889)));
	assign g3530 = (((!g2804) & (!g2845) & (g2810) & (g2868) & (!g3528) & (g3529)) + ((!g2804) & (g2845) & (!g2810) & (g2868) & (!g3528) & (g3529)) + ((!g2804) & (g2845) & (!g2810) & (g2868) & (g3528) & (g3529)) + ((!g2804) & (g2845) & (g2810) & (!g2868) & (!g3528) & (g3529)) + ((!g2804) & (g2845) & (g2810) & (g2868) & (!g3528) & (g3529)) + ((!g2804) & (g2845) & (g2810) & (g2868) & (g3528) & (g3529)) + ((g2804) & (!g2845) & (!g2810) & (g2868) & (!g3528) & (g3529)) + ((g2804) & (!g2845) & (g2810) & (g2868) & (!g3528) & (g3529)) + ((g2804) & (!g2845) & (g2810) & (g2868) & (g3528) & (g3529)) + ((g2804) & (g2845) & (!g2810) & (!g2868) & (!g3528) & (g3529)) + ((g2804) & (g2845) & (!g2810) & (g2868) & (!g3528) & (g3529)) + ((g2804) & (g2845) & (!g2810) & (g2868) & (g3528) & (g3529)) + ((g2804) & (g2845) & (g2810) & (!g2868) & (!g3528) & (g3529)) + ((g2804) & (g2845) & (g2810) & (!g2868) & (g3528) & (g3529)) + ((g2804) & (g2845) & (g2810) & (g2868) & (!g3528) & (g3529)) + ((g2804) & (g2845) & (g2810) & (g2868) & (g3528) & (g3529)));
	assign g3531 = (((g2885) & (g2889)));
	assign g3532 = (((!g2932) & (!g3003) & (!g2979) & (!g3007) & (!g3530) & (!g3531)) + ((!g2932) & (!g3003) & (!g2979) & (!g3007) & (!g3530) & (g3531)) + ((!g2932) & (!g3003) & (!g2979) & (!g3007) & (g3530) & (!g3531)) + ((!g2932) & (!g3003) & (!g2979) & (!g3007) & (g3530) & (g3531)) + ((!g2932) & (!g3003) & (!g2979) & (g3007) & (!g3530) & (!g3531)) + ((!g2932) & (!g3003) & (!g2979) & (g3007) & (!g3530) & (g3531)) + ((!g2932) & (!g3003) & (!g2979) & (g3007) & (g3530) & (!g3531)) + ((!g2932) & (!g3003) & (!g2979) & (g3007) & (g3530) & (g3531)) + ((!g2932) & (!g3003) & (g2979) & (!g3007) & (!g3530) & (!g3531)) + ((!g2932) & (!g3003) & (g2979) & (!g3007) & (!g3530) & (g3531)) + ((!g2932) & (!g3003) & (g2979) & (!g3007) & (g3530) & (!g3531)) + ((!g2932) & (!g3003) & (g2979) & (!g3007) & (g3530) & (g3531)) + ((!g2932) & (!g3003) & (g2979) & (g3007) & (!g3530) & (!g3531)) + ((!g2932) & (g3003) & (!g2979) & (!g3007) & (!g3530) & (!g3531)) + ((!g2932) & (g3003) & (!g2979) & (!g3007) & (!g3530) & (g3531)) + ((!g2932) & (g3003) & (!g2979) & (!g3007) & (g3530) & (!g3531)) + ((!g2932) & (g3003) & (!g2979) & (!g3007) & (g3530) & (g3531)) + ((!g2932) & (g3003) & (g2979) & (!g3007) & (!g3530) & (!g3531)) + ((g2932) & (!g3003) & (!g2979) & (!g3007) & (!g3530) & (!g3531)) + ((g2932) & (!g3003) & (!g2979) & (!g3007) & (!g3530) & (g3531)) + ((g2932) & (!g3003) & (!g2979) & (!g3007) & (g3530) & (!g3531)) + ((g2932) & (!g3003) & (!g2979) & (!g3007) & (g3530) & (g3531)) + ((g2932) & (!g3003) & (!g2979) & (g3007) & (!g3530) & (!g3531)) + ((g2932) & (!g3003) & (g2979) & (!g3007) & (!g3530) & (!g3531)) + ((g2932) & (!g3003) & (g2979) & (!g3007) & (!g3530) & (g3531)) + ((g2932) & (!g3003) & (g2979) & (!g3007) & (g3530) & (!g3531)) + ((g2932) & (!g3003) & (g2979) & (!g3007) & (g3530) & (g3531)) + ((g2932) & (g3003) & (!g2979) & (!g3007) & (!g3530) & (!g3531)));
	assign g3533 = (((!g1914) & (!g3038) & (!g3061) & (!g3532)) + ((!g1914) & (!g3038) & (g3061) & (g3532)) + ((!g1914) & (g3038) & (!g3061) & (g3532)) + ((!g1914) & (g3038) & (g3061) & (!g3532)));
	assign g3534 = (((!g830) & (!g1890) & (!g3516) & (!g3533) & (key[32])) + ((!g830) & (!g1890) & (!g3516) & (g3533) & (key[32])) + ((!g830) & (!g1890) & (g3516) & (!g3533) & (key[32])) + ((!g830) & (!g1890) & (g3516) & (g3533) & (key[32])) + ((!g830) & (g1890) & (!g3516) & (!g3533) & (key[32])) + ((!g830) & (g1890) & (!g3516) & (g3533) & (key[32])) + ((!g830) & (g1890) & (g3516) & (!g3533) & (key[32])) + ((!g830) & (g1890) & (g3516) & (g3533) & (key[32])) + ((g830) & (!g1890) & (!g3516) & (g3533) & (!key[32])) + ((g830) & (!g1890) & (!g3516) & (g3533) & (key[32])) + ((g830) & (!g1890) & (g3516) & (!g3533) & (!key[32])) + ((g830) & (!g1890) & (g3516) & (!g3533) & (key[32])) + ((g830) & (!g1890) & (g3516) & (g3533) & (!key[32])) + ((g830) & (!g1890) & (g3516) & (g3533) & (key[32])) + ((g830) & (g1890) & (!g3516) & (!g3533) & (!key[32])) + ((g830) & (g1890) & (!g3516) & (!g3533) & (key[32])));
	assign g3535 = (((!g1884) & (!g1977) & (g1979) & (!g1900) & (!g2028) & (g2074)) + ((!g1884) & (!g1977) & (g1979) & (!g1900) & (g2028) & (g2074)) + ((!g1884) & (!g1977) & (g1979) & (g1900) & (!g2028) & (g2074)) + ((!g1884) & (!g1977) & (g1979) & (g1900) & (g2028) & (g2074)) + ((!g1884) & (g1977) & (!g1979) & (!g1900) & (g2028) & (g2074)) + ((!g1884) & (g1977) & (!g1979) & (g1900) & (g2028) & (g2074)) + ((!g1884) & (g1977) & (g1979) & (!g1900) & (!g2028) & (g2074)) + ((!g1884) & (g1977) & (g1979) & (!g1900) & (g2028) & (!g2074)) + ((!g1884) & (g1977) & (g1979) & (!g1900) & (g2028) & (g2074)) + ((!g1884) & (g1977) & (g1979) & (g1900) & (!g2028) & (g2074)) + ((!g1884) & (g1977) & (g1979) & (g1900) & (g2028) & (!g2074)) + ((!g1884) & (g1977) & (g1979) & (g1900) & (g2028) & (g2074)) + ((g1884) & (!g1977) & (!g1979) & (g1900) & (g2028) & (g2074)) + ((g1884) & (!g1977) & (g1979) & (!g1900) & (!g2028) & (g2074)) + ((g1884) & (!g1977) & (g1979) & (!g1900) & (g2028) & (g2074)) + ((g1884) & (!g1977) & (g1979) & (g1900) & (!g2028) & (g2074)) + ((g1884) & (!g1977) & (g1979) & (g1900) & (g2028) & (!g2074)) + ((g1884) & (!g1977) & (g1979) & (g1900) & (g2028) & (g2074)) + ((g1884) & (g1977) & (!g1979) & (!g1900) & (g2028) & (g2074)) + ((g1884) & (g1977) & (!g1979) & (g1900) & (!g2028) & (g2074)) + ((g1884) & (g1977) & (!g1979) & (g1900) & (g2028) & (g2074)) + ((g1884) & (g1977) & (g1979) & (!g1900) & (!g2028) & (g2074)) + ((g1884) & (g1977) & (g1979) & (!g1900) & (g2028) & (!g2074)) + ((g1884) & (g1977) & (g1979) & (!g1900) & (g2028) & (g2074)) + ((g1884) & (g1977) & (g1979) & (g1900) & (!g2028) & (!g2074)) + ((g1884) & (g1977) & (g1979) & (g1900) & (!g2028) & (g2074)) + ((g1884) & (g1977) & (g1979) & (g1900) & (g2028) & (!g2074)) + ((g1884) & (g1977) & (g1979) & (g1900) & (g2028) & (g2074)));
	assign g3536 = (((!g1986) & (g2190)) + ((g1986) & (!g2190)));
	assign g3537 = (((!g1982) & (!g1984) & (g3535) & (g2110) & (g2156) & (g3536)) + ((!g1982) & (g1984) & (!g3535) & (!g2110) & (g2156) & (g3536)) + ((!g1982) & (g1984) & (!g3535) & (g2110) & (g2156) & (g3536)) + ((!g1982) & (g1984) & (g3535) & (!g2110) & (g2156) & (g3536)) + ((!g1982) & (g1984) & (g3535) & (g2110) & (!g2156) & (g3536)) + ((!g1982) & (g1984) & (g3535) & (g2110) & (g2156) & (g3536)) + ((g1982) & (!g1984) & (!g3535) & (g2110) & (g2156) & (g3536)) + ((g1982) & (!g1984) & (g3535) & (!g2110) & (g2156) & (g3536)) + ((g1982) & (!g1984) & (g3535) & (g2110) & (g2156) & (g3536)) + ((g1982) & (g1984) & (!g3535) & (!g2110) & (g2156) & (g3536)) + ((g1982) & (g1984) & (!g3535) & (g2110) & (!g2156) & (g3536)) + ((g1982) & (g1984) & (!g3535) & (g2110) & (g2156) & (g3536)) + ((g1982) & (g1984) & (g3535) & (!g2110) & (!g2156) & (g3536)) + ((g1982) & (g1984) & (g3535) & (!g2110) & (g2156) & (g3536)) + ((g1982) & (g1984) & (g3535) & (g2110) & (!g2156) & (g3536)) + ((g1982) & (g1984) & (g3535) & (g2110) & (g2156) & (g3536)));
	assign g3538 = (((g1986) & (g2190)));
	assign g3539 = (((!g1991) & (!g1993) & (!g3537) & (g3538) & (g2236) & (g2273)) + ((!g1991) & (!g1993) & (g3537) & (!g3538) & (g2236) & (g2273)) + ((!g1991) & (!g1993) & (g3537) & (g3538) & (g2236) & (g2273)) + ((!g1991) & (g1993) & (!g3537) & (!g3538) & (!g2236) & (g2273)) + ((!g1991) & (g1993) & (!g3537) & (!g3538) & (g2236) & (g2273)) + ((!g1991) & (g1993) & (!g3537) & (g3538) & (!g2236) & (g2273)) + ((!g1991) & (g1993) & (!g3537) & (g3538) & (g2236) & (!g2273)) + ((!g1991) & (g1993) & (!g3537) & (g3538) & (g2236) & (g2273)) + ((!g1991) & (g1993) & (g3537) & (!g3538) & (!g2236) & (g2273)) + ((!g1991) & (g1993) & (g3537) & (!g3538) & (g2236) & (!g2273)) + ((!g1991) & (g1993) & (g3537) & (!g3538) & (g2236) & (g2273)) + ((!g1991) & (g1993) & (g3537) & (g3538) & (!g2236) & (g2273)) + ((!g1991) & (g1993) & (g3537) & (g3538) & (g2236) & (!g2273)) + ((!g1991) & (g1993) & (g3537) & (g3538) & (g2236) & (g2273)) + ((g1991) & (!g1993) & (!g3537) & (!g3538) & (g2236) & (g2273)) + ((g1991) & (!g1993) & (!g3537) & (g3538) & (!g2236) & (g2273)) + ((g1991) & (!g1993) & (!g3537) & (g3538) & (g2236) & (g2273)) + ((g1991) & (!g1993) & (g3537) & (!g3538) & (!g2236) & (g2273)) + ((g1991) & (!g1993) & (g3537) & (!g3538) & (g2236) & (g2273)) + ((g1991) & (!g1993) & (g3537) & (g3538) & (!g2236) & (g2273)) + ((g1991) & (!g1993) & (g3537) & (g3538) & (g2236) & (g2273)) + ((g1991) & (g1993) & (!g3537) & (!g3538) & (!g2236) & (g2273)) + ((g1991) & (g1993) & (!g3537) & (!g3538) & (g2236) & (!g2273)) + ((g1991) & (g1993) & (!g3537) & (!g3538) & (g2236) & (g2273)) + ((g1991) & (g1993) & (!g3537) & (g3538) & (!g2236) & (!g2273)) + ((g1991) & (g1993) & (!g3537) & (g3538) & (!g2236) & (g2273)) + ((g1991) & (g1993) & (!g3537) & (g3538) & (g2236) & (!g2273)) + ((g1991) & (g1993) & (!g3537) & (g3538) & (g2236) & (g2273)) + ((g1991) & (g1993) & (g3537) & (!g3538) & (!g2236) & (!g2273)) + ((g1991) & (g1993) & (g3537) & (!g3538) & (!g2236) & (g2273)) + ((g1991) & (g1993) & (g3537) & (!g3538) & (g2236) & (!g2273)) + ((g1991) & (g1993) & (g3537) & (!g3538) & (g2236) & (g2273)) + ((g1991) & (g1993) & (g3537) & (g3538) & (!g2236) & (!g2273)) + ((g1991) & (g1993) & (g3537) & (g3538) & (!g2236) & (g2273)) + ((g1991) & (g1993) & (g3537) & (g3538) & (g2236) & (!g2273)) + ((g1991) & (g1993) & (g3537) & (g3538) & (g2236) & (g2273)));
	assign g3540 = (((!g1991) & (!g3537) & (!g3538) & (!g2236) & (!g5830) & (g5831)) + ((!g1991) & (!g3537) & (!g3538) & (g2236) & (!g5830) & (g5831)) + ((!g1991) & (!g3537) & (g3538) & (!g2236) & (!g5830) & (g5831)) + ((!g1991) & (!g3537) & (g3538) & (g2236) & (!g5830) & (g5831)) + ((!g1991) & (!g3537) & (g3538) & (g2236) & (g5830) & (g5831)) + ((!g1991) & (g3537) & (!g3538) & (!g2236) & (!g5830) & (g5831)) + ((!g1991) & (g3537) & (!g3538) & (g2236) & (!g5830) & (g5831)) + ((!g1991) & (g3537) & (!g3538) & (g2236) & (g5830) & (g5831)) + ((!g1991) & (g3537) & (g3538) & (!g2236) & (!g5830) & (g5831)) + ((!g1991) & (g3537) & (g3538) & (g2236) & (!g5830) & (g5831)) + ((!g1991) & (g3537) & (g3538) & (g2236) & (g5830) & (g5831)) + ((g1991) & (!g3537) & (!g3538) & (!g2236) & (!g5830) & (g5831)) + ((g1991) & (!g3537) & (!g3538) & (g2236) & (!g5830) & (g5831)) + ((g1991) & (!g3537) & (!g3538) & (g2236) & (g5830) & (g5831)) + ((g1991) & (!g3537) & (g3538) & (!g2236) & (!g5830) & (g5831)) + ((g1991) & (!g3537) & (g3538) & (!g2236) & (g5830) & (g5831)) + ((g1991) & (!g3537) & (g3538) & (g2236) & (!g5830) & (g5831)) + ((g1991) & (!g3537) & (g3538) & (g2236) & (g5830) & (g5831)) + ((g1991) & (g3537) & (!g3538) & (!g2236) & (!g5830) & (g5831)) + ((g1991) & (g3537) & (!g3538) & (!g2236) & (g5830) & (g5831)) + ((g1991) & (g3537) & (!g3538) & (g2236) & (!g5830) & (g5831)) + ((g1991) & (g3537) & (!g3538) & (g2236) & (g5830) & (g5831)) + ((g1991) & (g3537) & (g3538) & (!g2236) & (!g5830) & (g5831)) + ((g1991) & (g3537) & (g3538) & (!g2236) & (g5830) & (g5831)) + ((g1991) & (g3537) & (g3538) & (g2236) & (!g5830) & (g5831)) + ((g1991) & (g3537) & (g3538) & (g2236) & (g5830) & (g5831)));
	assign g3541 = (((g2001) & (g2402)));
	assign g3542 = (((!g2003) & (!g2005) & (!g3540) & (g3541) & (g2456) & (g2535)) + ((!g2003) & (!g2005) & (g3540) & (!g3541) & (g2456) & (g2535)) + ((!g2003) & (!g2005) & (g3540) & (g3541) & (g2456) & (g2535)) + ((!g2003) & (g2005) & (!g3540) & (!g3541) & (!g2456) & (g2535)) + ((!g2003) & (g2005) & (!g3540) & (!g3541) & (g2456) & (g2535)) + ((!g2003) & (g2005) & (!g3540) & (g3541) & (!g2456) & (g2535)) + ((!g2003) & (g2005) & (!g3540) & (g3541) & (g2456) & (!g2535)) + ((!g2003) & (g2005) & (!g3540) & (g3541) & (g2456) & (g2535)) + ((!g2003) & (g2005) & (g3540) & (!g3541) & (!g2456) & (g2535)) + ((!g2003) & (g2005) & (g3540) & (!g3541) & (g2456) & (!g2535)) + ((!g2003) & (g2005) & (g3540) & (!g3541) & (g2456) & (g2535)) + ((!g2003) & (g2005) & (g3540) & (g3541) & (!g2456) & (g2535)) + ((!g2003) & (g2005) & (g3540) & (g3541) & (g2456) & (!g2535)) + ((!g2003) & (g2005) & (g3540) & (g3541) & (g2456) & (g2535)) + ((g2003) & (!g2005) & (!g3540) & (!g3541) & (g2456) & (g2535)) + ((g2003) & (!g2005) & (!g3540) & (g3541) & (!g2456) & (g2535)) + ((g2003) & (!g2005) & (!g3540) & (g3541) & (g2456) & (g2535)) + ((g2003) & (!g2005) & (g3540) & (!g3541) & (!g2456) & (g2535)) + ((g2003) & (!g2005) & (g3540) & (!g3541) & (g2456) & (g2535)) + ((g2003) & (!g2005) & (g3540) & (g3541) & (!g2456) & (g2535)) + ((g2003) & (!g2005) & (g3540) & (g3541) & (g2456) & (g2535)) + ((g2003) & (g2005) & (!g3540) & (!g3541) & (!g2456) & (g2535)) + ((g2003) & (g2005) & (!g3540) & (!g3541) & (g2456) & (!g2535)) + ((g2003) & (g2005) & (!g3540) & (!g3541) & (g2456) & (g2535)) + ((g2003) & (g2005) & (!g3540) & (g3541) & (!g2456) & (!g2535)) + ((g2003) & (g2005) & (!g3540) & (g3541) & (!g2456) & (g2535)) + ((g2003) & (g2005) & (!g3540) & (g3541) & (g2456) & (!g2535)) + ((g2003) & (g2005) & (!g3540) & (g3541) & (g2456) & (g2535)) + ((g2003) & (g2005) & (g3540) & (!g3541) & (!g2456) & (!g2535)) + ((g2003) & (g2005) & (g3540) & (!g3541) & (!g2456) & (g2535)) + ((g2003) & (g2005) & (g3540) & (!g3541) & (g2456) & (!g2535)) + ((g2003) & (g2005) & (g3540) & (!g3541) & (g2456) & (g2535)) + ((g2003) & (g2005) & (g3540) & (g3541) & (!g2456) & (!g2535)) + ((g2003) & (g2005) & (g3540) & (g3541) & (!g2456) & (g2535)) + ((g2003) & (g2005) & (g3540) & (g3541) & (g2456) & (!g2535)) + ((g2003) & (g2005) & (g3540) & (g3541) & (g2456) & (g2535)));
	assign g3543 = (((!g2011) & (g3542) & (g2569)) + ((g2011) & (!g3542) & (g2569)) + ((g2011) & (g3542) & (!g2569)) + ((g2011) & (g3542) & (g2569)));
	assign g3544 = (((!g1890) & (!g1939) & (g1941) & (!g1894) & (!g2034) & (g2065)) + ((!g1890) & (!g1939) & (g1941) & (!g1894) & (g2034) & (g2065)) + ((!g1890) & (!g1939) & (g1941) & (g1894) & (!g2034) & (g2065)) + ((!g1890) & (!g1939) & (g1941) & (g1894) & (g2034) & (g2065)) + ((!g1890) & (g1939) & (!g1941) & (!g1894) & (g2034) & (g2065)) + ((!g1890) & (g1939) & (!g1941) & (g1894) & (g2034) & (g2065)) + ((!g1890) & (g1939) & (g1941) & (!g1894) & (!g2034) & (g2065)) + ((!g1890) & (g1939) & (g1941) & (!g1894) & (g2034) & (!g2065)) + ((!g1890) & (g1939) & (g1941) & (!g1894) & (g2034) & (g2065)) + ((!g1890) & (g1939) & (g1941) & (g1894) & (!g2034) & (g2065)) + ((!g1890) & (g1939) & (g1941) & (g1894) & (g2034) & (!g2065)) + ((!g1890) & (g1939) & (g1941) & (g1894) & (g2034) & (g2065)) + ((g1890) & (!g1939) & (!g1941) & (g1894) & (g2034) & (g2065)) + ((g1890) & (!g1939) & (g1941) & (!g1894) & (!g2034) & (g2065)) + ((g1890) & (!g1939) & (g1941) & (!g1894) & (g2034) & (g2065)) + ((g1890) & (!g1939) & (g1941) & (g1894) & (!g2034) & (g2065)) + ((g1890) & (!g1939) & (g1941) & (g1894) & (g2034) & (!g2065)) + ((g1890) & (!g1939) & (g1941) & (g1894) & (g2034) & (g2065)) + ((g1890) & (g1939) & (!g1941) & (!g1894) & (g2034) & (g2065)) + ((g1890) & (g1939) & (!g1941) & (g1894) & (!g2034) & (g2065)) + ((g1890) & (g1939) & (!g1941) & (g1894) & (g2034) & (g2065)) + ((g1890) & (g1939) & (g1941) & (!g1894) & (!g2034) & (g2065)) + ((g1890) & (g1939) & (g1941) & (!g1894) & (g2034) & (!g2065)) + ((g1890) & (g1939) & (g1941) & (!g1894) & (g2034) & (g2065)) + ((g1890) & (g1939) & (g1941) & (g1894) & (!g2034) & (!g2065)) + ((g1890) & (g1939) & (g1941) & (g1894) & (!g2034) & (g2065)) + ((g1890) & (g1939) & (g1941) & (g1894) & (g2034) & (!g2065)) + ((g1890) & (g1939) & (g1941) & (g1894) & (g2034) & (g2065)));
	assign g3545 = (((!g1948) & (g2196)) + ((g1948) & (!g2196)));
	assign g3546 = (((!g1944) & (!g1946) & (g2116) & (g2147) & (g3544) & (g3545)) + ((!g1944) & (g1946) & (!g2116) & (g2147) & (!g3544) & (g3545)) + ((!g1944) & (g1946) & (!g2116) & (g2147) & (g3544) & (g3545)) + ((!g1944) & (g1946) & (g2116) & (!g2147) & (g3544) & (g3545)) + ((!g1944) & (g1946) & (g2116) & (g2147) & (!g3544) & (g3545)) + ((!g1944) & (g1946) & (g2116) & (g2147) & (g3544) & (g3545)) + ((g1944) & (!g1946) & (!g2116) & (g2147) & (g3544) & (g3545)) + ((g1944) & (!g1946) & (g2116) & (g2147) & (!g3544) & (g3545)) + ((g1944) & (!g1946) & (g2116) & (g2147) & (g3544) & (g3545)) + ((g1944) & (g1946) & (!g2116) & (!g2147) & (g3544) & (g3545)) + ((g1944) & (g1946) & (!g2116) & (g2147) & (!g3544) & (g3545)) + ((g1944) & (g1946) & (!g2116) & (g2147) & (g3544) & (g3545)) + ((g1944) & (g1946) & (g2116) & (!g2147) & (!g3544) & (g3545)) + ((g1944) & (g1946) & (g2116) & (!g2147) & (g3544) & (g3545)) + ((g1944) & (g1946) & (g2116) & (g2147) & (!g3544) & (g3545)) + ((g1944) & (g1946) & (g2116) & (g2147) & (g3544) & (g3545)));
	assign g3547 = (((g1948) & (g2196)));
	assign g3548 = (((!g1953) & (!g1955) & (!g2227) & (!g2279) & (!g3546) & (!g3547)) + ((!g1953) & (!g1955) & (!g2227) & (!g2279) & (!g3546) & (g3547)) + ((!g1953) & (!g1955) & (!g2227) & (!g2279) & (g3546) & (!g3547)) + ((!g1953) & (!g1955) & (!g2227) & (!g2279) & (g3546) & (g3547)) + ((!g1953) & (!g1955) & (!g2227) & (g2279) & (!g3546) & (!g3547)) + ((!g1953) & (!g1955) & (!g2227) & (g2279) & (!g3546) & (g3547)) + ((!g1953) & (!g1955) & (!g2227) & (g2279) & (g3546) & (!g3547)) + ((!g1953) & (!g1955) & (!g2227) & (g2279) & (g3546) & (g3547)) + ((!g1953) & (!g1955) & (g2227) & (!g2279) & (!g3546) & (!g3547)) + ((!g1953) & (!g1955) & (g2227) & (!g2279) & (!g3546) & (g3547)) + ((!g1953) & (!g1955) & (g2227) & (!g2279) & (g3546) & (!g3547)) + ((!g1953) & (!g1955) & (g2227) & (!g2279) & (g3546) & (g3547)) + ((!g1953) & (!g1955) & (g2227) & (g2279) & (!g3546) & (!g3547)) + ((!g1953) & (g1955) & (!g2227) & (!g2279) & (!g3546) & (!g3547)) + ((!g1953) & (g1955) & (!g2227) & (!g2279) & (!g3546) & (g3547)) + ((!g1953) & (g1955) & (!g2227) & (!g2279) & (g3546) & (!g3547)) + ((!g1953) & (g1955) & (!g2227) & (!g2279) & (g3546) & (g3547)) + ((!g1953) & (g1955) & (g2227) & (!g2279) & (!g3546) & (!g3547)) + ((g1953) & (!g1955) & (!g2227) & (!g2279) & (!g3546) & (!g3547)) + ((g1953) & (!g1955) & (!g2227) & (!g2279) & (!g3546) & (g3547)) + ((g1953) & (!g1955) & (!g2227) & (!g2279) & (g3546) & (!g3547)) + ((g1953) & (!g1955) & (!g2227) & (!g2279) & (g3546) & (g3547)) + ((g1953) & (!g1955) & (!g2227) & (g2279) & (!g3546) & (!g3547)) + ((g1953) & (!g1955) & (g2227) & (!g2279) & (!g3546) & (!g3547)) + ((g1953) & (!g1955) & (g2227) & (!g2279) & (!g3546) & (g3547)) + ((g1953) & (!g1955) & (g2227) & (!g2279) & (g3546) & (!g3547)) + ((g1953) & (!g1955) & (g2227) & (!g2279) & (g3546) & (g3547)) + ((g1953) & (g1955) & (!g2227) & (!g2279) & (!g3546) & (!g3547)));
	assign g3549 = (((!g1958) & (!g1960) & (g2314) & (g2362) & (!g3548)) + ((!g1958) & (g1960) & (!g2314) & (g2362) & (!g3548)) + ((!g1958) & (g1960) & (!g2314) & (g2362) & (g3548)) + ((!g1958) & (g1960) & (g2314) & (!g2362) & (!g3548)) + ((!g1958) & (g1960) & (g2314) & (g2362) & (!g3548)) + ((!g1958) & (g1960) & (g2314) & (g2362) & (g3548)) + ((g1958) & (!g1960) & (!g2314) & (g2362) & (!g3548)) + ((g1958) & (!g1960) & (g2314) & (g2362) & (!g3548)) + ((g1958) & (!g1960) & (g2314) & (g2362) & (g3548)) + ((g1958) & (g1960) & (!g2314) & (!g2362) & (!g3548)) + ((g1958) & (g1960) & (!g2314) & (g2362) & (!g3548)) + ((g1958) & (g1960) & (!g2314) & (g2362) & (g3548)) + ((g1958) & (g1960) & (g2314) & (!g2362) & (!g3548)) + ((g1958) & (g1960) & (g2314) & (!g2362) & (g3548)) + ((g1958) & (g1960) & (g2314) & (g2362) & (!g3548)) + ((g1958) & (g1960) & (g2314) & (g2362) & (g3548)));
	assign g3550 = (((!g1969) & (g2529)) + ((g1969) & (!g2529)));
	assign g3551 = (((!g1962) & (!g1967) & (g2393) & (g2474) & (g3549) & (g3550)) + ((!g1962) & (g1967) & (!g2393) & (g2474) & (!g3549) & (g3550)) + ((!g1962) & (g1967) & (!g2393) & (g2474) & (g3549) & (g3550)) + ((!g1962) & (g1967) & (g2393) & (!g2474) & (g3549) & (g3550)) + ((!g1962) & (g1967) & (g2393) & (g2474) & (!g3549) & (g3550)) + ((!g1962) & (g1967) & (g2393) & (g2474) & (g3549) & (g3550)) + ((g1962) & (!g1967) & (!g2393) & (g2474) & (g3549) & (g3550)) + ((g1962) & (!g1967) & (g2393) & (g2474) & (!g3549) & (g3550)) + ((g1962) & (!g1967) & (g2393) & (g2474) & (g3549) & (g3550)) + ((g1962) & (g1967) & (!g2393) & (!g2474) & (g3549) & (g3550)) + ((g1962) & (g1967) & (!g2393) & (g2474) & (!g3549) & (g3550)) + ((g1962) & (g1967) & (!g2393) & (g2474) & (g3549) & (g3550)) + ((g1962) & (g1967) & (g2393) & (!g2474) & (!g3549) & (g3550)) + ((g1962) & (g1967) & (g2393) & (!g2474) & (g3549) & (g3550)) + ((g1962) & (g1967) & (g2393) & (g2474) & (!g3549) & (g3550)) + ((g1962) & (g1967) & (g2393) & (g2474) & (g3549) & (g3550)));
	assign g3552 = (((g1969) & (g2529)));
	assign g3553 = (((!g3551) & (!g3552)));
	assign g3554 = (((!g1972) & (!g1975) & (!g2578) & (g2617) & (!g3553)) + ((!g1972) & (!g1975) & (!g2578) & (g2617) & (g3553)) + ((!g1972) & (!g1975) & (g2578) & (!g2617) & (!g3553)) + ((!g1972) & (!g1975) & (g2578) & (g2617) & (g3553)) + ((!g1972) & (g1975) & (!g2578) & (!g2617) & (!g3553)) + ((!g1972) & (g1975) & (!g2578) & (!g2617) & (g3553)) + ((!g1972) & (g1975) & (g2578) & (!g2617) & (g3553)) + ((!g1972) & (g1975) & (g2578) & (g2617) & (!g3553)) + ((g1972) & (!g1975) & (!g2578) & (!g2617) & (!g3553)) + ((g1972) & (!g1975) & (!g2578) & (g2617) & (g3553)) + ((g1972) & (!g1975) & (g2578) & (!g2617) & (!g3553)) + ((g1972) & (!g1975) & (g2578) & (!g2617) & (g3553)) + ((g1972) & (g1975) & (!g2578) & (!g2617) & (g3553)) + ((g1972) & (g1975) & (!g2578) & (g2617) & (!g3553)) + ((g1972) & (g1975) & (g2578) & (g2617) & (!g3553)) + ((g1972) & (g1975) & (g2578) & (g2617) & (g3553)));
	assign g3555 = (((!g1886) & (!g2032) & (g2055) & (!g1902) & (!g2036) & (g2077)) + ((!g1886) & (!g2032) & (g2055) & (!g1902) & (g2036) & (g2077)) + ((!g1886) & (!g2032) & (g2055) & (g1902) & (!g2036) & (g2077)) + ((!g1886) & (!g2032) & (g2055) & (g1902) & (g2036) & (g2077)) + ((!g1886) & (g2032) & (!g2055) & (!g1902) & (g2036) & (g2077)) + ((!g1886) & (g2032) & (!g2055) & (g1902) & (g2036) & (g2077)) + ((!g1886) & (g2032) & (g2055) & (!g1902) & (!g2036) & (g2077)) + ((!g1886) & (g2032) & (g2055) & (!g1902) & (g2036) & (!g2077)) + ((!g1886) & (g2032) & (g2055) & (!g1902) & (g2036) & (g2077)) + ((!g1886) & (g2032) & (g2055) & (g1902) & (!g2036) & (g2077)) + ((!g1886) & (g2032) & (g2055) & (g1902) & (g2036) & (!g2077)) + ((!g1886) & (g2032) & (g2055) & (g1902) & (g2036) & (g2077)) + ((g1886) & (!g2032) & (!g2055) & (g1902) & (g2036) & (g2077)) + ((g1886) & (!g2032) & (g2055) & (!g1902) & (!g2036) & (g2077)) + ((g1886) & (!g2032) & (g2055) & (!g1902) & (g2036) & (g2077)) + ((g1886) & (!g2032) & (g2055) & (g1902) & (!g2036) & (g2077)) + ((g1886) & (!g2032) & (g2055) & (g1902) & (g2036) & (!g2077)) + ((g1886) & (!g2032) & (g2055) & (g1902) & (g2036) & (g2077)) + ((g1886) & (g2032) & (!g2055) & (!g1902) & (g2036) & (g2077)) + ((g1886) & (g2032) & (!g2055) & (g1902) & (!g2036) & (g2077)) + ((g1886) & (g2032) & (!g2055) & (g1902) & (g2036) & (g2077)) + ((g1886) & (g2032) & (g2055) & (!g1902) & (!g2036) & (g2077)) + ((g1886) & (g2032) & (g2055) & (!g1902) & (g2036) & (!g2077)) + ((g1886) & (g2032) & (g2055) & (!g1902) & (g2036) & (g2077)) + ((g1886) & (g2032) & (g2055) & (g1902) & (!g2036) & (!g2077)) + ((g1886) & (g2032) & (g2055) & (g1902) & (!g2036) & (g2077)) + ((g1886) & (g2032) & (g2055) & (g1902) & (g2036) & (!g2077)) + ((g1886) & (g2032) & (g2055) & (g1902) & (g2036) & (g2077)));
	assign g3556 = (((!g2194) & (g2198)) + ((g2194) & (!g2198)));
	assign g3557 = (((!g2114) & (!g2137) & (g3555) & (g2118) & (g2159) & (g3556)) + ((!g2114) & (g2137) & (!g3555) & (!g2118) & (g2159) & (g3556)) + ((!g2114) & (g2137) & (!g3555) & (g2118) & (g2159) & (g3556)) + ((!g2114) & (g2137) & (g3555) & (!g2118) & (g2159) & (g3556)) + ((!g2114) & (g2137) & (g3555) & (g2118) & (!g2159) & (g3556)) + ((!g2114) & (g2137) & (g3555) & (g2118) & (g2159) & (g3556)) + ((g2114) & (!g2137) & (!g3555) & (g2118) & (g2159) & (g3556)) + ((g2114) & (!g2137) & (g3555) & (!g2118) & (g2159) & (g3556)) + ((g2114) & (!g2137) & (g3555) & (g2118) & (g2159) & (g3556)) + ((g2114) & (g2137) & (!g3555) & (!g2118) & (g2159) & (g3556)) + ((g2114) & (g2137) & (!g3555) & (g2118) & (!g2159) & (g3556)) + ((g2114) & (g2137) & (!g3555) & (g2118) & (g2159) & (g3556)) + ((g2114) & (g2137) & (g3555) & (!g2118) & (!g2159) & (g3556)) + ((g2114) & (g2137) & (g3555) & (!g2118) & (g2159) & (g3556)) + ((g2114) & (g2137) & (g3555) & (g2118) & (!g2159) & (g3556)) + ((g2114) & (g2137) & (g3555) & (g2118) & (g2159) & (g3556)));
	assign g3558 = (((g2194) & (g2198)));
	assign g3559 = (((!g2217) & (!g2277) & (!g3557) & (!g3558) & (!g2239) & (!g2281)) + ((!g2217) & (!g2277) & (!g3557) & (!g3558) & (!g2239) & (g2281)) + ((!g2217) & (!g2277) & (!g3557) & (!g3558) & (g2239) & (!g2281)) + ((!g2217) & (!g2277) & (!g3557) & (!g3558) & (g2239) & (g2281)) + ((!g2217) & (!g2277) & (!g3557) & (g3558) & (!g2239) & (!g2281)) + ((!g2217) & (!g2277) & (!g3557) & (g3558) & (!g2239) & (g2281)) + ((!g2217) & (!g2277) & (!g3557) & (g3558) & (g2239) & (!g2281)) + ((!g2217) & (!g2277) & (g3557) & (!g3558) & (!g2239) & (!g2281)) + ((!g2217) & (!g2277) & (g3557) & (!g3558) & (!g2239) & (g2281)) + ((!g2217) & (!g2277) & (g3557) & (!g3558) & (g2239) & (!g2281)) + ((!g2217) & (!g2277) & (g3557) & (g3558) & (!g2239) & (!g2281)) + ((!g2217) & (!g2277) & (g3557) & (g3558) & (!g2239) & (g2281)) + ((!g2217) & (!g2277) & (g3557) & (g3558) & (g2239) & (!g2281)) + ((!g2217) & (g2277) & (!g3557) & (!g3558) & (!g2239) & (!g2281)) + ((!g2217) & (g2277) & (!g3557) & (!g3558) & (g2239) & (!g2281)) + ((!g2217) & (g2277) & (!g3557) & (g3558) & (!g2239) & (!g2281)) + ((!g2217) & (g2277) & (g3557) & (!g3558) & (!g2239) & (!g2281)) + ((!g2217) & (g2277) & (g3557) & (g3558) & (!g2239) & (!g2281)) + ((g2217) & (!g2277) & (!g3557) & (!g3558) & (!g2239) & (!g2281)) + ((g2217) & (!g2277) & (!g3557) & (!g3558) & (!g2239) & (g2281)) + ((g2217) & (!g2277) & (!g3557) & (!g3558) & (g2239) & (!g2281)) + ((g2217) & (!g2277) & (!g3557) & (g3558) & (!g2239) & (!g2281)) + ((g2217) & (!g2277) & (!g3557) & (g3558) & (g2239) & (!g2281)) + ((g2217) & (!g2277) & (g3557) & (!g3558) & (!g2239) & (!g2281)) + ((g2217) & (!g2277) & (g3557) & (!g3558) & (g2239) & (!g2281)) + ((g2217) & (!g2277) & (g3557) & (g3558) & (!g2239) & (!g2281)) + ((g2217) & (!g2277) & (g3557) & (g3558) & (g2239) & (!g2281)) + ((g2217) & (g2277) & (!g3557) & (!g3558) & (!g2239) & (!g2281)));
	assign g3560 = (((!g2217) & (!g3557) & (!g3558) & (!g2239) & (!g5788) & (g5789)) + ((!g2217) & (!g3557) & (!g3558) & (g2239) & (!g5788) & (g5789)) + ((!g2217) & (!g3557) & (g3558) & (!g2239) & (!g5788) & (g5789)) + ((!g2217) & (!g3557) & (g3558) & (g2239) & (!g5788) & (g5789)) + ((!g2217) & (!g3557) & (g3558) & (g2239) & (g5788) & (g5789)) + ((!g2217) & (g3557) & (!g3558) & (!g2239) & (!g5788) & (g5789)) + ((!g2217) & (g3557) & (!g3558) & (g2239) & (!g5788) & (g5789)) + ((!g2217) & (g3557) & (!g3558) & (g2239) & (g5788) & (g5789)) + ((!g2217) & (g3557) & (g3558) & (!g2239) & (!g5788) & (g5789)) + ((!g2217) & (g3557) & (g3558) & (g2239) & (!g5788) & (g5789)) + ((!g2217) & (g3557) & (g3558) & (g2239) & (g5788) & (g5789)) + ((g2217) & (!g3557) & (!g3558) & (!g2239) & (!g5788) & (g5789)) + ((g2217) & (!g3557) & (!g3558) & (g2239) & (!g5788) & (g5789)) + ((g2217) & (!g3557) & (!g3558) & (g2239) & (g5788) & (g5789)) + ((g2217) & (!g3557) & (g3558) & (!g2239) & (!g5788) & (g5789)) + ((g2217) & (!g3557) & (g3558) & (!g2239) & (g5788) & (g5789)) + ((g2217) & (!g3557) & (g3558) & (g2239) & (!g5788) & (g5789)) + ((g2217) & (!g3557) & (g3558) & (g2239) & (g5788) & (g5789)) + ((g2217) & (g3557) & (!g3558) & (!g2239) & (!g5788) & (g5789)) + ((g2217) & (g3557) & (!g3558) & (!g2239) & (g5788) & (g5789)) + ((g2217) & (g3557) & (!g3558) & (g2239) & (!g5788) & (g5789)) + ((g2217) & (g3557) & (!g3558) & (g2239) & (g5788) & (g5789)) + ((g2217) & (g3557) & (g3558) & (!g2239) & (!g5788) & (g5789)) + ((g2217) & (g3557) & (g3558) & (!g2239) & (g5788) & (g5789)) + ((g2217) & (g3557) & (g3558) & (g2239) & (!g5788) & (g5789)) + ((g2217) & (g3557) & (g3558) & (g2239) & (g5788) & (g5789)));
	assign g3561 = (((g2383) & (g2405)));
	assign g3562 = (((!g2468) & (!g2523) & (!g3560) & (!g3561) & (!g2480) & (!g2537)) + ((!g2468) & (!g2523) & (!g3560) & (!g3561) & (!g2480) & (g2537)) + ((!g2468) & (!g2523) & (!g3560) & (!g3561) & (g2480) & (!g2537)) + ((!g2468) & (!g2523) & (!g3560) & (!g3561) & (g2480) & (g2537)) + ((!g2468) & (!g2523) & (!g3560) & (g3561) & (!g2480) & (!g2537)) + ((!g2468) & (!g2523) & (!g3560) & (g3561) & (!g2480) & (g2537)) + ((!g2468) & (!g2523) & (!g3560) & (g3561) & (g2480) & (!g2537)) + ((!g2468) & (!g2523) & (g3560) & (!g3561) & (!g2480) & (!g2537)) + ((!g2468) & (!g2523) & (g3560) & (!g3561) & (!g2480) & (g2537)) + ((!g2468) & (!g2523) & (g3560) & (!g3561) & (g2480) & (!g2537)) + ((!g2468) & (!g2523) & (g3560) & (g3561) & (!g2480) & (!g2537)) + ((!g2468) & (!g2523) & (g3560) & (g3561) & (!g2480) & (g2537)) + ((!g2468) & (!g2523) & (g3560) & (g3561) & (g2480) & (!g2537)) + ((!g2468) & (g2523) & (!g3560) & (!g3561) & (!g2480) & (!g2537)) + ((!g2468) & (g2523) & (!g3560) & (!g3561) & (g2480) & (!g2537)) + ((!g2468) & (g2523) & (!g3560) & (g3561) & (!g2480) & (!g2537)) + ((!g2468) & (g2523) & (g3560) & (!g3561) & (!g2480) & (!g2537)) + ((!g2468) & (g2523) & (g3560) & (g3561) & (!g2480) & (!g2537)) + ((g2468) & (!g2523) & (!g3560) & (!g3561) & (!g2480) & (!g2537)) + ((g2468) & (!g2523) & (!g3560) & (!g3561) & (!g2480) & (g2537)) + ((g2468) & (!g2523) & (!g3560) & (!g3561) & (g2480) & (!g2537)) + ((g2468) & (!g2523) & (!g3560) & (g3561) & (!g2480) & (!g2537)) + ((g2468) & (!g2523) & (!g3560) & (g3561) & (g2480) & (!g2537)) + ((g2468) & (!g2523) & (g3560) & (!g3561) & (!g2480) & (!g2537)) + ((g2468) & (!g2523) & (g3560) & (!g3561) & (g2480) & (!g2537)) + ((g2468) & (!g2523) & (g3560) & (g3561) & (!g2480) & (!g2537)) + ((g2468) & (!g2523) & (g3560) & (g3561) & (g2480) & (!g2537)) + ((g2468) & (g2523) & (!g3560) & (!g3561) & (!g2480) & (!g2537)));
	assign g3563 = (((!g2663) & (g2667)) + ((g2663) & (!g2667)));
	assign g3564 = (((!g2575) & (!g2607) & (!g3562) & (g2581) & (g2629) & (g3563)) + ((!g2575) & (g2607) & (!g3562) & (!g2581) & (g2629) & (g3563)) + ((!g2575) & (g2607) & (!g3562) & (g2581) & (!g2629) & (g3563)) + ((!g2575) & (g2607) & (!g3562) & (g2581) & (g2629) & (g3563)) + ((!g2575) & (g2607) & (g3562) & (!g2581) & (g2629) & (g3563)) + ((!g2575) & (g2607) & (g3562) & (g2581) & (g2629) & (g3563)) + ((g2575) & (!g2607) & (!g3562) & (!g2581) & (g2629) & (g3563)) + ((g2575) & (!g2607) & (!g3562) & (g2581) & (g2629) & (g3563)) + ((g2575) & (!g2607) & (g3562) & (g2581) & (g2629) & (g3563)) + ((g2575) & (g2607) & (!g3562) & (!g2581) & (!g2629) & (g3563)) + ((g2575) & (g2607) & (!g3562) & (!g2581) & (g2629) & (g3563)) + ((g2575) & (g2607) & (!g3562) & (g2581) & (!g2629) & (g3563)) + ((g2575) & (g2607) & (!g3562) & (g2581) & (g2629) & (g3563)) + ((g2575) & (g2607) & (g3562) & (!g2581) & (g2629) & (g3563)) + ((g2575) & (g2607) & (g3562) & (g2581) & (!g2629) & (g3563)) + ((g2575) & (g2607) & (g3562) & (g2581) & (g2629) & (g3563)));
	assign g3565 = (((g2663) & (g2667)));
	assign g3566 = (((!g2690) & (!g2774) & (!g3564) & (!g3565) & (!g2728) & (!g2778)) + ((!g2690) & (!g2774) & (!g3564) & (!g3565) & (!g2728) & (g2778)) + ((!g2690) & (!g2774) & (!g3564) & (!g3565) & (g2728) & (!g2778)) + ((!g2690) & (!g2774) & (!g3564) & (!g3565) & (g2728) & (g2778)) + ((!g2690) & (!g2774) & (!g3564) & (g3565) & (!g2728) & (!g2778)) + ((!g2690) & (!g2774) & (!g3564) & (g3565) & (!g2728) & (g2778)) + ((!g2690) & (!g2774) & (!g3564) & (g3565) & (g2728) & (!g2778)) + ((!g2690) & (!g2774) & (g3564) & (!g3565) & (!g2728) & (!g2778)) + ((!g2690) & (!g2774) & (g3564) & (!g3565) & (!g2728) & (g2778)) + ((!g2690) & (!g2774) & (g3564) & (!g3565) & (g2728) & (!g2778)) + ((!g2690) & (!g2774) & (g3564) & (g3565) & (!g2728) & (!g2778)) + ((!g2690) & (!g2774) & (g3564) & (g3565) & (!g2728) & (g2778)) + ((!g2690) & (!g2774) & (g3564) & (g3565) & (g2728) & (!g2778)) + ((!g2690) & (g2774) & (!g3564) & (!g3565) & (!g2728) & (!g2778)) + ((!g2690) & (g2774) & (!g3564) & (!g3565) & (g2728) & (!g2778)) + ((!g2690) & (g2774) & (!g3564) & (g3565) & (!g2728) & (!g2778)) + ((!g2690) & (g2774) & (g3564) & (!g3565) & (!g2728) & (!g2778)) + ((!g2690) & (g2774) & (g3564) & (g3565) & (!g2728) & (!g2778)) + ((g2690) & (!g2774) & (!g3564) & (!g3565) & (!g2728) & (!g2778)) + ((g2690) & (!g2774) & (!g3564) & (!g3565) & (!g2728) & (g2778)) + ((g2690) & (!g2774) & (!g3564) & (!g3565) & (g2728) & (!g2778)) + ((g2690) & (!g2774) & (!g3564) & (g3565) & (!g2728) & (!g2778)) + ((g2690) & (!g2774) & (!g3564) & (g3565) & (g2728) & (!g2778)) + ((g2690) & (!g2774) & (g3564) & (!g3565) & (!g2728) & (!g2778)) + ((g2690) & (!g2774) & (g3564) & (!g3565) & (g2728) & (!g2778)) + ((g2690) & (!g2774) & (g3564) & (g3565) & (!g2728) & (!g2778)) + ((g2690) & (!g2774) & (g3564) & (g3565) & (g2728) & (!g2778)) + ((g2690) & (g2774) & (!g3564) & (!g3565) & (!g2728) & (!g2778)));
	assign g3567 = (((!g2881) & (g2895)) + ((g2881) & (!g2895)));
	assign g3568 = (((!g2797) & (!g2854) & (!g3566) & (g2819) & (g2860) & (g3567)) + ((!g2797) & (g2854) & (!g3566) & (!g2819) & (g2860) & (g3567)) + ((!g2797) & (g2854) & (!g3566) & (g2819) & (!g2860) & (g3567)) + ((!g2797) & (g2854) & (!g3566) & (g2819) & (g2860) & (g3567)) + ((!g2797) & (g2854) & (g3566) & (!g2819) & (g2860) & (g3567)) + ((!g2797) & (g2854) & (g3566) & (g2819) & (g2860) & (g3567)) + ((g2797) & (!g2854) & (!g3566) & (!g2819) & (g2860) & (g3567)) + ((g2797) & (!g2854) & (!g3566) & (g2819) & (g2860) & (g3567)) + ((g2797) & (!g2854) & (g3566) & (g2819) & (g2860) & (g3567)) + ((g2797) & (g2854) & (!g3566) & (!g2819) & (!g2860) & (g3567)) + ((g2797) & (g2854) & (!g3566) & (!g2819) & (g2860) & (g3567)) + ((g2797) & (g2854) & (!g3566) & (g2819) & (!g2860) & (g3567)) + ((g2797) & (g2854) & (!g3566) & (g2819) & (g2860) & (g3567)) + ((g2797) & (g2854) & (g3566) & (!g2819) & (g2860) & (g3567)) + ((g2797) & (g2854) & (g3566) & (g2819) & (!g2860) & (g3567)) + ((g2797) & (g2854) & (g3566) & (g2819) & (g2860) & (g3567)));
	assign g3569 = (((g2881) & (g2895)));
	assign g3570 = (((!g2950) & (!g2999) & (!g3568) & (!g3569) & (!g2962) & (!g3013)) + ((!g2950) & (!g2999) & (!g3568) & (!g3569) & (!g2962) & (g3013)) + ((!g2950) & (!g2999) & (!g3568) & (!g3569) & (g2962) & (!g3013)) + ((!g2950) & (!g2999) & (!g3568) & (!g3569) & (g2962) & (g3013)) + ((!g2950) & (!g2999) & (!g3568) & (g3569) & (!g2962) & (!g3013)) + ((!g2950) & (!g2999) & (!g3568) & (g3569) & (!g2962) & (g3013)) + ((!g2950) & (!g2999) & (!g3568) & (g3569) & (g2962) & (!g3013)) + ((!g2950) & (!g2999) & (g3568) & (!g3569) & (!g2962) & (!g3013)) + ((!g2950) & (!g2999) & (g3568) & (!g3569) & (!g2962) & (g3013)) + ((!g2950) & (!g2999) & (g3568) & (!g3569) & (g2962) & (!g3013)) + ((!g2950) & (!g2999) & (g3568) & (g3569) & (!g2962) & (!g3013)) + ((!g2950) & (!g2999) & (g3568) & (g3569) & (!g2962) & (g3013)) + ((!g2950) & (!g2999) & (g3568) & (g3569) & (g2962) & (!g3013)) + ((!g2950) & (g2999) & (!g3568) & (!g3569) & (!g2962) & (!g3013)) + ((!g2950) & (g2999) & (!g3568) & (!g3569) & (g2962) & (!g3013)) + ((!g2950) & (g2999) & (!g3568) & (g3569) & (!g2962) & (!g3013)) + ((!g2950) & (g2999) & (g3568) & (!g3569) & (!g2962) & (!g3013)) + ((!g2950) & (g2999) & (g3568) & (g3569) & (!g2962) & (!g3013)) + ((g2950) & (!g2999) & (!g3568) & (!g3569) & (!g2962) & (!g3013)) + ((g2950) & (!g2999) & (!g3568) & (!g3569) & (!g2962) & (g3013)) + ((g2950) & (!g2999) & (!g3568) & (!g3569) & (g2962) & (!g3013)) + ((g2950) & (!g2999) & (!g3568) & (g3569) & (!g2962) & (!g3013)) + ((g2950) & (!g2999) & (!g3568) & (g3569) & (g2962) & (!g3013)) + ((g2950) & (!g2999) & (g3568) & (!g3569) & (!g2962) & (!g3013)) + ((g2950) & (!g2999) & (g3568) & (!g3569) & (g2962) & (!g3013)) + ((g2950) & (!g2999) & (g3568) & (g3569) & (!g2962) & (!g3013)) + ((g2950) & (!g2999) & (g3568) & (g3569) & (g2962) & (!g3013)) + ((g2950) & (g2999) & (!g3568) & (!g3569) & (!g2962) & (!g3013)));
	assign g3571 = (((!g3047) & (!g3570) & (g3053)) + ((g3047) & (!g3570) & (!g3053)) + ((g3047) & (!g3570) & (g3053)) + ((g3047) & (g3570) & (g3053)));
	assign g3572 = (((!g1890) & (!g1939) & (g1941) & (!g1896) & (!g2041) & (g2068)) + ((!g1890) & (!g1939) & (g1941) & (!g1896) & (g2041) & (g2068)) + ((!g1890) & (!g1939) & (g1941) & (g1896) & (!g2041) & (g2068)) + ((!g1890) & (!g1939) & (g1941) & (g1896) & (g2041) & (g2068)) + ((!g1890) & (g1939) & (!g1941) & (!g1896) & (g2041) & (g2068)) + ((!g1890) & (g1939) & (!g1941) & (g1896) & (g2041) & (g2068)) + ((!g1890) & (g1939) & (g1941) & (!g1896) & (!g2041) & (g2068)) + ((!g1890) & (g1939) & (g1941) & (!g1896) & (g2041) & (!g2068)) + ((!g1890) & (g1939) & (g1941) & (!g1896) & (g2041) & (g2068)) + ((!g1890) & (g1939) & (g1941) & (g1896) & (!g2041) & (g2068)) + ((!g1890) & (g1939) & (g1941) & (g1896) & (g2041) & (!g2068)) + ((!g1890) & (g1939) & (g1941) & (g1896) & (g2041) & (g2068)) + ((g1890) & (!g1939) & (!g1941) & (g1896) & (g2041) & (g2068)) + ((g1890) & (!g1939) & (g1941) & (!g1896) & (!g2041) & (g2068)) + ((g1890) & (!g1939) & (g1941) & (!g1896) & (g2041) & (g2068)) + ((g1890) & (!g1939) & (g1941) & (g1896) & (!g2041) & (g2068)) + ((g1890) & (!g1939) & (g1941) & (g1896) & (g2041) & (!g2068)) + ((g1890) & (!g1939) & (g1941) & (g1896) & (g2041) & (g2068)) + ((g1890) & (g1939) & (!g1941) & (!g1896) & (g2041) & (g2068)) + ((g1890) & (g1939) & (!g1941) & (g1896) & (!g2041) & (g2068)) + ((g1890) & (g1939) & (!g1941) & (g1896) & (g2041) & (g2068)) + ((g1890) & (g1939) & (g1941) & (!g1896) & (!g2041) & (g2068)) + ((g1890) & (g1939) & (g1941) & (!g1896) & (g2041) & (!g2068)) + ((g1890) & (g1939) & (g1941) & (!g1896) & (g2041) & (g2068)) + ((g1890) & (g1939) & (g1941) & (g1896) & (!g2041) & (!g2068)) + ((g1890) & (g1939) & (g1941) & (g1896) & (!g2041) & (g2068)) + ((g1890) & (g1939) & (g1941) & (g1896) & (g2041) & (!g2068)) + ((g1890) & (g1939) & (g1941) & (g1896) & (g2041) & (g2068)));
	assign g3573 = (((!g1948) & (g2203)) + ((g1948) & (!g2203)));
	assign g3574 = (((!g1944) & (!g1946) & (g2123) & (g2150) & (g3572) & (g3573)) + ((!g1944) & (g1946) & (!g2123) & (g2150) & (!g3572) & (g3573)) + ((!g1944) & (g1946) & (!g2123) & (g2150) & (g3572) & (g3573)) + ((!g1944) & (g1946) & (g2123) & (!g2150) & (g3572) & (g3573)) + ((!g1944) & (g1946) & (g2123) & (g2150) & (!g3572) & (g3573)) + ((!g1944) & (g1946) & (g2123) & (g2150) & (g3572) & (g3573)) + ((g1944) & (!g1946) & (!g2123) & (g2150) & (g3572) & (g3573)) + ((g1944) & (!g1946) & (g2123) & (g2150) & (!g3572) & (g3573)) + ((g1944) & (!g1946) & (g2123) & (g2150) & (g3572) & (g3573)) + ((g1944) & (g1946) & (!g2123) & (!g2150) & (g3572) & (g3573)) + ((g1944) & (g1946) & (!g2123) & (g2150) & (!g3572) & (g3573)) + ((g1944) & (g1946) & (!g2123) & (g2150) & (g3572) & (g3573)) + ((g1944) & (g1946) & (g2123) & (!g2150) & (!g3572) & (g3573)) + ((g1944) & (g1946) & (g2123) & (!g2150) & (g3572) & (g3573)) + ((g1944) & (g1946) & (g2123) & (g2150) & (!g3572) & (g3573)) + ((g1944) & (g1946) & (g2123) & (g2150) & (g3572) & (g3573)));
	assign g3575 = (((g1948) & (g2203)));
	assign g3576 = (((!g1953) & (!g1955) & (!g2230) & (!g2286) & (!g3574) & (!g3575)) + ((!g1953) & (!g1955) & (!g2230) & (!g2286) & (!g3574) & (g3575)) + ((!g1953) & (!g1955) & (!g2230) & (!g2286) & (g3574) & (!g3575)) + ((!g1953) & (!g1955) & (!g2230) & (!g2286) & (g3574) & (g3575)) + ((!g1953) & (!g1955) & (!g2230) & (g2286) & (!g3574) & (!g3575)) + ((!g1953) & (!g1955) & (!g2230) & (g2286) & (!g3574) & (g3575)) + ((!g1953) & (!g1955) & (!g2230) & (g2286) & (g3574) & (!g3575)) + ((!g1953) & (!g1955) & (!g2230) & (g2286) & (g3574) & (g3575)) + ((!g1953) & (!g1955) & (g2230) & (!g2286) & (!g3574) & (!g3575)) + ((!g1953) & (!g1955) & (g2230) & (!g2286) & (!g3574) & (g3575)) + ((!g1953) & (!g1955) & (g2230) & (!g2286) & (g3574) & (!g3575)) + ((!g1953) & (!g1955) & (g2230) & (!g2286) & (g3574) & (g3575)) + ((!g1953) & (!g1955) & (g2230) & (g2286) & (!g3574) & (!g3575)) + ((!g1953) & (g1955) & (!g2230) & (!g2286) & (!g3574) & (!g3575)) + ((!g1953) & (g1955) & (!g2230) & (!g2286) & (!g3574) & (g3575)) + ((!g1953) & (g1955) & (!g2230) & (!g2286) & (g3574) & (!g3575)) + ((!g1953) & (g1955) & (!g2230) & (!g2286) & (g3574) & (g3575)) + ((!g1953) & (g1955) & (g2230) & (!g2286) & (!g3574) & (!g3575)) + ((g1953) & (!g1955) & (!g2230) & (!g2286) & (!g3574) & (!g3575)) + ((g1953) & (!g1955) & (!g2230) & (!g2286) & (!g3574) & (g3575)) + ((g1953) & (!g1955) & (!g2230) & (!g2286) & (g3574) & (!g3575)) + ((g1953) & (!g1955) & (!g2230) & (!g2286) & (g3574) & (g3575)) + ((g1953) & (!g1955) & (!g2230) & (g2286) & (!g3574) & (!g3575)) + ((g1953) & (!g1955) & (g2230) & (!g2286) & (!g3574) & (!g3575)) + ((g1953) & (!g1955) & (g2230) & (!g2286) & (!g3574) & (g3575)) + ((g1953) & (!g1955) & (g2230) & (!g2286) & (g3574) & (!g3575)) + ((g1953) & (!g1955) & (g2230) & (!g2286) & (g3574) & (g3575)) + ((g1953) & (g1955) & (!g2230) & (!g2286) & (!g3574) & (!g3575)));
	assign g3577 = (((!g1962) & (g2396)) + ((g1962) & (!g2396)));
	assign g3578 = (((!g1958) & (!g1960) & (g2317) & (g2369) & (!g3576) & (g3577)) + ((!g1958) & (g1960) & (!g2317) & (g2369) & (!g3576) & (g3577)) + ((!g1958) & (g1960) & (!g2317) & (g2369) & (g3576) & (g3577)) + ((!g1958) & (g1960) & (g2317) & (!g2369) & (!g3576) & (g3577)) + ((!g1958) & (g1960) & (g2317) & (g2369) & (!g3576) & (g3577)) + ((!g1958) & (g1960) & (g2317) & (g2369) & (g3576) & (g3577)) + ((g1958) & (!g1960) & (!g2317) & (g2369) & (!g3576) & (g3577)) + ((g1958) & (!g1960) & (g2317) & (g2369) & (!g3576) & (g3577)) + ((g1958) & (!g1960) & (g2317) & (g2369) & (g3576) & (g3577)) + ((g1958) & (g1960) & (!g2317) & (!g2369) & (!g3576) & (g3577)) + ((g1958) & (g1960) & (!g2317) & (g2369) & (!g3576) & (g3577)) + ((g1958) & (g1960) & (!g2317) & (g2369) & (g3576) & (g3577)) + ((g1958) & (g1960) & (g2317) & (!g2369) & (!g3576) & (g3577)) + ((g1958) & (g1960) & (g2317) & (!g2369) & (g3576) & (g3577)) + ((g1958) & (g1960) & (g2317) & (g2369) & (!g3576) & (g3577)) + ((g1958) & (g1960) & (g2317) & (g2369) & (g3576) & (g3577)));
	assign g3579 = (((g1962) & (g2396)));
	assign g3580 = (((!g1967) & (!g1969) & (!g2497) & (!g2531) & (!g3578) & (!g3579)) + ((!g1967) & (!g1969) & (!g2497) & (!g2531) & (!g3578) & (g3579)) + ((!g1967) & (!g1969) & (!g2497) & (!g2531) & (g3578) & (!g3579)) + ((!g1967) & (!g1969) & (!g2497) & (!g2531) & (g3578) & (g3579)) + ((!g1967) & (!g1969) & (!g2497) & (g2531) & (!g3578) & (!g3579)) + ((!g1967) & (!g1969) & (!g2497) & (g2531) & (!g3578) & (g3579)) + ((!g1967) & (!g1969) & (!g2497) & (g2531) & (g3578) & (!g3579)) + ((!g1967) & (!g1969) & (!g2497) & (g2531) & (g3578) & (g3579)) + ((!g1967) & (!g1969) & (g2497) & (!g2531) & (!g3578) & (!g3579)) + ((!g1967) & (!g1969) & (g2497) & (!g2531) & (!g3578) & (g3579)) + ((!g1967) & (!g1969) & (g2497) & (!g2531) & (g3578) & (!g3579)) + ((!g1967) & (!g1969) & (g2497) & (!g2531) & (g3578) & (g3579)) + ((!g1967) & (!g1969) & (g2497) & (g2531) & (!g3578) & (!g3579)) + ((!g1967) & (g1969) & (!g2497) & (!g2531) & (!g3578) & (!g3579)) + ((!g1967) & (g1969) & (!g2497) & (!g2531) & (!g3578) & (g3579)) + ((!g1967) & (g1969) & (!g2497) & (!g2531) & (g3578) & (!g3579)) + ((!g1967) & (g1969) & (!g2497) & (!g2531) & (g3578) & (g3579)) + ((!g1967) & (g1969) & (g2497) & (!g2531) & (!g3578) & (!g3579)) + ((g1967) & (!g1969) & (!g2497) & (!g2531) & (!g3578) & (!g3579)) + ((g1967) & (!g1969) & (!g2497) & (!g2531) & (!g3578) & (g3579)) + ((g1967) & (!g1969) & (!g2497) & (!g2531) & (g3578) & (!g3579)) + ((g1967) & (!g1969) & (!g2497) & (!g2531) & (g3578) & (g3579)) + ((g1967) & (!g1969) & (!g2497) & (g2531) & (!g3578) & (!g3579)) + ((g1967) & (!g1969) & (g2497) & (!g2531) & (!g3578) & (!g3579)) + ((g1967) & (!g1969) & (g2497) & (!g2531) & (!g3578) & (g3579)) + ((g1967) & (!g1969) & (g2497) & (!g2531) & (g3578) & (!g3579)) + ((g1967) & (!g1969) & (g2497) & (!g2531) & (g3578) & (g3579)) + ((g1967) & (g1969) & (!g2497) & (!g2531) & (!g3578) & (!g3579)));
	assign g3581 = (((!g2047) & (g2672)) + ((g2047) & (!g2672)));
	assign g3582 = (((!g1972) & (!g1975) & (g2589) & (g2620) & (!g3580) & (g3581)) + ((!g1972) & (g1975) & (!g2589) & (g2620) & (!g3580) & (g3581)) + ((!g1972) & (g1975) & (!g2589) & (g2620) & (g3580) & (g3581)) + ((!g1972) & (g1975) & (g2589) & (!g2620) & (!g3580) & (g3581)) + ((!g1972) & (g1975) & (g2589) & (g2620) & (!g3580) & (g3581)) + ((!g1972) & (g1975) & (g2589) & (g2620) & (g3580) & (g3581)) + ((g1972) & (!g1975) & (!g2589) & (g2620) & (!g3580) & (g3581)) + ((g1972) & (!g1975) & (g2589) & (g2620) & (!g3580) & (g3581)) + ((g1972) & (!g1975) & (g2589) & (g2620) & (g3580) & (g3581)) + ((g1972) & (g1975) & (!g2589) & (!g2620) & (!g3580) & (g3581)) + ((g1972) & (g1975) & (!g2589) & (g2620) & (!g3580) & (g3581)) + ((g1972) & (g1975) & (!g2589) & (g2620) & (g3580) & (g3581)) + ((g1972) & (g1975) & (g2589) & (!g2620) & (!g3580) & (g3581)) + ((g1972) & (g1975) & (g2589) & (!g2620) & (g3580) & (g3581)) + ((g1972) & (g1975) & (g2589) & (g2620) & (!g3580) & (g3581)) + ((g1972) & (g1975) & (g2589) & (g2620) & (g3580) & (g3581)));
	assign g3583 = (((g2047) & (g2672)));
	assign g3584 = (((!g2098) & (!g2129) & (!g2713) & (!g2783) & (!g3582) & (!g3583)) + ((!g2098) & (!g2129) & (!g2713) & (!g2783) & (!g3582) & (g3583)) + ((!g2098) & (!g2129) & (!g2713) & (!g2783) & (g3582) & (!g3583)) + ((!g2098) & (!g2129) & (!g2713) & (!g2783) & (g3582) & (g3583)) + ((!g2098) & (!g2129) & (!g2713) & (g2783) & (!g3582) & (!g3583)) + ((!g2098) & (!g2129) & (!g2713) & (g2783) & (!g3582) & (g3583)) + ((!g2098) & (!g2129) & (!g2713) & (g2783) & (g3582) & (!g3583)) + ((!g2098) & (!g2129) & (!g2713) & (g2783) & (g3582) & (g3583)) + ((!g2098) & (!g2129) & (g2713) & (!g2783) & (!g3582) & (!g3583)) + ((!g2098) & (!g2129) & (g2713) & (!g2783) & (!g3582) & (g3583)) + ((!g2098) & (!g2129) & (g2713) & (!g2783) & (g3582) & (!g3583)) + ((!g2098) & (!g2129) & (g2713) & (!g2783) & (g3582) & (g3583)) + ((!g2098) & (!g2129) & (g2713) & (g2783) & (!g3582) & (!g3583)) + ((!g2098) & (g2129) & (!g2713) & (!g2783) & (!g3582) & (!g3583)) + ((!g2098) & (g2129) & (!g2713) & (!g2783) & (!g3582) & (g3583)) + ((!g2098) & (g2129) & (!g2713) & (!g2783) & (g3582) & (!g3583)) + ((!g2098) & (g2129) & (!g2713) & (!g2783) & (g3582) & (g3583)) + ((!g2098) & (g2129) & (g2713) & (!g2783) & (!g3582) & (!g3583)) + ((g2098) & (!g2129) & (!g2713) & (!g2783) & (!g3582) & (!g3583)) + ((g2098) & (!g2129) & (!g2713) & (!g2783) & (!g3582) & (g3583)) + ((g2098) & (!g2129) & (!g2713) & (!g2783) & (g3582) & (!g3583)) + ((g2098) & (!g2129) & (!g2713) & (!g2783) & (g3582) & (g3583)) + ((g2098) & (!g2129) & (!g2713) & (g2783) & (!g3582) & (!g3583)) + ((g2098) & (!g2129) & (g2713) & (!g2783) & (!g3582) & (!g3583)) + ((g2098) & (!g2129) & (g2713) & (!g2783) & (!g3582) & (g3583)) + ((g2098) & (!g2129) & (g2713) & (!g2783) & (g3582) & (!g3583)) + ((g2098) & (!g2129) & (g2713) & (!g2783) & (g3582) & (g3583)) + ((g2098) & (g2129) & (!g2713) & (!g2783) & (!g3582) & (!g3583)));
	assign g3585 = (((!g2177) & (g2810) & (!g3584)) + ((g2177) & (!g2810) & (!g3584)) + ((g2177) & (g2810) & (!g3584)) + ((g2177) & (g2810) & (g3584)));
	assign g3586 = (((!g2210) & (!g2868) & (g3585)) + ((!g2210) & (g2868) & (!g3585)) + ((g2210) & (!g2868) & (!g3585)) + ((g2210) & (g2868) & (g3585)));
	assign g3587 = (((!g830) & (!g1894) & (!g7042) & (nonce[0])) + ((!g830) & (!g1894) & (g7042) & (nonce[0])) + ((!g830) & (g1894) & (!g7042) & (nonce[0])) + ((!g830) & (g1894) & (g7042) & (nonce[0])) + ((g830) & (!g1894) & (g7042) & (!nonce[0])) + ((g830) & (!g1894) & (g7042) & (nonce[0])) + ((g830) & (g1894) & (!g7042) & (!nonce[0])) + ((g830) & (g1894) & (!g7042) & (nonce[0])));
	assign g3588 = (((!g1888) & (!g1978) & (g1980) & (!g1904) & (!g2043) & (g2080)) + ((!g1888) & (!g1978) & (g1980) & (!g1904) & (g2043) & (g2080)) + ((!g1888) & (!g1978) & (g1980) & (g1904) & (!g2043) & (g2080)) + ((!g1888) & (!g1978) & (g1980) & (g1904) & (g2043) & (g2080)) + ((!g1888) & (g1978) & (!g1980) & (!g1904) & (g2043) & (g2080)) + ((!g1888) & (g1978) & (!g1980) & (g1904) & (g2043) & (g2080)) + ((!g1888) & (g1978) & (g1980) & (!g1904) & (!g2043) & (g2080)) + ((!g1888) & (g1978) & (g1980) & (!g1904) & (g2043) & (!g2080)) + ((!g1888) & (g1978) & (g1980) & (!g1904) & (g2043) & (g2080)) + ((!g1888) & (g1978) & (g1980) & (g1904) & (!g2043) & (g2080)) + ((!g1888) & (g1978) & (g1980) & (g1904) & (g2043) & (!g2080)) + ((!g1888) & (g1978) & (g1980) & (g1904) & (g2043) & (g2080)) + ((g1888) & (!g1978) & (!g1980) & (g1904) & (g2043) & (g2080)) + ((g1888) & (!g1978) & (g1980) & (!g1904) & (!g2043) & (g2080)) + ((g1888) & (!g1978) & (g1980) & (!g1904) & (g2043) & (g2080)) + ((g1888) & (!g1978) & (g1980) & (g1904) & (!g2043) & (g2080)) + ((g1888) & (!g1978) & (g1980) & (g1904) & (g2043) & (!g2080)) + ((g1888) & (!g1978) & (g1980) & (g1904) & (g2043) & (g2080)) + ((g1888) & (g1978) & (!g1980) & (!g1904) & (g2043) & (g2080)) + ((g1888) & (g1978) & (!g1980) & (g1904) & (!g2043) & (g2080)) + ((g1888) & (g1978) & (!g1980) & (g1904) & (g2043) & (g2080)) + ((g1888) & (g1978) & (g1980) & (!g1904) & (!g2043) & (g2080)) + ((g1888) & (g1978) & (g1980) & (!g1904) & (g2043) & (!g2080)) + ((g1888) & (g1978) & (g1980) & (!g1904) & (g2043) & (g2080)) + ((g1888) & (g1978) & (g1980) & (g1904) & (!g2043) & (!g2080)) + ((g1888) & (g1978) & (g1980) & (g1904) & (!g2043) & (g2080)) + ((g1888) & (g1978) & (g1980) & (g1904) & (g2043) & (!g2080)) + ((g1888) & (g1978) & (g1980) & (g1904) & (g2043) & (g2080)));
	assign g3589 = (((!g1987) & (g2205)) + ((g1987) & (!g2205)));
	assign g3590 = (((!g1983) & (!g1985) & (g3588) & (g2125) & (g2162) & (g3589)) + ((!g1983) & (g1985) & (!g3588) & (!g2125) & (g2162) & (g3589)) + ((!g1983) & (g1985) & (!g3588) & (g2125) & (g2162) & (g3589)) + ((!g1983) & (g1985) & (g3588) & (!g2125) & (g2162) & (g3589)) + ((!g1983) & (g1985) & (g3588) & (g2125) & (!g2162) & (g3589)) + ((!g1983) & (g1985) & (g3588) & (g2125) & (g2162) & (g3589)) + ((g1983) & (!g1985) & (!g3588) & (g2125) & (g2162) & (g3589)) + ((g1983) & (!g1985) & (g3588) & (!g2125) & (g2162) & (g3589)) + ((g1983) & (!g1985) & (g3588) & (g2125) & (g2162) & (g3589)) + ((g1983) & (g1985) & (!g3588) & (!g2125) & (g2162) & (g3589)) + ((g1983) & (g1985) & (!g3588) & (g2125) & (!g2162) & (g3589)) + ((g1983) & (g1985) & (!g3588) & (g2125) & (g2162) & (g3589)) + ((g1983) & (g1985) & (g3588) & (!g2125) & (!g2162) & (g3589)) + ((g1983) & (g1985) & (g3588) & (!g2125) & (g2162) & (g3589)) + ((g1983) & (g1985) & (g3588) & (g2125) & (!g2162) & (g3589)) + ((g1983) & (g1985) & (g3588) & (g2125) & (g2162) & (g3589)));
	assign g3591 = (((g1987) & (g2205)));
	assign g3592 = (((!g1992) & (!g1994) & (!g3590) & (!g3591) & (!g2242) & (!g2288)) + ((!g1992) & (!g1994) & (!g3590) & (!g3591) & (!g2242) & (g2288)) + ((!g1992) & (!g1994) & (!g3590) & (!g3591) & (g2242) & (!g2288)) + ((!g1992) & (!g1994) & (!g3590) & (!g3591) & (g2242) & (g2288)) + ((!g1992) & (!g1994) & (!g3590) & (g3591) & (!g2242) & (!g2288)) + ((!g1992) & (!g1994) & (!g3590) & (g3591) & (!g2242) & (g2288)) + ((!g1992) & (!g1994) & (!g3590) & (g3591) & (g2242) & (!g2288)) + ((!g1992) & (!g1994) & (g3590) & (!g3591) & (!g2242) & (!g2288)) + ((!g1992) & (!g1994) & (g3590) & (!g3591) & (!g2242) & (g2288)) + ((!g1992) & (!g1994) & (g3590) & (!g3591) & (g2242) & (!g2288)) + ((!g1992) & (!g1994) & (g3590) & (g3591) & (!g2242) & (!g2288)) + ((!g1992) & (!g1994) & (g3590) & (g3591) & (!g2242) & (g2288)) + ((!g1992) & (!g1994) & (g3590) & (g3591) & (g2242) & (!g2288)) + ((!g1992) & (g1994) & (!g3590) & (!g3591) & (!g2242) & (!g2288)) + ((!g1992) & (g1994) & (!g3590) & (!g3591) & (g2242) & (!g2288)) + ((!g1992) & (g1994) & (!g3590) & (g3591) & (!g2242) & (!g2288)) + ((!g1992) & (g1994) & (g3590) & (!g3591) & (!g2242) & (!g2288)) + ((!g1992) & (g1994) & (g3590) & (g3591) & (!g2242) & (!g2288)) + ((g1992) & (!g1994) & (!g3590) & (!g3591) & (!g2242) & (!g2288)) + ((g1992) & (!g1994) & (!g3590) & (!g3591) & (!g2242) & (g2288)) + ((g1992) & (!g1994) & (!g3590) & (!g3591) & (g2242) & (!g2288)) + ((g1992) & (!g1994) & (!g3590) & (g3591) & (!g2242) & (!g2288)) + ((g1992) & (!g1994) & (!g3590) & (g3591) & (g2242) & (!g2288)) + ((g1992) & (!g1994) & (g3590) & (!g3591) & (!g2242) & (!g2288)) + ((g1992) & (!g1994) & (g3590) & (!g3591) & (g2242) & (!g2288)) + ((g1992) & (!g1994) & (g3590) & (g3591) & (!g2242) & (!g2288)) + ((g1992) & (!g1994) & (g3590) & (g3591) & (g2242) & (!g2288)) + ((g1992) & (g1994) & (!g3590) & (!g3591) & (!g2242) & (!g2288)));
	assign g3593 = (((!g2002) & (g2408)) + ((g2002) & (!g2408)));
	assign g3594 = (((!g1997) & (!g1999) & (!g3592) & (g2329) & (g2371) & (g3593)) + ((!g1997) & (g1999) & (!g3592) & (!g2329) & (g2371) & (g3593)) + ((!g1997) & (g1999) & (!g3592) & (g2329) & (!g2371) & (g3593)) + ((!g1997) & (g1999) & (!g3592) & (g2329) & (g2371) & (g3593)) + ((!g1997) & (g1999) & (g3592) & (!g2329) & (g2371) & (g3593)) + ((!g1997) & (g1999) & (g3592) & (g2329) & (g2371) & (g3593)) + ((g1997) & (!g1999) & (!g3592) & (!g2329) & (g2371) & (g3593)) + ((g1997) & (!g1999) & (!g3592) & (g2329) & (g2371) & (g3593)) + ((g1997) & (!g1999) & (g3592) & (g2329) & (g2371) & (g3593)) + ((g1997) & (g1999) & (!g3592) & (!g2329) & (!g2371) & (g3593)) + ((g1997) & (g1999) & (!g3592) & (!g2329) & (g2371) & (g3593)) + ((g1997) & (g1999) & (!g3592) & (g2329) & (!g2371) & (g3593)) + ((g1997) & (g1999) & (!g3592) & (g2329) & (g2371) & (g3593)) + ((g1997) & (g1999) & (g3592) & (!g2329) & (g2371) & (g3593)) + ((g1997) & (g1999) & (g3592) & (g2329) & (!g2371) & (g3593)) + ((g1997) & (g1999) & (g3592) & (g2329) & (g2371) & (g3593)));
	assign g3595 = (((g2002) & (g2408)));
	assign g3596 = (((!g2004) & (!g2006) & (!g3594) & (!g3595) & (!g2503) & (!g2539)) + ((!g2004) & (!g2006) & (!g3594) & (!g3595) & (!g2503) & (g2539)) + ((!g2004) & (!g2006) & (!g3594) & (!g3595) & (g2503) & (!g2539)) + ((!g2004) & (!g2006) & (!g3594) & (!g3595) & (g2503) & (g2539)) + ((!g2004) & (!g2006) & (!g3594) & (g3595) & (!g2503) & (!g2539)) + ((!g2004) & (!g2006) & (!g3594) & (g3595) & (!g2503) & (g2539)) + ((!g2004) & (!g2006) & (!g3594) & (g3595) & (g2503) & (!g2539)) + ((!g2004) & (!g2006) & (g3594) & (!g3595) & (!g2503) & (!g2539)) + ((!g2004) & (!g2006) & (g3594) & (!g3595) & (!g2503) & (g2539)) + ((!g2004) & (!g2006) & (g3594) & (!g3595) & (g2503) & (!g2539)) + ((!g2004) & (!g2006) & (g3594) & (g3595) & (!g2503) & (!g2539)) + ((!g2004) & (!g2006) & (g3594) & (g3595) & (!g2503) & (g2539)) + ((!g2004) & (!g2006) & (g3594) & (g3595) & (g2503) & (!g2539)) + ((!g2004) & (g2006) & (!g3594) & (!g3595) & (!g2503) & (!g2539)) + ((!g2004) & (g2006) & (!g3594) & (!g3595) & (g2503) & (!g2539)) + ((!g2004) & (g2006) & (!g3594) & (g3595) & (!g2503) & (!g2539)) + ((!g2004) & (g2006) & (g3594) & (!g3595) & (!g2503) & (!g2539)) + ((!g2004) & (g2006) & (g3594) & (g3595) & (!g2503) & (!g2539)) + ((g2004) & (!g2006) & (!g3594) & (!g3595) & (!g2503) & (!g2539)) + ((g2004) & (!g2006) & (!g3594) & (!g3595) & (!g2503) & (g2539)) + ((g2004) & (!g2006) & (!g3594) & (!g3595) & (g2503) & (!g2539)) + ((g2004) & (!g2006) & (!g3594) & (g3595) & (!g2503) & (!g2539)) + ((g2004) & (!g2006) & (!g3594) & (g3595) & (g2503) & (!g2539)) + ((g2004) & (!g2006) & (g3594) & (!g3595) & (!g2503) & (!g2539)) + ((g2004) & (!g2006) & (g3594) & (!g3595) & (g2503) & (!g2539)) + ((g2004) & (!g2006) & (g3594) & (g3595) & (!g2503) & (!g2539)) + ((g2004) & (!g2006) & (g3594) & (g3595) & (g2503) & (!g2539)) + ((g2004) & (g2006) & (!g3594) & (!g3595) & (!g2503) & (!g2539)));
	assign g3597 = (((!g2052) & (g2674)) + ((g2052) & (!g2674)));
	assign g3598 = (((!g2012) & (!g2014) & (!g3596) & (g2592) & (g2632) & (g3597)) + ((!g2012) & (g2014) & (!g3596) & (!g2592) & (g2632) & (g3597)) + ((!g2012) & (g2014) & (!g3596) & (g2592) & (!g2632) & (g3597)) + ((!g2012) & (g2014) & (!g3596) & (g2592) & (g2632) & (g3597)) + ((!g2012) & (g2014) & (g3596) & (!g2592) & (g2632) & (g3597)) + ((!g2012) & (g2014) & (g3596) & (g2592) & (g2632) & (g3597)) + ((g2012) & (!g2014) & (!g3596) & (!g2592) & (g2632) & (g3597)) + ((g2012) & (!g2014) & (!g3596) & (g2592) & (g2632) & (g3597)) + ((g2012) & (!g2014) & (g3596) & (g2592) & (g2632) & (g3597)) + ((g2012) & (g2014) & (!g3596) & (!g2592) & (!g2632) & (g3597)) + ((g2012) & (g2014) & (!g3596) & (!g2592) & (g2632) & (g3597)) + ((g2012) & (g2014) & (!g3596) & (g2592) & (!g2632) & (g3597)) + ((g2012) & (g2014) & (!g3596) & (g2592) & (g2632) & (g3597)) + ((g2012) & (g2014) & (g3596) & (!g2592) & (g2632) & (g3597)) + ((g2012) & (g2014) & (g3596) & (g2592) & (!g2632) & (g3597)) + ((g2012) & (g2014) & (g3596) & (g2592) & (g2632) & (g3597)));
	assign g3599 = (((g2052) & (g2674)));
	assign g3600 = (((!g2101) & (!g2134) & (!g3598) & (!g3599) & (!g2733) & (!g2785)) + ((!g2101) & (!g2134) & (!g3598) & (!g3599) & (!g2733) & (g2785)) + ((!g2101) & (!g2134) & (!g3598) & (!g3599) & (g2733) & (!g2785)) + ((!g2101) & (!g2134) & (!g3598) & (!g3599) & (g2733) & (g2785)) + ((!g2101) & (!g2134) & (!g3598) & (g3599) & (!g2733) & (!g2785)) + ((!g2101) & (!g2134) & (!g3598) & (g3599) & (!g2733) & (g2785)) + ((!g2101) & (!g2134) & (!g3598) & (g3599) & (g2733) & (!g2785)) + ((!g2101) & (!g2134) & (g3598) & (!g3599) & (!g2733) & (!g2785)) + ((!g2101) & (!g2134) & (g3598) & (!g3599) & (!g2733) & (g2785)) + ((!g2101) & (!g2134) & (g3598) & (!g3599) & (g2733) & (!g2785)) + ((!g2101) & (!g2134) & (g3598) & (g3599) & (!g2733) & (!g2785)) + ((!g2101) & (!g2134) & (g3598) & (g3599) & (!g2733) & (g2785)) + ((!g2101) & (!g2134) & (g3598) & (g3599) & (g2733) & (!g2785)) + ((!g2101) & (g2134) & (!g3598) & (!g3599) & (!g2733) & (!g2785)) + ((!g2101) & (g2134) & (!g3598) & (!g3599) & (g2733) & (!g2785)) + ((!g2101) & (g2134) & (!g3598) & (g3599) & (!g2733) & (!g2785)) + ((!g2101) & (g2134) & (g3598) & (!g3599) & (!g2733) & (!g2785)) + ((!g2101) & (g2134) & (g3598) & (g3599) & (!g2733) & (!g2785)) + ((g2101) & (!g2134) & (!g3598) & (!g3599) & (!g2733) & (!g2785)) + ((g2101) & (!g2134) & (!g3598) & (!g3599) & (!g2733) & (g2785)) + ((g2101) & (!g2134) & (!g3598) & (!g3599) & (g2733) & (!g2785)) + ((g2101) & (!g2134) & (!g3598) & (g3599) & (!g2733) & (!g2785)) + ((g2101) & (!g2134) & (!g3598) & (g3599) & (g2733) & (!g2785)) + ((g2101) & (!g2134) & (g3598) & (!g3599) & (!g2733) & (!g2785)) + ((g2101) & (!g2134) & (g3598) & (!g3599) & (g2733) & (!g2785)) + ((g2101) & (!g2134) & (g3598) & (g3599) & (!g2733) & (!g2785)) + ((g2101) & (!g2134) & (g3598) & (g3599) & (g2733) & (!g2785)) + ((g2101) & (g2134) & (!g3598) & (!g3599) & (!g2733) & (!g2785)));
	assign g3601 = (((!g2181) & (!g3600) & (g2822)) + ((g2181) & (!g3600) & (!g2822)) + ((g2181) & (!g3600) & (g2822)) + ((g2181) & (g3600) & (g2822)));
	assign g3602 = (((!g1892) & (!g2026) & (g2062) & (!g1894) & (!g2034) & (g2065)) + ((!g1892) & (!g2026) & (g2062) & (!g1894) & (g2034) & (g2065)) + ((!g1892) & (!g2026) & (g2062) & (g1894) & (!g2034) & (g2065)) + ((!g1892) & (!g2026) & (g2062) & (g1894) & (g2034) & (g2065)) + ((!g1892) & (g2026) & (!g2062) & (!g1894) & (g2034) & (g2065)) + ((!g1892) & (g2026) & (!g2062) & (g1894) & (g2034) & (g2065)) + ((!g1892) & (g2026) & (g2062) & (!g1894) & (!g2034) & (g2065)) + ((!g1892) & (g2026) & (g2062) & (!g1894) & (g2034) & (!g2065)) + ((!g1892) & (g2026) & (g2062) & (!g1894) & (g2034) & (g2065)) + ((!g1892) & (g2026) & (g2062) & (g1894) & (!g2034) & (g2065)) + ((!g1892) & (g2026) & (g2062) & (g1894) & (g2034) & (!g2065)) + ((!g1892) & (g2026) & (g2062) & (g1894) & (g2034) & (g2065)) + ((g1892) & (!g2026) & (!g2062) & (g1894) & (g2034) & (g2065)) + ((g1892) & (!g2026) & (g2062) & (!g1894) & (!g2034) & (g2065)) + ((g1892) & (!g2026) & (g2062) & (!g1894) & (g2034) & (g2065)) + ((g1892) & (!g2026) & (g2062) & (g1894) & (!g2034) & (g2065)) + ((g1892) & (!g2026) & (g2062) & (g1894) & (g2034) & (!g2065)) + ((g1892) & (!g2026) & (g2062) & (g1894) & (g2034) & (g2065)) + ((g1892) & (g2026) & (!g2062) & (!g1894) & (g2034) & (g2065)) + ((g1892) & (g2026) & (!g2062) & (g1894) & (!g2034) & (g2065)) + ((g1892) & (g2026) & (!g2062) & (g1894) & (g2034) & (g2065)) + ((g1892) & (g2026) & (g2062) & (!g1894) & (!g2034) & (g2065)) + ((g1892) & (g2026) & (g2062) & (!g1894) & (g2034) & (!g2065)) + ((g1892) & (g2026) & (g2062) & (!g1894) & (g2034) & (g2065)) + ((g1892) & (g2026) & (g2062) & (g1894) & (!g2034) & (!g2065)) + ((g1892) & (g2026) & (g2062) & (g1894) & (!g2034) & (g2065)) + ((g1892) & (g2026) & (g2062) & (g1894) & (g2034) & (!g2065)) + ((g1892) & (g2026) & (g2062) & (g1894) & (g2034) & (g2065)));
	assign g3603 = (((!g2188) & (g2196)) + ((g2188) & (!g2196)));
	assign g3604 = (((!g2108) & (!g2144) & (g2116) & (g2147) & (g3602) & (g3603)) + ((!g2108) & (g2144) & (!g2116) & (g2147) & (!g3602) & (g3603)) + ((!g2108) & (g2144) & (!g2116) & (g2147) & (g3602) & (g3603)) + ((!g2108) & (g2144) & (g2116) & (!g2147) & (g3602) & (g3603)) + ((!g2108) & (g2144) & (g2116) & (g2147) & (!g3602) & (g3603)) + ((!g2108) & (g2144) & (g2116) & (g2147) & (g3602) & (g3603)) + ((g2108) & (!g2144) & (!g2116) & (g2147) & (g3602) & (g3603)) + ((g2108) & (!g2144) & (g2116) & (g2147) & (!g3602) & (g3603)) + ((g2108) & (!g2144) & (g2116) & (g2147) & (g3602) & (g3603)) + ((g2108) & (g2144) & (!g2116) & (!g2147) & (g3602) & (g3603)) + ((g2108) & (g2144) & (!g2116) & (g2147) & (!g3602) & (g3603)) + ((g2108) & (g2144) & (!g2116) & (g2147) & (g3602) & (g3603)) + ((g2108) & (g2144) & (g2116) & (!g2147) & (!g3602) & (g3603)) + ((g2108) & (g2144) & (g2116) & (!g2147) & (g3602) & (g3603)) + ((g2108) & (g2144) & (g2116) & (g2147) & (!g3602) & (g3603)) + ((g2108) & (g2144) & (g2116) & (g2147) & (g3602) & (g3603)));
	assign g3605 = (((g2188) & (g2196)));
	assign g3606 = (((!g2224) & (!g2271) & (!g2227) & (!g2279) & (!g3604) & (!g3605)) + ((!g2224) & (!g2271) & (!g2227) & (!g2279) & (!g3604) & (g3605)) + ((!g2224) & (!g2271) & (!g2227) & (!g2279) & (g3604) & (!g3605)) + ((!g2224) & (!g2271) & (!g2227) & (!g2279) & (g3604) & (g3605)) + ((!g2224) & (!g2271) & (!g2227) & (g2279) & (!g3604) & (!g3605)) + ((!g2224) & (!g2271) & (!g2227) & (g2279) & (!g3604) & (g3605)) + ((!g2224) & (!g2271) & (!g2227) & (g2279) & (g3604) & (!g3605)) + ((!g2224) & (!g2271) & (!g2227) & (g2279) & (g3604) & (g3605)) + ((!g2224) & (!g2271) & (g2227) & (!g2279) & (!g3604) & (!g3605)) + ((!g2224) & (!g2271) & (g2227) & (!g2279) & (!g3604) & (g3605)) + ((!g2224) & (!g2271) & (g2227) & (!g2279) & (g3604) & (!g3605)) + ((!g2224) & (!g2271) & (g2227) & (!g2279) & (g3604) & (g3605)) + ((!g2224) & (!g2271) & (g2227) & (g2279) & (!g3604) & (!g3605)) + ((!g2224) & (g2271) & (!g2227) & (!g2279) & (!g3604) & (!g3605)) + ((!g2224) & (g2271) & (!g2227) & (!g2279) & (!g3604) & (g3605)) + ((!g2224) & (g2271) & (!g2227) & (!g2279) & (g3604) & (!g3605)) + ((!g2224) & (g2271) & (!g2227) & (!g2279) & (g3604) & (g3605)) + ((!g2224) & (g2271) & (g2227) & (!g2279) & (!g3604) & (!g3605)) + ((g2224) & (!g2271) & (!g2227) & (!g2279) & (!g3604) & (!g3605)) + ((g2224) & (!g2271) & (!g2227) & (!g2279) & (!g3604) & (g3605)) + ((g2224) & (!g2271) & (!g2227) & (!g2279) & (g3604) & (!g3605)) + ((g2224) & (!g2271) & (!g2227) & (!g2279) & (g3604) & (g3605)) + ((g2224) & (!g2271) & (!g2227) & (g2279) & (!g3604) & (!g3605)) + ((g2224) & (!g2271) & (g2227) & (!g2279) & (!g3604) & (!g3605)) + ((g2224) & (!g2271) & (g2227) & (!g2279) & (!g3604) & (g3605)) + ((g2224) & (!g2271) & (g2227) & (!g2279) & (g3604) & (!g3605)) + ((g2224) & (!g2271) & (g2227) & (!g2279) & (g3604) & (g3605)) + ((g2224) & (g2271) & (!g2227) & (!g2279) & (!g3604) & (!g3605)));
	assign g3607 = (((!g2390) & (g2393)) + ((g2390) & (!g2393)));
	assign g3608 = (((!g2311) & (!g2354) & (g2314) & (g2362) & (!g3606) & (g3607)) + ((!g2311) & (g2354) & (!g2314) & (g2362) & (!g3606) & (g3607)) + ((!g2311) & (g2354) & (!g2314) & (g2362) & (g3606) & (g3607)) + ((!g2311) & (g2354) & (g2314) & (!g2362) & (!g3606) & (g3607)) + ((!g2311) & (g2354) & (g2314) & (g2362) & (!g3606) & (g3607)) + ((!g2311) & (g2354) & (g2314) & (g2362) & (g3606) & (g3607)) + ((g2311) & (!g2354) & (!g2314) & (g2362) & (!g3606) & (g3607)) + ((g2311) & (!g2354) & (g2314) & (g2362) & (!g3606) & (g3607)) + ((g2311) & (!g2354) & (g2314) & (g2362) & (g3606) & (g3607)) + ((g2311) & (g2354) & (!g2314) & (!g2362) & (!g3606) & (g3607)) + ((g2311) & (g2354) & (!g2314) & (g2362) & (!g3606) & (g3607)) + ((g2311) & (g2354) & (!g2314) & (g2362) & (g3606) & (g3607)) + ((g2311) & (g2354) & (g2314) & (!g2362) & (!g3606) & (g3607)) + ((g2311) & (g2354) & (g2314) & (!g2362) & (g3606) & (g3607)) + ((g2311) & (g2354) & (g2314) & (g2362) & (!g3606) & (g3607)) + ((g2311) & (g2354) & (g2314) & (g2362) & (g3606) & (g3607)));
	assign g3609 = (((g2390) & (g2393)));
	assign g3610 = (((!g2450) & (!g2527) & (!g2474) & (!g2529) & (!g3608) & (!g3609)) + ((!g2450) & (!g2527) & (!g2474) & (!g2529) & (!g3608) & (g3609)) + ((!g2450) & (!g2527) & (!g2474) & (!g2529) & (g3608) & (!g3609)) + ((!g2450) & (!g2527) & (!g2474) & (!g2529) & (g3608) & (g3609)) + ((!g2450) & (!g2527) & (!g2474) & (g2529) & (!g3608) & (!g3609)) + ((!g2450) & (!g2527) & (!g2474) & (g2529) & (!g3608) & (g3609)) + ((!g2450) & (!g2527) & (!g2474) & (g2529) & (g3608) & (!g3609)) + ((!g2450) & (!g2527) & (!g2474) & (g2529) & (g3608) & (g3609)) + ((!g2450) & (!g2527) & (g2474) & (!g2529) & (!g3608) & (!g3609)) + ((!g2450) & (!g2527) & (g2474) & (!g2529) & (!g3608) & (g3609)) + ((!g2450) & (!g2527) & (g2474) & (!g2529) & (g3608) & (!g3609)) + ((!g2450) & (!g2527) & (g2474) & (!g2529) & (g3608) & (g3609)) + ((!g2450) & (!g2527) & (g2474) & (g2529) & (!g3608) & (!g3609)) + ((!g2450) & (g2527) & (!g2474) & (!g2529) & (!g3608) & (!g3609)) + ((!g2450) & (g2527) & (!g2474) & (!g2529) & (!g3608) & (g3609)) + ((!g2450) & (g2527) & (!g2474) & (!g2529) & (g3608) & (!g3609)) + ((!g2450) & (g2527) & (!g2474) & (!g2529) & (g3608) & (g3609)) + ((!g2450) & (g2527) & (g2474) & (!g2529) & (!g3608) & (!g3609)) + ((g2450) & (!g2527) & (!g2474) & (!g2529) & (!g3608) & (!g3609)) + ((g2450) & (!g2527) & (!g2474) & (!g2529) & (!g3608) & (g3609)) + ((g2450) & (!g2527) & (!g2474) & (!g2529) & (g3608) & (!g3609)) + ((g2450) & (!g2527) & (!g2474) & (!g2529) & (g3608) & (g3609)) + ((g2450) & (!g2527) & (!g2474) & (g2529) & (!g3608) & (!g3609)) + ((g2450) & (!g2527) & (g2474) & (!g2529) & (!g3608) & (!g3609)) + ((g2450) & (!g2527) & (g2474) & (!g2529) & (!g3608) & (g3609)) + ((g2450) & (!g2527) & (g2474) & (!g2529) & (g3608) & (!g3609)) + ((g2450) & (!g2527) & (g2474) & (!g2529) & (g3608) & (g3609)) + ((g2450) & (g2527) & (!g2474) & (!g2529) & (!g3608) & (!g3609)));
	assign g3611 = (((!g2450) & (!g2474) & (!g3608) & (!g3609) & (!g5800) & (g5801)) + ((!g2450) & (!g2474) & (!g3608) & (g3609) & (!g5800) & (g5801)) + ((!g2450) & (!g2474) & (g3608) & (!g3609) & (!g5800) & (g5801)) + ((!g2450) & (!g2474) & (g3608) & (g3609) & (!g5800) & (g5801)) + ((!g2450) & (g2474) & (!g3608) & (!g3609) & (!g5800) & (g5801)) + ((!g2450) & (g2474) & (!g3608) & (g3609) & (!g5800) & (g5801)) + ((!g2450) & (g2474) & (!g3608) & (g3609) & (g5800) & (g5801)) + ((!g2450) & (g2474) & (g3608) & (!g3609) & (!g5800) & (g5801)) + ((!g2450) & (g2474) & (g3608) & (!g3609) & (g5800) & (g5801)) + ((!g2450) & (g2474) & (g3608) & (g3609) & (!g5800) & (g5801)) + ((!g2450) & (g2474) & (g3608) & (g3609) & (g5800) & (g5801)) + ((g2450) & (!g2474) & (!g3608) & (!g3609) & (!g5800) & (g5801)) + ((g2450) & (!g2474) & (!g3608) & (g3609) & (!g5800) & (g5801)) + ((g2450) & (!g2474) & (!g3608) & (g3609) & (g5800) & (g5801)) + ((g2450) & (!g2474) & (g3608) & (!g3609) & (!g5800) & (g5801)) + ((g2450) & (!g2474) & (g3608) & (!g3609) & (g5800) & (g5801)) + ((g2450) & (!g2474) & (g3608) & (g3609) & (!g5800) & (g5801)) + ((g2450) & (!g2474) & (g3608) & (g3609) & (g5800) & (g5801)) + ((g2450) & (g2474) & (!g3608) & (!g3609) & (!g5800) & (g5801)) + ((g2450) & (g2474) & (!g3608) & (!g3609) & (g5800) & (g5801)) + ((g2450) & (g2474) & (!g3608) & (g3609) & (!g5800) & (g5801)) + ((g2450) & (g2474) & (!g3608) & (g3609) & (g5800) & (g5801)) + ((g2450) & (g2474) & (g3608) & (!g3609) & (!g5800) & (g5801)) + ((g2450) & (g2474) & (g3608) & (!g3609) & (g5800) & (g5801)) + ((g2450) & (g2474) & (g3608) & (g3609) & (!g5800) & (g5801)) + ((g2450) & (g2474) & (g3608) & (g3609) & (g5800) & (g5801)));
	assign g3612 = (((g2657) & (g2665)));
	assign g3613 = (((!g2703) & (!g2768) & (!g2708) & (!g2776) & (!g3611) & (!g3612)) + ((!g2703) & (!g2768) & (!g2708) & (!g2776) & (!g3611) & (g3612)) + ((!g2703) & (!g2768) & (!g2708) & (!g2776) & (g3611) & (!g3612)) + ((!g2703) & (!g2768) & (!g2708) & (!g2776) & (g3611) & (g3612)) + ((!g2703) & (!g2768) & (!g2708) & (g2776) & (!g3611) & (!g3612)) + ((!g2703) & (!g2768) & (!g2708) & (g2776) & (!g3611) & (g3612)) + ((!g2703) & (!g2768) & (!g2708) & (g2776) & (g3611) & (!g3612)) + ((!g2703) & (!g2768) & (!g2708) & (g2776) & (g3611) & (g3612)) + ((!g2703) & (!g2768) & (g2708) & (!g2776) & (!g3611) & (!g3612)) + ((!g2703) & (!g2768) & (g2708) & (!g2776) & (!g3611) & (g3612)) + ((!g2703) & (!g2768) & (g2708) & (!g2776) & (g3611) & (!g3612)) + ((!g2703) & (!g2768) & (g2708) & (!g2776) & (g3611) & (g3612)) + ((!g2703) & (!g2768) & (g2708) & (g2776) & (!g3611) & (!g3612)) + ((!g2703) & (g2768) & (!g2708) & (!g2776) & (!g3611) & (!g3612)) + ((!g2703) & (g2768) & (!g2708) & (!g2776) & (!g3611) & (g3612)) + ((!g2703) & (g2768) & (!g2708) & (!g2776) & (g3611) & (!g3612)) + ((!g2703) & (g2768) & (!g2708) & (!g2776) & (g3611) & (g3612)) + ((!g2703) & (g2768) & (g2708) & (!g2776) & (!g3611) & (!g3612)) + ((g2703) & (!g2768) & (!g2708) & (!g2776) & (!g3611) & (!g3612)) + ((g2703) & (!g2768) & (!g2708) & (!g2776) & (!g3611) & (g3612)) + ((g2703) & (!g2768) & (!g2708) & (!g2776) & (g3611) & (!g3612)) + ((g2703) & (!g2768) & (!g2708) & (!g2776) & (g3611) & (g3612)) + ((g2703) & (!g2768) & (!g2708) & (g2776) & (!g3611) & (!g3612)) + ((g2703) & (!g2768) & (g2708) & (!g2776) & (!g3611) & (!g3612)) + ((g2703) & (!g2768) & (g2708) & (!g2776) & (!g3611) & (g3612)) + ((g2703) & (!g2768) & (g2708) & (!g2776) & (g3611) & (!g3612)) + ((g2703) & (!g2768) & (g2708) & (!g2776) & (g3611) & (g3612)) + ((g2703) & (g2768) & (!g2708) & (!g2776) & (!g3611) & (!g3612)));
	assign g3614 = (((!g2885) & (g2887)) + ((g2885) & (!g2887)));
	assign g3615 = (((!g2804) & (!g2845) & (g2807) & (g2857) & (!g3613) & (g3614)) + ((!g2804) & (g2845) & (!g2807) & (g2857) & (!g3613) & (g3614)) + ((!g2804) & (g2845) & (!g2807) & (g2857) & (g3613) & (g3614)) + ((!g2804) & (g2845) & (g2807) & (!g2857) & (!g3613) & (g3614)) + ((!g2804) & (g2845) & (g2807) & (g2857) & (!g3613) & (g3614)) + ((!g2804) & (g2845) & (g2807) & (g2857) & (g3613) & (g3614)) + ((g2804) & (!g2845) & (!g2807) & (g2857) & (!g3613) & (g3614)) + ((g2804) & (!g2845) & (g2807) & (g2857) & (!g3613) & (g3614)) + ((g2804) & (!g2845) & (g2807) & (g2857) & (g3613) & (g3614)) + ((g2804) & (g2845) & (!g2807) & (!g2857) & (!g3613) & (g3614)) + ((g2804) & (g2845) & (!g2807) & (g2857) & (!g3613) & (g3614)) + ((g2804) & (g2845) & (!g2807) & (g2857) & (g3613) & (g3614)) + ((g2804) & (g2845) & (g2807) & (!g2857) & (!g3613) & (g3614)) + ((g2804) & (g2845) & (g2807) & (!g2857) & (g3613) & (g3614)) + ((g2804) & (g2845) & (g2807) & (g2857) & (!g3613) & (g3614)) + ((g2804) & (g2845) & (g2807) & (g2857) & (g3613) & (g3614)));
	assign g3616 = (((g2885) & (g2887)));
	assign g3617 = (((!g2932) & (!g3003) & (!g3615) & (!g3616) & (!g2956) & (!g3005)) + ((!g2932) & (!g3003) & (!g3615) & (!g3616) & (!g2956) & (g3005)) + ((!g2932) & (!g3003) & (!g3615) & (!g3616) & (g2956) & (!g3005)) + ((!g2932) & (!g3003) & (!g3615) & (!g3616) & (g2956) & (g3005)) + ((!g2932) & (!g3003) & (!g3615) & (g3616) & (!g2956) & (!g3005)) + ((!g2932) & (!g3003) & (!g3615) & (g3616) & (!g2956) & (g3005)) + ((!g2932) & (!g3003) & (!g3615) & (g3616) & (g2956) & (!g3005)) + ((!g2932) & (!g3003) & (g3615) & (!g3616) & (!g2956) & (!g3005)) + ((!g2932) & (!g3003) & (g3615) & (!g3616) & (!g2956) & (g3005)) + ((!g2932) & (!g3003) & (g3615) & (!g3616) & (g2956) & (!g3005)) + ((!g2932) & (!g3003) & (g3615) & (g3616) & (!g2956) & (!g3005)) + ((!g2932) & (!g3003) & (g3615) & (g3616) & (!g2956) & (g3005)) + ((!g2932) & (!g3003) & (g3615) & (g3616) & (g2956) & (!g3005)) + ((!g2932) & (g3003) & (!g3615) & (!g3616) & (!g2956) & (!g3005)) + ((!g2932) & (g3003) & (!g3615) & (!g3616) & (g2956) & (!g3005)) + ((!g2932) & (g3003) & (!g3615) & (g3616) & (!g2956) & (!g3005)) + ((!g2932) & (g3003) & (g3615) & (!g3616) & (!g2956) & (!g3005)) + ((!g2932) & (g3003) & (g3615) & (g3616) & (!g2956) & (!g3005)) + ((g2932) & (!g3003) & (!g3615) & (!g3616) & (!g2956) & (!g3005)) + ((g2932) & (!g3003) & (!g3615) & (!g3616) & (!g2956) & (g3005)) + ((g2932) & (!g3003) & (!g3615) & (!g3616) & (g2956) & (!g3005)) + ((g2932) & (!g3003) & (!g3615) & (g3616) & (!g2956) & (!g3005)) + ((g2932) & (!g3003) & (!g3615) & (g3616) & (g2956) & (!g3005)) + ((g2932) & (!g3003) & (g3615) & (!g3616) & (!g2956) & (!g3005)) + ((g2932) & (!g3003) & (g3615) & (!g3616) & (g2956) & (!g3005)) + ((g2932) & (!g3003) & (g3615) & (g3616) & (!g2956) & (!g3005)) + ((g2932) & (!g3003) & (g3615) & (g3616) & (g2956) & (!g3005)) + ((g2932) & (g3003) & (!g3615) & (!g3616) & (!g2956) & (!g3005)));
	assign g3618 = (((!g3038) & (!g3617) & (g3050)) + ((g3038) & (!g3617) & (!g3050)) + ((g3038) & (!g3617) & (g3050)) + ((g3038) & (g3617) & (g3050)));
	assign g3619 = (((!g3618) & (g3078) & (g3080)) + ((g3618) & (!g3078) & (g3080)) + ((g3618) & (g3078) & (!g3080)) + ((g3618) & (g3078) & (g3080)));
	assign g3620 = (((!g830) & (!g1896) & (!g7029) & (key[224])) + ((!g830) & (!g1896) & (g7029) & (key[224])) + ((!g830) & (g1896) & (!g7029) & (key[224])) + ((!g830) & (g1896) & (g7029) & (key[224])) + ((g830) & (!g1896) & (g7029) & (!key[224])) + ((g830) & (!g1896) & (g7029) & (key[224])) + ((g830) & (g1896) & (!g7029) & (!key[224])) + ((g830) & (g1896) & (!g7029) & (key[224])));
	assign g3621 = (((!g1906) & (!g1940) & (g1942) & (!g828) & (!g864) & (g897)) + ((!g1906) & (!g1940) & (g1942) & (!g828) & (g864) & (g897)) + ((!g1906) & (!g1940) & (g1942) & (g828) & (!g864) & (g897)) + ((!g1906) & (!g1940) & (g1942) & (g828) & (g864) & (g897)) + ((!g1906) & (g1940) & (!g1942) & (!g828) & (g864) & (g897)) + ((!g1906) & (g1940) & (!g1942) & (g828) & (g864) & (g897)) + ((!g1906) & (g1940) & (g1942) & (!g828) & (!g864) & (g897)) + ((!g1906) & (g1940) & (g1942) & (!g828) & (g864) & (!g897)) + ((!g1906) & (g1940) & (g1942) & (!g828) & (g864) & (g897)) + ((!g1906) & (g1940) & (g1942) & (g828) & (!g864) & (g897)) + ((!g1906) & (g1940) & (g1942) & (g828) & (g864) & (!g897)) + ((!g1906) & (g1940) & (g1942) & (g828) & (g864) & (g897)) + ((g1906) & (!g1940) & (!g1942) & (g828) & (g864) & (g897)) + ((g1906) & (!g1940) & (g1942) & (!g828) & (!g864) & (g897)) + ((g1906) & (!g1940) & (g1942) & (!g828) & (g864) & (g897)) + ((g1906) & (!g1940) & (g1942) & (g828) & (!g864) & (g897)) + ((g1906) & (!g1940) & (g1942) & (g828) & (g864) & (!g897)) + ((g1906) & (!g1940) & (g1942) & (g828) & (g864) & (g897)) + ((g1906) & (g1940) & (!g1942) & (!g828) & (g864) & (g897)) + ((g1906) & (g1940) & (!g1942) & (g828) & (!g864) & (g897)) + ((g1906) & (g1940) & (!g1942) & (g828) & (g864) & (g897)) + ((g1906) & (g1940) & (g1942) & (!g828) & (!g864) & (g897)) + ((g1906) & (g1940) & (g1942) & (!g828) & (g864) & (!g897)) + ((g1906) & (g1940) & (g1942) & (!g828) & (g864) & (g897)) + ((g1906) & (g1940) & (g1942) & (g828) & (!g864) & (!g897)) + ((g1906) & (g1940) & (g1942) & (g828) & (!g864) & (g897)) + ((g1906) & (g1940) & (g1942) & (g828) & (g864) & (!g897)) + ((g1906) & (g1940) & (g1942) & (g828) & (g864) & (g897)));
	assign g3622 = (((!g1949) & (g998)) + ((g1949) & (!g998)));
	assign g3623 = (((!g1945) & (!g1947) & (g931) & (g964) & (g3621) & (g3622)) + ((!g1945) & (g1947) & (!g931) & (g964) & (!g3621) & (g3622)) + ((!g1945) & (g1947) & (!g931) & (g964) & (g3621) & (g3622)) + ((!g1945) & (g1947) & (g931) & (!g964) & (g3621) & (g3622)) + ((!g1945) & (g1947) & (g931) & (g964) & (!g3621) & (g3622)) + ((!g1945) & (g1947) & (g931) & (g964) & (g3621) & (g3622)) + ((g1945) & (!g1947) & (!g931) & (g964) & (g3621) & (g3622)) + ((g1945) & (!g1947) & (g931) & (g964) & (!g3621) & (g3622)) + ((g1945) & (!g1947) & (g931) & (g964) & (g3621) & (g3622)) + ((g1945) & (g1947) & (!g931) & (!g964) & (g3621) & (g3622)) + ((g1945) & (g1947) & (!g931) & (g964) & (!g3621) & (g3622)) + ((g1945) & (g1947) & (!g931) & (g964) & (g3621) & (g3622)) + ((g1945) & (g1947) & (g931) & (!g964) & (!g3621) & (g3622)) + ((g1945) & (g1947) & (g931) & (!g964) & (g3621) & (g3622)) + ((g1945) & (g1947) & (g931) & (g964) & (!g3621) & (g3622)) + ((g1945) & (g1947) & (g931) & (g964) & (g3621) & (g3622)));
	assign g3624 = (((g1949) & (g998)));
	assign g3625 = (((!g1954) & (!g1956) & (!g1031) & (!g1065) & (!g3623) & (!g3624)) + ((!g1954) & (!g1956) & (!g1031) & (!g1065) & (!g3623) & (g3624)) + ((!g1954) & (!g1956) & (!g1031) & (!g1065) & (g3623) & (!g3624)) + ((!g1954) & (!g1956) & (!g1031) & (!g1065) & (g3623) & (g3624)) + ((!g1954) & (!g1956) & (!g1031) & (g1065) & (!g3623) & (!g3624)) + ((!g1954) & (!g1956) & (!g1031) & (g1065) & (!g3623) & (g3624)) + ((!g1954) & (!g1956) & (!g1031) & (g1065) & (g3623) & (!g3624)) + ((!g1954) & (!g1956) & (!g1031) & (g1065) & (g3623) & (g3624)) + ((!g1954) & (!g1956) & (g1031) & (!g1065) & (!g3623) & (!g3624)) + ((!g1954) & (!g1956) & (g1031) & (!g1065) & (!g3623) & (g3624)) + ((!g1954) & (!g1956) & (g1031) & (!g1065) & (g3623) & (!g3624)) + ((!g1954) & (!g1956) & (g1031) & (!g1065) & (g3623) & (g3624)) + ((!g1954) & (!g1956) & (g1031) & (g1065) & (!g3623) & (!g3624)) + ((!g1954) & (g1956) & (!g1031) & (!g1065) & (!g3623) & (!g3624)) + ((!g1954) & (g1956) & (!g1031) & (!g1065) & (!g3623) & (g3624)) + ((!g1954) & (g1956) & (!g1031) & (!g1065) & (g3623) & (!g3624)) + ((!g1954) & (g1956) & (!g1031) & (!g1065) & (g3623) & (g3624)) + ((!g1954) & (g1956) & (g1031) & (!g1065) & (!g3623) & (!g3624)) + ((g1954) & (!g1956) & (!g1031) & (!g1065) & (!g3623) & (!g3624)) + ((g1954) & (!g1956) & (!g1031) & (!g1065) & (!g3623) & (g3624)) + ((g1954) & (!g1956) & (!g1031) & (!g1065) & (g3623) & (!g3624)) + ((g1954) & (!g1956) & (!g1031) & (!g1065) & (g3623) & (g3624)) + ((g1954) & (!g1956) & (!g1031) & (g1065) & (!g3623) & (!g3624)) + ((g1954) & (!g1956) & (g1031) & (!g1065) & (!g3623) & (!g3624)) + ((g1954) & (!g1956) & (g1031) & (!g1065) & (!g3623) & (g3624)) + ((g1954) & (!g1956) & (g1031) & (!g1065) & (g3623) & (!g3624)) + ((g1954) & (!g1956) & (g1031) & (!g1065) & (g3623) & (g3624)) + ((g1954) & (g1956) & (!g1031) & (!g1065) & (!g3623) & (!g3624)));
	assign g3626 = (((!g1963) & (g1165)) + ((g1963) & (!g1165)));
	assign g3627 = (((!g1959) & (!g1961) & (g1098) & (g1132) & (!g3625) & (g3626)) + ((!g1959) & (g1961) & (!g1098) & (g1132) & (!g3625) & (g3626)) + ((!g1959) & (g1961) & (!g1098) & (g1132) & (g3625) & (g3626)) + ((!g1959) & (g1961) & (g1098) & (!g1132) & (!g3625) & (g3626)) + ((!g1959) & (g1961) & (g1098) & (g1132) & (!g3625) & (g3626)) + ((!g1959) & (g1961) & (g1098) & (g1132) & (g3625) & (g3626)) + ((g1959) & (!g1961) & (!g1098) & (g1132) & (!g3625) & (g3626)) + ((g1959) & (!g1961) & (g1098) & (g1132) & (!g3625) & (g3626)) + ((g1959) & (!g1961) & (g1098) & (g1132) & (g3625) & (g3626)) + ((g1959) & (g1961) & (!g1098) & (!g1132) & (!g3625) & (g3626)) + ((g1959) & (g1961) & (!g1098) & (g1132) & (!g3625) & (g3626)) + ((g1959) & (g1961) & (!g1098) & (g1132) & (g3625) & (g3626)) + ((g1959) & (g1961) & (g1098) & (!g1132) & (!g3625) & (g3626)) + ((g1959) & (g1961) & (g1098) & (!g1132) & (g3625) & (g3626)) + ((g1959) & (g1961) & (g1098) & (g1132) & (!g3625) & (g3626)) + ((g1959) & (g1961) & (g1098) & (g1132) & (g3625) & (g3626)));
	assign g3628 = (((g1963) & (g1165)));
	assign g3629 = (((!g1968) & (!g1970) & (!g1199) & (!g1236) & (!g3627) & (!g3628)) + ((!g1968) & (!g1970) & (!g1199) & (!g1236) & (!g3627) & (g3628)) + ((!g1968) & (!g1970) & (!g1199) & (!g1236) & (g3627) & (!g3628)) + ((!g1968) & (!g1970) & (!g1199) & (!g1236) & (g3627) & (g3628)) + ((!g1968) & (!g1970) & (!g1199) & (g1236) & (!g3627) & (!g3628)) + ((!g1968) & (!g1970) & (!g1199) & (g1236) & (!g3627) & (g3628)) + ((!g1968) & (!g1970) & (!g1199) & (g1236) & (g3627) & (!g3628)) + ((!g1968) & (!g1970) & (!g1199) & (g1236) & (g3627) & (g3628)) + ((!g1968) & (!g1970) & (g1199) & (!g1236) & (!g3627) & (!g3628)) + ((!g1968) & (!g1970) & (g1199) & (!g1236) & (!g3627) & (g3628)) + ((!g1968) & (!g1970) & (g1199) & (!g1236) & (g3627) & (!g3628)) + ((!g1968) & (!g1970) & (g1199) & (!g1236) & (g3627) & (g3628)) + ((!g1968) & (!g1970) & (g1199) & (g1236) & (!g3627) & (!g3628)) + ((!g1968) & (g1970) & (!g1199) & (!g1236) & (!g3627) & (!g3628)) + ((!g1968) & (g1970) & (!g1199) & (!g1236) & (!g3627) & (g3628)) + ((!g1968) & (g1970) & (!g1199) & (!g1236) & (g3627) & (!g3628)) + ((!g1968) & (g1970) & (!g1199) & (!g1236) & (g3627) & (g3628)) + ((!g1968) & (g1970) & (g1199) & (!g1236) & (!g3627) & (!g3628)) + ((g1968) & (!g1970) & (!g1199) & (!g1236) & (!g3627) & (!g3628)) + ((g1968) & (!g1970) & (!g1199) & (!g1236) & (!g3627) & (g3628)) + ((g1968) & (!g1970) & (!g1199) & (!g1236) & (g3627) & (!g3628)) + ((g1968) & (!g1970) & (!g1199) & (!g1236) & (g3627) & (g3628)) + ((g1968) & (!g1970) & (!g1199) & (g1236) & (!g3627) & (!g3628)) + ((g1968) & (!g1970) & (g1199) & (!g1236) & (!g3627) & (!g3628)) + ((g1968) & (!g1970) & (g1199) & (!g1236) & (!g3627) & (g3628)) + ((g1968) & (!g1970) & (g1199) & (!g1236) & (g3627) & (!g3628)) + ((g1968) & (!g1970) & (g1199) & (!g1236) & (g3627) & (g3628)) + ((g1968) & (g1970) & (!g1199) & (!g1236) & (!g3627) & (!g3628)));
	assign g3630 = (((!g1968) & (!g1199) & (!g3627) & (!g3628) & (!g5803) & (g5804)) + ((!g1968) & (!g1199) & (!g3627) & (g3628) & (!g5803) & (g5804)) + ((!g1968) & (!g1199) & (g3627) & (!g3628) & (!g5803) & (g5804)) + ((!g1968) & (!g1199) & (g3627) & (g3628) & (!g5803) & (g5804)) + ((!g1968) & (g1199) & (!g3627) & (!g3628) & (!g5803) & (g5804)) + ((!g1968) & (g1199) & (!g3627) & (g3628) & (!g5803) & (g5804)) + ((!g1968) & (g1199) & (!g3627) & (g3628) & (g5803) & (g5804)) + ((!g1968) & (g1199) & (g3627) & (!g3628) & (!g5803) & (g5804)) + ((!g1968) & (g1199) & (g3627) & (!g3628) & (g5803) & (g5804)) + ((!g1968) & (g1199) & (g3627) & (g3628) & (!g5803) & (g5804)) + ((!g1968) & (g1199) & (g3627) & (g3628) & (g5803) & (g5804)) + ((g1968) & (!g1199) & (!g3627) & (!g3628) & (!g5803) & (g5804)) + ((g1968) & (!g1199) & (!g3627) & (g3628) & (!g5803) & (g5804)) + ((g1968) & (!g1199) & (!g3627) & (g3628) & (g5803) & (g5804)) + ((g1968) & (!g1199) & (g3627) & (!g3628) & (!g5803) & (g5804)) + ((g1968) & (!g1199) & (g3627) & (!g3628) & (g5803) & (g5804)) + ((g1968) & (!g1199) & (g3627) & (g3628) & (!g5803) & (g5804)) + ((g1968) & (!g1199) & (g3627) & (g3628) & (g5803) & (g5804)) + ((g1968) & (g1199) & (!g3627) & (!g3628) & (!g5803) & (g5804)) + ((g1968) & (g1199) & (!g3627) & (!g3628) & (g5803) & (g5804)) + ((g1968) & (g1199) & (!g3627) & (g3628) & (!g5803) & (g5804)) + ((g1968) & (g1199) & (!g3627) & (g3628) & (g5803) & (g5804)) + ((g1968) & (g1199) & (g3627) & (!g3628) & (!g5803) & (g5804)) + ((g1968) & (g1199) & (g3627) & (!g3628) & (g5803) & (g5804)) + ((g1968) & (g1199) & (g3627) & (g3628) & (!g5803) & (g5804)) + ((g1968) & (g1199) & (g3627) & (g3628) & (g5803) & (g5804)));
	assign g3631 = (((g2048) & (g1337)));
	assign g3632 = (((!g2099) & (!g2130) & (!g1370) & (!g1406) & (!g3630) & (!g3631)) + ((!g2099) & (!g2130) & (!g1370) & (!g1406) & (!g3630) & (g3631)) + ((!g2099) & (!g2130) & (!g1370) & (!g1406) & (g3630) & (!g3631)) + ((!g2099) & (!g2130) & (!g1370) & (!g1406) & (g3630) & (g3631)) + ((!g2099) & (!g2130) & (!g1370) & (g1406) & (!g3630) & (!g3631)) + ((!g2099) & (!g2130) & (!g1370) & (g1406) & (!g3630) & (g3631)) + ((!g2099) & (!g2130) & (!g1370) & (g1406) & (g3630) & (!g3631)) + ((!g2099) & (!g2130) & (!g1370) & (g1406) & (g3630) & (g3631)) + ((!g2099) & (!g2130) & (g1370) & (!g1406) & (!g3630) & (!g3631)) + ((!g2099) & (!g2130) & (g1370) & (!g1406) & (!g3630) & (g3631)) + ((!g2099) & (!g2130) & (g1370) & (!g1406) & (g3630) & (!g3631)) + ((!g2099) & (!g2130) & (g1370) & (!g1406) & (g3630) & (g3631)) + ((!g2099) & (!g2130) & (g1370) & (g1406) & (!g3630) & (!g3631)) + ((!g2099) & (g2130) & (!g1370) & (!g1406) & (!g3630) & (!g3631)) + ((!g2099) & (g2130) & (!g1370) & (!g1406) & (!g3630) & (g3631)) + ((!g2099) & (g2130) & (!g1370) & (!g1406) & (g3630) & (!g3631)) + ((!g2099) & (g2130) & (!g1370) & (!g1406) & (g3630) & (g3631)) + ((!g2099) & (g2130) & (g1370) & (!g1406) & (!g3630) & (!g3631)) + ((g2099) & (!g2130) & (!g1370) & (!g1406) & (!g3630) & (!g3631)) + ((g2099) & (!g2130) & (!g1370) & (!g1406) & (!g3630) & (g3631)) + ((g2099) & (!g2130) & (!g1370) & (!g1406) & (g3630) & (!g3631)) + ((g2099) & (!g2130) & (!g1370) & (!g1406) & (g3630) & (g3631)) + ((g2099) & (!g2130) & (!g1370) & (g1406) & (!g3630) & (!g3631)) + ((g2099) & (!g2130) & (g1370) & (!g1406) & (!g3630) & (!g3631)) + ((g2099) & (!g2130) & (g1370) & (!g1406) & (!g3630) & (g3631)) + ((g2099) & (!g2130) & (g1370) & (!g1406) & (g3630) & (!g3631)) + ((g2099) & (!g2130) & (g1370) & (!g1406) & (g3630) & (g3631)) + ((g2099) & (g2130) & (!g1370) & (!g1406) & (!g3630) & (!g3631)));
	assign g3633 = (((!g2257) & (g1507)) + ((g2257) & (!g1507)));
	assign g3634 = (((!g2178) & (!g2211) & (g1439) & (g1473) & (!g3632) & (g3633)) + ((!g2178) & (g2211) & (!g1439) & (g1473) & (!g3632) & (g3633)) + ((!g2178) & (g2211) & (!g1439) & (g1473) & (g3632) & (g3633)) + ((!g2178) & (g2211) & (g1439) & (!g1473) & (!g3632) & (g3633)) + ((!g2178) & (g2211) & (g1439) & (g1473) & (!g3632) & (g3633)) + ((!g2178) & (g2211) & (g1439) & (g1473) & (g3632) & (g3633)) + ((g2178) & (!g2211) & (!g1439) & (g1473) & (!g3632) & (g3633)) + ((g2178) & (!g2211) & (g1439) & (g1473) & (!g3632) & (g3633)) + ((g2178) & (!g2211) & (g1439) & (g1473) & (g3632) & (g3633)) + ((g2178) & (g2211) & (!g1439) & (!g1473) & (!g3632) & (g3633)) + ((g2178) & (g2211) & (!g1439) & (g1473) & (!g3632) & (g3633)) + ((g2178) & (g2211) & (!g1439) & (g1473) & (g3632) & (g3633)) + ((g2178) & (g2211) & (g1439) & (!g1473) & (!g3632) & (g3633)) + ((g2178) & (g2211) & (g1439) & (!g1473) & (g3632) & (g3633)) + ((g2178) & (g2211) & (g1439) & (g1473) & (!g3632) & (g3633)) + ((g2178) & (g2211) & (g1439) & (g1473) & (g3632) & (g3633)));
	assign g3635 = (((g2257) & (g1507)));
	assign g3636 = (((!g2296) & (!g2344) & (!g1540) & (!g1577) & (!g3634) & (!g3635)) + ((!g2296) & (!g2344) & (!g1540) & (!g1577) & (!g3634) & (g3635)) + ((!g2296) & (!g2344) & (!g1540) & (!g1577) & (g3634) & (!g3635)) + ((!g2296) & (!g2344) & (!g1540) & (!g1577) & (g3634) & (g3635)) + ((!g2296) & (!g2344) & (!g1540) & (g1577) & (!g3634) & (!g3635)) + ((!g2296) & (!g2344) & (!g1540) & (g1577) & (!g3634) & (g3635)) + ((!g2296) & (!g2344) & (!g1540) & (g1577) & (g3634) & (!g3635)) + ((!g2296) & (!g2344) & (!g1540) & (g1577) & (g3634) & (g3635)) + ((!g2296) & (!g2344) & (g1540) & (!g1577) & (!g3634) & (!g3635)) + ((!g2296) & (!g2344) & (g1540) & (!g1577) & (!g3634) & (g3635)) + ((!g2296) & (!g2344) & (g1540) & (!g1577) & (g3634) & (!g3635)) + ((!g2296) & (!g2344) & (g1540) & (!g1577) & (g3634) & (g3635)) + ((!g2296) & (!g2344) & (g1540) & (g1577) & (!g3634) & (!g3635)) + ((!g2296) & (g2344) & (!g1540) & (!g1577) & (!g3634) & (!g3635)) + ((!g2296) & (g2344) & (!g1540) & (!g1577) & (!g3634) & (g3635)) + ((!g2296) & (g2344) & (!g1540) & (!g1577) & (g3634) & (!g3635)) + ((!g2296) & (g2344) & (!g1540) & (!g1577) & (g3634) & (g3635)) + ((!g2296) & (g2344) & (g1540) & (!g1577) & (!g3634) & (!g3635)) + ((g2296) & (!g2344) & (!g1540) & (!g1577) & (!g3634) & (!g3635)) + ((g2296) & (!g2344) & (!g1540) & (!g1577) & (!g3634) & (g3635)) + ((g2296) & (!g2344) & (!g1540) & (!g1577) & (g3634) & (!g3635)) + ((g2296) & (!g2344) & (!g1540) & (!g1577) & (g3634) & (g3635)) + ((g2296) & (!g2344) & (!g1540) & (g1577) & (!g3634) & (!g3635)) + ((g2296) & (!g2344) & (g1540) & (!g1577) & (!g3634) & (!g3635)) + ((g2296) & (!g2344) & (g1540) & (!g1577) & (!g3634) & (g3635)) + ((g2296) & (!g2344) & (g1540) & (!g1577) & (g3634) & (!g3635)) + ((g2296) & (!g2344) & (g1540) & (!g1577) & (g3634) & (g3635)) + ((g2296) & (g2344) & (!g1540) & (!g1577) & (!g3634) & (!g3635)));
	assign g3637 = (((!g2377) & (g1610) & (!g3636)) + ((g2377) & (!g1610) & (!g3636)) + ((g2377) & (g1610) & (!g3636)) + ((g2377) & (g1610) & (g3636)));
	assign g3638 = (((!g1900) & (!g2028) & (g2074) & (!g1904) & (!g2043) & (g2080)) + ((!g1900) & (!g2028) & (g2074) & (!g1904) & (g2043) & (g2080)) + ((!g1900) & (!g2028) & (g2074) & (g1904) & (!g2043) & (g2080)) + ((!g1900) & (!g2028) & (g2074) & (g1904) & (g2043) & (g2080)) + ((!g1900) & (g2028) & (!g2074) & (!g1904) & (g2043) & (g2080)) + ((!g1900) & (g2028) & (!g2074) & (g1904) & (g2043) & (g2080)) + ((!g1900) & (g2028) & (g2074) & (!g1904) & (!g2043) & (g2080)) + ((!g1900) & (g2028) & (g2074) & (!g1904) & (g2043) & (!g2080)) + ((!g1900) & (g2028) & (g2074) & (!g1904) & (g2043) & (g2080)) + ((!g1900) & (g2028) & (g2074) & (g1904) & (!g2043) & (g2080)) + ((!g1900) & (g2028) & (g2074) & (g1904) & (g2043) & (!g2080)) + ((!g1900) & (g2028) & (g2074) & (g1904) & (g2043) & (g2080)) + ((g1900) & (!g2028) & (!g2074) & (g1904) & (g2043) & (g2080)) + ((g1900) & (!g2028) & (g2074) & (!g1904) & (!g2043) & (g2080)) + ((g1900) & (!g2028) & (g2074) & (!g1904) & (g2043) & (g2080)) + ((g1900) & (!g2028) & (g2074) & (g1904) & (!g2043) & (g2080)) + ((g1900) & (!g2028) & (g2074) & (g1904) & (g2043) & (!g2080)) + ((g1900) & (!g2028) & (g2074) & (g1904) & (g2043) & (g2080)) + ((g1900) & (g2028) & (!g2074) & (!g1904) & (g2043) & (g2080)) + ((g1900) & (g2028) & (!g2074) & (g1904) & (!g2043) & (g2080)) + ((g1900) & (g2028) & (!g2074) & (g1904) & (g2043) & (g2080)) + ((g1900) & (g2028) & (g2074) & (!g1904) & (!g2043) & (g2080)) + ((g1900) & (g2028) & (g2074) & (!g1904) & (g2043) & (!g2080)) + ((g1900) & (g2028) & (g2074) & (!g1904) & (g2043) & (g2080)) + ((g1900) & (g2028) & (g2074) & (g1904) & (!g2043) & (!g2080)) + ((g1900) & (g2028) & (g2074) & (g1904) & (!g2043) & (g2080)) + ((g1900) & (g2028) & (g2074) & (g1904) & (g2043) & (!g2080)) + ((g1900) & (g2028) & (g2074) & (g1904) & (g2043) & (g2080)));
	assign g3639 = (((!g2190) & (g2205)) + ((g2190) & (!g2205)));
	assign g3640 = (((!g2110) & (!g2156) & (g2125) & (g2162) & (g3638) & (g3639)) + ((!g2110) & (g2156) & (!g2125) & (g2162) & (!g3638) & (g3639)) + ((!g2110) & (g2156) & (!g2125) & (g2162) & (g3638) & (g3639)) + ((!g2110) & (g2156) & (g2125) & (!g2162) & (g3638) & (g3639)) + ((!g2110) & (g2156) & (g2125) & (g2162) & (!g3638) & (g3639)) + ((!g2110) & (g2156) & (g2125) & (g2162) & (g3638) & (g3639)) + ((g2110) & (!g2156) & (!g2125) & (g2162) & (g3638) & (g3639)) + ((g2110) & (!g2156) & (g2125) & (g2162) & (!g3638) & (g3639)) + ((g2110) & (!g2156) & (g2125) & (g2162) & (g3638) & (g3639)) + ((g2110) & (g2156) & (!g2125) & (!g2162) & (g3638) & (g3639)) + ((g2110) & (g2156) & (!g2125) & (g2162) & (!g3638) & (g3639)) + ((g2110) & (g2156) & (!g2125) & (g2162) & (g3638) & (g3639)) + ((g2110) & (g2156) & (g2125) & (!g2162) & (!g3638) & (g3639)) + ((g2110) & (g2156) & (g2125) & (!g2162) & (g3638) & (g3639)) + ((g2110) & (g2156) & (g2125) & (g2162) & (!g3638) & (g3639)) + ((g2110) & (g2156) & (g2125) & (g2162) & (g3638) & (g3639)));
	assign g3641 = (((g2190) & (g2205)));
	assign g3642 = (((!g2236) & (!g2273) & (!g2242) & (!g2288) & (!g3640) & (!g3641)) + ((!g2236) & (!g2273) & (!g2242) & (!g2288) & (!g3640) & (g3641)) + ((!g2236) & (!g2273) & (!g2242) & (!g2288) & (g3640) & (!g3641)) + ((!g2236) & (!g2273) & (!g2242) & (!g2288) & (g3640) & (g3641)) + ((!g2236) & (!g2273) & (!g2242) & (g2288) & (!g3640) & (!g3641)) + ((!g2236) & (!g2273) & (!g2242) & (g2288) & (!g3640) & (g3641)) + ((!g2236) & (!g2273) & (!g2242) & (g2288) & (g3640) & (!g3641)) + ((!g2236) & (!g2273) & (!g2242) & (g2288) & (g3640) & (g3641)) + ((!g2236) & (!g2273) & (g2242) & (!g2288) & (!g3640) & (!g3641)) + ((!g2236) & (!g2273) & (g2242) & (!g2288) & (!g3640) & (g3641)) + ((!g2236) & (!g2273) & (g2242) & (!g2288) & (g3640) & (!g3641)) + ((!g2236) & (!g2273) & (g2242) & (!g2288) & (g3640) & (g3641)) + ((!g2236) & (!g2273) & (g2242) & (g2288) & (!g3640) & (!g3641)) + ((!g2236) & (g2273) & (!g2242) & (!g2288) & (!g3640) & (!g3641)) + ((!g2236) & (g2273) & (!g2242) & (!g2288) & (!g3640) & (g3641)) + ((!g2236) & (g2273) & (!g2242) & (!g2288) & (g3640) & (!g3641)) + ((!g2236) & (g2273) & (!g2242) & (!g2288) & (g3640) & (g3641)) + ((!g2236) & (g2273) & (g2242) & (!g2288) & (!g3640) & (!g3641)) + ((g2236) & (!g2273) & (!g2242) & (!g2288) & (!g3640) & (!g3641)) + ((g2236) & (!g2273) & (!g2242) & (!g2288) & (!g3640) & (g3641)) + ((g2236) & (!g2273) & (!g2242) & (!g2288) & (g3640) & (!g3641)) + ((g2236) & (!g2273) & (!g2242) & (!g2288) & (g3640) & (g3641)) + ((g2236) & (!g2273) & (!g2242) & (g2288) & (!g3640) & (!g3641)) + ((g2236) & (!g2273) & (g2242) & (!g2288) & (!g3640) & (!g3641)) + ((g2236) & (!g2273) & (g2242) & (!g2288) & (!g3640) & (g3641)) + ((g2236) & (!g2273) & (g2242) & (!g2288) & (g3640) & (!g3641)) + ((g2236) & (!g2273) & (g2242) & (!g2288) & (g3640) & (g3641)) + ((g2236) & (g2273) & (!g2242) & (!g2288) & (!g3640) & (!g3641)));
	assign g3643 = (((!g2402) & (g2408)) + ((g2402) & (!g2408)));
	assign g3644 = (((!g2323) & (!g2356) & (g2329) & (g2371) & (!g3642) & (g3643)) + ((!g2323) & (g2356) & (!g2329) & (g2371) & (!g3642) & (g3643)) + ((!g2323) & (g2356) & (!g2329) & (g2371) & (g3642) & (g3643)) + ((!g2323) & (g2356) & (g2329) & (!g2371) & (!g3642) & (g3643)) + ((!g2323) & (g2356) & (g2329) & (g2371) & (!g3642) & (g3643)) + ((!g2323) & (g2356) & (g2329) & (g2371) & (g3642) & (g3643)) + ((g2323) & (!g2356) & (!g2329) & (g2371) & (!g3642) & (g3643)) + ((g2323) & (!g2356) & (g2329) & (g2371) & (!g3642) & (g3643)) + ((g2323) & (!g2356) & (g2329) & (g2371) & (g3642) & (g3643)) + ((g2323) & (g2356) & (!g2329) & (!g2371) & (!g3642) & (g3643)) + ((g2323) & (g2356) & (!g2329) & (g2371) & (!g3642) & (g3643)) + ((g2323) & (g2356) & (!g2329) & (g2371) & (g3642) & (g3643)) + ((g2323) & (g2356) & (g2329) & (!g2371) & (!g3642) & (g3643)) + ((g2323) & (g2356) & (g2329) & (!g2371) & (g3642) & (g3643)) + ((g2323) & (g2356) & (g2329) & (g2371) & (!g3642) & (g3643)) + ((g2323) & (g2356) & (g2329) & (g2371) & (g3642) & (g3643)));
	assign g3645 = (((g2402) & (g2408)));
	assign g3646 = (((!g2456) & (!g2535) & (!g2503) & (!g2539) & (!g3644) & (!g3645)) + ((!g2456) & (!g2535) & (!g2503) & (!g2539) & (!g3644) & (g3645)) + ((!g2456) & (!g2535) & (!g2503) & (!g2539) & (g3644) & (!g3645)) + ((!g2456) & (!g2535) & (!g2503) & (!g2539) & (g3644) & (g3645)) + ((!g2456) & (!g2535) & (!g2503) & (g2539) & (!g3644) & (!g3645)) + ((!g2456) & (!g2535) & (!g2503) & (g2539) & (!g3644) & (g3645)) + ((!g2456) & (!g2535) & (!g2503) & (g2539) & (g3644) & (!g3645)) + ((!g2456) & (!g2535) & (!g2503) & (g2539) & (g3644) & (g3645)) + ((!g2456) & (!g2535) & (g2503) & (!g2539) & (!g3644) & (!g3645)) + ((!g2456) & (!g2535) & (g2503) & (!g2539) & (!g3644) & (g3645)) + ((!g2456) & (!g2535) & (g2503) & (!g2539) & (g3644) & (!g3645)) + ((!g2456) & (!g2535) & (g2503) & (!g2539) & (g3644) & (g3645)) + ((!g2456) & (!g2535) & (g2503) & (g2539) & (!g3644) & (!g3645)) + ((!g2456) & (g2535) & (!g2503) & (!g2539) & (!g3644) & (!g3645)) + ((!g2456) & (g2535) & (!g2503) & (!g2539) & (!g3644) & (g3645)) + ((!g2456) & (g2535) & (!g2503) & (!g2539) & (g3644) & (!g3645)) + ((!g2456) & (g2535) & (!g2503) & (!g2539) & (g3644) & (g3645)) + ((!g2456) & (g2535) & (g2503) & (!g2539) & (!g3644) & (!g3645)) + ((g2456) & (!g2535) & (!g2503) & (!g2539) & (!g3644) & (!g3645)) + ((g2456) & (!g2535) & (!g2503) & (!g2539) & (!g3644) & (g3645)) + ((g2456) & (!g2535) & (!g2503) & (!g2539) & (g3644) & (!g3645)) + ((g2456) & (!g2535) & (!g2503) & (!g2539) & (g3644) & (g3645)) + ((g2456) & (!g2535) & (!g2503) & (g2539) & (!g3644) & (!g3645)) + ((g2456) & (!g2535) & (g2503) & (!g2539) & (!g3644) & (!g3645)) + ((g2456) & (!g2535) & (g2503) & (!g2539) & (!g3644) & (g3645)) + ((g2456) & (!g2535) & (g2503) & (!g2539) & (g3644) & (!g3645)) + ((g2456) & (!g2535) & (g2503) & (!g2539) & (g3644) & (g3645)) + ((g2456) & (g2535) & (!g2503) & (!g2539) & (!g3644) & (!g3645)));
	assign g3647 = (((!g2674) & (g2659)) + ((g2674) & (!g2659)));
	assign g3648 = (((!g2569) & (!g2626) & (g2592) & (g2632) & (!g3646) & (g3647)) + ((!g2569) & (g2626) & (!g2592) & (g2632) & (!g3646) & (g3647)) + ((!g2569) & (g2626) & (!g2592) & (g2632) & (g3646) & (g3647)) + ((!g2569) & (g2626) & (g2592) & (!g2632) & (!g3646) & (g3647)) + ((!g2569) & (g2626) & (g2592) & (g2632) & (!g3646) & (g3647)) + ((!g2569) & (g2626) & (g2592) & (g2632) & (g3646) & (g3647)) + ((g2569) & (!g2626) & (!g2592) & (g2632) & (!g3646) & (g3647)) + ((g2569) & (!g2626) & (g2592) & (g2632) & (!g3646) & (g3647)) + ((g2569) & (!g2626) & (g2592) & (g2632) & (g3646) & (g3647)) + ((g2569) & (g2626) & (!g2592) & (!g2632) & (!g3646) & (g3647)) + ((g2569) & (g2626) & (!g2592) & (g2632) & (!g3646) & (g3647)) + ((g2569) & (g2626) & (!g2592) & (g2632) & (g3646) & (g3647)) + ((g2569) & (g2626) & (g2592) & (!g2632) & (!g3646) & (g3647)) + ((g2569) & (g2626) & (g2592) & (!g2632) & (g3646) & (g3647)) + ((g2569) & (g2626) & (g2592) & (g2632) & (!g3646) & (g3647)) + ((g2569) & (g2626) & (g2592) & (g2632) & (g3646) & (g3647)));
	assign g3649 = (((g2674) & (g2659)));
	assign g3650 = (((!g2733) & (!g2785) & (!g3648) & (!g3649) & (!g2723) & (!g2770)) + ((!g2733) & (!g2785) & (!g3648) & (!g3649) & (!g2723) & (g2770)) + ((!g2733) & (!g2785) & (!g3648) & (!g3649) & (g2723) & (!g2770)) + ((!g2733) & (!g2785) & (!g3648) & (!g3649) & (g2723) & (g2770)) + ((!g2733) & (!g2785) & (!g3648) & (g3649) & (!g2723) & (!g2770)) + ((!g2733) & (!g2785) & (!g3648) & (g3649) & (!g2723) & (g2770)) + ((!g2733) & (!g2785) & (!g3648) & (g3649) & (g2723) & (!g2770)) + ((!g2733) & (!g2785) & (g3648) & (!g3649) & (!g2723) & (!g2770)) + ((!g2733) & (!g2785) & (g3648) & (!g3649) & (!g2723) & (g2770)) + ((!g2733) & (!g2785) & (g3648) & (!g3649) & (g2723) & (!g2770)) + ((!g2733) & (!g2785) & (g3648) & (g3649) & (!g2723) & (!g2770)) + ((!g2733) & (!g2785) & (g3648) & (g3649) & (!g2723) & (g2770)) + ((!g2733) & (!g2785) & (g3648) & (g3649) & (g2723) & (!g2770)) + ((!g2733) & (g2785) & (!g3648) & (!g3649) & (!g2723) & (!g2770)) + ((!g2733) & (g2785) & (!g3648) & (!g3649) & (g2723) & (!g2770)) + ((!g2733) & (g2785) & (!g3648) & (g3649) & (!g2723) & (!g2770)) + ((!g2733) & (g2785) & (g3648) & (!g3649) & (!g2723) & (!g2770)) + ((!g2733) & (g2785) & (g3648) & (g3649) & (!g2723) & (!g2770)) + ((g2733) & (!g2785) & (!g3648) & (!g3649) & (!g2723) & (!g2770)) + ((g2733) & (!g2785) & (!g3648) & (!g3649) & (!g2723) & (g2770)) + ((g2733) & (!g2785) & (!g3648) & (!g3649) & (g2723) & (!g2770)) + ((g2733) & (!g2785) & (!g3648) & (g3649) & (!g2723) & (!g2770)) + ((g2733) & (!g2785) & (!g3648) & (g3649) & (g2723) & (!g2770)) + ((g2733) & (!g2785) & (g3648) & (!g3649) & (!g2723) & (!g2770)) + ((g2733) & (!g2785) & (g3648) & (!g3649) & (g2723) & (!g2770)) + ((g2733) & (!g2785) & (g3648) & (g3649) & (!g2723) & (!g2770)) + ((g2733) & (!g2785) & (g3648) & (g3649) & (g2723) & (!g2770)) + ((g2733) & (g2785) & (!g3648) & (!g3649) & (!g2723) & (!g2770)));
	assign g3651 = (((!g2822) & (!g3650) & (g2816)) + ((g2822) & (!g3650) & (!g2816)) + ((g2822) & (!g3650) & (g2816)) + ((g2822) & (g3650) & (g2816)));
	assign g3652 = (((!g2871) & (!g3651) & (g2848)) + ((!g2871) & (g3651) & (!g2848)) + ((g2871) & (!g3651) & (!g2848)) + ((g2871) & (g3651) & (g2848)));
	assign g3653 = (((!g830) & (!g1898) & (!g7018) & (key[0])) + ((!g830) & (!g1898) & (g7018) & (key[0])) + ((!g830) & (g1898) & (!g7018) & (key[0])) + ((!g830) & (g1898) & (g7018) & (key[0])) + ((g830) & (!g1898) & (g7018) & (!key[0])) + ((g830) & (!g1898) & (g7018) & (key[0])) + ((g830) & (g1898) & (!g7018) & (!key[0])) + ((g830) & (g1898) & (!g7018) & (key[0])));
	assign g3654 = (((!g1884) & (!g1977) & (g1979) & (!g1908) & (!g2030) & (g2085)) + ((!g1884) & (!g1977) & (g1979) & (!g1908) & (g2030) & (g2085)) + ((!g1884) & (!g1977) & (g1979) & (g1908) & (!g2030) & (g2085)) + ((!g1884) & (!g1977) & (g1979) & (g1908) & (g2030) & (g2085)) + ((!g1884) & (g1977) & (!g1979) & (!g1908) & (g2030) & (g2085)) + ((!g1884) & (g1977) & (!g1979) & (g1908) & (g2030) & (g2085)) + ((!g1884) & (g1977) & (g1979) & (!g1908) & (!g2030) & (g2085)) + ((!g1884) & (g1977) & (g1979) & (!g1908) & (g2030) & (!g2085)) + ((!g1884) & (g1977) & (g1979) & (!g1908) & (g2030) & (g2085)) + ((!g1884) & (g1977) & (g1979) & (g1908) & (!g2030) & (g2085)) + ((!g1884) & (g1977) & (g1979) & (g1908) & (g2030) & (!g2085)) + ((!g1884) & (g1977) & (g1979) & (g1908) & (g2030) & (g2085)) + ((g1884) & (!g1977) & (!g1979) & (g1908) & (g2030) & (g2085)) + ((g1884) & (!g1977) & (g1979) & (!g1908) & (!g2030) & (g2085)) + ((g1884) & (!g1977) & (g1979) & (!g1908) & (g2030) & (g2085)) + ((g1884) & (!g1977) & (g1979) & (g1908) & (!g2030) & (g2085)) + ((g1884) & (!g1977) & (g1979) & (g1908) & (g2030) & (!g2085)) + ((g1884) & (!g1977) & (g1979) & (g1908) & (g2030) & (g2085)) + ((g1884) & (g1977) & (!g1979) & (!g1908) & (g2030) & (g2085)) + ((g1884) & (g1977) & (!g1979) & (g1908) & (!g2030) & (g2085)) + ((g1884) & (g1977) & (!g1979) & (g1908) & (g2030) & (g2085)) + ((g1884) & (g1977) & (g1979) & (!g1908) & (!g2030) & (g2085)) + ((g1884) & (g1977) & (g1979) & (!g1908) & (g2030) & (!g2085)) + ((g1884) & (g1977) & (g1979) & (!g1908) & (g2030) & (g2085)) + ((g1884) & (g1977) & (g1979) & (g1908) & (!g2030) & (!g2085)) + ((g1884) & (g1977) & (g1979) & (g1908) & (!g2030) & (g2085)) + ((g1884) & (g1977) & (g1979) & (g1908) & (g2030) & (!g2085)) + ((g1884) & (g1977) & (g1979) & (g1908) & (g2030) & (g2085)));
	assign g3655 = (((!g1986) & (g2192)) + ((g1986) & (!g2192)));
	assign g3656 = (((!g1982) & (!g1984) & (g2112) & (g2167) & (g3654) & (g3655)) + ((!g1982) & (g1984) & (!g2112) & (g2167) & (!g3654) & (g3655)) + ((!g1982) & (g1984) & (!g2112) & (g2167) & (g3654) & (g3655)) + ((!g1982) & (g1984) & (g2112) & (!g2167) & (g3654) & (g3655)) + ((!g1982) & (g1984) & (g2112) & (g2167) & (!g3654) & (g3655)) + ((!g1982) & (g1984) & (g2112) & (g2167) & (g3654) & (g3655)) + ((g1982) & (!g1984) & (!g2112) & (g2167) & (g3654) & (g3655)) + ((g1982) & (!g1984) & (g2112) & (g2167) & (!g3654) & (g3655)) + ((g1982) & (!g1984) & (g2112) & (g2167) & (g3654) & (g3655)) + ((g1982) & (g1984) & (!g2112) & (!g2167) & (g3654) & (g3655)) + ((g1982) & (g1984) & (!g2112) & (g2167) & (!g3654) & (g3655)) + ((g1982) & (g1984) & (!g2112) & (g2167) & (g3654) & (g3655)) + ((g1982) & (g1984) & (g2112) & (!g2167) & (!g3654) & (g3655)) + ((g1982) & (g1984) & (g2112) & (!g2167) & (g3654) & (g3655)) + ((g1982) & (g1984) & (g2112) & (g2167) & (!g3654) & (g3655)) + ((g1982) & (g1984) & (g2112) & (g2167) & (g3654) & (g3655)));
	assign g3657 = (((g1986) & (g2192)));
	assign g3658 = (((!g1991) & (!g1993) & (!g2247) & (!g2275) & (!g3656) & (!g3657)) + ((!g1991) & (!g1993) & (!g2247) & (!g2275) & (!g3656) & (g3657)) + ((!g1991) & (!g1993) & (!g2247) & (!g2275) & (g3656) & (!g3657)) + ((!g1991) & (!g1993) & (!g2247) & (!g2275) & (g3656) & (g3657)) + ((!g1991) & (!g1993) & (!g2247) & (g2275) & (!g3656) & (!g3657)) + ((!g1991) & (!g1993) & (!g2247) & (g2275) & (!g3656) & (g3657)) + ((!g1991) & (!g1993) & (!g2247) & (g2275) & (g3656) & (!g3657)) + ((!g1991) & (!g1993) & (!g2247) & (g2275) & (g3656) & (g3657)) + ((!g1991) & (!g1993) & (g2247) & (!g2275) & (!g3656) & (!g3657)) + ((!g1991) & (!g1993) & (g2247) & (!g2275) & (!g3656) & (g3657)) + ((!g1991) & (!g1993) & (g2247) & (!g2275) & (g3656) & (!g3657)) + ((!g1991) & (!g1993) & (g2247) & (!g2275) & (g3656) & (g3657)) + ((!g1991) & (!g1993) & (g2247) & (g2275) & (!g3656) & (!g3657)) + ((!g1991) & (g1993) & (!g2247) & (!g2275) & (!g3656) & (!g3657)) + ((!g1991) & (g1993) & (!g2247) & (!g2275) & (!g3656) & (g3657)) + ((!g1991) & (g1993) & (!g2247) & (!g2275) & (g3656) & (!g3657)) + ((!g1991) & (g1993) & (!g2247) & (!g2275) & (g3656) & (g3657)) + ((!g1991) & (g1993) & (g2247) & (!g2275) & (!g3656) & (!g3657)) + ((g1991) & (!g1993) & (!g2247) & (!g2275) & (!g3656) & (!g3657)) + ((g1991) & (!g1993) & (!g2247) & (!g2275) & (!g3656) & (g3657)) + ((g1991) & (!g1993) & (!g2247) & (!g2275) & (g3656) & (!g3657)) + ((g1991) & (!g1993) & (!g2247) & (!g2275) & (g3656) & (g3657)) + ((g1991) & (!g1993) & (!g2247) & (g2275) & (!g3656) & (!g3657)) + ((g1991) & (!g1993) & (g2247) & (!g2275) & (!g3656) & (!g3657)) + ((g1991) & (!g1993) & (g2247) & (!g2275) & (!g3656) & (g3657)) + ((g1991) & (!g1993) & (g2247) & (!g2275) & (g3656) & (!g3657)) + ((g1991) & (!g1993) & (g2247) & (!g2275) & (g3656) & (g3657)) + ((g1991) & (g1993) & (!g2247) & (!g2275) & (!g3656) & (!g3657)));
	assign g3659 = (((!g2001) & (g2413)) + ((g2001) & (!g2413)));
	assign g3660 = (((!g1996) & (!g1998) & (g2334) & (g2358) & (!g3658) & (g3659)) + ((!g1996) & (g1998) & (!g2334) & (g2358) & (!g3658) & (g3659)) + ((!g1996) & (g1998) & (!g2334) & (g2358) & (g3658) & (g3659)) + ((!g1996) & (g1998) & (g2334) & (!g2358) & (!g3658) & (g3659)) + ((!g1996) & (g1998) & (g2334) & (g2358) & (!g3658) & (g3659)) + ((!g1996) & (g1998) & (g2334) & (g2358) & (g3658) & (g3659)) + ((g1996) & (!g1998) & (!g2334) & (g2358) & (!g3658) & (g3659)) + ((g1996) & (!g1998) & (g2334) & (g2358) & (!g3658) & (g3659)) + ((g1996) & (!g1998) & (g2334) & (g2358) & (g3658) & (g3659)) + ((g1996) & (g1998) & (!g2334) & (!g2358) & (!g3658) & (g3659)) + ((g1996) & (g1998) & (!g2334) & (g2358) & (!g3658) & (g3659)) + ((g1996) & (g1998) & (!g2334) & (g2358) & (g3658) & (g3659)) + ((g1996) & (g1998) & (g2334) & (!g2358) & (!g3658) & (g3659)) + ((g1996) & (g1998) & (g2334) & (!g2358) & (g3658) & (g3659)) + ((g1996) & (g1998) & (g2334) & (g2358) & (!g3658) & (g3659)) + ((g1996) & (g1998) & (g2334) & (g2358) & (g3658) & (g3659)));
	assign g3661 = (((g2001) & (g2413)));
	assign g3662 = (((!g2003) & (!g2005) & (!g2462) & (!g2542) & (!g3660) & (!g3661)) + ((!g2003) & (!g2005) & (!g2462) & (!g2542) & (!g3660) & (g3661)) + ((!g2003) & (!g2005) & (!g2462) & (!g2542) & (g3660) & (!g3661)) + ((!g2003) & (!g2005) & (!g2462) & (!g2542) & (g3660) & (g3661)) + ((!g2003) & (!g2005) & (!g2462) & (g2542) & (!g3660) & (!g3661)) + ((!g2003) & (!g2005) & (!g2462) & (g2542) & (!g3660) & (g3661)) + ((!g2003) & (!g2005) & (!g2462) & (g2542) & (g3660) & (!g3661)) + ((!g2003) & (!g2005) & (!g2462) & (g2542) & (g3660) & (g3661)) + ((!g2003) & (!g2005) & (g2462) & (!g2542) & (!g3660) & (!g3661)) + ((!g2003) & (!g2005) & (g2462) & (!g2542) & (!g3660) & (g3661)) + ((!g2003) & (!g2005) & (g2462) & (!g2542) & (g3660) & (!g3661)) + ((!g2003) & (!g2005) & (g2462) & (!g2542) & (g3660) & (g3661)) + ((!g2003) & (!g2005) & (g2462) & (g2542) & (!g3660) & (!g3661)) + ((!g2003) & (g2005) & (!g2462) & (!g2542) & (!g3660) & (!g3661)) + ((!g2003) & (g2005) & (!g2462) & (!g2542) & (!g3660) & (g3661)) + ((!g2003) & (g2005) & (!g2462) & (!g2542) & (g3660) & (!g3661)) + ((!g2003) & (g2005) & (!g2462) & (!g2542) & (g3660) & (g3661)) + ((!g2003) & (g2005) & (g2462) & (!g2542) & (!g3660) & (!g3661)) + ((g2003) & (!g2005) & (!g2462) & (!g2542) & (!g3660) & (!g3661)) + ((g2003) & (!g2005) & (!g2462) & (!g2542) & (!g3660) & (g3661)) + ((g2003) & (!g2005) & (!g2462) & (!g2542) & (g3660) & (!g3661)) + ((g2003) & (!g2005) & (!g2462) & (!g2542) & (g3660) & (g3661)) + ((g2003) & (!g2005) & (!g2462) & (g2542) & (!g3660) & (!g3661)) + ((g2003) & (!g2005) & (g2462) & (!g2542) & (!g3660) & (!g3661)) + ((g2003) & (!g2005) & (g2462) & (!g2542) & (!g3660) & (g3661)) + ((g2003) & (!g2005) & (g2462) & (!g2542) & (g3660) & (!g3661)) + ((g2003) & (!g2005) & (g2462) & (!g2542) & (g3660) & (g3661)) + ((g2003) & (g2005) & (!g2462) & (!g2542) & (!g3660) & (!g3661)));
	assign g3663 = (((!g2051) & (g2661)) + ((g2051) & (!g2661)));
	assign g3664 = (((!g2011) & (!g2013) & (g2572) & (g2637) & (!g3662) & (g3663)) + ((!g2011) & (g2013) & (!g2572) & (g2637) & (!g3662) & (g3663)) + ((!g2011) & (g2013) & (!g2572) & (g2637) & (g3662) & (g3663)) + ((!g2011) & (g2013) & (g2572) & (!g2637) & (!g3662) & (g3663)) + ((!g2011) & (g2013) & (g2572) & (g2637) & (!g3662) & (g3663)) + ((!g2011) & (g2013) & (g2572) & (g2637) & (g3662) & (g3663)) + ((g2011) & (!g2013) & (!g2572) & (g2637) & (!g3662) & (g3663)) + ((g2011) & (!g2013) & (g2572) & (g2637) & (!g3662) & (g3663)) + ((g2011) & (!g2013) & (g2572) & (g2637) & (g3662) & (g3663)) + ((g2011) & (g2013) & (!g2572) & (!g2637) & (!g3662) & (g3663)) + ((g2011) & (g2013) & (!g2572) & (g2637) & (!g3662) & (g3663)) + ((g2011) & (g2013) & (!g2572) & (g2637) & (g3662) & (g3663)) + ((g2011) & (g2013) & (g2572) & (!g2637) & (!g3662) & (g3663)) + ((g2011) & (g2013) & (g2572) & (!g2637) & (g3662) & (g3663)) + ((g2011) & (g2013) & (g2572) & (g2637) & (!g3662) & (g3663)) + ((g2011) & (g2013) & (g2572) & (g2637) & (g3662) & (g3663)));
	assign g3665 = (((g2051) & (g2661)));
	assign g3666 = (((!g2100) & (!g2133) & (!g2742) & (!g2772) & (!g3664) & (!g3665)) + ((!g2100) & (!g2133) & (!g2742) & (!g2772) & (!g3664) & (g3665)) + ((!g2100) & (!g2133) & (!g2742) & (!g2772) & (g3664) & (!g3665)) + ((!g2100) & (!g2133) & (!g2742) & (!g2772) & (g3664) & (g3665)) + ((!g2100) & (!g2133) & (!g2742) & (g2772) & (!g3664) & (!g3665)) + ((!g2100) & (!g2133) & (!g2742) & (g2772) & (!g3664) & (g3665)) + ((!g2100) & (!g2133) & (!g2742) & (g2772) & (g3664) & (!g3665)) + ((!g2100) & (!g2133) & (!g2742) & (g2772) & (g3664) & (g3665)) + ((!g2100) & (!g2133) & (g2742) & (!g2772) & (!g3664) & (!g3665)) + ((!g2100) & (!g2133) & (g2742) & (!g2772) & (!g3664) & (g3665)) + ((!g2100) & (!g2133) & (g2742) & (!g2772) & (g3664) & (!g3665)) + ((!g2100) & (!g2133) & (g2742) & (!g2772) & (g3664) & (g3665)) + ((!g2100) & (!g2133) & (g2742) & (g2772) & (!g3664) & (!g3665)) + ((!g2100) & (g2133) & (!g2742) & (!g2772) & (!g3664) & (!g3665)) + ((!g2100) & (g2133) & (!g2742) & (!g2772) & (!g3664) & (g3665)) + ((!g2100) & (g2133) & (!g2742) & (!g2772) & (g3664) & (!g3665)) + ((!g2100) & (g2133) & (!g2742) & (!g2772) & (g3664) & (g3665)) + ((!g2100) & (g2133) & (g2742) & (!g2772) & (!g3664) & (!g3665)) + ((g2100) & (!g2133) & (!g2742) & (!g2772) & (!g3664) & (!g3665)) + ((g2100) & (!g2133) & (!g2742) & (!g2772) & (!g3664) & (g3665)) + ((g2100) & (!g2133) & (!g2742) & (!g2772) & (g3664) & (!g3665)) + ((g2100) & (!g2133) & (!g2742) & (!g2772) & (g3664) & (g3665)) + ((g2100) & (!g2133) & (!g2742) & (g2772) & (!g3664) & (!g3665)) + ((g2100) & (!g2133) & (g2742) & (!g2772) & (!g3664) & (!g3665)) + ((g2100) & (!g2133) & (g2742) & (!g2772) & (!g3664) & (g3665)) + ((g2100) & (!g2133) & (g2742) & (!g2772) & (g3664) & (!g3665)) + ((g2100) & (!g2133) & (g2742) & (!g2772) & (g3664) & (g3665)) + ((g2100) & (g2133) & (!g2742) & (!g2772) & (!g3664) & (!g3665)));
	assign g3667 = (((!g2180) & (g2827) & (!g3666)) + ((g2180) & (!g2827) & (!g3666)) + ((g2180) & (g2827) & (!g3666)) + ((g2180) & (g2827) & (g3666)));
	assign g3668 = (((!g2212) & (!g2851) & (g3667)) + ((!g2212) & (g2851) & (!g3667)) + ((g2212) & (!g2851) & (!g3667)) + ((g2212) & (g2851) & (g3667)));
	assign g3669 = (((!g1898) & (!g2022) & (g2071) & (!g1902) & (!g2036) & (g2077)) + ((!g1898) & (!g2022) & (g2071) & (!g1902) & (g2036) & (g2077)) + ((!g1898) & (!g2022) & (g2071) & (g1902) & (!g2036) & (g2077)) + ((!g1898) & (!g2022) & (g2071) & (g1902) & (g2036) & (g2077)) + ((!g1898) & (g2022) & (!g2071) & (!g1902) & (g2036) & (g2077)) + ((!g1898) & (g2022) & (!g2071) & (g1902) & (g2036) & (g2077)) + ((!g1898) & (g2022) & (g2071) & (!g1902) & (!g2036) & (g2077)) + ((!g1898) & (g2022) & (g2071) & (!g1902) & (g2036) & (!g2077)) + ((!g1898) & (g2022) & (g2071) & (!g1902) & (g2036) & (g2077)) + ((!g1898) & (g2022) & (g2071) & (g1902) & (!g2036) & (g2077)) + ((!g1898) & (g2022) & (g2071) & (g1902) & (g2036) & (!g2077)) + ((!g1898) & (g2022) & (g2071) & (g1902) & (g2036) & (g2077)) + ((g1898) & (!g2022) & (!g2071) & (g1902) & (g2036) & (g2077)) + ((g1898) & (!g2022) & (g2071) & (!g1902) & (!g2036) & (g2077)) + ((g1898) & (!g2022) & (g2071) & (!g1902) & (g2036) & (g2077)) + ((g1898) & (!g2022) & (g2071) & (g1902) & (!g2036) & (g2077)) + ((g1898) & (!g2022) & (g2071) & (g1902) & (g2036) & (!g2077)) + ((g1898) & (!g2022) & (g2071) & (g1902) & (g2036) & (g2077)) + ((g1898) & (g2022) & (!g2071) & (!g1902) & (g2036) & (g2077)) + ((g1898) & (g2022) & (!g2071) & (g1902) & (!g2036) & (g2077)) + ((g1898) & (g2022) & (!g2071) & (g1902) & (g2036) & (g2077)) + ((g1898) & (g2022) & (g2071) & (!g1902) & (!g2036) & (g2077)) + ((g1898) & (g2022) & (g2071) & (!g1902) & (g2036) & (!g2077)) + ((g1898) & (g2022) & (g2071) & (!g1902) & (g2036) & (g2077)) + ((g1898) & (g2022) & (g2071) & (g1902) & (!g2036) & (!g2077)) + ((g1898) & (g2022) & (g2071) & (g1902) & (!g2036) & (g2077)) + ((g1898) & (g2022) & (g2071) & (g1902) & (g2036) & (!g2077)) + ((g1898) & (g2022) & (g2071) & (g1902) & (g2036) & (g2077)));
	assign g3670 = (((!g2184) & (g2198)) + ((g2184) & (!g2198)));
	assign g3671 = (((!g2104) & (!g2153) & (g2118) & (g2159) & (g3669) & (g3670)) + ((!g2104) & (g2153) & (!g2118) & (g2159) & (!g3669) & (g3670)) + ((!g2104) & (g2153) & (!g2118) & (g2159) & (g3669) & (g3670)) + ((!g2104) & (g2153) & (g2118) & (!g2159) & (g3669) & (g3670)) + ((!g2104) & (g2153) & (g2118) & (g2159) & (!g3669) & (g3670)) + ((!g2104) & (g2153) & (g2118) & (g2159) & (g3669) & (g3670)) + ((g2104) & (!g2153) & (!g2118) & (g2159) & (g3669) & (g3670)) + ((g2104) & (!g2153) & (g2118) & (g2159) & (!g3669) & (g3670)) + ((g2104) & (!g2153) & (g2118) & (g2159) & (g3669) & (g3670)) + ((g2104) & (g2153) & (!g2118) & (!g2159) & (g3669) & (g3670)) + ((g2104) & (g2153) & (!g2118) & (g2159) & (!g3669) & (g3670)) + ((g2104) & (g2153) & (!g2118) & (g2159) & (g3669) & (g3670)) + ((g2104) & (g2153) & (g2118) & (!g2159) & (!g3669) & (g3670)) + ((g2104) & (g2153) & (g2118) & (!g2159) & (g3669) & (g3670)) + ((g2104) & (g2153) & (g2118) & (g2159) & (!g3669) & (g3670)) + ((g2104) & (g2153) & (g2118) & (g2159) & (g3669) & (g3670)));
	assign g3672 = (((g2184) & (g2198)));
	assign g3673 = (((!g2233) & (!g2267) & (!g2239) & (!g2281) & (!g3671) & (!g3672)) + ((!g2233) & (!g2267) & (!g2239) & (!g2281) & (!g3671) & (g3672)) + ((!g2233) & (!g2267) & (!g2239) & (!g2281) & (g3671) & (!g3672)) + ((!g2233) & (!g2267) & (!g2239) & (!g2281) & (g3671) & (g3672)) + ((!g2233) & (!g2267) & (!g2239) & (g2281) & (!g3671) & (!g3672)) + ((!g2233) & (!g2267) & (!g2239) & (g2281) & (!g3671) & (g3672)) + ((!g2233) & (!g2267) & (!g2239) & (g2281) & (g3671) & (!g3672)) + ((!g2233) & (!g2267) & (!g2239) & (g2281) & (g3671) & (g3672)) + ((!g2233) & (!g2267) & (g2239) & (!g2281) & (!g3671) & (!g3672)) + ((!g2233) & (!g2267) & (g2239) & (!g2281) & (!g3671) & (g3672)) + ((!g2233) & (!g2267) & (g2239) & (!g2281) & (g3671) & (!g3672)) + ((!g2233) & (!g2267) & (g2239) & (!g2281) & (g3671) & (g3672)) + ((!g2233) & (!g2267) & (g2239) & (g2281) & (!g3671) & (!g3672)) + ((!g2233) & (g2267) & (!g2239) & (!g2281) & (!g3671) & (!g3672)) + ((!g2233) & (g2267) & (!g2239) & (!g2281) & (!g3671) & (g3672)) + ((!g2233) & (g2267) & (!g2239) & (!g2281) & (g3671) & (!g3672)) + ((!g2233) & (g2267) & (!g2239) & (!g2281) & (g3671) & (g3672)) + ((!g2233) & (g2267) & (g2239) & (!g2281) & (!g3671) & (!g3672)) + ((g2233) & (!g2267) & (!g2239) & (!g2281) & (!g3671) & (!g3672)) + ((g2233) & (!g2267) & (!g2239) & (!g2281) & (!g3671) & (g3672)) + ((g2233) & (!g2267) & (!g2239) & (!g2281) & (g3671) & (!g3672)) + ((g2233) & (!g2267) & (!g2239) & (!g2281) & (g3671) & (g3672)) + ((g2233) & (!g2267) & (!g2239) & (g2281) & (!g3671) & (!g3672)) + ((g2233) & (!g2267) & (g2239) & (!g2281) & (!g3671) & (!g3672)) + ((g2233) & (!g2267) & (g2239) & (!g2281) & (!g3671) & (g3672)) + ((g2233) & (!g2267) & (g2239) & (!g2281) & (g3671) & (!g3672)) + ((g2233) & (!g2267) & (g2239) & (!g2281) & (g3671) & (g3672)) + ((g2233) & (g2267) & (!g2239) & (!g2281) & (!g3671) & (!g3672)));
	assign g3674 = (((!g2399) & (g2405)) + ((g2399) & (!g2405)));
	assign g3675 = (((!g2320) & (!g2350) & (g2326) & (g2364) & (!g3673) & (g3674)) + ((!g2320) & (g2350) & (!g2326) & (g2364) & (!g3673) & (g3674)) + ((!g2320) & (g2350) & (!g2326) & (g2364) & (g3673) & (g3674)) + ((!g2320) & (g2350) & (g2326) & (!g2364) & (!g3673) & (g3674)) + ((!g2320) & (g2350) & (g2326) & (g2364) & (!g3673) & (g3674)) + ((!g2320) & (g2350) & (g2326) & (g2364) & (g3673) & (g3674)) + ((g2320) & (!g2350) & (!g2326) & (g2364) & (!g3673) & (g3674)) + ((g2320) & (!g2350) & (g2326) & (g2364) & (!g3673) & (g3674)) + ((g2320) & (!g2350) & (g2326) & (g2364) & (g3673) & (g3674)) + ((g2320) & (g2350) & (!g2326) & (!g2364) & (!g3673) & (g3674)) + ((g2320) & (g2350) & (!g2326) & (g2364) & (!g3673) & (g3674)) + ((g2320) & (g2350) & (!g2326) & (g2364) & (g3673) & (g3674)) + ((g2320) & (g2350) & (g2326) & (!g2364) & (!g3673) & (g3674)) + ((g2320) & (g2350) & (g2326) & (!g2364) & (g3673) & (g3674)) + ((g2320) & (g2350) & (g2326) & (g2364) & (!g3673) & (g3674)) + ((g2320) & (g2350) & (g2326) & (g2364) & (g3673) & (g3674)));
	assign g3676 = (((g2399) & (g2405)));
	assign g3677 = (((!g2434) & (!g2533) & (!g2480) & (!g2537) & (!g3675) & (!g3676)) + ((!g2434) & (!g2533) & (!g2480) & (!g2537) & (!g3675) & (g3676)) + ((!g2434) & (!g2533) & (!g2480) & (!g2537) & (g3675) & (!g3676)) + ((!g2434) & (!g2533) & (!g2480) & (!g2537) & (g3675) & (g3676)) + ((!g2434) & (!g2533) & (!g2480) & (g2537) & (!g3675) & (!g3676)) + ((!g2434) & (!g2533) & (!g2480) & (g2537) & (!g3675) & (g3676)) + ((!g2434) & (!g2533) & (!g2480) & (g2537) & (g3675) & (!g3676)) + ((!g2434) & (!g2533) & (!g2480) & (g2537) & (g3675) & (g3676)) + ((!g2434) & (!g2533) & (g2480) & (!g2537) & (!g3675) & (!g3676)) + ((!g2434) & (!g2533) & (g2480) & (!g2537) & (!g3675) & (g3676)) + ((!g2434) & (!g2533) & (g2480) & (!g2537) & (g3675) & (!g3676)) + ((!g2434) & (!g2533) & (g2480) & (!g2537) & (g3675) & (g3676)) + ((!g2434) & (!g2533) & (g2480) & (g2537) & (!g3675) & (!g3676)) + ((!g2434) & (g2533) & (!g2480) & (!g2537) & (!g3675) & (!g3676)) + ((!g2434) & (g2533) & (!g2480) & (!g2537) & (!g3675) & (g3676)) + ((!g2434) & (g2533) & (!g2480) & (!g2537) & (g3675) & (!g3676)) + ((!g2434) & (g2533) & (!g2480) & (!g2537) & (g3675) & (g3676)) + ((!g2434) & (g2533) & (g2480) & (!g2537) & (!g3675) & (!g3676)) + ((g2434) & (!g2533) & (!g2480) & (!g2537) & (!g3675) & (!g3676)) + ((g2434) & (!g2533) & (!g2480) & (!g2537) & (!g3675) & (g3676)) + ((g2434) & (!g2533) & (!g2480) & (!g2537) & (g3675) & (!g3676)) + ((g2434) & (!g2533) & (!g2480) & (!g2537) & (g3675) & (g3676)) + ((g2434) & (!g2533) & (!g2480) & (g2537) & (!g3675) & (!g3676)) + ((g2434) & (!g2533) & (g2480) & (!g2537) & (!g3675) & (!g3676)) + ((g2434) & (!g2533) & (g2480) & (!g2537) & (!g3675) & (g3676)) + ((g2434) & (!g2533) & (g2480) & (!g2537) & (g3675) & (!g3676)) + ((g2434) & (!g2533) & (g2480) & (!g2537) & (g3675) & (g3676)) + ((g2434) & (g2533) & (!g2480) & (!g2537) & (!g3675) & (!g3676)));
	assign g3678 = (((!g2434) & (!g2480) & (!g3675) & (!g3676) & (!g5806) & (g5807)) + ((!g2434) & (!g2480) & (!g3675) & (g3676) & (!g5806) & (g5807)) + ((!g2434) & (!g2480) & (g3675) & (!g3676) & (!g5806) & (g5807)) + ((!g2434) & (!g2480) & (g3675) & (g3676) & (!g5806) & (g5807)) + ((!g2434) & (g2480) & (!g3675) & (!g3676) & (!g5806) & (g5807)) + ((!g2434) & (g2480) & (!g3675) & (g3676) & (!g5806) & (g5807)) + ((!g2434) & (g2480) & (!g3675) & (g3676) & (g5806) & (g5807)) + ((!g2434) & (g2480) & (g3675) & (!g3676) & (!g5806) & (g5807)) + ((!g2434) & (g2480) & (g3675) & (!g3676) & (g5806) & (g5807)) + ((!g2434) & (g2480) & (g3675) & (g3676) & (!g5806) & (g5807)) + ((!g2434) & (g2480) & (g3675) & (g3676) & (g5806) & (g5807)) + ((g2434) & (!g2480) & (!g3675) & (!g3676) & (!g5806) & (g5807)) + ((g2434) & (!g2480) & (!g3675) & (g3676) & (!g5806) & (g5807)) + ((g2434) & (!g2480) & (!g3675) & (g3676) & (g5806) & (g5807)) + ((g2434) & (!g2480) & (g3675) & (!g3676) & (!g5806) & (g5807)) + ((g2434) & (!g2480) & (g3675) & (!g3676) & (g5806) & (g5807)) + ((g2434) & (!g2480) & (g3675) & (g3676) & (!g5806) & (g5807)) + ((g2434) & (!g2480) & (g3675) & (g3676) & (g5806) & (g5807)) + ((g2434) & (g2480) & (!g3675) & (!g3676) & (!g5806) & (g5807)) + ((g2434) & (g2480) & (!g3675) & (!g3676) & (g5806) & (g5807)) + ((g2434) & (g2480) & (!g3675) & (g3676) & (!g5806) & (g5807)) + ((g2434) & (g2480) & (!g3675) & (g3676) & (g5806) & (g5807)) + ((g2434) & (g2480) & (g3675) & (!g3676) & (!g5806) & (g5807)) + ((g2434) & (g2480) & (g3675) & (!g3676) & (g5806) & (g5807)) + ((g2434) & (g2480) & (g3675) & (g3676) & (!g5806) & (g5807)) + ((g2434) & (g2480) & (g3675) & (g3676) & (g5806) & (g5807)));
	assign g3679 = (((g2653) & (g2667)));
	assign g3680 = (((!g2718) & (!g2764) & (!g2728) & (!g2778) & (!g3678) & (!g3679)) + ((!g2718) & (!g2764) & (!g2728) & (!g2778) & (!g3678) & (g3679)) + ((!g2718) & (!g2764) & (!g2728) & (!g2778) & (g3678) & (!g3679)) + ((!g2718) & (!g2764) & (!g2728) & (!g2778) & (g3678) & (g3679)) + ((!g2718) & (!g2764) & (!g2728) & (g2778) & (!g3678) & (!g3679)) + ((!g2718) & (!g2764) & (!g2728) & (g2778) & (!g3678) & (g3679)) + ((!g2718) & (!g2764) & (!g2728) & (g2778) & (g3678) & (!g3679)) + ((!g2718) & (!g2764) & (!g2728) & (g2778) & (g3678) & (g3679)) + ((!g2718) & (!g2764) & (g2728) & (!g2778) & (!g3678) & (!g3679)) + ((!g2718) & (!g2764) & (g2728) & (!g2778) & (!g3678) & (g3679)) + ((!g2718) & (!g2764) & (g2728) & (!g2778) & (g3678) & (!g3679)) + ((!g2718) & (!g2764) & (g2728) & (!g2778) & (g3678) & (g3679)) + ((!g2718) & (!g2764) & (g2728) & (g2778) & (!g3678) & (!g3679)) + ((!g2718) & (g2764) & (!g2728) & (!g2778) & (!g3678) & (!g3679)) + ((!g2718) & (g2764) & (!g2728) & (!g2778) & (!g3678) & (g3679)) + ((!g2718) & (g2764) & (!g2728) & (!g2778) & (g3678) & (!g3679)) + ((!g2718) & (g2764) & (!g2728) & (!g2778) & (g3678) & (g3679)) + ((!g2718) & (g2764) & (g2728) & (!g2778) & (!g3678) & (!g3679)) + ((g2718) & (!g2764) & (!g2728) & (!g2778) & (!g3678) & (!g3679)) + ((g2718) & (!g2764) & (!g2728) & (!g2778) & (!g3678) & (g3679)) + ((g2718) & (!g2764) & (!g2728) & (!g2778) & (g3678) & (!g3679)) + ((g2718) & (!g2764) & (!g2728) & (!g2778) & (g3678) & (g3679)) + ((g2718) & (!g2764) & (!g2728) & (g2778) & (!g3678) & (!g3679)) + ((g2718) & (!g2764) & (g2728) & (!g2778) & (!g3678) & (!g3679)) + ((g2718) & (!g2764) & (g2728) & (!g2778) & (!g3678) & (g3679)) + ((g2718) & (!g2764) & (g2728) & (!g2778) & (g3678) & (!g3679)) + ((g2718) & (!g2764) & (g2728) & (!g2778) & (g3678) & (g3679)) + ((g2718) & (g2764) & (!g2728) & (!g2778) & (!g3678) & (!g3679)));
	assign g3681 = (((!g2891) & (g2895)) + ((g2891) & (!g2895)));
	assign g3682 = (((!g2813) & (!g2838) & (g2819) & (g2860) & (!g3680) & (g3681)) + ((!g2813) & (g2838) & (!g2819) & (g2860) & (!g3680) & (g3681)) + ((!g2813) & (g2838) & (!g2819) & (g2860) & (g3680) & (g3681)) + ((!g2813) & (g2838) & (g2819) & (!g2860) & (!g3680) & (g3681)) + ((!g2813) & (g2838) & (g2819) & (g2860) & (!g3680) & (g3681)) + ((!g2813) & (g2838) & (g2819) & (g2860) & (g3680) & (g3681)) + ((g2813) & (!g2838) & (!g2819) & (g2860) & (!g3680) & (g3681)) + ((g2813) & (!g2838) & (g2819) & (g2860) & (!g3680) & (g3681)) + ((g2813) & (!g2838) & (g2819) & (g2860) & (g3680) & (g3681)) + ((g2813) & (g2838) & (!g2819) & (!g2860) & (!g3680) & (g3681)) + ((g2813) & (g2838) & (!g2819) & (g2860) & (!g3680) & (g3681)) + ((g2813) & (g2838) & (!g2819) & (g2860) & (g3680) & (g3681)) + ((g2813) & (g2838) & (g2819) & (!g2860) & (!g3680) & (g3681)) + ((g2813) & (g2838) & (g2819) & (!g2860) & (g3680) & (g3681)) + ((g2813) & (g2838) & (g2819) & (g2860) & (!g3680) & (g3681)) + ((g2813) & (g2838) & (g2819) & (g2860) & (g3680) & (g3681)));
	assign g3683 = (((g2891) & (g2895)));
	assign g3684 = (((!g2916) & (!g3009) & (!g2962) & (!g3013) & (!g3682) & (!g3683)) + ((!g2916) & (!g3009) & (!g2962) & (!g3013) & (!g3682) & (g3683)) + ((!g2916) & (!g3009) & (!g2962) & (!g3013) & (g3682) & (!g3683)) + ((!g2916) & (!g3009) & (!g2962) & (!g3013) & (g3682) & (g3683)) + ((!g2916) & (!g3009) & (!g2962) & (g3013) & (!g3682) & (!g3683)) + ((!g2916) & (!g3009) & (!g2962) & (g3013) & (!g3682) & (g3683)) + ((!g2916) & (!g3009) & (!g2962) & (g3013) & (g3682) & (!g3683)) + ((!g2916) & (!g3009) & (!g2962) & (g3013) & (g3682) & (g3683)) + ((!g2916) & (!g3009) & (g2962) & (!g3013) & (!g3682) & (!g3683)) + ((!g2916) & (!g3009) & (g2962) & (!g3013) & (!g3682) & (g3683)) + ((!g2916) & (!g3009) & (g2962) & (!g3013) & (g3682) & (!g3683)) + ((!g2916) & (!g3009) & (g2962) & (!g3013) & (g3682) & (g3683)) + ((!g2916) & (!g3009) & (g2962) & (g3013) & (!g3682) & (!g3683)) + ((!g2916) & (g3009) & (!g2962) & (!g3013) & (!g3682) & (!g3683)) + ((!g2916) & (g3009) & (!g2962) & (!g3013) & (!g3682) & (g3683)) + ((!g2916) & (g3009) & (!g2962) & (!g3013) & (g3682) & (!g3683)) + ((!g2916) & (g3009) & (!g2962) & (!g3013) & (g3682) & (g3683)) + ((!g2916) & (g3009) & (g2962) & (!g3013) & (!g3682) & (!g3683)) + ((g2916) & (!g3009) & (!g2962) & (!g3013) & (!g3682) & (!g3683)) + ((g2916) & (!g3009) & (!g2962) & (!g3013) & (!g3682) & (g3683)) + ((g2916) & (!g3009) & (!g2962) & (!g3013) & (g3682) & (!g3683)) + ((g2916) & (!g3009) & (!g2962) & (!g3013) & (g3682) & (g3683)) + ((g2916) & (!g3009) & (!g2962) & (g3013) & (!g3682) & (!g3683)) + ((g2916) & (!g3009) & (g2962) & (!g3013) & (!g3682) & (!g3683)) + ((g2916) & (!g3009) & (g2962) & (!g3013) & (!g3682) & (g3683)) + ((g2916) & (!g3009) & (g2962) & (!g3013) & (g3682) & (!g3683)) + ((g2916) & (!g3009) & (g2962) & (!g3013) & (g3682) & (g3683)) + ((g2916) & (g3009) & (!g2962) & (!g3013) & (!g3682) & (!g3683)));
	assign g3685 = (((!g3031) & (g3053) & (!g3684)) + ((g3031) & (!g3053) & (!g3684)) + ((g3031) & (g3053) & (!g3684)) + ((g3031) & (g3053) & (g3684)));
	assign g3686 = (((!g3088) & (!g3128) & (!g3685) & (!g3084) & (g3106)) + ((!g3088) & (!g3128) & (!g3685) & (g3084) & (g3106)) + ((!g3088) & (!g3128) & (g3685) & (!g3084) & (g3106)) + ((!g3088) & (!g3128) & (g3685) & (g3084) & (!g3106)) + ((!g3088) & (g3128) & (!g3685) & (!g3084) & (!g3106)) + ((!g3088) & (g3128) & (!g3685) & (g3084) & (!g3106)) + ((!g3088) & (g3128) & (g3685) & (!g3084) & (!g3106)) + ((!g3088) & (g3128) & (g3685) & (g3084) & (g3106)) + ((g3088) & (!g3128) & (!g3685) & (!g3084) & (g3106)) + ((g3088) & (!g3128) & (!g3685) & (g3084) & (!g3106)) + ((g3088) & (!g3128) & (g3685) & (!g3084) & (!g3106)) + ((g3088) & (!g3128) & (g3685) & (g3084) & (!g3106)) + ((g3088) & (g3128) & (!g3685) & (!g3084) & (!g3106)) + ((g3088) & (g3128) & (!g3685) & (g3084) & (g3106)) + ((g3088) & (g3128) & (g3685) & (!g3084) & (g3106)) + ((g3088) & (g3128) & (g3685) & (g3084) & (g3106)));
	assign g8277 = (((!g5560) & (g5569) & (!g3687)) + ((!g5560) & (g5569) & (g3687)) + ((g5560) & (!g5569) & (g3687)) + ((g5560) & (g5569) & (g3687)));
	assign g3688 = (((!g830) & (!g1914) & (!g1900) & (!g3668) & (!g3686) & (g3687)) + ((!g830) & (!g1914) & (!g1900) & (!g3668) & (g3686) & (g3687)) + ((!g830) & (!g1914) & (!g1900) & (g3668) & (!g3686) & (g3687)) + ((!g830) & (!g1914) & (!g1900) & (g3668) & (g3686) & (g3687)) + ((!g830) & (!g1914) & (g1900) & (!g3668) & (!g3686) & (g3687)) + ((!g830) & (!g1914) & (g1900) & (!g3668) & (g3686) & (g3687)) + ((!g830) & (!g1914) & (g1900) & (g3668) & (!g3686) & (g3687)) + ((!g830) & (!g1914) & (g1900) & (g3668) & (g3686) & (g3687)) + ((!g830) & (g1914) & (!g1900) & (!g3668) & (!g3686) & (g3687)) + ((!g830) & (g1914) & (!g1900) & (!g3668) & (g3686) & (g3687)) + ((!g830) & (g1914) & (!g1900) & (g3668) & (!g3686) & (g3687)) + ((!g830) & (g1914) & (!g1900) & (g3668) & (g3686) & (g3687)) + ((!g830) & (g1914) & (g1900) & (!g3668) & (!g3686) & (g3687)) + ((!g830) & (g1914) & (g1900) & (!g3668) & (g3686) & (g3687)) + ((!g830) & (g1914) & (g1900) & (g3668) & (!g3686) & (g3687)) + ((!g830) & (g1914) & (g1900) & (g3668) & (g3686) & (g3687)) + ((g830) & (!g1914) & (!g1900) & (!g3668) & (g3686) & (!g3687)) + ((g830) & (!g1914) & (!g1900) & (!g3668) & (g3686) & (g3687)) + ((g830) & (!g1914) & (!g1900) & (g3668) & (g3686) & (!g3687)) + ((g830) & (!g1914) & (!g1900) & (g3668) & (g3686) & (g3687)) + ((g830) & (!g1914) & (g1900) & (!g3668) & (!g3686) & (!g3687)) + ((g830) & (!g1914) & (g1900) & (!g3668) & (!g3686) & (g3687)) + ((g830) & (!g1914) & (g1900) & (g3668) & (!g3686) & (!g3687)) + ((g830) & (!g1914) & (g1900) & (g3668) & (!g3686) & (g3687)) + ((g830) & (g1914) & (!g1900) & (g3668) & (!g3686) & (!g3687)) + ((g830) & (g1914) & (!g1900) & (g3668) & (!g3686) & (g3687)) + ((g830) & (g1914) & (!g1900) & (g3668) & (g3686) & (!g3687)) + ((g830) & (g1914) & (!g1900) & (g3668) & (g3686) & (g3687)) + ((g830) & (g1914) & (g1900) & (!g3668) & (!g3686) & (!g3687)) + ((g830) & (g1914) & (g1900) & (!g3668) & (!g3686) & (g3687)) + ((g830) & (g1914) & (g1900) & (!g3668) & (g3686) & (!g3687)) + ((g830) & (g1914) & (g1900) & (!g3668) & (g3686) & (g3687)));
	assign g3689 = (((!g1886) & (!g2032) & (g2055) & (!g1910) & (!g2038) & (g2088)) + ((!g1886) & (!g2032) & (g2055) & (!g1910) & (g2038) & (g2088)) + ((!g1886) & (!g2032) & (g2055) & (g1910) & (!g2038) & (g2088)) + ((!g1886) & (!g2032) & (g2055) & (g1910) & (g2038) & (g2088)) + ((!g1886) & (g2032) & (!g2055) & (!g1910) & (g2038) & (g2088)) + ((!g1886) & (g2032) & (!g2055) & (g1910) & (g2038) & (g2088)) + ((!g1886) & (g2032) & (g2055) & (!g1910) & (!g2038) & (g2088)) + ((!g1886) & (g2032) & (g2055) & (!g1910) & (g2038) & (!g2088)) + ((!g1886) & (g2032) & (g2055) & (!g1910) & (g2038) & (g2088)) + ((!g1886) & (g2032) & (g2055) & (g1910) & (!g2038) & (g2088)) + ((!g1886) & (g2032) & (g2055) & (g1910) & (g2038) & (!g2088)) + ((!g1886) & (g2032) & (g2055) & (g1910) & (g2038) & (g2088)) + ((g1886) & (!g2032) & (!g2055) & (g1910) & (g2038) & (g2088)) + ((g1886) & (!g2032) & (g2055) & (!g1910) & (!g2038) & (g2088)) + ((g1886) & (!g2032) & (g2055) & (!g1910) & (g2038) & (g2088)) + ((g1886) & (!g2032) & (g2055) & (g1910) & (!g2038) & (g2088)) + ((g1886) & (!g2032) & (g2055) & (g1910) & (g2038) & (!g2088)) + ((g1886) & (!g2032) & (g2055) & (g1910) & (g2038) & (g2088)) + ((g1886) & (g2032) & (!g2055) & (!g1910) & (g2038) & (g2088)) + ((g1886) & (g2032) & (!g2055) & (g1910) & (!g2038) & (g2088)) + ((g1886) & (g2032) & (!g2055) & (g1910) & (g2038) & (g2088)) + ((g1886) & (g2032) & (g2055) & (!g1910) & (!g2038) & (g2088)) + ((g1886) & (g2032) & (g2055) & (!g1910) & (g2038) & (!g2088)) + ((g1886) & (g2032) & (g2055) & (!g1910) & (g2038) & (g2088)) + ((g1886) & (g2032) & (g2055) & (g1910) & (!g2038) & (!g2088)) + ((g1886) & (g2032) & (g2055) & (g1910) & (!g2038) & (g2088)) + ((g1886) & (g2032) & (g2055) & (g1910) & (g2038) & (!g2088)) + ((g1886) & (g2032) & (g2055) & (g1910) & (g2038) & (g2088)));
	assign g3690 = (((!g2194) & (g2200)) + ((g2194) & (!g2200)));
	assign g3691 = (((!g2114) & (!g2137) & (g2120) & (g2170) & (g3689) & (g3690)) + ((!g2114) & (g2137) & (!g2120) & (g2170) & (!g3689) & (g3690)) + ((!g2114) & (g2137) & (!g2120) & (g2170) & (g3689) & (g3690)) + ((!g2114) & (g2137) & (g2120) & (!g2170) & (g3689) & (g3690)) + ((!g2114) & (g2137) & (g2120) & (g2170) & (!g3689) & (g3690)) + ((!g2114) & (g2137) & (g2120) & (g2170) & (g3689) & (g3690)) + ((g2114) & (!g2137) & (!g2120) & (g2170) & (g3689) & (g3690)) + ((g2114) & (!g2137) & (g2120) & (g2170) & (!g3689) & (g3690)) + ((g2114) & (!g2137) & (g2120) & (g2170) & (g3689) & (g3690)) + ((g2114) & (g2137) & (!g2120) & (!g2170) & (g3689) & (g3690)) + ((g2114) & (g2137) & (!g2120) & (g2170) & (!g3689) & (g3690)) + ((g2114) & (g2137) & (!g2120) & (g2170) & (g3689) & (g3690)) + ((g2114) & (g2137) & (g2120) & (!g2170) & (!g3689) & (g3690)) + ((g2114) & (g2137) & (g2120) & (!g2170) & (g3689) & (g3690)) + ((g2114) & (g2137) & (g2120) & (g2170) & (!g3689) & (g3690)) + ((g2114) & (g2137) & (g2120) & (g2170) & (g3689) & (g3690)));
	assign g3692 = (((g2194) & (g2200)));
	assign g3693 = (((!g2217) & (!g2277) & (g2250) & (g2283) & (!g3691) & (g3692)) + ((!g2217) & (!g2277) & (g2250) & (g2283) & (g3691) & (!g3692)) + ((!g2217) & (!g2277) & (g2250) & (g2283) & (g3691) & (g3692)) + ((!g2217) & (g2277) & (!g2250) & (g2283) & (!g3691) & (!g3692)) + ((!g2217) & (g2277) & (!g2250) & (g2283) & (!g3691) & (g3692)) + ((!g2217) & (g2277) & (!g2250) & (g2283) & (g3691) & (!g3692)) + ((!g2217) & (g2277) & (!g2250) & (g2283) & (g3691) & (g3692)) + ((!g2217) & (g2277) & (g2250) & (!g2283) & (!g3691) & (g3692)) + ((!g2217) & (g2277) & (g2250) & (!g2283) & (g3691) & (!g3692)) + ((!g2217) & (g2277) & (g2250) & (!g2283) & (g3691) & (g3692)) + ((!g2217) & (g2277) & (g2250) & (g2283) & (!g3691) & (!g3692)) + ((!g2217) & (g2277) & (g2250) & (g2283) & (!g3691) & (g3692)) + ((!g2217) & (g2277) & (g2250) & (g2283) & (g3691) & (!g3692)) + ((!g2217) & (g2277) & (g2250) & (g2283) & (g3691) & (g3692)) + ((g2217) & (!g2277) & (!g2250) & (g2283) & (!g3691) & (g3692)) + ((g2217) & (!g2277) & (!g2250) & (g2283) & (g3691) & (!g3692)) + ((g2217) & (!g2277) & (!g2250) & (g2283) & (g3691) & (g3692)) + ((g2217) & (!g2277) & (g2250) & (g2283) & (!g3691) & (!g3692)) + ((g2217) & (!g2277) & (g2250) & (g2283) & (!g3691) & (g3692)) + ((g2217) & (!g2277) & (g2250) & (g2283) & (g3691) & (!g3692)) + ((g2217) & (!g2277) & (g2250) & (g2283) & (g3691) & (g3692)) + ((g2217) & (g2277) & (!g2250) & (!g2283) & (!g3691) & (g3692)) + ((g2217) & (g2277) & (!g2250) & (!g2283) & (g3691) & (!g3692)) + ((g2217) & (g2277) & (!g2250) & (!g2283) & (g3691) & (g3692)) + ((g2217) & (g2277) & (!g2250) & (g2283) & (!g3691) & (!g3692)) + ((g2217) & (g2277) & (!g2250) & (g2283) & (!g3691) & (g3692)) + ((g2217) & (g2277) & (!g2250) & (g2283) & (g3691) & (!g3692)) + ((g2217) & (g2277) & (!g2250) & (g2283) & (g3691) & (g3692)) + ((g2217) & (g2277) & (g2250) & (!g2283) & (!g3691) & (!g3692)) + ((g2217) & (g2277) & (g2250) & (!g2283) & (!g3691) & (g3692)) + ((g2217) & (g2277) & (g2250) & (!g2283) & (g3691) & (!g3692)) + ((g2217) & (g2277) & (g2250) & (!g2283) & (g3691) & (g3692)) + ((g2217) & (g2277) & (g2250) & (g2283) & (!g3691) & (!g3692)) + ((g2217) & (g2277) & (g2250) & (g2283) & (!g3691) & (g3692)) + ((g2217) & (g2277) & (g2250) & (g2283) & (g3691) & (!g3692)) + ((g2217) & (g2277) & (g2250) & (g2283) & (g3691) & (g3692)));
	assign g3694 = (((!g2383) & (g2416)) + ((g2383) & (!g2416)));
	assign g3695 = (((!g2304) & (!g2360) & (g2337) & (g2366) & (g3693) & (g3694)) + ((!g2304) & (g2360) & (!g2337) & (g2366) & (!g3693) & (g3694)) + ((!g2304) & (g2360) & (!g2337) & (g2366) & (g3693) & (g3694)) + ((!g2304) & (g2360) & (g2337) & (!g2366) & (g3693) & (g3694)) + ((!g2304) & (g2360) & (g2337) & (g2366) & (!g3693) & (g3694)) + ((!g2304) & (g2360) & (g2337) & (g2366) & (g3693) & (g3694)) + ((g2304) & (!g2360) & (!g2337) & (g2366) & (g3693) & (g3694)) + ((g2304) & (!g2360) & (g2337) & (g2366) & (!g3693) & (g3694)) + ((g2304) & (!g2360) & (g2337) & (g2366) & (g3693) & (g3694)) + ((g2304) & (g2360) & (!g2337) & (!g2366) & (g3693) & (g3694)) + ((g2304) & (g2360) & (!g2337) & (g2366) & (!g3693) & (g3694)) + ((g2304) & (g2360) & (!g2337) & (g2366) & (g3693) & (g3694)) + ((g2304) & (g2360) & (g2337) & (!g2366) & (!g3693) & (g3694)) + ((g2304) & (g2360) & (g2337) & (!g2366) & (g3693) & (g3694)) + ((g2304) & (g2360) & (g2337) & (g2366) & (!g3693) & (g3694)) + ((g2304) & (g2360) & (g2337) & (g2366) & (g3693) & (g3694)));
	assign g3696 = (((g2383) & (g2416)));
	assign g3697 = (((!g2468) & (!g2523) & (g2486) & (g2544) & (!g3695) & (g3696)) + ((!g2468) & (!g2523) & (g2486) & (g2544) & (g3695) & (!g3696)) + ((!g2468) & (!g2523) & (g2486) & (g2544) & (g3695) & (g3696)) + ((!g2468) & (g2523) & (!g2486) & (g2544) & (!g3695) & (!g3696)) + ((!g2468) & (g2523) & (!g2486) & (g2544) & (!g3695) & (g3696)) + ((!g2468) & (g2523) & (!g2486) & (g2544) & (g3695) & (!g3696)) + ((!g2468) & (g2523) & (!g2486) & (g2544) & (g3695) & (g3696)) + ((!g2468) & (g2523) & (g2486) & (!g2544) & (!g3695) & (g3696)) + ((!g2468) & (g2523) & (g2486) & (!g2544) & (g3695) & (!g3696)) + ((!g2468) & (g2523) & (g2486) & (!g2544) & (g3695) & (g3696)) + ((!g2468) & (g2523) & (g2486) & (g2544) & (!g3695) & (!g3696)) + ((!g2468) & (g2523) & (g2486) & (g2544) & (!g3695) & (g3696)) + ((!g2468) & (g2523) & (g2486) & (g2544) & (g3695) & (!g3696)) + ((!g2468) & (g2523) & (g2486) & (g2544) & (g3695) & (g3696)) + ((g2468) & (!g2523) & (!g2486) & (g2544) & (!g3695) & (g3696)) + ((g2468) & (!g2523) & (!g2486) & (g2544) & (g3695) & (!g3696)) + ((g2468) & (!g2523) & (!g2486) & (g2544) & (g3695) & (g3696)) + ((g2468) & (!g2523) & (g2486) & (g2544) & (!g3695) & (!g3696)) + ((g2468) & (!g2523) & (g2486) & (g2544) & (!g3695) & (g3696)) + ((g2468) & (!g2523) & (g2486) & (g2544) & (g3695) & (!g3696)) + ((g2468) & (!g2523) & (g2486) & (g2544) & (g3695) & (g3696)) + ((g2468) & (g2523) & (!g2486) & (!g2544) & (!g3695) & (g3696)) + ((g2468) & (g2523) & (!g2486) & (!g2544) & (g3695) & (!g3696)) + ((g2468) & (g2523) & (!g2486) & (!g2544) & (g3695) & (g3696)) + ((g2468) & (g2523) & (!g2486) & (g2544) & (!g3695) & (!g3696)) + ((g2468) & (g2523) & (!g2486) & (g2544) & (!g3695) & (g3696)) + ((g2468) & (g2523) & (!g2486) & (g2544) & (g3695) & (!g3696)) + ((g2468) & (g2523) & (!g2486) & (g2544) & (g3695) & (g3696)) + ((g2468) & (g2523) & (g2486) & (!g2544) & (!g3695) & (!g3696)) + ((g2468) & (g2523) & (g2486) & (!g2544) & (!g3695) & (g3696)) + ((g2468) & (g2523) & (g2486) & (!g2544) & (g3695) & (!g3696)) + ((g2468) & (g2523) & (g2486) & (!g2544) & (g3695) & (g3696)) + ((g2468) & (g2523) & (g2486) & (g2544) & (!g3695) & (!g3696)) + ((g2468) & (g2523) & (g2486) & (g2544) & (!g3695) & (g3696)) + ((g2468) & (g2523) & (g2486) & (g2544) & (g3695) & (!g3696)) + ((g2468) & (g2523) & (g2486) & (g2544) & (g3695) & (g3696)));
	assign g3698 = (((!g2575) & (g2584) & (g3697)) + ((g2575) & (!g2584) & (g3697)) + ((g2575) & (g2584) & (!g3697)) + ((g2575) & (g2584) & (g3697)));
	assign g3699 = (((!g1898) & (!g2022) & (g2071) & (!g1904) & (!g2043) & (g2080)) + ((!g1898) & (!g2022) & (g2071) & (!g1904) & (g2043) & (g2080)) + ((!g1898) & (!g2022) & (g2071) & (g1904) & (!g2043) & (g2080)) + ((!g1898) & (!g2022) & (g2071) & (g1904) & (g2043) & (g2080)) + ((!g1898) & (g2022) & (!g2071) & (!g1904) & (g2043) & (g2080)) + ((!g1898) & (g2022) & (!g2071) & (g1904) & (g2043) & (g2080)) + ((!g1898) & (g2022) & (g2071) & (!g1904) & (!g2043) & (g2080)) + ((!g1898) & (g2022) & (g2071) & (!g1904) & (g2043) & (!g2080)) + ((!g1898) & (g2022) & (g2071) & (!g1904) & (g2043) & (g2080)) + ((!g1898) & (g2022) & (g2071) & (g1904) & (!g2043) & (g2080)) + ((!g1898) & (g2022) & (g2071) & (g1904) & (g2043) & (!g2080)) + ((!g1898) & (g2022) & (g2071) & (g1904) & (g2043) & (g2080)) + ((g1898) & (!g2022) & (!g2071) & (g1904) & (g2043) & (g2080)) + ((g1898) & (!g2022) & (g2071) & (!g1904) & (!g2043) & (g2080)) + ((g1898) & (!g2022) & (g2071) & (!g1904) & (g2043) & (g2080)) + ((g1898) & (!g2022) & (g2071) & (g1904) & (!g2043) & (g2080)) + ((g1898) & (!g2022) & (g2071) & (g1904) & (g2043) & (!g2080)) + ((g1898) & (!g2022) & (g2071) & (g1904) & (g2043) & (g2080)) + ((g1898) & (g2022) & (!g2071) & (!g1904) & (g2043) & (g2080)) + ((g1898) & (g2022) & (!g2071) & (g1904) & (!g2043) & (g2080)) + ((g1898) & (g2022) & (!g2071) & (g1904) & (g2043) & (g2080)) + ((g1898) & (g2022) & (g2071) & (!g1904) & (!g2043) & (g2080)) + ((g1898) & (g2022) & (g2071) & (!g1904) & (g2043) & (!g2080)) + ((g1898) & (g2022) & (g2071) & (!g1904) & (g2043) & (g2080)) + ((g1898) & (g2022) & (g2071) & (g1904) & (!g2043) & (!g2080)) + ((g1898) & (g2022) & (g2071) & (g1904) & (!g2043) & (g2080)) + ((g1898) & (g2022) & (g2071) & (g1904) & (g2043) & (!g2080)) + ((g1898) & (g2022) & (g2071) & (g1904) & (g2043) & (g2080)));
	assign g3700 = (((!g2184) & (g2205)) + ((g2184) & (!g2205)));
	assign g3701 = (((!g2104) & (!g2153) & (g2125) & (g2162) & (g3699) & (g3700)) + ((!g2104) & (g2153) & (!g2125) & (g2162) & (!g3699) & (g3700)) + ((!g2104) & (g2153) & (!g2125) & (g2162) & (g3699) & (g3700)) + ((!g2104) & (g2153) & (g2125) & (!g2162) & (g3699) & (g3700)) + ((!g2104) & (g2153) & (g2125) & (g2162) & (!g3699) & (g3700)) + ((!g2104) & (g2153) & (g2125) & (g2162) & (g3699) & (g3700)) + ((g2104) & (!g2153) & (!g2125) & (g2162) & (g3699) & (g3700)) + ((g2104) & (!g2153) & (g2125) & (g2162) & (!g3699) & (g3700)) + ((g2104) & (!g2153) & (g2125) & (g2162) & (g3699) & (g3700)) + ((g2104) & (g2153) & (!g2125) & (!g2162) & (g3699) & (g3700)) + ((g2104) & (g2153) & (!g2125) & (g2162) & (!g3699) & (g3700)) + ((g2104) & (g2153) & (!g2125) & (g2162) & (g3699) & (g3700)) + ((g2104) & (g2153) & (g2125) & (!g2162) & (!g3699) & (g3700)) + ((g2104) & (g2153) & (g2125) & (!g2162) & (g3699) & (g3700)) + ((g2104) & (g2153) & (g2125) & (g2162) & (!g3699) & (g3700)) + ((g2104) & (g2153) & (g2125) & (g2162) & (g3699) & (g3700)));
	assign g3702 = (((g2184) & (g2205)));
	assign g3703 = (((!g2233) & (!g2267) & (!g2242) & (!g2288) & (!g3701) & (!g3702)) + ((!g2233) & (!g2267) & (!g2242) & (!g2288) & (!g3701) & (g3702)) + ((!g2233) & (!g2267) & (!g2242) & (!g2288) & (g3701) & (!g3702)) + ((!g2233) & (!g2267) & (!g2242) & (!g2288) & (g3701) & (g3702)) + ((!g2233) & (!g2267) & (!g2242) & (g2288) & (!g3701) & (!g3702)) + ((!g2233) & (!g2267) & (!g2242) & (g2288) & (!g3701) & (g3702)) + ((!g2233) & (!g2267) & (!g2242) & (g2288) & (g3701) & (!g3702)) + ((!g2233) & (!g2267) & (!g2242) & (g2288) & (g3701) & (g3702)) + ((!g2233) & (!g2267) & (g2242) & (!g2288) & (!g3701) & (!g3702)) + ((!g2233) & (!g2267) & (g2242) & (!g2288) & (!g3701) & (g3702)) + ((!g2233) & (!g2267) & (g2242) & (!g2288) & (g3701) & (!g3702)) + ((!g2233) & (!g2267) & (g2242) & (!g2288) & (g3701) & (g3702)) + ((!g2233) & (!g2267) & (g2242) & (g2288) & (!g3701) & (!g3702)) + ((!g2233) & (g2267) & (!g2242) & (!g2288) & (!g3701) & (!g3702)) + ((!g2233) & (g2267) & (!g2242) & (!g2288) & (!g3701) & (g3702)) + ((!g2233) & (g2267) & (!g2242) & (!g2288) & (g3701) & (!g3702)) + ((!g2233) & (g2267) & (!g2242) & (!g2288) & (g3701) & (g3702)) + ((!g2233) & (g2267) & (g2242) & (!g2288) & (!g3701) & (!g3702)) + ((g2233) & (!g2267) & (!g2242) & (!g2288) & (!g3701) & (!g3702)) + ((g2233) & (!g2267) & (!g2242) & (!g2288) & (!g3701) & (g3702)) + ((g2233) & (!g2267) & (!g2242) & (!g2288) & (g3701) & (!g3702)) + ((g2233) & (!g2267) & (!g2242) & (!g2288) & (g3701) & (g3702)) + ((g2233) & (!g2267) & (!g2242) & (g2288) & (!g3701) & (!g3702)) + ((g2233) & (!g2267) & (g2242) & (!g2288) & (!g3701) & (!g3702)) + ((g2233) & (!g2267) & (g2242) & (!g2288) & (!g3701) & (g3702)) + ((g2233) & (!g2267) & (g2242) & (!g2288) & (g3701) & (!g3702)) + ((g2233) & (!g2267) & (g2242) & (!g2288) & (g3701) & (g3702)) + ((g2233) & (g2267) & (!g2242) & (!g2288) & (!g3701) & (!g3702)));
	assign g3704 = (((!g2320) & (!g2350) & (g2329) & (g2371) & (!g3703)) + ((!g2320) & (g2350) & (!g2329) & (g2371) & (!g3703)) + ((!g2320) & (g2350) & (!g2329) & (g2371) & (g3703)) + ((!g2320) & (g2350) & (g2329) & (!g2371) & (!g3703)) + ((!g2320) & (g2350) & (g2329) & (g2371) & (!g3703)) + ((!g2320) & (g2350) & (g2329) & (g2371) & (g3703)) + ((g2320) & (!g2350) & (!g2329) & (g2371) & (!g3703)) + ((g2320) & (!g2350) & (g2329) & (g2371) & (!g3703)) + ((g2320) & (!g2350) & (g2329) & (g2371) & (g3703)) + ((g2320) & (g2350) & (!g2329) & (!g2371) & (!g3703)) + ((g2320) & (g2350) & (!g2329) & (g2371) & (!g3703)) + ((g2320) & (g2350) & (!g2329) & (g2371) & (g3703)) + ((g2320) & (g2350) & (g2329) & (!g2371) & (!g3703)) + ((g2320) & (g2350) & (g2329) & (!g2371) & (g3703)) + ((g2320) & (g2350) & (g2329) & (g2371) & (!g3703)) + ((g2320) & (g2350) & (g2329) & (g2371) & (g3703)));
	assign g3705 = (((!g2533) & (g2539)) + ((g2533) & (!g2539)));
	assign g3706 = (((!g2399) & (!g2434) & (g2408) & (g2503) & (g3704) & (g3705)) + ((!g2399) & (g2434) & (!g2408) & (g2503) & (!g3704) & (g3705)) + ((!g2399) & (g2434) & (!g2408) & (g2503) & (g3704) & (g3705)) + ((!g2399) & (g2434) & (g2408) & (!g2503) & (g3704) & (g3705)) + ((!g2399) & (g2434) & (g2408) & (g2503) & (!g3704) & (g3705)) + ((!g2399) & (g2434) & (g2408) & (g2503) & (g3704) & (g3705)) + ((g2399) & (!g2434) & (!g2408) & (g2503) & (g3704) & (g3705)) + ((g2399) & (!g2434) & (g2408) & (g2503) & (!g3704) & (g3705)) + ((g2399) & (!g2434) & (g2408) & (g2503) & (g3704) & (g3705)) + ((g2399) & (g2434) & (!g2408) & (!g2503) & (g3704) & (g3705)) + ((g2399) & (g2434) & (!g2408) & (g2503) & (!g3704) & (g3705)) + ((g2399) & (g2434) & (!g2408) & (g2503) & (g3704) & (g3705)) + ((g2399) & (g2434) & (g2408) & (!g2503) & (!g3704) & (g3705)) + ((g2399) & (g2434) & (g2408) & (!g2503) & (g3704) & (g3705)) + ((g2399) & (g2434) & (g2408) & (g2503) & (!g3704) & (g3705)) + ((g2399) & (g2434) & (g2408) & (g2503) & (g3704) & (g3705)));
	assign g3707 = (((g2533) & (g2539)));
	assign g3708 = (((!g3706) & (!g3707)));
	assign g3709 = (((!g2559) & (!g2623) & (!g2592) & (g2632) & (!g3708)) + ((!g2559) & (!g2623) & (!g2592) & (g2632) & (g3708)) + ((!g2559) & (!g2623) & (g2592) & (!g2632) & (!g3708)) + ((!g2559) & (!g2623) & (g2592) & (g2632) & (g3708)) + ((!g2559) & (g2623) & (!g2592) & (!g2632) & (!g3708)) + ((!g2559) & (g2623) & (!g2592) & (!g2632) & (g3708)) + ((!g2559) & (g2623) & (g2592) & (!g2632) & (g3708)) + ((!g2559) & (g2623) & (g2592) & (g2632) & (!g3708)) + ((g2559) & (!g2623) & (!g2592) & (!g2632) & (!g3708)) + ((g2559) & (!g2623) & (!g2592) & (g2632) & (g3708)) + ((g2559) & (!g2623) & (g2592) & (!g2632) & (!g3708)) + ((g2559) & (!g2623) & (g2592) & (!g2632) & (g3708)) + ((g2559) & (g2623) & (!g2592) & (!g2632) & (g3708)) + ((g2559) & (g2623) & (!g2592) & (g2632) & (!g3708)) + ((g2559) & (g2623) & (g2592) & (g2632) & (!g3708)) + ((g2559) & (g2623) & (g2592) & (g2632) & (g3708)));
	assign g3710 = (((!g1888) & (!g1978) & (g1980) & (!g1912) & (!g2045) & (g2091)) + ((!g1888) & (!g1978) & (g1980) & (!g1912) & (g2045) & (g2091)) + ((!g1888) & (!g1978) & (g1980) & (g1912) & (!g2045) & (g2091)) + ((!g1888) & (!g1978) & (g1980) & (g1912) & (g2045) & (g2091)) + ((!g1888) & (g1978) & (!g1980) & (!g1912) & (g2045) & (g2091)) + ((!g1888) & (g1978) & (!g1980) & (g1912) & (g2045) & (g2091)) + ((!g1888) & (g1978) & (g1980) & (!g1912) & (!g2045) & (g2091)) + ((!g1888) & (g1978) & (g1980) & (!g1912) & (g2045) & (!g2091)) + ((!g1888) & (g1978) & (g1980) & (!g1912) & (g2045) & (g2091)) + ((!g1888) & (g1978) & (g1980) & (g1912) & (!g2045) & (g2091)) + ((!g1888) & (g1978) & (g1980) & (g1912) & (g2045) & (!g2091)) + ((!g1888) & (g1978) & (g1980) & (g1912) & (g2045) & (g2091)) + ((g1888) & (!g1978) & (!g1980) & (g1912) & (g2045) & (g2091)) + ((g1888) & (!g1978) & (g1980) & (!g1912) & (!g2045) & (g2091)) + ((g1888) & (!g1978) & (g1980) & (!g1912) & (g2045) & (g2091)) + ((g1888) & (!g1978) & (g1980) & (g1912) & (!g2045) & (g2091)) + ((g1888) & (!g1978) & (g1980) & (g1912) & (g2045) & (!g2091)) + ((g1888) & (!g1978) & (g1980) & (g1912) & (g2045) & (g2091)) + ((g1888) & (g1978) & (!g1980) & (!g1912) & (g2045) & (g2091)) + ((g1888) & (g1978) & (!g1980) & (g1912) & (!g2045) & (g2091)) + ((g1888) & (g1978) & (!g1980) & (g1912) & (g2045) & (g2091)) + ((g1888) & (g1978) & (g1980) & (!g1912) & (!g2045) & (g2091)) + ((g1888) & (g1978) & (g1980) & (!g1912) & (g2045) & (!g2091)) + ((g1888) & (g1978) & (g1980) & (!g1912) & (g2045) & (g2091)) + ((g1888) & (g1978) & (g1980) & (g1912) & (!g2045) & (!g2091)) + ((g1888) & (g1978) & (g1980) & (g1912) & (!g2045) & (g2091)) + ((g1888) & (g1978) & (g1980) & (g1912) & (g2045) & (!g2091)) + ((g1888) & (g1978) & (g1980) & (g1912) & (g2045) & (g2091)));
	assign g3711 = (((!g1987) & (g2207)) + ((g1987) & (!g2207)));
	assign g3712 = (((!g1983) & (!g1985) & (g2127) & (g2173) & (g3710) & (g3711)) + ((!g1983) & (g1985) & (!g2127) & (g2173) & (!g3710) & (g3711)) + ((!g1983) & (g1985) & (!g2127) & (g2173) & (g3710) & (g3711)) + ((!g1983) & (g1985) & (g2127) & (!g2173) & (g3710) & (g3711)) + ((!g1983) & (g1985) & (g2127) & (g2173) & (!g3710) & (g3711)) + ((!g1983) & (g1985) & (g2127) & (g2173) & (g3710) & (g3711)) + ((g1983) & (!g1985) & (!g2127) & (g2173) & (g3710) & (g3711)) + ((g1983) & (!g1985) & (g2127) & (g2173) & (!g3710) & (g3711)) + ((g1983) & (!g1985) & (g2127) & (g2173) & (g3710) & (g3711)) + ((g1983) & (g1985) & (!g2127) & (!g2173) & (g3710) & (g3711)) + ((g1983) & (g1985) & (!g2127) & (g2173) & (!g3710) & (g3711)) + ((g1983) & (g1985) & (!g2127) & (g2173) & (g3710) & (g3711)) + ((g1983) & (g1985) & (g2127) & (!g2173) & (!g3710) & (g3711)) + ((g1983) & (g1985) & (g2127) & (!g2173) & (g3710) & (g3711)) + ((g1983) & (g1985) & (g2127) & (g2173) & (!g3710) & (g3711)) + ((g1983) & (g1985) & (g2127) & (g2173) & (g3710) & (g3711)));
	assign g3713 = (((g1987) & (g2207)));
	assign g3714 = (((!g1992) & (!g1994) & (!g2253) & (!g2290) & (!g3712) & (!g3713)) + ((!g1992) & (!g1994) & (!g2253) & (!g2290) & (!g3712) & (g3713)) + ((!g1992) & (!g1994) & (!g2253) & (!g2290) & (g3712) & (!g3713)) + ((!g1992) & (!g1994) & (!g2253) & (!g2290) & (g3712) & (g3713)) + ((!g1992) & (!g1994) & (!g2253) & (g2290) & (!g3712) & (!g3713)) + ((!g1992) & (!g1994) & (!g2253) & (g2290) & (!g3712) & (g3713)) + ((!g1992) & (!g1994) & (!g2253) & (g2290) & (g3712) & (!g3713)) + ((!g1992) & (!g1994) & (!g2253) & (g2290) & (g3712) & (g3713)) + ((!g1992) & (!g1994) & (g2253) & (!g2290) & (!g3712) & (!g3713)) + ((!g1992) & (!g1994) & (g2253) & (!g2290) & (!g3712) & (g3713)) + ((!g1992) & (!g1994) & (g2253) & (!g2290) & (g3712) & (!g3713)) + ((!g1992) & (!g1994) & (g2253) & (!g2290) & (g3712) & (g3713)) + ((!g1992) & (!g1994) & (g2253) & (g2290) & (!g3712) & (!g3713)) + ((!g1992) & (g1994) & (!g2253) & (!g2290) & (!g3712) & (!g3713)) + ((!g1992) & (g1994) & (!g2253) & (!g2290) & (!g3712) & (g3713)) + ((!g1992) & (g1994) & (!g2253) & (!g2290) & (g3712) & (!g3713)) + ((!g1992) & (g1994) & (!g2253) & (!g2290) & (g3712) & (g3713)) + ((!g1992) & (g1994) & (g2253) & (!g2290) & (!g3712) & (!g3713)) + ((g1992) & (!g1994) & (!g2253) & (!g2290) & (!g3712) & (!g3713)) + ((g1992) & (!g1994) & (!g2253) & (!g2290) & (!g3712) & (g3713)) + ((g1992) & (!g1994) & (!g2253) & (!g2290) & (g3712) & (!g3713)) + ((g1992) & (!g1994) & (!g2253) & (!g2290) & (g3712) & (g3713)) + ((g1992) & (!g1994) & (!g2253) & (g2290) & (!g3712) & (!g3713)) + ((g1992) & (!g1994) & (g2253) & (!g2290) & (!g3712) & (!g3713)) + ((g1992) & (!g1994) & (g2253) & (!g2290) & (!g3712) & (g3713)) + ((g1992) & (!g1994) & (g2253) & (!g2290) & (g3712) & (!g3713)) + ((g1992) & (!g1994) & (g2253) & (!g2290) & (g3712) & (g3713)) + ((g1992) & (g1994) & (!g2253) & (!g2290) & (!g3712) & (!g3713)));
	assign g3715 = (((!g2002) & (g2419)) + ((g2002) & (!g2419)));
	assign g3716 = (((!g1997) & (!g1999) & (g2340) & (g2373) & (!g3714) & (g3715)) + ((!g1997) & (g1999) & (!g2340) & (g2373) & (!g3714) & (g3715)) + ((!g1997) & (g1999) & (!g2340) & (g2373) & (g3714) & (g3715)) + ((!g1997) & (g1999) & (g2340) & (!g2373) & (!g3714) & (g3715)) + ((!g1997) & (g1999) & (g2340) & (g2373) & (!g3714) & (g3715)) + ((!g1997) & (g1999) & (g2340) & (g2373) & (g3714) & (g3715)) + ((g1997) & (!g1999) & (!g2340) & (g2373) & (!g3714) & (g3715)) + ((g1997) & (!g1999) & (g2340) & (g2373) & (!g3714) & (g3715)) + ((g1997) & (!g1999) & (g2340) & (g2373) & (g3714) & (g3715)) + ((g1997) & (g1999) & (!g2340) & (!g2373) & (!g3714) & (g3715)) + ((g1997) & (g1999) & (!g2340) & (g2373) & (!g3714) & (g3715)) + ((g1997) & (g1999) & (!g2340) & (g2373) & (g3714) & (g3715)) + ((g1997) & (g1999) & (g2340) & (!g2373) & (!g3714) & (g3715)) + ((g1997) & (g1999) & (g2340) & (!g2373) & (g3714) & (g3715)) + ((g1997) & (g1999) & (g2340) & (g2373) & (!g3714) & (g3715)) + ((g1997) & (g1999) & (g2340) & (g2373) & (g3714) & (g3715)));
	assign g3717 = (((g2002) & (g2419)));
	assign g3718 = (((!g2004) & (!g2006) & (!g2509) & (!g2546) & (!g3716) & (!g3717)) + ((!g2004) & (!g2006) & (!g2509) & (!g2546) & (!g3716) & (g3717)) + ((!g2004) & (!g2006) & (!g2509) & (!g2546) & (g3716) & (!g3717)) + ((!g2004) & (!g2006) & (!g2509) & (!g2546) & (g3716) & (g3717)) + ((!g2004) & (!g2006) & (!g2509) & (g2546) & (!g3716) & (!g3717)) + ((!g2004) & (!g2006) & (!g2509) & (g2546) & (!g3716) & (g3717)) + ((!g2004) & (!g2006) & (!g2509) & (g2546) & (g3716) & (!g3717)) + ((!g2004) & (!g2006) & (!g2509) & (g2546) & (g3716) & (g3717)) + ((!g2004) & (!g2006) & (g2509) & (!g2546) & (!g3716) & (!g3717)) + ((!g2004) & (!g2006) & (g2509) & (!g2546) & (!g3716) & (g3717)) + ((!g2004) & (!g2006) & (g2509) & (!g2546) & (g3716) & (!g3717)) + ((!g2004) & (!g2006) & (g2509) & (!g2546) & (g3716) & (g3717)) + ((!g2004) & (!g2006) & (g2509) & (g2546) & (!g3716) & (!g3717)) + ((!g2004) & (g2006) & (!g2509) & (!g2546) & (!g3716) & (!g3717)) + ((!g2004) & (g2006) & (!g2509) & (!g2546) & (!g3716) & (g3717)) + ((!g2004) & (g2006) & (!g2509) & (!g2546) & (g3716) & (!g3717)) + ((!g2004) & (g2006) & (!g2509) & (!g2546) & (g3716) & (g3717)) + ((!g2004) & (g2006) & (g2509) & (!g2546) & (!g3716) & (!g3717)) + ((g2004) & (!g2006) & (!g2509) & (!g2546) & (!g3716) & (!g3717)) + ((g2004) & (!g2006) & (!g2509) & (!g2546) & (!g3716) & (g3717)) + ((g2004) & (!g2006) & (!g2509) & (!g2546) & (g3716) & (!g3717)) + ((g2004) & (!g2006) & (!g2509) & (!g2546) & (g3716) & (g3717)) + ((g2004) & (!g2006) & (!g2509) & (g2546) & (!g3716) & (!g3717)) + ((g2004) & (!g2006) & (g2509) & (!g2546) & (!g3716) & (!g3717)) + ((g2004) & (!g2006) & (g2509) & (!g2546) & (!g3716) & (g3717)) + ((g2004) & (!g2006) & (g2509) & (!g2546) & (g3716) & (!g3717)) + ((g2004) & (!g2006) & (g2509) & (!g2546) & (g3716) & (g3717)) + ((g2004) & (g2006) & (!g2509) & (!g2546) & (!g3716) & (!g3717)));
	assign g3719 = (((!g2004) & (!g2509) & (!g3716) & (!g3717) & (!g5818) & (g5819)) + ((!g2004) & (!g2509) & (!g3716) & (g3717) & (!g5818) & (g5819)) + ((!g2004) & (!g2509) & (g3716) & (!g3717) & (!g5818) & (g5819)) + ((!g2004) & (!g2509) & (g3716) & (g3717) & (!g5818) & (g5819)) + ((!g2004) & (g2509) & (!g3716) & (!g3717) & (!g5818) & (g5819)) + ((!g2004) & (g2509) & (!g3716) & (g3717) & (!g5818) & (g5819)) + ((!g2004) & (g2509) & (!g3716) & (g3717) & (g5818) & (g5819)) + ((!g2004) & (g2509) & (g3716) & (!g3717) & (!g5818) & (g5819)) + ((!g2004) & (g2509) & (g3716) & (!g3717) & (g5818) & (g5819)) + ((!g2004) & (g2509) & (g3716) & (g3717) & (!g5818) & (g5819)) + ((!g2004) & (g2509) & (g3716) & (g3717) & (g5818) & (g5819)) + ((g2004) & (!g2509) & (!g3716) & (!g3717) & (!g5818) & (g5819)) + ((g2004) & (!g2509) & (!g3716) & (g3717) & (!g5818) & (g5819)) + ((g2004) & (!g2509) & (!g3716) & (g3717) & (g5818) & (g5819)) + ((g2004) & (!g2509) & (g3716) & (!g3717) & (!g5818) & (g5819)) + ((g2004) & (!g2509) & (g3716) & (!g3717) & (g5818) & (g5819)) + ((g2004) & (!g2509) & (g3716) & (g3717) & (!g5818) & (g5819)) + ((g2004) & (!g2509) & (g3716) & (g3717) & (g5818) & (g5819)) + ((g2004) & (g2509) & (!g3716) & (!g3717) & (!g5818) & (g5819)) + ((g2004) & (g2509) & (!g3716) & (!g3717) & (g5818) & (g5819)) + ((g2004) & (g2509) & (!g3716) & (g3717) & (!g5818) & (g5819)) + ((g2004) & (g2509) & (!g3716) & (g3717) & (g5818) & (g5819)) + ((g2004) & (g2509) & (g3716) & (!g3717) & (!g5818) & (g5819)) + ((g2004) & (g2509) & (g3716) & (!g3717) & (g5818) & (g5819)) + ((g2004) & (g2509) & (g3716) & (g3717) & (!g5818) & (g5819)) + ((g2004) & (g2509) & (g3716) & (g3717) & (g5818) & (g5819)));
	assign g3720 = (((g2052) & (g2676)));
	assign g3721 = (((!g2101) & (!g2134) & (!g2752) & (!g2787) & (!g3719) & (!g3720)) + ((!g2101) & (!g2134) & (!g2752) & (!g2787) & (!g3719) & (g3720)) + ((!g2101) & (!g2134) & (!g2752) & (!g2787) & (g3719) & (!g3720)) + ((!g2101) & (!g2134) & (!g2752) & (!g2787) & (g3719) & (g3720)) + ((!g2101) & (!g2134) & (!g2752) & (g2787) & (!g3719) & (!g3720)) + ((!g2101) & (!g2134) & (!g2752) & (g2787) & (!g3719) & (g3720)) + ((!g2101) & (!g2134) & (!g2752) & (g2787) & (g3719) & (!g3720)) + ((!g2101) & (!g2134) & (!g2752) & (g2787) & (g3719) & (g3720)) + ((!g2101) & (!g2134) & (g2752) & (!g2787) & (!g3719) & (!g3720)) + ((!g2101) & (!g2134) & (g2752) & (!g2787) & (!g3719) & (g3720)) + ((!g2101) & (!g2134) & (g2752) & (!g2787) & (g3719) & (!g3720)) + ((!g2101) & (!g2134) & (g2752) & (!g2787) & (g3719) & (g3720)) + ((!g2101) & (!g2134) & (g2752) & (g2787) & (!g3719) & (!g3720)) + ((!g2101) & (g2134) & (!g2752) & (!g2787) & (!g3719) & (!g3720)) + ((!g2101) & (g2134) & (!g2752) & (!g2787) & (!g3719) & (g3720)) + ((!g2101) & (g2134) & (!g2752) & (!g2787) & (g3719) & (!g3720)) + ((!g2101) & (g2134) & (!g2752) & (!g2787) & (g3719) & (g3720)) + ((!g2101) & (g2134) & (g2752) & (!g2787) & (!g3719) & (!g3720)) + ((g2101) & (!g2134) & (!g2752) & (!g2787) & (!g3719) & (!g3720)) + ((g2101) & (!g2134) & (!g2752) & (!g2787) & (!g3719) & (g3720)) + ((g2101) & (!g2134) & (!g2752) & (!g2787) & (g3719) & (!g3720)) + ((g2101) & (!g2134) & (!g2752) & (!g2787) & (g3719) & (g3720)) + ((g2101) & (!g2134) & (!g2752) & (g2787) & (!g3719) & (!g3720)) + ((g2101) & (!g2134) & (g2752) & (!g2787) & (!g3719) & (!g3720)) + ((g2101) & (!g2134) & (g2752) & (!g2787) & (!g3719) & (g3720)) + ((g2101) & (!g2134) & (g2752) & (!g2787) & (g3719) & (!g3720)) + ((g2101) & (!g2134) & (g2752) & (!g2787) & (g3719) & (g3720)) + ((g2101) & (g2134) & (!g2752) & (!g2787) & (!g3719) & (!g3720)));
	assign g3722 = (((!g2263) & (g2904)) + ((g2263) & (!g2904)));
	assign g3723 = (((!g2181) & (!g2213) & (g2833) & (g2874) & (!g3721) & (g3722)) + ((!g2181) & (g2213) & (!g2833) & (g2874) & (!g3721) & (g3722)) + ((!g2181) & (g2213) & (!g2833) & (g2874) & (g3721) & (g3722)) + ((!g2181) & (g2213) & (g2833) & (!g2874) & (!g3721) & (g3722)) + ((!g2181) & (g2213) & (g2833) & (g2874) & (!g3721) & (g3722)) + ((!g2181) & (g2213) & (g2833) & (g2874) & (g3721) & (g3722)) + ((g2181) & (!g2213) & (!g2833) & (g2874) & (!g3721) & (g3722)) + ((g2181) & (!g2213) & (g2833) & (g2874) & (!g3721) & (g3722)) + ((g2181) & (!g2213) & (g2833) & (g2874) & (g3721) & (g3722)) + ((g2181) & (g2213) & (!g2833) & (!g2874) & (!g3721) & (g3722)) + ((g2181) & (g2213) & (!g2833) & (g2874) & (!g3721) & (g3722)) + ((g2181) & (g2213) & (!g2833) & (g2874) & (g3721) & (g3722)) + ((g2181) & (g2213) & (g2833) & (!g2874) & (!g3721) & (g3722)) + ((g2181) & (g2213) & (g2833) & (!g2874) & (g3721) & (g3722)) + ((g2181) & (g2213) & (g2833) & (g2874) & (!g3721) & (g3722)) + ((g2181) & (g2213) & (g2833) & (g2874) & (g3721) & (g3722)));
	assign g3724 = (((g2263) & (g2904)));
	assign g3725 = (((!g2299) & (!g2348) & (!g2991) & (!g3022) & (!g3723) & (!g3724)) + ((!g2299) & (!g2348) & (!g2991) & (!g3022) & (!g3723) & (g3724)) + ((!g2299) & (!g2348) & (!g2991) & (!g3022) & (g3723) & (!g3724)) + ((!g2299) & (!g2348) & (!g2991) & (!g3022) & (g3723) & (g3724)) + ((!g2299) & (!g2348) & (!g2991) & (g3022) & (!g3723) & (!g3724)) + ((!g2299) & (!g2348) & (!g2991) & (g3022) & (!g3723) & (g3724)) + ((!g2299) & (!g2348) & (!g2991) & (g3022) & (g3723) & (!g3724)) + ((!g2299) & (!g2348) & (!g2991) & (g3022) & (g3723) & (g3724)) + ((!g2299) & (!g2348) & (g2991) & (!g3022) & (!g3723) & (!g3724)) + ((!g2299) & (!g2348) & (g2991) & (!g3022) & (!g3723) & (g3724)) + ((!g2299) & (!g2348) & (g2991) & (!g3022) & (g3723) & (!g3724)) + ((!g2299) & (!g2348) & (g2991) & (!g3022) & (g3723) & (g3724)) + ((!g2299) & (!g2348) & (g2991) & (g3022) & (!g3723) & (!g3724)) + ((!g2299) & (g2348) & (!g2991) & (!g3022) & (!g3723) & (!g3724)) + ((!g2299) & (g2348) & (!g2991) & (!g3022) & (!g3723) & (g3724)) + ((!g2299) & (g2348) & (!g2991) & (!g3022) & (g3723) & (!g3724)) + ((!g2299) & (g2348) & (!g2991) & (!g3022) & (g3723) & (g3724)) + ((!g2299) & (g2348) & (g2991) & (!g3022) & (!g3723) & (!g3724)) + ((g2299) & (!g2348) & (!g2991) & (!g3022) & (!g3723) & (!g3724)) + ((g2299) & (!g2348) & (!g2991) & (!g3022) & (!g3723) & (g3724)) + ((g2299) & (!g2348) & (!g2991) & (!g3022) & (g3723) & (!g3724)) + ((g2299) & (!g2348) & (!g2991) & (!g3022) & (g3723) & (g3724)) + ((g2299) & (!g2348) & (!g2991) & (g3022) & (!g3723) & (!g3724)) + ((g2299) & (!g2348) & (g2991) & (!g3022) & (!g3723) & (!g3724)) + ((g2299) & (!g2348) & (g2991) & (!g3022) & (!g3723) & (g3724)) + ((g2299) & (!g2348) & (g2991) & (!g3022) & (g3723) & (!g3724)) + ((g2299) & (!g2348) & (g2991) & (!g3022) & (g3723) & (g3724)) + ((g2299) & (g2348) & (!g2991) & (!g3022) & (!g3723) & (!g3724)));
	assign g3726 = (((g1914) & (!g2379) & (!g3067) & (!g3725)) + ((g1914) & (!g2379) & (g3067) & (g3725)) + ((g1914) & (g2379) & (!g3067) & (g3725)) + ((g1914) & (g2379) & (g3067) & (!g3725)));
	assign g3727 = (((!g1900) & (!g2028) & (g2074) & (!g1902) & (!g2036) & (g2077)) + ((!g1900) & (!g2028) & (g2074) & (!g1902) & (g2036) & (g2077)) + ((!g1900) & (!g2028) & (g2074) & (g1902) & (!g2036) & (g2077)) + ((!g1900) & (!g2028) & (g2074) & (g1902) & (g2036) & (g2077)) + ((!g1900) & (g2028) & (!g2074) & (!g1902) & (g2036) & (g2077)) + ((!g1900) & (g2028) & (!g2074) & (g1902) & (g2036) & (g2077)) + ((!g1900) & (g2028) & (g2074) & (!g1902) & (!g2036) & (g2077)) + ((!g1900) & (g2028) & (g2074) & (!g1902) & (g2036) & (!g2077)) + ((!g1900) & (g2028) & (g2074) & (!g1902) & (g2036) & (g2077)) + ((!g1900) & (g2028) & (g2074) & (g1902) & (!g2036) & (g2077)) + ((!g1900) & (g2028) & (g2074) & (g1902) & (g2036) & (!g2077)) + ((!g1900) & (g2028) & (g2074) & (g1902) & (g2036) & (g2077)) + ((g1900) & (!g2028) & (!g2074) & (g1902) & (g2036) & (g2077)) + ((g1900) & (!g2028) & (g2074) & (!g1902) & (!g2036) & (g2077)) + ((g1900) & (!g2028) & (g2074) & (!g1902) & (g2036) & (g2077)) + ((g1900) & (!g2028) & (g2074) & (g1902) & (!g2036) & (g2077)) + ((g1900) & (!g2028) & (g2074) & (g1902) & (g2036) & (!g2077)) + ((g1900) & (!g2028) & (g2074) & (g1902) & (g2036) & (g2077)) + ((g1900) & (g2028) & (!g2074) & (!g1902) & (g2036) & (g2077)) + ((g1900) & (g2028) & (!g2074) & (g1902) & (!g2036) & (g2077)) + ((g1900) & (g2028) & (!g2074) & (g1902) & (g2036) & (g2077)) + ((g1900) & (g2028) & (g2074) & (!g1902) & (!g2036) & (g2077)) + ((g1900) & (g2028) & (g2074) & (!g1902) & (g2036) & (!g2077)) + ((g1900) & (g2028) & (g2074) & (!g1902) & (g2036) & (g2077)) + ((g1900) & (g2028) & (g2074) & (g1902) & (!g2036) & (!g2077)) + ((g1900) & (g2028) & (g2074) & (g1902) & (!g2036) & (g2077)) + ((g1900) & (g2028) & (g2074) & (g1902) & (g2036) & (!g2077)) + ((g1900) & (g2028) & (g2074) & (g1902) & (g2036) & (g2077)));
	assign g3728 = (((!g2190) & (g2198)) + ((g2190) & (!g2198)));
	assign g3729 = (((!g2110) & (!g2156) & (g2118) & (g2159) & (g3727) & (g3728)) + ((!g2110) & (g2156) & (!g2118) & (g2159) & (!g3727) & (g3728)) + ((!g2110) & (g2156) & (!g2118) & (g2159) & (g3727) & (g3728)) + ((!g2110) & (g2156) & (g2118) & (!g2159) & (g3727) & (g3728)) + ((!g2110) & (g2156) & (g2118) & (g2159) & (!g3727) & (g3728)) + ((!g2110) & (g2156) & (g2118) & (g2159) & (g3727) & (g3728)) + ((g2110) & (!g2156) & (!g2118) & (g2159) & (g3727) & (g3728)) + ((g2110) & (!g2156) & (g2118) & (g2159) & (!g3727) & (g3728)) + ((g2110) & (!g2156) & (g2118) & (g2159) & (g3727) & (g3728)) + ((g2110) & (g2156) & (!g2118) & (!g2159) & (g3727) & (g3728)) + ((g2110) & (g2156) & (!g2118) & (g2159) & (!g3727) & (g3728)) + ((g2110) & (g2156) & (!g2118) & (g2159) & (g3727) & (g3728)) + ((g2110) & (g2156) & (g2118) & (!g2159) & (!g3727) & (g3728)) + ((g2110) & (g2156) & (g2118) & (!g2159) & (g3727) & (g3728)) + ((g2110) & (g2156) & (g2118) & (g2159) & (!g3727) & (g3728)) + ((g2110) & (g2156) & (g2118) & (g2159) & (g3727) & (g3728)));
	assign g3730 = (((g2190) & (g2198)));
	assign g3731 = (((!g2236) & (!g2273) & (!g2239) & (!g2281) & (!g3729) & (!g3730)) + ((!g2236) & (!g2273) & (!g2239) & (!g2281) & (!g3729) & (g3730)) + ((!g2236) & (!g2273) & (!g2239) & (!g2281) & (g3729) & (!g3730)) + ((!g2236) & (!g2273) & (!g2239) & (!g2281) & (g3729) & (g3730)) + ((!g2236) & (!g2273) & (!g2239) & (g2281) & (!g3729) & (!g3730)) + ((!g2236) & (!g2273) & (!g2239) & (g2281) & (!g3729) & (g3730)) + ((!g2236) & (!g2273) & (!g2239) & (g2281) & (g3729) & (!g3730)) + ((!g2236) & (!g2273) & (!g2239) & (g2281) & (g3729) & (g3730)) + ((!g2236) & (!g2273) & (g2239) & (!g2281) & (!g3729) & (!g3730)) + ((!g2236) & (!g2273) & (g2239) & (!g2281) & (!g3729) & (g3730)) + ((!g2236) & (!g2273) & (g2239) & (!g2281) & (g3729) & (!g3730)) + ((!g2236) & (!g2273) & (g2239) & (!g2281) & (g3729) & (g3730)) + ((!g2236) & (!g2273) & (g2239) & (g2281) & (!g3729) & (!g3730)) + ((!g2236) & (g2273) & (!g2239) & (!g2281) & (!g3729) & (!g3730)) + ((!g2236) & (g2273) & (!g2239) & (!g2281) & (!g3729) & (g3730)) + ((!g2236) & (g2273) & (!g2239) & (!g2281) & (g3729) & (!g3730)) + ((!g2236) & (g2273) & (!g2239) & (!g2281) & (g3729) & (g3730)) + ((!g2236) & (g2273) & (g2239) & (!g2281) & (!g3729) & (!g3730)) + ((g2236) & (!g2273) & (!g2239) & (!g2281) & (!g3729) & (!g3730)) + ((g2236) & (!g2273) & (!g2239) & (!g2281) & (!g3729) & (g3730)) + ((g2236) & (!g2273) & (!g2239) & (!g2281) & (g3729) & (!g3730)) + ((g2236) & (!g2273) & (!g2239) & (!g2281) & (g3729) & (g3730)) + ((g2236) & (!g2273) & (!g2239) & (g2281) & (!g3729) & (!g3730)) + ((g2236) & (!g2273) & (g2239) & (!g2281) & (!g3729) & (!g3730)) + ((g2236) & (!g2273) & (g2239) & (!g2281) & (!g3729) & (g3730)) + ((g2236) & (!g2273) & (g2239) & (!g2281) & (g3729) & (!g3730)) + ((g2236) & (!g2273) & (g2239) & (!g2281) & (g3729) & (g3730)) + ((g2236) & (g2273) & (!g2239) & (!g2281) & (!g3729) & (!g3730)));
	assign g3732 = (((!g2402) & (g2405)) + ((g2402) & (!g2405)));
	assign g3733 = (((!g2323) & (!g2356) & (g2326) & (g2364) & (!g3731) & (g3732)) + ((!g2323) & (g2356) & (!g2326) & (g2364) & (!g3731) & (g3732)) + ((!g2323) & (g2356) & (!g2326) & (g2364) & (g3731) & (g3732)) + ((!g2323) & (g2356) & (g2326) & (!g2364) & (!g3731) & (g3732)) + ((!g2323) & (g2356) & (g2326) & (g2364) & (!g3731) & (g3732)) + ((!g2323) & (g2356) & (g2326) & (g2364) & (g3731) & (g3732)) + ((g2323) & (!g2356) & (!g2326) & (g2364) & (!g3731) & (g3732)) + ((g2323) & (!g2356) & (g2326) & (g2364) & (!g3731) & (g3732)) + ((g2323) & (!g2356) & (g2326) & (g2364) & (g3731) & (g3732)) + ((g2323) & (g2356) & (!g2326) & (!g2364) & (!g3731) & (g3732)) + ((g2323) & (g2356) & (!g2326) & (g2364) & (!g3731) & (g3732)) + ((g2323) & (g2356) & (!g2326) & (g2364) & (g3731) & (g3732)) + ((g2323) & (g2356) & (g2326) & (!g2364) & (!g3731) & (g3732)) + ((g2323) & (g2356) & (g2326) & (!g2364) & (g3731) & (g3732)) + ((g2323) & (g2356) & (g2326) & (g2364) & (!g3731) & (g3732)) + ((g2323) & (g2356) & (g2326) & (g2364) & (g3731) & (g3732)));
	assign g3734 = (((g2402) & (g2405)));
	assign g3735 = (((!g2456) & (!g2535) & (!g2480) & (!g2537) & (!g3733) & (!g3734)) + ((!g2456) & (!g2535) & (!g2480) & (!g2537) & (!g3733) & (g3734)) + ((!g2456) & (!g2535) & (!g2480) & (!g2537) & (g3733) & (!g3734)) + ((!g2456) & (!g2535) & (!g2480) & (!g2537) & (g3733) & (g3734)) + ((!g2456) & (!g2535) & (!g2480) & (g2537) & (!g3733) & (!g3734)) + ((!g2456) & (!g2535) & (!g2480) & (g2537) & (!g3733) & (g3734)) + ((!g2456) & (!g2535) & (!g2480) & (g2537) & (g3733) & (!g3734)) + ((!g2456) & (!g2535) & (!g2480) & (g2537) & (g3733) & (g3734)) + ((!g2456) & (!g2535) & (g2480) & (!g2537) & (!g3733) & (!g3734)) + ((!g2456) & (!g2535) & (g2480) & (!g2537) & (!g3733) & (g3734)) + ((!g2456) & (!g2535) & (g2480) & (!g2537) & (g3733) & (!g3734)) + ((!g2456) & (!g2535) & (g2480) & (!g2537) & (g3733) & (g3734)) + ((!g2456) & (!g2535) & (g2480) & (g2537) & (!g3733) & (!g3734)) + ((!g2456) & (g2535) & (!g2480) & (!g2537) & (!g3733) & (!g3734)) + ((!g2456) & (g2535) & (!g2480) & (!g2537) & (!g3733) & (g3734)) + ((!g2456) & (g2535) & (!g2480) & (!g2537) & (g3733) & (!g3734)) + ((!g2456) & (g2535) & (!g2480) & (!g2537) & (g3733) & (g3734)) + ((!g2456) & (g2535) & (g2480) & (!g2537) & (!g3733) & (!g3734)) + ((g2456) & (!g2535) & (!g2480) & (!g2537) & (!g3733) & (!g3734)) + ((g2456) & (!g2535) & (!g2480) & (!g2537) & (!g3733) & (g3734)) + ((g2456) & (!g2535) & (!g2480) & (!g2537) & (g3733) & (!g3734)) + ((g2456) & (!g2535) & (!g2480) & (!g2537) & (g3733) & (g3734)) + ((g2456) & (!g2535) & (!g2480) & (g2537) & (!g3733) & (!g3734)) + ((g2456) & (!g2535) & (g2480) & (!g2537) & (!g3733) & (!g3734)) + ((g2456) & (!g2535) & (g2480) & (!g2537) & (!g3733) & (g3734)) + ((g2456) & (!g2535) & (g2480) & (!g2537) & (g3733) & (!g3734)) + ((g2456) & (!g2535) & (g2480) & (!g2537) & (g3733) & (g3734)) + ((g2456) & (g2535) & (!g2480) & (!g2537) & (!g3733) & (!g3734)));
	assign g3736 = (((!g2456) & (!g2480) & (!g3733) & (!g3734) & (!g5821) & (g5822)) + ((!g2456) & (!g2480) & (!g3733) & (g3734) & (!g5821) & (g5822)) + ((!g2456) & (!g2480) & (g3733) & (!g3734) & (!g5821) & (g5822)) + ((!g2456) & (!g2480) & (g3733) & (g3734) & (!g5821) & (g5822)) + ((!g2456) & (g2480) & (!g3733) & (!g3734) & (!g5821) & (g5822)) + ((!g2456) & (g2480) & (!g3733) & (g3734) & (!g5821) & (g5822)) + ((!g2456) & (g2480) & (!g3733) & (g3734) & (g5821) & (g5822)) + ((!g2456) & (g2480) & (g3733) & (!g3734) & (!g5821) & (g5822)) + ((!g2456) & (g2480) & (g3733) & (!g3734) & (g5821) & (g5822)) + ((!g2456) & (g2480) & (g3733) & (g3734) & (!g5821) & (g5822)) + ((!g2456) & (g2480) & (g3733) & (g3734) & (g5821) & (g5822)) + ((g2456) & (!g2480) & (!g3733) & (!g3734) & (!g5821) & (g5822)) + ((g2456) & (!g2480) & (!g3733) & (g3734) & (!g5821) & (g5822)) + ((g2456) & (!g2480) & (!g3733) & (g3734) & (g5821) & (g5822)) + ((g2456) & (!g2480) & (g3733) & (!g3734) & (!g5821) & (g5822)) + ((g2456) & (!g2480) & (g3733) & (!g3734) & (g5821) & (g5822)) + ((g2456) & (!g2480) & (g3733) & (g3734) & (!g5821) & (g5822)) + ((g2456) & (!g2480) & (g3733) & (g3734) & (g5821) & (g5822)) + ((g2456) & (g2480) & (!g3733) & (!g3734) & (!g5821) & (g5822)) + ((g2456) & (g2480) & (!g3733) & (!g3734) & (g5821) & (g5822)) + ((g2456) & (g2480) & (!g3733) & (g3734) & (!g5821) & (g5822)) + ((g2456) & (g2480) & (!g3733) & (g3734) & (g5821) & (g5822)) + ((g2456) & (g2480) & (g3733) & (!g3734) & (!g5821) & (g5822)) + ((g2456) & (g2480) & (g3733) & (!g3734) & (g5821) & (g5822)) + ((g2456) & (g2480) & (g3733) & (g3734) & (!g5821) & (g5822)) + ((g2456) & (g2480) & (g3733) & (g3734) & (g5821) & (g5822)));
	assign g3737 = (((g2667) & (g2659)));
	assign g3738 = (((!g2728) & (!g2778) & (!g2723) & (!g2770) & (!g3736) & (!g3737)) + ((!g2728) & (!g2778) & (!g2723) & (!g2770) & (!g3736) & (g3737)) + ((!g2728) & (!g2778) & (!g2723) & (!g2770) & (g3736) & (!g3737)) + ((!g2728) & (!g2778) & (!g2723) & (!g2770) & (g3736) & (g3737)) + ((!g2728) & (!g2778) & (!g2723) & (g2770) & (!g3736) & (!g3737)) + ((!g2728) & (!g2778) & (!g2723) & (g2770) & (!g3736) & (g3737)) + ((!g2728) & (!g2778) & (!g2723) & (g2770) & (g3736) & (!g3737)) + ((!g2728) & (!g2778) & (!g2723) & (g2770) & (g3736) & (g3737)) + ((!g2728) & (!g2778) & (g2723) & (!g2770) & (!g3736) & (!g3737)) + ((!g2728) & (!g2778) & (g2723) & (!g2770) & (!g3736) & (g3737)) + ((!g2728) & (!g2778) & (g2723) & (!g2770) & (g3736) & (!g3737)) + ((!g2728) & (!g2778) & (g2723) & (!g2770) & (g3736) & (g3737)) + ((!g2728) & (!g2778) & (g2723) & (g2770) & (!g3736) & (!g3737)) + ((!g2728) & (g2778) & (!g2723) & (!g2770) & (!g3736) & (!g3737)) + ((!g2728) & (g2778) & (!g2723) & (!g2770) & (!g3736) & (g3737)) + ((!g2728) & (g2778) & (!g2723) & (!g2770) & (g3736) & (!g3737)) + ((!g2728) & (g2778) & (!g2723) & (!g2770) & (g3736) & (g3737)) + ((!g2728) & (g2778) & (g2723) & (!g2770) & (!g3736) & (!g3737)) + ((g2728) & (!g2778) & (!g2723) & (!g2770) & (!g3736) & (!g3737)) + ((g2728) & (!g2778) & (!g2723) & (!g2770) & (!g3736) & (g3737)) + ((g2728) & (!g2778) & (!g2723) & (!g2770) & (g3736) & (!g3737)) + ((g2728) & (!g2778) & (!g2723) & (!g2770) & (g3736) & (g3737)) + ((g2728) & (!g2778) & (!g2723) & (g2770) & (!g3736) & (!g3737)) + ((g2728) & (!g2778) & (g2723) & (!g2770) & (!g3736) & (!g3737)) + ((g2728) & (!g2778) & (g2723) & (!g2770) & (!g3736) & (g3737)) + ((g2728) & (!g2778) & (g2723) & (!g2770) & (g3736) & (!g3737)) + ((g2728) & (!g2778) & (g2723) & (!g2770) & (g3736) & (g3737)) + ((g2728) & (g2778) & (!g2723) & (!g2770) & (!g3736) & (!g3737)));
	assign g3739 = (((!g2895) & (g2893)) + ((g2895) & (!g2893)));
	assign g3740 = (((!g2819) & (!g2860) & (g2816) & (g2848) & (!g3738) & (g3739)) + ((!g2819) & (g2860) & (!g2816) & (g2848) & (!g3738) & (g3739)) + ((!g2819) & (g2860) & (!g2816) & (g2848) & (g3738) & (g3739)) + ((!g2819) & (g2860) & (g2816) & (!g2848) & (!g3738) & (g3739)) + ((!g2819) & (g2860) & (g2816) & (g2848) & (!g3738) & (g3739)) + ((!g2819) & (g2860) & (g2816) & (g2848) & (g3738) & (g3739)) + ((g2819) & (!g2860) & (!g2816) & (g2848) & (!g3738) & (g3739)) + ((g2819) & (!g2860) & (g2816) & (g2848) & (!g3738) & (g3739)) + ((g2819) & (!g2860) & (g2816) & (g2848) & (g3738) & (g3739)) + ((g2819) & (g2860) & (!g2816) & (!g2848) & (!g3738) & (g3739)) + ((g2819) & (g2860) & (!g2816) & (g2848) & (!g3738) & (g3739)) + ((g2819) & (g2860) & (!g2816) & (g2848) & (g3738) & (g3739)) + ((g2819) & (g2860) & (g2816) & (!g2848) & (!g3738) & (g3739)) + ((g2819) & (g2860) & (g2816) & (!g2848) & (g3738) & (g3739)) + ((g2819) & (g2860) & (g2816) & (g2848) & (!g3738) & (g3739)) + ((g2819) & (g2860) & (g2816) & (g2848) & (g3738) & (g3739)));
	assign g3741 = (((g2895) & (g2893)));
	assign g3742 = (((!g2962) & (!g3013) & (!g3740) & (!g3741) & (!g2938) & (!g3011)) + ((!g2962) & (!g3013) & (!g3740) & (!g3741) & (!g2938) & (g3011)) + ((!g2962) & (!g3013) & (!g3740) & (!g3741) & (g2938) & (!g3011)) + ((!g2962) & (!g3013) & (!g3740) & (!g3741) & (g2938) & (g3011)) + ((!g2962) & (!g3013) & (!g3740) & (g3741) & (!g2938) & (!g3011)) + ((!g2962) & (!g3013) & (!g3740) & (g3741) & (!g2938) & (g3011)) + ((!g2962) & (!g3013) & (!g3740) & (g3741) & (g2938) & (!g3011)) + ((!g2962) & (!g3013) & (g3740) & (!g3741) & (!g2938) & (!g3011)) + ((!g2962) & (!g3013) & (g3740) & (!g3741) & (!g2938) & (g3011)) + ((!g2962) & (!g3013) & (g3740) & (!g3741) & (g2938) & (!g3011)) + ((!g2962) & (!g3013) & (g3740) & (g3741) & (!g2938) & (!g3011)) + ((!g2962) & (!g3013) & (g3740) & (g3741) & (!g2938) & (g3011)) + ((!g2962) & (!g3013) & (g3740) & (g3741) & (g2938) & (!g3011)) + ((!g2962) & (g3013) & (!g3740) & (!g3741) & (!g2938) & (!g3011)) + ((!g2962) & (g3013) & (!g3740) & (!g3741) & (g2938) & (!g3011)) + ((!g2962) & (g3013) & (!g3740) & (g3741) & (!g2938) & (!g3011)) + ((!g2962) & (g3013) & (g3740) & (!g3741) & (!g2938) & (!g3011)) + ((!g2962) & (g3013) & (g3740) & (g3741) & (!g2938) & (!g3011)) + ((g2962) & (!g3013) & (!g3740) & (!g3741) & (!g2938) & (!g3011)) + ((g2962) & (!g3013) & (!g3740) & (!g3741) & (!g2938) & (g3011)) + ((g2962) & (!g3013) & (!g3740) & (!g3741) & (g2938) & (!g3011)) + ((g2962) & (!g3013) & (!g3740) & (g3741) & (!g2938) & (!g3011)) + ((g2962) & (!g3013) & (!g3740) & (g3741) & (g2938) & (!g3011)) + ((g2962) & (!g3013) & (g3740) & (!g3741) & (!g2938) & (!g3011)) + ((g2962) & (!g3013) & (g3740) & (!g3741) & (g2938) & (!g3011)) + ((g2962) & (!g3013) & (g3740) & (g3741) & (!g2938) & (!g3011)) + ((g2962) & (!g3013) & (g3740) & (g3741) & (g2938) & (!g3011)) + ((g2962) & (g3013) & (!g3740) & (!g3741) & (!g2938) & (!g3011)));
	assign g3743 = (((!g1914) & (!g3053) & (!g3742) & (!g3041)) + ((!g1914) & (!g3053) & (g3742) & (g3041)) + ((!g1914) & (g3053) & (!g3742) & (g3041)) + ((!g1914) & (g3053) & (g3742) & (!g3041)));
	assign g3744 = (((!g830) & (!g1904) & (!g3726) & (!g3743) & (key[192])) + ((!g830) & (!g1904) & (!g3726) & (g3743) & (key[192])) + ((!g830) & (!g1904) & (g3726) & (!g3743) & (key[192])) + ((!g830) & (!g1904) & (g3726) & (g3743) & (key[192])) + ((!g830) & (g1904) & (!g3726) & (!g3743) & (key[192])) + ((!g830) & (g1904) & (!g3726) & (g3743) & (key[192])) + ((!g830) & (g1904) & (g3726) & (!g3743) & (key[192])) + ((!g830) & (g1904) & (g3726) & (g3743) & (key[192])) + ((g830) & (!g1904) & (!g3726) & (g3743) & (!key[192])) + ((g830) & (!g1904) & (!g3726) & (g3743) & (key[192])) + ((g830) & (!g1904) & (g3726) & (!g3743) & (!key[192])) + ((g830) & (!g1904) & (g3726) & (!g3743) & (key[192])) + ((g830) & (!g1904) & (g3726) & (g3743) & (!key[192])) + ((g830) & (!g1904) & (g3726) & (g3743) & (key[192])) + ((g830) & (g1904) & (!g3726) & (!g3743) & (!key[192])) + ((g830) & (g1904) & (!g3726) & (!g3743) & (key[192])));
	assign g3745 = (((!g1890) & (!g1939) & (g1941) & (!g1898) & (!g2022) & (g2071)) + ((!g1890) & (!g1939) & (g1941) & (!g1898) & (g2022) & (g2071)) + ((!g1890) & (!g1939) & (g1941) & (g1898) & (!g2022) & (g2071)) + ((!g1890) & (!g1939) & (g1941) & (g1898) & (g2022) & (g2071)) + ((!g1890) & (g1939) & (!g1941) & (!g1898) & (g2022) & (g2071)) + ((!g1890) & (g1939) & (!g1941) & (g1898) & (g2022) & (g2071)) + ((!g1890) & (g1939) & (g1941) & (!g1898) & (!g2022) & (g2071)) + ((!g1890) & (g1939) & (g1941) & (!g1898) & (g2022) & (!g2071)) + ((!g1890) & (g1939) & (g1941) & (!g1898) & (g2022) & (g2071)) + ((!g1890) & (g1939) & (g1941) & (g1898) & (!g2022) & (g2071)) + ((!g1890) & (g1939) & (g1941) & (g1898) & (g2022) & (!g2071)) + ((!g1890) & (g1939) & (g1941) & (g1898) & (g2022) & (g2071)) + ((g1890) & (!g1939) & (!g1941) & (g1898) & (g2022) & (g2071)) + ((g1890) & (!g1939) & (g1941) & (!g1898) & (!g2022) & (g2071)) + ((g1890) & (!g1939) & (g1941) & (!g1898) & (g2022) & (g2071)) + ((g1890) & (!g1939) & (g1941) & (g1898) & (!g2022) & (g2071)) + ((g1890) & (!g1939) & (g1941) & (g1898) & (g2022) & (!g2071)) + ((g1890) & (!g1939) & (g1941) & (g1898) & (g2022) & (g2071)) + ((g1890) & (g1939) & (!g1941) & (!g1898) & (g2022) & (g2071)) + ((g1890) & (g1939) & (!g1941) & (g1898) & (!g2022) & (g2071)) + ((g1890) & (g1939) & (!g1941) & (g1898) & (g2022) & (g2071)) + ((g1890) & (g1939) & (g1941) & (!g1898) & (!g2022) & (g2071)) + ((g1890) & (g1939) & (g1941) & (!g1898) & (g2022) & (!g2071)) + ((g1890) & (g1939) & (g1941) & (!g1898) & (g2022) & (g2071)) + ((g1890) & (g1939) & (g1941) & (g1898) & (!g2022) & (!g2071)) + ((g1890) & (g1939) & (g1941) & (g1898) & (!g2022) & (g2071)) + ((g1890) & (g1939) & (g1941) & (g1898) & (g2022) & (!g2071)) + ((g1890) & (g1939) & (g1941) & (g1898) & (g2022) & (g2071)));
	assign g3746 = (((!g1948) & (g2184)) + ((g1948) & (!g2184)));
	assign g3747 = (((!g1944) & (!g1946) & (g2104) & (g2153) & (g3745) & (g3746)) + ((!g1944) & (g1946) & (!g2104) & (g2153) & (!g3745) & (g3746)) + ((!g1944) & (g1946) & (!g2104) & (g2153) & (g3745) & (g3746)) + ((!g1944) & (g1946) & (g2104) & (!g2153) & (g3745) & (g3746)) + ((!g1944) & (g1946) & (g2104) & (g2153) & (!g3745) & (g3746)) + ((!g1944) & (g1946) & (g2104) & (g2153) & (g3745) & (g3746)) + ((g1944) & (!g1946) & (!g2104) & (g2153) & (g3745) & (g3746)) + ((g1944) & (!g1946) & (g2104) & (g2153) & (!g3745) & (g3746)) + ((g1944) & (!g1946) & (g2104) & (g2153) & (g3745) & (g3746)) + ((g1944) & (g1946) & (!g2104) & (!g2153) & (g3745) & (g3746)) + ((g1944) & (g1946) & (!g2104) & (g2153) & (!g3745) & (g3746)) + ((g1944) & (g1946) & (!g2104) & (g2153) & (g3745) & (g3746)) + ((g1944) & (g1946) & (g2104) & (!g2153) & (!g3745) & (g3746)) + ((g1944) & (g1946) & (g2104) & (!g2153) & (g3745) & (g3746)) + ((g1944) & (g1946) & (g2104) & (g2153) & (!g3745) & (g3746)) + ((g1944) & (g1946) & (g2104) & (g2153) & (g3745) & (g3746)));
	assign g3748 = (((g1948) & (g2184)));
	assign g3749 = (((!g1953) & (!g1955) & (!g2233) & (!g2267) & (!g3747) & (!g3748)) + ((!g1953) & (!g1955) & (!g2233) & (!g2267) & (!g3747) & (g3748)) + ((!g1953) & (!g1955) & (!g2233) & (!g2267) & (g3747) & (!g3748)) + ((!g1953) & (!g1955) & (!g2233) & (!g2267) & (g3747) & (g3748)) + ((!g1953) & (!g1955) & (!g2233) & (g2267) & (!g3747) & (!g3748)) + ((!g1953) & (!g1955) & (!g2233) & (g2267) & (!g3747) & (g3748)) + ((!g1953) & (!g1955) & (!g2233) & (g2267) & (g3747) & (!g3748)) + ((!g1953) & (!g1955) & (!g2233) & (g2267) & (g3747) & (g3748)) + ((!g1953) & (!g1955) & (g2233) & (!g2267) & (!g3747) & (!g3748)) + ((!g1953) & (!g1955) & (g2233) & (!g2267) & (!g3747) & (g3748)) + ((!g1953) & (!g1955) & (g2233) & (!g2267) & (g3747) & (!g3748)) + ((!g1953) & (!g1955) & (g2233) & (!g2267) & (g3747) & (g3748)) + ((!g1953) & (!g1955) & (g2233) & (g2267) & (!g3747) & (!g3748)) + ((!g1953) & (g1955) & (!g2233) & (!g2267) & (!g3747) & (!g3748)) + ((!g1953) & (g1955) & (!g2233) & (!g2267) & (!g3747) & (g3748)) + ((!g1953) & (g1955) & (!g2233) & (!g2267) & (g3747) & (!g3748)) + ((!g1953) & (g1955) & (!g2233) & (!g2267) & (g3747) & (g3748)) + ((!g1953) & (g1955) & (g2233) & (!g2267) & (!g3747) & (!g3748)) + ((g1953) & (!g1955) & (!g2233) & (!g2267) & (!g3747) & (!g3748)) + ((g1953) & (!g1955) & (!g2233) & (!g2267) & (!g3747) & (g3748)) + ((g1953) & (!g1955) & (!g2233) & (!g2267) & (g3747) & (!g3748)) + ((g1953) & (!g1955) & (!g2233) & (!g2267) & (g3747) & (g3748)) + ((g1953) & (!g1955) & (!g2233) & (g2267) & (!g3747) & (!g3748)) + ((g1953) & (!g1955) & (g2233) & (!g2267) & (!g3747) & (!g3748)) + ((g1953) & (!g1955) & (g2233) & (!g2267) & (!g3747) & (g3748)) + ((g1953) & (!g1955) & (g2233) & (!g2267) & (g3747) & (!g3748)) + ((g1953) & (!g1955) & (g2233) & (!g2267) & (g3747) & (g3748)) + ((g1953) & (g1955) & (!g2233) & (!g2267) & (!g3747) & (!g3748)));
	assign g3750 = (((!g1962) & (g2399)) + ((g1962) & (!g2399)));
	assign g3751 = (((!g1958) & (!g1960) & (g2320) & (g2350) & (!g3749) & (g3750)) + ((!g1958) & (g1960) & (!g2320) & (g2350) & (!g3749) & (g3750)) + ((!g1958) & (g1960) & (!g2320) & (g2350) & (g3749) & (g3750)) + ((!g1958) & (g1960) & (g2320) & (!g2350) & (!g3749) & (g3750)) + ((!g1958) & (g1960) & (g2320) & (g2350) & (!g3749) & (g3750)) + ((!g1958) & (g1960) & (g2320) & (g2350) & (g3749) & (g3750)) + ((g1958) & (!g1960) & (!g2320) & (g2350) & (!g3749) & (g3750)) + ((g1958) & (!g1960) & (g2320) & (g2350) & (!g3749) & (g3750)) + ((g1958) & (!g1960) & (g2320) & (g2350) & (g3749) & (g3750)) + ((g1958) & (g1960) & (!g2320) & (!g2350) & (!g3749) & (g3750)) + ((g1958) & (g1960) & (!g2320) & (g2350) & (!g3749) & (g3750)) + ((g1958) & (g1960) & (!g2320) & (g2350) & (g3749) & (g3750)) + ((g1958) & (g1960) & (g2320) & (!g2350) & (!g3749) & (g3750)) + ((g1958) & (g1960) & (g2320) & (!g2350) & (g3749) & (g3750)) + ((g1958) & (g1960) & (g2320) & (g2350) & (!g3749) & (g3750)) + ((g1958) & (g1960) & (g2320) & (g2350) & (g3749) & (g3750)));
	assign g3752 = (((g1962) & (g2399)));
	assign g3753 = (((!g1967) & (!g1969) & (!g2434) & (!g2533) & (!g3751) & (!g3752)) + ((!g1967) & (!g1969) & (!g2434) & (!g2533) & (!g3751) & (g3752)) + ((!g1967) & (!g1969) & (!g2434) & (!g2533) & (g3751) & (!g3752)) + ((!g1967) & (!g1969) & (!g2434) & (!g2533) & (g3751) & (g3752)) + ((!g1967) & (!g1969) & (!g2434) & (g2533) & (!g3751) & (!g3752)) + ((!g1967) & (!g1969) & (!g2434) & (g2533) & (!g3751) & (g3752)) + ((!g1967) & (!g1969) & (!g2434) & (g2533) & (g3751) & (!g3752)) + ((!g1967) & (!g1969) & (!g2434) & (g2533) & (g3751) & (g3752)) + ((!g1967) & (!g1969) & (g2434) & (!g2533) & (!g3751) & (!g3752)) + ((!g1967) & (!g1969) & (g2434) & (!g2533) & (!g3751) & (g3752)) + ((!g1967) & (!g1969) & (g2434) & (!g2533) & (g3751) & (!g3752)) + ((!g1967) & (!g1969) & (g2434) & (!g2533) & (g3751) & (g3752)) + ((!g1967) & (!g1969) & (g2434) & (g2533) & (!g3751) & (!g3752)) + ((!g1967) & (g1969) & (!g2434) & (!g2533) & (!g3751) & (!g3752)) + ((!g1967) & (g1969) & (!g2434) & (!g2533) & (!g3751) & (g3752)) + ((!g1967) & (g1969) & (!g2434) & (!g2533) & (g3751) & (!g3752)) + ((!g1967) & (g1969) & (!g2434) & (!g2533) & (g3751) & (g3752)) + ((!g1967) & (g1969) & (g2434) & (!g2533) & (!g3751) & (!g3752)) + ((g1967) & (!g1969) & (!g2434) & (!g2533) & (!g3751) & (!g3752)) + ((g1967) & (!g1969) & (!g2434) & (!g2533) & (!g3751) & (g3752)) + ((g1967) & (!g1969) & (!g2434) & (!g2533) & (g3751) & (!g3752)) + ((g1967) & (!g1969) & (!g2434) & (!g2533) & (g3751) & (g3752)) + ((g1967) & (!g1969) & (!g2434) & (g2533) & (!g3751) & (!g3752)) + ((g1967) & (!g1969) & (g2434) & (!g2533) & (!g3751) & (!g3752)) + ((g1967) & (!g1969) & (g2434) & (!g2533) & (!g3751) & (g3752)) + ((g1967) & (!g1969) & (g2434) & (!g2533) & (g3751) & (!g3752)) + ((g1967) & (!g1969) & (g2434) & (!g2533) & (g3751) & (g3752)) + ((g1967) & (g1969) & (!g2434) & (!g2533) & (!g3751) & (!g3752)));
	assign g3754 = (((!g2047) & (g2653)) + ((g2047) & (!g2653)));
	assign g3755 = (((!g1972) & (!g1975) & (g2559) & (g2623) & (!g3753) & (g3754)) + ((!g1972) & (g1975) & (!g2559) & (g2623) & (!g3753) & (g3754)) + ((!g1972) & (g1975) & (!g2559) & (g2623) & (g3753) & (g3754)) + ((!g1972) & (g1975) & (g2559) & (!g2623) & (!g3753) & (g3754)) + ((!g1972) & (g1975) & (g2559) & (g2623) & (!g3753) & (g3754)) + ((!g1972) & (g1975) & (g2559) & (g2623) & (g3753) & (g3754)) + ((g1972) & (!g1975) & (!g2559) & (g2623) & (!g3753) & (g3754)) + ((g1972) & (!g1975) & (g2559) & (g2623) & (!g3753) & (g3754)) + ((g1972) & (!g1975) & (g2559) & (g2623) & (g3753) & (g3754)) + ((g1972) & (g1975) & (!g2559) & (!g2623) & (!g3753) & (g3754)) + ((g1972) & (g1975) & (!g2559) & (g2623) & (!g3753) & (g3754)) + ((g1972) & (g1975) & (!g2559) & (g2623) & (g3753) & (g3754)) + ((g1972) & (g1975) & (g2559) & (!g2623) & (!g3753) & (g3754)) + ((g1972) & (g1975) & (g2559) & (!g2623) & (g3753) & (g3754)) + ((g1972) & (g1975) & (g2559) & (g2623) & (!g3753) & (g3754)) + ((g1972) & (g1975) & (g2559) & (g2623) & (g3753) & (g3754)));
	assign g3756 = (((g2047) & (g2653)));
	assign g3757 = (((!g2098) & (!g2129) & (!g2718) & (!g2764) & (!g3755) & (!g3756)) + ((!g2098) & (!g2129) & (!g2718) & (!g2764) & (!g3755) & (g3756)) + ((!g2098) & (!g2129) & (!g2718) & (!g2764) & (g3755) & (!g3756)) + ((!g2098) & (!g2129) & (!g2718) & (!g2764) & (g3755) & (g3756)) + ((!g2098) & (!g2129) & (!g2718) & (g2764) & (!g3755) & (!g3756)) + ((!g2098) & (!g2129) & (!g2718) & (g2764) & (!g3755) & (g3756)) + ((!g2098) & (!g2129) & (!g2718) & (g2764) & (g3755) & (!g3756)) + ((!g2098) & (!g2129) & (!g2718) & (g2764) & (g3755) & (g3756)) + ((!g2098) & (!g2129) & (g2718) & (!g2764) & (!g3755) & (!g3756)) + ((!g2098) & (!g2129) & (g2718) & (!g2764) & (!g3755) & (g3756)) + ((!g2098) & (!g2129) & (g2718) & (!g2764) & (g3755) & (!g3756)) + ((!g2098) & (!g2129) & (g2718) & (!g2764) & (g3755) & (g3756)) + ((!g2098) & (!g2129) & (g2718) & (g2764) & (!g3755) & (!g3756)) + ((!g2098) & (g2129) & (!g2718) & (!g2764) & (!g3755) & (!g3756)) + ((!g2098) & (g2129) & (!g2718) & (!g2764) & (!g3755) & (g3756)) + ((!g2098) & (g2129) & (!g2718) & (!g2764) & (g3755) & (!g3756)) + ((!g2098) & (g2129) & (!g2718) & (!g2764) & (g3755) & (g3756)) + ((!g2098) & (g2129) & (g2718) & (!g2764) & (!g3755) & (!g3756)) + ((g2098) & (!g2129) & (!g2718) & (!g2764) & (!g3755) & (!g3756)) + ((g2098) & (!g2129) & (!g2718) & (!g2764) & (!g3755) & (g3756)) + ((g2098) & (!g2129) & (!g2718) & (!g2764) & (g3755) & (!g3756)) + ((g2098) & (!g2129) & (!g2718) & (!g2764) & (g3755) & (g3756)) + ((g2098) & (!g2129) & (!g2718) & (g2764) & (!g3755) & (!g3756)) + ((g2098) & (!g2129) & (g2718) & (!g2764) & (!g3755) & (!g3756)) + ((g2098) & (!g2129) & (g2718) & (!g2764) & (!g3755) & (g3756)) + ((g2098) & (!g2129) & (g2718) & (!g2764) & (g3755) & (!g3756)) + ((g2098) & (!g2129) & (g2718) & (!g2764) & (g3755) & (g3756)) + ((g2098) & (g2129) & (!g2718) & (!g2764) & (!g3755) & (!g3756)));
	assign g3758 = (((!g2177) & (g2813) & (!g3757)) + ((g2177) & (!g2813) & (!g3757)) + ((g2177) & (g2813) & (!g3757)) + ((g2177) & (g2813) & (g3757)));
	assign g3759 = (((!g1908) & (!g2030) & (g2085) & (!g1912) & (!g2045) & (g2091)) + ((!g1908) & (!g2030) & (g2085) & (!g1912) & (g2045) & (g2091)) + ((!g1908) & (!g2030) & (g2085) & (g1912) & (!g2045) & (g2091)) + ((!g1908) & (!g2030) & (g2085) & (g1912) & (g2045) & (g2091)) + ((!g1908) & (g2030) & (!g2085) & (!g1912) & (g2045) & (g2091)) + ((!g1908) & (g2030) & (!g2085) & (g1912) & (g2045) & (g2091)) + ((!g1908) & (g2030) & (g2085) & (!g1912) & (!g2045) & (g2091)) + ((!g1908) & (g2030) & (g2085) & (!g1912) & (g2045) & (!g2091)) + ((!g1908) & (g2030) & (g2085) & (!g1912) & (g2045) & (g2091)) + ((!g1908) & (g2030) & (g2085) & (g1912) & (!g2045) & (g2091)) + ((!g1908) & (g2030) & (g2085) & (g1912) & (g2045) & (!g2091)) + ((!g1908) & (g2030) & (g2085) & (g1912) & (g2045) & (g2091)) + ((g1908) & (!g2030) & (!g2085) & (g1912) & (g2045) & (g2091)) + ((g1908) & (!g2030) & (g2085) & (!g1912) & (!g2045) & (g2091)) + ((g1908) & (!g2030) & (g2085) & (!g1912) & (g2045) & (g2091)) + ((g1908) & (!g2030) & (g2085) & (g1912) & (!g2045) & (g2091)) + ((g1908) & (!g2030) & (g2085) & (g1912) & (g2045) & (!g2091)) + ((g1908) & (!g2030) & (g2085) & (g1912) & (g2045) & (g2091)) + ((g1908) & (g2030) & (!g2085) & (!g1912) & (g2045) & (g2091)) + ((g1908) & (g2030) & (!g2085) & (g1912) & (!g2045) & (g2091)) + ((g1908) & (g2030) & (!g2085) & (g1912) & (g2045) & (g2091)) + ((g1908) & (g2030) & (g2085) & (!g1912) & (!g2045) & (g2091)) + ((g1908) & (g2030) & (g2085) & (!g1912) & (g2045) & (!g2091)) + ((g1908) & (g2030) & (g2085) & (!g1912) & (g2045) & (g2091)) + ((g1908) & (g2030) & (g2085) & (g1912) & (!g2045) & (!g2091)) + ((g1908) & (g2030) & (g2085) & (g1912) & (!g2045) & (g2091)) + ((g1908) & (g2030) & (g2085) & (g1912) & (g2045) & (!g2091)) + ((g1908) & (g2030) & (g2085) & (g1912) & (g2045) & (g2091)));
	assign g3760 = (((!g2192) & (g2207)) + ((g2192) & (!g2207)));
	assign g3761 = (((!g2112) & (!g2167) & (g2127) & (g2173) & (g3759) & (g3760)) + ((!g2112) & (g2167) & (!g2127) & (g2173) & (!g3759) & (g3760)) + ((!g2112) & (g2167) & (!g2127) & (g2173) & (g3759) & (g3760)) + ((!g2112) & (g2167) & (g2127) & (!g2173) & (g3759) & (g3760)) + ((!g2112) & (g2167) & (g2127) & (g2173) & (!g3759) & (g3760)) + ((!g2112) & (g2167) & (g2127) & (g2173) & (g3759) & (g3760)) + ((g2112) & (!g2167) & (!g2127) & (g2173) & (g3759) & (g3760)) + ((g2112) & (!g2167) & (g2127) & (g2173) & (!g3759) & (g3760)) + ((g2112) & (!g2167) & (g2127) & (g2173) & (g3759) & (g3760)) + ((g2112) & (g2167) & (!g2127) & (!g2173) & (g3759) & (g3760)) + ((g2112) & (g2167) & (!g2127) & (g2173) & (!g3759) & (g3760)) + ((g2112) & (g2167) & (!g2127) & (g2173) & (g3759) & (g3760)) + ((g2112) & (g2167) & (g2127) & (!g2173) & (!g3759) & (g3760)) + ((g2112) & (g2167) & (g2127) & (!g2173) & (g3759) & (g3760)) + ((g2112) & (g2167) & (g2127) & (g2173) & (!g3759) & (g3760)) + ((g2112) & (g2167) & (g2127) & (g2173) & (g3759) & (g3760)));
	assign g3762 = (((g2192) & (g2207)));
	assign g3763 = (((!g2247) & (!g2275) & (!g2253) & (!g2290) & (!g3761) & (!g3762)) + ((!g2247) & (!g2275) & (!g2253) & (!g2290) & (!g3761) & (g3762)) + ((!g2247) & (!g2275) & (!g2253) & (!g2290) & (g3761) & (!g3762)) + ((!g2247) & (!g2275) & (!g2253) & (!g2290) & (g3761) & (g3762)) + ((!g2247) & (!g2275) & (!g2253) & (g2290) & (!g3761) & (!g3762)) + ((!g2247) & (!g2275) & (!g2253) & (g2290) & (!g3761) & (g3762)) + ((!g2247) & (!g2275) & (!g2253) & (g2290) & (g3761) & (!g3762)) + ((!g2247) & (!g2275) & (!g2253) & (g2290) & (g3761) & (g3762)) + ((!g2247) & (!g2275) & (g2253) & (!g2290) & (!g3761) & (!g3762)) + ((!g2247) & (!g2275) & (g2253) & (!g2290) & (!g3761) & (g3762)) + ((!g2247) & (!g2275) & (g2253) & (!g2290) & (g3761) & (!g3762)) + ((!g2247) & (!g2275) & (g2253) & (!g2290) & (g3761) & (g3762)) + ((!g2247) & (!g2275) & (g2253) & (g2290) & (!g3761) & (!g3762)) + ((!g2247) & (g2275) & (!g2253) & (!g2290) & (!g3761) & (!g3762)) + ((!g2247) & (g2275) & (!g2253) & (!g2290) & (!g3761) & (g3762)) + ((!g2247) & (g2275) & (!g2253) & (!g2290) & (g3761) & (!g3762)) + ((!g2247) & (g2275) & (!g2253) & (!g2290) & (g3761) & (g3762)) + ((!g2247) & (g2275) & (g2253) & (!g2290) & (!g3761) & (!g3762)) + ((g2247) & (!g2275) & (!g2253) & (!g2290) & (!g3761) & (!g3762)) + ((g2247) & (!g2275) & (!g2253) & (!g2290) & (!g3761) & (g3762)) + ((g2247) & (!g2275) & (!g2253) & (!g2290) & (g3761) & (!g3762)) + ((g2247) & (!g2275) & (!g2253) & (!g2290) & (g3761) & (g3762)) + ((g2247) & (!g2275) & (!g2253) & (g2290) & (!g3761) & (!g3762)) + ((g2247) & (!g2275) & (g2253) & (!g2290) & (!g3761) & (!g3762)) + ((g2247) & (!g2275) & (g2253) & (!g2290) & (!g3761) & (g3762)) + ((g2247) & (!g2275) & (g2253) & (!g2290) & (g3761) & (!g3762)) + ((g2247) & (!g2275) & (g2253) & (!g2290) & (g3761) & (g3762)) + ((g2247) & (g2275) & (!g2253) & (!g2290) & (!g3761) & (!g3762)));
	assign g3764 = (((!g2413) & (g2419)) + ((g2413) & (!g2419)));
	assign g3765 = (((!g2334) & (!g2358) & (g2340) & (g2373) & (!g3763) & (g3764)) + ((!g2334) & (g2358) & (!g2340) & (g2373) & (!g3763) & (g3764)) + ((!g2334) & (g2358) & (!g2340) & (g2373) & (g3763) & (g3764)) + ((!g2334) & (g2358) & (g2340) & (!g2373) & (!g3763) & (g3764)) + ((!g2334) & (g2358) & (g2340) & (g2373) & (!g3763) & (g3764)) + ((!g2334) & (g2358) & (g2340) & (g2373) & (g3763) & (g3764)) + ((g2334) & (!g2358) & (!g2340) & (g2373) & (!g3763) & (g3764)) + ((g2334) & (!g2358) & (g2340) & (g2373) & (!g3763) & (g3764)) + ((g2334) & (!g2358) & (g2340) & (g2373) & (g3763) & (g3764)) + ((g2334) & (g2358) & (!g2340) & (!g2373) & (!g3763) & (g3764)) + ((g2334) & (g2358) & (!g2340) & (g2373) & (!g3763) & (g3764)) + ((g2334) & (g2358) & (!g2340) & (g2373) & (g3763) & (g3764)) + ((g2334) & (g2358) & (g2340) & (!g2373) & (!g3763) & (g3764)) + ((g2334) & (g2358) & (g2340) & (!g2373) & (g3763) & (g3764)) + ((g2334) & (g2358) & (g2340) & (g2373) & (!g3763) & (g3764)) + ((g2334) & (g2358) & (g2340) & (g2373) & (g3763) & (g3764)));
	assign g3766 = (((g2413) & (g2419)));
	assign g3767 = (((!g2462) & (!g2542) & (!g2509) & (!g2546) & (!g3765) & (!g3766)) + ((!g2462) & (!g2542) & (!g2509) & (!g2546) & (!g3765) & (g3766)) + ((!g2462) & (!g2542) & (!g2509) & (!g2546) & (g3765) & (!g3766)) + ((!g2462) & (!g2542) & (!g2509) & (!g2546) & (g3765) & (g3766)) + ((!g2462) & (!g2542) & (!g2509) & (g2546) & (!g3765) & (!g3766)) + ((!g2462) & (!g2542) & (!g2509) & (g2546) & (!g3765) & (g3766)) + ((!g2462) & (!g2542) & (!g2509) & (g2546) & (g3765) & (!g3766)) + ((!g2462) & (!g2542) & (!g2509) & (g2546) & (g3765) & (g3766)) + ((!g2462) & (!g2542) & (g2509) & (!g2546) & (!g3765) & (!g3766)) + ((!g2462) & (!g2542) & (g2509) & (!g2546) & (!g3765) & (g3766)) + ((!g2462) & (!g2542) & (g2509) & (!g2546) & (g3765) & (!g3766)) + ((!g2462) & (!g2542) & (g2509) & (!g2546) & (g3765) & (g3766)) + ((!g2462) & (!g2542) & (g2509) & (g2546) & (!g3765) & (!g3766)) + ((!g2462) & (g2542) & (!g2509) & (!g2546) & (!g3765) & (!g3766)) + ((!g2462) & (g2542) & (!g2509) & (!g2546) & (!g3765) & (g3766)) + ((!g2462) & (g2542) & (!g2509) & (!g2546) & (g3765) & (!g3766)) + ((!g2462) & (g2542) & (!g2509) & (!g2546) & (g3765) & (g3766)) + ((!g2462) & (g2542) & (g2509) & (!g2546) & (!g3765) & (!g3766)) + ((g2462) & (!g2542) & (!g2509) & (!g2546) & (!g3765) & (!g3766)) + ((g2462) & (!g2542) & (!g2509) & (!g2546) & (!g3765) & (g3766)) + ((g2462) & (!g2542) & (!g2509) & (!g2546) & (g3765) & (!g3766)) + ((g2462) & (!g2542) & (!g2509) & (!g2546) & (g3765) & (g3766)) + ((g2462) & (!g2542) & (!g2509) & (g2546) & (!g3765) & (!g3766)) + ((g2462) & (!g2542) & (g2509) & (!g2546) & (!g3765) & (!g3766)) + ((g2462) & (!g2542) & (g2509) & (!g2546) & (!g3765) & (g3766)) + ((g2462) & (!g2542) & (g2509) & (!g2546) & (g3765) & (!g3766)) + ((g2462) & (!g2542) & (g2509) & (!g2546) & (g3765) & (g3766)) + ((g2462) & (g2542) & (!g2509) & (!g2546) & (!g3765) & (!g3766)));
	assign g3768 = (((!g2462) & (!g2509) & (!g3765) & (!g3766) & (!g5809) & (g5810)) + ((!g2462) & (!g2509) & (!g3765) & (g3766) & (!g5809) & (g5810)) + ((!g2462) & (!g2509) & (g3765) & (!g3766) & (!g5809) & (g5810)) + ((!g2462) & (!g2509) & (g3765) & (g3766) & (!g5809) & (g5810)) + ((!g2462) & (g2509) & (!g3765) & (!g3766) & (!g5809) & (g5810)) + ((!g2462) & (g2509) & (!g3765) & (g3766) & (!g5809) & (g5810)) + ((!g2462) & (g2509) & (!g3765) & (g3766) & (g5809) & (g5810)) + ((!g2462) & (g2509) & (g3765) & (!g3766) & (!g5809) & (g5810)) + ((!g2462) & (g2509) & (g3765) & (!g3766) & (g5809) & (g5810)) + ((!g2462) & (g2509) & (g3765) & (g3766) & (!g5809) & (g5810)) + ((!g2462) & (g2509) & (g3765) & (g3766) & (g5809) & (g5810)) + ((g2462) & (!g2509) & (!g3765) & (!g3766) & (!g5809) & (g5810)) + ((g2462) & (!g2509) & (!g3765) & (g3766) & (!g5809) & (g5810)) + ((g2462) & (!g2509) & (!g3765) & (g3766) & (g5809) & (g5810)) + ((g2462) & (!g2509) & (g3765) & (!g3766) & (!g5809) & (g5810)) + ((g2462) & (!g2509) & (g3765) & (!g3766) & (g5809) & (g5810)) + ((g2462) & (!g2509) & (g3765) & (g3766) & (!g5809) & (g5810)) + ((g2462) & (!g2509) & (g3765) & (g3766) & (g5809) & (g5810)) + ((g2462) & (g2509) & (!g3765) & (!g3766) & (!g5809) & (g5810)) + ((g2462) & (g2509) & (!g3765) & (!g3766) & (g5809) & (g5810)) + ((g2462) & (g2509) & (!g3765) & (g3766) & (!g5809) & (g5810)) + ((g2462) & (g2509) & (!g3765) & (g3766) & (g5809) & (g5810)) + ((g2462) & (g2509) & (g3765) & (!g3766) & (!g5809) & (g5810)) + ((g2462) & (g2509) & (g3765) & (!g3766) & (g5809) & (g5810)) + ((g2462) & (g2509) & (g3765) & (g3766) & (!g5809) & (g5810)) + ((g2462) & (g2509) & (g3765) & (g3766) & (g5809) & (g5810)));
	assign g3769 = (((g2661) & (g2676)));
	assign g3770 = (((!g2742) & (!g2772) & (!g2752) & (!g2787) & (!g3768) & (!g3769)) + ((!g2742) & (!g2772) & (!g2752) & (!g2787) & (!g3768) & (g3769)) + ((!g2742) & (!g2772) & (!g2752) & (!g2787) & (g3768) & (!g3769)) + ((!g2742) & (!g2772) & (!g2752) & (!g2787) & (g3768) & (g3769)) + ((!g2742) & (!g2772) & (!g2752) & (g2787) & (!g3768) & (!g3769)) + ((!g2742) & (!g2772) & (!g2752) & (g2787) & (!g3768) & (g3769)) + ((!g2742) & (!g2772) & (!g2752) & (g2787) & (g3768) & (!g3769)) + ((!g2742) & (!g2772) & (!g2752) & (g2787) & (g3768) & (g3769)) + ((!g2742) & (!g2772) & (g2752) & (!g2787) & (!g3768) & (!g3769)) + ((!g2742) & (!g2772) & (g2752) & (!g2787) & (!g3768) & (g3769)) + ((!g2742) & (!g2772) & (g2752) & (!g2787) & (g3768) & (!g3769)) + ((!g2742) & (!g2772) & (g2752) & (!g2787) & (g3768) & (g3769)) + ((!g2742) & (!g2772) & (g2752) & (g2787) & (!g3768) & (!g3769)) + ((!g2742) & (g2772) & (!g2752) & (!g2787) & (!g3768) & (!g3769)) + ((!g2742) & (g2772) & (!g2752) & (!g2787) & (!g3768) & (g3769)) + ((!g2742) & (g2772) & (!g2752) & (!g2787) & (g3768) & (!g3769)) + ((!g2742) & (g2772) & (!g2752) & (!g2787) & (g3768) & (g3769)) + ((!g2742) & (g2772) & (g2752) & (!g2787) & (!g3768) & (!g3769)) + ((g2742) & (!g2772) & (!g2752) & (!g2787) & (!g3768) & (!g3769)) + ((g2742) & (!g2772) & (!g2752) & (!g2787) & (!g3768) & (g3769)) + ((g2742) & (!g2772) & (!g2752) & (!g2787) & (g3768) & (!g3769)) + ((g2742) & (!g2772) & (!g2752) & (!g2787) & (g3768) & (g3769)) + ((g2742) & (!g2772) & (!g2752) & (g2787) & (!g3768) & (!g3769)) + ((g2742) & (!g2772) & (g2752) & (!g2787) & (!g3768) & (!g3769)) + ((g2742) & (!g2772) & (g2752) & (!g2787) & (!g3768) & (g3769)) + ((g2742) & (!g2772) & (g2752) & (!g2787) & (g3768) & (!g3769)) + ((g2742) & (!g2772) & (g2752) & (!g2787) & (g3768) & (g3769)) + ((g2742) & (g2772) & (!g2752) & (!g2787) & (!g3768) & (!g3769)));
	assign g3771 = (((!g2900) & (g2904)) + ((g2900) & (!g2904)));
	assign g3772 = (((!g2827) & (!g2851) & (g2833) & (g2874) & (!g3770) & (g3771)) + ((!g2827) & (g2851) & (!g2833) & (g2874) & (!g3770) & (g3771)) + ((!g2827) & (g2851) & (!g2833) & (g2874) & (g3770) & (g3771)) + ((!g2827) & (g2851) & (g2833) & (!g2874) & (!g3770) & (g3771)) + ((!g2827) & (g2851) & (g2833) & (g2874) & (!g3770) & (g3771)) + ((!g2827) & (g2851) & (g2833) & (g2874) & (g3770) & (g3771)) + ((g2827) & (!g2851) & (!g2833) & (g2874) & (!g3770) & (g3771)) + ((g2827) & (!g2851) & (g2833) & (g2874) & (!g3770) & (g3771)) + ((g2827) & (!g2851) & (g2833) & (g2874) & (g3770) & (g3771)) + ((g2827) & (g2851) & (!g2833) & (!g2874) & (!g3770) & (g3771)) + ((g2827) & (g2851) & (!g2833) & (g2874) & (!g3770) & (g3771)) + ((g2827) & (g2851) & (!g2833) & (g2874) & (g3770) & (g3771)) + ((g2827) & (g2851) & (g2833) & (!g2874) & (!g3770) & (g3771)) + ((g2827) & (g2851) & (g2833) & (!g2874) & (g3770) & (g3771)) + ((g2827) & (g2851) & (g2833) & (g2874) & (!g3770) & (g3771)) + ((g2827) & (g2851) & (g2833) & (g2874) & (g3770) & (g3771)));
	assign g3773 = (((g2900) & (g2904)));
	assign g3774 = (((!g2944) & (!g3018) & (!g2991) & (!g3022) & (!g3772) & (!g3773)) + ((!g2944) & (!g3018) & (!g2991) & (!g3022) & (!g3772) & (g3773)) + ((!g2944) & (!g3018) & (!g2991) & (!g3022) & (g3772) & (!g3773)) + ((!g2944) & (!g3018) & (!g2991) & (!g3022) & (g3772) & (g3773)) + ((!g2944) & (!g3018) & (!g2991) & (g3022) & (!g3772) & (!g3773)) + ((!g2944) & (!g3018) & (!g2991) & (g3022) & (!g3772) & (g3773)) + ((!g2944) & (!g3018) & (!g2991) & (g3022) & (g3772) & (!g3773)) + ((!g2944) & (!g3018) & (!g2991) & (g3022) & (g3772) & (g3773)) + ((!g2944) & (!g3018) & (g2991) & (!g3022) & (!g3772) & (!g3773)) + ((!g2944) & (!g3018) & (g2991) & (!g3022) & (!g3772) & (g3773)) + ((!g2944) & (!g3018) & (g2991) & (!g3022) & (g3772) & (!g3773)) + ((!g2944) & (!g3018) & (g2991) & (!g3022) & (g3772) & (g3773)) + ((!g2944) & (!g3018) & (g2991) & (g3022) & (!g3772) & (!g3773)) + ((!g2944) & (g3018) & (!g2991) & (!g3022) & (!g3772) & (!g3773)) + ((!g2944) & (g3018) & (!g2991) & (!g3022) & (!g3772) & (g3773)) + ((!g2944) & (g3018) & (!g2991) & (!g3022) & (g3772) & (!g3773)) + ((!g2944) & (g3018) & (!g2991) & (!g3022) & (g3772) & (g3773)) + ((!g2944) & (g3018) & (g2991) & (!g3022) & (!g3772) & (!g3773)) + ((g2944) & (!g3018) & (!g2991) & (!g3022) & (!g3772) & (!g3773)) + ((g2944) & (!g3018) & (!g2991) & (!g3022) & (!g3772) & (g3773)) + ((g2944) & (!g3018) & (!g2991) & (!g3022) & (g3772) & (!g3773)) + ((g2944) & (!g3018) & (!g2991) & (!g3022) & (g3772) & (g3773)) + ((g2944) & (!g3018) & (!g2991) & (g3022) & (!g3772) & (!g3773)) + ((g2944) & (!g3018) & (g2991) & (!g3022) & (!g3772) & (!g3773)) + ((g2944) & (!g3018) & (g2991) & (!g3022) & (!g3772) & (g3773)) + ((g2944) & (!g3018) & (g2991) & (!g3022) & (g3772) & (!g3773)) + ((g2944) & (!g3018) & (g2991) & (!g3022) & (g3772) & (g3773)) + ((g2944) & (g3018) & (!g2991) & (!g3022) & (!g3772) & (!g3773)));
	assign g3775 = (((!g3044) & (g3067) & (!g3774)) + ((g3044) & (!g3067) & (!g3774)) + ((g3044) & (g3067) & (!g3774)) + ((g3044) & (g3067) & (g3774)));
	assign g3776 = (((!g3097) & (g3775) & (g3093)) + ((g3097) & (!g3775) & (g3093)) + ((g3097) & (g3775) & (!g3093)) + ((g3097) & (g3775) & (g3093)));
	assign g3777 = (((!g830) & (!g1906) & (!g6999) & (key[64])) + ((!g830) & (!g1906) & (g6999) & (key[64])) + ((!g830) & (g1906) & (!g6999) & (key[64])) + ((!g830) & (g1906) & (g6999) & (key[64])) + ((g830) & (!g1906) & (g6999) & (!key[64])) + ((g830) & (!g1906) & (g6999) & (key[64])) + ((g830) & (g1906) & (!g6999) & (!key[64])) + ((g830) & (g1906) & (!g6999) & (key[64])));
	assign g3778 = (((!g1892) & (!g2026) & (g2062) & (!g1900) & (!g2028) & (g2074)) + ((!g1892) & (!g2026) & (g2062) & (!g1900) & (g2028) & (g2074)) + ((!g1892) & (!g2026) & (g2062) & (g1900) & (!g2028) & (g2074)) + ((!g1892) & (!g2026) & (g2062) & (g1900) & (g2028) & (g2074)) + ((!g1892) & (g2026) & (!g2062) & (!g1900) & (g2028) & (g2074)) + ((!g1892) & (g2026) & (!g2062) & (g1900) & (g2028) & (g2074)) + ((!g1892) & (g2026) & (g2062) & (!g1900) & (!g2028) & (g2074)) + ((!g1892) & (g2026) & (g2062) & (!g1900) & (g2028) & (!g2074)) + ((!g1892) & (g2026) & (g2062) & (!g1900) & (g2028) & (g2074)) + ((!g1892) & (g2026) & (g2062) & (g1900) & (!g2028) & (g2074)) + ((!g1892) & (g2026) & (g2062) & (g1900) & (g2028) & (!g2074)) + ((!g1892) & (g2026) & (g2062) & (g1900) & (g2028) & (g2074)) + ((g1892) & (!g2026) & (!g2062) & (g1900) & (g2028) & (g2074)) + ((g1892) & (!g2026) & (g2062) & (!g1900) & (!g2028) & (g2074)) + ((g1892) & (!g2026) & (g2062) & (!g1900) & (g2028) & (g2074)) + ((g1892) & (!g2026) & (g2062) & (g1900) & (!g2028) & (g2074)) + ((g1892) & (!g2026) & (g2062) & (g1900) & (g2028) & (!g2074)) + ((g1892) & (!g2026) & (g2062) & (g1900) & (g2028) & (g2074)) + ((g1892) & (g2026) & (!g2062) & (!g1900) & (g2028) & (g2074)) + ((g1892) & (g2026) & (!g2062) & (g1900) & (!g2028) & (g2074)) + ((g1892) & (g2026) & (!g2062) & (g1900) & (g2028) & (g2074)) + ((g1892) & (g2026) & (g2062) & (!g1900) & (!g2028) & (g2074)) + ((g1892) & (g2026) & (g2062) & (!g1900) & (g2028) & (!g2074)) + ((g1892) & (g2026) & (g2062) & (!g1900) & (g2028) & (g2074)) + ((g1892) & (g2026) & (g2062) & (g1900) & (!g2028) & (!g2074)) + ((g1892) & (g2026) & (g2062) & (g1900) & (!g2028) & (g2074)) + ((g1892) & (g2026) & (g2062) & (g1900) & (g2028) & (!g2074)) + ((g1892) & (g2026) & (g2062) & (g1900) & (g2028) & (g2074)));
	assign g3779 = (((!g2188) & (g2190)) + ((g2188) & (!g2190)));
	assign g3780 = (((!g2108) & (!g2144) & (g2110) & (g2156) & (g3778) & (g3779)) + ((!g2108) & (g2144) & (!g2110) & (g2156) & (!g3778) & (g3779)) + ((!g2108) & (g2144) & (!g2110) & (g2156) & (g3778) & (g3779)) + ((!g2108) & (g2144) & (g2110) & (!g2156) & (g3778) & (g3779)) + ((!g2108) & (g2144) & (g2110) & (g2156) & (!g3778) & (g3779)) + ((!g2108) & (g2144) & (g2110) & (g2156) & (g3778) & (g3779)) + ((g2108) & (!g2144) & (!g2110) & (g2156) & (g3778) & (g3779)) + ((g2108) & (!g2144) & (g2110) & (g2156) & (!g3778) & (g3779)) + ((g2108) & (!g2144) & (g2110) & (g2156) & (g3778) & (g3779)) + ((g2108) & (g2144) & (!g2110) & (!g2156) & (g3778) & (g3779)) + ((g2108) & (g2144) & (!g2110) & (g2156) & (!g3778) & (g3779)) + ((g2108) & (g2144) & (!g2110) & (g2156) & (g3778) & (g3779)) + ((g2108) & (g2144) & (g2110) & (!g2156) & (!g3778) & (g3779)) + ((g2108) & (g2144) & (g2110) & (!g2156) & (g3778) & (g3779)) + ((g2108) & (g2144) & (g2110) & (g2156) & (!g3778) & (g3779)) + ((g2108) & (g2144) & (g2110) & (g2156) & (g3778) & (g3779)));
	assign g3781 = (((g2188) & (g2190)));
	assign g3782 = (((!g2224) & (!g2271) & (!g2236) & (!g2273) & (!g3780) & (!g3781)) + ((!g2224) & (!g2271) & (!g2236) & (!g2273) & (!g3780) & (g3781)) + ((!g2224) & (!g2271) & (!g2236) & (!g2273) & (g3780) & (!g3781)) + ((!g2224) & (!g2271) & (!g2236) & (!g2273) & (g3780) & (g3781)) + ((!g2224) & (!g2271) & (!g2236) & (g2273) & (!g3780) & (!g3781)) + ((!g2224) & (!g2271) & (!g2236) & (g2273) & (!g3780) & (g3781)) + ((!g2224) & (!g2271) & (!g2236) & (g2273) & (g3780) & (!g3781)) + ((!g2224) & (!g2271) & (!g2236) & (g2273) & (g3780) & (g3781)) + ((!g2224) & (!g2271) & (g2236) & (!g2273) & (!g3780) & (!g3781)) + ((!g2224) & (!g2271) & (g2236) & (!g2273) & (!g3780) & (g3781)) + ((!g2224) & (!g2271) & (g2236) & (!g2273) & (g3780) & (!g3781)) + ((!g2224) & (!g2271) & (g2236) & (!g2273) & (g3780) & (g3781)) + ((!g2224) & (!g2271) & (g2236) & (g2273) & (!g3780) & (!g3781)) + ((!g2224) & (g2271) & (!g2236) & (!g2273) & (!g3780) & (!g3781)) + ((!g2224) & (g2271) & (!g2236) & (!g2273) & (!g3780) & (g3781)) + ((!g2224) & (g2271) & (!g2236) & (!g2273) & (g3780) & (!g3781)) + ((!g2224) & (g2271) & (!g2236) & (!g2273) & (g3780) & (g3781)) + ((!g2224) & (g2271) & (g2236) & (!g2273) & (!g3780) & (!g3781)) + ((g2224) & (!g2271) & (!g2236) & (!g2273) & (!g3780) & (!g3781)) + ((g2224) & (!g2271) & (!g2236) & (!g2273) & (!g3780) & (g3781)) + ((g2224) & (!g2271) & (!g2236) & (!g2273) & (g3780) & (!g3781)) + ((g2224) & (!g2271) & (!g2236) & (!g2273) & (g3780) & (g3781)) + ((g2224) & (!g2271) & (!g2236) & (g2273) & (!g3780) & (!g3781)) + ((g2224) & (!g2271) & (g2236) & (!g2273) & (!g3780) & (!g3781)) + ((g2224) & (!g2271) & (g2236) & (!g2273) & (!g3780) & (g3781)) + ((g2224) & (!g2271) & (g2236) & (!g2273) & (g3780) & (!g3781)) + ((g2224) & (!g2271) & (g2236) & (!g2273) & (g3780) & (g3781)) + ((g2224) & (g2271) & (!g2236) & (!g2273) & (!g3780) & (!g3781)));
	assign g3783 = (((!g2390) & (g2402)) + ((g2390) & (!g2402)));
	assign g3784 = (((!g2311) & (!g2354) & (g2323) & (g2356) & (!g3782) & (g3783)) + ((!g2311) & (g2354) & (!g2323) & (g2356) & (!g3782) & (g3783)) + ((!g2311) & (g2354) & (!g2323) & (g2356) & (g3782) & (g3783)) + ((!g2311) & (g2354) & (g2323) & (!g2356) & (!g3782) & (g3783)) + ((!g2311) & (g2354) & (g2323) & (g2356) & (!g3782) & (g3783)) + ((!g2311) & (g2354) & (g2323) & (g2356) & (g3782) & (g3783)) + ((g2311) & (!g2354) & (!g2323) & (g2356) & (!g3782) & (g3783)) + ((g2311) & (!g2354) & (g2323) & (g2356) & (!g3782) & (g3783)) + ((g2311) & (!g2354) & (g2323) & (g2356) & (g3782) & (g3783)) + ((g2311) & (g2354) & (!g2323) & (!g2356) & (!g3782) & (g3783)) + ((g2311) & (g2354) & (!g2323) & (g2356) & (!g3782) & (g3783)) + ((g2311) & (g2354) & (!g2323) & (g2356) & (g3782) & (g3783)) + ((g2311) & (g2354) & (g2323) & (!g2356) & (!g3782) & (g3783)) + ((g2311) & (g2354) & (g2323) & (!g2356) & (g3782) & (g3783)) + ((g2311) & (g2354) & (g2323) & (g2356) & (!g3782) & (g3783)) + ((g2311) & (g2354) & (g2323) & (g2356) & (g3782) & (g3783)));
	assign g3785 = (((g2390) & (g2402)));
	assign g3786 = (((!g2450) & (!g2527) & (!g2456) & (!g2535) & (!g3784) & (!g3785)) + ((!g2450) & (!g2527) & (!g2456) & (!g2535) & (!g3784) & (g3785)) + ((!g2450) & (!g2527) & (!g2456) & (!g2535) & (g3784) & (!g3785)) + ((!g2450) & (!g2527) & (!g2456) & (!g2535) & (g3784) & (g3785)) + ((!g2450) & (!g2527) & (!g2456) & (g2535) & (!g3784) & (!g3785)) + ((!g2450) & (!g2527) & (!g2456) & (g2535) & (!g3784) & (g3785)) + ((!g2450) & (!g2527) & (!g2456) & (g2535) & (g3784) & (!g3785)) + ((!g2450) & (!g2527) & (!g2456) & (g2535) & (g3784) & (g3785)) + ((!g2450) & (!g2527) & (g2456) & (!g2535) & (!g3784) & (!g3785)) + ((!g2450) & (!g2527) & (g2456) & (!g2535) & (!g3784) & (g3785)) + ((!g2450) & (!g2527) & (g2456) & (!g2535) & (g3784) & (!g3785)) + ((!g2450) & (!g2527) & (g2456) & (!g2535) & (g3784) & (g3785)) + ((!g2450) & (!g2527) & (g2456) & (g2535) & (!g3784) & (!g3785)) + ((!g2450) & (g2527) & (!g2456) & (!g2535) & (!g3784) & (!g3785)) + ((!g2450) & (g2527) & (!g2456) & (!g2535) & (!g3784) & (g3785)) + ((!g2450) & (g2527) & (!g2456) & (!g2535) & (g3784) & (!g3785)) + ((!g2450) & (g2527) & (!g2456) & (!g2535) & (g3784) & (g3785)) + ((!g2450) & (g2527) & (g2456) & (!g2535) & (!g3784) & (!g3785)) + ((g2450) & (!g2527) & (!g2456) & (!g2535) & (!g3784) & (!g3785)) + ((g2450) & (!g2527) & (!g2456) & (!g2535) & (!g3784) & (g3785)) + ((g2450) & (!g2527) & (!g2456) & (!g2535) & (g3784) & (!g3785)) + ((g2450) & (!g2527) & (!g2456) & (!g2535) & (g3784) & (g3785)) + ((g2450) & (!g2527) & (!g2456) & (g2535) & (!g3784) & (!g3785)) + ((g2450) & (!g2527) & (g2456) & (!g2535) & (!g3784) & (!g3785)) + ((g2450) & (!g2527) & (g2456) & (!g2535) & (!g3784) & (g3785)) + ((g2450) & (!g2527) & (g2456) & (!g2535) & (g3784) & (!g3785)) + ((g2450) & (!g2527) & (g2456) & (!g2535) & (g3784) & (g3785)) + ((g2450) & (g2527) & (!g2456) & (!g2535) & (!g3784) & (!g3785)));
	assign g3787 = (((!g2450) & (!g2456) & (!g3784) & (!g3785) & (!g5812) & (g5813)) + ((!g2450) & (!g2456) & (!g3784) & (g3785) & (!g5812) & (g5813)) + ((!g2450) & (!g2456) & (g3784) & (!g3785) & (!g5812) & (g5813)) + ((!g2450) & (!g2456) & (g3784) & (g3785) & (!g5812) & (g5813)) + ((!g2450) & (g2456) & (!g3784) & (!g3785) & (!g5812) & (g5813)) + ((!g2450) & (g2456) & (!g3784) & (g3785) & (!g5812) & (g5813)) + ((!g2450) & (g2456) & (!g3784) & (g3785) & (g5812) & (g5813)) + ((!g2450) & (g2456) & (g3784) & (!g3785) & (!g5812) & (g5813)) + ((!g2450) & (g2456) & (g3784) & (!g3785) & (g5812) & (g5813)) + ((!g2450) & (g2456) & (g3784) & (g3785) & (!g5812) & (g5813)) + ((!g2450) & (g2456) & (g3784) & (g3785) & (g5812) & (g5813)) + ((g2450) & (!g2456) & (!g3784) & (!g3785) & (!g5812) & (g5813)) + ((g2450) & (!g2456) & (!g3784) & (g3785) & (!g5812) & (g5813)) + ((g2450) & (!g2456) & (!g3784) & (g3785) & (g5812) & (g5813)) + ((g2450) & (!g2456) & (g3784) & (!g3785) & (!g5812) & (g5813)) + ((g2450) & (!g2456) & (g3784) & (!g3785) & (g5812) & (g5813)) + ((g2450) & (!g2456) & (g3784) & (g3785) & (!g5812) & (g5813)) + ((g2450) & (!g2456) & (g3784) & (g3785) & (g5812) & (g5813)) + ((g2450) & (g2456) & (!g3784) & (!g3785) & (!g5812) & (g5813)) + ((g2450) & (g2456) & (!g3784) & (!g3785) & (g5812) & (g5813)) + ((g2450) & (g2456) & (!g3784) & (g3785) & (!g5812) & (g5813)) + ((g2450) & (g2456) & (!g3784) & (g3785) & (g5812) & (g5813)) + ((g2450) & (g2456) & (g3784) & (!g3785) & (!g5812) & (g5813)) + ((g2450) & (g2456) & (g3784) & (!g3785) & (g5812) & (g5813)) + ((g2450) & (g2456) & (g3784) & (g3785) & (!g5812) & (g5813)) + ((g2450) & (g2456) & (g3784) & (g3785) & (g5812) & (g5813)));
	assign g3788 = (((g2657) & (g2659)));
	assign g3789 = (((!g2703) & (!g2768) & (!g2723) & (!g2770) & (!g3787) & (!g3788)) + ((!g2703) & (!g2768) & (!g2723) & (!g2770) & (!g3787) & (g3788)) + ((!g2703) & (!g2768) & (!g2723) & (!g2770) & (g3787) & (!g3788)) + ((!g2703) & (!g2768) & (!g2723) & (!g2770) & (g3787) & (g3788)) + ((!g2703) & (!g2768) & (!g2723) & (g2770) & (!g3787) & (!g3788)) + ((!g2703) & (!g2768) & (!g2723) & (g2770) & (!g3787) & (g3788)) + ((!g2703) & (!g2768) & (!g2723) & (g2770) & (g3787) & (!g3788)) + ((!g2703) & (!g2768) & (!g2723) & (g2770) & (g3787) & (g3788)) + ((!g2703) & (!g2768) & (g2723) & (!g2770) & (!g3787) & (!g3788)) + ((!g2703) & (!g2768) & (g2723) & (!g2770) & (!g3787) & (g3788)) + ((!g2703) & (!g2768) & (g2723) & (!g2770) & (g3787) & (!g3788)) + ((!g2703) & (!g2768) & (g2723) & (!g2770) & (g3787) & (g3788)) + ((!g2703) & (!g2768) & (g2723) & (g2770) & (!g3787) & (!g3788)) + ((!g2703) & (g2768) & (!g2723) & (!g2770) & (!g3787) & (!g3788)) + ((!g2703) & (g2768) & (!g2723) & (!g2770) & (!g3787) & (g3788)) + ((!g2703) & (g2768) & (!g2723) & (!g2770) & (g3787) & (!g3788)) + ((!g2703) & (g2768) & (!g2723) & (!g2770) & (g3787) & (g3788)) + ((!g2703) & (g2768) & (g2723) & (!g2770) & (!g3787) & (!g3788)) + ((g2703) & (!g2768) & (!g2723) & (!g2770) & (!g3787) & (!g3788)) + ((g2703) & (!g2768) & (!g2723) & (!g2770) & (!g3787) & (g3788)) + ((g2703) & (!g2768) & (!g2723) & (!g2770) & (g3787) & (!g3788)) + ((g2703) & (!g2768) & (!g2723) & (!g2770) & (g3787) & (g3788)) + ((g2703) & (!g2768) & (!g2723) & (g2770) & (!g3787) & (!g3788)) + ((g2703) & (!g2768) & (g2723) & (!g2770) & (!g3787) & (!g3788)) + ((g2703) & (!g2768) & (g2723) & (!g2770) & (!g3787) & (g3788)) + ((g2703) & (!g2768) & (g2723) & (!g2770) & (g3787) & (!g3788)) + ((g2703) & (!g2768) & (g2723) & (!g2770) & (g3787) & (g3788)) + ((g2703) & (g2768) & (!g2723) & (!g2770) & (!g3787) & (!g3788)));
	assign g3790 = (((!g2885) & (g2893)) + ((g2885) & (!g2893)));
	assign g3791 = (((!g2804) & (!g2845) & (g2816) & (g2848) & (!g3789) & (g3790)) + ((!g2804) & (g2845) & (!g2816) & (g2848) & (!g3789) & (g3790)) + ((!g2804) & (g2845) & (!g2816) & (g2848) & (g3789) & (g3790)) + ((!g2804) & (g2845) & (g2816) & (!g2848) & (!g3789) & (g3790)) + ((!g2804) & (g2845) & (g2816) & (g2848) & (!g3789) & (g3790)) + ((!g2804) & (g2845) & (g2816) & (g2848) & (g3789) & (g3790)) + ((g2804) & (!g2845) & (!g2816) & (g2848) & (!g3789) & (g3790)) + ((g2804) & (!g2845) & (g2816) & (g2848) & (!g3789) & (g3790)) + ((g2804) & (!g2845) & (g2816) & (g2848) & (g3789) & (g3790)) + ((g2804) & (g2845) & (!g2816) & (!g2848) & (!g3789) & (g3790)) + ((g2804) & (g2845) & (!g2816) & (g2848) & (!g3789) & (g3790)) + ((g2804) & (g2845) & (!g2816) & (g2848) & (g3789) & (g3790)) + ((g2804) & (g2845) & (g2816) & (!g2848) & (!g3789) & (g3790)) + ((g2804) & (g2845) & (g2816) & (!g2848) & (g3789) & (g3790)) + ((g2804) & (g2845) & (g2816) & (g2848) & (!g3789) & (g3790)) + ((g2804) & (g2845) & (g2816) & (g2848) & (g3789) & (g3790)));
	assign g3792 = (((g2885) & (g2893)));
	assign g3793 = (((!g2932) & (!g3003) & (!g2938) & (!g3011) & (!g3791) & (!g3792)) + ((!g2932) & (!g3003) & (!g2938) & (!g3011) & (!g3791) & (g3792)) + ((!g2932) & (!g3003) & (!g2938) & (!g3011) & (g3791) & (!g3792)) + ((!g2932) & (!g3003) & (!g2938) & (!g3011) & (g3791) & (g3792)) + ((!g2932) & (!g3003) & (!g2938) & (g3011) & (!g3791) & (!g3792)) + ((!g2932) & (!g3003) & (!g2938) & (g3011) & (!g3791) & (g3792)) + ((!g2932) & (!g3003) & (!g2938) & (g3011) & (g3791) & (!g3792)) + ((!g2932) & (!g3003) & (!g2938) & (g3011) & (g3791) & (g3792)) + ((!g2932) & (!g3003) & (g2938) & (!g3011) & (!g3791) & (!g3792)) + ((!g2932) & (!g3003) & (g2938) & (!g3011) & (!g3791) & (g3792)) + ((!g2932) & (!g3003) & (g2938) & (!g3011) & (g3791) & (!g3792)) + ((!g2932) & (!g3003) & (g2938) & (!g3011) & (g3791) & (g3792)) + ((!g2932) & (!g3003) & (g2938) & (g3011) & (!g3791) & (!g3792)) + ((!g2932) & (g3003) & (!g2938) & (!g3011) & (!g3791) & (!g3792)) + ((!g2932) & (g3003) & (!g2938) & (!g3011) & (!g3791) & (g3792)) + ((!g2932) & (g3003) & (!g2938) & (!g3011) & (g3791) & (!g3792)) + ((!g2932) & (g3003) & (!g2938) & (!g3011) & (g3791) & (g3792)) + ((!g2932) & (g3003) & (g2938) & (!g3011) & (!g3791) & (!g3792)) + ((g2932) & (!g3003) & (!g2938) & (!g3011) & (!g3791) & (!g3792)) + ((g2932) & (!g3003) & (!g2938) & (!g3011) & (!g3791) & (g3792)) + ((g2932) & (!g3003) & (!g2938) & (!g3011) & (g3791) & (!g3792)) + ((g2932) & (!g3003) & (!g2938) & (!g3011) & (g3791) & (g3792)) + ((g2932) & (!g3003) & (!g2938) & (g3011) & (!g3791) & (!g3792)) + ((g2932) & (!g3003) & (g2938) & (!g3011) & (!g3791) & (!g3792)) + ((g2932) & (!g3003) & (g2938) & (!g3011) & (!g3791) & (g3792)) + ((g2932) & (!g3003) & (g2938) & (!g3011) & (g3791) & (!g3792)) + ((g2932) & (!g3003) & (g2938) & (!g3011) & (g3791) & (g3792)) + ((g2932) & (g3003) & (!g2938) & (!g3011) & (!g3791) & (!g3792)));
	assign g3794 = (((!g3038) & (g3041) & (!g3793)) + ((g3038) & (!g3041) & (!g3793)) + ((g3038) & (g3041) & (!g3793)) + ((g3038) & (g3041) & (g3793)));
	assign g3795 = (((!g1906) & (!g1940) & (g1942) & (!g1910) & (!g2038) & (g2088)) + ((!g1906) & (!g1940) & (g1942) & (!g1910) & (g2038) & (g2088)) + ((!g1906) & (!g1940) & (g1942) & (g1910) & (!g2038) & (g2088)) + ((!g1906) & (!g1940) & (g1942) & (g1910) & (g2038) & (g2088)) + ((!g1906) & (g1940) & (!g1942) & (!g1910) & (g2038) & (g2088)) + ((!g1906) & (g1940) & (!g1942) & (g1910) & (g2038) & (g2088)) + ((!g1906) & (g1940) & (g1942) & (!g1910) & (!g2038) & (g2088)) + ((!g1906) & (g1940) & (g1942) & (!g1910) & (g2038) & (!g2088)) + ((!g1906) & (g1940) & (g1942) & (!g1910) & (g2038) & (g2088)) + ((!g1906) & (g1940) & (g1942) & (g1910) & (!g2038) & (g2088)) + ((!g1906) & (g1940) & (g1942) & (g1910) & (g2038) & (!g2088)) + ((!g1906) & (g1940) & (g1942) & (g1910) & (g2038) & (g2088)) + ((g1906) & (!g1940) & (!g1942) & (g1910) & (g2038) & (g2088)) + ((g1906) & (!g1940) & (g1942) & (!g1910) & (!g2038) & (g2088)) + ((g1906) & (!g1940) & (g1942) & (!g1910) & (g2038) & (g2088)) + ((g1906) & (!g1940) & (g1942) & (g1910) & (!g2038) & (g2088)) + ((g1906) & (!g1940) & (g1942) & (g1910) & (g2038) & (!g2088)) + ((g1906) & (!g1940) & (g1942) & (g1910) & (g2038) & (g2088)) + ((g1906) & (g1940) & (!g1942) & (!g1910) & (g2038) & (g2088)) + ((g1906) & (g1940) & (!g1942) & (g1910) & (!g2038) & (g2088)) + ((g1906) & (g1940) & (!g1942) & (g1910) & (g2038) & (g2088)) + ((g1906) & (g1940) & (g1942) & (!g1910) & (!g2038) & (g2088)) + ((g1906) & (g1940) & (g1942) & (!g1910) & (g2038) & (!g2088)) + ((g1906) & (g1940) & (g1942) & (!g1910) & (g2038) & (g2088)) + ((g1906) & (g1940) & (g1942) & (g1910) & (!g2038) & (!g2088)) + ((g1906) & (g1940) & (g1942) & (g1910) & (!g2038) & (g2088)) + ((g1906) & (g1940) & (g1942) & (g1910) & (g2038) & (!g2088)) + ((g1906) & (g1940) & (g1942) & (g1910) & (g2038) & (g2088)));
	assign g3796 = (((!g1949) & (g2200)) + ((g1949) & (!g2200)));
	assign g3797 = (((!g1945) & (!g1947) & (g2120) & (g2170) & (g3795) & (g3796)) + ((!g1945) & (g1947) & (!g2120) & (g2170) & (!g3795) & (g3796)) + ((!g1945) & (g1947) & (!g2120) & (g2170) & (g3795) & (g3796)) + ((!g1945) & (g1947) & (g2120) & (!g2170) & (g3795) & (g3796)) + ((!g1945) & (g1947) & (g2120) & (g2170) & (!g3795) & (g3796)) + ((!g1945) & (g1947) & (g2120) & (g2170) & (g3795) & (g3796)) + ((g1945) & (!g1947) & (!g2120) & (g2170) & (g3795) & (g3796)) + ((g1945) & (!g1947) & (g2120) & (g2170) & (!g3795) & (g3796)) + ((g1945) & (!g1947) & (g2120) & (g2170) & (g3795) & (g3796)) + ((g1945) & (g1947) & (!g2120) & (!g2170) & (g3795) & (g3796)) + ((g1945) & (g1947) & (!g2120) & (g2170) & (!g3795) & (g3796)) + ((g1945) & (g1947) & (!g2120) & (g2170) & (g3795) & (g3796)) + ((g1945) & (g1947) & (g2120) & (!g2170) & (!g3795) & (g3796)) + ((g1945) & (g1947) & (g2120) & (!g2170) & (g3795) & (g3796)) + ((g1945) & (g1947) & (g2120) & (g2170) & (!g3795) & (g3796)) + ((g1945) & (g1947) & (g2120) & (g2170) & (g3795) & (g3796)));
	assign g3798 = (((g1949) & (g2200)));
	assign g3799 = (((!g1954) & (!g1956) & (!g2250) & (!g2283) & (!g3797) & (!g3798)) + ((!g1954) & (!g1956) & (!g2250) & (!g2283) & (!g3797) & (g3798)) + ((!g1954) & (!g1956) & (!g2250) & (!g2283) & (g3797) & (!g3798)) + ((!g1954) & (!g1956) & (!g2250) & (!g2283) & (g3797) & (g3798)) + ((!g1954) & (!g1956) & (!g2250) & (g2283) & (!g3797) & (!g3798)) + ((!g1954) & (!g1956) & (!g2250) & (g2283) & (!g3797) & (g3798)) + ((!g1954) & (!g1956) & (!g2250) & (g2283) & (g3797) & (!g3798)) + ((!g1954) & (!g1956) & (!g2250) & (g2283) & (g3797) & (g3798)) + ((!g1954) & (!g1956) & (g2250) & (!g2283) & (!g3797) & (!g3798)) + ((!g1954) & (!g1956) & (g2250) & (!g2283) & (!g3797) & (g3798)) + ((!g1954) & (!g1956) & (g2250) & (!g2283) & (g3797) & (!g3798)) + ((!g1954) & (!g1956) & (g2250) & (!g2283) & (g3797) & (g3798)) + ((!g1954) & (!g1956) & (g2250) & (g2283) & (!g3797) & (!g3798)) + ((!g1954) & (g1956) & (!g2250) & (!g2283) & (!g3797) & (!g3798)) + ((!g1954) & (g1956) & (!g2250) & (!g2283) & (!g3797) & (g3798)) + ((!g1954) & (g1956) & (!g2250) & (!g2283) & (g3797) & (!g3798)) + ((!g1954) & (g1956) & (!g2250) & (!g2283) & (g3797) & (g3798)) + ((!g1954) & (g1956) & (g2250) & (!g2283) & (!g3797) & (!g3798)) + ((g1954) & (!g1956) & (!g2250) & (!g2283) & (!g3797) & (!g3798)) + ((g1954) & (!g1956) & (!g2250) & (!g2283) & (!g3797) & (g3798)) + ((g1954) & (!g1956) & (!g2250) & (!g2283) & (g3797) & (!g3798)) + ((g1954) & (!g1956) & (!g2250) & (!g2283) & (g3797) & (g3798)) + ((g1954) & (!g1956) & (!g2250) & (g2283) & (!g3797) & (!g3798)) + ((g1954) & (!g1956) & (g2250) & (!g2283) & (!g3797) & (!g3798)) + ((g1954) & (!g1956) & (g2250) & (!g2283) & (!g3797) & (g3798)) + ((g1954) & (!g1956) & (g2250) & (!g2283) & (g3797) & (!g3798)) + ((g1954) & (!g1956) & (g2250) & (!g2283) & (g3797) & (g3798)) + ((g1954) & (g1956) & (!g2250) & (!g2283) & (!g3797) & (!g3798)));
	assign g3800 = (((!g1963) & (g2416)) + ((g1963) & (!g2416)));
	assign g3801 = (((!g1959) & (!g1961) & (g2337) & (g2366) & (!g3799) & (g3800)) + ((!g1959) & (g1961) & (!g2337) & (g2366) & (!g3799) & (g3800)) + ((!g1959) & (g1961) & (!g2337) & (g2366) & (g3799) & (g3800)) + ((!g1959) & (g1961) & (g2337) & (!g2366) & (!g3799) & (g3800)) + ((!g1959) & (g1961) & (g2337) & (g2366) & (!g3799) & (g3800)) + ((!g1959) & (g1961) & (g2337) & (g2366) & (g3799) & (g3800)) + ((g1959) & (!g1961) & (!g2337) & (g2366) & (!g3799) & (g3800)) + ((g1959) & (!g1961) & (g2337) & (g2366) & (!g3799) & (g3800)) + ((g1959) & (!g1961) & (g2337) & (g2366) & (g3799) & (g3800)) + ((g1959) & (g1961) & (!g2337) & (!g2366) & (!g3799) & (g3800)) + ((g1959) & (g1961) & (!g2337) & (g2366) & (!g3799) & (g3800)) + ((g1959) & (g1961) & (!g2337) & (g2366) & (g3799) & (g3800)) + ((g1959) & (g1961) & (g2337) & (!g2366) & (!g3799) & (g3800)) + ((g1959) & (g1961) & (g2337) & (!g2366) & (g3799) & (g3800)) + ((g1959) & (g1961) & (g2337) & (g2366) & (!g3799) & (g3800)) + ((g1959) & (g1961) & (g2337) & (g2366) & (g3799) & (g3800)));
	assign g3802 = (((g1963) & (g2416)));
	assign g3803 = (((!g1968) & (!g1970) & (!g2486) & (!g2544) & (!g3801) & (!g3802)) + ((!g1968) & (!g1970) & (!g2486) & (!g2544) & (!g3801) & (g3802)) + ((!g1968) & (!g1970) & (!g2486) & (!g2544) & (g3801) & (!g3802)) + ((!g1968) & (!g1970) & (!g2486) & (!g2544) & (g3801) & (g3802)) + ((!g1968) & (!g1970) & (!g2486) & (g2544) & (!g3801) & (!g3802)) + ((!g1968) & (!g1970) & (!g2486) & (g2544) & (!g3801) & (g3802)) + ((!g1968) & (!g1970) & (!g2486) & (g2544) & (g3801) & (!g3802)) + ((!g1968) & (!g1970) & (!g2486) & (g2544) & (g3801) & (g3802)) + ((!g1968) & (!g1970) & (g2486) & (!g2544) & (!g3801) & (!g3802)) + ((!g1968) & (!g1970) & (g2486) & (!g2544) & (!g3801) & (g3802)) + ((!g1968) & (!g1970) & (g2486) & (!g2544) & (g3801) & (!g3802)) + ((!g1968) & (!g1970) & (g2486) & (!g2544) & (g3801) & (g3802)) + ((!g1968) & (!g1970) & (g2486) & (g2544) & (!g3801) & (!g3802)) + ((!g1968) & (g1970) & (!g2486) & (!g2544) & (!g3801) & (!g3802)) + ((!g1968) & (g1970) & (!g2486) & (!g2544) & (!g3801) & (g3802)) + ((!g1968) & (g1970) & (!g2486) & (!g2544) & (g3801) & (!g3802)) + ((!g1968) & (g1970) & (!g2486) & (!g2544) & (g3801) & (g3802)) + ((!g1968) & (g1970) & (g2486) & (!g2544) & (!g3801) & (!g3802)) + ((g1968) & (!g1970) & (!g2486) & (!g2544) & (!g3801) & (!g3802)) + ((g1968) & (!g1970) & (!g2486) & (!g2544) & (!g3801) & (g3802)) + ((g1968) & (!g1970) & (!g2486) & (!g2544) & (g3801) & (!g3802)) + ((g1968) & (!g1970) & (!g2486) & (!g2544) & (g3801) & (g3802)) + ((g1968) & (!g1970) & (!g2486) & (g2544) & (!g3801) & (!g3802)) + ((g1968) & (!g1970) & (g2486) & (!g2544) & (!g3801) & (!g3802)) + ((g1968) & (!g1970) & (g2486) & (!g2544) & (!g3801) & (g3802)) + ((g1968) & (!g1970) & (g2486) & (!g2544) & (g3801) & (!g3802)) + ((g1968) & (!g1970) & (g2486) & (!g2544) & (g3801) & (g3802)) + ((g1968) & (g1970) & (!g2486) & (!g2544) & (!g3801) & (!g3802)));
	assign g3804 = (((!g2048) & (g2669)) + ((g2048) & (!g2669)));
	assign g3805 = (((!g1973) & (!g1976) & (g2584) & (g2640) & (!g3803) & (g3804)) + ((!g1973) & (g1976) & (!g2584) & (g2640) & (!g3803) & (g3804)) + ((!g1973) & (g1976) & (!g2584) & (g2640) & (g3803) & (g3804)) + ((!g1973) & (g1976) & (g2584) & (!g2640) & (!g3803) & (g3804)) + ((!g1973) & (g1976) & (g2584) & (g2640) & (!g3803) & (g3804)) + ((!g1973) & (g1976) & (g2584) & (g2640) & (g3803) & (g3804)) + ((g1973) & (!g1976) & (!g2584) & (g2640) & (!g3803) & (g3804)) + ((g1973) & (!g1976) & (g2584) & (g2640) & (!g3803) & (g3804)) + ((g1973) & (!g1976) & (g2584) & (g2640) & (g3803) & (g3804)) + ((g1973) & (g1976) & (!g2584) & (!g2640) & (!g3803) & (g3804)) + ((g1973) & (g1976) & (!g2584) & (g2640) & (!g3803) & (g3804)) + ((g1973) & (g1976) & (!g2584) & (g2640) & (g3803) & (g3804)) + ((g1973) & (g1976) & (g2584) & (!g2640) & (!g3803) & (g3804)) + ((g1973) & (g1976) & (g2584) & (!g2640) & (g3803) & (g3804)) + ((g1973) & (g1976) & (g2584) & (g2640) & (!g3803) & (g3804)) + ((g1973) & (g1976) & (g2584) & (g2640) & (g3803) & (g3804)));
	assign g3806 = (((g2048) & (g2669)));
	assign g3807 = (((!g2099) & (!g2130) & (!g2747) & (!g2780) & (!g3805) & (!g3806)) + ((!g2099) & (!g2130) & (!g2747) & (!g2780) & (!g3805) & (g3806)) + ((!g2099) & (!g2130) & (!g2747) & (!g2780) & (g3805) & (!g3806)) + ((!g2099) & (!g2130) & (!g2747) & (!g2780) & (g3805) & (g3806)) + ((!g2099) & (!g2130) & (!g2747) & (g2780) & (!g3805) & (!g3806)) + ((!g2099) & (!g2130) & (!g2747) & (g2780) & (!g3805) & (g3806)) + ((!g2099) & (!g2130) & (!g2747) & (g2780) & (g3805) & (!g3806)) + ((!g2099) & (!g2130) & (!g2747) & (g2780) & (g3805) & (g3806)) + ((!g2099) & (!g2130) & (g2747) & (!g2780) & (!g3805) & (!g3806)) + ((!g2099) & (!g2130) & (g2747) & (!g2780) & (!g3805) & (g3806)) + ((!g2099) & (!g2130) & (g2747) & (!g2780) & (g3805) & (!g3806)) + ((!g2099) & (!g2130) & (g2747) & (!g2780) & (g3805) & (g3806)) + ((!g2099) & (!g2130) & (g2747) & (g2780) & (!g3805) & (!g3806)) + ((!g2099) & (g2130) & (!g2747) & (!g2780) & (!g3805) & (!g3806)) + ((!g2099) & (g2130) & (!g2747) & (!g2780) & (!g3805) & (g3806)) + ((!g2099) & (g2130) & (!g2747) & (!g2780) & (g3805) & (!g3806)) + ((!g2099) & (g2130) & (!g2747) & (!g2780) & (g3805) & (g3806)) + ((!g2099) & (g2130) & (g2747) & (!g2780) & (!g3805) & (!g3806)) + ((g2099) & (!g2130) & (!g2747) & (!g2780) & (!g3805) & (!g3806)) + ((g2099) & (!g2130) & (!g2747) & (!g2780) & (!g3805) & (g3806)) + ((g2099) & (!g2130) & (!g2747) & (!g2780) & (g3805) & (!g3806)) + ((g2099) & (!g2130) & (!g2747) & (!g2780) & (g3805) & (g3806)) + ((g2099) & (!g2130) & (!g2747) & (g2780) & (!g3805) & (!g3806)) + ((g2099) & (!g2130) & (g2747) & (!g2780) & (!g3805) & (!g3806)) + ((g2099) & (!g2130) & (g2747) & (!g2780) & (!g3805) & (g3806)) + ((g2099) & (!g2130) & (g2747) & (!g2780) & (g3805) & (!g3806)) + ((g2099) & (!g2130) & (g2747) & (!g2780) & (g3805) & (g3806)) + ((g2099) & (g2130) & (!g2747) & (!g2780) & (!g3805) & (!g3806)));
	assign g3808 = (((!g2178) & (g2830) & (!g3807)) + ((g2178) & (!g2830) & (!g3807)) + ((g2178) & (g2830) & (!g3807)) + ((g2178) & (g2830) & (g3807)));
	assign g3809 = (((!g2211) & (!g2863) & (g3808)) + ((!g2211) & (g2863) & (!g3808)) + ((g2211) & (!g2863) & (!g3808)) + ((g2211) & (g2863) & (g3808)));
	assign g3810 = (((!g830) & (!g1908) & (!g6988) & (key[128])) + ((!g830) & (!g1908) & (g6988) & (key[128])) + ((!g830) & (g1908) & (!g6988) & (key[128])) + ((!g830) & (g1908) & (g6988) & (key[128])) + ((g830) & (!g1908) & (g6988) & (!key[128])) + ((g830) & (!g1908) & (g6988) & (key[128])) + ((g830) & (g1908) & (!g6988) & (!key[128])) + ((g830) & (g1908) & (!g6988) & (key[128])));
	assign g3811 = (((!g1894) & (!g2034) & (g2065) & (!g1902) & (!g2036) & (g2077)) + ((!g1894) & (!g2034) & (g2065) & (!g1902) & (g2036) & (g2077)) + ((!g1894) & (!g2034) & (g2065) & (g1902) & (!g2036) & (g2077)) + ((!g1894) & (!g2034) & (g2065) & (g1902) & (g2036) & (g2077)) + ((!g1894) & (g2034) & (!g2065) & (!g1902) & (g2036) & (g2077)) + ((!g1894) & (g2034) & (!g2065) & (g1902) & (g2036) & (g2077)) + ((!g1894) & (g2034) & (g2065) & (!g1902) & (!g2036) & (g2077)) + ((!g1894) & (g2034) & (g2065) & (!g1902) & (g2036) & (!g2077)) + ((!g1894) & (g2034) & (g2065) & (!g1902) & (g2036) & (g2077)) + ((!g1894) & (g2034) & (g2065) & (g1902) & (!g2036) & (g2077)) + ((!g1894) & (g2034) & (g2065) & (g1902) & (g2036) & (!g2077)) + ((!g1894) & (g2034) & (g2065) & (g1902) & (g2036) & (g2077)) + ((g1894) & (!g2034) & (!g2065) & (g1902) & (g2036) & (g2077)) + ((g1894) & (!g2034) & (g2065) & (!g1902) & (!g2036) & (g2077)) + ((g1894) & (!g2034) & (g2065) & (!g1902) & (g2036) & (g2077)) + ((g1894) & (!g2034) & (g2065) & (g1902) & (!g2036) & (g2077)) + ((g1894) & (!g2034) & (g2065) & (g1902) & (g2036) & (!g2077)) + ((g1894) & (!g2034) & (g2065) & (g1902) & (g2036) & (g2077)) + ((g1894) & (g2034) & (!g2065) & (!g1902) & (g2036) & (g2077)) + ((g1894) & (g2034) & (!g2065) & (g1902) & (!g2036) & (g2077)) + ((g1894) & (g2034) & (!g2065) & (g1902) & (g2036) & (g2077)) + ((g1894) & (g2034) & (g2065) & (!g1902) & (!g2036) & (g2077)) + ((g1894) & (g2034) & (g2065) & (!g1902) & (g2036) & (!g2077)) + ((g1894) & (g2034) & (g2065) & (!g1902) & (g2036) & (g2077)) + ((g1894) & (g2034) & (g2065) & (g1902) & (!g2036) & (!g2077)) + ((g1894) & (g2034) & (g2065) & (g1902) & (!g2036) & (g2077)) + ((g1894) & (g2034) & (g2065) & (g1902) & (g2036) & (!g2077)) + ((g1894) & (g2034) & (g2065) & (g1902) & (g2036) & (g2077)));
	assign g3812 = (((!g2196) & (g2198)) + ((g2196) & (!g2198)));
	assign g3813 = (((!g2116) & (!g2147) & (g2118) & (g2159) & (g3811) & (g3812)) + ((!g2116) & (g2147) & (!g2118) & (g2159) & (!g3811) & (g3812)) + ((!g2116) & (g2147) & (!g2118) & (g2159) & (g3811) & (g3812)) + ((!g2116) & (g2147) & (g2118) & (!g2159) & (g3811) & (g3812)) + ((!g2116) & (g2147) & (g2118) & (g2159) & (!g3811) & (g3812)) + ((!g2116) & (g2147) & (g2118) & (g2159) & (g3811) & (g3812)) + ((g2116) & (!g2147) & (!g2118) & (g2159) & (g3811) & (g3812)) + ((g2116) & (!g2147) & (g2118) & (g2159) & (!g3811) & (g3812)) + ((g2116) & (!g2147) & (g2118) & (g2159) & (g3811) & (g3812)) + ((g2116) & (g2147) & (!g2118) & (!g2159) & (g3811) & (g3812)) + ((g2116) & (g2147) & (!g2118) & (g2159) & (!g3811) & (g3812)) + ((g2116) & (g2147) & (!g2118) & (g2159) & (g3811) & (g3812)) + ((g2116) & (g2147) & (g2118) & (!g2159) & (!g3811) & (g3812)) + ((g2116) & (g2147) & (g2118) & (!g2159) & (g3811) & (g3812)) + ((g2116) & (g2147) & (g2118) & (g2159) & (!g3811) & (g3812)) + ((g2116) & (g2147) & (g2118) & (g2159) & (g3811) & (g3812)));
	assign g3814 = (((g2196) & (g2198)));
	assign g3815 = (((!g2227) & (!g2279) & (!g2239) & (!g2281) & (!g3813) & (!g3814)) + ((!g2227) & (!g2279) & (!g2239) & (!g2281) & (!g3813) & (g3814)) + ((!g2227) & (!g2279) & (!g2239) & (!g2281) & (g3813) & (!g3814)) + ((!g2227) & (!g2279) & (!g2239) & (!g2281) & (g3813) & (g3814)) + ((!g2227) & (!g2279) & (!g2239) & (g2281) & (!g3813) & (!g3814)) + ((!g2227) & (!g2279) & (!g2239) & (g2281) & (!g3813) & (g3814)) + ((!g2227) & (!g2279) & (!g2239) & (g2281) & (g3813) & (!g3814)) + ((!g2227) & (!g2279) & (!g2239) & (g2281) & (g3813) & (g3814)) + ((!g2227) & (!g2279) & (g2239) & (!g2281) & (!g3813) & (!g3814)) + ((!g2227) & (!g2279) & (g2239) & (!g2281) & (!g3813) & (g3814)) + ((!g2227) & (!g2279) & (g2239) & (!g2281) & (g3813) & (!g3814)) + ((!g2227) & (!g2279) & (g2239) & (!g2281) & (g3813) & (g3814)) + ((!g2227) & (!g2279) & (g2239) & (g2281) & (!g3813) & (!g3814)) + ((!g2227) & (g2279) & (!g2239) & (!g2281) & (!g3813) & (!g3814)) + ((!g2227) & (g2279) & (!g2239) & (!g2281) & (!g3813) & (g3814)) + ((!g2227) & (g2279) & (!g2239) & (!g2281) & (g3813) & (!g3814)) + ((!g2227) & (g2279) & (!g2239) & (!g2281) & (g3813) & (g3814)) + ((!g2227) & (g2279) & (g2239) & (!g2281) & (!g3813) & (!g3814)) + ((g2227) & (!g2279) & (!g2239) & (!g2281) & (!g3813) & (!g3814)) + ((g2227) & (!g2279) & (!g2239) & (!g2281) & (!g3813) & (g3814)) + ((g2227) & (!g2279) & (!g2239) & (!g2281) & (g3813) & (!g3814)) + ((g2227) & (!g2279) & (!g2239) & (!g2281) & (g3813) & (g3814)) + ((g2227) & (!g2279) & (!g2239) & (g2281) & (!g3813) & (!g3814)) + ((g2227) & (!g2279) & (g2239) & (!g2281) & (!g3813) & (!g3814)) + ((g2227) & (!g2279) & (g2239) & (!g2281) & (!g3813) & (g3814)) + ((g2227) & (!g2279) & (g2239) & (!g2281) & (g3813) & (!g3814)) + ((g2227) & (!g2279) & (g2239) & (!g2281) & (g3813) & (g3814)) + ((g2227) & (g2279) & (!g2239) & (!g2281) & (!g3813) & (!g3814)));
	assign g3816 = (((!g2393) & (g2405)) + ((g2393) & (!g2405)));
	assign g3817 = (((!g2314) & (!g2362) & (g2326) & (g2364) & (!g3815) & (g3816)) + ((!g2314) & (g2362) & (!g2326) & (g2364) & (!g3815) & (g3816)) + ((!g2314) & (g2362) & (!g2326) & (g2364) & (g3815) & (g3816)) + ((!g2314) & (g2362) & (g2326) & (!g2364) & (!g3815) & (g3816)) + ((!g2314) & (g2362) & (g2326) & (g2364) & (!g3815) & (g3816)) + ((!g2314) & (g2362) & (g2326) & (g2364) & (g3815) & (g3816)) + ((g2314) & (!g2362) & (!g2326) & (g2364) & (!g3815) & (g3816)) + ((g2314) & (!g2362) & (g2326) & (g2364) & (!g3815) & (g3816)) + ((g2314) & (!g2362) & (g2326) & (g2364) & (g3815) & (g3816)) + ((g2314) & (g2362) & (!g2326) & (!g2364) & (!g3815) & (g3816)) + ((g2314) & (g2362) & (!g2326) & (g2364) & (!g3815) & (g3816)) + ((g2314) & (g2362) & (!g2326) & (g2364) & (g3815) & (g3816)) + ((g2314) & (g2362) & (g2326) & (!g2364) & (!g3815) & (g3816)) + ((g2314) & (g2362) & (g2326) & (!g2364) & (g3815) & (g3816)) + ((g2314) & (g2362) & (g2326) & (g2364) & (!g3815) & (g3816)) + ((g2314) & (g2362) & (g2326) & (g2364) & (g3815) & (g3816)));
	assign g3818 = (((g2393) & (g2405)));
	assign g3819 = (((!g2474) & (!g2529) & (!g2480) & (!g2537) & (!g3817) & (!g3818)) + ((!g2474) & (!g2529) & (!g2480) & (!g2537) & (!g3817) & (g3818)) + ((!g2474) & (!g2529) & (!g2480) & (!g2537) & (g3817) & (!g3818)) + ((!g2474) & (!g2529) & (!g2480) & (!g2537) & (g3817) & (g3818)) + ((!g2474) & (!g2529) & (!g2480) & (g2537) & (!g3817) & (!g3818)) + ((!g2474) & (!g2529) & (!g2480) & (g2537) & (!g3817) & (g3818)) + ((!g2474) & (!g2529) & (!g2480) & (g2537) & (g3817) & (!g3818)) + ((!g2474) & (!g2529) & (!g2480) & (g2537) & (g3817) & (g3818)) + ((!g2474) & (!g2529) & (g2480) & (!g2537) & (!g3817) & (!g3818)) + ((!g2474) & (!g2529) & (g2480) & (!g2537) & (!g3817) & (g3818)) + ((!g2474) & (!g2529) & (g2480) & (!g2537) & (g3817) & (!g3818)) + ((!g2474) & (!g2529) & (g2480) & (!g2537) & (g3817) & (g3818)) + ((!g2474) & (!g2529) & (g2480) & (g2537) & (!g3817) & (!g3818)) + ((!g2474) & (g2529) & (!g2480) & (!g2537) & (!g3817) & (!g3818)) + ((!g2474) & (g2529) & (!g2480) & (!g2537) & (!g3817) & (g3818)) + ((!g2474) & (g2529) & (!g2480) & (!g2537) & (g3817) & (!g3818)) + ((!g2474) & (g2529) & (!g2480) & (!g2537) & (g3817) & (g3818)) + ((!g2474) & (g2529) & (g2480) & (!g2537) & (!g3817) & (!g3818)) + ((g2474) & (!g2529) & (!g2480) & (!g2537) & (!g3817) & (!g3818)) + ((g2474) & (!g2529) & (!g2480) & (!g2537) & (!g3817) & (g3818)) + ((g2474) & (!g2529) & (!g2480) & (!g2537) & (g3817) & (!g3818)) + ((g2474) & (!g2529) & (!g2480) & (!g2537) & (g3817) & (g3818)) + ((g2474) & (!g2529) & (!g2480) & (g2537) & (!g3817) & (!g3818)) + ((g2474) & (!g2529) & (g2480) & (!g2537) & (!g3817) & (!g3818)) + ((g2474) & (!g2529) & (g2480) & (!g2537) & (!g3817) & (g3818)) + ((g2474) & (!g2529) & (g2480) & (!g2537) & (g3817) & (!g3818)) + ((g2474) & (!g2529) & (g2480) & (!g2537) & (g3817) & (g3818)) + ((g2474) & (g2529) & (!g2480) & (!g2537) & (!g3817) & (!g3818)));
	assign g3820 = (((!g2474) & (!g2480) & (!g3817) & (!g3818) & (!g5824) & (g5825)) + ((!g2474) & (!g2480) & (!g3817) & (g3818) & (!g5824) & (g5825)) + ((!g2474) & (!g2480) & (g3817) & (!g3818) & (!g5824) & (g5825)) + ((!g2474) & (!g2480) & (g3817) & (g3818) & (!g5824) & (g5825)) + ((!g2474) & (g2480) & (!g3817) & (!g3818) & (!g5824) & (g5825)) + ((!g2474) & (g2480) & (!g3817) & (g3818) & (!g5824) & (g5825)) + ((!g2474) & (g2480) & (!g3817) & (g3818) & (g5824) & (g5825)) + ((!g2474) & (g2480) & (g3817) & (!g3818) & (!g5824) & (g5825)) + ((!g2474) & (g2480) & (g3817) & (!g3818) & (g5824) & (g5825)) + ((!g2474) & (g2480) & (g3817) & (g3818) & (!g5824) & (g5825)) + ((!g2474) & (g2480) & (g3817) & (g3818) & (g5824) & (g5825)) + ((g2474) & (!g2480) & (!g3817) & (!g3818) & (!g5824) & (g5825)) + ((g2474) & (!g2480) & (!g3817) & (g3818) & (!g5824) & (g5825)) + ((g2474) & (!g2480) & (!g3817) & (g3818) & (g5824) & (g5825)) + ((g2474) & (!g2480) & (g3817) & (!g3818) & (!g5824) & (g5825)) + ((g2474) & (!g2480) & (g3817) & (!g3818) & (g5824) & (g5825)) + ((g2474) & (!g2480) & (g3817) & (g3818) & (!g5824) & (g5825)) + ((g2474) & (!g2480) & (g3817) & (g3818) & (g5824) & (g5825)) + ((g2474) & (g2480) & (!g3817) & (!g3818) & (!g5824) & (g5825)) + ((g2474) & (g2480) & (!g3817) & (!g3818) & (g5824) & (g5825)) + ((g2474) & (g2480) & (!g3817) & (g3818) & (!g5824) & (g5825)) + ((g2474) & (g2480) & (!g3817) & (g3818) & (g5824) & (g5825)) + ((g2474) & (g2480) & (g3817) & (!g3818) & (!g5824) & (g5825)) + ((g2474) & (g2480) & (g3817) & (!g3818) & (g5824) & (g5825)) + ((g2474) & (g2480) & (g3817) & (g3818) & (!g5824) & (g5825)) + ((g2474) & (g2480) & (g3817) & (g3818) & (g5824) & (g5825)));
	assign g3821 = (((g2665) & (g2667)));
	assign g3822 = (((!g2708) & (!g2776) & (!g2728) & (!g2778) & (!g3820) & (!g3821)) + ((!g2708) & (!g2776) & (!g2728) & (!g2778) & (!g3820) & (g3821)) + ((!g2708) & (!g2776) & (!g2728) & (!g2778) & (g3820) & (!g3821)) + ((!g2708) & (!g2776) & (!g2728) & (!g2778) & (g3820) & (g3821)) + ((!g2708) & (!g2776) & (!g2728) & (g2778) & (!g3820) & (!g3821)) + ((!g2708) & (!g2776) & (!g2728) & (g2778) & (!g3820) & (g3821)) + ((!g2708) & (!g2776) & (!g2728) & (g2778) & (g3820) & (!g3821)) + ((!g2708) & (!g2776) & (!g2728) & (g2778) & (g3820) & (g3821)) + ((!g2708) & (!g2776) & (g2728) & (!g2778) & (!g3820) & (!g3821)) + ((!g2708) & (!g2776) & (g2728) & (!g2778) & (!g3820) & (g3821)) + ((!g2708) & (!g2776) & (g2728) & (!g2778) & (g3820) & (!g3821)) + ((!g2708) & (!g2776) & (g2728) & (!g2778) & (g3820) & (g3821)) + ((!g2708) & (!g2776) & (g2728) & (g2778) & (!g3820) & (!g3821)) + ((!g2708) & (g2776) & (!g2728) & (!g2778) & (!g3820) & (!g3821)) + ((!g2708) & (g2776) & (!g2728) & (!g2778) & (!g3820) & (g3821)) + ((!g2708) & (g2776) & (!g2728) & (!g2778) & (g3820) & (!g3821)) + ((!g2708) & (g2776) & (!g2728) & (!g2778) & (g3820) & (g3821)) + ((!g2708) & (g2776) & (g2728) & (!g2778) & (!g3820) & (!g3821)) + ((g2708) & (!g2776) & (!g2728) & (!g2778) & (!g3820) & (!g3821)) + ((g2708) & (!g2776) & (!g2728) & (!g2778) & (!g3820) & (g3821)) + ((g2708) & (!g2776) & (!g2728) & (!g2778) & (g3820) & (!g3821)) + ((g2708) & (!g2776) & (!g2728) & (!g2778) & (g3820) & (g3821)) + ((g2708) & (!g2776) & (!g2728) & (g2778) & (!g3820) & (!g3821)) + ((g2708) & (!g2776) & (g2728) & (!g2778) & (!g3820) & (!g3821)) + ((g2708) & (!g2776) & (g2728) & (!g2778) & (!g3820) & (g3821)) + ((g2708) & (!g2776) & (g2728) & (!g2778) & (g3820) & (!g3821)) + ((g2708) & (!g2776) & (g2728) & (!g2778) & (g3820) & (g3821)) + ((g2708) & (g2776) & (!g2728) & (!g2778) & (!g3820) & (!g3821)));
	assign g3823 = (((!g2895) & (g2887)) + ((g2895) & (!g2887)));
	assign g3824 = (((!g2807) & (!g2857) & (g2819) & (g2860) & (!g3822) & (g3823)) + ((!g2807) & (g2857) & (!g2819) & (g2860) & (!g3822) & (g3823)) + ((!g2807) & (g2857) & (!g2819) & (g2860) & (g3822) & (g3823)) + ((!g2807) & (g2857) & (g2819) & (!g2860) & (!g3822) & (g3823)) + ((!g2807) & (g2857) & (g2819) & (g2860) & (!g3822) & (g3823)) + ((!g2807) & (g2857) & (g2819) & (g2860) & (g3822) & (g3823)) + ((g2807) & (!g2857) & (!g2819) & (g2860) & (!g3822) & (g3823)) + ((g2807) & (!g2857) & (g2819) & (g2860) & (!g3822) & (g3823)) + ((g2807) & (!g2857) & (g2819) & (g2860) & (g3822) & (g3823)) + ((g2807) & (g2857) & (!g2819) & (!g2860) & (!g3822) & (g3823)) + ((g2807) & (g2857) & (!g2819) & (g2860) & (!g3822) & (g3823)) + ((g2807) & (g2857) & (!g2819) & (g2860) & (g3822) & (g3823)) + ((g2807) & (g2857) & (g2819) & (!g2860) & (!g3822) & (g3823)) + ((g2807) & (g2857) & (g2819) & (!g2860) & (g3822) & (g3823)) + ((g2807) & (g2857) & (g2819) & (g2860) & (!g3822) & (g3823)) + ((g2807) & (g2857) & (g2819) & (g2860) & (g3822) & (g3823)));
	assign g3825 = (((g2895) & (g2887)));
	assign g3826 = (((!g2962) & (!g3013) & (!g2956) & (!g3005) & (!g3824) & (!g3825)) + ((!g2962) & (!g3013) & (!g2956) & (!g3005) & (!g3824) & (g3825)) + ((!g2962) & (!g3013) & (!g2956) & (!g3005) & (g3824) & (!g3825)) + ((!g2962) & (!g3013) & (!g2956) & (!g3005) & (g3824) & (g3825)) + ((!g2962) & (!g3013) & (!g2956) & (g3005) & (!g3824) & (!g3825)) + ((!g2962) & (!g3013) & (!g2956) & (g3005) & (!g3824) & (g3825)) + ((!g2962) & (!g3013) & (!g2956) & (g3005) & (g3824) & (!g3825)) + ((!g2962) & (!g3013) & (!g2956) & (g3005) & (g3824) & (g3825)) + ((!g2962) & (!g3013) & (g2956) & (!g3005) & (!g3824) & (!g3825)) + ((!g2962) & (!g3013) & (g2956) & (!g3005) & (!g3824) & (g3825)) + ((!g2962) & (!g3013) & (g2956) & (!g3005) & (g3824) & (!g3825)) + ((!g2962) & (!g3013) & (g2956) & (!g3005) & (g3824) & (g3825)) + ((!g2962) & (!g3013) & (g2956) & (g3005) & (!g3824) & (!g3825)) + ((!g2962) & (g3013) & (!g2956) & (!g3005) & (!g3824) & (!g3825)) + ((!g2962) & (g3013) & (!g2956) & (!g3005) & (!g3824) & (g3825)) + ((!g2962) & (g3013) & (!g2956) & (!g3005) & (g3824) & (!g3825)) + ((!g2962) & (g3013) & (!g2956) & (!g3005) & (g3824) & (g3825)) + ((!g2962) & (g3013) & (g2956) & (!g3005) & (!g3824) & (!g3825)) + ((g2962) & (!g3013) & (!g2956) & (!g3005) & (!g3824) & (!g3825)) + ((g2962) & (!g3013) & (!g2956) & (!g3005) & (!g3824) & (g3825)) + ((g2962) & (!g3013) & (!g2956) & (!g3005) & (g3824) & (!g3825)) + ((g2962) & (!g3013) & (!g2956) & (!g3005) & (g3824) & (g3825)) + ((g2962) & (!g3013) & (!g2956) & (g3005) & (!g3824) & (!g3825)) + ((g2962) & (!g3013) & (g2956) & (!g3005) & (!g3824) & (!g3825)) + ((g2962) & (!g3013) & (g2956) & (!g3005) & (!g3824) & (g3825)) + ((g2962) & (!g3013) & (g2956) & (!g3005) & (g3824) & (!g3825)) + ((g2962) & (!g3013) & (g2956) & (!g3005) & (g3824) & (g3825)) + ((g2962) & (g3013) & (!g2956) & (!g3005) & (!g3824) & (!g3825)));
	assign g3827 = (((g1914) & (!g3053) & (!g3050) & (!g3826)) + ((g1914) & (!g3053) & (g3050) & (g3826)) + ((g1914) & (g3053) & (!g3050) & (g3826)) + ((g1914) & (g3053) & (g3050) & (!g3826)));
	assign g3828 = (((!g1906) & (!g1940) & (g1942) & (!g1912) & (!g2045) & (g2091)) + ((!g1906) & (!g1940) & (g1942) & (!g1912) & (g2045) & (g2091)) + ((!g1906) & (!g1940) & (g1942) & (g1912) & (!g2045) & (g2091)) + ((!g1906) & (!g1940) & (g1942) & (g1912) & (g2045) & (g2091)) + ((!g1906) & (g1940) & (!g1942) & (!g1912) & (g2045) & (g2091)) + ((!g1906) & (g1940) & (!g1942) & (g1912) & (g2045) & (g2091)) + ((!g1906) & (g1940) & (g1942) & (!g1912) & (!g2045) & (g2091)) + ((!g1906) & (g1940) & (g1942) & (!g1912) & (g2045) & (!g2091)) + ((!g1906) & (g1940) & (g1942) & (!g1912) & (g2045) & (g2091)) + ((!g1906) & (g1940) & (g1942) & (g1912) & (!g2045) & (g2091)) + ((!g1906) & (g1940) & (g1942) & (g1912) & (g2045) & (!g2091)) + ((!g1906) & (g1940) & (g1942) & (g1912) & (g2045) & (g2091)) + ((g1906) & (!g1940) & (!g1942) & (g1912) & (g2045) & (g2091)) + ((g1906) & (!g1940) & (g1942) & (!g1912) & (!g2045) & (g2091)) + ((g1906) & (!g1940) & (g1942) & (!g1912) & (g2045) & (g2091)) + ((g1906) & (!g1940) & (g1942) & (g1912) & (!g2045) & (g2091)) + ((g1906) & (!g1940) & (g1942) & (g1912) & (g2045) & (!g2091)) + ((g1906) & (!g1940) & (g1942) & (g1912) & (g2045) & (g2091)) + ((g1906) & (g1940) & (!g1942) & (!g1912) & (g2045) & (g2091)) + ((g1906) & (g1940) & (!g1942) & (g1912) & (!g2045) & (g2091)) + ((g1906) & (g1940) & (!g1942) & (g1912) & (g2045) & (g2091)) + ((g1906) & (g1940) & (g1942) & (!g1912) & (!g2045) & (g2091)) + ((g1906) & (g1940) & (g1942) & (!g1912) & (g2045) & (!g2091)) + ((g1906) & (g1940) & (g1942) & (!g1912) & (g2045) & (g2091)) + ((g1906) & (g1940) & (g1942) & (g1912) & (!g2045) & (!g2091)) + ((g1906) & (g1940) & (g1942) & (g1912) & (!g2045) & (g2091)) + ((g1906) & (g1940) & (g1942) & (g1912) & (g2045) & (!g2091)) + ((g1906) & (g1940) & (g1942) & (g1912) & (g2045) & (g2091)));
	assign g3829 = (((!g1949) & (g2207)) + ((g1949) & (!g2207)));
	assign g3830 = (((!g1945) & (!g1947) & (g2127) & (g2173) & (g3828) & (g3829)) + ((!g1945) & (g1947) & (!g2127) & (g2173) & (!g3828) & (g3829)) + ((!g1945) & (g1947) & (!g2127) & (g2173) & (g3828) & (g3829)) + ((!g1945) & (g1947) & (g2127) & (!g2173) & (g3828) & (g3829)) + ((!g1945) & (g1947) & (g2127) & (g2173) & (!g3828) & (g3829)) + ((!g1945) & (g1947) & (g2127) & (g2173) & (g3828) & (g3829)) + ((g1945) & (!g1947) & (!g2127) & (g2173) & (g3828) & (g3829)) + ((g1945) & (!g1947) & (g2127) & (g2173) & (!g3828) & (g3829)) + ((g1945) & (!g1947) & (g2127) & (g2173) & (g3828) & (g3829)) + ((g1945) & (g1947) & (!g2127) & (!g2173) & (g3828) & (g3829)) + ((g1945) & (g1947) & (!g2127) & (g2173) & (!g3828) & (g3829)) + ((g1945) & (g1947) & (!g2127) & (g2173) & (g3828) & (g3829)) + ((g1945) & (g1947) & (g2127) & (!g2173) & (!g3828) & (g3829)) + ((g1945) & (g1947) & (g2127) & (!g2173) & (g3828) & (g3829)) + ((g1945) & (g1947) & (g2127) & (g2173) & (!g3828) & (g3829)) + ((g1945) & (g1947) & (g2127) & (g2173) & (g3828) & (g3829)));
	assign g3831 = (((g1949) & (g2207)));
	assign g3832 = (((!g1954) & (!g1956) & (!g2253) & (!g2290) & (!g3830) & (!g3831)) + ((!g1954) & (!g1956) & (!g2253) & (!g2290) & (!g3830) & (g3831)) + ((!g1954) & (!g1956) & (!g2253) & (!g2290) & (g3830) & (!g3831)) + ((!g1954) & (!g1956) & (!g2253) & (!g2290) & (g3830) & (g3831)) + ((!g1954) & (!g1956) & (!g2253) & (g2290) & (!g3830) & (!g3831)) + ((!g1954) & (!g1956) & (!g2253) & (g2290) & (!g3830) & (g3831)) + ((!g1954) & (!g1956) & (!g2253) & (g2290) & (g3830) & (!g3831)) + ((!g1954) & (!g1956) & (!g2253) & (g2290) & (g3830) & (g3831)) + ((!g1954) & (!g1956) & (g2253) & (!g2290) & (!g3830) & (!g3831)) + ((!g1954) & (!g1956) & (g2253) & (!g2290) & (!g3830) & (g3831)) + ((!g1954) & (!g1956) & (g2253) & (!g2290) & (g3830) & (!g3831)) + ((!g1954) & (!g1956) & (g2253) & (!g2290) & (g3830) & (g3831)) + ((!g1954) & (!g1956) & (g2253) & (g2290) & (!g3830) & (!g3831)) + ((!g1954) & (g1956) & (!g2253) & (!g2290) & (!g3830) & (!g3831)) + ((!g1954) & (g1956) & (!g2253) & (!g2290) & (!g3830) & (g3831)) + ((!g1954) & (g1956) & (!g2253) & (!g2290) & (g3830) & (!g3831)) + ((!g1954) & (g1956) & (!g2253) & (!g2290) & (g3830) & (g3831)) + ((!g1954) & (g1956) & (g2253) & (!g2290) & (!g3830) & (!g3831)) + ((g1954) & (!g1956) & (!g2253) & (!g2290) & (!g3830) & (!g3831)) + ((g1954) & (!g1956) & (!g2253) & (!g2290) & (!g3830) & (g3831)) + ((g1954) & (!g1956) & (!g2253) & (!g2290) & (g3830) & (!g3831)) + ((g1954) & (!g1956) & (!g2253) & (!g2290) & (g3830) & (g3831)) + ((g1954) & (!g1956) & (!g2253) & (g2290) & (!g3830) & (!g3831)) + ((g1954) & (!g1956) & (g2253) & (!g2290) & (!g3830) & (!g3831)) + ((g1954) & (!g1956) & (g2253) & (!g2290) & (!g3830) & (g3831)) + ((g1954) & (!g1956) & (g2253) & (!g2290) & (g3830) & (!g3831)) + ((g1954) & (!g1956) & (g2253) & (!g2290) & (g3830) & (g3831)) + ((g1954) & (g1956) & (!g2253) & (!g2290) & (!g3830) & (!g3831)));
	assign g3833 = (((!g1963) & (g2419)) + ((g1963) & (!g2419)));
	assign g3834 = (((!g1959) & (!g1961) & (g2340) & (g2373) & (!g3832) & (g3833)) + ((!g1959) & (g1961) & (!g2340) & (g2373) & (!g3832) & (g3833)) + ((!g1959) & (g1961) & (!g2340) & (g2373) & (g3832) & (g3833)) + ((!g1959) & (g1961) & (g2340) & (!g2373) & (!g3832) & (g3833)) + ((!g1959) & (g1961) & (g2340) & (g2373) & (!g3832) & (g3833)) + ((!g1959) & (g1961) & (g2340) & (g2373) & (g3832) & (g3833)) + ((g1959) & (!g1961) & (!g2340) & (g2373) & (!g3832) & (g3833)) + ((g1959) & (!g1961) & (g2340) & (g2373) & (!g3832) & (g3833)) + ((g1959) & (!g1961) & (g2340) & (g2373) & (g3832) & (g3833)) + ((g1959) & (g1961) & (!g2340) & (!g2373) & (!g3832) & (g3833)) + ((g1959) & (g1961) & (!g2340) & (g2373) & (!g3832) & (g3833)) + ((g1959) & (g1961) & (!g2340) & (g2373) & (g3832) & (g3833)) + ((g1959) & (g1961) & (g2340) & (!g2373) & (!g3832) & (g3833)) + ((g1959) & (g1961) & (g2340) & (!g2373) & (g3832) & (g3833)) + ((g1959) & (g1961) & (g2340) & (g2373) & (!g3832) & (g3833)) + ((g1959) & (g1961) & (g2340) & (g2373) & (g3832) & (g3833)));
	assign g3835 = (((g1963) & (g2419)));
	assign g3836 = (((!g1968) & (!g1970) & (!g2509) & (!g2546) & (!g3834) & (!g3835)) + ((!g1968) & (!g1970) & (!g2509) & (!g2546) & (!g3834) & (g3835)) + ((!g1968) & (!g1970) & (!g2509) & (!g2546) & (g3834) & (!g3835)) + ((!g1968) & (!g1970) & (!g2509) & (!g2546) & (g3834) & (g3835)) + ((!g1968) & (!g1970) & (!g2509) & (g2546) & (!g3834) & (!g3835)) + ((!g1968) & (!g1970) & (!g2509) & (g2546) & (!g3834) & (g3835)) + ((!g1968) & (!g1970) & (!g2509) & (g2546) & (g3834) & (!g3835)) + ((!g1968) & (!g1970) & (!g2509) & (g2546) & (g3834) & (g3835)) + ((!g1968) & (!g1970) & (g2509) & (!g2546) & (!g3834) & (!g3835)) + ((!g1968) & (!g1970) & (g2509) & (!g2546) & (!g3834) & (g3835)) + ((!g1968) & (!g1970) & (g2509) & (!g2546) & (g3834) & (!g3835)) + ((!g1968) & (!g1970) & (g2509) & (!g2546) & (g3834) & (g3835)) + ((!g1968) & (!g1970) & (g2509) & (g2546) & (!g3834) & (!g3835)) + ((!g1968) & (g1970) & (!g2509) & (!g2546) & (!g3834) & (!g3835)) + ((!g1968) & (g1970) & (!g2509) & (!g2546) & (!g3834) & (g3835)) + ((!g1968) & (g1970) & (!g2509) & (!g2546) & (g3834) & (!g3835)) + ((!g1968) & (g1970) & (!g2509) & (!g2546) & (g3834) & (g3835)) + ((!g1968) & (g1970) & (g2509) & (!g2546) & (!g3834) & (!g3835)) + ((g1968) & (!g1970) & (!g2509) & (!g2546) & (!g3834) & (!g3835)) + ((g1968) & (!g1970) & (!g2509) & (!g2546) & (!g3834) & (g3835)) + ((g1968) & (!g1970) & (!g2509) & (!g2546) & (g3834) & (!g3835)) + ((g1968) & (!g1970) & (!g2509) & (!g2546) & (g3834) & (g3835)) + ((g1968) & (!g1970) & (!g2509) & (g2546) & (!g3834) & (!g3835)) + ((g1968) & (!g1970) & (g2509) & (!g2546) & (!g3834) & (!g3835)) + ((g1968) & (!g1970) & (g2509) & (!g2546) & (!g3834) & (g3835)) + ((g1968) & (!g1970) & (g2509) & (!g2546) & (g3834) & (!g3835)) + ((g1968) & (!g1970) & (g2509) & (!g2546) & (g3834) & (g3835)) + ((g1968) & (g1970) & (!g2509) & (!g2546) & (!g3834) & (!g3835)));
	assign g3837 = (((!g1968) & (!g2509) & (!g3834) & (!g3835) & (!g5827) & (g5828)) + ((!g1968) & (!g2509) & (!g3834) & (g3835) & (!g5827) & (g5828)) + ((!g1968) & (!g2509) & (g3834) & (!g3835) & (!g5827) & (g5828)) + ((!g1968) & (!g2509) & (g3834) & (g3835) & (!g5827) & (g5828)) + ((!g1968) & (g2509) & (!g3834) & (!g3835) & (!g5827) & (g5828)) + ((!g1968) & (g2509) & (!g3834) & (g3835) & (!g5827) & (g5828)) + ((!g1968) & (g2509) & (!g3834) & (g3835) & (g5827) & (g5828)) + ((!g1968) & (g2509) & (g3834) & (!g3835) & (!g5827) & (g5828)) + ((!g1968) & (g2509) & (g3834) & (!g3835) & (g5827) & (g5828)) + ((!g1968) & (g2509) & (g3834) & (g3835) & (!g5827) & (g5828)) + ((!g1968) & (g2509) & (g3834) & (g3835) & (g5827) & (g5828)) + ((g1968) & (!g2509) & (!g3834) & (!g3835) & (!g5827) & (g5828)) + ((g1968) & (!g2509) & (!g3834) & (g3835) & (!g5827) & (g5828)) + ((g1968) & (!g2509) & (!g3834) & (g3835) & (g5827) & (g5828)) + ((g1968) & (!g2509) & (g3834) & (!g3835) & (!g5827) & (g5828)) + ((g1968) & (!g2509) & (g3834) & (!g3835) & (g5827) & (g5828)) + ((g1968) & (!g2509) & (g3834) & (g3835) & (!g5827) & (g5828)) + ((g1968) & (!g2509) & (g3834) & (g3835) & (g5827) & (g5828)) + ((g1968) & (g2509) & (!g3834) & (!g3835) & (!g5827) & (g5828)) + ((g1968) & (g2509) & (!g3834) & (!g3835) & (g5827) & (g5828)) + ((g1968) & (g2509) & (!g3834) & (g3835) & (!g5827) & (g5828)) + ((g1968) & (g2509) & (!g3834) & (g3835) & (g5827) & (g5828)) + ((g1968) & (g2509) & (g3834) & (!g3835) & (!g5827) & (g5828)) + ((g1968) & (g2509) & (g3834) & (!g3835) & (g5827) & (g5828)) + ((g1968) & (g2509) & (g3834) & (g3835) & (!g5827) & (g5828)) + ((g1968) & (g2509) & (g3834) & (g3835) & (g5827) & (g5828)));
	assign g3838 = (((g2048) & (g2676)));
	assign g3839 = (((!g2099) & (!g2130) & (!g2752) & (!g2787) & (!g3837) & (!g3838)) + ((!g2099) & (!g2130) & (!g2752) & (!g2787) & (!g3837) & (g3838)) + ((!g2099) & (!g2130) & (!g2752) & (!g2787) & (g3837) & (!g3838)) + ((!g2099) & (!g2130) & (!g2752) & (!g2787) & (g3837) & (g3838)) + ((!g2099) & (!g2130) & (!g2752) & (g2787) & (!g3837) & (!g3838)) + ((!g2099) & (!g2130) & (!g2752) & (g2787) & (!g3837) & (g3838)) + ((!g2099) & (!g2130) & (!g2752) & (g2787) & (g3837) & (!g3838)) + ((!g2099) & (!g2130) & (!g2752) & (g2787) & (g3837) & (g3838)) + ((!g2099) & (!g2130) & (g2752) & (!g2787) & (!g3837) & (!g3838)) + ((!g2099) & (!g2130) & (g2752) & (!g2787) & (!g3837) & (g3838)) + ((!g2099) & (!g2130) & (g2752) & (!g2787) & (g3837) & (!g3838)) + ((!g2099) & (!g2130) & (g2752) & (!g2787) & (g3837) & (g3838)) + ((!g2099) & (!g2130) & (g2752) & (g2787) & (!g3837) & (!g3838)) + ((!g2099) & (g2130) & (!g2752) & (!g2787) & (!g3837) & (!g3838)) + ((!g2099) & (g2130) & (!g2752) & (!g2787) & (!g3837) & (g3838)) + ((!g2099) & (g2130) & (!g2752) & (!g2787) & (g3837) & (!g3838)) + ((!g2099) & (g2130) & (!g2752) & (!g2787) & (g3837) & (g3838)) + ((!g2099) & (g2130) & (g2752) & (!g2787) & (!g3837) & (!g3838)) + ((g2099) & (!g2130) & (!g2752) & (!g2787) & (!g3837) & (!g3838)) + ((g2099) & (!g2130) & (!g2752) & (!g2787) & (!g3837) & (g3838)) + ((g2099) & (!g2130) & (!g2752) & (!g2787) & (g3837) & (!g3838)) + ((g2099) & (!g2130) & (!g2752) & (!g2787) & (g3837) & (g3838)) + ((g2099) & (!g2130) & (!g2752) & (g2787) & (!g3837) & (!g3838)) + ((g2099) & (!g2130) & (g2752) & (!g2787) & (!g3837) & (!g3838)) + ((g2099) & (!g2130) & (g2752) & (!g2787) & (!g3837) & (g3838)) + ((g2099) & (!g2130) & (g2752) & (!g2787) & (g3837) & (!g3838)) + ((g2099) & (!g2130) & (g2752) & (!g2787) & (g3837) & (g3838)) + ((g2099) & (g2130) & (!g2752) & (!g2787) & (!g3837) & (!g3838)));
	assign g3840 = (((!g2257) & (g2904)) + ((g2257) & (!g2904)));
	assign g3841 = (((!g2178) & (!g2211) & (g2833) & (g2874) & (!g3839) & (g3840)) + ((!g2178) & (g2211) & (!g2833) & (g2874) & (!g3839) & (g3840)) + ((!g2178) & (g2211) & (!g2833) & (g2874) & (g3839) & (g3840)) + ((!g2178) & (g2211) & (g2833) & (!g2874) & (!g3839) & (g3840)) + ((!g2178) & (g2211) & (g2833) & (g2874) & (!g3839) & (g3840)) + ((!g2178) & (g2211) & (g2833) & (g2874) & (g3839) & (g3840)) + ((g2178) & (!g2211) & (!g2833) & (g2874) & (!g3839) & (g3840)) + ((g2178) & (!g2211) & (g2833) & (g2874) & (!g3839) & (g3840)) + ((g2178) & (!g2211) & (g2833) & (g2874) & (g3839) & (g3840)) + ((g2178) & (g2211) & (!g2833) & (!g2874) & (!g3839) & (g3840)) + ((g2178) & (g2211) & (!g2833) & (g2874) & (!g3839) & (g3840)) + ((g2178) & (g2211) & (!g2833) & (g2874) & (g3839) & (g3840)) + ((g2178) & (g2211) & (g2833) & (!g2874) & (!g3839) & (g3840)) + ((g2178) & (g2211) & (g2833) & (!g2874) & (g3839) & (g3840)) + ((g2178) & (g2211) & (g2833) & (g2874) & (!g3839) & (g3840)) + ((g2178) & (g2211) & (g2833) & (g2874) & (g3839) & (g3840)));
	assign g3842 = (((g2257) & (g2904)));
	assign g3843 = (((!g2296) & (!g2344) & (!g2991) & (!g3022) & (!g3841) & (!g3842)) + ((!g2296) & (!g2344) & (!g2991) & (!g3022) & (!g3841) & (g3842)) + ((!g2296) & (!g2344) & (!g2991) & (!g3022) & (g3841) & (!g3842)) + ((!g2296) & (!g2344) & (!g2991) & (!g3022) & (g3841) & (g3842)) + ((!g2296) & (!g2344) & (!g2991) & (g3022) & (!g3841) & (!g3842)) + ((!g2296) & (!g2344) & (!g2991) & (g3022) & (!g3841) & (g3842)) + ((!g2296) & (!g2344) & (!g2991) & (g3022) & (g3841) & (!g3842)) + ((!g2296) & (!g2344) & (!g2991) & (g3022) & (g3841) & (g3842)) + ((!g2296) & (!g2344) & (g2991) & (!g3022) & (!g3841) & (!g3842)) + ((!g2296) & (!g2344) & (g2991) & (!g3022) & (!g3841) & (g3842)) + ((!g2296) & (!g2344) & (g2991) & (!g3022) & (g3841) & (!g3842)) + ((!g2296) & (!g2344) & (g2991) & (!g3022) & (g3841) & (g3842)) + ((!g2296) & (!g2344) & (g2991) & (g3022) & (!g3841) & (!g3842)) + ((!g2296) & (g2344) & (!g2991) & (!g3022) & (!g3841) & (!g3842)) + ((!g2296) & (g2344) & (!g2991) & (!g3022) & (!g3841) & (g3842)) + ((!g2296) & (g2344) & (!g2991) & (!g3022) & (g3841) & (!g3842)) + ((!g2296) & (g2344) & (!g2991) & (!g3022) & (g3841) & (g3842)) + ((!g2296) & (g2344) & (g2991) & (!g3022) & (!g3841) & (!g3842)) + ((g2296) & (!g2344) & (!g2991) & (!g3022) & (!g3841) & (!g3842)) + ((g2296) & (!g2344) & (!g2991) & (!g3022) & (!g3841) & (g3842)) + ((g2296) & (!g2344) & (!g2991) & (!g3022) & (g3841) & (!g3842)) + ((g2296) & (!g2344) & (!g2991) & (!g3022) & (g3841) & (g3842)) + ((g2296) & (!g2344) & (!g2991) & (g3022) & (!g3841) & (!g3842)) + ((g2296) & (!g2344) & (g2991) & (!g3022) & (!g3841) & (!g3842)) + ((g2296) & (!g2344) & (g2991) & (!g3022) & (!g3841) & (g3842)) + ((g2296) & (!g2344) & (g2991) & (!g3022) & (g3841) & (!g3842)) + ((g2296) & (!g2344) & (g2991) & (!g3022) & (g3841) & (g3842)) + ((g2296) & (g2344) & (!g2991) & (!g3022) & (!g3841) & (!g3842)));
	assign g3844 = (((!g1914) & (!g2377) & (!g3067) & (!g3843)) + ((!g1914) & (!g2377) & (g3067) & (g3843)) + ((!g1914) & (g2377) & (!g3067) & (g3843)) + ((!g1914) & (g2377) & (g3067) & (!g3843)));
	assign g3845 = (((!g830) & (!g1910) & (!g3827) & (!g3844) & (nonce[32])) + ((!g830) & (!g1910) & (!g3827) & (g3844) & (nonce[32])) + ((!g830) & (!g1910) & (g3827) & (!g3844) & (nonce[32])) + ((!g830) & (!g1910) & (g3827) & (g3844) & (nonce[32])) + ((!g830) & (g1910) & (!g3827) & (!g3844) & (nonce[32])) + ((!g830) & (g1910) & (!g3827) & (g3844) & (nonce[32])) + ((!g830) & (g1910) & (g3827) & (!g3844) & (nonce[32])) + ((!g830) & (g1910) & (g3827) & (g3844) & (nonce[32])) + ((g830) & (!g1910) & (!g3827) & (g3844) & (!nonce[32])) + ((g830) & (!g1910) & (!g3827) & (g3844) & (nonce[32])) + ((g830) & (!g1910) & (g3827) & (!g3844) & (!nonce[32])) + ((g830) & (!g1910) & (g3827) & (!g3844) & (nonce[32])) + ((g830) & (!g1910) & (g3827) & (g3844) & (!nonce[32])) + ((g830) & (!g1910) & (g3827) & (g3844) & (nonce[32])) + ((g830) & (g1910) & (!g3827) & (!g3844) & (!nonce[32])) + ((g830) & (g1910) & (!g3827) & (!g3844) & (nonce[32])));
	assign g3846 = (((!g1896) & (!g2041) & (g2068) & (!g1904) & (!g2043) & (g2080)) + ((!g1896) & (!g2041) & (g2068) & (!g1904) & (g2043) & (g2080)) + ((!g1896) & (!g2041) & (g2068) & (g1904) & (!g2043) & (g2080)) + ((!g1896) & (!g2041) & (g2068) & (g1904) & (g2043) & (g2080)) + ((!g1896) & (g2041) & (!g2068) & (!g1904) & (g2043) & (g2080)) + ((!g1896) & (g2041) & (!g2068) & (g1904) & (g2043) & (g2080)) + ((!g1896) & (g2041) & (g2068) & (!g1904) & (!g2043) & (g2080)) + ((!g1896) & (g2041) & (g2068) & (!g1904) & (g2043) & (!g2080)) + ((!g1896) & (g2041) & (g2068) & (!g1904) & (g2043) & (g2080)) + ((!g1896) & (g2041) & (g2068) & (g1904) & (!g2043) & (g2080)) + ((!g1896) & (g2041) & (g2068) & (g1904) & (g2043) & (!g2080)) + ((!g1896) & (g2041) & (g2068) & (g1904) & (g2043) & (g2080)) + ((g1896) & (!g2041) & (!g2068) & (g1904) & (g2043) & (g2080)) + ((g1896) & (!g2041) & (g2068) & (!g1904) & (!g2043) & (g2080)) + ((g1896) & (!g2041) & (g2068) & (!g1904) & (g2043) & (g2080)) + ((g1896) & (!g2041) & (g2068) & (g1904) & (!g2043) & (g2080)) + ((g1896) & (!g2041) & (g2068) & (g1904) & (g2043) & (!g2080)) + ((g1896) & (!g2041) & (g2068) & (g1904) & (g2043) & (g2080)) + ((g1896) & (g2041) & (!g2068) & (!g1904) & (g2043) & (g2080)) + ((g1896) & (g2041) & (!g2068) & (g1904) & (!g2043) & (g2080)) + ((g1896) & (g2041) & (!g2068) & (g1904) & (g2043) & (g2080)) + ((g1896) & (g2041) & (g2068) & (!g1904) & (!g2043) & (g2080)) + ((g1896) & (g2041) & (g2068) & (!g1904) & (g2043) & (!g2080)) + ((g1896) & (g2041) & (g2068) & (!g1904) & (g2043) & (g2080)) + ((g1896) & (g2041) & (g2068) & (g1904) & (!g2043) & (!g2080)) + ((g1896) & (g2041) & (g2068) & (g1904) & (!g2043) & (g2080)) + ((g1896) & (g2041) & (g2068) & (g1904) & (g2043) & (!g2080)) + ((g1896) & (g2041) & (g2068) & (g1904) & (g2043) & (g2080)));
	assign g3847 = (((!g2203) & (g2205)) + ((g2203) & (!g2205)));
	assign g3848 = (((!g2123) & (!g2150) & (g2125) & (g2162) & (g3846) & (g3847)) + ((!g2123) & (g2150) & (!g2125) & (g2162) & (!g3846) & (g3847)) + ((!g2123) & (g2150) & (!g2125) & (g2162) & (g3846) & (g3847)) + ((!g2123) & (g2150) & (g2125) & (!g2162) & (g3846) & (g3847)) + ((!g2123) & (g2150) & (g2125) & (g2162) & (!g3846) & (g3847)) + ((!g2123) & (g2150) & (g2125) & (g2162) & (g3846) & (g3847)) + ((g2123) & (!g2150) & (!g2125) & (g2162) & (g3846) & (g3847)) + ((g2123) & (!g2150) & (g2125) & (g2162) & (!g3846) & (g3847)) + ((g2123) & (!g2150) & (g2125) & (g2162) & (g3846) & (g3847)) + ((g2123) & (g2150) & (!g2125) & (!g2162) & (g3846) & (g3847)) + ((g2123) & (g2150) & (!g2125) & (g2162) & (!g3846) & (g3847)) + ((g2123) & (g2150) & (!g2125) & (g2162) & (g3846) & (g3847)) + ((g2123) & (g2150) & (g2125) & (!g2162) & (!g3846) & (g3847)) + ((g2123) & (g2150) & (g2125) & (!g2162) & (g3846) & (g3847)) + ((g2123) & (g2150) & (g2125) & (g2162) & (!g3846) & (g3847)) + ((g2123) & (g2150) & (g2125) & (g2162) & (g3846) & (g3847)));
	assign g3849 = (((g2203) & (g2205)));
	assign g3850 = (((!g2230) & (!g2286) & (g2242) & (g2288) & (!g3848) & (g3849)) + ((!g2230) & (!g2286) & (g2242) & (g2288) & (g3848) & (!g3849)) + ((!g2230) & (!g2286) & (g2242) & (g2288) & (g3848) & (g3849)) + ((!g2230) & (g2286) & (!g2242) & (g2288) & (!g3848) & (!g3849)) + ((!g2230) & (g2286) & (!g2242) & (g2288) & (!g3848) & (g3849)) + ((!g2230) & (g2286) & (!g2242) & (g2288) & (g3848) & (!g3849)) + ((!g2230) & (g2286) & (!g2242) & (g2288) & (g3848) & (g3849)) + ((!g2230) & (g2286) & (g2242) & (!g2288) & (!g3848) & (g3849)) + ((!g2230) & (g2286) & (g2242) & (!g2288) & (g3848) & (!g3849)) + ((!g2230) & (g2286) & (g2242) & (!g2288) & (g3848) & (g3849)) + ((!g2230) & (g2286) & (g2242) & (g2288) & (!g3848) & (!g3849)) + ((!g2230) & (g2286) & (g2242) & (g2288) & (!g3848) & (g3849)) + ((!g2230) & (g2286) & (g2242) & (g2288) & (g3848) & (!g3849)) + ((!g2230) & (g2286) & (g2242) & (g2288) & (g3848) & (g3849)) + ((g2230) & (!g2286) & (!g2242) & (g2288) & (!g3848) & (g3849)) + ((g2230) & (!g2286) & (!g2242) & (g2288) & (g3848) & (!g3849)) + ((g2230) & (!g2286) & (!g2242) & (g2288) & (g3848) & (g3849)) + ((g2230) & (!g2286) & (g2242) & (g2288) & (!g3848) & (!g3849)) + ((g2230) & (!g2286) & (g2242) & (g2288) & (!g3848) & (g3849)) + ((g2230) & (!g2286) & (g2242) & (g2288) & (g3848) & (!g3849)) + ((g2230) & (!g2286) & (g2242) & (g2288) & (g3848) & (g3849)) + ((g2230) & (g2286) & (!g2242) & (!g2288) & (!g3848) & (g3849)) + ((g2230) & (g2286) & (!g2242) & (!g2288) & (g3848) & (!g3849)) + ((g2230) & (g2286) & (!g2242) & (!g2288) & (g3848) & (g3849)) + ((g2230) & (g2286) & (!g2242) & (g2288) & (!g3848) & (!g3849)) + ((g2230) & (g2286) & (!g2242) & (g2288) & (!g3848) & (g3849)) + ((g2230) & (g2286) & (!g2242) & (g2288) & (g3848) & (!g3849)) + ((g2230) & (g2286) & (!g2242) & (g2288) & (g3848) & (g3849)) + ((g2230) & (g2286) & (g2242) & (!g2288) & (!g3848) & (!g3849)) + ((g2230) & (g2286) & (g2242) & (!g2288) & (!g3848) & (g3849)) + ((g2230) & (g2286) & (g2242) & (!g2288) & (g3848) & (!g3849)) + ((g2230) & (g2286) & (g2242) & (!g2288) & (g3848) & (g3849)) + ((g2230) & (g2286) & (g2242) & (g2288) & (!g3848) & (!g3849)) + ((g2230) & (g2286) & (g2242) & (g2288) & (!g3848) & (g3849)) + ((g2230) & (g2286) & (g2242) & (g2288) & (g3848) & (!g3849)) + ((g2230) & (g2286) & (g2242) & (g2288) & (g3848) & (g3849)));
	assign g3851 = (((!g2396) & (g2408)) + ((g2396) & (!g2408)));
	assign g3852 = (((!g2317) & (!g2369) & (g2329) & (g2371) & (g3850) & (g3851)) + ((!g2317) & (g2369) & (!g2329) & (g2371) & (!g3850) & (g3851)) + ((!g2317) & (g2369) & (!g2329) & (g2371) & (g3850) & (g3851)) + ((!g2317) & (g2369) & (g2329) & (!g2371) & (g3850) & (g3851)) + ((!g2317) & (g2369) & (g2329) & (g2371) & (!g3850) & (g3851)) + ((!g2317) & (g2369) & (g2329) & (g2371) & (g3850) & (g3851)) + ((g2317) & (!g2369) & (!g2329) & (g2371) & (g3850) & (g3851)) + ((g2317) & (!g2369) & (g2329) & (g2371) & (!g3850) & (g3851)) + ((g2317) & (!g2369) & (g2329) & (g2371) & (g3850) & (g3851)) + ((g2317) & (g2369) & (!g2329) & (!g2371) & (g3850) & (g3851)) + ((g2317) & (g2369) & (!g2329) & (g2371) & (!g3850) & (g3851)) + ((g2317) & (g2369) & (!g2329) & (g2371) & (g3850) & (g3851)) + ((g2317) & (g2369) & (g2329) & (!g2371) & (!g3850) & (g3851)) + ((g2317) & (g2369) & (g2329) & (!g2371) & (g3850) & (g3851)) + ((g2317) & (g2369) & (g2329) & (g2371) & (!g3850) & (g3851)) + ((g2317) & (g2369) & (g2329) & (g2371) & (g3850) & (g3851)));
	assign g3853 = (((g2396) & (g2408)));
	assign g3854 = (((!g2497) & (!g2531) & (g2503) & (g2539) & (!g3852) & (g3853)) + ((!g2497) & (!g2531) & (g2503) & (g2539) & (g3852) & (!g3853)) + ((!g2497) & (!g2531) & (g2503) & (g2539) & (g3852) & (g3853)) + ((!g2497) & (g2531) & (!g2503) & (g2539) & (!g3852) & (!g3853)) + ((!g2497) & (g2531) & (!g2503) & (g2539) & (!g3852) & (g3853)) + ((!g2497) & (g2531) & (!g2503) & (g2539) & (g3852) & (!g3853)) + ((!g2497) & (g2531) & (!g2503) & (g2539) & (g3852) & (g3853)) + ((!g2497) & (g2531) & (g2503) & (!g2539) & (!g3852) & (g3853)) + ((!g2497) & (g2531) & (g2503) & (!g2539) & (g3852) & (!g3853)) + ((!g2497) & (g2531) & (g2503) & (!g2539) & (g3852) & (g3853)) + ((!g2497) & (g2531) & (g2503) & (g2539) & (!g3852) & (!g3853)) + ((!g2497) & (g2531) & (g2503) & (g2539) & (!g3852) & (g3853)) + ((!g2497) & (g2531) & (g2503) & (g2539) & (g3852) & (!g3853)) + ((!g2497) & (g2531) & (g2503) & (g2539) & (g3852) & (g3853)) + ((g2497) & (!g2531) & (!g2503) & (g2539) & (!g3852) & (g3853)) + ((g2497) & (!g2531) & (!g2503) & (g2539) & (g3852) & (!g3853)) + ((g2497) & (!g2531) & (!g2503) & (g2539) & (g3852) & (g3853)) + ((g2497) & (!g2531) & (g2503) & (g2539) & (!g3852) & (!g3853)) + ((g2497) & (!g2531) & (g2503) & (g2539) & (!g3852) & (g3853)) + ((g2497) & (!g2531) & (g2503) & (g2539) & (g3852) & (!g3853)) + ((g2497) & (!g2531) & (g2503) & (g2539) & (g3852) & (g3853)) + ((g2497) & (g2531) & (!g2503) & (!g2539) & (!g3852) & (g3853)) + ((g2497) & (g2531) & (!g2503) & (!g2539) & (g3852) & (!g3853)) + ((g2497) & (g2531) & (!g2503) & (!g2539) & (g3852) & (g3853)) + ((g2497) & (g2531) & (!g2503) & (g2539) & (!g3852) & (!g3853)) + ((g2497) & (g2531) & (!g2503) & (g2539) & (!g3852) & (g3853)) + ((g2497) & (g2531) & (!g2503) & (g2539) & (g3852) & (!g3853)) + ((g2497) & (g2531) & (!g2503) & (g2539) & (g3852) & (g3853)) + ((g2497) & (g2531) & (g2503) & (!g2539) & (!g3852) & (!g3853)) + ((g2497) & (g2531) & (g2503) & (!g2539) & (!g3852) & (g3853)) + ((g2497) & (g2531) & (g2503) & (!g2539) & (g3852) & (!g3853)) + ((g2497) & (g2531) & (g2503) & (!g2539) & (g3852) & (g3853)) + ((g2497) & (g2531) & (g2503) & (g2539) & (!g3852) & (!g3853)) + ((g2497) & (g2531) & (g2503) & (g2539) & (!g3852) & (g3853)) + ((g2497) & (g2531) & (g2503) & (g2539) & (g3852) & (!g3853)) + ((g2497) & (g2531) & (g2503) & (g2539) & (g3852) & (g3853)));
	assign g3855 = (((!g2589) & (g2592) & (g3854)) + ((g2589) & (!g2592) & (g3854)) + ((g2589) & (g2592) & (!g3854)) + ((g2589) & (g2592) & (g3854)));
	assign g3856 = (((!g1908) & (!g2030) & (g2085) & (!g1910) & (!g2038) & (g2088)) + ((!g1908) & (!g2030) & (g2085) & (!g1910) & (g2038) & (g2088)) + ((!g1908) & (!g2030) & (g2085) & (g1910) & (!g2038) & (g2088)) + ((!g1908) & (!g2030) & (g2085) & (g1910) & (g2038) & (g2088)) + ((!g1908) & (g2030) & (!g2085) & (!g1910) & (g2038) & (g2088)) + ((!g1908) & (g2030) & (!g2085) & (g1910) & (g2038) & (g2088)) + ((!g1908) & (g2030) & (g2085) & (!g1910) & (!g2038) & (g2088)) + ((!g1908) & (g2030) & (g2085) & (!g1910) & (g2038) & (!g2088)) + ((!g1908) & (g2030) & (g2085) & (!g1910) & (g2038) & (g2088)) + ((!g1908) & (g2030) & (g2085) & (g1910) & (!g2038) & (g2088)) + ((!g1908) & (g2030) & (g2085) & (g1910) & (g2038) & (!g2088)) + ((!g1908) & (g2030) & (g2085) & (g1910) & (g2038) & (g2088)) + ((g1908) & (!g2030) & (!g2085) & (g1910) & (g2038) & (g2088)) + ((g1908) & (!g2030) & (g2085) & (!g1910) & (!g2038) & (g2088)) + ((g1908) & (!g2030) & (g2085) & (!g1910) & (g2038) & (g2088)) + ((g1908) & (!g2030) & (g2085) & (g1910) & (!g2038) & (g2088)) + ((g1908) & (!g2030) & (g2085) & (g1910) & (g2038) & (!g2088)) + ((g1908) & (!g2030) & (g2085) & (g1910) & (g2038) & (g2088)) + ((g1908) & (g2030) & (!g2085) & (!g1910) & (g2038) & (g2088)) + ((g1908) & (g2030) & (!g2085) & (g1910) & (!g2038) & (g2088)) + ((g1908) & (g2030) & (!g2085) & (g1910) & (g2038) & (g2088)) + ((g1908) & (g2030) & (g2085) & (!g1910) & (!g2038) & (g2088)) + ((g1908) & (g2030) & (g2085) & (!g1910) & (g2038) & (!g2088)) + ((g1908) & (g2030) & (g2085) & (!g1910) & (g2038) & (g2088)) + ((g1908) & (g2030) & (g2085) & (g1910) & (!g2038) & (!g2088)) + ((g1908) & (g2030) & (g2085) & (g1910) & (!g2038) & (g2088)) + ((g1908) & (g2030) & (g2085) & (g1910) & (g2038) & (!g2088)) + ((g1908) & (g2030) & (g2085) & (g1910) & (g2038) & (g2088)));
	assign g3857 = (((!g2192) & (g2200)) + ((g2192) & (!g2200)));
	assign g3858 = (((!g2112) & (!g2167) & (g2120) & (g2170) & (g3856) & (g3857)) + ((!g2112) & (g2167) & (!g2120) & (g2170) & (!g3856) & (g3857)) + ((!g2112) & (g2167) & (!g2120) & (g2170) & (g3856) & (g3857)) + ((!g2112) & (g2167) & (g2120) & (!g2170) & (g3856) & (g3857)) + ((!g2112) & (g2167) & (g2120) & (g2170) & (!g3856) & (g3857)) + ((!g2112) & (g2167) & (g2120) & (g2170) & (g3856) & (g3857)) + ((g2112) & (!g2167) & (!g2120) & (g2170) & (g3856) & (g3857)) + ((g2112) & (!g2167) & (g2120) & (g2170) & (!g3856) & (g3857)) + ((g2112) & (!g2167) & (g2120) & (g2170) & (g3856) & (g3857)) + ((g2112) & (g2167) & (!g2120) & (!g2170) & (g3856) & (g3857)) + ((g2112) & (g2167) & (!g2120) & (g2170) & (!g3856) & (g3857)) + ((g2112) & (g2167) & (!g2120) & (g2170) & (g3856) & (g3857)) + ((g2112) & (g2167) & (g2120) & (!g2170) & (!g3856) & (g3857)) + ((g2112) & (g2167) & (g2120) & (!g2170) & (g3856) & (g3857)) + ((g2112) & (g2167) & (g2120) & (g2170) & (!g3856) & (g3857)) + ((g2112) & (g2167) & (g2120) & (g2170) & (g3856) & (g3857)));
	assign g3859 = (((g2192) & (g2200)));
	assign g3860 = (((!g2247) & (!g2275) & (!g2250) & (!g2283) & (!g3858) & (!g3859)) + ((!g2247) & (!g2275) & (!g2250) & (!g2283) & (!g3858) & (g3859)) + ((!g2247) & (!g2275) & (!g2250) & (!g2283) & (g3858) & (!g3859)) + ((!g2247) & (!g2275) & (!g2250) & (!g2283) & (g3858) & (g3859)) + ((!g2247) & (!g2275) & (!g2250) & (g2283) & (!g3858) & (!g3859)) + ((!g2247) & (!g2275) & (!g2250) & (g2283) & (!g3858) & (g3859)) + ((!g2247) & (!g2275) & (!g2250) & (g2283) & (g3858) & (!g3859)) + ((!g2247) & (!g2275) & (!g2250) & (g2283) & (g3858) & (g3859)) + ((!g2247) & (!g2275) & (g2250) & (!g2283) & (!g3858) & (!g3859)) + ((!g2247) & (!g2275) & (g2250) & (!g2283) & (!g3858) & (g3859)) + ((!g2247) & (!g2275) & (g2250) & (!g2283) & (g3858) & (!g3859)) + ((!g2247) & (!g2275) & (g2250) & (!g2283) & (g3858) & (g3859)) + ((!g2247) & (!g2275) & (g2250) & (g2283) & (!g3858) & (!g3859)) + ((!g2247) & (g2275) & (!g2250) & (!g2283) & (!g3858) & (!g3859)) + ((!g2247) & (g2275) & (!g2250) & (!g2283) & (!g3858) & (g3859)) + ((!g2247) & (g2275) & (!g2250) & (!g2283) & (g3858) & (!g3859)) + ((!g2247) & (g2275) & (!g2250) & (!g2283) & (g3858) & (g3859)) + ((!g2247) & (g2275) & (g2250) & (!g2283) & (!g3858) & (!g3859)) + ((g2247) & (!g2275) & (!g2250) & (!g2283) & (!g3858) & (!g3859)) + ((g2247) & (!g2275) & (!g2250) & (!g2283) & (!g3858) & (g3859)) + ((g2247) & (!g2275) & (!g2250) & (!g2283) & (g3858) & (!g3859)) + ((g2247) & (!g2275) & (!g2250) & (!g2283) & (g3858) & (g3859)) + ((g2247) & (!g2275) & (!g2250) & (g2283) & (!g3858) & (!g3859)) + ((g2247) & (!g2275) & (g2250) & (!g2283) & (!g3858) & (!g3859)) + ((g2247) & (!g2275) & (g2250) & (!g2283) & (!g3858) & (g3859)) + ((g2247) & (!g2275) & (g2250) & (!g2283) & (g3858) & (!g3859)) + ((g2247) & (!g2275) & (g2250) & (!g2283) & (g3858) & (g3859)) + ((g2247) & (g2275) & (!g2250) & (!g2283) & (!g3858) & (!g3859)));
	assign g3861 = (((!g2334) & (!g2358) & (g2337) & (g2366) & (!g3860)) + ((!g2334) & (g2358) & (!g2337) & (g2366) & (!g3860)) + ((!g2334) & (g2358) & (!g2337) & (g2366) & (g3860)) + ((!g2334) & (g2358) & (g2337) & (!g2366) & (!g3860)) + ((!g2334) & (g2358) & (g2337) & (g2366) & (!g3860)) + ((!g2334) & (g2358) & (g2337) & (g2366) & (g3860)) + ((g2334) & (!g2358) & (!g2337) & (g2366) & (!g3860)) + ((g2334) & (!g2358) & (g2337) & (g2366) & (!g3860)) + ((g2334) & (!g2358) & (g2337) & (g2366) & (g3860)) + ((g2334) & (g2358) & (!g2337) & (!g2366) & (!g3860)) + ((g2334) & (g2358) & (!g2337) & (g2366) & (!g3860)) + ((g2334) & (g2358) & (!g2337) & (g2366) & (g3860)) + ((g2334) & (g2358) & (g2337) & (!g2366) & (!g3860)) + ((g2334) & (g2358) & (g2337) & (!g2366) & (g3860)) + ((g2334) & (g2358) & (g2337) & (g2366) & (!g3860)) + ((g2334) & (g2358) & (g2337) & (g2366) & (g3860)));
	assign g3862 = (((!g2542) & (g2544)) + ((g2542) & (!g2544)));
	assign g3863 = (((!g2413) & (!g2462) & (g2416) & (g2486) & (g3861) & (g3862)) + ((!g2413) & (g2462) & (!g2416) & (g2486) & (!g3861) & (g3862)) + ((!g2413) & (g2462) & (!g2416) & (g2486) & (g3861) & (g3862)) + ((!g2413) & (g2462) & (g2416) & (!g2486) & (g3861) & (g3862)) + ((!g2413) & (g2462) & (g2416) & (g2486) & (!g3861) & (g3862)) + ((!g2413) & (g2462) & (g2416) & (g2486) & (g3861) & (g3862)) + ((g2413) & (!g2462) & (!g2416) & (g2486) & (g3861) & (g3862)) + ((g2413) & (!g2462) & (g2416) & (g2486) & (!g3861) & (g3862)) + ((g2413) & (!g2462) & (g2416) & (g2486) & (g3861) & (g3862)) + ((g2413) & (g2462) & (!g2416) & (!g2486) & (g3861) & (g3862)) + ((g2413) & (g2462) & (!g2416) & (g2486) & (!g3861) & (g3862)) + ((g2413) & (g2462) & (!g2416) & (g2486) & (g3861) & (g3862)) + ((g2413) & (g2462) & (g2416) & (!g2486) & (!g3861) & (g3862)) + ((g2413) & (g2462) & (g2416) & (!g2486) & (g3861) & (g3862)) + ((g2413) & (g2462) & (g2416) & (g2486) & (!g3861) & (g3862)) + ((g2413) & (g2462) & (g2416) & (g2486) & (g3861) & (g3862)));
	assign g3864 = (((g2542) & (g2544)));
	assign g3865 = (((!g3863) & (!g3864)));
	assign g3866 = (((!g2572) & (!g2637) & (!g2584) & (g2640) & (!g3865)) + ((!g2572) & (!g2637) & (!g2584) & (g2640) & (g3865)) + ((!g2572) & (!g2637) & (g2584) & (!g2640) & (!g3865)) + ((!g2572) & (!g2637) & (g2584) & (g2640) & (g3865)) + ((!g2572) & (g2637) & (!g2584) & (!g2640) & (!g3865)) + ((!g2572) & (g2637) & (!g2584) & (!g2640) & (g3865)) + ((!g2572) & (g2637) & (g2584) & (!g2640) & (g3865)) + ((!g2572) & (g2637) & (g2584) & (g2640) & (!g3865)) + ((g2572) & (!g2637) & (!g2584) & (!g2640) & (!g3865)) + ((g2572) & (!g2637) & (!g2584) & (g2640) & (g3865)) + ((g2572) & (!g2637) & (g2584) & (!g2640) & (!g3865)) + ((g2572) & (!g2637) & (g2584) & (!g2640) & (g3865)) + ((g2572) & (g2637) & (!g2584) & (!g2640) & (g3865)) + ((g2572) & (g2637) & (!g2584) & (g2640) & (!g3865)) + ((g2572) & (g2637) & (g2584) & (g2640) & (!g3865)) + ((g2572) & (g2637) & (g2584) & (g2640) & (g3865)));
	assign g3867 = (((g831) & (!g1914) & (!g1921) & (!g1922) & (!g1930) & (!g1933)) + ((g831) & (!g1914) & (!g1921) & (!g1922) & (!g1930) & (g1933)) + ((g831) & (!g1914) & (!g1921) & (!g1922) & (g1930) & (!g1933)) + ((g831) & (!g1914) & (!g1921) & (!g1922) & (g1930) & (g1933)) + ((g831) & (!g1914) & (!g1921) & (g1922) & (!g1930) & (!g1933)) + ((g831) & (!g1914) & (!g1921) & (g1922) & (!g1930) & (g1933)) + ((g831) & (!g1914) & (!g1921) & (g1922) & (g1930) & (!g1933)) + ((g831) & (!g1914) & (!g1921) & (g1922) & (g1930) & (g1933)) + ((g831) & (!g1914) & (g1921) & (!g1922) & (!g1930) & (!g1933)) + ((g831) & (!g1914) & (g1921) & (!g1922) & (!g1930) & (g1933)) + ((g831) & (!g1914) & (g1921) & (!g1922) & (g1930) & (!g1933)) + ((g831) & (!g1914) & (g1921) & (!g1922) & (g1930) & (g1933)) + ((g831) & (!g1914) & (g1921) & (g1922) & (!g1930) & (!g1933)) + ((g831) & (!g1914) & (g1921) & (g1922) & (!g1930) & (g1933)) + ((g831) & (!g1914) & (g1921) & (g1922) & (g1930) & (!g1933)) + ((g831) & (!g1914) & (g1921) & (g1922) & (g1930) & (g1933)) + ((g831) & (g1914) & (!g1921) & (!g1922) & (!g1930) & (!g1933)) + ((g831) & (g1914) & (!g1921) & (!g1922) & (!g1930) & (g1933)) + ((g831) & (g1914) & (!g1921) & (!g1922) & (g1930) & (!g1933)) + ((g831) & (g1914) & (!g1921) & (!g1922) & (g1930) & (g1933)) + ((g831) & (g1914) & (!g1921) & (g1922) & (!g1930) & (!g1933)) + ((g831) & (g1914) & (!g1921) & (g1922) & (!g1930) & (g1933)) + ((g831) & (g1914) & (!g1921) & (g1922) & (g1930) & (!g1933)) + ((g831) & (g1914) & (!g1921) & (g1922) & (g1930) & (g1933)) + ((g831) & (g1914) & (g1921) & (!g1922) & (!g1930) & (!g1933)) + ((g831) & (g1914) & (g1921) & (!g1922) & (!g1930) & (g1933)) + ((g831) & (g1914) & (g1921) & (!g1922) & (g1930) & (!g1933)) + ((g831) & (g1914) & (g1921) & (!g1922) & (g1930) & (g1933)) + ((g831) & (g1914) & (g1921) & (g1922) & (g1930) & (g1933)));
	assign g3868 = (((!g1914) & (g1920) & (g1922) & (g3867)) + ((g1914) & (!g1920) & (!g1922) & (g3867)) + ((g1914) & (!g1920) & (g1922) & (g3867)) + ((g1914) & (g1920) & (!g1922) & (g3867)));
	assign g3869 = (((!reset) & (!g827) & (g830)));
	assign g3870 = (((g1914) & (g1918) & (g1920) & (g1922)));
	assign g3871 = (((g1917) & (g3870)));
	assign g3872 = (((!g1915) & (g1916) & (g3867) & (g3871)) + ((g1915) & (!g1916) & (g3867) & (!g3871)) + ((g1915) & (!g1916) & (g3867) & (g3871)) + ((g1915) & (g1916) & (g3867) & (!g3871)));
	assign g3873 = (((!g1916) & (g3867) & (g3871)) + ((g1916) & (g3867) & (!g3871)));
	assign g3874 = (((!g1917) & (g3867) & (g3870)) + ((g1917) & (g3867) & (!g3870)));
	assign g3875 = (((!g1914) & (g1918) & (!g1920) & (!g1922) & (g3867)) + ((!g1914) & (g1918) & (!g1920) & (g1922) & (g3867)) + ((!g1914) & (g1918) & (g1920) & (!g1922) & (g3867)) + ((!g1914) & (g1918) & (g1920) & (g1922) & (g3867)) + ((g1914) & (!g1918) & (g1920) & (g1922) & (g3867)) + ((g1914) & (g1918) & (!g1920) & (!g1922) & (g3867)) + ((g1914) & (g1918) & (!g1920) & (g1922) & (g3867)) + ((g1914) & (g1918) & (g1920) & (!g1922) & (g3867)));
	assign g3876 = (((!g1915) & (!g1916) & (g1919) & (g3867) & (!g3871)) + ((!g1915) & (!g1916) & (g1919) & (g3867) & (g3871)) + ((!g1915) & (g1916) & (g1919) & (g3867) & (!g3871)) + ((!g1915) & (g1916) & (g1919) & (g3867) & (g3871)) + ((g1915) & (!g1916) & (g1919) & (g3867) & (!g3871)) + ((g1915) & (!g1916) & (g1919) & (g3867) & (g3871)) + ((g1915) & (g1916) & (!g1919) & (g3867) & (g3871)) + ((g1915) & (g1916) & (g1919) & (g3867) & (!g3871)));
	assign g3877 = (((!g1920) & (g3867)));
	assign g3878 = (((!g1920) & (g1922) & (g3867)) + ((g1920) & (!g1922) & (g3867)));
	assign g3879 = (((g831) & (!g1924) & (g1925) & (g1931) & (g1932)) + ((g831) & (g1924) & (!g1925) & (!g1931) & (!g1932)) + ((g831) & (g1924) & (!g1925) & (!g1931) & (g1932)) + ((g831) & (g1924) & (!g1925) & (g1931) & (!g1932)) + ((g831) & (g1924) & (!g1925) & (g1931) & (g1932)) + ((g831) & (g1924) & (g1925) & (!g1931) & (!g1932)) + ((g831) & (g1924) & (g1925) & (!g1931) & (g1932)) + ((g831) & (g1924) & (g1925) & (g1931) & (!g1932)));
	assign g3880 = (((!reset) & (!g827) & (!g830) & (!g3867)) + ((!reset) & (!g827) & (!g830) & (g3867)) + ((!reset) & (!g827) & (g830) & (g3867)) + ((!reset) & (g827) & (!g830) & (!g3867)) + ((!reset) & (g827) & (!g830) & (g3867)) + ((!reset) & (g827) & (g830) & (!g3867)) + ((!reset) & (g827) & (g830) & (g3867)) + ((reset) & (!g827) & (!g830) & (!g3867)) + ((reset) & (!g827) & (!g830) & (g3867)) + ((reset) & (!g827) & (g830) & (!g3867)) + ((reset) & (!g827) & (g830) & (g3867)) + ((reset) & (g827) & (!g830) & (!g3867)) + ((reset) & (g827) & (!g830) & (g3867)) + ((reset) & (g827) & (g830) & (!g3867)) + ((reset) & (g827) & (g830) & (g3867)));
	assign g3881 = (((g831) & (!g1925) & (g1932)) + ((g831) & (g1925) & (!g1932)));
	assign g3882 = (((g1924) & (g1925) & (g1931) & (g1932)));
	assign g3883 = (((g1929) & (g3882)));
	assign g3884 = (((g831) & (!g1926) & (g1927) & (g1928) & (g3883)) + ((g831) & (g1926) & (!g1927) & (!g1928) & (!g3883)) + ((g831) & (g1926) & (!g1927) & (!g1928) & (g3883)) + ((g831) & (g1926) & (!g1927) & (g1928) & (!g3883)) + ((g831) & (g1926) & (!g1927) & (g1928) & (g3883)) + ((g831) & (g1926) & (g1927) & (!g1928) & (!g3883)) + ((g831) & (g1926) & (g1927) & (!g1928) & (g3883)) + ((g831) & (g1926) & (g1927) & (g1928) & (!g3883)));
	assign g3885 = (((g831) & (!g1927) & (g1928) & (g3883)) + ((g831) & (g1927) & (!g1928) & (!g3883)) + ((g831) & (g1927) & (!g1928) & (g3883)) + ((g831) & (g1927) & (g1928) & (!g3883)));
	assign g3886 = (((g831) & (!g1928) & (g3883)) + ((g831) & (g1928) & (!g3883)));
	assign g3887 = (((g831) & (!g1929) & (g3882)) + ((g831) & (g1929) & (!g3882)));
	assign g3888 = (((g831) & (!g1925) & (g1931) & (!g1932)) + ((g831) & (!g1925) & (g1931) & (g1932)) + ((g831) & (g1925) & (!g1931) & (g1932)) + ((g831) & (g1925) & (g1931) & (!g1932)));
	assign g3889 = (((g831) & (!g1932)));
	assign g3890 = (((!g34) & (!g35) & (g36) & (!g1935)) + ((!g34) & (!g35) & (g36) & (g1935)) + ((!g34) & (g35) & (g36) & (!g1935)) + ((!g34) & (g35) & (g36) & (g1935)) + ((g34) & (g35) & (g36) & (g1935)));
	assign g3891 = (((!g1610) & (!g3515) & (g3031)) + ((g1610) & (!g3515) & (!g3031)) + ((g1610) & (!g3515) & (g3031)) + ((g1610) & (g3515) & (g3031)));
	assign g3892 = (((g1914) & (!g1644) & (!g3084) & (g3891)) + ((g1914) & (!g1644) & (g3084) & (!g3891)) + ((g1914) & (g1644) & (!g3084) & (!g3891)) + ((g1914) & (g1644) & (g3084) & (g3891)));
	assign g3893 = (((!g3038) & (g3061) & (!g3532)) + ((g3038) & (!g3061) & (!g3532)) + ((g3038) & (g3061) & (!g3532)) + ((g3038) & (g3061) & (g3532)));
	assign g3894 = (((!g1914) & (!g3082) & (!g3078) & (g3893)) + ((!g1914) & (!g3082) & (g3078) & (!g3893)) + ((!g1914) & (g3082) & (!g3078) & (!g3893)) + ((!g1914) & (g3082) & (g3078) & (g3893)));
	assign g3895 = (((!g830) & (!g1939) & (!g3892) & (!g3894) & (key[33])) + ((!g830) & (!g1939) & (!g3892) & (g3894) & (key[33])) + ((!g830) & (!g1939) & (g3892) & (!g3894) & (key[33])) + ((!g830) & (!g1939) & (g3892) & (g3894) & (key[33])) + ((!g830) & (g1939) & (!g3892) & (!g3894) & (key[33])) + ((!g830) & (g1939) & (!g3892) & (g3894) & (key[33])) + ((!g830) & (g1939) & (g3892) & (!g3894) & (key[33])) + ((!g830) & (g1939) & (g3892) & (g3894) & (key[33])) + ((g830) & (!g1939) & (!g3892) & (g3894) & (!key[33])) + ((g830) & (!g1939) & (!g3892) & (g3894) & (key[33])) + ((g830) & (!g1939) & (g3892) & (!g3894) & (!key[33])) + ((g830) & (!g1939) & (g3892) & (!g3894) & (key[33])) + ((g830) & (!g1939) & (g3892) & (g3894) & (!key[33])) + ((g830) & (!g1939) & (g3892) & (g3894) & (key[33])) + ((g830) & (g1939) & (!g3892) & (!g3894) & (!key[33])) + ((g830) & (g1939) & (!g3892) & (!g3894) & (key[33])));
	assign g3896 = (((!g2210) & (!g2256) & (!g2838) & (g2891) & (!g3758)) + ((!g2210) & (!g2256) & (!g2838) & (g2891) & (g3758)) + ((!g2210) & (!g2256) & (g2838) & (!g2891) & (g3758)) + ((!g2210) & (!g2256) & (g2838) & (g2891) & (!g3758)) + ((!g2210) & (g2256) & (!g2838) & (!g2891) & (!g3758)) + ((!g2210) & (g2256) & (!g2838) & (!g2891) & (g3758)) + ((!g2210) & (g2256) & (g2838) & (!g2891) & (!g3758)) + ((!g2210) & (g2256) & (g2838) & (g2891) & (g3758)) + ((g2210) & (!g2256) & (!g2838) & (!g2891) & (g3758)) + ((g2210) & (!g2256) & (!g2838) & (g2891) & (!g3758)) + ((g2210) & (!g2256) & (g2838) & (!g2891) & (!g3758)) + ((g2210) & (!g2256) & (g2838) & (!g2891) & (g3758)) + ((g2210) & (g2256) & (!g2838) & (!g2891) & (!g3758)) + ((g2210) & (g2256) & (!g2838) & (g2891) & (g3758)) + ((g2210) & (g2256) & (g2838) & (g2891) & (!g3758)) + ((g2210) & (g2256) & (g2838) & (g2891) & (g3758)));
	assign g3897 = (((!g3142) & (g3119)) + ((g3142) & (!g3119)));
	assign g3898 = (((!g3044) & (!g3067) & (g3097) & (!g3774) & (g3093) & (g3897)) + ((!g3044) & (!g3067) & (g3097) & (g3774) & (g3093) & (g3897)) + ((!g3044) & (g3067) & (!g3097) & (!g3774) & (g3093) & (g3897)) + ((!g3044) & (g3067) & (g3097) & (!g3774) & (!g3093) & (g3897)) + ((!g3044) & (g3067) & (g3097) & (!g3774) & (g3093) & (g3897)) + ((!g3044) & (g3067) & (g3097) & (g3774) & (g3093) & (g3897)) + ((g3044) & (!g3067) & (!g3097) & (!g3774) & (g3093) & (g3897)) + ((g3044) & (!g3067) & (g3097) & (!g3774) & (!g3093) & (g3897)) + ((g3044) & (!g3067) & (g3097) & (!g3774) & (g3093) & (g3897)) + ((g3044) & (!g3067) & (g3097) & (g3774) & (g3093) & (g3897)) + ((g3044) & (g3067) & (!g3097) & (!g3774) & (g3093) & (g3897)) + ((g3044) & (g3067) & (!g3097) & (g3774) & (g3093) & (g3897)) + ((g3044) & (g3067) & (g3097) & (!g3774) & (!g3093) & (g3897)) + ((g3044) & (g3067) & (g3097) & (!g3774) & (g3093) & (g3897)) + ((g3044) & (g3067) & (g3097) & (g3774) & (!g3093) & (g3897)) + ((g3044) & (g3067) & (g3097) & (g3774) & (g3093) & (g3897)));
	assign g3899 = (((g3142) & (g3119)));
	assign g3900 = (((!g3898) & (!g3899) & (!g3168) & (g3172)) + ((!g3898) & (!g3899) & (g3168) & (!g3172)) + ((!g3898) & (g3899) & (!g3168) & (!g3172)) + ((!g3898) & (g3899) & (g3168) & (g3172)) + ((g3898) & (!g3899) & (!g3168) & (!g3172)) + ((g3898) & (!g3899) & (g3168) & (g3172)) + ((g3898) & (g3899) & (!g3168) & (!g3172)) + ((g3898) & (g3899) & (g3168) & (g3172)));
	assign g3901 = (((!g830) & (!g1914) & (!g1940) & (!g3896) & (!g3900) & (key[65])) + ((!g830) & (!g1914) & (!g1940) & (!g3896) & (g3900) & (key[65])) + ((!g830) & (!g1914) & (!g1940) & (g3896) & (!g3900) & (key[65])) + ((!g830) & (!g1914) & (!g1940) & (g3896) & (g3900) & (key[65])) + ((!g830) & (!g1914) & (g1940) & (!g3896) & (!g3900) & (key[65])) + ((!g830) & (!g1914) & (g1940) & (!g3896) & (g3900) & (key[65])) + ((!g830) & (!g1914) & (g1940) & (g3896) & (!g3900) & (key[65])) + ((!g830) & (!g1914) & (g1940) & (g3896) & (g3900) & (key[65])) + ((!g830) & (g1914) & (!g1940) & (!g3896) & (!g3900) & (key[65])) + ((!g830) & (g1914) & (!g1940) & (!g3896) & (g3900) & (key[65])) + ((!g830) & (g1914) & (!g1940) & (g3896) & (!g3900) & (key[65])) + ((!g830) & (g1914) & (!g1940) & (g3896) & (g3900) & (key[65])) + ((!g830) & (g1914) & (g1940) & (!g3896) & (!g3900) & (key[65])) + ((!g830) & (g1914) & (g1940) & (!g3896) & (g3900) & (key[65])) + ((!g830) & (g1914) & (g1940) & (g3896) & (!g3900) & (key[65])) + ((!g830) & (g1914) & (g1940) & (g3896) & (g3900) & (key[65])) + ((g830) & (!g1914) & (!g1940) & (!g3896) & (g3900) & (!key[65])) + ((g830) & (!g1914) & (!g1940) & (!g3896) & (g3900) & (key[65])) + ((g830) & (!g1914) & (!g1940) & (g3896) & (g3900) & (!key[65])) + ((g830) & (!g1914) & (!g1940) & (g3896) & (g3900) & (key[65])) + ((g830) & (!g1914) & (g1940) & (!g3896) & (!g3900) & (!key[65])) + ((g830) & (!g1914) & (g1940) & (!g3896) & (!g3900) & (key[65])) + ((g830) & (!g1914) & (g1940) & (g3896) & (!g3900) & (!key[65])) + ((g830) & (!g1914) & (g1940) & (g3896) & (!g3900) & (key[65])) + ((g830) & (g1914) & (!g1940) & (g3896) & (!g3900) & (!key[65])) + ((g830) & (g1914) & (!g1940) & (g3896) & (!g3900) & (key[65])) + ((g830) & (g1914) & (!g1940) & (g3896) & (g3900) & (!key[65])) + ((g830) & (g1914) & (!g1940) & (g3896) & (g3900) & (key[65])) + ((g830) & (g1914) & (g1940) & (!g3896) & (!g3900) & (!key[65])) + ((g830) & (g1914) & (g1940) & (!g3896) & (!g3900) & (key[65])) + ((g830) & (g1914) & (g1940) & (!g3896) & (g3900) & (!key[65])) + ((g830) & (g1914) & (g1940) & (!g3896) & (g3900) & (key[65])));
	assign g3902 = (((!g1644) & (!g1677) & (!g3084) & (g3106) & (!g3891)) + ((!g1644) & (!g1677) & (!g3084) & (g3106) & (g3891)) + ((!g1644) & (!g1677) & (g3084) & (!g3106) & (g3891)) + ((!g1644) & (!g1677) & (g3084) & (g3106) & (!g3891)) + ((!g1644) & (g1677) & (!g3084) & (!g3106) & (!g3891)) + ((!g1644) & (g1677) & (!g3084) & (!g3106) & (g3891)) + ((!g1644) & (g1677) & (g3084) & (!g3106) & (!g3891)) + ((!g1644) & (g1677) & (g3084) & (g3106) & (g3891)) + ((g1644) & (!g1677) & (!g3084) & (!g3106) & (g3891)) + ((g1644) & (!g1677) & (!g3084) & (g3106) & (!g3891)) + ((g1644) & (!g1677) & (g3084) & (!g3106) & (!g3891)) + ((g1644) & (!g1677) & (g3084) & (!g3106) & (g3891)) + ((g1644) & (g1677) & (!g3084) & (!g3106) & (!g3891)) + ((g1644) & (g1677) & (!g3084) & (g3106) & (g3891)) + ((g1644) & (g1677) & (g3084) & (g3106) & (!g3891)) + ((g1644) & (g1677) & (g3084) & (g3106) & (g3891)));
	assign g3903 = (((!g3082) & (!g3136) & (!g3078) & (g3113) & (!g3893)) + ((!g3082) & (!g3136) & (!g3078) & (g3113) & (g3893)) + ((!g3082) & (!g3136) & (g3078) & (!g3113) & (g3893)) + ((!g3082) & (!g3136) & (g3078) & (g3113) & (!g3893)) + ((!g3082) & (g3136) & (!g3078) & (!g3113) & (!g3893)) + ((!g3082) & (g3136) & (!g3078) & (!g3113) & (g3893)) + ((!g3082) & (g3136) & (g3078) & (!g3113) & (!g3893)) + ((!g3082) & (g3136) & (g3078) & (g3113) & (g3893)) + ((g3082) & (!g3136) & (!g3078) & (!g3113) & (g3893)) + ((g3082) & (!g3136) & (!g3078) & (g3113) & (!g3893)) + ((g3082) & (!g3136) & (g3078) & (!g3113) & (!g3893)) + ((g3082) & (!g3136) & (g3078) & (!g3113) & (g3893)) + ((g3082) & (g3136) & (!g3078) & (!g3113) & (!g3893)) + ((g3082) & (g3136) & (!g3078) & (g3113) & (g3893)) + ((g3082) & (g3136) & (g3078) & (g3113) & (!g3893)) + ((g3082) & (g3136) & (g3078) & (g3113) & (g3893)));
	assign g3904 = (((!g830) & (!g1914) & (!g1941) & (!g3902) & (!g3903) & (key[34])) + ((!g830) & (!g1914) & (!g1941) & (!g3902) & (g3903) & (key[34])) + ((!g830) & (!g1914) & (!g1941) & (g3902) & (!g3903) & (key[34])) + ((!g830) & (!g1914) & (!g1941) & (g3902) & (g3903) & (key[34])) + ((!g830) & (!g1914) & (g1941) & (!g3902) & (!g3903) & (key[34])) + ((!g830) & (!g1914) & (g1941) & (!g3902) & (g3903) & (key[34])) + ((!g830) & (!g1914) & (g1941) & (g3902) & (!g3903) & (key[34])) + ((!g830) & (!g1914) & (g1941) & (g3902) & (g3903) & (key[34])) + ((!g830) & (g1914) & (!g1941) & (!g3902) & (!g3903) & (key[34])) + ((!g830) & (g1914) & (!g1941) & (!g3902) & (g3903) & (key[34])) + ((!g830) & (g1914) & (!g1941) & (g3902) & (!g3903) & (key[34])) + ((!g830) & (g1914) & (!g1941) & (g3902) & (g3903) & (key[34])) + ((!g830) & (g1914) & (g1941) & (!g3902) & (!g3903) & (key[34])) + ((!g830) & (g1914) & (g1941) & (!g3902) & (g3903) & (key[34])) + ((!g830) & (g1914) & (g1941) & (g3902) & (!g3903) & (key[34])) + ((!g830) & (g1914) & (g1941) & (g3902) & (g3903) & (key[34])) + ((g830) & (!g1914) & (!g1941) & (!g3902) & (g3903) & (!key[34])) + ((g830) & (!g1914) & (!g1941) & (!g3902) & (g3903) & (key[34])) + ((g830) & (!g1914) & (!g1941) & (g3902) & (g3903) & (!key[34])) + ((g830) & (!g1914) & (!g1941) & (g3902) & (g3903) & (key[34])) + ((g830) & (!g1914) & (g1941) & (!g3902) & (!g3903) & (!key[34])) + ((g830) & (!g1914) & (g1941) & (!g3902) & (!g3903) & (key[34])) + ((g830) & (!g1914) & (g1941) & (g3902) & (!g3903) & (!key[34])) + ((g830) & (!g1914) & (g1941) & (g3902) & (!g3903) & (key[34])) + ((g830) & (g1914) & (!g1941) & (g3902) & (!g3903) & (!key[34])) + ((g830) & (g1914) & (!g1941) & (g3902) & (!g3903) & (key[34])) + ((g830) & (g1914) & (!g1941) & (g3902) & (g3903) & (!key[34])) + ((g830) & (g1914) & (!g1941) & (g3902) & (g3903) & (key[34])) + ((g830) & (g1914) & (g1941) & (!g3902) & (!g3903) & (!key[34])) + ((g830) & (g1914) & (g1941) & (!g3902) & (!g3903) & (key[34])) + ((g830) & (g1914) & (g1941) & (!g3902) & (g3903) & (!key[34])) + ((g830) & (g1914) & (g1941) & (!g3902) & (g3903) & (key[34])));
	assign g3905 = (((!g2256) & (g2891)) + ((g2256) & (!g2891)));
	assign g3906 = (((!g2177) & (!g2210) & (g2813) & (g2838) & (!g3757) & (g3905)) + ((!g2177) & (g2210) & (!g2813) & (g2838) & (!g3757) & (g3905)) + ((!g2177) & (g2210) & (!g2813) & (g2838) & (g3757) & (g3905)) + ((!g2177) & (g2210) & (g2813) & (!g2838) & (!g3757) & (g3905)) + ((!g2177) & (g2210) & (g2813) & (g2838) & (!g3757) & (g3905)) + ((!g2177) & (g2210) & (g2813) & (g2838) & (g3757) & (g3905)) + ((g2177) & (!g2210) & (!g2813) & (g2838) & (!g3757) & (g3905)) + ((g2177) & (!g2210) & (g2813) & (g2838) & (!g3757) & (g3905)) + ((g2177) & (!g2210) & (g2813) & (g2838) & (g3757) & (g3905)) + ((g2177) & (g2210) & (!g2813) & (!g2838) & (!g3757) & (g3905)) + ((g2177) & (g2210) & (!g2813) & (g2838) & (!g3757) & (g3905)) + ((g2177) & (g2210) & (!g2813) & (g2838) & (g3757) & (g3905)) + ((g2177) & (g2210) & (g2813) & (!g2838) & (!g3757) & (g3905)) + ((g2177) & (g2210) & (g2813) & (!g2838) & (g3757) & (g3905)) + ((g2177) & (g2210) & (g2813) & (g2838) & (!g3757) & (g3905)) + ((g2177) & (g2210) & (g2813) & (g2838) & (g3757) & (g3905)));
	assign g3907 = (((g2256) & (g2891)));
	assign g3908 = (((!g2295) & (!g2916) & (!g3906) & (g3907)) + ((!g2295) & (!g2916) & (g3906) & (!g3907)) + ((!g2295) & (!g2916) & (g3906) & (g3907)) + ((!g2295) & (g2916) & (!g3906) & (!g3907)) + ((g2295) & (!g2916) & (!g3906) & (!g3907)) + ((g2295) & (g2916) & (!g3906) & (g3907)) + ((g2295) & (g2916) & (g3906) & (!g3907)) + ((g2295) & (g2916) & (g3906) & (g3907)));
	assign g3909 = (((!g3898) & (!g3899) & (!g3168) & (!g3172)) + ((!g3898) & (!g3899) & (!g3168) & (g3172)) + ((!g3898) & (!g3899) & (g3168) & (!g3172)) + ((!g3898) & (g3899) & (!g3168) & (!g3172)) + ((g3898) & (!g3899) & (!g3168) & (!g3172)) + ((g3898) & (g3899) & (!g3168) & (!g3172)));
	assign g3910 = (((!g1914) & (!g3213) & (!g3908) & (!g3909) & (!g3190)) + ((!g1914) & (!g3213) & (!g3908) & (g3909) & (g3190)) + ((!g1914) & (!g3213) & (g3908) & (!g3909) & (!g3190)) + ((!g1914) & (!g3213) & (g3908) & (g3909) & (g3190)) + ((!g1914) & (g3213) & (!g3908) & (!g3909) & (g3190)) + ((!g1914) & (g3213) & (!g3908) & (g3909) & (!g3190)) + ((!g1914) & (g3213) & (g3908) & (!g3909) & (g3190)) + ((!g1914) & (g3213) & (g3908) & (g3909) & (!g3190)) + ((g1914) & (!g3213) & (g3908) & (!g3909) & (!g3190)) + ((g1914) & (!g3213) & (g3908) & (!g3909) & (g3190)) + ((g1914) & (!g3213) & (g3908) & (g3909) & (!g3190)) + ((g1914) & (!g3213) & (g3908) & (g3909) & (g3190)) + ((g1914) & (g3213) & (g3908) & (!g3909) & (!g3190)) + ((g1914) & (g3213) & (g3908) & (!g3909) & (g3190)) + ((g1914) & (g3213) & (g3908) & (g3909) & (!g3190)) + ((g1914) & (g3213) & (g3908) & (g3909) & (g3190)));
	assign g3911 = (((!g830) & (!g1942) & (!g3910) & (key[66])) + ((!g830) & (!g1942) & (g3910) & (key[66])) + ((!g830) & (g1942) & (!g3910) & (key[66])) + ((!g830) & (g1942) & (g3910) & (key[66])) + ((g830) & (!g1942) & (g3910) & (!key[66])) + ((g830) & (!g1942) & (g3910) & (key[66])) + ((g830) & (g1942) & (!g3910) & (!key[66])) + ((g830) & (g1942) & (!g3910) & (key[66])));
	assign g3912 = (((!g1677) & (g3106)) + ((g1677) & (!g3106)));
	assign g3913 = (((!g1610) & (!g1644) & (!g3515) & (g3031) & (g3084) & (g3912)) + ((!g1610) & (g1644) & (!g3515) & (!g3031) & (g3084) & (g3912)) + ((!g1610) & (g1644) & (!g3515) & (g3031) & (!g3084) & (g3912)) + ((!g1610) & (g1644) & (!g3515) & (g3031) & (g3084) & (g3912)) + ((!g1610) & (g1644) & (g3515) & (!g3031) & (g3084) & (g3912)) + ((!g1610) & (g1644) & (g3515) & (g3031) & (g3084) & (g3912)) + ((g1610) & (!g1644) & (!g3515) & (!g3031) & (g3084) & (g3912)) + ((g1610) & (!g1644) & (!g3515) & (g3031) & (g3084) & (g3912)) + ((g1610) & (!g1644) & (g3515) & (g3031) & (g3084) & (g3912)) + ((g1610) & (g1644) & (!g3515) & (!g3031) & (!g3084) & (g3912)) + ((g1610) & (g1644) & (!g3515) & (!g3031) & (g3084) & (g3912)) + ((g1610) & (g1644) & (!g3515) & (g3031) & (!g3084) & (g3912)) + ((g1610) & (g1644) & (!g3515) & (g3031) & (g3084) & (g3912)) + ((g1610) & (g1644) & (g3515) & (!g3031) & (g3084) & (g3912)) + ((g1610) & (g1644) & (g3515) & (g3031) & (!g3084) & (g3912)) + ((g1610) & (g1644) & (g3515) & (g3031) & (g3084) & (g3912)));
	assign g3914 = (((g1677) & (g3106)));
	assign g3915 = (((!g1711) & (!g3159) & (!g3913) & (g3914)) + ((!g1711) & (!g3159) & (g3913) & (!g3914)) + ((!g1711) & (!g3159) & (g3913) & (g3914)) + ((!g1711) & (g3159) & (!g3913) & (!g3914)) + ((g1711) & (!g3159) & (!g3913) & (!g3914)) + ((g1711) & (g3159) & (!g3913) & (g3914)) + ((g1711) & (g3159) & (g3913) & (!g3914)) + ((g1711) & (g3159) & (g3913) & (g3914)));
	assign g3916 = (((!g3136) & (g3113)) + ((g3136) & (!g3113)));
	assign g3917 = (((!g3038) & (!g3061) & (g3082) & (!g3532) & (g3078) & (g3916)) + ((!g3038) & (!g3061) & (g3082) & (g3532) & (g3078) & (g3916)) + ((!g3038) & (g3061) & (!g3082) & (!g3532) & (g3078) & (g3916)) + ((!g3038) & (g3061) & (g3082) & (!g3532) & (!g3078) & (g3916)) + ((!g3038) & (g3061) & (g3082) & (!g3532) & (g3078) & (g3916)) + ((!g3038) & (g3061) & (g3082) & (g3532) & (g3078) & (g3916)) + ((g3038) & (!g3061) & (!g3082) & (!g3532) & (g3078) & (g3916)) + ((g3038) & (!g3061) & (g3082) & (!g3532) & (!g3078) & (g3916)) + ((g3038) & (!g3061) & (g3082) & (!g3532) & (g3078) & (g3916)) + ((g3038) & (!g3061) & (g3082) & (g3532) & (g3078) & (g3916)) + ((g3038) & (g3061) & (!g3082) & (!g3532) & (g3078) & (g3916)) + ((g3038) & (g3061) & (!g3082) & (g3532) & (g3078) & (g3916)) + ((g3038) & (g3061) & (g3082) & (!g3532) & (!g3078) & (g3916)) + ((g3038) & (g3061) & (g3082) & (!g3532) & (g3078) & (g3916)) + ((g3038) & (g3061) & (g3082) & (g3532) & (!g3078) & (g3916)) + ((g3038) & (g3061) & (g3082) & (g3532) & (g3078) & (g3916)));
	assign g3918 = (((g3136) & (g3113)));
	assign g3919 = (((!g3153) & (!g3157) & (!g3917) & (g3918)) + ((!g3153) & (!g3157) & (g3917) & (!g3918)) + ((!g3153) & (!g3157) & (g3917) & (g3918)) + ((!g3153) & (g3157) & (!g3917) & (!g3918)) + ((g3153) & (!g3157) & (!g3917) & (!g3918)) + ((g3153) & (g3157) & (!g3917) & (g3918)) + ((g3153) & (g3157) & (g3917) & (!g3918)) + ((g3153) & (g3157) & (g3917) & (g3918)));
	assign g3920 = (((!g830) & (!g1914) & (!g1944) & (!g3915) & (!g3919) & (key[35])) + ((!g830) & (!g1914) & (!g1944) & (!g3915) & (g3919) & (key[35])) + ((!g830) & (!g1914) & (!g1944) & (g3915) & (!g3919) & (key[35])) + ((!g830) & (!g1914) & (!g1944) & (g3915) & (g3919) & (key[35])) + ((!g830) & (!g1914) & (g1944) & (!g3915) & (!g3919) & (key[35])) + ((!g830) & (!g1914) & (g1944) & (!g3915) & (g3919) & (key[35])) + ((!g830) & (!g1914) & (g1944) & (g3915) & (!g3919) & (key[35])) + ((!g830) & (!g1914) & (g1944) & (g3915) & (g3919) & (key[35])) + ((!g830) & (g1914) & (!g1944) & (!g3915) & (!g3919) & (key[35])) + ((!g830) & (g1914) & (!g1944) & (!g3915) & (g3919) & (key[35])) + ((!g830) & (g1914) & (!g1944) & (g3915) & (!g3919) & (key[35])) + ((!g830) & (g1914) & (!g1944) & (g3915) & (g3919) & (key[35])) + ((!g830) & (g1914) & (g1944) & (!g3915) & (!g3919) & (key[35])) + ((!g830) & (g1914) & (g1944) & (!g3915) & (g3919) & (key[35])) + ((!g830) & (g1914) & (g1944) & (g3915) & (!g3919) & (key[35])) + ((!g830) & (g1914) & (g1944) & (g3915) & (g3919) & (key[35])) + ((g830) & (!g1914) & (!g1944) & (!g3915) & (g3919) & (!key[35])) + ((g830) & (!g1914) & (!g1944) & (!g3915) & (g3919) & (key[35])) + ((g830) & (!g1914) & (!g1944) & (g3915) & (g3919) & (!key[35])) + ((g830) & (!g1914) & (!g1944) & (g3915) & (g3919) & (key[35])) + ((g830) & (!g1914) & (g1944) & (!g3915) & (!g3919) & (!key[35])) + ((g830) & (!g1914) & (g1944) & (!g3915) & (!g3919) & (key[35])) + ((g830) & (!g1914) & (g1944) & (g3915) & (!g3919) & (!key[35])) + ((g830) & (!g1914) & (g1944) & (g3915) & (!g3919) & (key[35])) + ((g830) & (g1914) & (!g1944) & (g3915) & (!g3919) & (!key[35])) + ((g830) & (g1914) & (!g1944) & (g3915) & (!g3919) & (key[35])) + ((g830) & (g1914) & (!g1944) & (g3915) & (g3919) & (!key[35])) + ((g830) & (g1914) & (!g1944) & (g3915) & (g3919) & (key[35])) + ((g830) & (g1914) & (g1944) & (!g3915) & (!g3919) & (!key[35])) + ((g830) & (g1914) & (g1944) & (!g3915) & (!g3919) & (key[35])) + ((g830) & (g1914) & (g1944) & (!g3915) & (g3919) & (!key[35])) + ((g830) & (g1914) & (g1944) & (!g3915) & (g3919) & (key[35])));
	assign g3921 = (((!g2295) & (!g2343) & (!g2916) & (g3009) & (!g3906) & (!g3907)) + ((!g2295) & (!g2343) & (!g2916) & (g3009) & (!g3906) & (g3907)) + ((!g2295) & (!g2343) & (!g2916) & (g3009) & (g3906) & (!g3907)) + ((!g2295) & (!g2343) & (!g2916) & (g3009) & (g3906) & (g3907)) + ((!g2295) & (!g2343) & (g2916) & (!g3009) & (!g3906) & (g3907)) + ((!g2295) & (!g2343) & (g2916) & (!g3009) & (g3906) & (!g3907)) + ((!g2295) & (!g2343) & (g2916) & (!g3009) & (g3906) & (g3907)) + ((!g2295) & (!g2343) & (g2916) & (g3009) & (!g3906) & (!g3907)) + ((!g2295) & (g2343) & (!g2916) & (!g3009) & (!g3906) & (!g3907)) + ((!g2295) & (g2343) & (!g2916) & (!g3009) & (!g3906) & (g3907)) + ((!g2295) & (g2343) & (!g2916) & (!g3009) & (g3906) & (!g3907)) + ((!g2295) & (g2343) & (!g2916) & (!g3009) & (g3906) & (g3907)) + ((!g2295) & (g2343) & (g2916) & (!g3009) & (!g3906) & (!g3907)) + ((!g2295) & (g2343) & (g2916) & (g3009) & (!g3906) & (g3907)) + ((!g2295) & (g2343) & (g2916) & (g3009) & (g3906) & (!g3907)) + ((!g2295) & (g2343) & (g2916) & (g3009) & (g3906) & (g3907)) + ((g2295) & (!g2343) & (!g2916) & (!g3009) & (!g3906) & (g3907)) + ((g2295) & (!g2343) & (!g2916) & (!g3009) & (g3906) & (!g3907)) + ((g2295) & (!g2343) & (!g2916) & (!g3009) & (g3906) & (g3907)) + ((g2295) & (!g2343) & (!g2916) & (g3009) & (!g3906) & (!g3907)) + ((g2295) & (!g2343) & (g2916) & (!g3009) & (!g3906) & (!g3907)) + ((g2295) & (!g2343) & (g2916) & (!g3009) & (!g3906) & (g3907)) + ((g2295) & (!g2343) & (g2916) & (!g3009) & (g3906) & (!g3907)) + ((g2295) & (!g2343) & (g2916) & (!g3009) & (g3906) & (g3907)) + ((g2295) & (g2343) & (!g2916) & (!g3009) & (!g3906) & (!g3907)) + ((g2295) & (g2343) & (!g2916) & (g3009) & (!g3906) & (g3907)) + ((g2295) & (g2343) & (!g2916) & (g3009) & (g3906) & (!g3907)) + ((g2295) & (g2343) & (!g2916) & (g3009) & (g3906) & (g3907)) + ((g2295) & (g2343) & (g2916) & (g3009) & (!g3906) & (!g3907)) + ((g2295) & (g2343) & (g2916) & (g3009) & (!g3906) & (g3907)) + ((g2295) & (g2343) & (g2916) & (g3009) & (g3906) & (!g3907)) + ((g2295) & (g2343) & (g2916) & (g3009) & (g3906) & (g3907)));
	assign g3922 = (((!g3898) & (!g3899) & (!g3168) & (!g3172) & (!g3213) & (!g3190)) + ((!g3898) & (!g3899) & (!g3168) & (!g3172) & (!g3213) & (g3190)) + ((!g3898) & (!g3899) & (!g3168) & (!g3172) & (g3213) & (!g3190)) + ((!g3898) & (!g3899) & (!g3168) & (g3172) & (!g3213) & (!g3190)) + ((!g3898) & (!g3899) & (!g3168) & (g3172) & (!g3213) & (g3190)) + ((!g3898) & (!g3899) & (!g3168) & (g3172) & (g3213) & (!g3190)) + ((!g3898) & (!g3899) & (g3168) & (!g3172) & (!g3213) & (!g3190)) + ((!g3898) & (!g3899) & (g3168) & (!g3172) & (!g3213) & (g3190)) + ((!g3898) & (!g3899) & (g3168) & (!g3172) & (g3213) & (!g3190)) + ((!g3898) & (!g3899) & (g3168) & (g3172) & (!g3213) & (!g3190)) + ((!g3898) & (g3899) & (!g3168) & (!g3172) & (!g3213) & (!g3190)) + ((!g3898) & (g3899) & (!g3168) & (!g3172) & (!g3213) & (g3190)) + ((!g3898) & (g3899) & (!g3168) & (!g3172) & (g3213) & (!g3190)) + ((!g3898) & (g3899) & (!g3168) & (g3172) & (!g3213) & (!g3190)) + ((!g3898) & (g3899) & (g3168) & (!g3172) & (!g3213) & (!g3190)) + ((!g3898) & (g3899) & (g3168) & (g3172) & (!g3213) & (!g3190)) + ((g3898) & (!g3899) & (!g3168) & (!g3172) & (!g3213) & (!g3190)) + ((g3898) & (!g3899) & (!g3168) & (!g3172) & (!g3213) & (g3190)) + ((g3898) & (!g3899) & (!g3168) & (!g3172) & (g3213) & (!g3190)) + ((g3898) & (!g3899) & (!g3168) & (g3172) & (!g3213) & (!g3190)) + ((g3898) & (!g3899) & (g3168) & (!g3172) & (!g3213) & (!g3190)) + ((g3898) & (!g3899) & (g3168) & (g3172) & (!g3213) & (!g3190)) + ((g3898) & (g3899) & (!g3168) & (!g3172) & (!g3213) & (!g3190)) + ((g3898) & (g3899) & (!g3168) & (!g3172) & (!g3213) & (g3190)) + ((g3898) & (g3899) & (!g3168) & (!g3172) & (g3213) & (!g3190)) + ((g3898) & (g3899) & (!g3168) & (g3172) & (!g3213) & (!g3190)) + ((g3898) & (g3899) & (g3168) & (!g3172) & (!g3213) & (!g3190)) + ((g3898) & (g3899) & (g3168) & (g3172) & (!g3213) & (!g3190)));
	assign g3923 = (((!g1914) & (!g3921) & (!g3922) & (!g3274) & (!g3284)) + ((!g1914) & (!g3921) & (!g3922) & (g3274) & (g3284)) + ((!g1914) & (!g3921) & (g3922) & (!g3274) & (g3284)) + ((!g1914) & (!g3921) & (g3922) & (g3274) & (!g3284)) + ((!g1914) & (g3921) & (!g3922) & (!g3274) & (!g3284)) + ((!g1914) & (g3921) & (!g3922) & (g3274) & (g3284)) + ((!g1914) & (g3921) & (g3922) & (!g3274) & (g3284)) + ((!g1914) & (g3921) & (g3922) & (g3274) & (!g3284)) + ((g1914) & (g3921) & (!g3922) & (!g3274) & (!g3284)) + ((g1914) & (g3921) & (!g3922) & (!g3274) & (g3284)) + ((g1914) & (g3921) & (!g3922) & (g3274) & (!g3284)) + ((g1914) & (g3921) & (!g3922) & (g3274) & (g3284)) + ((g1914) & (g3921) & (g3922) & (!g3274) & (!g3284)) + ((g1914) & (g3921) & (g3922) & (!g3274) & (g3284)) + ((g1914) & (g3921) & (g3922) & (g3274) & (!g3284)) + ((g1914) & (g3921) & (g3922) & (g3274) & (g3284)));
	assign g3924 = (((!g830) & (!g1945) & (!g3923) & (key[67])) + ((!g830) & (!g1945) & (g3923) & (key[67])) + ((!g830) & (g1945) & (!g3923) & (key[67])) + ((!g830) & (g1945) & (g3923) & (key[67])) + ((g830) & (!g1945) & (g3923) & (!key[67])) + ((g830) & (!g1945) & (g3923) & (key[67])) + ((g830) & (g1945) & (!g3923) & (!key[67])) + ((g830) & (g1945) & (!g3923) & (key[67])));
	assign g3925 = (((!g1711) & (!g3159) & (!g3913) & (!g3914)) + ((!g1711) & (!g3159) & (!g3913) & (g3914)) + ((!g1711) & (!g3159) & (g3913) & (!g3914)) + ((!g1711) & (!g3159) & (g3913) & (g3914)) + ((!g1711) & (g3159) & (!g3913) & (!g3914)) + ((g1711) & (!g3159) & (!g3913) & (!g3914)));
	assign g3926 = (((g1914) & (!g1744) & (!g3177) & (!g3925)) + ((g1914) & (!g1744) & (g3177) & (g3925)) + ((g1914) & (g1744) & (!g3177) & (g3925)) + ((g1914) & (g1744) & (g3177) & (!g3925)));
	assign g3927 = (((!g3153) & (!g3157) & (!g3917) & (!g3918)) + ((!g3153) & (!g3157) & (!g3917) & (g3918)) + ((!g3153) & (!g3157) & (g3917) & (!g3918)) + ((!g3153) & (!g3157) & (g3917) & (g3918)) + ((!g3153) & (g3157) & (!g3917) & (!g3918)) + ((g3153) & (!g3157) & (!g3917) & (!g3918)));
	assign g3928 = (((!g1914) & (!g3207) & (!g3184) & (!g3927)) + ((!g1914) & (!g3207) & (g3184) & (g3927)) + ((!g1914) & (g3207) & (!g3184) & (g3927)) + ((!g1914) & (g3207) & (g3184) & (!g3927)));
	assign g3929 = (((!g830) & (!g1946) & (!g3926) & (!g3928) & (key[36])) + ((!g830) & (!g1946) & (!g3926) & (g3928) & (key[36])) + ((!g830) & (!g1946) & (g3926) & (!g3928) & (key[36])) + ((!g830) & (!g1946) & (g3926) & (g3928) & (key[36])) + ((!g830) & (g1946) & (!g3926) & (!g3928) & (key[36])) + ((!g830) & (g1946) & (!g3926) & (g3928) & (key[36])) + ((!g830) & (g1946) & (g3926) & (!g3928) & (key[36])) + ((!g830) & (g1946) & (g3926) & (g3928) & (key[36])) + ((g830) & (!g1946) & (!g3926) & (g3928) & (!key[36])) + ((g830) & (!g1946) & (!g3926) & (g3928) & (key[36])) + ((g830) & (!g1946) & (g3926) & (!g3928) & (!key[36])) + ((g830) & (!g1946) & (g3926) & (!g3928) & (key[36])) + ((g830) & (!g1946) & (g3926) & (g3928) & (!key[36])) + ((g830) & (!g1946) & (g3926) & (g3928) & (key[36])) + ((g830) & (g1946) & (!g3926) & (!g3928) & (!key[36])) + ((g830) & (g1946) & (!g3926) & (!g3928) & (key[36])));
	assign g3930 = (((!g2295) & (!g2343) & (!g2916) & (!g3009) & (!g3906) & (!g3907)) + ((!g2295) & (!g2343) & (!g2916) & (!g3009) & (!g3906) & (g3907)) + ((!g2295) & (!g2343) & (!g2916) & (!g3009) & (g3906) & (!g3907)) + ((!g2295) & (!g2343) & (!g2916) & (!g3009) & (g3906) & (g3907)) + ((!g2295) & (!g2343) & (!g2916) & (g3009) & (!g3906) & (!g3907)) + ((!g2295) & (!g2343) & (!g2916) & (g3009) & (!g3906) & (g3907)) + ((!g2295) & (!g2343) & (!g2916) & (g3009) & (g3906) & (!g3907)) + ((!g2295) & (!g2343) & (!g2916) & (g3009) & (g3906) & (g3907)) + ((!g2295) & (!g2343) & (g2916) & (!g3009) & (!g3906) & (!g3907)) + ((!g2295) & (!g2343) & (g2916) & (!g3009) & (!g3906) & (g3907)) + ((!g2295) & (!g2343) & (g2916) & (!g3009) & (g3906) & (!g3907)) + ((!g2295) & (!g2343) & (g2916) & (!g3009) & (g3906) & (g3907)) + ((!g2295) & (!g2343) & (g2916) & (g3009) & (!g3906) & (!g3907)) + ((!g2295) & (g2343) & (!g2916) & (!g3009) & (!g3906) & (!g3907)) + ((!g2295) & (g2343) & (!g2916) & (!g3009) & (!g3906) & (g3907)) + ((!g2295) & (g2343) & (!g2916) & (!g3009) & (g3906) & (!g3907)) + ((!g2295) & (g2343) & (!g2916) & (!g3009) & (g3906) & (g3907)) + ((!g2295) & (g2343) & (g2916) & (!g3009) & (!g3906) & (!g3907)) + ((g2295) & (!g2343) & (!g2916) & (!g3009) & (!g3906) & (!g3907)) + ((g2295) & (!g2343) & (!g2916) & (!g3009) & (!g3906) & (g3907)) + ((g2295) & (!g2343) & (!g2916) & (!g3009) & (g3906) & (!g3907)) + ((g2295) & (!g2343) & (!g2916) & (!g3009) & (g3906) & (g3907)) + ((g2295) & (!g2343) & (!g2916) & (g3009) & (!g3906) & (!g3907)) + ((g2295) & (!g2343) & (g2916) & (!g3009) & (!g3906) & (!g3907)) + ((g2295) & (!g2343) & (g2916) & (!g3009) & (!g3906) & (g3907)) + ((g2295) & (!g2343) & (g2916) & (!g3009) & (g3906) & (!g3907)) + ((g2295) & (!g2343) & (g2916) & (!g3009) & (g3906) & (g3907)) + ((g2295) & (g2343) & (!g2916) & (!g3009) & (!g3906) & (!g3907)));
	assign g3931 = (((!g2376) & (!g3031) & (!g3930)) + ((!g2376) & (g3031) & (g3930)) + ((g2376) & (!g3031) & (g3930)) + ((g2376) & (g3031) & (!g3930)));
	assign g3932 = (((!g3922) & (!g3274) & (!g3284) & (!g3314) & (g3299)) + ((!g3922) & (!g3274) & (!g3284) & (g3314) & (!g3299)) + ((!g3922) & (!g3274) & (g3284) & (!g3314) & (!g3299)) + ((!g3922) & (!g3274) & (g3284) & (g3314) & (g3299)) + ((!g3922) & (g3274) & (!g3284) & (!g3314) & (!g3299)) + ((!g3922) & (g3274) & (!g3284) & (g3314) & (g3299)) + ((!g3922) & (g3274) & (g3284) & (!g3314) & (!g3299)) + ((!g3922) & (g3274) & (g3284) & (g3314) & (g3299)) + ((g3922) & (!g3274) & (!g3284) & (!g3314) & (g3299)) + ((g3922) & (!g3274) & (!g3284) & (g3314) & (!g3299)) + ((g3922) & (!g3274) & (g3284) & (!g3314) & (g3299)) + ((g3922) & (!g3274) & (g3284) & (g3314) & (!g3299)) + ((g3922) & (g3274) & (!g3284) & (!g3314) & (g3299)) + ((g3922) & (g3274) & (!g3284) & (g3314) & (!g3299)) + ((g3922) & (g3274) & (g3284) & (!g3314) & (!g3299)) + ((g3922) & (g3274) & (g3284) & (g3314) & (g3299)));
	assign g3933 = (((!g830) & (!g1914) & (!g1947) & (!g3931) & (!g3932) & (key[68])) + ((!g830) & (!g1914) & (!g1947) & (!g3931) & (g3932) & (key[68])) + ((!g830) & (!g1914) & (!g1947) & (g3931) & (!g3932) & (key[68])) + ((!g830) & (!g1914) & (!g1947) & (g3931) & (g3932) & (key[68])) + ((!g830) & (!g1914) & (g1947) & (!g3931) & (!g3932) & (key[68])) + ((!g830) & (!g1914) & (g1947) & (!g3931) & (g3932) & (key[68])) + ((!g830) & (!g1914) & (g1947) & (g3931) & (!g3932) & (key[68])) + ((!g830) & (!g1914) & (g1947) & (g3931) & (g3932) & (key[68])) + ((!g830) & (g1914) & (!g1947) & (!g3931) & (!g3932) & (key[68])) + ((!g830) & (g1914) & (!g1947) & (!g3931) & (g3932) & (key[68])) + ((!g830) & (g1914) & (!g1947) & (g3931) & (!g3932) & (key[68])) + ((!g830) & (g1914) & (!g1947) & (g3931) & (g3932) & (key[68])) + ((!g830) & (g1914) & (g1947) & (!g3931) & (!g3932) & (key[68])) + ((!g830) & (g1914) & (g1947) & (!g3931) & (g3932) & (key[68])) + ((!g830) & (g1914) & (g1947) & (g3931) & (!g3932) & (key[68])) + ((!g830) & (g1914) & (g1947) & (g3931) & (g3932) & (key[68])) + ((g830) & (!g1914) & (!g1947) & (!g3931) & (g3932) & (!key[68])) + ((g830) & (!g1914) & (!g1947) & (!g3931) & (g3932) & (key[68])) + ((g830) & (!g1914) & (!g1947) & (g3931) & (g3932) & (!key[68])) + ((g830) & (!g1914) & (!g1947) & (g3931) & (g3932) & (key[68])) + ((g830) & (!g1914) & (g1947) & (!g3931) & (!g3932) & (!key[68])) + ((g830) & (!g1914) & (g1947) & (!g3931) & (!g3932) & (key[68])) + ((g830) & (!g1914) & (g1947) & (g3931) & (!g3932) & (!key[68])) + ((g830) & (!g1914) & (g1947) & (g3931) & (!g3932) & (key[68])) + ((g830) & (g1914) & (!g1947) & (g3931) & (!g3932) & (!key[68])) + ((g830) & (g1914) & (!g1947) & (g3931) & (!g3932) & (key[68])) + ((g830) & (g1914) & (!g1947) & (g3931) & (g3932) & (!key[68])) + ((g830) & (g1914) & (!g1947) & (g3931) & (g3932) & (key[68])) + ((g830) & (g1914) & (g1947) & (!g3931) & (!g3932) & (!key[68])) + ((g830) & (g1914) & (g1947) & (!g3931) & (!g3932) & (key[68])) + ((g830) & (g1914) & (g1947) & (!g3931) & (g3932) & (!key[68])) + ((g830) & (g1914) & (g1947) & (!g3931) & (g3932) & (key[68])));
	assign g3934 = (((!g1711) & (!g1744) & (!g3159) & (!g3177) & (!g3913) & (!g3914)) + ((!g1711) & (!g1744) & (!g3159) & (!g3177) & (!g3913) & (g3914)) + ((!g1711) & (!g1744) & (!g3159) & (!g3177) & (g3913) & (!g3914)) + ((!g1711) & (!g1744) & (!g3159) & (!g3177) & (g3913) & (g3914)) + ((!g1711) & (!g1744) & (!g3159) & (g3177) & (!g3913) & (!g3914)) + ((!g1711) & (!g1744) & (!g3159) & (g3177) & (!g3913) & (g3914)) + ((!g1711) & (!g1744) & (!g3159) & (g3177) & (g3913) & (!g3914)) + ((!g1711) & (!g1744) & (!g3159) & (g3177) & (g3913) & (g3914)) + ((!g1711) & (!g1744) & (g3159) & (!g3177) & (!g3913) & (!g3914)) + ((!g1711) & (!g1744) & (g3159) & (!g3177) & (!g3913) & (g3914)) + ((!g1711) & (!g1744) & (g3159) & (!g3177) & (g3913) & (!g3914)) + ((!g1711) & (!g1744) & (g3159) & (!g3177) & (g3913) & (g3914)) + ((!g1711) & (!g1744) & (g3159) & (g3177) & (!g3913) & (!g3914)) + ((!g1711) & (g1744) & (!g3159) & (!g3177) & (!g3913) & (!g3914)) + ((!g1711) & (g1744) & (!g3159) & (!g3177) & (!g3913) & (g3914)) + ((!g1711) & (g1744) & (!g3159) & (!g3177) & (g3913) & (!g3914)) + ((!g1711) & (g1744) & (!g3159) & (!g3177) & (g3913) & (g3914)) + ((!g1711) & (g1744) & (g3159) & (!g3177) & (!g3913) & (!g3914)) + ((g1711) & (!g1744) & (!g3159) & (!g3177) & (!g3913) & (!g3914)) + ((g1711) & (!g1744) & (!g3159) & (!g3177) & (!g3913) & (g3914)) + ((g1711) & (!g1744) & (!g3159) & (!g3177) & (g3913) & (!g3914)) + ((g1711) & (!g1744) & (!g3159) & (!g3177) & (g3913) & (g3914)) + ((g1711) & (!g1744) & (!g3159) & (g3177) & (!g3913) & (!g3914)) + ((g1711) & (!g1744) & (g3159) & (!g3177) & (!g3913) & (!g3914)) + ((g1711) & (!g1744) & (g3159) & (!g3177) & (!g3913) & (g3914)) + ((g1711) & (!g1744) & (g3159) & (!g3177) & (g3913) & (!g3914)) + ((g1711) & (!g1744) & (g3159) & (!g3177) & (g3913) & (g3914)) + ((g1711) & (g1744) & (!g3159) & (!g3177) & (!g3913) & (!g3914)));
	assign g3935 = (((g1914) & (!g1778) & (!g3250) & (!g3934)) + ((g1914) & (!g1778) & (g3250) & (g3934)) + ((g1914) & (g1778) & (!g3250) & (g3934)) + ((g1914) & (g1778) & (g3250) & (!g3934)));
	assign g3936 = (((!g3153) & (!g3157) & (!g3207) & (!g3184) & (!g3917) & (!g3918)) + ((!g3153) & (!g3157) & (!g3207) & (!g3184) & (!g3917) & (g3918)) + ((!g3153) & (!g3157) & (!g3207) & (!g3184) & (g3917) & (!g3918)) + ((!g3153) & (!g3157) & (!g3207) & (!g3184) & (g3917) & (g3918)) + ((!g3153) & (!g3157) & (!g3207) & (g3184) & (!g3917) & (!g3918)) + ((!g3153) & (!g3157) & (!g3207) & (g3184) & (!g3917) & (g3918)) + ((!g3153) & (!g3157) & (!g3207) & (g3184) & (g3917) & (!g3918)) + ((!g3153) & (!g3157) & (!g3207) & (g3184) & (g3917) & (g3918)) + ((!g3153) & (!g3157) & (g3207) & (!g3184) & (!g3917) & (!g3918)) + ((!g3153) & (!g3157) & (g3207) & (!g3184) & (!g3917) & (g3918)) + ((!g3153) & (!g3157) & (g3207) & (!g3184) & (g3917) & (!g3918)) + ((!g3153) & (!g3157) & (g3207) & (!g3184) & (g3917) & (g3918)) + ((!g3153) & (g3157) & (!g3207) & (!g3184) & (!g3917) & (!g3918)) + ((!g3153) & (g3157) & (!g3207) & (!g3184) & (!g3917) & (g3918)) + ((!g3153) & (g3157) & (!g3207) & (!g3184) & (g3917) & (!g3918)) + ((!g3153) & (g3157) & (!g3207) & (!g3184) & (g3917) & (g3918)) + ((!g3153) & (g3157) & (!g3207) & (g3184) & (!g3917) & (!g3918)) + ((!g3153) & (g3157) & (g3207) & (!g3184) & (!g3917) & (!g3918)) + ((g3153) & (!g3157) & (!g3207) & (!g3184) & (!g3917) & (!g3918)) + ((g3153) & (!g3157) & (!g3207) & (!g3184) & (!g3917) & (g3918)) + ((g3153) & (!g3157) & (!g3207) & (!g3184) & (g3917) & (!g3918)) + ((g3153) & (!g3157) & (!g3207) & (!g3184) & (g3917) & (g3918)) + ((g3153) & (!g3157) & (!g3207) & (g3184) & (!g3917) & (!g3918)) + ((g3153) & (!g3157) & (g3207) & (!g3184) & (!g3917) & (!g3918)) + ((g3153) & (g3157) & (!g3207) & (!g3184) & (!g3917) & (!g3918)) + ((g3153) & (g3157) & (!g3207) & (!g3184) & (!g3917) & (g3918)) + ((g3153) & (g3157) & (!g3207) & (!g3184) & (g3917) & (!g3918)) + ((g3153) & (g3157) & (!g3207) & (!g3184) & (g3917) & (g3918)));
	assign g3937 = (((!g1914) & (!g3235) & (!g3245) & (!g3936)) + ((!g1914) & (!g3235) & (g3245) & (g3936)) + ((!g1914) & (g3235) & (!g3245) & (g3936)) + ((!g1914) & (g3235) & (g3245) & (!g3936)));
	assign g3938 = (((!g830) & (!g1948) & (!g3935) & (!g3937) & (key[37])) + ((!g830) & (!g1948) & (!g3935) & (g3937) & (key[37])) + ((!g830) & (!g1948) & (g3935) & (!g3937) & (key[37])) + ((!g830) & (!g1948) & (g3935) & (g3937) & (key[37])) + ((!g830) & (g1948) & (!g3935) & (!g3937) & (key[37])) + ((!g830) & (g1948) & (!g3935) & (g3937) & (key[37])) + ((!g830) & (g1948) & (g3935) & (!g3937) & (key[37])) + ((!g830) & (g1948) & (g3935) & (g3937) & (key[37])) + ((g830) & (!g1948) & (!g3935) & (g3937) & (!key[37])) + ((g830) & (!g1948) & (!g3935) & (g3937) & (key[37])) + ((g830) & (!g1948) & (g3935) & (!g3937) & (!key[37])) + ((g830) & (!g1948) & (g3935) & (!g3937) & (key[37])) + ((g830) & (!g1948) & (g3935) & (g3937) & (!key[37])) + ((g830) & (!g1948) & (g3935) & (g3937) & (key[37])) + ((g830) & (g1948) & (!g3935) & (!g3937) & (!key[37])) + ((g830) & (g1948) & (!g3935) & (!g3937) & (key[37])));
	assign g3939 = (((!g2376) & (g3031) & (!g3930)) + ((g2376) & (!g3031) & (!g3930)) + ((g2376) & (g3031) & (!g3930)) + ((g2376) & (g3031) & (g3930)));
	assign g3940 = (((!g3922) & (!g3274) & (!g3284) & (g3314) & (g3299)) + ((!g3922) & (!g3274) & (g3284) & (!g3314) & (g3299)) + ((!g3922) & (!g3274) & (g3284) & (g3314) & (!g3299)) + ((!g3922) & (!g3274) & (g3284) & (g3314) & (g3299)) + ((!g3922) & (g3274) & (!g3284) & (!g3314) & (g3299)) + ((!g3922) & (g3274) & (!g3284) & (g3314) & (!g3299)) + ((!g3922) & (g3274) & (!g3284) & (g3314) & (g3299)) + ((!g3922) & (g3274) & (g3284) & (!g3314) & (g3299)) + ((!g3922) & (g3274) & (g3284) & (g3314) & (!g3299)) + ((!g3922) & (g3274) & (g3284) & (g3314) & (g3299)) + ((g3922) & (!g3274) & (!g3284) & (g3314) & (g3299)) + ((g3922) & (!g3274) & (g3284) & (g3314) & (g3299)) + ((g3922) & (g3274) & (!g3284) & (g3314) & (g3299)) + ((g3922) & (g3274) & (g3284) & (!g3314) & (g3299)) + ((g3922) & (g3274) & (g3284) & (g3314) & (!g3299)) + ((g3922) & (g3274) & (g3284) & (g3314) & (g3299)));
	assign g3941 = (((!g830) & (key[69]) & (!g1914) & (!g3940) & (!g3939) & (!g5665)) + ((!g830) & (key[69]) & (!g1914) & (!g3940) & (!g3939) & (g5665)) + ((!g830) & (key[69]) & (!g1914) & (!g3940) & (g3939) & (!g5665)) + ((!g830) & (key[69]) & (!g1914) & (!g3940) & (g3939) & (g5665)) + ((!g830) & (key[69]) & (!g1914) & (g3940) & (!g3939) & (!g5665)) + ((!g830) & (key[69]) & (!g1914) & (g3940) & (!g3939) & (g5665)) + ((!g830) & (key[69]) & (!g1914) & (g3940) & (g3939) & (!g5665)) + ((!g830) & (key[69]) & (!g1914) & (g3940) & (g3939) & (g5665)) + ((!g830) & (key[69]) & (g1914) & (!g3940) & (!g3939) & (!g5665)) + ((!g830) & (key[69]) & (g1914) & (!g3940) & (!g3939) & (g5665)) + ((!g830) & (key[69]) & (g1914) & (!g3940) & (g3939) & (!g5665)) + ((!g830) & (key[69]) & (g1914) & (!g3940) & (g3939) & (g5665)) + ((!g830) & (key[69]) & (g1914) & (g3940) & (!g3939) & (!g5665)) + ((!g830) & (key[69]) & (g1914) & (g3940) & (!g3939) & (g5665)) + ((!g830) & (key[69]) & (g1914) & (g3940) & (g3939) & (!g5665)) + ((!g830) & (key[69]) & (g1914) & (g3940) & (g3939) & (g5665)) + ((g830) & (!key[69]) & (!g1914) & (!g3940) & (!g3939) & (!g5665)) + ((g830) & (!key[69]) & (!g1914) & (!g3940) & (g3939) & (!g5665)) + ((g830) & (!key[69]) & (!g1914) & (g3940) & (!g3939) & (g5665)) + ((g830) & (!key[69]) & (!g1914) & (g3940) & (g3939) & (g5665)) + ((g830) & (!key[69]) & (g1914) & (!g3940) & (!g3939) & (!g5665)) + ((g830) & (!key[69]) & (g1914) & (!g3940) & (g3939) & (g5665)) + ((g830) & (!key[69]) & (g1914) & (g3940) & (!g3939) & (!g5665)) + ((g830) & (!key[69]) & (g1914) & (g3940) & (g3939) & (g5665)) + ((g830) & (key[69]) & (!g1914) & (!g3940) & (!g3939) & (!g5665)) + ((g830) & (key[69]) & (!g1914) & (!g3940) & (g3939) & (!g5665)) + ((g830) & (key[69]) & (!g1914) & (g3940) & (!g3939) & (g5665)) + ((g830) & (key[69]) & (!g1914) & (g3940) & (g3939) & (g5665)) + ((g830) & (key[69]) & (g1914) & (!g3940) & (!g3939) & (!g5665)) + ((g830) & (key[69]) & (g1914) & (!g3940) & (g3939) & (g5665)) + ((g830) & (key[69]) & (g1914) & (g3940) & (!g3939) & (!g5665)) + ((g830) & (key[69]) & (g1914) & (g3940) & (g3939) & (g5665)));
	assign g3942 = (((!g1778) & (!g1814) & (!g3250) & (g3291) & (!g3934)) + ((!g1778) & (!g1814) & (!g3250) & (g3291) & (g3934)) + ((!g1778) & (!g1814) & (g3250) & (!g3291) & (!g3934)) + ((!g1778) & (!g1814) & (g3250) & (g3291) & (g3934)) + ((!g1778) & (g1814) & (!g3250) & (!g3291) & (!g3934)) + ((!g1778) & (g1814) & (!g3250) & (!g3291) & (g3934)) + ((!g1778) & (g1814) & (g3250) & (!g3291) & (g3934)) + ((!g1778) & (g1814) & (g3250) & (g3291) & (!g3934)) + ((g1778) & (!g1814) & (!g3250) & (!g3291) & (!g3934)) + ((g1778) & (!g1814) & (!g3250) & (g3291) & (g3934)) + ((g1778) & (!g1814) & (g3250) & (!g3291) & (!g3934)) + ((g1778) & (!g1814) & (g3250) & (!g3291) & (g3934)) + ((g1778) & (g1814) & (!g3250) & (!g3291) & (g3934)) + ((g1778) & (g1814) & (!g3250) & (g3291) & (!g3934)) + ((g1778) & (g1814) & (g3250) & (g3291) & (!g3934)) + ((g1778) & (g1814) & (g3250) & (g3291) & (g3934)));
	assign g3943 = (((!g3235) & (!g3245) & (!g3310) & (g3295) & (!g3936)) + ((!g3235) & (!g3245) & (!g3310) & (g3295) & (g3936)) + ((!g3235) & (!g3245) & (g3310) & (!g3295) & (!g3936)) + ((!g3235) & (!g3245) & (g3310) & (!g3295) & (g3936)) + ((!g3235) & (g3245) & (!g3310) & (!g3295) & (!g3936)) + ((!g3235) & (g3245) & (!g3310) & (g3295) & (g3936)) + ((!g3235) & (g3245) & (g3310) & (!g3295) & (g3936)) + ((!g3235) & (g3245) & (g3310) & (g3295) & (!g3936)) + ((g3235) & (!g3245) & (!g3310) & (!g3295) & (!g3936)) + ((g3235) & (!g3245) & (!g3310) & (g3295) & (g3936)) + ((g3235) & (!g3245) & (g3310) & (!g3295) & (g3936)) + ((g3235) & (!g3245) & (g3310) & (g3295) & (!g3936)) + ((g3235) & (g3245) & (!g3310) & (!g3295) & (!g3936)) + ((g3235) & (g3245) & (!g3310) & (!g3295) & (g3936)) + ((g3235) & (g3245) & (g3310) & (g3295) & (!g3936)) + ((g3235) & (g3245) & (g3310) & (g3295) & (g3936)));
	assign g3944 = (((!g830) & (!g1914) & (!g1953) & (!g3942) & (!g3943) & (key[38])) + ((!g830) & (!g1914) & (!g1953) & (!g3942) & (g3943) & (key[38])) + ((!g830) & (!g1914) & (!g1953) & (g3942) & (!g3943) & (key[38])) + ((!g830) & (!g1914) & (!g1953) & (g3942) & (g3943) & (key[38])) + ((!g830) & (!g1914) & (g1953) & (!g3942) & (!g3943) & (key[38])) + ((!g830) & (!g1914) & (g1953) & (!g3942) & (g3943) & (key[38])) + ((!g830) & (!g1914) & (g1953) & (g3942) & (!g3943) & (key[38])) + ((!g830) & (!g1914) & (g1953) & (g3942) & (g3943) & (key[38])) + ((!g830) & (g1914) & (!g1953) & (!g3942) & (!g3943) & (key[38])) + ((!g830) & (g1914) & (!g1953) & (!g3942) & (g3943) & (key[38])) + ((!g830) & (g1914) & (!g1953) & (g3942) & (!g3943) & (key[38])) + ((!g830) & (g1914) & (!g1953) & (g3942) & (g3943) & (key[38])) + ((!g830) & (g1914) & (g1953) & (!g3942) & (!g3943) & (key[38])) + ((!g830) & (g1914) & (g1953) & (!g3942) & (g3943) & (key[38])) + ((!g830) & (g1914) & (g1953) & (g3942) & (!g3943) & (key[38])) + ((!g830) & (g1914) & (g1953) & (g3942) & (g3943) & (key[38])) + ((g830) & (!g1914) & (!g1953) & (!g3942) & (g3943) & (!key[38])) + ((g830) & (!g1914) & (!g1953) & (!g3942) & (g3943) & (key[38])) + ((g830) & (!g1914) & (!g1953) & (g3942) & (g3943) & (!key[38])) + ((g830) & (!g1914) & (!g1953) & (g3942) & (g3943) & (key[38])) + ((g830) & (!g1914) & (g1953) & (!g3942) & (!g3943) & (!key[38])) + ((g830) & (!g1914) & (g1953) & (!g3942) & (!g3943) & (key[38])) + ((g830) & (!g1914) & (g1953) & (g3942) & (!g3943) & (!key[38])) + ((g830) & (!g1914) & (g1953) & (g3942) & (!g3943) & (key[38])) + ((g830) & (g1914) & (!g1953) & (g3942) & (!g3943) & (!key[38])) + ((g830) & (g1914) & (!g1953) & (g3942) & (!g3943) & (key[38])) + ((g830) & (g1914) & (!g1953) & (g3942) & (g3943) & (!key[38])) + ((g830) & (g1914) & (!g1953) & (g3942) & (g3943) & (key[38])) + ((g830) & (g1914) & (g1953) & (!g3942) & (!g3943) & (!key[38])) + ((g830) & (g1914) & (g1953) & (!g3942) & (!g3943) & (key[38])) + ((g830) & (g1914) & (g1953) & (!g3942) & (g3943) & (!key[38])) + ((g830) & (g1914) & (g1953) & (!g3942) & (g3943) & (key[38])));
	assign g3945 = (((!g2423) & (!g2515) & (!g3084) & (g3106) & (!g3939)) + ((!g2423) & (!g2515) & (!g3084) & (g3106) & (g3939)) + ((!g2423) & (!g2515) & (g3084) & (!g3106) & (g3939)) + ((!g2423) & (!g2515) & (g3084) & (g3106) & (!g3939)) + ((!g2423) & (g2515) & (!g3084) & (!g3106) & (!g3939)) + ((!g2423) & (g2515) & (!g3084) & (!g3106) & (g3939)) + ((!g2423) & (g2515) & (g3084) & (!g3106) & (!g3939)) + ((!g2423) & (g2515) & (g3084) & (g3106) & (g3939)) + ((g2423) & (!g2515) & (!g3084) & (!g3106) & (g3939)) + ((g2423) & (!g2515) & (!g3084) & (g3106) & (!g3939)) + ((g2423) & (!g2515) & (g3084) & (!g3106) & (!g3939)) + ((g2423) & (!g2515) & (g3084) & (!g3106) & (g3939)) + ((g2423) & (g2515) & (!g3084) & (!g3106) & (!g3939)) + ((g2423) & (g2515) & (!g3084) & (g3106) & (g3939)) + ((g2423) & (g2515) & (g3084) & (g3106) & (!g3939)) + ((g2423) & (g2515) & (g3084) & (g3106) & (g3939)));
	assign g3946 = (((!g3940) & (!g3353) & (!g3359) & (!g3389) & (g3374)) + ((!g3940) & (!g3353) & (!g3359) & (g3389) & (!g3374)) + ((!g3940) & (!g3353) & (g3359) & (!g3389) & (g3374)) + ((!g3940) & (!g3353) & (g3359) & (g3389) & (!g3374)) + ((!g3940) & (g3353) & (!g3359) & (!g3389) & (g3374)) + ((!g3940) & (g3353) & (!g3359) & (g3389) & (!g3374)) + ((!g3940) & (g3353) & (g3359) & (!g3389) & (!g3374)) + ((!g3940) & (g3353) & (g3359) & (g3389) & (g3374)) + ((g3940) & (!g3353) & (!g3359) & (!g3389) & (g3374)) + ((g3940) & (!g3353) & (!g3359) & (g3389) & (!g3374)) + ((g3940) & (!g3353) & (g3359) & (!g3389) & (!g3374)) + ((g3940) & (!g3353) & (g3359) & (g3389) & (g3374)) + ((g3940) & (g3353) & (!g3359) & (!g3389) & (!g3374)) + ((g3940) & (g3353) & (!g3359) & (g3389) & (g3374)) + ((g3940) & (g3353) & (g3359) & (!g3389) & (!g3374)) + ((g3940) & (g3353) & (g3359) & (g3389) & (g3374)));
	assign g3947 = (((!g830) & (!g1914) & (!g1954) & (!g3945) & (!g3946) & (key[70])) + ((!g830) & (!g1914) & (!g1954) & (!g3945) & (g3946) & (key[70])) + ((!g830) & (!g1914) & (!g1954) & (g3945) & (!g3946) & (key[70])) + ((!g830) & (!g1914) & (!g1954) & (g3945) & (g3946) & (key[70])) + ((!g830) & (!g1914) & (g1954) & (!g3945) & (!g3946) & (key[70])) + ((!g830) & (!g1914) & (g1954) & (!g3945) & (g3946) & (key[70])) + ((!g830) & (!g1914) & (g1954) & (g3945) & (!g3946) & (key[70])) + ((!g830) & (!g1914) & (g1954) & (g3945) & (g3946) & (key[70])) + ((!g830) & (g1914) & (!g1954) & (!g3945) & (!g3946) & (key[70])) + ((!g830) & (g1914) & (!g1954) & (!g3945) & (g3946) & (key[70])) + ((!g830) & (g1914) & (!g1954) & (g3945) & (!g3946) & (key[70])) + ((!g830) & (g1914) & (!g1954) & (g3945) & (g3946) & (key[70])) + ((!g830) & (g1914) & (g1954) & (!g3945) & (!g3946) & (key[70])) + ((!g830) & (g1914) & (g1954) & (!g3945) & (g3946) & (key[70])) + ((!g830) & (g1914) & (g1954) & (g3945) & (!g3946) & (key[70])) + ((!g830) & (g1914) & (g1954) & (g3945) & (g3946) & (key[70])) + ((g830) & (!g1914) & (!g1954) & (!g3945) & (g3946) & (!key[70])) + ((g830) & (!g1914) & (!g1954) & (!g3945) & (g3946) & (key[70])) + ((g830) & (!g1914) & (!g1954) & (g3945) & (g3946) & (!key[70])) + ((g830) & (!g1914) & (!g1954) & (g3945) & (g3946) & (key[70])) + ((g830) & (!g1914) & (g1954) & (!g3945) & (!g3946) & (!key[70])) + ((g830) & (!g1914) & (g1954) & (!g3945) & (!g3946) & (key[70])) + ((g830) & (!g1914) & (g1954) & (g3945) & (!g3946) & (!key[70])) + ((g830) & (!g1914) & (g1954) & (g3945) & (!g3946) & (key[70])) + ((g830) & (g1914) & (!g1954) & (g3945) & (!g3946) & (!key[70])) + ((g830) & (g1914) & (!g1954) & (g3945) & (!g3946) & (key[70])) + ((g830) & (g1914) & (!g1954) & (g3945) & (g3946) & (!key[70])) + ((g830) & (g1914) & (!g1954) & (g3945) & (g3946) & (key[70])) + ((g830) & (g1914) & (g1954) & (!g3945) & (!g3946) & (!key[70])) + ((g830) & (g1914) & (g1954) & (!g3945) & (!g3946) & (key[70])) + ((g830) & (g1914) & (g1954) & (!g3945) & (g3946) & (!key[70])) + ((g830) & (g1914) & (g1954) & (!g3945) & (g3946) & (key[70])));
	assign g3948 = (((!g1778) & (!g1814) & (g3250) & (g3291) & (!g3934)) + ((!g1778) & (g1814) & (!g3250) & (g3291) & (!g3934)) + ((!g1778) & (g1814) & (!g3250) & (g3291) & (g3934)) + ((!g1778) & (g1814) & (g3250) & (!g3291) & (!g3934)) + ((!g1778) & (g1814) & (g3250) & (g3291) & (!g3934)) + ((!g1778) & (g1814) & (g3250) & (g3291) & (g3934)) + ((g1778) & (!g1814) & (!g3250) & (g3291) & (!g3934)) + ((g1778) & (!g1814) & (g3250) & (g3291) & (!g3934)) + ((g1778) & (!g1814) & (g3250) & (g3291) & (g3934)) + ((g1778) & (g1814) & (!g3250) & (!g3291) & (!g3934)) + ((g1778) & (g1814) & (!g3250) & (g3291) & (!g3934)) + ((g1778) & (g1814) & (!g3250) & (g3291) & (g3934)) + ((g1778) & (g1814) & (g3250) & (!g3291) & (!g3934)) + ((g1778) & (g1814) & (g3250) & (!g3291) & (g3934)) + ((g1778) & (g1814) & (g3250) & (g3291) & (!g3934)) + ((g1778) & (g1814) & (g3250) & (g3291) & (g3934)));
	assign g3949 = (((!g3235) & (!g3245) & (g3310) & (g3295) & (!g3936)) + ((!g3235) & (!g3245) & (g3310) & (g3295) & (g3936)) + ((!g3235) & (g3245) & (!g3310) & (g3295) & (!g3936)) + ((!g3235) & (g3245) & (g3310) & (!g3295) & (!g3936)) + ((!g3235) & (g3245) & (g3310) & (g3295) & (!g3936)) + ((!g3235) & (g3245) & (g3310) & (g3295) & (g3936)) + ((g3235) & (!g3245) & (!g3310) & (g3295) & (!g3936)) + ((g3235) & (!g3245) & (g3310) & (!g3295) & (!g3936)) + ((g3235) & (!g3245) & (g3310) & (g3295) & (!g3936)) + ((g3235) & (!g3245) & (g3310) & (g3295) & (g3936)) + ((g3235) & (g3245) & (!g3310) & (g3295) & (!g3936)) + ((g3235) & (g3245) & (!g3310) & (g3295) & (g3936)) + ((g3235) & (g3245) & (g3310) & (!g3295) & (!g3936)) + ((g3235) & (g3245) & (g3310) & (!g3295) & (g3936)) + ((g3235) & (g3245) & (g3310) & (g3295) & (!g3936)) + ((g3235) & (g3245) & (g3310) & (g3295) & (g3936)));
	assign g3950 = (((!g830) & (key[39]) & (!g1914) & (!g3948) & (!g3949) & (!g5672)) + ((!g830) & (key[39]) & (!g1914) & (!g3948) & (!g3949) & (g5672)) + ((!g830) & (key[39]) & (!g1914) & (!g3948) & (g3949) & (!g5672)) + ((!g830) & (key[39]) & (!g1914) & (!g3948) & (g3949) & (g5672)) + ((!g830) & (key[39]) & (!g1914) & (g3948) & (!g3949) & (!g5672)) + ((!g830) & (key[39]) & (!g1914) & (g3948) & (!g3949) & (g5672)) + ((!g830) & (key[39]) & (!g1914) & (g3948) & (g3949) & (!g5672)) + ((!g830) & (key[39]) & (!g1914) & (g3948) & (g3949) & (g5672)) + ((!g830) & (key[39]) & (g1914) & (!g3948) & (!g3949) & (!g5672)) + ((!g830) & (key[39]) & (g1914) & (!g3948) & (!g3949) & (g5672)) + ((!g830) & (key[39]) & (g1914) & (!g3948) & (g3949) & (!g5672)) + ((!g830) & (key[39]) & (g1914) & (!g3948) & (g3949) & (g5672)) + ((!g830) & (key[39]) & (g1914) & (g3948) & (!g3949) & (!g5672)) + ((!g830) & (key[39]) & (g1914) & (g3948) & (!g3949) & (g5672)) + ((!g830) & (key[39]) & (g1914) & (g3948) & (g3949) & (!g5672)) + ((!g830) & (key[39]) & (g1914) & (g3948) & (g3949) & (g5672)) + ((g830) & (!key[39]) & (!g1914) & (!g3948) & (!g3949) & (!g5672)) + ((g830) & (!key[39]) & (!g1914) & (!g3948) & (g3949) & (g5672)) + ((g830) & (!key[39]) & (!g1914) & (g3948) & (!g3949) & (!g5672)) + ((g830) & (!key[39]) & (!g1914) & (g3948) & (g3949) & (g5672)) + ((g830) & (!key[39]) & (g1914) & (!g3948) & (!g3949) & (!g5672)) + ((g830) & (!key[39]) & (g1914) & (!g3948) & (g3949) & (!g5672)) + ((g830) & (!key[39]) & (g1914) & (g3948) & (!g3949) & (g5672)) + ((g830) & (!key[39]) & (g1914) & (g3948) & (g3949) & (g5672)) + ((g830) & (key[39]) & (!g1914) & (!g3948) & (!g3949) & (!g5672)) + ((g830) & (key[39]) & (!g1914) & (!g3948) & (g3949) & (g5672)) + ((g830) & (key[39]) & (!g1914) & (g3948) & (!g3949) & (!g5672)) + ((g830) & (key[39]) & (!g1914) & (g3948) & (g3949) & (g5672)) + ((g830) & (key[39]) & (g1914) & (!g3948) & (!g3949) & (!g5672)) + ((g830) & (key[39]) & (g1914) & (!g3948) & (g3949) & (!g5672)) + ((g830) & (key[39]) & (g1914) & (g3948) & (!g3949) & (g5672)) + ((g830) & (key[39]) & (g1914) & (g3948) & (g3949) & (g5672)));
	assign g3951 = (((!g2515) & (g3106)) + ((g2515) & (!g3106)));
	assign g3952 = (((!g2376) & (!g2423) & (g3031) & (g3084) & (!g3930) & (g3951)) + ((!g2376) & (g2423) & (!g3031) & (g3084) & (!g3930) & (g3951)) + ((!g2376) & (g2423) & (!g3031) & (g3084) & (g3930) & (g3951)) + ((!g2376) & (g2423) & (g3031) & (!g3084) & (!g3930) & (g3951)) + ((!g2376) & (g2423) & (g3031) & (g3084) & (!g3930) & (g3951)) + ((!g2376) & (g2423) & (g3031) & (g3084) & (g3930) & (g3951)) + ((g2376) & (!g2423) & (!g3031) & (g3084) & (!g3930) & (g3951)) + ((g2376) & (!g2423) & (g3031) & (g3084) & (!g3930) & (g3951)) + ((g2376) & (!g2423) & (g3031) & (g3084) & (g3930) & (g3951)) + ((g2376) & (g2423) & (!g3031) & (!g3084) & (!g3930) & (g3951)) + ((g2376) & (g2423) & (!g3031) & (g3084) & (!g3930) & (g3951)) + ((g2376) & (g2423) & (!g3031) & (g3084) & (g3930) & (g3951)) + ((g2376) & (g2423) & (g3031) & (!g3084) & (!g3930) & (g3951)) + ((g2376) & (g2423) & (g3031) & (!g3084) & (g3930) & (g3951)) + ((g2376) & (g2423) & (g3031) & (g3084) & (!g3930) & (g3951)) + ((g2376) & (g2423) & (g3031) & (g3084) & (g3930) & (g3951)));
	assign g3953 = (((g2515) & (g3106)));
	assign g3954 = (((!g2551) & (!g3159) & (!g3952) & (g3953)) + ((!g2551) & (!g3159) & (g3952) & (!g3953)) + ((!g2551) & (!g3159) & (g3952) & (g3953)) + ((!g2551) & (g3159) & (!g3952) & (!g3953)) + ((g2551) & (!g3159) & (!g3952) & (!g3953)) + ((g2551) & (g3159) & (!g3952) & (g3953)) + ((g2551) & (g3159) & (g3952) & (!g3953)) + ((g2551) & (g3159) & (g3952) & (g3953)));
	assign g3955 = (((!g1847) & (!g1881) & (!g3339) & (g3366) & (!g3948)) + ((!g1847) & (!g1881) & (!g3339) & (g3366) & (g3948)) + ((!g1847) & (!g1881) & (g3339) & (!g3366) & (g3948)) + ((!g1847) & (!g1881) & (g3339) & (g3366) & (!g3948)) + ((!g1847) & (g1881) & (!g3339) & (!g3366) & (!g3948)) + ((!g1847) & (g1881) & (!g3339) & (!g3366) & (g3948)) + ((!g1847) & (g1881) & (g3339) & (!g3366) & (!g3948)) + ((!g1847) & (g1881) & (g3339) & (g3366) & (g3948)) + ((g1847) & (!g1881) & (!g3339) & (!g3366) & (g3948)) + ((g1847) & (!g1881) & (!g3339) & (g3366) & (!g3948)) + ((g1847) & (!g1881) & (g3339) & (!g3366) & (!g3948)) + ((g1847) & (!g1881) & (g3339) & (!g3366) & (g3948)) + ((g1847) & (g1881) & (!g3339) & (!g3366) & (!g3948)) + ((g1847) & (g1881) & (!g3339) & (g3366) & (g3948)) + ((g1847) & (g1881) & (g3339) & (g3366) & (!g3948)) + ((g1847) & (g1881) & (g3339) & (g3366) & (g3948)));
	assign g3956 = (((!g3330) & (!g3336) & (!g3385) & (g3370) & (!g3949)) + ((!g3330) & (!g3336) & (!g3385) & (g3370) & (g3949)) + ((!g3330) & (!g3336) & (g3385) & (!g3370) & (!g3949)) + ((!g3330) & (!g3336) & (g3385) & (!g3370) & (g3949)) + ((!g3330) & (g3336) & (!g3385) & (!g3370) & (g3949)) + ((!g3330) & (g3336) & (!g3385) & (g3370) & (!g3949)) + ((!g3330) & (g3336) & (g3385) & (!g3370) & (!g3949)) + ((!g3330) & (g3336) & (g3385) & (g3370) & (g3949)) + ((g3330) & (!g3336) & (!g3385) & (!g3370) & (g3949)) + ((g3330) & (!g3336) & (!g3385) & (g3370) & (!g3949)) + ((g3330) & (!g3336) & (g3385) & (!g3370) & (!g3949)) + ((g3330) & (!g3336) & (g3385) & (g3370) & (g3949)) + ((g3330) & (g3336) & (!g3385) & (!g3370) & (!g3949)) + ((g3330) & (g3336) & (!g3385) & (!g3370) & (g3949)) + ((g3330) & (g3336) & (g3385) & (g3370) & (!g3949)) + ((g3330) & (g3336) & (g3385) & (g3370) & (g3949)));
	assign g3957 = (((!g830) & (!g1914) & (!g1958) & (!g3955) & (!g3956) & (key[40])) + ((!g830) & (!g1914) & (!g1958) & (!g3955) & (g3956) & (key[40])) + ((!g830) & (!g1914) & (!g1958) & (g3955) & (!g3956) & (key[40])) + ((!g830) & (!g1914) & (!g1958) & (g3955) & (g3956) & (key[40])) + ((!g830) & (!g1914) & (g1958) & (!g3955) & (!g3956) & (key[40])) + ((!g830) & (!g1914) & (g1958) & (!g3955) & (g3956) & (key[40])) + ((!g830) & (!g1914) & (g1958) & (g3955) & (!g3956) & (key[40])) + ((!g830) & (!g1914) & (g1958) & (g3955) & (g3956) & (key[40])) + ((!g830) & (g1914) & (!g1958) & (!g3955) & (!g3956) & (key[40])) + ((!g830) & (g1914) & (!g1958) & (!g3955) & (g3956) & (key[40])) + ((!g830) & (g1914) & (!g1958) & (g3955) & (!g3956) & (key[40])) + ((!g830) & (g1914) & (!g1958) & (g3955) & (g3956) & (key[40])) + ((!g830) & (g1914) & (g1958) & (!g3955) & (!g3956) & (key[40])) + ((!g830) & (g1914) & (g1958) & (!g3955) & (g3956) & (key[40])) + ((!g830) & (g1914) & (g1958) & (g3955) & (!g3956) & (key[40])) + ((!g830) & (g1914) & (g1958) & (g3955) & (g3956) & (key[40])) + ((g830) & (!g1914) & (!g1958) & (!g3955) & (g3956) & (!key[40])) + ((g830) & (!g1914) & (!g1958) & (!g3955) & (g3956) & (key[40])) + ((g830) & (!g1914) & (!g1958) & (g3955) & (g3956) & (!key[40])) + ((g830) & (!g1914) & (!g1958) & (g3955) & (g3956) & (key[40])) + ((g830) & (!g1914) & (g1958) & (!g3955) & (!g3956) & (!key[40])) + ((g830) & (!g1914) & (g1958) & (!g3955) & (!g3956) & (key[40])) + ((g830) & (!g1914) & (g1958) & (g3955) & (!g3956) & (!key[40])) + ((g830) & (!g1914) & (g1958) & (g3955) & (!g3956) & (key[40])) + ((g830) & (g1914) & (!g1958) & (g3955) & (!g3956) & (!key[40])) + ((g830) & (g1914) & (!g1958) & (g3955) & (!g3956) & (key[40])) + ((g830) & (g1914) & (!g1958) & (g3955) & (g3956) & (!key[40])) + ((g830) & (g1914) & (!g1958) & (g3955) & (g3956) & (key[40])) + ((g830) & (g1914) & (g1958) & (!g3955) & (!g3956) & (!key[40])) + ((g830) & (g1914) & (g1958) & (!g3955) & (!g3956) & (key[40])) + ((g830) & (g1914) & (g1958) & (!g3955) & (g3956) & (!key[40])) + ((g830) & (g1914) & (g1958) & (!g3955) & (g3956) & (key[40])));
	assign g3958 = (((!g2551) & (!g3159) & (!g3952) & (!g3953)) + ((!g2551) & (!g3159) & (!g3952) & (g3953)) + ((!g2551) & (!g3159) & (g3952) & (!g3953)) + ((!g2551) & (!g3159) & (g3952) & (g3953)) + ((!g2551) & (g3159) & (!g3952) & (!g3953)) + ((g2551) & (!g3159) & (!g3952) & (!g3953)));
	assign g3959 = (((!g1908) & (!g2030) & (!g1912) & (g2045)) + ((!g1908) & (!g2030) & (g1912) & (g2045)) + ((!g1908) & (g2030) & (!g1912) & (!g2045)) + ((!g1908) & (g2030) & (g1912) & (!g2045)) + ((g1908) & (!g2030) & (!g1912) & (g2045)) + ((g1908) & (!g2030) & (g1912) & (!g2045)) + ((g1908) & (g2030) & (!g1912) & (!g2045)) + ((g1908) & (g2030) & (g1912) & (g2045)));
	assign g3960 = (((!g1914) & (!g2598) & (!g3177) & (!g3958) & (g3959)) + ((!g1914) & (!g2598) & (!g3177) & (g3958) & (g3959)) + ((!g1914) & (!g2598) & (g3177) & (!g3958) & (g3959)) + ((!g1914) & (!g2598) & (g3177) & (g3958) & (g3959)) + ((!g1914) & (g2598) & (!g3177) & (!g3958) & (g3959)) + ((!g1914) & (g2598) & (!g3177) & (g3958) & (g3959)) + ((!g1914) & (g2598) & (g3177) & (!g3958) & (g3959)) + ((!g1914) & (g2598) & (g3177) & (g3958) & (g3959)) + ((g1914) & (!g2598) & (!g3177) & (!g3958) & (!g3959)) + ((g1914) & (!g2598) & (!g3177) & (!g3958) & (g3959)) + ((g1914) & (!g2598) & (g3177) & (g3958) & (!g3959)) + ((g1914) & (!g2598) & (g3177) & (g3958) & (g3959)) + ((g1914) & (g2598) & (!g3177) & (g3958) & (!g3959)) + ((g1914) & (g2598) & (!g3177) & (g3958) & (g3959)) + ((g1914) & (g2598) & (g3177) & (!g3958) & (!g3959)) + ((g1914) & (g2598) & (g3177) & (!g3958) & (g3959)));
	assign g3961 = (((!g830) & (!g1959) & (!g3960) & (key[72])) + ((!g830) & (!g1959) & (g3960) & (key[72])) + ((!g830) & (g1959) & (!g3960) & (key[72])) + ((!g830) & (g1959) & (g3960) & (key[72])) + ((g830) & (!g1959) & (g3960) & (!key[72])) + ((g830) & (!g1959) & (g3960) & (key[72])) + ((g830) & (g1959) & (!g3960) & (!key[72])) + ((g830) & (g1959) & (!g3960) & (key[72])));
	assign g3962 = (((!g1914) & (!g828) & (!g1892) & (g1896) & (!g1898)) + ((!g1914) & (!g828) & (!g1892) & (g1896) & (g1898)) + ((!g1914) & (!g828) & (g1892) & (!g1896) & (!g1898)) + ((!g1914) & (!g828) & (g1892) & (!g1896) & (g1898)) + ((!g1914) & (g828) & (!g1892) & (g1896) & (!g1898)) + ((!g1914) & (g828) & (!g1892) & (g1896) & (g1898)) + ((!g1914) & (g828) & (g1892) & (!g1896) & (!g1898)) + ((!g1914) & (g828) & (g1892) & (!g1896) & (g1898)) + ((g1914) & (!g828) & (!g1892) & (!g1896) & (g1898)) + ((g1914) & (!g828) & (!g1892) & (g1896) & (g1898)) + ((g1914) & (!g828) & (g1892) & (!g1896) & (g1898)) + ((g1914) & (!g828) & (g1892) & (g1896) & (g1898)) + ((g1914) & (g828) & (!g1892) & (!g1896) & (!g1898)) + ((g1914) & (g828) & (!g1892) & (g1896) & (!g1898)) + ((g1914) & (g828) & (g1892) & (!g1896) & (!g1898)) + ((g1914) & (g828) & (g1892) & (g1896) & (!g1898)));
	assign g3963 = (((!g830) & (!g1960) & (!g3962) & (key[41])) + ((!g830) & (!g1960) & (g3962) & (key[41])) + ((!g830) & (g1960) & (!g3962) & (key[41])) + ((!g830) & (g1960) & (g3962) & (key[41])) + ((g830) & (!g1960) & (g3962) & (!key[41])) + ((g830) & (!g1960) & (g3962) & (key[41])) + ((g830) & (g1960) & (!g3962) & (!key[41])) + ((g830) & (g1960) & (!g3962) & (key[41])));
	assign g3964 = (((!g2551) & (!g2598) & (!g3159) & (!g3177) & (!g3952) & (!g3953)) + ((!g2551) & (!g2598) & (!g3159) & (!g3177) & (!g3952) & (g3953)) + ((!g2551) & (!g2598) & (!g3159) & (!g3177) & (g3952) & (!g3953)) + ((!g2551) & (!g2598) & (!g3159) & (!g3177) & (g3952) & (g3953)) + ((!g2551) & (!g2598) & (!g3159) & (g3177) & (!g3952) & (!g3953)) + ((!g2551) & (!g2598) & (!g3159) & (g3177) & (!g3952) & (g3953)) + ((!g2551) & (!g2598) & (!g3159) & (g3177) & (g3952) & (!g3953)) + ((!g2551) & (!g2598) & (!g3159) & (g3177) & (g3952) & (g3953)) + ((!g2551) & (!g2598) & (g3159) & (!g3177) & (!g3952) & (!g3953)) + ((!g2551) & (!g2598) & (g3159) & (!g3177) & (!g3952) & (g3953)) + ((!g2551) & (!g2598) & (g3159) & (!g3177) & (g3952) & (!g3953)) + ((!g2551) & (!g2598) & (g3159) & (!g3177) & (g3952) & (g3953)) + ((!g2551) & (!g2598) & (g3159) & (g3177) & (!g3952) & (!g3953)) + ((!g2551) & (g2598) & (!g3159) & (!g3177) & (!g3952) & (!g3953)) + ((!g2551) & (g2598) & (!g3159) & (!g3177) & (!g3952) & (g3953)) + ((!g2551) & (g2598) & (!g3159) & (!g3177) & (g3952) & (!g3953)) + ((!g2551) & (g2598) & (!g3159) & (!g3177) & (g3952) & (g3953)) + ((!g2551) & (g2598) & (g3159) & (!g3177) & (!g3952) & (!g3953)) + ((g2551) & (!g2598) & (!g3159) & (!g3177) & (!g3952) & (!g3953)) + ((g2551) & (!g2598) & (!g3159) & (!g3177) & (!g3952) & (g3953)) + ((g2551) & (!g2598) & (!g3159) & (!g3177) & (g3952) & (!g3953)) + ((g2551) & (!g2598) & (!g3159) & (!g3177) & (g3952) & (g3953)) + ((g2551) & (!g2598) & (!g3159) & (g3177) & (!g3952) & (!g3953)) + ((g2551) & (!g2598) & (g3159) & (!g3177) & (!g3952) & (!g3953)) + ((g2551) & (!g2598) & (g3159) & (!g3177) & (!g3952) & (g3953)) + ((g2551) & (!g2598) & (g3159) & (!g3177) & (g3952) & (!g3953)) + ((g2551) & (!g2598) & (g3159) & (!g3177) & (g3952) & (g3953)) + ((g2551) & (g2598) & (!g3159) & (!g3177) & (!g3952) & (!g3953)));
	assign g3965 = (((!g1908) & (!g2030) & (!g2085) & (!g1912) & (!g2045) & (g2091)) + ((!g1908) & (!g2030) & (!g2085) & (!g1912) & (g2045) & (g2091)) + ((!g1908) & (!g2030) & (!g2085) & (g1912) & (!g2045) & (g2091)) + ((!g1908) & (!g2030) & (!g2085) & (g1912) & (g2045) & (g2091)) + ((!g1908) & (!g2030) & (g2085) & (!g1912) & (!g2045) & (!g2091)) + ((!g1908) & (!g2030) & (g2085) & (!g1912) & (g2045) & (!g2091)) + ((!g1908) & (!g2030) & (g2085) & (g1912) & (!g2045) & (!g2091)) + ((!g1908) & (!g2030) & (g2085) & (g1912) & (g2045) & (!g2091)) + ((!g1908) & (g2030) & (!g2085) & (!g1912) & (!g2045) & (g2091)) + ((!g1908) & (g2030) & (!g2085) & (!g1912) & (g2045) & (!g2091)) + ((!g1908) & (g2030) & (!g2085) & (g1912) & (!g2045) & (g2091)) + ((!g1908) & (g2030) & (!g2085) & (g1912) & (g2045) & (!g2091)) + ((!g1908) & (g2030) & (g2085) & (!g1912) & (!g2045) & (!g2091)) + ((!g1908) & (g2030) & (g2085) & (!g1912) & (g2045) & (g2091)) + ((!g1908) & (g2030) & (g2085) & (g1912) & (!g2045) & (!g2091)) + ((!g1908) & (g2030) & (g2085) & (g1912) & (g2045) & (g2091)) + ((g1908) & (!g2030) & (!g2085) & (!g1912) & (!g2045) & (g2091)) + ((g1908) & (!g2030) & (!g2085) & (!g1912) & (g2045) & (g2091)) + ((g1908) & (!g2030) & (!g2085) & (g1912) & (!g2045) & (g2091)) + ((g1908) & (!g2030) & (!g2085) & (g1912) & (g2045) & (!g2091)) + ((g1908) & (!g2030) & (g2085) & (!g1912) & (!g2045) & (!g2091)) + ((g1908) & (!g2030) & (g2085) & (!g1912) & (g2045) & (!g2091)) + ((g1908) & (!g2030) & (g2085) & (g1912) & (!g2045) & (!g2091)) + ((g1908) & (!g2030) & (g2085) & (g1912) & (g2045) & (g2091)) + ((g1908) & (g2030) & (!g2085) & (!g1912) & (!g2045) & (g2091)) + ((g1908) & (g2030) & (!g2085) & (!g1912) & (g2045) & (!g2091)) + ((g1908) & (g2030) & (!g2085) & (g1912) & (!g2045) & (!g2091)) + ((g1908) & (g2030) & (!g2085) & (g1912) & (g2045) & (!g2091)) + ((g1908) & (g2030) & (g2085) & (!g1912) & (!g2045) & (!g2091)) + ((g1908) & (g2030) & (g2085) & (!g1912) & (g2045) & (g2091)) + ((g1908) & (g2030) & (g2085) & (g1912) & (!g2045) & (g2091)) + ((g1908) & (g2030) & (g2085) & (g1912) & (g2045) & (g2091)));
	assign g3966 = (((!g1914) & (!g2647) & (!g3250) & (!g3964) & (g3965)) + ((!g1914) & (!g2647) & (!g3250) & (g3964) & (g3965)) + ((!g1914) & (!g2647) & (g3250) & (!g3964) & (g3965)) + ((!g1914) & (!g2647) & (g3250) & (g3964) & (g3965)) + ((!g1914) & (g2647) & (!g3250) & (!g3964) & (g3965)) + ((!g1914) & (g2647) & (!g3250) & (g3964) & (g3965)) + ((!g1914) & (g2647) & (g3250) & (!g3964) & (g3965)) + ((!g1914) & (g2647) & (g3250) & (g3964) & (g3965)) + ((g1914) & (!g2647) & (!g3250) & (!g3964) & (!g3965)) + ((g1914) & (!g2647) & (!g3250) & (!g3964) & (g3965)) + ((g1914) & (!g2647) & (g3250) & (g3964) & (!g3965)) + ((g1914) & (!g2647) & (g3250) & (g3964) & (g3965)) + ((g1914) & (g2647) & (!g3250) & (g3964) & (!g3965)) + ((g1914) & (g2647) & (!g3250) & (g3964) & (g3965)) + ((g1914) & (g2647) & (g3250) & (!g3964) & (!g3965)) + ((g1914) & (g2647) & (g3250) & (!g3964) & (g3965)));
	assign g3967 = (((!g830) & (!g1961) & (!g3966) & (key[73])) + ((!g830) & (!g1961) & (g3966) & (key[73])) + ((!g830) & (g1961) & (!g3966) & (key[73])) + ((!g830) & (g1961) & (g3966) & (key[73])) + ((g830) & (!g1961) & (g3966) & (!key[73])) + ((g830) & (!g1961) & (g3966) & (key[73])) + ((g830) & (g1961) & (!g3966) & (!key[73])) + ((g830) & (g1961) & (!g3966) & (key[73])));
	assign g3968 = (((g1914) & (!g828) & (!g864) & (!g1898) & (g2022)) + ((g1914) & (!g828) & (!g864) & (g1898) & (g2022)) + ((g1914) & (!g828) & (g864) & (!g1898) & (!g2022)) + ((g1914) & (!g828) & (g864) & (g1898) & (!g2022)) + ((g1914) & (g828) & (!g864) & (!g1898) & (g2022)) + ((g1914) & (g828) & (!g864) & (g1898) & (!g2022)) + ((g1914) & (g828) & (g864) & (!g1898) & (!g2022)) + ((g1914) & (g828) & (g864) & (g1898) & (g2022)));
	assign g3969 = (((!g1914) & (!g1892) & (!g2026) & (!g1896) & (g2041)) + ((!g1914) & (!g1892) & (!g2026) & (g1896) & (g2041)) + ((!g1914) & (!g1892) & (g2026) & (!g1896) & (!g2041)) + ((!g1914) & (!g1892) & (g2026) & (g1896) & (!g2041)) + ((!g1914) & (g1892) & (!g2026) & (!g1896) & (g2041)) + ((!g1914) & (g1892) & (!g2026) & (g1896) & (!g2041)) + ((!g1914) & (g1892) & (g2026) & (!g1896) & (!g2041)) + ((!g1914) & (g1892) & (g2026) & (g1896) & (g2041)));
	assign g3970 = (((!g830) & (!g1962) & (!g3968) & (!g3969) & (key[42])) + ((!g830) & (!g1962) & (!g3968) & (g3969) & (key[42])) + ((!g830) & (!g1962) & (g3968) & (!g3969) & (key[42])) + ((!g830) & (!g1962) & (g3968) & (g3969) & (key[42])) + ((!g830) & (g1962) & (!g3968) & (!g3969) & (key[42])) + ((!g830) & (g1962) & (!g3968) & (g3969) & (key[42])) + ((!g830) & (g1962) & (g3968) & (!g3969) & (key[42])) + ((!g830) & (g1962) & (g3968) & (g3969) & (key[42])) + ((g830) & (!g1962) & (!g3968) & (g3969) & (!key[42])) + ((g830) & (!g1962) & (!g3968) & (g3969) & (key[42])) + ((g830) & (!g1962) & (g3968) & (!g3969) & (!key[42])) + ((g830) & (!g1962) & (g3968) & (!g3969) & (key[42])) + ((g830) & (!g1962) & (g3968) & (g3969) & (!key[42])) + ((g830) & (!g1962) & (g3968) & (g3969) & (key[42])) + ((g830) & (g1962) & (!g3968) & (!g3969) & (!key[42])) + ((g830) & (g1962) & (!g3968) & (!g3969) & (key[42])));
	assign g3971 = (((!g2647) & (!g2678) & (!g3250) & (g3291) & (!g3964)) + ((!g2647) & (!g2678) & (!g3250) & (g3291) & (g3964)) + ((!g2647) & (!g2678) & (g3250) & (!g3291) & (!g3964)) + ((!g2647) & (!g2678) & (g3250) & (g3291) & (g3964)) + ((!g2647) & (g2678) & (!g3250) & (!g3291) & (!g3964)) + ((!g2647) & (g2678) & (!g3250) & (!g3291) & (g3964)) + ((!g2647) & (g2678) & (g3250) & (!g3291) & (g3964)) + ((!g2647) & (g2678) & (g3250) & (g3291) & (!g3964)) + ((g2647) & (!g2678) & (!g3250) & (!g3291) & (!g3964)) + ((g2647) & (!g2678) & (!g3250) & (g3291) & (g3964)) + ((g2647) & (!g2678) & (g3250) & (!g3291) & (!g3964)) + ((g2647) & (!g2678) & (g3250) & (!g3291) & (g3964)) + ((g2647) & (g2678) & (!g3250) & (!g3291) & (g3964)) + ((g2647) & (g2678) & (!g3250) & (g3291) & (!g3964)) + ((g2647) & (g2678) & (g3250) & (g3291) & (!g3964)) + ((g2647) & (g2678) & (g3250) & (g3291) & (g3964)));
	assign g3972 = (((!g2112) & (!g2127) & (g3759)) + ((!g2112) & (g2127) & (!g3759)) + ((g2112) & (!g2127) & (!g3759)) + ((g2112) & (g2127) & (g3759)));
	assign g3973 = (((!g830) & (!g1914) & (!g1963) & (!g3971) & (!g3972) & (key[74])) + ((!g830) & (!g1914) & (!g1963) & (!g3971) & (g3972) & (key[74])) + ((!g830) & (!g1914) & (!g1963) & (g3971) & (!g3972) & (key[74])) + ((!g830) & (!g1914) & (!g1963) & (g3971) & (g3972) & (key[74])) + ((!g830) & (!g1914) & (g1963) & (!g3971) & (!g3972) & (key[74])) + ((!g830) & (!g1914) & (g1963) & (!g3971) & (g3972) & (key[74])) + ((!g830) & (!g1914) & (g1963) & (g3971) & (!g3972) & (key[74])) + ((!g830) & (!g1914) & (g1963) & (g3971) & (g3972) & (key[74])) + ((!g830) & (g1914) & (!g1963) & (!g3971) & (!g3972) & (key[74])) + ((!g830) & (g1914) & (!g1963) & (!g3971) & (g3972) & (key[74])) + ((!g830) & (g1914) & (!g1963) & (g3971) & (!g3972) & (key[74])) + ((!g830) & (g1914) & (!g1963) & (g3971) & (g3972) & (key[74])) + ((!g830) & (g1914) & (g1963) & (!g3971) & (!g3972) & (key[74])) + ((!g830) & (g1914) & (g1963) & (!g3971) & (g3972) & (key[74])) + ((!g830) & (g1914) & (g1963) & (g3971) & (!g3972) & (key[74])) + ((!g830) & (g1914) & (g1963) & (g3971) & (g3972) & (key[74])) + ((g830) & (!g1914) & (!g1963) & (!g3971) & (g3972) & (!key[74])) + ((g830) & (!g1914) & (!g1963) & (!g3971) & (g3972) & (key[74])) + ((g830) & (!g1914) & (!g1963) & (g3971) & (g3972) & (!key[74])) + ((g830) & (!g1914) & (!g1963) & (g3971) & (g3972) & (key[74])) + ((g830) & (!g1914) & (g1963) & (!g3971) & (!g3972) & (!key[74])) + ((g830) & (!g1914) & (g1963) & (!g3971) & (!g3972) & (key[74])) + ((g830) & (!g1914) & (g1963) & (g3971) & (!g3972) & (!key[74])) + ((g830) & (!g1914) & (g1963) & (g3971) & (!g3972) & (key[74])) + ((g830) & (g1914) & (!g1963) & (g3971) & (!g3972) & (!key[74])) + ((g830) & (g1914) & (!g1963) & (g3971) & (!g3972) & (key[74])) + ((g830) & (g1914) & (!g1963) & (g3971) & (g3972) & (!key[74])) + ((g830) & (g1914) & (!g1963) & (g3971) & (g3972) & (key[74])) + ((g830) & (g1914) & (g1963) & (!g3971) & (!g3972) & (!key[74])) + ((g830) & (g1914) & (g1963) & (!g3971) & (!g3972) & (key[74])) + ((g830) & (g1914) & (g1963) & (!g3971) & (g3972) & (!key[74])) + ((g830) & (g1914) & (g1963) & (!g3971) & (g3972) & (key[74])));
	assign g3974 = (((!g828) & (g864) & (!g1898) & (g2022)) + ((!g828) & (g864) & (g1898) & (g2022)) + ((g828) & (!g864) & (g1898) & (g2022)) + ((g828) & (g864) & (!g1898) & (g2022)) + ((g828) & (g864) & (g1898) & (!g2022)) + ((g828) & (g864) & (g1898) & (g2022)));
	assign g3975 = (((g1914) & (!g897) & (!g3974) & (g2071)) + ((g1914) & (!g897) & (g3974) & (!g2071)) + ((g1914) & (g897) & (!g3974) & (!g2071)) + ((g1914) & (g897) & (g3974) & (g2071)));
	assign g3976 = (((!g1892) & (g2026) & (!g1896) & (g2041)) + ((!g1892) & (g2026) & (g1896) & (g2041)) + ((g1892) & (!g2026) & (g1896) & (g2041)) + ((g1892) & (g2026) & (!g1896) & (g2041)) + ((g1892) & (g2026) & (g1896) & (!g2041)) + ((g1892) & (g2026) & (g1896) & (g2041)));
	assign g3977 = (((!g1914) & (!g2062) & (!g2068) & (g3976)) + ((!g1914) & (!g2062) & (g2068) & (!g3976)) + ((!g1914) & (g2062) & (!g2068) & (!g3976)) + ((!g1914) & (g2062) & (g2068) & (g3976)));
	assign g3978 = (((!g830) & (!g1967) & (!g3975) & (!g3977) & (key[43])) + ((!g830) & (!g1967) & (!g3975) & (g3977) & (key[43])) + ((!g830) & (!g1967) & (g3975) & (!g3977) & (key[43])) + ((!g830) & (!g1967) & (g3975) & (g3977) & (key[43])) + ((!g830) & (g1967) & (!g3975) & (!g3977) & (key[43])) + ((!g830) & (g1967) & (!g3975) & (g3977) & (key[43])) + ((!g830) & (g1967) & (g3975) & (!g3977) & (key[43])) + ((!g830) & (g1967) & (g3975) & (g3977) & (key[43])) + ((g830) & (!g1967) & (!g3975) & (g3977) & (!key[43])) + ((g830) & (!g1967) & (!g3975) & (g3977) & (key[43])) + ((g830) & (!g1967) & (g3975) & (!g3977) & (!key[43])) + ((g830) & (!g1967) & (g3975) & (!g3977) & (key[43])) + ((g830) & (!g1967) & (g3975) & (g3977) & (!key[43])) + ((g830) & (!g1967) & (g3975) & (g3977) & (key[43])) + ((g830) & (g1967) & (!g3975) & (!g3977) & (!key[43])) + ((g830) & (g1967) & (!g3975) & (!g3977) & (key[43])));
	assign g3979 = (((!g2647) & (!g2678) & (g3250) & (g3291) & (!g3964)) + ((!g2647) & (g2678) & (!g3250) & (g3291) & (!g3964)) + ((!g2647) & (g2678) & (!g3250) & (g3291) & (g3964)) + ((!g2647) & (g2678) & (g3250) & (!g3291) & (!g3964)) + ((!g2647) & (g2678) & (g3250) & (g3291) & (!g3964)) + ((!g2647) & (g2678) & (g3250) & (g3291) & (g3964)) + ((g2647) & (!g2678) & (!g3250) & (g3291) & (!g3964)) + ((g2647) & (!g2678) & (g3250) & (g3291) & (!g3964)) + ((g2647) & (!g2678) & (g3250) & (g3291) & (g3964)) + ((g2647) & (g2678) & (!g3250) & (!g3291) & (!g3964)) + ((g2647) & (g2678) & (!g3250) & (g3291) & (!g3964)) + ((g2647) & (g2678) & (!g3250) & (g3291) & (g3964)) + ((g2647) & (g2678) & (g3250) & (!g3291) & (!g3964)) + ((g2647) & (g2678) & (g3250) & (!g3291) & (g3964)) + ((g2647) & (g2678) & (g3250) & (g3291) & (!g3964)) + ((g2647) & (g2678) & (g3250) & (g3291) & (g3964)));
	assign g3980 = (((!g2112) & (g2127) & (g3759)) + ((g2112) & (!g2127) & (g3759)) + ((g2112) & (g2127) & (!g3759)) + ((g2112) & (g2127) & (g3759)));
	assign g3981 = (((!g830) & (key[75]) & (!g1914) & (!g3979) & (!g2167) & (!g5677)) + ((!g830) & (key[75]) & (!g1914) & (!g3979) & (!g2167) & (g5677)) + ((!g830) & (key[75]) & (!g1914) & (!g3979) & (g2167) & (!g5677)) + ((!g830) & (key[75]) & (!g1914) & (!g3979) & (g2167) & (g5677)) + ((!g830) & (key[75]) & (!g1914) & (g3979) & (!g2167) & (!g5677)) + ((!g830) & (key[75]) & (!g1914) & (g3979) & (!g2167) & (g5677)) + ((!g830) & (key[75]) & (!g1914) & (g3979) & (g2167) & (!g5677)) + ((!g830) & (key[75]) & (!g1914) & (g3979) & (g2167) & (g5677)) + ((!g830) & (key[75]) & (g1914) & (!g3979) & (!g2167) & (!g5677)) + ((!g830) & (key[75]) & (g1914) & (!g3979) & (!g2167) & (g5677)) + ((!g830) & (key[75]) & (g1914) & (!g3979) & (g2167) & (!g5677)) + ((!g830) & (key[75]) & (g1914) & (!g3979) & (g2167) & (g5677)) + ((!g830) & (key[75]) & (g1914) & (g3979) & (!g2167) & (!g5677)) + ((!g830) & (key[75]) & (g1914) & (g3979) & (!g2167) & (g5677)) + ((!g830) & (key[75]) & (g1914) & (g3979) & (g2167) & (!g5677)) + ((!g830) & (key[75]) & (g1914) & (g3979) & (g2167) & (g5677)) + ((g830) & (!key[75]) & (!g1914) & (!g3979) & (!g2167) & (!g5677)) + ((g830) & (!key[75]) & (!g1914) & (!g3979) & (g2167) & (g5677)) + ((g830) & (!key[75]) & (!g1914) & (g3979) & (!g2167) & (!g5677)) + ((g830) & (!key[75]) & (!g1914) & (g3979) & (g2167) & (g5677)) + ((g830) & (!key[75]) & (g1914) & (!g3979) & (!g2167) & (!g5677)) + ((g830) & (!key[75]) & (g1914) & (!g3979) & (g2167) & (!g5677)) + ((g830) & (!key[75]) & (g1914) & (g3979) & (!g2167) & (g5677)) + ((g830) & (!key[75]) & (g1914) & (g3979) & (g2167) & (g5677)) + ((g830) & (key[75]) & (!g1914) & (!g3979) & (!g2167) & (!g5677)) + ((g830) & (key[75]) & (!g1914) & (!g3979) & (g2167) & (g5677)) + ((g830) & (key[75]) & (!g1914) & (g3979) & (!g2167) & (!g5677)) + ((g830) & (key[75]) & (!g1914) & (g3979) & (g2167) & (g5677)) + ((g830) & (key[75]) & (g1914) & (!g3979) & (!g2167) & (!g5677)) + ((g830) & (key[75]) & (g1914) & (!g3979) & (g2167) & (!g5677)) + ((g830) & (key[75]) & (g1914) & (g3979) & (!g2167) & (g5677)) + ((g830) & (key[75]) & (g1914) & (g3979) & (g2167) & (g5677)));
	assign g3982 = (((!g931) & (!g3500) & (g2104)) + ((!g931) & (g3500) & (!g2104)) + ((g931) & (!g3500) & (!g2104)) + ((g931) & (g3500) & (g2104)));
	assign g3983 = (((!g2108) & (!g2123) & (g3517)) + ((!g2108) & (g2123) & (!g3517)) + ((g2108) & (!g2123) & (!g3517)) + ((g2108) & (g2123) & (g3517)));
	assign g3984 = (((!g830) & (!g1914) & (!g1969) & (!g3982) & (!g3983) & (key[44])) + ((!g830) & (!g1914) & (!g1969) & (!g3982) & (g3983) & (key[44])) + ((!g830) & (!g1914) & (!g1969) & (g3982) & (!g3983) & (key[44])) + ((!g830) & (!g1914) & (!g1969) & (g3982) & (g3983) & (key[44])) + ((!g830) & (!g1914) & (g1969) & (!g3982) & (!g3983) & (key[44])) + ((!g830) & (!g1914) & (g1969) & (!g3982) & (g3983) & (key[44])) + ((!g830) & (!g1914) & (g1969) & (g3982) & (!g3983) & (key[44])) + ((!g830) & (!g1914) & (g1969) & (g3982) & (g3983) & (key[44])) + ((!g830) & (g1914) & (!g1969) & (!g3982) & (!g3983) & (key[44])) + ((!g830) & (g1914) & (!g1969) & (!g3982) & (g3983) & (key[44])) + ((!g830) & (g1914) & (!g1969) & (g3982) & (!g3983) & (key[44])) + ((!g830) & (g1914) & (!g1969) & (g3982) & (g3983) & (key[44])) + ((!g830) & (g1914) & (g1969) & (!g3982) & (!g3983) & (key[44])) + ((!g830) & (g1914) & (g1969) & (!g3982) & (g3983) & (key[44])) + ((!g830) & (g1914) & (g1969) & (g3982) & (!g3983) & (key[44])) + ((!g830) & (g1914) & (g1969) & (g3982) & (g3983) & (key[44])) + ((g830) & (!g1914) & (!g1969) & (!g3982) & (g3983) & (!key[44])) + ((g830) & (!g1914) & (!g1969) & (!g3982) & (g3983) & (key[44])) + ((g830) & (!g1914) & (!g1969) & (g3982) & (g3983) & (!key[44])) + ((g830) & (!g1914) & (!g1969) & (g3982) & (g3983) & (key[44])) + ((g830) & (!g1914) & (g1969) & (!g3982) & (!g3983) & (!key[44])) + ((g830) & (!g1914) & (g1969) & (!g3982) & (!g3983) & (key[44])) + ((g830) & (!g1914) & (g1969) & (g3982) & (!g3983) & (!key[44])) + ((g830) & (!g1914) & (g1969) & (g3982) & (!g3983) & (key[44])) + ((g830) & (g1914) & (!g1969) & (g3982) & (!g3983) & (!key[44])) + ((g830) & (g1914) & (!g1969) & (g3982) & (!g3983) & (key[44])) + ((g830) & (g1914) & (!g1969) & (g3982) & (g3983) & (!key[44])) + ((g830) & (g1914) & (!g1969) & (g3982) & (g3983) & (key[44])) + ((g830) & (g1914) & (g1969) & (!g3982) & (!g3983) & (!key[44])) + ((g830) & (g1914) & (g1969) & (!g3982) & (!g3983) & (key[44])) + ((g830) & (g1914) & (g1969) & (!g3982) & (g3983) & (!key[44])) + ((g830) & (g1914) & (g1969) & (!g3982) & (g3983) & (key[44])));
	assign g3985 = (((!g931) & (g3500) & (g2104)) + ((g931) & (!g3500) & (g2104)) + ((g931) & (g3500) & (!g2104)) + ((g931) & (g3500) & (g2104)));
	assign g3986 = (((g1914) & (!g964) & (!g3985) & (g2153)) + ((g1914) & (!g964) & (g3985) & (!g2153)) + ((g1914) & (g964) & (!g3985) & (!g2153)) + ((g1914) & (g964) & (g3985) & (g2153)));
	assign g3987 = (((!g2108) & (g2123) & (g3517)) + ((g2108) & (!g2123) & (g3517)) + ((g2108) & (g2123) & (!g3517)) + ((g2108) & (g2123) & (g3517)));
	assign g3988 = (((!g1914) & (!g2144) & (!g2150) & (g3987)) + ((!g1914) & (!g2144) & (g2150) & (!g3987)) + ((!g1914) & (g2144) & (!g2150) & (!g3987)) + ((!g1914) & (g2144) & (g2150) & (g3987)));
	assign g3989 = (((!g830) & (!g1972) & (!g3986) & (!g3988) & (key[45])) + ((!g830) & (!g1972) & (!g3986) & (g3988) & (key[45])) + ((!g830) & (!g1972) & (g3986) & (!g3988) & (key[45])) + ((!g830) & (!g1972) & (g3986) & (g3988) & (key[45])) + ((!g830) & (g1972) & (!g3986) & (!g3988) & (key[45])) + ((!g830) & (g1972) & (!g3986) & (g3988) & (key[45])) + ((!g830) & (g1972) & (g3986) & (!g3988) & (key[45])) + ((!g830) & (g1972) & (g3986) & (g3988) & (key[45])) + ((g830) & (!g1972) & (!g3986) & (g3988) & (!key[45])) + ((g830) & (!g1972) & (!g3986) & (g3988) & (key[45])) + ((g830) & (!g1972) & (g3986) & (!g3988) & (!key[45])) + ((g830) & (!g1972) & (g3986) & (!g3988) & (key[45])) + ((g830) & (!g1972) & (g3986) & (g3988) & (!key[45])) + ((g830) & (!g1972) & (g3986) & (g3988) & (key[45])) + ((g830) & (g1972) & (!g3986) & (!g3988) & (!key[45])) + ((g830) & (g1972) & (!g3986) & (!g3988) & (key[45])));
	assign g3990 = (((!g3761) & (g3762)) + ((g3761) & (!g3762)) + ((g3761) & (g3762)));
	assign g3991 = (((!g1914) & (!g1890) & (!g2247) & (!g2253) & (!g1898) & (g3990)) + ((!g1914) & (!g1890) & (!g2247) & (!g2253) & (g1898) & (g3990)) + ((!g1914) & (!g1890) & (!g2247) & (g2253) & (!g1898) & (!g3990)) + ((!g1914) & (!g1890) & (!g2247) & (g2253) & (g1898) & (!g3990)) + ((!g1914) & (!g1890) & (g2247) & (!g2253) & (!g1898) & (!g3990)) + ((!g1914) & (!g1890) & (g2247) & (!g2253) & (g1898) & (!g3990)) + ((!g1914) & (!g1890) & (g2247) & (g2253) & (!g1898) & (g3990)) + ((!g1914) & (!g1890) & (g2247) & (g2253) & (g1898) & (g3990)) + ((!g1914) & (g1890) & (!g2247) & (!g2253) & (!g1898) & (g3990)) + ((!g1914) & (g1890) & (!g2247) & (!g2253) & (g1898) & (g3990)) + ((!g1914) & (g1890) & (!g2247) & (g2253) & (!g1898) & (!g3990)) + ((!g1914) & (g1890) & (!g2247) & (g2253) & (g1898) & (!g3990)) + ((!g1914) & (g1890) & (g2247) & (!g2253) & (!g1898) & (!g3990)) + ((!g1914) & (g1890) & (g2247) & (!g2253) & (g1898) & (!g3990)) + ((!g1914) & (g1890) & (g2247) & (g2253) & (!g1898) & (g3990)) + ((!g1914) & (g1890) & (g2247) & (g2253) & (g1898) & (g3990)) + ((g1914) & (!g1890) & (!g2247) & (!g2253) & (g1898) & (!g3990)) + ((g1914) & (!g1890) & (!g2247) & (!g2253) & (g1898) & (g3990)) + ((g1914) & (!g1890) & (!g2247) & (g2253) & (g1898) & (!g3990)) + ((g1914) & (!g1890) & (!g2247) & (g2253) & (g1898) & (g3990)) + ((g1914) & (!g1890) & (g2247) & (!g2253) & (g1898) & (!g3990)) + ((g1914) & (!g1890) & (g2247) & (!g2253) & (g1898) & (g3990)) + ((g1914) & (!g1890) & (g2247) & (g2253) & (g1898) & (!g3990)) + ((g1914) & (!g1890) & (g2247) & (g2253) & (g1898) & (g3990)) + ((g1914) & (g1890) & (!g2247) & (!g2253) & (!g1898) & (!g3990)) + ((g1914) & (g1890) & (!g2247) & (!g2253) & (!g1898) & (g3990)) + ((g1914) & (g1890) & (!g2247) & (g2253) & (!g1898) & (!g3990)) + ((g1914) & (g1890) & (!g2247) & (g2253) & (!g1898) & (g3990)) + ((g1914) & (g1890) & (g2247) & (!g2253) & (!g1898) & (!g3990)) + ((g1914) & (g1890) & (g2247) & (!g2253) & (!g1898) & (g3990)) + ((g1914) & (g1890) & (g2247) & (g2253) & (!g1898) & (!g3990)) + ((g1914) & (g1890) & (g2247) & (g2253) & (!g1898) & (g3990)));
	assign g3992 = (((!g830) & (!g1973) & (!g3991) & (key[77])) + ((!g830) & (!g1973) & (g3991) & (key[77])) + ((!g830) & (g1973) & (!g3991) & (key[77])) + ((!g830) & (g1973) & (g3991) & (key[77])) + ((g830) & (!g1973) & (g3991) & (!key[77])) + ((g830) & (!g1973) & (g3991) & (key[77])) + ((g830) & (g1973) & (!g3991) & (!key[77])) + ((g830) & (g1973) & (!g3991) & (key[77])));
	assign g3993 = (((!g964) & (!g998) & (!g3985) & (!g2153) & (g2184)) + ((!g964) & (!g998) & (!g3985) & (g2153) & (g2184)) + ((!g964) & (!g998) & (g3985) & (!g2153) & (g2184)) + ((!g964) & (!g998) & (g3985) & (g2153) & (!g2184)) + ((!g964) & (g998) & (!g3985) & (!g2153) & (!g2184)) + ((!g964) & (g998) & (!g3985) & (g2153) & (!g2184)) + ((!g964) & (g998) & (g3985) & (!g2153) & (!g2184)) + ((!g964) & (g998) & (g3985) & (g2153) & (g2184)) + ((g964) & (!g998) & (!g3985) & (!g2153) & (g2184)) + ((g964) & (!g998) & (!g3985) & (g2153) & (!g2184)) + ((g964) & (!g998) & (g3985) & (!g2153) & (!g2184)) + ((g964) & (!g998) & (g3985) & (g2153) & (!g2184)) + ((g964) & (g998) & (!g3985) & (!g2153) & (!g2184)) + ((g964) & (g998) & (!g3985) & (g2153) & (g2184)) + ((g964) & (g998) & (g3985) & (!g2153) & (g2184)) + ((g964) & (g998) & (g3985) & (g2153) & (g2184)));
	assign g3994 = (((!g2144) & (!g2188) & (!g2150) & (g2203) & (!g3987)) + ((!g2144) & (!g2188) & (!g2150) & (g2203) & (g3987)) + ((!g2144) & (!g2188) & (g2150) & (!g2203) & (g3987)) + ((!g2144) & (!g2188) & (g2150) & (g2203) & (!g3987)) + ((!g2144) & (g2188) & (!g2150) & (!g2203) & (!g3987)) + ((!g2144) & (g2188) & (!g2150) & (!g2203) & (g3987)) + ((!g2144) & (g2188) & (g2150) & (!g2203) & (!g3987)) + ((!g2144) & (g2188) & (g2150) & (g2203) & (g3987)) + ((g2144) & (!g2188) & (!g2150) & (!g2203) & (g3987)) + ((g2144) & (!g2188) & (!g2150) & (g2203) & (!g3987)) + ((g2144) & (!g2188) & (g2150) & (!g2203) & (!g3987)) + ((g2144) & (!g2188) & (g2150) & (!g2203) & (g3987)) + ((g2144) & (g2188) & (!g2150) & (!g2203) & (!g3987)) + ((g2144) & (g2188) & (!g2150) & (g2203) & (g3987)) + ((g2144) & (g2188) & (g2150) & (g2203) & (!g3987)) + ((g2144) & (g2188) & (g2150) & (g2203) & (g3987)));
	assign g3995 = (((!g830) & (!g1914) & (!g1975) & (!g3993) & (!g3994) & (key[46])) + ((!g830) & (!g1914) & (!g1975) & (!g3993) & (g3994) & (key[46])) + ((!g830) & (!g1914) & (!g1975) & (g3993) & (!g3994) & (key[46])) + ((!g830) & (!g1914) & (!g1975) & (g3993) & (g3994) & (key[46])) + ((!g830) & (!g1914) & (g1975) & (!g3993) & (!g3994) & (key[46])) + ((!g830) & (!g1914) & (g1975) & (!g3993) & (g3994) & (key[46])) + ((!g830) & (!g1914) & (g1975) & (g3993) & (!g3994) & (key[46])) + ((!g830) & (!g1914) & (g1975) & (g3993) & (g3994) & (key[46])) + ((!g830) & (g1914) & (!g1975) & (!g3993) & (!g3994) & (key[46])) + ((!g830) & (g1914) & (!g1975) & (!g3993) & (g3994) & (key[46])) + ((!g830) & (g1914) & (!g1975) & (g3993) & (!g3994) & (key[46])) + ((!g830) & (g1914) & (!g1975) & (g3993) & (g3994) & (key[46])) + ((!g830) & (g1914) & (g1975) & (!g3993) & (!g3994) & (key[46])) + ((!g830) & (g1914) & (g1975) & (!g3993) & (g3994) & (key[46])) + ((!g830) & (g1914) & (g1975) & (g3993) & (!g3994) & (key[46])) + ((!g830) & (g1914) & (g1975) & (g3993) & (g3994) & (key[46])) + ((g830) & (!g1914) & (!g1975) & (!g3993) & (g3994) & (!key[46])) + ((g830) & (!g1914) & (!g1975) & (!g3993) & (g3994) & (key[46])) + ((g830) & (!g1914) & (!g1975) & (g3993) & (g3994) & (!key[46])) + ((g830) & (!g1914) & (!g1975) & (g3993) & (g3994) & (key[46])) + ((g830) & (!g1914) & (g1975) & (!g3993) & (!g3994) & (!key[46])) + ((g830) & (!g1914) & (g1975) & (!g3993) & (!g3994) & (key[46])) + ((g830) & (!g1914) & (g1975) & (g3993) & (!g3994) & (!key[46])) + ((g830) & (!g1914) & (g1975) & (g3993) & (!g3994) & (key[46])) + ((g830) & (g1914) & (!g1975) & (g3993) & (!g3994) & (!key[46])) + ((g830) & (g1914) & (!g1975) & (g3993) & (!g3994) & (key[46])) + ((g830) & (g1914) & (!g1975) & (g3993) & (g3994) & (!key[46])) + ((g830) & (g1914) & (!g1975) & (g3993) & (g3994) & (key[46])) + ((g830) & (g1914) & (g1975) & (!g3993) & (!g3994) & (!key[46])) + ((g830) & (g1914) & (g1975) & (!g3993) & (!g3994) & (key[46])) + ((g830) & (g1914) & (g1975) & (!g3993) & (g3994) & (!key[46])) + ((g830) & (g1914) & (g1975) & (!g3993) & (g3994) & (key[46])));
	assign g3996 = (((!g1890) & (!g1939) & (!g1898) & (g2022)) + ((!g1890) & (!g1939) & (g1898) & (g2022)) + ((!g1890) & (g1939) & (!g1898) & (!g2022)) + ((!g1890) & (g1939) & (g1898) & (!g2022)) + ((g1890) & (!g1939) & (!g1898) & (g2022)) + ((g1890) & (!g1939) & (g1898) & (!g2022)) + ((g1890) & (g1939) & (!g1898) & (!g2022)) + ((g1890) & (g1939) & (g1898) & (g2022)));
	assign g3997 = (((!g830) & (!g1976) & (!g6950) & (key[78])) + ((!g830) & (!g1976) & (g6950) & (key[78])) + ((!g830) & (g1976) & (!g6950) & (key[78])) + ((!g830) & (g1976) & (g6950) & (key[78])) + ((g830) & (!g1976) & (g6950) & (!key[78])) + ((g830) & (!g1976) & (g6950) & (key[78])) + ((g830) & (g1976) & (!g6950) & (!key[78])) + ((g830) & (g1976) & (!g6950) & (key[78])));
	assign g3998 = (((!g3408) & (!g3038) & (g3044)) + ((!g3408) & (g3038) & (!g3044)) + ((!g3408) & (g3038) & (g3044)) + ((g3408) & (g3038) & (g3044)));
	assign g3999 = (((!g1610) & (!g3425) & (g3047)) + ((g1610) & (!g3425) & (!g3047)) + ((g1610) & (!g3425) & (g3047)) + ((g1610) & (g3425) & (g3047)));
	assign g8278 = (((!g5560) & (g5570) & (!g4000)) + ((!g5560) & (g5570) & (g4000)) + ((g5560) & (!g5570) & (g4000)) + ((g5560) & (g5570) & (g4000)));
	assign g4001 = (((!g830) & (!g1977) & (!g6937) & (g4000)) + ((!g830) & (!g1977) & (g6937) & (g4000)) + ((!g830) & (g1977) & (!g6937) & (g4000)) + ((!g830) & (g1977) & (g6937) & (g4000)) + ((g830) & (!g1977) & (g6937) & (!g4000)) + ((g830) & (!g1977) & (g6937) & (g4000)) + ((g830) & (g1977) & (!g6937) & (!g4000)) + ((g830) & (g1977) & (!g6937) & (g4000)));
	assign g4002 = (((!g3136) & (g3142)) + ((g3136) & (!g3142)));
	assign g4003 = (((!g3481) & (!g3061) & (!g3067) & (g3082) & (g3097) & (g4002)) + ((!g3481) & (!g3061) & (g3067) & (!g3082) & (g3097) & (g4002)) + ((!g3481) & (!g3061) & (g3067) & (g3082) & (!g3097) & (g4002)) + ((!g3481) & (!g3061) & (g3067) & (g3082) & (g3097) & (g4002)) + ((!g3481) & (g3061) & (!g3067) & (!g3082) & (g3097) & (g4002)) + ((!g3481) & (g3061) & (!g3067) & (g3082) & (!g3097) & (g4002)) + ((!g3481) & (g3061) & (!g3067) & (g3082) & (g3097) & (g4002)) + ((!g3481) & (g3061) & (g3067) & (!g3082) & (g3097) & (g4002)) + ((!g3481) & (g3061) & (g3067) & (g3082) & (!g3097) & (g4002)) + ((!g3481) & (g3061) & (g3067) & (g3082) & (g3097) & (g4002)) + ((g3481) & (!g3061) & (!g3067) & (g3082) & (g3097) & (g4002)) + ((g3481) & (!g3061) & (g3067) & (g3082) & (g3097) & (g4002)) + ((g3481) & (g3061) & (!g3067) & (g3082) & (g3097) & (g4002)) + ((g3481) & (g3061) & (g3067) & (!g3082) & (g3097) & (g4002)) + ((g3481) & (g3061) & (g3067) & (g3082) & (!g3097) & (g4002)) + ((g3481) & (g3061) & (g3067) & (g3082) & (g3097) & (g4002)));
	assign g4004 = (((g3136) & (g3142)));
	assign g4005 = (((!g3172) & (!g4003) & (!g4004) & (g3157)) + ((!g3172) & (!g4003) & (g4004) & (!g3157)) + ((!g3172) & (g4003) & (!g4004) & (!g3157)) + ((!g3172) & (g4003) & (g4004) & (!g3157)) + ((g3172) & (!g4003) & (!g4004) & (!g3157)) + ((g3172) & (!g4003) & (g4004) & (g3157)) + ((g3172) & (g4003) & (!g4004) & (g3157)) + ((g3172) & (g4003) & (g4004) & (g3157)));
	assign g4006 = (((!g2212) & (!g2262) & (!g2854) & (g2881) & (!g3496)) + ((!g2212) & (!g2262) & (!g2854) & (g2881) & (g3496)) + ((!g2212) & (!g2262) & (g2854) & (!g2881) & (g3496)) + ((!g2212) & (!g2262) & (g2854) & (g2881) & (!g3496)) + ((!g2212) & (g2262) & (!g2854) & (!g2881) & (!g3496)) + ((!g2212) & (g2262) & (!g2854) & (!g2881) & (g3496)) + ((!g2212) & (g2262) & (g2854) & (!g2881) & (!g3496)) + ((!g2212) & (g2262) & (g2854) & (g2881) & (g3496)) + ((g2212) & (!g2262) & (!g2854) & (!g2881) & (g3496)) + ((g2212) & (!g2262) & (!g2854) & (g2881) & (!g3496)) + ((g2212) & (!g2262) & (g2854) & (!g2881) & (!g3496)) + ((g2212) & (!g2262) & (g2854) & (!g2881) & (g3496)) + ((g2212) & (g2262) & (!g2854) & (!g2881) & (!g3496)) + ((g2212) & (g2262) & (!g2854) & (g2881) & (g3496)) + ((g2212) & (g2262) & (g2854) & (g2881) & (!g3496)) + ((g2212) & (g2262) & (g2854) & (g2881) & (g3496)));
	assign g4007 = (((!g830) & (!g1914) & (!g1978) & (!g4005) & (!g4006) & (key[161])) + ((!g830) & (!g1914) & (!g1978) & (!g4005) & (g4006) & (key[161])) + ((!g830) & (!g1914) & (!g1978) & (g4005) & (!g4006) & (key[161])) + ((!g830) & (!g1914) & (!g1978) & (g4005) & (g4006) & (key[161])) + ((!g830) & (!g1914) & (g1978) & (!g4005) & (!g4006) & (key[161])) + ((!g830) & (!g1914) & (g1978) & (!g4005) & (g4006) & (key[161])) + ((!g830) & (!g1914) & (g1978) & (g4005) & (!g4006) & (key[161])) + ((!g830) & (!g1914) & (g1978) & (g4005) & (g4006) & (key[161])) + ((!g830) & (g1914) & (!g1978) & (!g4005) & (!g4006) & (key[161])) + ((!g830) & (g1914) & (!g1978) & (!g4005) & (g4006) & (key[161])) + ((!g830) & (g1914) & (!g1978) & (g4005) & (!g4006) & (key[161])) + ((!g830) & (g1914) & (!g1978) & (g4005) & (g4006) & (key[161])) + ((!g830) & (g1914) & (g1978) & (!g4005) & (!g4006) & (key[161])) + ((!g830) & (g1914) & (g1978) & (!g4005) & (g4006) & (key[161])) + ((!g830) & (g1914) & (g1978) & (g4005) & (!g4006) & (key[161])) + ((!g830) & (g1914) & (g1978) & (g4005) & (g4006) & (key[161])) + ((g830) & (!g1914) & (!g1978) & (!g4005) & (g4006) & (!key[161])) + ((g830) & (!g1914) & (!g1978) & (!g4005) & (g4006) & (key[161])) + ((g830) & (!g1914) & (!g1978) & (g4005) & (g4006) & (!key[161])) + ((g830) & (!g1914) & (!g1978) & (g4005) & (g4006) & (key[161])) + ((g830) & (!g1914) & (g1978) & (!g4005) & (!g4006) & (!key[161])) + ((g830) & (!g1914) & (g1978) & (!g4005) & (!g4006) & (key[161])) + ((g830) & (!g1914) & (g1978) & (g4005) & (!g4006) & (!key[161])) + ((g830) & (!g1914) & (g1978) & (g4005) & (!g4006) & (key[161])) + ((g830) & (g1914) & (!g1978) & (g4005) & (!g4006) & (!key[161])) + ((g830) & (g1914) & (!g1978) & (g4005) & (!g4006) & (key[161])) + ((g830) & (g1914) & (!g1978) & (g4005) & (g4006) & (!key[161])) + ((g830) & (g1914) & (!g1978) & (g4005) & (g4006) & (key[161])) + ((g830) & (g1914) & (g1978) & (!g4005) & (!g4006) & (!key[161])) + ((g830) & (g1914) & (g1978) & (!g4005) & (!g4006) & (key[161])) + ((g830) & (g1914) & (g1978) & (!g4005) & (g4006) & (!key[161])) + ((g830) & (g1914) & (g1978) & (!g4005) & (g4006) & (key[161])));
	assign g4008 = (((!g3078) & (!g3113) & (!g3093) & (g3119) & (!g3998)) + ((!g3078) & (!g3113) & (!g3093) & (g3119) & (g3998)) + ((!g3078) & (!g3113) & (g3093) & (!g3119) & (g3998)) + ((!g3078) & (!g3113) & (g3093) & (g3119) & (!g3998)) + ((!g3078) & (g3113) & (!g3093) & (!g3119) & (!g3998)) + ((!g3078) & (g3113) & (!g3093) & (!g3119) & (g3998)) + ((!g3078) & (g3113) & (g3093) & (!g3119) & (!g3998)) + ((!g3078) & (g3113) & (g3093) & (g3119) & (g3998)) + ((g3078) & (!g3113) & (!g3093) & (!g3119) & (g3998)) + ((g3078) & (!g3113) & (!g3093) & (g3119) & (!g3998)) + ((g3078) & (!g3113) & (g3093) & (!g3119) & (!g3998)) + ((g3078) & (!g3113) & (g3093) & (!g3119) & (g3998)) + ((g3078) & (g3113) & (!g3093) & (!g3119) & (!g3998)) + ((g3078) & (g3113) & (!g3093) & (g3119) & (g3998)) + ((g3078) & (g3113) & (g3093) & (g3119) & (!g3998)) + ((g3078) & (g3113) & (g3093) & (g3119) & (g3998)));
	assign g4009 = (((!g1644) & (!g1677) & (!g3074) & (g3122) & (!g3999)) + ((!g1644) & (!g1677) & (!g3074) & (g3122) & (g3999)) + ((!g1644) & (!g1677) & (g3074) & (!g3122) & (g3999)) + ((!g1644) & (!g1677) & (g3074) & (g3122) & (!g3999)) + ((!g1644) & (g1677) & (!g3074) & (!g3122) & (!g3999)) + ((!g1644) & (g1677) & (!g3074) & (!g3122) & (g3999)) + ((!g1644) & (g1677) & (g3074) & (!g3122) & (!g3999)) + ((!g1644) & (g1677) & (g3074) & (g3122) & (g3999)) + ((g1644) & (!g1677) & (!g3074) & (!g3122) & (g3999)) + ((g1644) & (!g1677) & (!g3074) & (g3122) & (!g3999)) + ((g1644) & (!g1677) & (g3074) & (!g3122) & (!g3999)) + ((g1644) & (!g1677) & (g3074) & (!g3122) & (g3999)) + ((g1644) & (g1677) & (!g3074) & (!g3122) & (!g3999)) + ((g1644) & (g1677) & (!g3074) & (g3122) & (g3999)) + ((g1644) & (g1677) & (g3074) & (g3122) & (!g3999)) + ((g1644) & (g1677) & (g3074) & (g3122) & (g3999)));
	assign g8279 = (((!g5560) & (g5571) & (!g4010)) + ((!g5560) & (g5571) & (g4010)) + ((g5560) & (!g5571) & (g4010)) + ((g5560) & (g5571) & (g4010)));
	assign g4011 = (((!g830) & (!g1914) & (!g1979) & (!g4008) & (!g4009) & (g4010)) + ((!g830) & (!g1914) & (!g1979) & (!g4008) & (g4009) & (g4010)) + ((!g830) & (!g1914) & (!g1979) & (g4008) & (!g4009) & (g4010)) + ((!g830) & (!g1914) & (!g1979) & (g4008) & (g4009) & (g4010)) + ((!g830) & (!g1914) & (g1979) & (!g4008) & (!g4009) & (g4010)) + ((!g830) & (!g1914) & (g1979) & (!g4008) & (g4009) & (g4010)) + ((!g830) & (!g1914) & (g1979) & (g4008) & (!g4009) & (g4010)) + ((!g830) & (!g1914) & (g1979) & (g4008) & (g4009) & (g4010)) + ((!g830) & (g1914) & (!g1979) & (!g4008) & (!g4009) & (g4010)) + ((!g830) & (g1914) & (!g1979) & (!g4008) & (g4009) & (g4010)) + ((!g830) & (g1914) & (!g1979) & (g4008) & (!g4009) & (g4010)) + ((!g830) & (g1914) & (!g1979) & (g4008) & (g4009) & (g4010)) + ((!g830) & (g1914) & (g1979) & (!g4008) & (!g4009) & (g4010)) + ((!g830) & (g1914) & (g1979) & (!g4008) & (g4009) & (g4010)) + ((!g830) & (g1914) & (g1979) & (g4008) & (!g4009) & (g4010)) + ((!g830) & (g1914) & (g1979) & (g4008) & (g4009) & (g4010)) + ((g830) & (!g1914) & (!g1979) & (!g4008) & (g4009) & (!g4010)) + ((g830) & (!g1914) & (!g1979) & (!g4008) & (g4009) & (g4010)) + ((g830) & (!g1914) & (!g1979) & (g4008) & (g4009) & (!g4010)) + ((g830) & (!g1914) & (!g1979) & (g4008) & (g4009) & (g4010)) + ((g830) & (!g1914) & (g1979) & (!g4008) & (!g4009) & (!g4010)) + ((g830) & (!g1914) & (g1979) & (!g4008) & (!g4009) & (g4010)) + ((g830) & (!g1914) & (g1979) & (g4008) & (!g4009) & (!g4010)) + ((g830) & (!g1914) & (g1979) & (g4008) & (!g4009) & (g4010)) + ((g830) & (g1914) & (!g1979) & (g4008) & (!g4009) & (!g4010)) + ((g830) & (g1914) & (!g1979) & (g4008) & (!g4009) & (g4010)) + ((g830) & (g1914) & (!g1979) & (g4008) & (g4009) & (!g4010)) + ((g830) & (g1914) & (!g1979) & (g4008) & (g4009) & (g4010)) + ((g830) & (g1914) & (g1979) & (!g4008) & (!g4009) & (!g4010)) + ((g830) & (g1914) & (g1979) & (!g4008) & (!g4009) & (g4010)) + ((g830) & (g1914) & (g1979) & (!g4008) & (g4009) & (!g4010)) + ((g830) & (g1914) & (g1979) & (!g4008) & (g4009) & (g4010)));
	assign g4012 = (((!g3172) & (!g4003) & (!g4004) & (!g3157)) + ((!g3172) & (!g4003) & (!g4004) & (g3157)) + ((!g3172) & (!g4003) & (g4004) & (!g3157)) + ((!g3172) & (g4003) & (!g4004) & (!g3157)) + ((!g3172) & (g4003) & (g4004) & (!g3157)) + ((g3172) & (!g4003) & (!g4004) & (!g3157)));
	assign g4013 = (((!g2262) & (g2881)) + ((g2262) & (!g2881)));
	assign g4014 = (((!g2180) & (!g2212) & (g2797) & (g2854) & (!g3495) & (g4013)) + ((!g2180) & (g2212) & (!g2797) & (g2854) & (!g3495) & (g4013)) + ((!g2180) & (g2212) & (!g2797) & (g2854) & (g3495) & (g4013)) + ((!g2180) & (g2212) & (g2797) & (!g2854) & (!g3495) & (g4013)) + ((!g2180) & (g2212) & (g2797) & (g2854) & (!g3495) & (g4013)) + ((!g2180) & (g2212) & (g2797) & (g2854) & (g3495) & (g4013)) + ((g2180) & (!g2212) & (!g2797) & (g2854) & (!g3495) & (g4013)) + ((g2180) & (!g2212) & (g2797) & (g2854) & (!g3495) & (g4013)) + ((g2180) & (!g2212) & (g2797) & (g2854) & (g3495) & (g4013)) + ((g2180) & (g2212) & (!g2797) & (!g2854) & (!g3495) & (g4013)) + ((g2180) & (g2212) & (!g2797) & (g2854) & (!g3495) & (g4013)) + ((g2180) & (g2212) & (!g2797) & (g2854) & (g3495) & (g4013)) + ((g2180) & (g2212) & (g2797) & (!g2854) & (!g3495) & (g4013)) + ((g2180) & (g2212) & (g2797) & (!g2854) & (g3495) & (g4013)) + ((g2180) & (g2212) & (g2797) & (g2854) & (!g3495) & (g4013)) + ((g2180) & (g2212) & (g2797) & (g2854) & (g3495) & (g4013)));
	assign g4015 = (((g2262) & (g2881)));
	assign g4016 = (((!g2298) & (!g2950) & (!g4014) & (g4015)) + ((!g2298) & (!g2950) & (g4014) & (!g4015)) + ((!g2298) & (!g2950) & (g4014) & (g4015)) + ((!g2298) & (g2950) & (!g4014) & (!g4015)) + ((g2298) & (!g2950) & (!g4014) & (!g4015)) + ((g2298) & (g2950) & (!g4014) & (g4015)) + ((g2298) & (g2950) & (g4014) & (!g4015)) + ((g2298) & (g2950) & (g4014) & (g4015)));
	assign g4017 = (((!g1914) & (!g4012) & (!g3207) & (!g3213) & (g4016)) + ((!g1914) & (!g4012) & (!g3207) & (g3213) & (g4016)) + ((!g1914) & (!g4012) & (g3207) & (!g3213) & (g4016)) + ((!g1914) & (!g4012) & (g3207) & (g3213) & (g4016)) + ((!g1914) & (g4012) & (!g3207) & (!g3213) & (g4016)) + ((!g1914) & (g4012) & (!g3207) & (g3213) & (g4016)) + ((!g1914) & (g4012) & (g3207) & (!g3213) & (g4016)) + ((!g1914) & (g4012) & (g3207) & (g3213) & (g4016)) + ((g1914) & (!g4012) & (!g3207) & (!g3213) & (!g4016)) + ((g1914) & (!g4012) & (!g3207) & (!g3213) & (g4016)) + ((g1914) & (!g4012) & (g3207) & (g3213) & (!g4016)) + ((g1914) & (!g4012) & (g3207) & (g3213) & (g4016)) + ((g1914) & (g4012) & (!g3207) & (g3213) & (!g4016)) + ((g1914) & (g4012) & (!g3207) & (g3213) & (g4016)) + ((g1914) & (g4012) & (g3207) & (!g3213) & (!g4016)) + ((g1914) & (g4012) & (g3207) & (!g3213) & (g4016)));
	assign g4018 = (((!g830) & (!g1980) & (!g4017) & (key[162])) + ((!g830) & (!g1980) & (g4017) & (key[162])) + ((!g830) & (g1980) & (!g4017) & (key[162])) + ((!g830) & (g1980) & (g4017) & (key[162])) + ((g830) & (!g1980) & (g4017) & (!key[162])) + ((g830) & (!g1980) & (g4017) & (key[162])) + ((g830) & (g1980) & (!g4017) & (!key[162])) + ((g830) & (g1980) & (!g4017) & (key[162])));
	assign g4019 = (((!g3113) & (g3119)) + ((g3113) & (!g3119)));
	assign g4020 = (((!g3408) & (!g3038) & (!g3044) & (g3078) & (g3093) & (g4019)) + ((!g3408) & (!g3038) & (g3044) & (!g3078) & (g3093) & (g4019)) + ((!g3408) & (!g3038) & (g3044) & (g3078) & (!g3093) & (g4019)) + ((!g3408) & (!g3038) & (g3044) & (g3078) & (g3093) & (g4019)) + ((!g3408) & (g3038) & (!g3044) & (!g3078) & (g3093) & (g4019)) + ((!g3408) & (g3038) & (!g3044) & (g3078) & (!g3093) & (g4019)) + ((!g3408) & (g3038) & (!g3044) & (g3078) & (g3093) & (g4019)) + ((!g3408) & (g3038) & (g3044) & (!g3078) & (g3093) & (g4019)) + ((!g3408) & (g3038) & (g3044) & (g3078) & (!g3093) & (g4019)) + ((!g3408) & (g3038) & (g3044) & (g3078) & (g3093) & (g4019)) + ((g3408) & (!g3038) & (!g3044) & (g3078) & (g3093) & (g4019)) + ((g3408) & (!g3038) & (g3044) & (g3078) & (g3093) & (g4019)) + ((g3408) & (g3038) & (!g3044) & (g3078) & (g3093) & (g4019)) + ((g3408) & (g3038) & (g3044) & (!g3078) & (g3093) & (g4019)) + ((g3408) & (g3038) & (g3044) & (g3078) & (!g3093) & (g4019)) + ((g3408) & (g3038) & (g3044) & (g3078) & (g3093) & (g4019)));
	assign g4021 = (((g3113) & (g3119)));
	assign g4022 = (((!g3168) & (!g3153) & (!g4020) & (g4021)) + ((!g3168) & (!g3153) & (g4020) & (!g4021)) + ((!g3168) & (!g3153) & (g4020) & (g4021)) + ((!g3168) & (g3153) & (!g4020) & (!g4021)) + ((g3168) & (!g3153) & (!g4020) & (!g4021)) + ((g3168) & (g3153) & (!g4020) & (g4021)) + ((g3168) & (g3153) & (g4020) & (!g4021)) + ((g3168) & (g3153) & (g4020) & (g4021)));
	assign g4023 = (((!g1677) & (g3122)) + ((g1677) & (!g3122)));
	assign g4024 = (((!g1610) & (!g1644) & (!g3425) & (g3047) & (g3074) & (g4023)) + ((!g1610) & (g1644) & (!g3425) & (!g3047) & (g3074) & (g4023)) + ((!g1610) & (g1644) & (!g3425) & (g3047) & (!g3074) & (g4023)) + ((!g1610) & (g1644) & (!g3425) & (g3047) & (g3074) & (g4023)) + ((!g1610) & (g1644) & (g3425) & (!g3047) & (g3074) & (g4023)) + ((!g1610) & (g1644) & (g3425) & (g3047) & (g3074) & (g4023)) + ((g1610) & (!g1644) & (!g3425) & (!g3047) & (g3074) & (g4023)) + ((g1610) & (!g1644) & (!g3425) & (g3047) & (g3074) & (g4023)) + ((g1610) & (!g1644) & (g3425) & (g3047) & (g3074) & (g4023)) + ((g1610) & (g1644) & (!g3425) & (!g3047) & (!g3074) & (g4023)) + ((g1610) & (g1644) & (!g3425) & (!g3047) & (g3074) & (g4023)) + ((g1610) & (g1644) & (!g3425) & (g3047) & (!g3074) & (g4023)) + ((g1610) & (g1644) & (!g3425) & (g3047) & (g3074) & (g4023)) + ((g1610) & (g1644) & (g3425) & (!g3047) & (g3074) & (g4023)) + ((g1610) & (g1644) & (g3425) & (g3047) & (!g3074) & (g4023)) + ((g1610) & (g1644) & (g3425) & (g3047) & (g3074) & (g4023)));
	assign g4025 = (((g1677) & (g3122)));
	assign g4026 = (((!g1711) & (!g3149) & (!g4024) & (g4025)) + ((!g1711) & (!g3149) & (g4024) & (!g4025)) + ((!g1711) & (!g3149) & (g4024) & (g4025)) + ((!g1711) & (g3149) & (!g4024) & (!g4025)) + ((g1711) & (!g3149) & (!g4024) & (!g4025)) + ((g1711) & (g3149) & (!g4024) & (g4025)) + ((g1711) & (g3149) & (g4024) & (!g4025)) + ((g1711) & (g3149) & (g4024) & (g4025)));
	assign g8280 = (((!g5560) & (g5572) & (!g4027)) + ((!g5560) & (g5572) & (g4027)) + ((g5560) & (!g5572) & (g4027)) + ((g5560) & (g5572) & (g4027)));
	assign g4028 = (((!g830) & (!g1914) & (!g1982) & (!g4022) & (!g4026) & (g4027)) + ((!g830) & (!g1914) & (!g1982) & (!g4022) & (g4026) & (g4027)) + ((!g830) & (!g1914) & (!g1982) & (g4022) & (!g4026) & (g4027)) + ((!g830) & (!g1914) & (!g1982) & (g4022) & (g4026) & (g4027)) + ((!g830) & (!g1914) & (g1982) & (!g4022) & (!g4026) & (g4027)) + ((!g830) & (!g1914) & (g1982) & (!g4022) & (g4026) & (g4027)) + ((!g830) & (!g1914) & (g1982) & (g4022) & (!g4026) & (g4027)) + ((!g830) & (!g1914) & (g1982) & (g4022) & (g4026) & (g4027)) + ((!g830) & (g1914) & (!g1982) & (!g4022) & (!g4026) & (g4027)) + ((!g830) & (g1914) & (!g1982) & (!g4022) & (g4026) & (g4027)) + ((!g830) & (g1914) & (!g1982) & (g4022) & (!g4026) & (g4027)) + ((!g830) & (g1914) & (!g1982) & (g4022) & (g4026) & (g4027)) + ((!g830) & (g1914) & (g1982) & (!g4022) & (!g4026) & (g4027)) + ((!g830) & (g1914) & (g1982) & (!g4022) & (g4026) & (g4027)) + ((!g830) & (g1914) & (g1982) & (g4022) & (!g4026) & (g4027)) + ((!g830) & (g1914) & (g1982) & (g4022) & (g4026) & (g4027)) + ((g830) & (!g1914) & (!g1982) & (!g4022) & (g4026) & (!g4027)) + ((g830) & (!g1914) & (!g1982) & (!g4022) & (g4026) & (g4027)) + ((g830) & (!g1914) & (!g1982) & (g4022) & (g4026) & (!g4027)) + ((g830) & (!g1914) & (!g1982) & (g4022) & (g4026) & (g4027)) + ((g830) & (!g1914) & (g1982) & (!g4022) & (!g4026) & (!g4027)) + ((g830) & (!g1914) & (g1982) & (!g4022) & (!g4026) & (g4027)) + ((g830) & (!g1914) & (g1982) & (g4022) & (!g4026) & (!g4027)) + ((g830) & (!g1914) & (g1982) & (g4022) & (!g4026) & (g4027)) + ((g830) & (g1914) & (!g1982) & (g4022) & (!g4026) & (!g4027)) + ((g830) & (g1914) & (!g1982) & (g4022) & (!g4026) & (g4027)) + ((g830) & (g1914) & (!g1982) & (g4022) & (g4026) & (!g4027)) + ((g830) & (g1914) & (!g1982) & (g4022) & (g4026) & (g4027)) + ((g830) & (g1914) & (g1982) & (!g4022) & (!g4026) & (!g4027)) + ((g830) & (g1914) & (g1982) & (!g4022) & (!g4026) & (g4027)) + ((g830) & (g1914) & (g1982) & (!g4022) & (g4026) & (!g4027)) + ((g830) & (g1914) & (g1982) & (!g4022) & (g4026) & (g4027)));
	assign g4029 = (((!g3172) & (!g4003) & (!g4004) & (!g3157) & (!g3207) & (!g3213)) + ((!g3172) & (!g4003) & (!g4004) & (!g3157) & (!g3207) & (g3213)) + ((!g3172) & (!g4003) & (!g4004) & (!g3157) & (g3207) & (!g3213)) + ((!g3172) & (!g4003) & (!g4004) & (g3157) & (!g3207) & (!g3213)) + ((!g3172) & (!g4003) & (!g4004) & (g3157) & (!g3207) & (g3213)) + ((!g3172) & (!g4003) & (!g4004) & (g3157) & (g3207) & (!g3213)) + ((!g3172) & (!g4003) & (g4004) & (!g3157) & (!g3207) & (!g3213)) + ((!g3172) & (!g4003) & (g4004) & (!g3157) & (!g3207) & (g3213)) + ((!g3172) & (!g4003) & (g4004) & (!g3157) & (g3207) & (!g3213)) + ((!g3172) & (!g4003) & (g4004) & (g3157) & (!g3207) & (!g3213)) + ((!g3172) & (g4003) & (!g4004) & (!g3157) & (!g3207) & (!g3213)) + ((!g3172) & (g4003) & (!g4004) & (!g3157) & (!g3207) & (g3213)) + ((!g3172) & (g4003) & (!g4004) & (!g3157) & (g3207) & (!g3213)) + ((!g3172) & (g4003) & (!g4004) & (g3157) & (!g3207) & (!g3213)) + ((!g3172) & (g4003) & (g4004) & (!g3157) & (!g3207) & (!g3213)) + ((!g3172) & (g4003) & (g4004) & (!g3157) & (!g3207) & (g3213)) + ((!g3172) & (g4003) & (g4004) & (!g3157) & (g3207) & (!g3213)) + ((!g3172) & (g4003) & (g4004) & (g3157) & (!g3207) & (!g3213)) + ((g3172) & (!g4003) & (!g4004) & (!g3157) & (!g3207) & (!g3213)) + ((g3172) & (!g4003) & (!g4004) & (!g3157) & (!g3207) & (g3213)) + ((g3172) & (!g4003) & (!g4004) & (!g3157) & (g3207) & (!g3213)) + ((g3172) & (!g4003) & (!g4004) & (g3157) & (!g3207) & (!g3213)) + ((g3172) & (!g4003) & (g4004) & (!g3157) & (!g3207) & (!g3213)) + ((g3172) & (!g4003) & (g4004) & (g3157) & (!g3207) & (!g3213)) + ((g3172) & (g4003) & (!g4004) & (!g3157) & (!g3207) & (!g3213)) + ((g3172) & (g4003) & (!g4004) & (g3157) & (!g3207) & (!g3213)) + ((g3172) & (g4003) & (g4004) & (!g3157) & (!g3207) & (!g3213)) + ((g3172) & (g4003) & (g4004) & (g3157) & (!g3207) & (!g3213)));
	assign g4030 = (((!g2298) & (!g2347) & (!g2950) & (g2999) & (!g4014) & (!g4015)) + ((!g2298) & (!g2347) & (!g2950) & (g2999) & (!g4014) & (g4015)) + ((!g2298) & (!g2347) & (!g2950) & (g2999) & (g4014) & (!g4015)) + ((!g2298) & (!g2347) & (!g2950) & (g2999) & (g4014) & (g4015)) + ((!g2298) & (!g2347) & (g2950) & (!g2999) & (!g4014) & (g4015)) + ((!g2298) & (!g2347) & (g2950) & (!g2999) & (g4014) & (!g4015)) + ((!g2298) & (!g2347) & (g2950) & (!g2999) & (g4014) & (g4015)) + ((!g2298) & (!g2347) & (g2950) & (g2999) & (!g4014) & (!g4015)) + ((!g2298) & (g2347) & (!g2950) & (!g2999) & (!g4014) & (!g4015)) + ((!g2298) & (g2347) & (!g2950) & (!g2999) & (!g4014) & (g4015)) + ((!g2298) & (g2347) & (!g2950) & (!g2999) & (g4014) & (!g4015)) + ((!g2298) & (g2347) & (!g2950) & (!g2999) & (g4014) & (g4015)) + ((!g2298) & (g2347) & (g2950) & (!g2999) & (!g4014) & (!g4015)) + ((!g2298) & (g2347) & (g2950) & (g2999) & (!g4014) & (g4015)) + ((!g2298) & (g2347) & (g2950) & (g2999) & (g4014) & (!g4015)) + ((!g2298) & (g2347) & (g2950) & (g2999) & (g4014) & (g4015)) + ((g2298) & (!g2347) & (!g2950) & (!g2999) & (!g4014) & (g4015)) + ((g2298) & (!g2347) & (!g2950) & (!g2999) & (g4014) & (!g4015)) + ((g2298) & (!g2347) & (!g2950) & (!g2999) & (g4014) & (g4015)) + ((g2298) & (!g2347) & (!g2950) & (g2999) & (!g4014) & (!g4015)) + ((g2298) & (!g2347) & (g2950) & (!g2999) & (!g4014) & (!g4015)) + ((g2298) & (!g2347) & (g2950) & (!g2999) & (!g4014) & (g4015)) + ((g2298) & (!g2347) & (g2950) & (!g2999) & (g4014) & (!g4015)) + ((g2298) & (!g2347) & (g2950) & (!g2999) & (g4014) & (g4015)) + ((g2298) & (g2347) & (!g2950) & (!g2999) & (!g4014) & (!g4015)) + ((g2298) & (g2347) & (!g2950) & (g2999) & (!g4014) & (g4015)) + ((g2298) & (g2347) & (!g2950) & (g2999) & (g4014) & (!g4015)) + ((g2298) & (g2347) & (!g2950) & (g2999) & (g4014) & (g4015)) + ((g2298) & (g2347) & (g2950) & (g2999) & (!g4014) & (!g4015)) + ((g2298) & (g2347) & (g2950) & (g2999) & (!g4014) & (g4015)) + ((g2298) & (g2347) & (g2950) & (g2999) & (g4014) & (!g4015)) + ((g2298) & (g2347) & (g2950) & (g2999) & (g4014) & (g4015)));
	assign g4031 = (((!g1914) & (!g3284) & (!g4029) & (!g3245) & (g4030)) + ((!g1914) & (!g3284) & (!g4029) & (g3245) & (g4030)) + ((!g1914) & (!g3284) & (g4029) & (!g3245) & (g4030)) + ((!g1914) & (!g3284) & (g4029) & (g3245) & (g4030)) + ((!g1914) & (g3284) & (!g4029) & (!g3245) & (g4030)) + ((!g1914) & (g3284) & (!g4029) & (g3245) & (g4030)) + ((!g1914) & (g3284) & (g4029) & (!g3245) & (g4030)) + ((!g1914) & (g3284) & (g4029) & (g3245) & (g4030)) + ((g1914) & (!g3284) & (!g4029) & (!g3245) & (!g4030)) + ((g1914) & (!g3284) & (!g4029) & (!g3245) & (g4030)) + ((g1914) & (!g3284) & (g4029) & (g3245) & (!g4030)) + ((g1914) & (!g3284) & (g4029) & (g3245) & (g4030)) + ((g1914) & (g3284) & (!g4029) & (g3245) & (!g4030)) + ((g1914) & (g3284) & (!g4029) & (g3245) & (g4030)) + ((g1914) & (g3284) & (g4029) & (!g3245) & (!g4030)) + ((g1914) & (g3284) & (g4029) & (!g3245) & (g4030)));
	assign g4032 = (((!g830) & (!g1983) & (!g4031) & (key[163])) + ((!g830) & (!g1983) & (g4031) & (key[163])) + ((!g830) & (g1983) & (!g4031) & (key[163])) + ((!g830) & (g1983) & (g4031) & (key[163])) + ((g830) & (!g1983) & (g4031) & (!key[163])) + ((g830) & (!g1983) & (g4031) & (key[163])) + ((g830) & (g1983) & (!g4031) & (!key[163])) + ((g830) & (g1983) & (!g4031) & (key[163])));
	assign g4033 = (((!g3168) & (!g3153) & (!g4020) & (!g4021)) + ((!g3168) & (!g3153) & (!g4020) & (g4021)) + ((!g3168) & (!g3153) & (g4020) & (!g4021)) + ((!g3168) & (!g3153) & (g4020) & (g4021)) + ((!g3168) & (g3153) & (!g4020) & (!g4021)) + ((g3168) & (!g3153) & (!g4020) & (!g4021)));
	assign g4034 = (((!g1711) & (!g1744) & (!g3149) & (g3193) & (!g4024) & (!g4025)) + ((!g1711) & (!g1744) & (!g3149) & (g3193) & (!g4024) & (g4025)) + ((!g1711) & (!g1744) & (!g3149) & (g3193) & (g4024) & (!g4025)) + ((!g1711) & (!g1744) & (!g3149) & (g3193) & (g4024) & (g4025)) + ((!g1711) & (!g1744) & (g3149) & (!g3193) & (!g4024) & (g4025)) + ((!g1711) & (!g1744) & (g3149) & (!g3193) & (g4024) & (!g4025)) + ((!g1711) & (!g1744) & (g3149) & (!g3193) & (g4024) & (g4025)) + ((!g1711) & (!g1744) & (g3149) & (g3193) & (!g4024) & (!g4025)) + ((!g1711) & (g1744) & (!g3149) & (!g3193) & (!g4024) & (!g4025)) + ((!g1711) & (g1744) & (!g3149) & (!g3193) & (!g4024) & (g4025)) + ((!g1711) & (g1744) & (!g3149) & (!g3193) & (g4024) & (!g4025)) + ((!g1711) & (g1744) & (!g3149) & (!g3193) & (g4024) & (g4025)) + ((!g1711) & (g1744) & (g3149) & (!g3193) & (!g4024) & (!g4025)) + ((!g1711) & (g1744) & (g3149) & (g3193) & (!g4024) & (g4025)) + ((!g1711) & (g1744) & (g3149) & (g3193) & (g4024) & (!g4025)) + ((!g1711) & (g1744) & (g3149) & (g3193) & (g4024) & (g4025)) + ((g1711) & (!g1744) & (!g3149) & (!g3193) & (!g4024) & (g4025)) + ((g1711) & (!g1744) & (!g3149) & (!g3193) & (g4024) & (!g4025)) + ((g1711) & (!g1744) & (!g3149) & (!g3193) & (g4024) & (g4025)) + ((g1711) & (!g1744) & (!g3149) & (g3193) & (!g4024) & (!g4025)) + ((g1711) & (!g1744) & (g3149) & (!g3193) & (!g4024) & (!g4025)) + ((g1711) & (!g1744) & (g3149) & (!g3193) & (!g4024) & (g4025)) + ((g1711) & (!g1744) & (g3149) & (!g3193) & (g4024) & (!g4025)) + ((g1711) & (!g1744) & (g3149) & (!g3193) & (g4024) & (g4025)) + ((g1711) & (g1744) & (!g3149) & (!g3193) & (!g4024) & (!g4025)) + ((g1711) & (g1744) & (!g3149) & (g3193) & (!g4024) & (g4025)) + ((g1711) & (g1744) & (!g3149) & (g3193) & (g4024) & (!g4025)) + ((g1711) & (g1744) & (!g3149) & (g3193) & (g4024) & (g4025)) + ((g1711) & (g1744) & (g3149) & (g3193) & (!g4024) & (!g4025)) + ((g1711) & (g1744) & (g3149) & (g3193) & (!g4024) & (g4025)) + ((g1711) & (g1744) & (g3149) & (g3193) & (g4024) & (!g4025)) + ((g1711) & (g1744) & (g3149) & (g3193) & (g4024) & (g4025)));
	assign g4035 = (((!g1914) & (!g3184) & (!g3190) & (!g4033) & (g4034)) + ((!g1914) & (!g3184) & (!g3190) & (g4033) & (g4034)) + ((!g1914) & (!g3184) & (g3190) & (!g4033) & (g4034)) + ((!g1914) & (!g3184) & (g3190) & (g4033) & (g4034)) + ((!g1914) & (g3184) & (!g3190) & (!g4033) & (g4034)) + ((!g1914) & (g3184) & (!g3190) & (g4033) & (g4034)) + ((!g1914) & (g3184) & (g3190) & (!g4033) & (g4034)) + ((!g1914) & (g3184) & (g3190) & (g4033) & (g4034)) + ((g1914) & (!g3184) & (!g3190) & (!g4033) & (!g4034)) + ((g1914) & (!g3184) & (!g3190) & (!g4033) & (g4034)) + ((g1914) & (!g3184) & (g3190) & (g4033) & (!g4034)) + ((g1914) & (!g3184) & (g3190) & (g4033) & (g4034)) + ((g1914) & (g3184) & (!g3190) & (g4033) & (!g4034)) + ((g1914) & (g3184) & (!g3190) & (g4033) & (g4034)) + ((g1914) & (g3184) & (g3190) & (!g4033) & (!g4034)) + ((g1914) & (g3184) & (g3190) & (!g4033) & (g4034)));
	assign g8281 = (((!g5560) & (g5573) & (!g4036)) + ((!g5560) & (g5573) & (g4036)) + ((g5560) & (!g5573) & (g4036)) + ((g5560) & (g5573) & (g4036)));
	assign g4037 = (((!g830) & (!g1984) & (!g4035) & (g4036)) + ((!g830) & (!g1984) & (g4035) & (g4036)) + ((!g830) & (g1984) & (!g4035) & (g4036)) + ((!g830) & (g1984) & (g4035) & (g4036)) + ((g830) & (!g1984) & (g4035) & (!g4036)) + ((g830) & (!g1984) & (g4035) & (g4036)) + ((g830) & (g1984) & (!g4035) & (!g4036)) + ((g830) & (g1984) & (!g4035) & (g4036)));
	assign g4038 = (((!g3284) & (!g4029) & (!g3245) & (!g3310) & (g3314)) + ((!g3284) & (!g4029) & (!g3245) & (g3310) & (!g3314)) + ((!g3284) & (!g4029) & (g3245) & (!g3310) & (!g3314)) + ((!g3284) & (!g4029) & (g3245) & (g3310) & (g3314)) + ((!g3284) & (g4029) & (!g3245) & (!g3310) & (g3314)) + ((!g3284) & (g4029) & (!g3245) & (g3310) & (!g3314)) + ((!g3284) & (g4029) & (g3245) & (!g3310) & (g3314)) + ((!g3284) & (g4029) & (g3245) & (g3310) & (!g3314)) + ((g3284) & (!g4029) & (!g3245) & (!g3310) & (!g3314)) + ((g3284) & (!g4029) & (!g3245) & (g3310) & (g3314)) + ((g3284) & (!g4029) & (g3245) & (!g3310) & (!g3314)) + ((g3284) & (!g4029) & (g3245) & (g3310) & (g3314)) + ((g3284) & (g4029) & (!g3245) & (!g3310) & (g3314)) + ((g3284) & (g4029) & (!g3245) & (g3310) & (!g3314)) + ((g3284) & (g4029) & (g3245) & (!g3310) & (!g3314)) + ((g3284) & (g4029) & (g3245) & (g3310) & (g3314)));
	assign g4039 = (((!g2298) & (!g2347) & (!g2950) & (!g2999) & (!g4014) & (!g4015)) + ((!g2298) & (!g2347) & (!g2950) & (!g2999) & (!g4014) & (g4015)) + ((!g2298) & (!g2347) & (!g2950) & (!g2999) & (g4014) & (!g4015)) + ((!g2298) & (!g2347) & (!g2950) & (!g2999) & (g4014) & (g4015)) + ((!g2298) & (!g2347) & (!g2950) & (g2999) & (!g4014) & (!g4015)) + ((!g2298) & (!g2347) & (!g2950) & (g2999) & (!g4014) & (g4015)) + ((!g2298) & (!g2347) & (!g2950) & (g2999) & (g4014) & (!g4015)) + ((!g2298) & (!g2347) & (!g2950) & (g2999) & (g4014) & (g4015)) + ((!g2298) & (!g2347) & (g2950) & (!g2999) & (!g4014) & (!g4015)) + ((!g2298) & (!g2347) & (g2950) & (!g2999) & (!g4014) & (g4015)) + ((!g2298) & (!g2347) & (g2950) & (!g2999) & (g4014) & (!g4015)) + ((!g2298) & (!g2347) & (g2950) & (!g2999) & (g4014) & (g4015)) + ((!g2298) & (!g2347) & (g2950) & (g2999) & (!g4014) & (!g4015)) + ((!g2298) & (g2347) & (!g2950) & (!g2999) & (!g4014) & (!g4015)) + ((!g2298) & (g2347) & (!g2950) & (!g2999) & (!g4014) & (g4015)) + ((!g2298) & (g2347) & (!g2950) & (!g2999) & (g4014) & (!g4015)) + ((!g2298) & (g2347) & (!g2950) & (!g2999) & (g4014) & (g4015)) + ((!g2298) & (g2347) & (g2950) & (!g2999) & (!g4014) & (!g4015)) + ((g2298) & (!g2347) & (!g2950) & (!g2999) & (!g4014) & (!g4015)) + ((g2298) & (!g2347) & (!g2950) & (!g2999) & (!g4014) & (g4015)) + ((g2298) & (!g2347) & (!g2950) & (!g2999) & (g4014) & (!g4015)) + ((g2298) & (!g2347) & (!g2950) & (!g2999) & (g4014) & (g4015)) + ((g2298) & (!g2347) & (!g2950) & (g2999) & (!g4014) & (!g4015)) + ((g2298) & (!g2347) & (g2950) & (!g2999) & (!g4014) & (!g4015)) + ((g2298) & (!g2347) & (g2950) & (!g2999) & (!g4014) & (g4015)) + ((g2298) & (!g2347) & (g2950) & (!g2999) & (g4014) & (!g4015)) + ((g2298) & (!g2347) & (g2950) & (!g2999) & (g4014) & (g4015)) + ((g2298) & (g2347) & (!g2950) & (!g2999) & (!g4014) & (!g4015)));
	assign g4040 = (((!g2378) & (!g3047) & (!g4039)) + ((!g2378) & (g3047) & (g4039)) + ((g2378) & (!g3047) & (g4039)) + ((g2378) & (g3047) & (!g4039)));
	assign g4041 = (((!g830) & (!g1914) & (!g1985) & (!g4038) & (!g4040) & (key[164])) + ((!g830) & (!g1914) & (!g1985) & (!g4038) & (g4040) & (key[164])) + ((!g830) & (!g1914) & (!g1985) & (g4038) & (!g4040) & (key[164])) + ((!g830) & (!g1914) & (!g1985) & (g4038) & (g4040) & (key[164])) + ((!g830) & (!g1914) & (g1985) & (!g4038) & (!g4040) & (key[164])) + ((!g830) & (!g1914) & (g1985) & (!g4038) & (g4040) & (key[164])) + ((!g830) & (!g1914) & (g1985) & (g4038) & (!g4040) & (key[164])) + ((!g830) & (!g1914) & (g1985) & (g4038) & (g4040) & (key[164])) + ((!g830) & (g1914) & (!g1985) & (!g4038) & (!g4040) & (key[164])) + ((!g830) & (g1914) & (!g1985) & (!g4038) & (g4040) & (key[164])) + ((!g830) & (g1914) & (!g1985) & (g4038) & (!g4040) & (key[164])) + ((!g830) & (g1914) & (!g1985) & (g4038) & (g4040) & (key[164])) + ((!g830) & (g1914) & (g1985) & (!g4038) & (!g4040) & (key[164])) + ((!g830) & (g1914) & (g1985) & (!g4038) & (g4040) & (key[164])) + ((!g830) & (g1914) & (g1985) & (g4038) & (!g4040) & (key[164])) + ((!g830) & (g1914) & (g1985) & (g4038) & (g4040) & (key[164])) + ((g830) & (!g1914) & (!g1985) & (!g4038) & (g4040) & (!key[164])) + ((g830) & (!g1914) & (!g1985) & (!g4038) & (g4040) & (key[164])) + ((g830) & (!g1914) & (!g1985) & (g4038) & (g4040) & (!key[164])) + ((g830) & (!g1914) & (!g1985) & (g4038) & (g4040) & (key[164])) + ((g830) & (!g1914) & (g1985) & (!g4038) & (!g4040) & (!key[164])) + ((g830) & (!g1914) & (g1985) & (!g4038) & (!g4040) & (key[164])) + ((g830) & (!g1914) & (g1985) & (g4038) & (!g4040) & (!key[164])) + ((g830) & (!g1914) & (g1985) & (g4038) & (!g4040) & (key[164])) + ((g830) & (g1914) & (!g1985) & (g4038) & (!g4040) & (!key[164])) + ((g830) & (g1914) & (!g1985) & (g4038) & (!g4040) & (key[164])) + ((g830) & (g1914) & (!g1985) & (g4038) & (g4040) & (!key[164])) + ((g830) & (g1914) & (!g1985) & (g4038) & (g4040) & (key[164])) + ((g830) & (g1914) & (g1985) & (!g4038) & (!g4040) & (!key[164])) + ((g830) & (g1914) & (g1985) & (!g4038) & (!g4040) & (key[164])) + ((g830) & (g1914) & (g1985) & (!g4038) & (g4040) & (!key[164])) + ((g830) & (g1914) & (g1985) & (!g4038) & (g4040) & (key[164])));
	assign g4042 = (((!g3168) & (!g3153) & (!g3184) & (!g3190) & (!g4020) & (!g4021)) + ((!g3168) & (!g3153) & (!g3184) & (!g3190) & (!g4020) & (g4021)) + ((!g3168) & (!g3153) & (!g3184) & (!g3190) & (g4020) & (!g4021)) + ((!g3168) & (!g3153) & (!g3184) & (!g3190) & (g4020) & (g4021)) + ((!g3168) & (!g3153) & (!g3184) & (g3190) & (!g4020) & (!g4021)) + ((!g3168) & (!g3153) & (!g3184) & (g3190) & (!g4020) & (g4021)) + ((!g3168) & (!g3153) & (!g3184) & (g3190) & (g4020) & (!g4021)) + ((!g3168) & (!g3153) & (!g3184) & (g3190) & (g4020) & (g4021)) + ((!g3168) & (!g3153) & (g3184) & (!g3190) & (!g4020) & (!g4021)) + ((!g3168) & (!g3153) & (g3184) & (!g3190) & (!g4020) & (g4021)) + ((!g3168) & (!g3153) & (g3184) & (!g3190) & (g4020) & (!g4021)) + ((!g3168) & (!g3153) & (g3184) & (!g3190) & (g4020) & (g4021)) + ((!g3168) & (g3153) & (!g3184) & (!g3190) & (!g4020) & (!g4021)) + ((!g3168) & (g3153) & (!g3184) & (!g3190) & (!g4020) & (g4021)) + ((!g3168) & (g3153) & (!g3184) & (!g3190) & (g4020) & (!g4021)) + ((!g3168) & (g3153) & (!g3184) & (!g3190) & (g4020) & (g4021)) + ((!g3168) & (g3153) & (!g3184) & (g3190) & (!g4020) & (!g4021)) + ((!g3168) & (g3153) & (g3184) & (!g3190) & (!g4020) & (!g4021)) + ((g3168) & (!g3153) & (!g3184) & (!g3190) & (!g4020) & (!g4021)) + ((g3168) & (!g3153) & (!g3184) & (!g3190) & (!g4020) & (g4021)) + ((g3168) & (!g3153) & (!g3184) & (!g3190) & (g4020) & (!g4021)) + ((g3168) & (!g3153) & (!g3184) & (!g3190) & (g4020) & (g4021)) + ((g3168) & (!g3153) & (!g3184) & (g3190) & (!g4020) & (!g4021)) + ((g3168) & (!g3153) & (g3184) & (!g3190) & (!g4020) & (!g4021)) + ((g3168) & (g3153) & (!g3184) & (!g3190) & (!g4020) & (!g4021)) + ((g3168) & (g3153) & (!g3184) & (!g3190) & (!g4020) & (g4021)) + ((g3168) & (g3153) & (!g3184) & (!g3190) & (g4020) & (!g4021)) + ((g3168) & (g3153) & (!g3184) & (!g3190) & (g4020) & (g4021)));
	assign g4043 = (((g1914) & (!g3274) & (!g3235) & (!g4042)) + ((g1914) & (!g3274) & (g3235) & (g4042)) + ((g1914) & (g3274) & (!g3235) & (g4042)) + ((g1914) & (g3274) & (g3235) & (!g4042)));
	assign g4044 = (((!g1711) & (!g1744) & (!g3149) & (!g3193) & (!g4024) & (!g4025)) + ((!g1711) & (!g1744) & (!g3149) & (!g3193) & (!g4024) & (g4025)) + ((!g1711) & (!g1744) & (!g3149) & (!g3193) & (g4024) & (!g4025)) + ((!g1711) & (!g1744) & (!g3149) & (!g3193) & (g4024) & (g4025)) + ((!g1711) & (!g1744) & (!g3149) & (g3193) & (!g4024) & (!g4025)) + ((!g1711) & (!g1744) & (!g3149) & (g3193) & (!g4024) & (g4025)) + ((!g1711) & (!g1744) & (!g3149) & (g3193) & (g4024) & (!g4025)) + ((!g1711) & (!g1744) & (!g3149) & (g3193) & (g4024) & (g4025)) + ((!g1711) & (!g1744) & (g3149) & (!g3193) & (!g4024) & (!g4025)) + ((!g1711) & (!g1744) & (g3149) & (!g3193) & (!g4024) & (g4025)) + ((!g1711) & (!g1744) & (g3149) & (!g3193) & (g4024) & (!g4025)) + ((!g1711) & (!g1744) & (g3149) & (!g3193) & (g4024) & (g4025)) + ((!g1711) & (!g1744) & (g3149) & (g3193) & (!g4024) & (!g4025)) + ((!g1711) & (g1744) & (!g3149) & (!g3193) & (!g4024) & (!g4025)) + ((!g1711) & (g1744) & (!g3149) & (!g3193) & (!g4024) & (g4025)) + ((!g1711) & (g1744) & (!g3149) & (!g3193) & (g4024) & (!g4025)) + ((!g1711) & (g1744) & (!g3149) & (!g3193) & (g4024) & (g4025)) + ((!g1711) & (g1744) & (g3149) & (!g3193) & (!g4024) & (!g4025)) + ((g1711) & (!g1744) & (!g3149) & (!g3193) & (!g4024) & (!g4025)) + ((g1711) & (!g1744) & (!g3149) & (!g3193) & (!g4024) & (g4025)) + ((g1711) & (!g1744) & (!g3149) & (!g3193) & (g4024) & (!g4025)) + ((g1711) & (!g1744) & (!g3149) & (!g3193) & (g4024) & (g4025)) + ((g1711) & (!g1744) & (!g3149) & (g3193) & (!g4024) & (!g4025)) + ((g1711) & (!g1744) & (g3149) & (!g3193) & (!g4024) & (!g4025)) + ((g1711) & (!g1744) & (g3149) & (!g3193) & (!g4024) & (g4025)) + ((g1711) & (!g1744) & (g3149) & (!g3193) & (g4024) & (!g4025)) + ((g1711) & (!g1744) & (g3149) & (!g3193) & (g4024) & (g4025)) + ((g1711) & (g1744) & (!g3149) & (!g3193) & (!g4024) & (!g4025)));
	assign g4045 = (((!g1914) & (!g1778) & (!g3222) & (!g4044)) + ((!g1914) & (!g1778) & (g3222) & (g4044)) + ((!g1914) & (g1778) & (!g3222) & (g4044)) + ((!g1914) & (g1778) & (g3222) & (!g4044)));
	assign g8282 = (((!g5560) & (g5574) & (!g4046)) + ((!g5560) & (g5574) & (g4046)) + ((g5560) & (!g5574) & (g4046)) + ((g5560) & (g5574) & (g4046)));
	assign g4047 = (((!g830) & (!g1986) & (!g4043) & (!g4045) & (g4046)) + ((!g830) & (!g1986) & (!g4043) & (g4045) & (g4046)) + ((!g830) & (!g1986) & (g4043) & (!g4045) & (g4046)) + ((!g830) & (!g1986) & (g4043) & (g4045) & (g4046)) + ((!g830) & (g1986) & (!g4043) & (!g4045) & (g4046)) + ((!g830) & (g1986) & (!g4043) & (g4045) & (g4046)) + ((!g830) & (g1986) & (g4043) & (!g4045) & (g4046)) + ((!g830) & (g1986) & (g4043) & (g4045) & (g4046)) + ((g830) & (!g1986) & (!g4043) & (g4045) & (!g4046)) + ((g830) & (!g1986) & (!g4043) & (g4045) & (g4046)) + ((g830) & (!g1986) & (g4043) & (!g4045) & (!g4046)) + ((g830) & (!g1986) & (g4043) & (!g4045) & (g4046)) + ((g830) & (!g1986) & (g4043) & (g4045) & (!g4046)) + ((g830) & (!g1986) & (g4043) & (g4045) & (g4046)) + ((g830) & (g1986) & (!g4043) & (!g4045) & (!g4046)) + ((g830) & (g1986) & (!g4043) & (!g4045) & (g4046)));
	assign g4048 = (((!g3172) & (!g4003) & (!g4004) & (!g3157) & (!g5776) & (!g5777)) + ((!g3172) & (!g4003) & (!g4004) & (g3157) & (!g5776) & (!g5777)) + ((!g3172) & (!g4003) & (g4004) & (!g3157) & (!g5776) & (!g5777)) + ((!g3172) & (!g4003) & (g4004) & (g3157) & (!g5776) & (!g5777)) + ((!g3172) & (!g4003) & (g4004) & (g3157) & (!g5776) & (g5777)) + ((!g3172) & (g4003) & (!g4004) & (!g3157) & (!g5776) & (!g5777)) + ((!g3172) & (g4003) & (!g4004) & (g3157) & (!g5776) & (!g5777)) + ((!g3172) & (g4003) & (!g4004) & (g3157) & (!g5776) & (g5777)) + ((!g3172) & (g4003) & (g4004) & (!g3157) & (!g5776) & (!g5777)) + ((!g3172) & (g4003) & (g4004) & (g3157) & (!g5776) & (!g5777)) + ((!g3172) & (g4003) & (g4004) & (g3157) & (!g5776) & (g5777)) + ((g3172) & (!g4003) & (!g4004) & (!g3157) & (!g5776) & (!g5777)) + ((g3172) & (!g4003) & (!g4004) & (g3157) & (!g5776) & (!g5777)) + ((g3172) & (!g4003) & (!g4004) & (g3157) & (!g5776) & (g5777)) + ((g3172) & (!g4003) & (g4004) & (!g3157) & (!g5776) & (!g5777)) + ((g3172) & (!g4003) & (g4004) & (!g3157) & (!g5776) & (g5777)) + ((g3172) & (!g4003) & (g4004) & (g3157) & (!g5776) & (!g5777)) + ((g3172) & (!g4003) & (g4004) & (g3157) & (!g5776) & (g5777)) + ((g3172) & (g4003) & (!g4004) & (!g3157) & (!g5776) & (!g5777)) + ((g3172) & (g4003) & (!g4004) & (!g3157) & (!g5776) & (g5777)) + ((g3172) & (g4003) & (!g4004) & (g3157) & (!g5776) & (!g5777)) + ((g3172) & (g4003) & (!g4004) & (g3157) & (!g5776) & (g5777)) + ((g3172) & (g4003) & (g4004) & (!g3157) & (!g5776) & (!g5777)) + ((g3172) & (g4003) & (g4004) & (!g3157) & (!g5776) & (g5777)) + ((g3172) & (g4003) & (g4004) & (g3157) & (!g5776) & (!g5777)) + ((g3172) & (g4003) & (g4004) & (g3157) & (!g5776) & (g5777)));
	assign g4049 = (((!g2378) & (g3047) & (!g4039)) + ((g2378) & (!g3047) & (!g4039)) + ((g2378) & (g3047) & (!g4039)) + ((g2378) & (g3047) & (g4039)));
	assign g4050 = (((!g830) & (key[165]) & (!g1914) & (!g4048) & (!g4049) & (!g5670)) + ((!g830) & (key[165]) & (!g1914) & (!g4048) & (!g4049) & (g5670)) + ((!g830) & (key[165]) & (!g1914) & (!g4048) & (g4049) & (!g5670)) + ((!g830) & (key[165]) & (!g1914) & (!g4048) & (g4049) & (g5670)) + ((!g830) & (key[165]) & (!g1914) & (g4048) & (!g4049) & (!g5670)) + ((!g830) & (key[165]) & (!g1914) & (g4048) & (!g4049) & (g5670)) + ((!g830) & (key[165]) & (!g1914) & (g4048) & (g4049) & (!g5670)) + ((!g830) & (key[165]) & (!g1914) & (g4048) & (g4049) & (g5670)) + ((!g830) & (key[165]) & (g1914) & (!g4048) & (!g4049) & (!g5670)) + ((!g830) & (key[165]) & (g1914) & (!g4048) & (!g4049) & (g5670)) + ((!g830) & (key[165]) & (g1914) & (!g4048) & (g4049) & (!g5670)) + ((!g830) & (key[165]) & (g1914) & (!g4048) & (g4049) & (g5670)) + ((!g830) & (key[165]) & (g1914) & (g4048) & (!g4049) & (!g5670)) + ((!g830) & (key[165]) & (g1914) & (g4048) & (!g4049) & (g5670)) + ((!g830) & (key[165]) & (g1914) & (g4048) & (g4049) & (!g5670)) + ((!g830) & (key[165]) & (g1914) & (g4048) & (g4049) & (g5670)) + ((g830) & (!key[165]) & (!g1914) & (!g4048) & (!g4049) & (!g5670)) + ((g830) & (!key[165]) & (!g1914) & (!g4048) & (g4049) & (g5670)) + ((g830) & (!key[165]) & (!g1914) & (g4048) & (!g4049) & (!g5670)) + ((g830) & (!key[165]) & (!g1914) & (g4048) & (g4049) & (g5670)) + ((g830) & (!key[165]) & (g1914) & (!g4048) & (!g4049) & (!g5670)) + ((g830) & (!key[165]) & (g1914) & (!g4048) & (g4049) & (!g5670)) + ((g830) & (!key[165]) & (g1914) & (g4048) & (!g4049) & (g5670)) + ((g830) & (!key[165]) & (g1914) & (g4048) & (g4049) & (g5670)) + ((g830) & (key[165]) & (!g1914) & (!g4048) & (!g4049) & (!g5670)) + ((g830) & (key[165]) & (!g1914) & (!g4048) & (g4049) & (g5670)) + ((g830) & (key[165]) & (!g1914) & (g4048) & (!g4049) & (!g5670)) + ((g830) & (key[165]) & (!g1914) & (g4048) & (g4049) & (g5670)) + ((g830) & (key[165]) & (g1914) & (!g4048) & (!g4049) & (!g5670)) + ((g830) & (key[165]) & (g1914) & (!g4048) & (g4049) & (!g5670)) + ((g830) & (key[165]) & (g1914) & (g4048) & (!g4049) & (g5670)) + ((g830) & (key[165]) & (g1914) & (g4048) & (g4049) & (g5670)));
	assign g4051 = (((!g3274) & (!g3235) & (!g3295) & (g3299) & (!g4042)) + ((!g3274) & (!g3235) & (!g3295) & (g3299) & (g4042)) + ((!g3274) & (!g3235) & (g3295) & (!g3299) & (!g4042)) + ((!g3274) & (!g3235) & (g3295) & (!g3299) & (g4042)) + ((!g3274) & (g3235) & (!g3295) & (!g3299) & (!g4042)) + ((!g3274) & (g3235) & (!g3295) & (g3299) & (g4042)) + ((!g3274) & (g3235) & (g3295) & (!g3299) & (g4042)) + ((!g3274) & (g3235) & (g3295) & (g3299) & (!g4042)) + ((g3274) & (!g3235) & (!g3295) & (!g3299) & (!g4042)) + ((g3274) & (!g3235) & (!g3295) & (g3299) & (g4042)) + ((g3274) & (!g3235) & (g3295) & (!g3299) & (g4042)) + ((g3274) & (!g3235) & (g3295) & (g3299) & (!g4042)) + ((g3274) & (g3235) & (!g3295) & (!g3299) & (!g4042)) + ((g3274) & (g3235) & (!g3295) & (!g3299) & (g4042)) + ((g3274) & (g3235) & (g3295) & (g3299) & (!g4042)) + ((g3274) & (g3235) & (g3295) & (g3299) & (g4042)));
	assign g4052 = (((!g1778) & (!g1814) & (!g3222) & (g3301) & (!g4044)) + ((!g1778) & (!g1814) & (!g3222) & (g3301) & (g4044)) + ((!g1778) & (!g1814) & (g3222) & (!g3301) & (!g4044)) + ((!g1778) & (!g1814) & (g3222) & (g3301) & (g4044)) + ((!g1778) & (g1814) & (!g3222) & (!g3301) & (!g4044)) + ((!g1778) & (g1814) & (!g3222) & (!g3301) & (g4044)) + ((!g1778) & (g1814) & (g3222) & (!g3301) & (g4044)) + ((!g1778) & (g1814) & (g3222) & (g3301) & (!g4044)) + ((g1778) & (!g1814) & (!g3222) & (!g3301) & (!g4044)) + ((g1778) & (!g1814) & (!g3222) & (g3301) & (g4044)) + ((g1778) & (!g1814) & (g3222) & (!g3301) & (!g4044)) + ((g1778) & (!g1814) & (g3222) & (!g3301) & (g4044)) + ((g1778) & (g1814) & (!g3222) & (!g3301) & (g4044)) + ((g1778) & (g1814) & (!g3222) & (g3301) & (!g4044)) + ((g1778) & (g1814) & (g3222) & (g3301) & (!g4044)) + ((g1778) & (g1814) & (g3222) & (g3301) & (g4044)));
	assign g8283 = (((!g5560) & (g5575) & (!g4053)) + ((!g5560) & (g5575) & (g4053)) + ((g5560) & (!g5575) & (g4053)) + ((g5560) & (g5575) & (g4053)));
	assign g4054 = (((!g830) & (!g1914) & (!g1991) & (!g4051) & (!g4052) & (g4053)) + ((!g830) & (!g1914) & (!g1991) & (!g4051) & (g4052) & (g4053)) + ((!g830) & (!g1914) & (!g1991) & (g4051) & (!g4052) & (g4053)) + ((!g830) & (!g1914) & (!g1991) & (g4051) & (g4052) & (g4053)) + ((!g830) & (!g1914) & (g1991) & (!g4051) & (!g4052) & (g4053)) + ((!g830) & (!g1914) & (g1991) & (!g4051) & (g4052) & (g4053)) + ((!g830) & (!g1914) & (g1991) & (g4051) & (!g4052) & (g4053)) + ((!g830) & (!g1914) & (g1991) & (g4051) & (g4052) & (g4053)) + ((!g830) & (g1914) & (!g1991) & (!g4051) & (!g4052) & (g4053)) + ((!g830) & (g1914) & (!g1991) & (!g4051) & (g4052) & (g4053)) + ((!g830) & (g1914) & (!g1991) & (g4051) & (!g4052) & (g4053)) + ((!g830) & (g1914) & (!g1991) & (g4051) & (g4052) & (g4053)) + ((!g830) & (g1914) & (g1991) & (!g4051) & (!g4052) & (g4053)) + ((!g830) & (g1914) & (g1991) & (!g4051) & (g4052) & (g4053)) + ((!g830) & (g1914) & (g1991) & (g4051) & (!g4052) & (g4053)) + ((!g830) & (g1914) & (g1991) & (g4051) & (g4052) & (g4053)) + ((g830) & (!g1914) & (!g1991) & (!g4051) & (g4052) & (!g4053)) + ((g830) & (!g1914) & (!g1991) & (!g4051) & (g4052) & (g4053)) + ((g830) & (!g1914) & (!g1991) & (g4051) & (g4052) & (!g4053)) + ((g830) & (!g1914) & (!g1991) & (g4051) & (g4052) & (g4053)) + ((g830) & (!g1914) & (g1991) & (!g4051) & (!g4052) & (!g4053)) + ((g830) & (!g1914) & (g1991) & (!g4051) & (!g4052) & (g4053)) + ((g830) & (!g1914) & (g1991) & (g4051) & (!g4052) & (!g4053)) + ((g830) & (!g1914) & (g1991) & (g4051) & (!g4052) & (g4053)) + ((g830) & (g1914) & (!g1991) & (g4051) & (!g4052) & (!g4053)) + ((g830) & (g1914) & (!g1991) & (g4051) & (!g4052) & (g4053)) + ((g830) & (g1914) & (!g1991) & (g4051) & (g4052) & (!g4053)) + ((g830) & (g1914) & (!g1991) & (g4051) & (g4052) & (g4053)) + ((g830) & (g1914) & (g1991) & (!g4051) & (!g4052) & (!g4053)) + ((g830) & (g1914) & (g1991) & (!g4051) & (!g4052) & (g4053)) + ((g830) & (g1914) & (g1991) & (!g4051) & (g4052) & (!g4053)) + ((g830) & (g1914) & (g1991) & (!g4051) & (g4052) & (g4053)));
	assign g4055 = (((!g3359) & (!g4048) & (!g3336) & (!g3385) & (g3389)) + ((!g3359) & (!g4048) & (!g3336) & (g3385) & (!g3389)) + ((!g3359) & (!g4048) & (g3336) & (!g3385) & (g3389)) + ((!g3359) & (!g4048) & (g3336) & (g3385) & (!g3389)) + ((!g3359) & (g4048) & (!g3336) & (!g3385) & (g3389)) + ((!g3359) & (g4048) & (!g3336) & (g3385) & (!g3389)) + ((!g3359) & (g4048) & (g3336) & (!g3385) & (!g3389)) + ((!g3359) & (g4048) & (g3336) & (g3385) & (g3389)) + ((g3359) & (!g4048) & (!g3336) & (!g3385) & (g3389)) + ((g3359) & (!g4048) & (!g3336) & (g3385) & (!g3389)) + ((g3359) & (!g4048) & (g3336) & (!g3385) & (!g3389)) + ((g3359) & (!g4048) & (g3336) & (g3385) & (g3389)) + ((g3359) & (g4048) & (!g3336) & (!g3385) & (!g3389)) + ((g3359) & (g4048) & (!g3336) & (g3385) & (g3389)) + ((g3359) & (g4048) & (g3336) & (!g3385) & (!g3389)) + ((g3359) & (g4048) & (g3336) & (g3385) & (g3389)));
	assign g4056 = (((!g2426) & (!g2518) & (!g3074) & (g3122) & (!g4049)) + ((!g2426) & (!g2518) & (!g3074) & (g3122) & (g4049)) + ((!g2426) & (!g2518) & (g3074) & (!g3122) & (g4049)) + ((!g2426) & (!g2518) & (g3074) & (g3122) & (!g4049)) + ((!g2426) & (g2518) & (!g3074) & (!g3122) & (!g4049)) + ((!g2426) & (g2518) & (!g3074) & (!g3122) & (g4049)) + ((!g2426) & (g2518) & (g3074) & (!g3122) & (!g4049)) + ((!g2426) & (g2518) & (g3074) & (g3122) & (g4049)) + ((g2426) & (!g2518) & (!g3074) & (!g3122) & (g4049)) + ((g2426) & (!g2518) & (!g3074) & (g3122) & (!g4049)) + ((g2426) & (!g2518) & (g3074) & (!g3122) & (!g4049)) + ((g2426) & (!g2518) & (g3074) & (!g3122) & (g4049)) + ((g2426) & (g2518) & (!g3074) & (!g3122) & (!g4049)) + ((g2426) & (g2518) & (!g3074) & (g3122) & (g4049)) + ((g2426) & (g2518) & (g3074) & (g3122) & (!g4049)) + ((g2426) & (g2518) & (g3074) & (g3122) & (g4049)));
	assign g4057 = (((!g830) & (!g1914) & (!g1992) & (!g4055) & (!g4056) & (key[166])) + ((!g830) & (!g1914) & (!g1992) & (!g4055) & (g4056) & (key[166])) + ((!g830) & (!g1914) & (!g1992) & (g4055) & (!g4056) & (key[166])) + ((!g830) & (!g1914) & (!g1992) & (g4055) & (g4056) & (key[166])) + ((!g830) & (!g1914) & (g1992) & (!g4055) & (!g4056) & (key[166])) + ((!g830) & (!g1914) & (g1992) & (!g4055) & (g4056) & (key[166])) + ((!g830) & (!g1914) & (g1992) & (g4055) & (!g4056) & (key[166])) + ((!g830) & (!g1914) & (g1992) & (g4055) & (g4056) & (key[166])) + ((!g830) & (g1914) & (!g1992) & (!g4055) & (!g4056) & (key[166])) + ((!g830) & (g1914) & (!g1992) & (!g4055) & (g4056) & (key[166])) + ((!g830) & (g1914) & (!g1992) & (g4055) & (!g4056) & (key[166])) + ((!g830) & (g1914) & (!g1992) & (g4055) & (g4056) & (key[166])) + ((!g830) & (g1914) & (g1992) & (!g4055) & (!g4056) & (key[166])) + ((!g830) & (g1914) & (g1992) & (!g4055) & (g4056) & (key[166])) + ((!g830) & (g1914) & (g1992) & (g4055) & (!g4056) & (key[166])) + ((!g830) & (g1914) & (g1992) & (g4055) & (g4056) & (key[166])) + ((g830) & (!g1914) & (!g1992) & (!g4055) & (g4056) & (!key[166])) + ((g830) & (!g1914) & (!g1992) & (!g4055) & (g4056) & (key[166])) + ((g830) & (!g1914) & (!g1992) & (g4055) & (g4056) & (!key[166])) + ((g830) & (!g1914) & (!g1992) & (g4055) & (g4056) & (key[166])) + ((g830) & (!g1914) & (g1992) & (!g4055) & (!g4056) & (!key[166])) + ((g830) & (!g1914) & (g1992) & (!g4055) & (!g4056) & (key[166])) + ((g830) & (!g1914) & (g1992) & (g4055) & (!g4056) & (!key[166])) + ((g830) & (!g1914) & (g1992) & (g4055) & (!g4056) & (key[166])) + ((g830) & (g1914) & (!g1992) & (g4055) & (!g4056) & (!key[166])) + ((g830) & (g1914) & (!g1992) & (g4055) & (!g4056) & (key[166])) + ((g830) & (g1914) & (!g1992) & (g4055) & (g4056) & (!key[166])) + ((g830) & (g1914) & (!g1992) & (g4055) & (g4056) & (key[166])) + ((g830) & (g1914) & (g1992) & (!g4055) & (!g4056) & (!key[166])) + ((g830) & (g1914) & (g1992) & (!g4055) & (!g4056) & (key[166])) + ((g830) & (g1914) & (g1992) & (!g4055) & (g4056) & (!key[166])) + ((g830) & (g1914) & (g1992) & (!g4055) & (g4056) & (key[166])));
	assign g4058 = (((!g3274) & (!g3235) & (g3295) & (g3299) & (!g4042)) + ((!g3274) & (!g3235) & (g3295) & (g3299) & (g4042)) + ((!g3274) & (g3235) & (!g3295) & (g3299) & (!g4042)) + ((!g3274) & (g3235) & (g3295) & (!g3299) & (!g4042)) + ((!g3274) & (g3235) & (g3295) & (g3299) & (!g4042)) + ((!g3274) & (g3235) & (g3295) & (g3299) & (g4042)) + ((g3274) & (!g3235) & (!g3295) & (g3299) & (!g4042)) + ((g3274) & (!g3235) & (g3295) & (!g3299) & (!g4042)) + ((g3274) & (!g3235) & (g3295) & (g3299) & (!g4042)) + ((g3274) & (!g3235) & (g3295) & (g3299) & (g4042)) + ((g3274) & (g3235) & (!g3295) & (g3299) & (!g4042)) + ((g3274) & (g3235) & (!g3295) & (g3299) & (g4042)) + ((g3274) & (g3235) & (g3295) & (!g3299) & (!g4042)) + ((g3274) & (g3235) & (g3295) & (!g3299) & (g4042)) + ((g3274) & (g3235) & (g3295) & (g3299) & (!g4042)) + ((g3274) & (g3235) & (g3295) & (g3299) & (g4042)));
	assign g4059 = (((!g1778) & (!g1814) & (g3222) & (g3301) & (!g4044)) + ((!g1778) & (g1814) & (!g3222) & (g3301) & (!g4044)) + ((!g1778) & (g1814) & (!g3222) & (g3301) & (g4044)) + ((!g1778) & (g1814) & (g3222) & (!g3301) & (!g4044)) + ((!g1778) & (g1814) & (g3222) & (g3301) & (!g4044)) + ((!g1778) & (g1814) & (g3222) & (g3301) & (g4044)) + ((g1778) & (!g1814) & (!g3222) & (g3301) & (!g4044)) + ((g1778) & (!g1814) & (g3222) & (g3301) & (!g4044)) + ((g1778) & (!g1814) & (g3222) & (g3301) & (g4044)) + ((g1778) & (g1814) & (!g3222) & (!g3301) & (!g4044)) + ((g1778) & (g1814) & (!g3222) & (g3301) & (!g4044)) + ((g1778) & (g1814) & (!g3222) & (g3301) & (g4044)) + ((g1778) & (g1814) & (g3222) & (!g3301) & (!g4044)) + ((g1778) & (g1814) & (g3222) & (!g3301) & (g4044)) + ((g1778) & (g1814) & (g3222) & (g3301) & (!g4044)) + ((g1778) & (g1814) & (g3222) & (g3301) & (g4044)));
	assign g8284 = (((!g5560) & (g5576) & (!g4060)) + ((!g5560) & (g5576) & (g4060)) + ((g5560) & (!g5576) & (g4060)) + ((g5560) & (g5576) & (g4060)));
	assign g4061 = (((!g830) & (g4060) & (!g1914) & (!g4058) & (!g4059) & (!g5673)) + ((!g830) & (g4060) & (!g1914) & (!g4058) & (!g4059) & (g5673)) + ((!g830) & (g4060) & (!g1914) & (!g4058) & (g4059) & (!g5673)) + ((!g830) & (g4060) & (!g1914) & (!g4058) & (g4059) & (g5673)) + ((!g830) & (g4060) & (!g1914) & (g4058) & (!g4059) & (!g5673)) + ((!g830) & (g4060) & (!g1914) & (g4058) & (!g4059) & (g5673)) + ((!g830) & (g4060) & (!g1914) & (g4058) & (g4059) & (!g5673)) + ((!g830) & (g4060) & (!g1914) & (g4058) & (g4059) & (g5673)) + ((!g830) & (g4060) & (g1914) & (!g4058) & (!g4059) & (!g5673)) + ((!g830) & (g4060) & (g1914) & (!g4058) & (!g4059) & (g5673)) + ((!g830) & (g4060) & (g1914) & (!g4058) & (g4059) & (!g5673)) + ((!g830) & (g4060) & (g1914) & (!g4058) & (g4059) & (g5673)) + ((!g830) & (g4060) & (g1914) & (g4058) & (!g4059) & (!g5673)) + ((!g830) & (g4060) & (g1914) & (g4058) & (!g4059) & (g5673)) + ((!g830) & (g4060) & (g1914) & (g4058) & (g4059) & (!g5673)) + ((!g830) & (g4060) & (g1914) & (g4058) & (g4059) & (g5673)) + ((g830) & (!g4060) & (!g1914) & (!g4058) & (!g4059) & (!g5673)) + ((g830) & (!g4060) & (!g1914) & (!g4058) & (g4059) & (g5673)) + ((g830) & (!g4060) & (!g1914) & (g4058) & (!g4059) & (!g5673)) + ((g830) & (!g4060) & (!g1914) & (g4058) & (g4059) & (g5673)) + ((g830) & (!g4060) & (g1914) & (!g4058) & (!g4059) & (!g5673)) + ((g830) & (!g4060) & (g1914) & (!g4058) & (g4059) & (!g5673)) + ((g830) & (!g4060) & (g1914) & (g4058) & (!g4059) & (g5673)) + ((g830) & (!g4060) & (g1914) & (g4058) & (g4059) & (g5673)) + ((g830) & (g4060) & (!g1914) & (!g4058) & (!g4059) & (!g5673)) + ((g830) & (g4060) & (!g1914) & (!g4058) & (g4059) & (g5673)) + ((g830) & (g4060) & (!g1914) & (g4058) & (!g4059) & (!g5673)) + ((g830) & (g4060) & (!g1914) & (g4058) & (g4059) & (g5673)) + ((g830) & (g4060) & (g1914) & (!g4058) & (!g4059) & (!g5673)) + ((g830) & (g4060) & (g1914) & (!g4058) & (g4059) & (!g5673)) + ((g830) & (g4060) & (g1914) & (g4058) & (!g4059) & (g5673)) + ((g830) & (g4060) & (g1914) & (g4058) & (g4059) & (g5673)));
	assign g4062 = (((!g2518) & (g3122)) + ((g2518) & (!g3122)));
	assign g4063 = (((!g2378) & (!g2426) & (g3047) & (g3074) & (!g4039) & (g4062)) + ((!g2378) & (g2426) & (!g3047) & (g3074) & (!g4039) & (g4062)) + ((!g2378) & (g2426) & (!g3047) & (g3074) & (g4039) & (g4062)) + ((!g2378) & (g2426) & (g3047) & (!g3074) & (!g4039) & (g4062)) + ((!g2378) & (g2426) & (g3047) & (g3074) & (!g4039) & (g4062)) + ((!g2378) & (g2426) & (g3047) & (g3074) & (g4039) & (g4062)) + ((g2378) & (!g2426) & (!g3047) & (g3074) & (!g4039) & (g4062)) + ((g2378) & (!g2426) & (g3047) & (g3074) & (!g4039) & (g4062)) + ((g2378) & (!g2426) & (g3047) & (g3074) & (g4039) & (g4062)) + ((g2378) & (g2426) & (!g3047) & (!g3074) & (!g4039) & (g4062)) + ((g2378) & (g2426) & (!g3047) & (g3074) & (!g4039) & (g4062)) + ((g2378) & (g2426) & (!g3047) & (g3074) & (g4039) & (g4062)) + ((g2378) & (g2426) & (g3047) & (!g3074) & (!g4039) & (g4062)) + ((g2378) & (g2426) & (g3047) & (!g3074) & (g4039) & (g4062)) + ((g2378) & (g2426) & (g3047) & (g3074) & (!g4039) & (g4062)) + ((g2378) & (g2426) & (g3047) & (g3074) & (g4039) & (g4062)));
	assign g4064 = (((g2518) & (g3122)));
	assign g4065 = (((!g2555) & (!g3149) & (!g4063) & (g4064)) + ((!g2555) & (!g3149) & (g4063) & (!g4064)) + ((!g2555) & (!g3149) & (g4063) & (g4064)) + ((!g2555) & (g3149) & (!g4063) & (!g4064)) + ((g2555) & (!g3149) & (!g4063) & (!g4064)) + ((g2555) & (g3149) & (!g4063) & (g4064)) + ((g2555) & (g3149) & (g4063) & (!g4064)) + ((g2555) & (g3149) & (g4063) & (g4064)));
	assign g4066 = (((!g3353) & (!g3330) & (!g3370) & (g3374) & (!g4058)) + ((!g3353) & (!g3330) & (!g3370) & (g3374) & (g4058)) + ((!g3353) & (!g3330) & (g3370) & (!g3374) & (!g4058)) + ((!g3353) & (!g3330) & (g3370) & (!g3374) & (g4058)) + ((!g3353) & (g3330) & (!g3370) & (!g3374) & (g4058)) + ((!g3353) & (g3330) & (!g3370) & (g3374) & (!g4058)) + ((!g3353) & (g3330) & (g3370) & (!g3374) & (!g4058)) + ((!g3353) & (g3330) & (g3370) & (g3374) & (g4058)) + ((g3353) & (!g3330) & (!g3370) & (!g3374) & (g4058)) + ((g3353) & (!g3330) & (!g3370) & (g3374) & (!g4058)) + ((g3353) & (!g3330) & (g3370) & (!g3374) & (!g4058)) + ((g3353) & (!g3330) & (g3370) & (g3374) & (g4058)) + ((g3353) & (g3330) & (!g3370) & (!g3374) & (!g4058)) + ((g3353) & (g3330) & (!g3370) & (!g3374) & (g4058)) + ((g3353) & (g3330) & (g3370) & (g3374) & (!g4058)) + ((g3353) & (g3330) & (g3370) & (g3374) & (g4058)));
	assign g4067 = (((!g1847) & (!g1881) & (!g3323) & (g3376) & (!g4059)) + ((!g1847) & (!g1881) & (!g3323) & (g3376) & (g4059)) + ((!g1847) & (!g1881) & (g3323) & (!g3376) & (g4059)) + ((!g1847) & (!g1881) & (g3323) & (g3376) & (!g4059)) + ((!g1847) & (g1881) & (!g3323) & (!g3376) & (!g4059)) + ((!g1847) & (g1881) & (!g3323) & (!g3376) & (g4059)) + ((!g1847) & (g1881) & (g3323) & (!g3376) & (!g4059)) + ((!g1847) & (g1881) & (g3323) & (g3376) & (g4059)) + ((g1847) & (!g1881) & (!g3323) & (!g3376) & (g4059)) + ((g1847) & (!g1881) & (!g3323) & (g3376) & (!g4059)) + ((g1847) & (!g1881) & (g3323) & (!g3376) & (!g4059)) + ((g1847) & (!g1881) & (g3323) & (!g3376) & (g4059)) + ((g1847) & (g1881) & (!g3323) & (!g3376) & (!g4059)) + ((g1847) & (g1881) & (!g3323) & (g3376) & (g4059)) + ((g1847) & (g1881) & (g3323) & (g3376) & (!g4059)) + ((g1847) & (g1881) & (g3323) & (g3376) & (g4059)));
	assign g8285 = (((!g5560) & (g5577) & (!g4068)) + ((!g5560) & (g5577) & (g4068)) + ((g5560) & (!g5577) & (g4068)) + ((g5560) & (g5577) & (g4068)));
	assign g4069 = (((!g830) & (!g1914) & (!g1996) & (!g4066) & (!g4067) & (g4068)) + ((!g830) & (!g1914) & (!g1996) & (!g4066) & (g4067) & (g4068)) + ((!g830) & (!g1914) & (!g1996) & (g4066) & (!g4067) & (g4068)) + ((!g830) & (!g1914) & (!g1996) & (g4066) & (g4067) & (g4068)) + ((!g830) & (!g1914) & (g1996) & (!g4066) & (!g4067) & (g4068)) + ((!g830) & (!g1914) & (g1996) & (!g4066) & (g4067) & (g4068)) + ((!g830) & (!g1914) & (g1996) & (g4066) & (!g4067) & (g4068)) + ((!g830) & (!g1914) & (g1996) & (g4066) & (g4067) & (g4068)) + ((!g830) & (g1914) & (!g1996) & (!g4066) & (!g4067) & (g4068)) + ((!g830) & (g1914) & (!g1996) & (!g4066) & (g4067) & (g4068)) + ((!g830) & (g1914) & (!g1996) & (g4066) & (!g4067) & (g4068)) + ((!g830) & (g1914) & (!g1996) & (g4066) & (g4067) & (g4068)) + ((!g830) & (g1914) & (g1996) & (!g4066) & (!g4067) & (g4068)) + ((!g830) & (g1914) & (g1996) & (!g4066) & (g4067) & (g4068)) + ((!g830) & (g1914) & (g1996) & (g4066) & (!g4067) & (g4068)) + ((!g830) & (g1914) & (g1996) & (g4066) & (g4067) & (g4068)) + ((g830) & (!g1914) & (!g1996) & (!g4066) & (g4067) & (!g4068)) + ((g830) & (!g1914) & (!g1996) & (!g4066) & (g4067) & (g4068)) + ((g830) & (!g1914) & (!g1996) & (g4066) & (g4067) & (!g4068)) + ((g830) & (!g1914) & (!g1996) & (g4066) & (g4067) & (g4068)) + ((g830) & (!g1914) & (g1996) & (!g4066) & (!g4067) & (!g4068)) + ((g830) & (!g1914) & (g1996) & (!g4066) & (!g4067) & (g4068)) + ((g830) & (!g1914) & (g1996) & (g4066) & (!g4067) & (!g4068)) + ((g830) & (!g1914) & (g1996) & (g4066) & (!g4067) & (g4068)) + ((g830) & (g1914) & (!g1996) & (g4066) & (!g4067) & (!g4068)) + ((g830) & (g1914) & (!g1996) & (g4066) & (!g4067) & (g4068)) + ((g830) & (g1914) & (!g1996) & (g4066) & (g4067) & (!g4068)) + ((g830) & (g1914) & (!g1996) & (g4066) & (g4067) & (g4068)) + ((g830) & (g1914) & (g1996) & (!g4066) & (!g4067) & (!g4068)) + ((g830) & (g1914) & (g1996) & (!g4066) & (!g4067) & (g4068)) + ((g830) & (g1914) & (g1996) & (!g4066) & (g4067) & (!g4068)) + ((g830) & (g1914) & (g1996) & (!g4066) & (g4067) & (g4068)));
	assign g4070 = (((!g1896) & (!g1912) & (!g2041) & (g2045)) + ((!g1896) & (!g1912) & (g2041) & (!g2045)) + ((!g1896) & (g1912) & (!g2041) & (g2045)) + ((!g1896) & (g1912) & (g2041) & (!g2045)) + ((g1896) & (!g1912) & (!g2041) & (g2045)) + ((g1896) & (!g1912) & (g2041) & (!g2045)) + ((g1896) & (g1912) & (!g2041) & (!g2045)) + ((g1896) & (g1912) & (g2041) & (g2045)));
	assign g4071 = (((!g2555) & (!g3149) & (!g4063) & (!g4064)) + ((!g2555) & (!g3149) & (!g4063) & (g4064)) + ((!g2555) & (!g3149) & (g4063) & (!g4064)) + ((!g2555) & (!g3149) & (g4063) & (g4064)) + ((!g2555) & (g3149) & (!g4063) & (!g4064)) + ((g2555) & (!g3149) & (!g4063) & (!g4064)));
	assign g4072 = (((!g1914) & (!g2601) & (!g3193) & (!g4070) & (!g4071)) + ((!g1914) & (!g2601) & (!g3193) & (g4070) & (!g4071)) + ((!g1914) & (!g2601) & (g3193) & (!g4070) & (g4071)) + ((!g1914) & (!g2601) & (g3193) & (g4070) & (g4071)) + ((!g1914) & (g2601) & (!g3193) & (!g4070) & (g4071)) + ((!g1914) & (g2601) & (!g3193) & (g4070) & (g4071)) + ((!g1914) & (g2601) & (g3193) & (!g4070) & (!g4071)) + ((!g1914) & (g2601) & (g3193) & (g4070) & (!g4071)) + ((g1914) & (!g2601) & (!g3193) & (g4070) & (!g4071)) + ((g1914) & (!g2601) & (!g3193) & (g4070) & (g4071)) + ((g1914) & (!g2601) & (g3193) & (g4070) & (!g4071)) + ((g1914) & (!g2601) & (g3193) & (g4070) & (g4071)) + ((g1914) & (g2601) & (!g3193) & (g4070) & (!g4071)) + ((g1914) & (g2601) & (!g3193) & (g4070) & (g4071)) + ((g1914) & (g2601) & (g3193) & (g4070) & (!g4071)) + ((g1914) & (g2601) & (g3193) & (g4070) & (g4071)));
	assign g4073 = (((!g830) & (!g1997) & (!g4072) & (key[168])) + ((!g830) & (!g1997) & (g4072) & (key[168])) + ((!g830) & (g1997) & (!g4072) & (key[168])) + ((!g830) & (g1997) & (g4072) & (key[168])) + ((g830) & (!g1997) & (g4072) & (!key[168])) + ((g830) & (!g1997) & (g4072) & (key[168])) + ((g830) & (g1997) & (!g4072) & (!key[168])) + ((g830) & (g1997) & (!g4072) & (key[168])));
	assign g4074 = (((!g1914) & (!g828) & (!g1892) & (!g1908) & (g1886)) + ((!g1914) & (!g828) & (!g1892) & (g1908) & (g1886)) + ((!g1914) & (!g828) & (g1892) & (!g1908) & (g1886)) + ((!g1914) & (!g828) & (g1892) & (g1908) & (g1886)) + ((!g1914) & (g828) & (!g1892) & (!g1908) & (!g1886)) + ((!g1914) & (g828) & (!g1892) & (g1908) & (!g1886)) + ((!g1914) & (g828) & (g1892) & (!g1908) & (!g1886)) + ((!g1914) & (g828) & (g1892) & (g1908) & (!g1886)) + ((g1914) & (!g828) & (!g1892) & (g1908) & (!g1886)) + ((g1914) & (!g828) & (!g1892) & (g1908) & (g1886)) + ((g1914) & (!g828) & (g1892) & (!g1908) & (!g1886)) + ((g1914) & (!g828) & (g1892) & (!g1908) & (g1886)) + ((g1914) & (g828) & (!g1892) & (g1908) & (!g1886)) + ((g1914) & (g828) & (!g1892) & (g1908) & (g1886)) + ((g1914) & (g828) & (g1892) & (!g1908) & (!g1886)) + ((g1914) & (g828) & (g1892) & (!g1908) & (g1886)));
	assign g8286 = (((!g5560) & (g5578) & (!g4075)) + ((!g5560) & (g5578) & (g4075)) + ((g5560) & (!g5578) & (g4075)) + ((g5560) & (g5578) & (g4075)));
	assign g4076 = (((!g830) & (!g1998) & (!g4074) & (g4075)) + ((!g830) & (!g1998) & (g4074) & (g4075)) + ((!g830) & (g1998) & (!g4074) & (g4075)) + ((!g830) & (g1998) & (g4074) & (g4075)) + ((g830) & (!g1998) & (g4074) & (!g4075)) + ((g830) & (!g1998) & (g4074) & (g4075)) + ((g830) & (g1998) & (!g4074) & (!g4075)) + ((g830) & (g1998) & (!g4074) & (g4075)));
	assign g4077 = (((!g1896) & (!g1912) & (!g2041) & (!g2045) & (!g2068) & (g2091)) + ((!g1896) & (!g1912) & (!g2041) & (!g2045) & (g2068) & (!g2091)) + ((!g1896) & (!g1912) & (!g2041) & (g2045) & (!g2068) & (g2091)) + ((!g1896) & (!g1912) & (!g2041) & (g2045) & (g2068) & (!g2091)) + ((!g1896) & (!g1912) & (g2041) & (!g2045) & (!g2068) & (g2091)) + ((!g1896) & (!g1912) & (g2041) & (!g2045) & (g2068) & (!g2091)) + ((!g1896) & (!g1912) & (g2041) & (g2045) & (!g2068) & (!g2091)) + ((!g1896) & (!g1912) & (g2041) & (g2045) & (g2068) & (g2091)) + ((!g1896) & (g1912) & (!g2041) & (!g2045) & (!g2068) & (g2091)) + ((!g1896) & (g1912) & (!g2041) & (!g2045) & (g2068) & (!g2091)) + ((!g1896) & (g1912) & (!g2041) & (g2045) & (!g2068) & (g2091)) + ((!g1896) & (g1912) & (!g2041) & (g2045) & (g2068) & (!g2091)) + ((!g1896) & (g1912) & (g2041) & (!g2045) & (!g2068) & (g2091)) + ((!g1896) & (g1912) & (g2041) & (!g2045) & (g2068) & (!g2091)) + ((!g1896) & (g1912) & (g2041) & (g2045) & (!g2068) & (!g2091)) + ((!g1896) & (g1912) & (g2041) & (g2045) & (g2068) & (g2091)) + ((g1896) & (!g1912) & (!g2041) & (!g2045) & (!g2068) & (g2091)) + ((g1896) & (!g1912) & (!g2041) & (!g2045) & (g2068) & (!g2091)) + ((g1896) & (!g1912) & (!g2041) & (g2045) & (!g2068) & (g2091)) + ((g1896) & (!g1912) & (!g2041) & (g2045) & (g2068) & (!g2091)) + ((g1896) & (!g1912) & (g2041) & (!g2045) & (!g2068) & (g2091)) + ((g1896) & (!g1912) & (g2041) & (!g2045) & (g2068) & (!g2091)) + ((g1896) & (!g1912) & (g2041) & (g2045) & (!g2068) & (!g2091)) + ((g1896) & (!g1912) & (g2041) & (g2045) & (g2068) & (g2091)) + ((g1896) & (g1912) & (!g2041) & (!g2045) & (!g2068) & (g2091)) + ((g1896) & (g1912) & (!g2041) & (!g2045) & (g2068) & (!g2091)) + ((g1896) & (g1912) & (!g2041) & (g2045) & (!g2068) & (!g2091)) + ((g1896) & (g1912) & (!g2041) & (g2045) & (g2068) & (g2091)) + ((g1896) & (g1912) & (g2041) & (!g2045) & (!g2068) & (!g2091)) + ((g1896) & (g1912) & (g2041) & (!g2045) & (g2068) & (g2091)) + ((g1896) & (g1912) & (g2041) & (g2045) & (!g2068) & (!g2091)) + ((g1896) & (g1912) & (g2041) & (g2045) & (g2068) & (g2091)));
	assign g4078 = (((!g2555) & (!g2601) & (!g3149) & (!g3193) & (!g4063) & (!g4064)) + ((!g2555) & (!g2601) & (!g3149) & (!g3193) & (!g4063) & (g4064)) + ((!g2555) & (!g2601) & (!g3149) & (!g3193) & (g4063) & (!g4064)) + ((!g2555) & (!g2601) & (!g3149) & (!g3193) & (g4063) & (g4064)) + ((!g2555) & (!g2601) & (!g3149) & (g3193) & (!g4063) & (!g4064)) + ((!g2555) & (!g2601) & (!g3149) & (g3193) & (!g4063) & (g4064)) + ((!g2555) & (!g2601) & (!g3149) & (g3193) & (g4063) & (!g4064)) + ((!g2555) & (!g2601) & (!g3149) & (g3193) & (g4063) & (g4064)) + ((!g2555) & (!g2601) & (g3149) & (!g3193) & (!g4063) & (!g4064)) + ((!g2555) & (!g2601) & (g3149) & (!g3193) & (!g4063) & (g4064)) + ((!g2555) & (!g2601) & (g3149) & (!g3193) & (g4063) & (!g4064)) + ((!g2555) & (!g2601) & (g3149) & (!g3193) & (g4063) & (g4064)) + ((!g2555) & (!g2601) & (g3149) & (g3193) & (!g4063) & (!g4064)) + ((!g2555) & (g2601) & (!g3149) & (!g3193) & (!g4063) & (!g4064)) + ((!g2555) & (g2601) & (!g3149) & (!g3193) & (!g4063) & (g4064)) + ((!g2555) & (g2601) & (!g3149) & (!g3193) & (g4063) & (!g4064)) + ((!g2555) & (g2601) & (!g3149) & (!g3193) & (g4063) & (g4064)) + ((!g2555) & (g2601) & (g3149) & (!g3193) & (!g4063) & (!g4064)) + ((g2555) & (!g2601) & (!g3149) & (!g3193) & (!g4063) & (!g4064)) + ((g2555) & (!g2601) & (!g3149) & (!g3193) & (!g4063) & (g4064)) + ((g2555) & (!g2601) & (!g3149) & (!g3193) & (g4063) & (!g4064)) + ((g2555) & (!g2601) & (!g3149) & (!g3193) & (g4063) & (g4064)) + ((g2555) & (!g2601) & (!g3149) & (g3193) & (!g4063) & (!g4064)) + ((g2555) & (!g2601) & (g3149) & (!g3193) & (!g4063) & (!g4064)) + ((g2555) & (!g2601) & (g3149) & (!g3193) & (!g4063) & (g4064)) + ((g2555) & (!g2601) & (g3149) & (!g3193) & (g4063) & (!g4064)) + ((g2555) & (!g2601) & (g3149) & (!g3193) & (g4063) & (g4064)) + ((g2555) & (g2601) & (!g3149) & (!g3193) & (!g4063) & (!g4064)));
	assign g4079 = (((!g1914) & (!g2649) & (!g3222) & (!g4077) & (!g4078)) + ((!g1914) & (!g2649) & (!g3222) & (g4077) & (!g4078)) + ((!g1914) & (!g2649) & (g3222) & (!g4077) & (g4078)) + ((!g1914) & (!g2649) & (g3222) & (g4077) & (g4078)) + ((!g1914) & (g2649) & (!g3222) & (!g4077) & (g4078)) + ((!g1914) & (g2649) & (!g3222) & (g4077) & (g4078)) + ((!g1914) & (g2649) & (g3222) & (!g4077) & (!g4078)) + ((!g1914) & (g2649) & (g3222) & (g4077) & (!g4078)) + ((g1914) & (!g2649) & (!g3222) & (g4077) & (!g4078)) + ((g1914) & (!g2649) & (!g3222) & (g4077) & (g4078)) + ((g1914) & (!g2649) & (g3222) & (g4077) & (!g4078)) + ((g1914) & (!g2649) & (g3222) & (g4077) & (g4078)) + ((g1914) & (g2649) & (!g3222) & (g4077) & (!g4078)) + ((g1914) & (g2649) & (!g3222) & (g4077) & (g4078)) + ((g1914) & (g2649) & (g3222) & (g4077) & (!g4078)) + ((g1914) & (g2649) & (g3222) & (g4077) & (g4078)));
	assign g4080 = (((!g830) & (!g1999) & (!g4079) & (key[169])) + ((!g830) & (!g1999) & (g4079) & (key[169])) + ((!g830) & (g1999) & (!g4079) & (key[169])) + ((!g830) & (g1999) & (g4079) & (key[169])) + ((g830) & (!g1999) & (g4079) & (!key[169])) + ((g830) & (!g1999) & (g4079) & (key[169])) + ((g830) & (g1999) & (!g4079) & (!key[169])) + ((g830) & (g1999) & (!g4079) & (key[169])));
	assign g4081 = (((g1914) & (!g1892) & (!g1908) & (!g2026) & (g2030)) + ((g1914) & (!g1892) & (!g1908) & (g2026) & (!g2030)) + ((g1914) & (!g1892) & (g1908) & (!g2026) & (g2030)) + ((g1914) & (!g1892) & (g1908) & (g2026) & (!g2030)) + ((g1914) & (g1892) & (!g1908) & (!g2026) & (g2030)) + ((g1914) & (g1892) & (!g1908) & (g2026) & (!g2030)) + ((g1914) & (g1892) & (g1908) & (!g2026) & (!g2030)) + ((g1914) & (g1892) & (g1908) & (g2026) & (g2030)));
	assign g4082 = (((!g1914) & (!g828) & (!g864) & (!g1886) & (g2032)) + ((!g1914) & (!g828) & (!g864) & (g1886) & (g2032)) + ((!g1914) & (!g828) & (g864) & (!g1886) & (!g2032)) + ((!g1914) & (!g828) & (g864) & (g1886) & (!g2032)) + ((!g1914) & (g828) & (!g864) & (!g1886) & (g2032)) + ((!g1914) & (g828) & (!g864) & (g1886) & (!g2032)) + ((!g1914) & (g828) & (g864) & (!g1886) & (!g2032)) + ((!g1914) & (g828) & (g864) & (g1886) & (g2032)));
	assign g8287 = (((!g5560) & (g5579) & (!g4083)) + ((!g5560) & (g5579) & (g4083)) + ((g5560) & (!g5579) & (g4083)) + ((g5560) & (g5579) & (g4083)));
	assign g4084 = (((!g830) & (!g2001) & (!g4081) & (!g4082) & (g4083)) + ((!g830) & (!g2001) & (!g4081) & (g4082) & (g4083)) + ((!g830) & (!g2001) & (g4081) & (!g4082) & (g4083)) + ((!g830) & (!g2001) & (g4081) & (g4082) & (g4083)) + ((!g830) & (g2001) & (!g4081) & (!g4082) & (g4083)) + ((!g830) & (g2001) & (!g4081) & (g4082) & (g4083)) + ((!g830) & (g2001) & (g4081) & (!g4082) & (g4083)) + ((!g830) & (g2001) & (g4081) & (g4082) & (g4083)) + ((g830) & (!g2001) & (!g4081) & (g4082) & (!g4083)) + ((g830) & (!g2001) & (!g4081) & (g4082) & (g4083)) + ((g830) & (!g2001) & (g4081) & (!g4082) & (!g4083)) + ((g830) & (!g2001) & (g4081) & (!g4082) & (g4083)) + ((g830) & (!g2001) & (g4081) & (g4082) & (!g4083)) + ((g830) & (!g2001) & (g4081) & (g4082) & (g4083)) + ((g830) & (g2001) & (!g4081) & (!g4082) & (!g4083)) + ((g830) & (g2001) & (!g4081) & (!g4082) & (g4083)));
	assign g4085 = (((!g3465) & (!g2123) & (g2127)) + ((!g3465) & (g2123) & (!g2127)) + ((g3465) & (!g2123) & (!g2127)) + ((g3465) & (g2123) & (g2127)));
	assign g4086 = (((!g2649) & (!g2683) & (!g3222) & (g3301) & (!g4078)) + ((!g2649) & (!g2683) & (!g3222) & (g3301) & (g4078)) + ((!g2649) & (!g2683) & (g3222) & (!g3301) & (!g4078)) + ((!g2649) & (!g2683) & (g3222) & (g3301) & (g4078)) + ((!g2649) & (g2683) & (!g3222) & (!g3301) & (!g4078)) + ((!g2649) & (g2683) & (!g3222) & (!g3301) & (g4078)) + ((!g2649) & (g2683) & (g3222) & (!g3301) & (g4078)) + ((!g2649) & (g2683) & (g3222) & (g3301) & (!g4078)) + ((g2649) & (!g2683) & (!g3222) & (!g3301) & (!g4078)) + ((g2649) & (!g2683) & (!g3222) & (g3301) & (g4078)) + ((g2649) & (!g2683) & (g3222) & (!g3301) & (!g4078)) + ((g2649) & (!g2683) & (g3222) & (!g3301) & (g4078)) + ((g2649) & (g2683) & (!g3222) & (!g3301) & (g4078)) + ((g2649) & (g2683) & (!g3222) & (g3301) & (!g4078)) + ((g2649) & (g2683) & (g3222) & (g3301) & (!g4078)) + ((g2649) & (g2683) & (g3222) & (g3301) & (g4078)));
	assign g4087 = (((!g830) & (!g1914) & (!g2002) & (!g4085) & (!g4086) & (key[170])) + ((!g830) & (!g1914) & (!g2002) & (!g4085) & (g4086) & (key[170])) + ((!g830) & (!g1914) & (!g2002) & (g4085) & (!g4086) & (key[170])) + ((!g830) & (!g1914) & (!g2002) & (g4085) & (g4086) & (key[170])) + ((!g830) & (!g1914) & (g2002) & (!g4085) & (!g4086) & (key[170])) + ((!g830) & (!g1914) & (g2002) & (!g4085) & (g4086) & (key[170])) + ((!g830) & (!g1914) & (g2002) & (g4085) & (!g4086) & (key[170])) + ((!g830) & (!g1914) & (g2002) & (g4085) & (g4086) & (key[170])) + ((!g830) & (g1914) & (!g2002) & (!g4085) & (!g4086) & (key[170])) + ((!g830) & (g1914) & (!g2002) & (!g4085) & (g4086) & (key[170])) + ((!g830) & (g1914) & (!g2002) & (g4085) & (!g4086) & (key[170])) + ((!g830) & (g1914) & (!g2002) & (g4085) & (g4086) & (key[170])) + ((!g830) & (g1914) & (g2002) & (!g4085) & (!g4086) & (key[170])) + ((!g830) & (g1914) & (g2002) & (!g4085) & (g4086) & (key[170])) + ((!g830) & (g1914) & (g2002) & (g4085) & (!g4086) & (key[170])) + ((!g830) & (g1914) & (g2002) & (g4085) & (g4086) & (key[170])) + ((g830) & (!g1914) & (!g2002) & (!g4085) & (g4086) & (!key[170])) + ((g830) & (!g1914) & (!g2002) & (!g4085) & (g4086) & (key[170])) + ((g830) & (!g1914) & (!g2002) & (g4085) & (g4086) & (!key[170])) + ((g830) & (!g1914) & (!g2002) & (g4085) & (g4086) & (key[170])) + ((g830) & (!g1914) & (g2002) & (!g4085) & (!g4086) & (!key[170])) + ((g830) & (!g1914) & (g2002) & (!g4085) & (!g4086) & (key[170])) + ((g830) & (!g1914) & (g2002) & (g4085) & (!g4086) & (!key[170])) + ((g830) & (!g1914) & (g2002) & (g4085) & (!g4086) & (key[170])) + ((g830) & (g1914) & (!g2002) & (g4085) & (!g4086) & (!key[170])) + ((g830) & (g1914) & (!g2002) & (g4085) & (!g4086) & (key[170])) + ((g830) & (g1914) & (!g2002) & (g4085) & (g4086) & (!key[170])) + ((g830) & (g1914) & (!g2002) & (g4085) & (g4086) & (key[170])) + ((g830) & (g1914) & (g2002) & (!g4085) & (!g4086) & (!key[170])) + ((g830) & (g1914) & (g2002) & (!g4085) & (!g4086) & (key[170])) + ((g830) & (g1914) & (g2002) & (!g4085) & (g4086) & (!key[170])) + ((g830) & (g1914) & (g2002) & (!g4085) & (g4086) & (key[170])));
	assign g4088 = (((!g828) & (g864) & (!g1886) & (g2032)) + ((!g828) & (g864) & (g1886) & (g2032)) + ((g828) & (!g864) & (g1886) & (g2032)) + ((g828) & (g864) & (!g1886) & (g2032)) + ((g828) & (g864) & (g1886) & (!g2032)) + ((g828) & (g864) & (g1886) & (g2032)));
	assign g4089 = (((!g1892) & (!g1908) & (!g2026) & (!g2030) & (!g2062) & (g2085)) + ((!g1892) & (!g1908) & (!g2026) & (!g2030) & (g2062) & (!g2085)) + ((!g1892) & (!g1908) & (!g2026) & (g2030) & (!g2062) & (g2085)) + ((!g1892) & (!g1908) & (!g2026) & (g2030) & (g2062) & (!g2085)) + ((!g1892) & (!g1908) & (g2026) & (!g2030) & (!g2062) & (g2085)) + ((!g1892) & (!g1908) & (g2026) & (!g2030) & (g2062) & (!g2085)) + ((!g1892) & (!g1908) & (g2026) & (g2030) & (!g2062) & (!g2085)) + ((!g1892) & (!g1908) & (g2026) & (g2030) & (g2062) & (g2085)) + ((!g1892) & (g1908) & (!g2026) & (!g2030) & (!g2062) & (g2085)) + ((!g1892) & (g1908) & (!g2026) & (!g2030) & (g2062) & (!g2085)) + ((!g1892) & (g1908) & (!g2026) & (g2030) & (!g2062) & (g2085)) + ((!g1892) & (g1908) & (!g2026) & (g2030) & (g2062) & (!g2085)) + ((!g1892) & (g1908) & (g2026) & (!g2030) & (!g2062) & (g2085)) + ((!g1892) & (g1908) & (g2026) & (!g2030) & (g2062) & (!g2085)) + ((!g1892) & (g1908) & (g2026) & (g2030) & (!g2062) & (!g2085)) + ((!g1892) & (g1908) & (g2026) & (g2030) & (g2062) & (g2085)) + ((g1892) & (!g1908) & (!g2026) & (!g2030) & (!g2062) & (g2085)) + ((g1892) & (!g1908) & (!g2026) & (!g2030) & (g2062) & (!g2085)) + ((g1892) & (!g1908) & (!g2026) & (g2030) & (!g2062) & (g2085)) + ((g1892) & (!g1908) & (!g2026) & (g2030) & (g2062) & (!g2085)) + ((g1892) & (!g1908) & (g2026) & (!g2030) & (!g2062) & (g2085)) + ((g1892) & (!g1908) & (g2026) & (!g2030) & (g2062) & (!g2085)) + ((g1892) & (!g1908) & (g2026) & (g2030) & (!g2062) & (!g2085)) + ((g1892) & (!g1908) & (g2026) & (g2030) & (g2062) & (g2085)) + ((g1892) & (g1908) & (!g2026) & (!g2030) & (!g2062) & (g2085)) + ((g1892) & (g1908) & (!g2026) & (!g2030) & (g2062) & (!g2085)) + ((g1892) & (g1908) & (!g2026) & (g2030) & (!g2062) & (!g2085)) + ((g1892) & (g1908) & (!g2026) & (g2030) & (g2062) & (g2085)) + ((g1892) & (g1908) & (g2026) & (!g2030) & (!g2062) & (!g2085)) + ((g1892) & (g1908) & (g2026) & (!g2030) & (g2062) & (g2085)) + ((g1892) & (g1908) & (g2026) & (g2030) & (!g2062) & (!g2085)) + ((g1892) & (g1908) & (g2026) & (g2030) & (g2062) & (g2085)));
	assign g4090 = (((!g1914) & (!g897) & (!g4088) & (g2055) & (!g4089)) + ((!g1914) & (!g897) & (!g4088) & (g2055) & (g4089)) + ((!g1914) & (!g897) & (g4088) & (!g2055) & (!g4089)) + ((!g1914) & (!g897) & (g4088) & (!g2055) & (g4089)) + ((!g1914) & (g897) & (!g4088) & (!g2055) & (!g4089)) + ((!g1914) & (g897) & (!g4088) & (!g2055) & (g4089)) + ((!g1914) & (g897) & (g4088) & (g2055) & (!g4089)) + ((!g1914) & (g897) & (g4088) & (g2055) & (g4089)) + ((g1914) & (!g897) & (!g4088) & (!g2055) & (g4089)) + ((g1914) & (!g897) & (!g4088) & (g2055) & (g4089)) + ((g1914) & (!g897) & (g4088) & (!g2055) & (g4089)) + ((g1914) & (!g897) & (g4088) & (g2055) & (g4089)) + ((g1914) & (g897) & (!g4088) & (!g2055) & (g4089)) + ((g1914) & (g897) & (!g4088) & (g2055) & (g4089)) + ((g1914) & (g897) & (g4088) & (!g2055) & (g4089)) + ((g1914) & (g897) & (g4088) & (g2055) & (g4089)));
	assign g8288 = (((!g5560) & (g5580) & (!g4091)) + ((!g5560) & (g5580) & (g4091)) + ((g5560) & (!g5580) & (g4091)) + ((g5560) & (g5580) & (g4091)));
	assign g4092 = (((!g830) & (!g2003) & (!g4090) & (g4091)) + ((!g830) & (!g2003) & (g4090) & (g4091)) + ((!g830) & (g2003) & (!g4090) & (g4091)) + ((!g830) & (g2003) & (g4090) & (g4091)) + ((g830) & (!g2003) & (g4090) & (!g4091)) + ((g830) & (!g2003) & (g4090) & (g4091)) + ((g830) & (g2003) & (!g4090) & (!g4091)) + ((g830) & (g2003) & (!g4090) & (g4091)));
	assign g4093 = (((!g3465) & (g2123) & (g2127)) + ((g3465) & (!g2123) & (g2127)) + ((g3465) & (g2123) & (!g2127)) + ((g3465) & (g2123) & (g2127)));
	assign g4094 = (((!g2649) & (!g2683) & (g3222) & (g3301) & (!g4078)) + ((!g2649) & (g2683) & (!g3222) & (g3301) & (!g4078)) + ((!g2649) & (g2683) & (!g3222) & (g3301) & (g4078)) + ((!g2649) & (g2683) & (g3222) & (!g3301) & (!g4078)) + ((!g2649) & (g2683) & (g3222) & (g3301) & (!g4078)) + ((!g2649) & (g2683) & (g3222) & (g3301) & (g4078)) + ((g2649) & (!g2683) & (!g3222) & (g3301) & (!g4078)) + ((g2649) & (!g2683) & (g3222) & (g3301) & (!g4078)) + ((g2649) & (!g2683) & (g3222) & (g3301) & (g4078)) + ((g2649) & (g2683) & (!g3222) & (!g3301) & (!g4078)) + ((g2649) & (g2683) & (!g3222) & (g3301) & (!g4078)) + ((g2649) & (g2683) & (!g3222) & (g3301) & (g4078)) + ((g2649) & (g2683) & (g3222) & (!g3301) & (!g4078)) + ((g2649) & (g2683) & (g3222) & (!g3301) & (g4078)) + ((g2649) & (g2683) & (g3222) & (g3301) & (!g4078)) + ((g2649) & (g2683) & (g3222) & (g3301) & (g4078)));
	assign g4095 = (((!g830) & (key[171]) & (!g1914) & (!g4094) & (!g4093) & (!g5682)) + ((!g830) & (key[171]) & (!g1914) & (!g4094) & (!g4093) & (g5682)) + ((!g830) & (key[171]) & (!g1914) & (!g4094) & (g4093) & (!g5682)) + ((!g830) & (key[171]) & (!g1914) & (!g4094) & (g4093) & (g5682)) + ((!g830) & (key[171]) & (!g1914) & (g4094) & (!g4093) & (!g5682)) + ((!g830) & (key[171]) & (!g1914) & (g4094) & (!g4093) & (g5682)) + ((!g830) & (key[171]) & (!g1914) & (g4094) & (g4093) & (!g5682)) + ((!g830) & (key[171]) & (!g1914) & (g4094) & (g4093) & (g5682)) + ((!g830) & (key[171]) & (g1914) & (!g4094) & (!g4093) & (!g5682)) + ((!g830) & (key[171]) & (g1914) & (!g4094) & (!g4093) & (g5682)) + ((!g830) & (key[171]) & (g1914) & (!g4094) & (g4093) & (!g5682)) + ((!g830) & (key[171]) & (g1914) & (!g4094) & (g4093) & (g5682)) + ((!g830) & (key[171]) & (g1914) & (g4094) & (!g4093) & (!g5682)) + ((!g830) & (key[171]) & (g1914) & (g4094) & (!g4093) & (g5682)) + ((!g830) & (key[171]) & (g1914) & (g4094) & (g4093) & (!g5682)) + ((!g830) & (key[171]) & (g1914) & (g4094) & (g4093) & (g5682)) + ((g830) & (!key[171]) & (!g1914) & (!g4094) & (!g4093) & (!g5682)) + ((g830) & (!key[171]) & (!g1914) & (!g4094) & (g4093) & (!g5682)) + ((g830) & (!key[171]) & (!g1914) & (g4094) & (!g4093) & (g5682)) + ((g830) & (!key[171]) & (!g1914) & (g4094) & (g4093) & (g5682)) + ((g830) & (!key[171]) & (g1914) & (!g4094) & (!g4093) & (!g5682)) + ((g830) & (!key[171]) & (g1914) & (!g4094) & (g4093) & (g5682)) + ((g830) & (!key[171]) & (g1914) & (g4094) & (!g4093) & (!g5682)) + ((g830) & (!key[171]) & (g1914) & (g4094) & (g4093) & (g5682)) + ((g830) & (key[171]) & (!g1914) & (!g4094) & (!g4093) & (!g5682)) + ((g830) & (key[171]) & (!g1914) & (!g4094) & (g4093) & (!g5682)) + ((g830) & (key[171]) & (!g1914) & (g4094) & (!g4093) & (g5682)) + ((g830) & (key[171]) & (!g1914) & (g4094) & (g4093) & (g5682)) + ((g830) & (key[171]) & (g1914) & (!g4094) & (!g4093) & (!g5682)) + ((g830) & (key[171]) & (g1914) & (!g4094) & (g4093) & (g5682)) + ((g830) & (key[171]) & (g1914) & (g4094) & (!g4093) & (!g5682)) + ((g830) & (key[171]) & (g1914) & (g4094) & (g4093) & (g5682)));
	assign g4096 = (((!g3392) & (!g2108) & (g2112)) + ((!g3392) & (g2108) & (!g2112)) + ((g3392) & (!g2108) & (!g2112)) + ((g3392) & (g2108) & (g2112)));
	assign g4097 = (((!g931) & (!g3410) & (g2114)) + ((!g931) & (g3410) & (!g2114)) + ((g931) & (!g3410) & (!g2114)) + ((g931) & (g3410) & (g2114)));
	assign g8289 = (((!g5560) & (g5581) & (!g4098)) + ((!g5560) & (g5581) & (g4098)) + ((g5560) & (!g5581) & (g4098)) + ((g5560) & (g5581) & (g4098)));
	assign g4099 = (((!g830) & (!g1914) & (!g2005) & (!g4096) & (!g4097) & (g4098)) + ((!g830) & (!g1914) & (!g2005) & (!g4096) & (g4097) & (g4098)) + ((!g830) & (!g1914) & (!g2005) & (g4096) & (!g4097) & (g4098)) + ((!g830) & (!g1914) & (!g2005) & (g4096) & (g4097) & (g4098)) + ((!g830) & (!g1914) & (g2005) & (!g4096) & (!g4097) & (g4098)) + ((!g830) & (!g1914) & (g2005) & (!g4096) & (g4097) & (g4098)) + ((!g830) & (!g1914) & (g2005) & (g4096) & (!g4097) & (g4098)) + ((!g830) & (!g1914) & (g2005) & (g4096) & (g4097) & (g4098)) + ((!g830) & (g1914) & (!g2005) & (!g4096) & (!g4097) & (g4098)) + ((!g830) & (g1914) & (!g2005) & (!g4096) & (g4097) & (g4098)) + ((!g830) & (g1914) & (!g2005) & (g4096) & (!g4097) & (g4098)) + ((!g830) & (g1914) & (!g2005) & (g4096) & (g4097) & (g4098)) + ((!g830) & (g1914) & (g2005) & (!g4096) & (!g4097) & (g4098)) + ((!g830) & (g1914) & (g2005) & (!g4096) & (g4097) & (g4098)) + ((!g830) & (g1914) & (g2005) & (g4096) & (!g4097) & (g4098)) + ((!g830) & (g1914) & (g2005) & (g4096) & (g4097) & (g4098)) + ((g830) & (!g1914) & (!g2005) & (!g4096) & (g4097) & (!g4098)) + ((g830) & (!g1914) & (!g2005) & (!g4096) & (g4097) & (g4098)) + ((g830) & (!g1914) & (!g2005) & (g4096) & (g4097) & (!g4098)) + ((g830) & (!g1914) & (!g2005) & (g4096) & (g4097) & (g4098)) + ((g830) & (!g1914) & (g2005) & (!g4096) & (!g4097) & (!g4098)) + ((g830) & (!g1914) & (g2005) & (!g4096) & (!g4097) & (g4098)) + ((g830) & (!g1914) & (g2005) & (g4096) & (!g4097) & (!g4098)) + ((g830) & (!g1914) & (g2005) & (g4096) & (!g4097) & (g4098)) + ((g830) & (g1914) & (!g2005) & (g4096) & (!g4097) & (!g4098)) + ((g830) & (g1914) & (!g2005) & (g4096) & (!g4097) & (g4098)) + ((g830) & (g1914) & (!g2005) & (g4096) & (g4097) & (!g4098)) + ((g830) & (g1914) & (!g2005) & (g4096) & (g4097) & (g4098)) + ((g830) & (g1914) & (g2005) & (!g4096) & (!g4097) & (!g4098)) + ((g830) & (g1914) & (g2005) & (!g4096) & (!g4097) & (g4098)) + ((g830) & (g1914) & (g2005) & (!g4096) & (g4097) & (!g4098)) + ((g830) & (g1914) & (g2005) & (!g4096) & (g4097) & (g4098)));
	assign g4100 = (((!g931) & (g3410) & (g2114)) + ((g931) & (!g3410) & (g2114)) + ((g931) & (g3410) & (!g2114)) + ((g931) & (g3410) & (g2114)));
	assign g4101 = (((!g3392) & (g2108) & (g2112)) + ((g3392) & (!g2108) & (g2112)) + ((g3392) & (g2108) & (!g2112)) + ((g3392) & (g2108) & (g2112)));
	assign g4102 = (((!g4101) & (!g2144) & (g2167)) + ((!g4101) & (g2144) & (!g2167)) + ((g4101) & (!g2144) & (!g2167)) + ((g4101) & (g2144) & (g2167)));
	assign g4103 = (((!g1914) & (!g964) & (!g4100) & (g2137) & (!g4102)) + ((!g1914) & (!g964) & (!g4100) & (g2137) & (g4102)) + ((!g1914) & (!g964) & (g4100) & (!g2137) & (!g4102)) + ((!g1914) & (!g964) & (g4100) & (!g2137) & (g4102)) + ((!g1914) & (g964) & (!g4100) & (!g2137) & (!g4102)) + ((!g1914) & (g964) & (!g4100) & (!g2137) & (g4102)) + ((!g1914) & (g964) & (g4100) & (g2137) & (!g4102)) + ((!g1914) & (g964) & (g4100) & (g2137) & (g4102)) + ((g1914) & (!g964) & (!g4100) & (!g2137) & (g4102)) + ((g1914) & (!g964) & (!g4100) & (g2137) & (g4102)) + ((g1914) & (!g964) & (g4100) & (!g2137) & (g4102)) + ((g1914) & (!g964) & (g4100) & (g2137) & (g4102)) + ((g1914) & (g964) & (!g4100) & (!g2137) & (g4102)) + ((g1914) & (g964) & (!g4100) & (g2137) & (g4102)) + ((g1914) & (g964) & (g4100) & (!g2137) & (g4102)) + ((g1914) & (g964) & (g4100) & (g2137) & (g4102)));
	assign g8290 = (((!g5560) & (g5582) & (!g4104)) + ((!g5560) & (g5582) & (g4104)) + ((g5560) & (!g5582) & (g4104)) + ((g5560) & (g5582) & (g4104)));
	assign g4105 = (((!g830) & (!g2011) & (!g4103) & (g4104)) + ((!g830) & (!g2011) & (g4103) & (g4104)) + ((!g830) & (g2011) & (!g4103) & (g4104)) + ((!g830) & (g2011) & (g4103) & (g4104)) + ((g830) & (!g2011) & (g4103) & (!g4104)) + ((g830) & (!g2011) & (g4103) & (g4104)) + ((g830) & (g2011) & (!g4103) & (!g4104)) + ((g830) & (g2011) & (!g4103) & (g4104)));
	assign g4106 = (((!g3467) & (g3468)) + ((g3467) & (!g3468)) + ((g3467) & (g3468)));
	assign g4107 = (((!g1914) & (!g1884) & (g1886) & (!g4106) & (!g2230) & (!g2253)) + ((!g1914) & (!g1884) & (g1886) & (!g4106) & (!g2230) & (g2253)) + ((!g1914) & (!g1884) & (g1886) & (!g4106) & (g2230) & (!g2253)) + ((!g1914) & (!g1884) & (g1886) & (!g4106) & (g2230) & (g2253)) + ((!g1914) & (!g1884) & (g1886) & (g4106) & (!g2230) & (!g2253)) + ((!g1914) & (!g1884) & (g1886) & (g4106) & (!g2230) & (g2253)) + ((!g1914) & (!g1884) & (g1886) & (g4106) & (g2230) & (!g2253)) + ((!g1914) & (!g1884) & (g1886) & (g4106) & (g2230) & (g2253)) + ((!g1914) & (g1884) & (!g1886) & (!g4106) & (!g2230) & (!g2253)) + ((!g1914) & (g1884) & (!g1886) & (!g4106) & (!g2230) & (g2253)) + ((!g1914) & (g1884) & (!g1886) & (!g4106) & (g2230) & (!g2253)) + ((!g1914) & (g1884) & (!g1886) & (!g4106) & (g2230) & (g2253)) + ((!g1914) & (g1884) & (!g1886) & (g4106) & (!g2230) & (!g2253)) + ((!g1914) & (g1884) & (!g1886) & (g4106) & (!g2230) & (g2253)) + ((!g1914) & (g1884) & (!g1886) & (g4106) & (g2230) & (!g2253)) + ((!g1914) & (g1884) & (!g1886) & (g4106) & (g2230) & (g2253)) + ((g1914) & (!g1884) & (!g1886) & (!g4106) & (!g2230) & (g2253)) + ((g1914) & (!g1884) & (!g1886) & (!g4106) & (g2230) & (!g2253)) + ((g1914) & (!g1884) & (!g1886) & (g4106) & (!g2230) & (!g2253)) + ((g1914) & (!g1884) & (!g1886) & (g4106) & (g2230) & (g2253)) + ((g1914) & (!g1884) & (g1886) & (!g4106) & (!g2230) & (g2253)) + ((g1914) & (!g1884) & (g1886) & (!g4106) & (g2230) & (!g2253)) + ((g1914) & (!g1884) & (g1886) & (g4106) & (!g2230) & (!g2253)) + ((g1914) & (!g1884) & (g1886) & (g4106) & (g2230) & (g2253)) + ((g1914) & (g1884) & (!g1886) & (!g4106) & (!g2230) & (g2253)) + ((g1914) & (g1884) & (!g1886) & (!g4106) & (g2230) & (!g2253)) + ((g1914) & (g1884) & (!g1886) & (g4106) & (!g2230) & (!g2253)) + ((g1914) & (g1884) & (!g1886) & (g4106) & (g2230) & (g2253)) + ((g1914) & (g1884) & (g1886) & (!g4106) & (!g2230) & (g2253)) + ((g1914) & (g1884) & (g1886) & (!g4106) & (g2230) & (!g2253)) + ((g1914) & (g1884) & (g1886) & (g4106) & (!g2230) & (!g2253)) + ((g1914) & (g1884) & (g1886) & (g4106) & (g2230) & (g2253)));
	assign g4108 = (((!g830) & (!g2012) & (!g4107) & (key[173])) + ((!g830) & (!g2012) & (g4107) & (key[173])) + ((!g830) & (g2012) & (!g4107) & (key[173])) + ((!g830) & (g2012) & (g4107) & (key[173])) + ((g830) & (!g2012) & (g4107) & (!key[173])) + ((g830) & (!g2012) & (g4107) & (key[173])) + ((g830) & (g2012) & (!g4107) & (!key[173])) + ((g830) & (g2012) & (!g4107) & (key[173])));
	assign g4109 = (((!g4101) & (!g2144) & (!g2167) & (!g2188) & (g2192)) + ((!g4101) & (!g2144) & (!g2167) & (g2188) & (!g2192)) + ((!g4101) & (!g2144) & (g2167) & (!g2188) & (g2192)) + ((!g4101) & (!g2144) & (g2167) & (g2188) & (!g2192)) + ((!g4101) & (g2144) & (!g2167) & (!g2188) & (g2192)) + ((!g4101) & (g2144) & (!g2167) & (g2188) & (!g2192)) + ((!g4101) & (g2144) & (g2167) & (!g2188) & (!g2192)) + ((!g4101) & (g2144) & (g2167) & (g2188) & (g2192)) + ((g4101) & (!g2144) & (!g2167) & (!g2188) & (g2192)) + ((g4101) & (!g2144) & (!g2167) & (g2188) & (!g2192)) + ((g4101) & (!g2144) & (g2167) & (!g2188) & (!g2192)) + ((g4101) & (!g2144) & (g2167) & (g2188) & (g2192)) + ((g4101) & (g2144) & (!g2167) & (!g2188) & (!g2192)) + ((g4101) & (g2144) & (!g2167) & (g2188) & (g2192)) + ((g4101) & (g2144) & (g2167) & (!g2188) & (!g2192)) + ((g4101) & (g2144) & (g2167) & (g2188) & (g2192)));
	assign g8291 = (((!g5560) & (g5584) & (!g4110)) + ((!g5560) & (g5584) & (g4110)) + ((g5560) & (!g5584) & (g4110)) + ((g5560) & (g5584) & (g4110)));
	assign g4111 = (((!g830) & (!g2013) & (!g6905) & (g4110)) + ((!g830) & (!g2013) & (g6905) & (g4110)) + ((!g830) & (g2013) & (!g6905) & (g4110)) + ((!g830) & (g2013) & (g6905) & (g4110)) + ((g830) & (!g2013) & (g6905) & (!g4110)) + ((g830) & (!g2013) & (g6905) & (g4110)) + ((g830) & (g2013) & (!g6905) & (!g4110)) + ((g830) & (g2013) & (!g6905) & (g4110)));
	assign g4112 = (((!g1884) & (!g1977) & (!g1886) & (g2032)) + ((!g1884) & (!g1977) & (g1886) & (g2032)) + ((!g1884) & (g1977) & (!g1886) & (!g2032)) + ((!g1884) & (g1977) & (g1886) & (!g2032)) + ((g1884) & (!g1977) & (!g1886) & (g2032)) + ((g1884) & (!g1977) & (g1886) & (!g2032)) + ((g1884) & (g1977) & (!g1886) & (!g2032)) + ((g1884) & (g1977) & (g1886) & (g2032)));
	assign g4113 = (((!g830) & (!g2014) & (!g6894) & (key[174])) + ((!g830) & (!g2014) & (g6894) & (key[174])) + ((!g830) & (g2014) & (!g6894) & (key[174])) + ((!g830) & (g2014) & (g6894) & (key[174])) + ((g830) & (!g2014) & (g6894) & (!key[174])) + ((g830) & (!g2014) & (g6894) & (key[174])) + ((g830) & (g2014) & (!g6894) & (!key[174])) + ((g830) & (g2014) & (!g6894) & (key[174])));
	assign g4114 = (((!g2516) & (g1677)) + ((g2516) & (!g1677)));
	assign g4115 = (((!g2377) & (!g2424) & (g1610) & (g1644) & (!g3636) & (g4114)) + ((!g2377) & (g2424) & (!g1610) & (g1644) & (!g3636) & (g4114)) + ((!g2377) & (g2424) & (!g1610) & (g1644) & (g3636) & (g4114)) + ((!g2377) & (g2424) & (g1610) & (!g1644) & (!g3636) & (g4114)) + ((!g2377) & (g2424) & (g1610) & (g1644) & (!g3636) & (g4114)) + ((!g2377) & (g2424) & (g1610) & (g1644) & (g3636) & (g4114)) + ((g2377) & (!g2424) & (!g1610) & (g1644) & (!g3636) & (g4114)) + ((g2377) & (!g2424) & (g1610) & (g1644) & (!g3636) & (g4114)) + ((g2377) & (!g2424) & (g1610) & (g1644) & (g3636) & (g4114)) + ((g2377) & (g2424) & (!g1610) & (!g1644) & (!g3636) & (g4114)) + ((g2377) & (g2424) & (!g1610) & (g1644) & (!g3636) & (g4114)) + ((g2377) & (g2424) & (!g1610) & (g1644) & (g3636) & (g4114)) + ((g2377) & (g2424) & (g1610) & (!g1644) & (!g3636) & (g4114)) + ((g2377) & (g2424) & (g1610) & (!g1644) & (g3636) & (g4114)) + ((g2377) & (g2424) & (g1610) & (g1644) & (!g3636) & (g4114)) + ((g2377) & (g2424) & (g1610) & (g1644) & (g3636) & (g4114)));
	assign g4116 = (((g2516) & (g1677)));
	assign g4117 = (((!g2552) & (!g1711) & (!g4115) & (g4116)) + ((!g2552) & (!g1711) & (g4115) & (!g4116)) + ((!g2552) & (!g1711) & (g4115) & (g4116)) + ((!g2552) & (g1711) & (!g4115) & (!g4116)) + ((g2552) & (!g1711) & (!g4115) & (!g4116)) + ((g2552) & (g1711) & (!g4115) & (g4116)) + ((g2552) & (g1711) & (g4115) & (!g4116)) + ((g2552) & (g1711) & (g4115) & (g4116)));
	assign g4118 = (((!g2871) & (!g3651) & (!g2848) & (!g2893) & (g2897)) + ((!g2871) & (!g3651) & (!g2848) & (g2893) & (!g2897)) + ((!g2871) & (!g3651) & (g2848) & (!g2893) & (g2897)) + ((!g2871) & (!g3651) & (g2848) & (g2893) & (!g2897)) + ((!g2871) & (g3651) & (!g2848) & (!g2893) & (g2897)) + ((!g2871) & (g3651) & (!g2848) & (g2893) & (!g2897)) + ((!g2871) & (g3651) & (g2848) & (!g2893) & (!g2897)) + ((!g2871) & (g3651) & (g2848) & (g2893) & (g2897)) + ((g2871) & (!g3651) & (!g2848) & (!g2893) & (g2897)) + ((g2871) & (!g3651) & (!g2848) & (g2893) & (!g2897)) + ((g2871) & (!g3651) & (g2848) & (!g2893) & (!g2897)) + ((g2871) & (!g3651) & (g2848) & (g2893) & (g2897)) + ((g2871) & (g3651) & (!g2848) & (!g2893) & (!g2897)) + ((g2871) & (g3651) & (!g2848) & (g2893) & (g2897)) + ((g2871) & (g3651) & (g2848) & (!g2893) & (!g2897)) + ((g2871) & (g3651) & (g2848) & (g2893) & (g2897)));
	assign g4119 = (((!g830) & (!g1914) & (!g2022) & (!g4117) & (!g4118) & (key[1])) + ((!g830) & (!g1914) & (!g2022) & (!g4117) & (g4118) & (key[1])) + ((!g830) & (!g1914) & (!g2022) & (g4117) & (!g4118) & (key[1])) + ((!g830) & (!g1914) & (!g2022) & (g4117) & (g4118) & (key[1])) + ((!g830) & (!g1914) & (g2022) & (!g4117) & (!g4118) & (key[1])) + ((!g830) & (!g1914) & (g2022) & (!g4117) & (g4118) & (key[1])) + ((!g830) & (!g1914) & (g2022) & (g4117) & (!g4118) & (key[1])) + ((!g830) & (!g1914) & (g2022) & (g4117) & (g4118) & (key[1])) + ((!g830) & (g1914) & (!g2022) & (!g4117) & (!g4118) & (key[1])) + ((!g830) & (g1914) & (!g2022) & (!g4117) & (g4118) & (key[1])) + ((!g830) & (g1914) & (!g2022) & (g4117) & (!g4118) & (key[1])) + ((!g830) & (g1914) & (!g2022) & (g4117) & (g4118) & (key[1])) + ((!g830) & (g1914) & (g2022) & (!g4117) & (!g4118) & (key[1])) + ((!g830) & (g1914) & (g2022) & (!g4117) & (g4118) & (key[1])) + ((!g830) & (g1914) & (g2022) & (g4117) & (!g4118) & (key[1])) + ((!g830) & (g1914) & (g2022) & (g4117) & (g4118) & (key[1])) + ((g830) & (!g1914) & (!g2022) & (!g4117) & (g4118) & (!key[1])) + ((g830) & (!g1914) & (!g2022) & (!g4117) & (g4118) & (key[1])) + ((g830) & (!g1914) & (!g2022) & (g4117) & (g4118) & (!key[1])) + ((g830) & (!g1914) & (!g2022) & (g4117) & (g4118) & (key[1])) + ((g830) & (!g1914) & (g2022) & (!g4117) & (!g4118) & (!key[1])) + ((g830) & (!g1914) & (g2022) & (!g4117) & (!g4118) & (key[1])) + ((g830) & (!g1914) & (g2022) & (g4117) & (!g4118) & (!key[1])) + ((g830) & (!g1914) & (g2022) & (g4117) & (!g4118) & (key[1])) + ((g830) & (g1914) & (!g2022) & (g4117) & (!g4118) & (!key[1])) + ((g830) & (g1914) & (!g2022) & (g4117) & (!g4118) & (key[1])) + ((g830) & (g1914) & (!g2022) & (g4117) & (g4118) & (!key[1])) + ((g830) & (g1914) & (!g2022) & (g4117) & (g4118) & (key[1])) + ((g830) & (g1914) & (g2022) & (!g4117) & (!g4118) & (!key[1])) + ((g830) & (g1914) & (g2022) & (!g4117) & (!g4118) & (key[1])) + ((g830) & (g1914) & (g2022) & (!g4117) & (g4118) & (!key[1])) + ((g830) & (g1914) & (g2022) & (!g4117) & (g4118) & (key[1])));
	assign g4120 = (((!g2013) & (!g2051) & (!g3543) & (!g2626) & (g2659)) + ((!g2013) & (!g2051) & (!g3543) & (g2626) & (g2659)) + ((!g2013) & (!g2051) & (g3543) & (!g2626) & (g2659)) + ((!g2013) & (!g2051) & (g3543) & (g2626) & (!g2659)) + ((!g2013) & (g2051) & (!g3543) & (!g2626) & (!g2659)) + ((!g2013) & (g2051) & (!g3543) & (g2626) & (!g2659)) + ((!g2013) & (g2051) & (g3543) & (!g2626) & (!g2659)) + ((!g2013) & (g2051) & (g3543) & (g2626) & (g2659)) + ((g2013) & (!g2051) & (!g3543) & (!g2626) & (g2659)) + ((g2013) & (!g2051) & (!g3543) & (g2626) & (!g2659)) + ((g2013) & (!g2051) & (g3543) & (!g2626) & (!g2659)) + ((g2013) & (!g2051) & (g3543) & (g2626) & (!g2659)) + ((g2013) & (g2051) & (!g3543) & (!g2626) & (!g2659)) + ((g2013) & (g2051) & (!g3543) & (g2626) & (g2659)) + ((g2013) & (g2051) & (g3543) & (!g2626) & (g2659)) + ((g2013) & (g2051) & (g3543) & (g2626) & (g2659)));
	assign g4121 = (((!g1972) & (!g1975) & (g2578) & (g2617) & (!g3551) & (g3552)) + ((!g1972) & (!g1975) & (g2578) & (g2617) & (g3551) & (!g3552)) + ((!g1972) & (!g1975) & (g2578) & (g2617) & (g3551) & (g3552)) + ((!g1972) & (g1975) & (!g2578) & (g2617) & (!g3551) & (!g3552)) + ((!g1972) & (g1975) & (!g2578) & (g2617) & (!g3551) & (g3552)) + ((!g1972) & (g1975) & (!g2578) & (g2617) & (g3551) & (!g3552)) + ((!g1972) & (g1975) & (!g2578) & (g2617) & (g3551) & (g3552)) + ((!g1972) & (g1975) & (g2578) & (!g2617) & (!g3551) & (g3552)) + ((!g1972) & (g1975) & (g2578) & (!g2617) & (g3551) & (!g3552)) + ((!g1972) & (g1975) & (g2578) & (!g2617) & (g3551) & (g3552)) + ((!g1972) & (g1975) & (g2578) & (g2617) & (!g3551) & (!g3552)) + ((!g1972) & (g1975) & (g2578) & (g2617) & (!g3551) & (g3552)) + ((!g1972) & (g1975) & (g2578) & (g2617) & (g3551) & (!g3552)) + ((!g1972) & (g1975) & (g2578) & (g2617) & (g3551) & (g3552)) + ((g1972) & (!g1975) & (!g2578) & (g2617) & (!g3551) & (g3552)) + ((g1972) & (!g1975) & (!g2578) & (g2617) & (g3551) & (!g3552)) + ((g1972) & (!g1975) & (!g2578) & (g2617) & (g3551) & (g3552)) + ((g1972) & (!g1975) & (g2578) & (g2617) & (!g3551) & (!g3552)) + ((g1972) & (!g1975) & (g2578) & (g2617) & (!g3551) & (g3552)) + ((g1972) & (!g1975) & (g2578) & (g2617) & (g3551) & (!g3552)) + ((g1972) & (!g1975) & (g2578) & (g2617) & (g3551) & (g3552)) + ((g1972) & (g1975) & (!g2578) & (!g2617) & (!g3551) & (g3552)) + ((g1972) & (g1975) & (!g2578) & (!g2617) & (g3551) & (!g3552)) + ((g1972) & (g1975) & (!g2578) & (!g2617) & (g3551) & (g3552)) + ((g1972) & (g1975) & (!g2578) & (g2617) & (!g3551) & (!g3552)) + ((g1972) & (g1975) & (!g2578) & (g2617) & (!g3551) & (g3552)) + ((g1972) & (g1975) & (!g2578) & (g2617) & (g3551) & (!g3552)) + ((g1972) & (g1975) & (!g2578) & (g2617) & (g3551) & (g3552)) + ((g1972) & (g1975) & (g2578) & (!g2617) & (!g3551) & (!g3552)) + ((g1972) & (g1975) & (g2578) & (!g2617) & (!g3551) & (g3552)) + ((g1972) & (g1975) & (g2578) & (!g2617) & (g3551) & (!g3552)) + ((g1972) & (g1975) & (g2578) & (!g2617) & (g3551) & (g3552)) + ((g1972) & (g1975) & (g2578) & (g2617) & (!g3551) & (!g3552)) + ((g1972) & (g1975) & (g2578) & (g2617) & (!g3551) & (g3552)) + ((g1972) & (g1975) & (g2578) & (g2617) & (g3551) & (!g3552)) + ((g1972) & (g1975) & (g2578) & (g2617) & (g3551) & (g3552)));
	assign g4122 = (((!g2212) & (!g2262) & (!g2851) & (g2900) & (!g3667)) + ((!g2212) & (!g2262) & (!g2851) & (g2900) & (g3667)) + ((!g2212) & (!g2262) & (g2851) & (!g2900) & (g3667)) + ((!g2212) & (!g2262) & (g2851) & (g2900) & (!g3667)) + ((!g2212) & (g2262) & (!g2851) & (!g2900) & (!g3667)) + ((!g2212) & (g2262) & (!g2851) & (!g2900) & (g3667)) + ((!g2212) & (g2262) & (g2851) & (!g2900) & (!g3667)) + ((!g2212) & (g2262) & (g2851) & (g2900) & (g3667)) + ((g2212) & (!g2262) & (!g2851) & (!g2900) & (g3667)) + ((g2212) & (!g2262) & (!g2851) & (g2900) & (!g3667)) + ((g2212) & (!g2262) & (g2851) & (!g2900) & (!g3667)) + ((g2212) & (!g2262) & (g2851) & (!g2900) & (g3667)) + ((g2212) & (g2262) & (!g2851) & (!g2900) & (!g3667)) + ((g2212) & (g2262) & (!g2851) & (g2900) & (g3667)) + ((g2212) & (g2262) & (g2851) & (g2900) & (!g3667)) + ((g2212) & (g2262) & (g2851) & (g2900) & (g3667)));
	assign g4123 = (((!g3128) & (g3106)) + ((g3128) & (!g3106)));
	assign g4124 = (((!g3031) & (!g3053) & (g3088) & (!g3684) & (g3084) & (g4123)) + ((!g3031) & (!g3053) & (g3088) & (g3684) & (g3084) & (g4123)) + ((!g3031) & (g3053) & (!g3088) & (!g3684) & (g3084) & (g4123)) + ((!g3031) & (g3053) & (g3088) & (!g3684) & (!g3084) & (g4123)) + ((!g3031) & (g3053) & (g3088) & (!g3684) & (g3084) & (g4123)) + ((!g3031) & (g3053) & (g3088) & (g3684) & (g3084) & (g4123)) + ((g3031) & (!g3053) & (!g3088) & (!g3684) & (g3084) & (g4123)) + ((g3031) & (!g3053) & (g3088) & (!g3684) & (!g3084) & (g4123)) + ((g3031) & (!g3053) & (g3088) & (!g3684) & (g3084) & (g4123)) + ((g3031) & (!g3053) & (g3088) & (g3684) & (g3084) & (g4123)) + ((g3031) & (g3053) & (!g3088) & (!g3684) & (g3084) & (g4123)) + ((g3031) & (g3053) & (!g3088) & (g3684) & (g3084) & (g4123)) + ((g3031) & (g3053) & (g3088) & (!g3684) & (!g3084) & (g4123)) + ((g3031) & (g3053) & (g3088) & (!g3684) & (g3084) & (g4123)) + ((g3031) & (g3053) & (g3088) & (g3684) & (!g3084) & (g4123)) + ((g3031) & (g3053) & (g3088) & (g3684) & (g3084) & (g4123)));
	assign g4125 = (((g3128) & (g3106)));
	assign g4126 = (((!g4124) & (!g4125) & (!g3159) & (g3163)) + ((!g4124) & (!g4125) & (g3159) & (!g3163)) + ((!g4124) & (g4125) & (!g3159) & (!g3163)) + ((!g4124) & (g4125) & (g3159) & (g3163)) + ((g4124) & (!g4125) & (!g3159) & (!g3163)) + ((g4124) & (!g4125) & (g3159) & (g3163)) + ((g4124) & (g4125) & (!g3159) & (!g3163)) + ((g4124) & (g4125) & (g3159) & (g3163)));
	assign g8292 = (((!g5560) & (g5585) & (!g4127)) + ((!g5560) & (g5585) & (g4127)) + ((g5560) & (!g5585) & (g4127)) + ((g5560) & (g5585) & (g4127)));
	assign g4128 = (((!g830) & (!g1914) & (!g2028) & (!g4122) & (!g4126) & (g4127)) + ((!g830) & (!g1914) & (!g2028) & (!g4122) & (g4126) & (g4127)) + ((!g830) & (!g1914) & (!g2028) & (g4122) & (!g4126) & (g4127)) + ((!g830) & (!g1914) & (!g2028) & (g4122) & (g4126) & (g4127)) + ((!g830) & (!g1914) & (g2028) & (!g4122) & (!g4126) & (g4127)) + ((!g830) & (!g1914) & (g2028) & (!g4122) & (g4126) & (g4127)) + ((!g830) & (!g1914) & (g2028) & (g4122) & (!g4126) & (g4127)) + ((!g830) & (!g1914) & (g2028) & (g4122) & (g4126) & (g4127)) + ((!g830) & (g1914) & (!g2028) & (!g4122) & (!g4126) & (g4127)) + ((!g830) & (g1914) & (!g2028) & (!g4122) & (g4126) & (g4127)) + ((!g830) & (g1914) & (!g2028) & (g4122) & (!g4126) & (g4127)) + ((!g830) & (g1914) & (!g2028) & (g4122) & (g4126) & (g4127)) + ((!g830) & (g1914) & (g2028) & (!g4122) & (!g4126) & (g4127)) + ((!g830) & (g1914) & (g2028) & (!g4122) & (g4126) & (g4127)) + ((!g830) & (g1914) & (g2028) & (g4122) & (!g4126) & (g4127)) + ((!g830) & (g1914) & (g2028) & (g4122) & (g4126) & (g4127)) + ((g830) & (!g1914) & (!g2028) & (!g4122) & (g4126) & (!g4127)) + ((g830) & (!g1914) & (!g2028) & (!g4122) & (g4126) & (g4127)) + ((g830) & (!g1914) & (!g2028) & (g4122) & (g4126) & (!g4127)) + ((g830) & (!g1914) & (!g2028) & (g4122) & (g4126) & (g4127)) + ((g830) & (!g1914) & (g2028) & (!g4122) & (!g4126) & (!g4127)) + ((g830) & (!g1914) & (g2028) & (!g4122) & (!g4126) & (g4127)) + ((g830) & (!g1914) & (g2028) & (g4122) & (!g4126) & (!g4127)) + ((g830) & (!g1914) & (g2028) & (g4122) & (!g4126) & (g4127)) + ((g830) & (g1914) & (!g2028) & (g4122) & (!g4126) & (!g4127)) + ((g830) & (g1914) & (!g2028) & (g4122) & (!g4126) & (g4127)) + ((g830) & (g1914) & (!g2028) & (g4122) & (g4126) & (!g4127)) + ((g830) & (g1914) & (!g2028) & (g4122) & (g4126) & (g4127)) + ((g830) & (g1914) & (g2028) & (!g4122) & (!g4126) & (!g4127)) + ((g830) & (g1914) & (g2028) & (!g4122) & (!g4126) & (g4127)) + ((g830) & (g1914) & (g2028) & (!g4122) & (g4126) & (!g4127)) + ((g830) & (g1914) & (g2028) & (!g4122) & (g4126) & (g4127)));
	assign g4129 = (((!g3113) & (g3116)) + ((g3113) & (!g3116)));
	assign g4130 = (((!g3038) & (!g3078) & (g3041) & (!g3793) & (g3086) & (g4129)) + ((!g3038) & (g3078) & (!g3041) & (!g3793) & (g3086) & (g4129)) + ((!g3038) & (g3078) & (!g3041) & (g3793) & (g3086) & (g4129)) + ((!g3038) & (g3078) & (g3041) & (!g3793) & (!g3086) & (g4129)) + ((!g3038) & (g3078) & (g3041) & (!g3793) & (g3086) & (g4129)) + ((!g3038) & (g3078) & (g3041) & (g3793) & (g3086) & (g4129)) + ((g3038) & (!g3078) & (!g3041) & (!g3793) & (g3086) & (g4129)) + ((g3038) & (!g3078) & (g3041) & (!g3793) & (g3086) & (g4129)) + ((g3038) & (!g3078) & (g3041) & (g3793) & (g3086) & (g4129)) + ((g3038) & (g3078) & (!g3041) & (!g3793) & (!g3086) & (g4129)) + ((g3038) & (g3078) & (!g3041) & (!g3793) & (g3086) & (g4129)) + ((g3038) & (g3078) & (!g3041) & (g3793) & (g3086) & (g4129)) + ((g3038) & (g3078) & (g3041) & (!g3793) & (!g3086) & (g4129)) + ((g3038) & (g3078) & (g3041) & (!g3793) & (g3086) & (g4129)) + ((g3038) & (g3078) & (g3041) & (g3793) & (!g3086) & (g4129)) + ((g3038) & (g3078) & (g3041) & (g3793) & (g3086) & (g4129)));
	assign g4131 = (((g3113) & (g3116)));
	assign g4132 = (((!g4130) & (!g4131) & (!g3153) & (g3161)) + ((!g4130) & (!g4131) & (g3153) & (!g3161)) + ((!g4130) & (g4131) & (!g3153) & (!g3161)) + ((!g4130) & (g4131) & (g3153) & (g3161)) + ((g4130) & (!g4131) & (!g3153) & (!g3161)) + ((g4130) & (!g4131) & (g3153) & (g3161)) + ((g4130) & (g4131) & (!g3153) & (!g3161)) + ((g4130) & (g4131) & (g3153) & (g3161)));
	assign g4133 = (((!g2211) & (!g2257) & (!g2863) & (!g3808) & (g2902)) + ((!g2211) & (!g2257) & (!g2863) & (g3808) & (g2902)) + ((!g2211) & (!g2257) & (g2863) & (!g3808) & (g2902)) + ((!g2211) & (!g2257) & (g2863) & (g3808) & (!g2902)) + ((!g2211) & (g2257) & (!g2863) & (!g3808) & (!g2902)) + ((!g2211) & (g2257) & (!g2863) & (g3808) & (!g2902)) + ((!g2211) & (g2257) & (g2863) & (!g3808) & (!g2902)) + ((!g2211) & (g2257) & (g2863) & (g3808) & (g2902)) + ((g2211) & (!g2257) & (!g2863) & (!g3808) & (g2902)) + ((g2211) & (!g2257) & (!g2863) & (g3808) & (!g2902)) + ((g2211) & (!g2257) & (g2863) & (!g3808) & (!g2902)) + ((g2211) & (!g2257) & (g2863) & (g3808) & (!g2902)) + ((g2211) & (g2257) & (!g2863) & (!g3808) & (!g2902)) + ((g2211) & (g2257) & (!g2863) & (g3808) & (g2902)) + ((g2211) & (g2257) & (g2863) & (!g3808) & (g2902)) + ((g2211) & (g2257) & (g2863) & (g3808) & (g2902)));
	assign g4134 = (((!g830) & (!g1914) & (!g2030) & (!g4132) & (!g4133) & (key[129])) + ((!g830) & (!g1914) & (!g2030) & (!g4132) & (g4133) & (key[129])) + ((!g830) & (!g1914) & (!g2030) & (g4132) & (!g4133) & (key[129])) + ((!g830) & (!g1914) & (!g2030) & (g4132) & (g4133) & (key[129])) + ((!g830) & (!g1914) & (g2030) & (!g4132) & (!g4133) & (key[129])) + ((!g830) & (!g1914) & (g2030) & (!g4132) & (g4133) & (key[129])) + ((!g830) & (!g1914) & (g2030) & (g4132) & (!g4133) & (key[129])) + ((!g830) & (!g1914) & (g2030) & (g4132) & (g4133) & (key[129])) + ((!g830) & (g1914) & (!g2030) & (!g4132) & (!g4133) & (key[129])) + ((!g830) & (g1914) & (!g2030) & (!g4132) & (g4133) & (key[129])) + ((!g830) & (g1914) & (!g2030) & (g4132) & (!g4133) & (key[129])) + ((!g830) & (g1914) & (!g2030) & (g4132) & (g4133) & (key[129])) + ((!g830) & (g1914) & (g2030) & (!g4132) & (!g4133) & (key[129])) + ((!g830) & (g1914) & (g2030) & (!g4132) & (g4133) & (key[129])) + ((!g830) & (g1914) & (g2030) & (g4132) & (!g4133) & (key[129])) + ((!g830) & (g1914) & (g2030) & (g4132) & (g4133) & (key[129])) + ((g830) & (!g1914) & (!g2030) & (!g4132) & (g4133) & (!key[129])) + ((g830) & (!g1914) & (!g2030) & (!g4132) & (g4133) & (key[129])) + ((g830) & (!g1914) & (!g2030) & (g4132) & (g4133) & (!key[129])) + ((g830) & (!g1914) & (!g2030) & (g4132) & (g4133) & (key[129])) + ((g830) & (!g1914) & (g2030) & (!g4132) & (!g4133) & (!key[129])) + ((g830) & (!g1914) & (g2030) & (!g4132) & (!g4133) & (key[129])) + ((g830) & (!g1914) & (g2030) & (g4132) & (!g4133) & (!key[129])) + ((g830) & (!g1914) & (g2030) & (g4132) & (!g4133) & (key[129])) + ((g830) & (g1914) & (!g2030) & (g4132) & (!g4133) & (!key[129])) + ((g830) & (g1914) & (!g2030) & (g4132) & (!g4133) & (key[129])) + ((g830) & (g1914) & (!g2030) & (g4132) & (g4133) & (!key[129])) + ((g830) & (g1914) & (!g2030) & (g4132) & (g4133) & (key[129])) + ((g830) & (g1914) & (g2030) & (!g4132) & (!g4133) & (!key[129])) + ((g830) & (g1914) & (g2030) & (!g4132) & (!g4133) & (key[129])) + ((g830) & (g1914) & (g2030) & (!g4132) & (g4133) & (!key[129])) + ((g830) & (g1914) & (g2030) & (!g4132) & (g4133) & (key[129])));
	assign g4135 = (((!g3443) & (!g2857) & (!g2863) & (!g2887) & (g2902)) + ((!g3443) & (!g2857) & (!g2863) & (g2887) & (!g2902)) + ((!g3443) & (!g2857) & (g2863) & (!g2887) & (g2902)) + ((!g3443) & (!g2857) & (g2863) & (g2887) & (!g2902)) + ((!g3443) & (g2857) & (!g2863) & (!g2887) & (g2902)) + ((!g3443) & (g2857) & (!g2863) & (g2887) & (!g2902)) + ((!g3443) & (g2857) & (g2863) & (!g2887) & (!g2902)) + ((!g3443) & (g2857) & (g2863) & (g2887) & (g2902)) + ((g3443) & (!g2857) & (!g2863) & (!g2887) & (g2902)) + ((g3443) & (!g2857) & (!g2863) & (g2887) & (!g2902)) + ((g3443) & (!g2857) & (g2863) & (!g2887) & (!g2902)) + ((g3443) & (!g2857) & (g2863) & (g2887) & (g2902)) + ((g3443) & (g2857) & (!g2863) & (!g2887) & (!g2902)) + ((g3443) & (g2857) & (!g2863) & (g2887) & (g2902)) + ((g3443) & (g2857) & (g2863) & (!g2887) & (!g2902)) + ((g3443) & (g2857) & (g2863) & (g2887) & (g2902)));
	assign g4136 = (((!g2519) & (g1677)) + ((g2519) & (!g1677)));
	assign g4137 = (((!g2379) & (!g2427) & (g1610) & (g1644) & (!g3459) & (g4136)) + ((!g2379) & (g2427) & (!g1610) & (g1644) & (!g3459) & (g4136)) + ((!g2379) & (g2427) & (!g1610) & (g1644) & (g3459) & (g4136)) + ((!g2379) & (g2427) & (g1610) & (!g1644) & (!g3459) & (g4136)) + ((!g2379) & (g2427) & (g1610) & (g1644) & (!g3459) & (g4136)) + ((!g2379) & (g2427) & (g1610) & (g1644) & (g3459) & (g4136)) + ((g2379) & (!g2427) & (!g1610) & (g1644) & (!g3459) & (g4136)) + ((g2379) & (!g2427) & (g1610) & (g1644) & (!g3459) & (g4136)) + ((g2379) & (!g2427) & (g1610) & (g1644) & (g3459) & (g4136)) + ((g2379) & (g2427) & (!g1610) & (!g1644) & (!g3459) & (g4136)) + ((g2379) & (g2427) & (!g1610) & (g1644) & (!g3459) & (g4136)) + ((g2379) & (g2427) & (!g1610) & (g1644) & (g3459) & (g4136)) + ((g2379) & (g2427) & (g1610) & (!g1644) & (!g3459) & (g4136)) + ((g2379) & (g2427) & (g1610) & (!g1644) & (g3459) & (g4136)) + ((g2379) & (g2427) & (g1610) & (g1644) & (!g3459) & (g4136)) + ((g2379) & (g2427) & (g1610) & (g1644) & (g3459) & (g4136)));
	assign g4138 = (((g2519) & (g1677)));
	assign g4139 = (((!g2556) & (!g1711) & (!g4137) & (g4138)) + ((!g2556) & (!g1711) & (g4137) & (!g4138)) + ((!g2556) & (!g1711) & (g4137) & (g4138)) + ((!g2556) & (g1711) & (!g4137) & (!g4138)) + ((g2556) & (!g1711) & (!g4137) & (!g4138)) + ((g2556) & (g1711) & (!g4137) & (g4138)) + ((g2556) & (g1711) & (g4137) & (!g4138)) + ((g2556) & (g1711) & (g4137) & (g4138)));
	assign g4140 = (((!g830) & (!g1914) & (!g2032) & (!g4135) & (!g4139) & (key[97])) + ((!g830) & (!g1914) & (!g2032) & (!g4135) & (g4139) & (key[97])) + ((!g830) & (!g1914) & (!g2032) & (g4135) & (!g4139) & (key[97])) + ((!g830) & (!g1914) & (!g2032) & (g4135) & (g4139) & (key[97])) + ((!g830) & (!g1914) & (g2032) & (!g4135) & (!g4139) & (key[97])) + ((!g830) & (!g1914) & (g2032) & (!g4135) & (g4139) & (key[97])) + ((!g830) & (!g1914) & (g2032) & (g4135) & (!g4139) & (key[97])) + ((!g830) & (!g1914) & (g2032) & (g4135) & (g4139) & (key[97])) + ((!g830) & (g1914) & (!g2032) & (!g4135) & (!g4139) & (key[97])) + ((!g830) & (g1914) & (!g2032) & (!g4135) & (g4139) & (key[97])) + ((!g830) & (g1914) & (!g2032) & (g4135) & (!g4139) & (key[97])) + ((!g830) & (g1914) & (!g2032) & (g4135) & (g4139) & (key[97])) + ((!g830) & (g1914) & (g2032) & (!g4135) & (!g4139) & (key[97])) + ((!g830) & (g1914) & (g2032) & (!g4135) & (g4139) & (key[97])) + ((!g830) & (g1914) & (g2032) & (g4135) & (!g4139) & (key[97])) + ((!g830) & (g1914) & (g2032) & (g4135) & (g4139) & (key[97])) + ((g830) & (!g1914) & (!g2032) & (!g4135) & (g4139) & (!key[97])) + ((g830) & (!g1914) & (!g2032) & (!g4135) & (g4139) & (key[97])) + ((g830) & (!g1914) & (!g2032) & (g4135) & (g4139) & (!key[97])) + ((g830) & (!g1914) & (!g2032) & (g4135) & (g4139) & (key[97])) + ((g830) & (!g1914) & (g2032) & (!g4135) & (!g4139) & (!key[97])) + ((g830) & (!g1914) & (g2032) & (!g4135) & (!g4139) & (key[97])) + ((g830) & (!g1914) & (g2032) & (g4135) & (!g4139) & (!key[97])) + ((g830) & (!g1914) & (g2032) & (g4135) & (!g4139) & (key[97])) + ((g830) & (g1914) & (!g2032) & (g4135) & (!g4139) & (!key[97])) + ((g830) & (g1914) & (!g2032) & (g4135) & (!g4139) & (key[97])) + ((g830) & (g1914) & (!g2032) & (g4135) & (g4139) & (!key[97])) + ((g830) & (g1914) & (!g2032) & (g4135) & (g4139) & (key[97])) + ((g830) & (g1914) & (g2032) & (!g4135) & (!g4139) & (!key[97])) + ((g830) & (g1914) & (g2032) & (!g4135) & (!g4139) & (key[97])) + ((g830) & (g1914) & (g2032) & (!g4135) & (g4139) & (!key[97])) + ((g830) & (g1914) & (g2032) & (!g4135) & (g4139) & (key[97])));
	assign g4141 = (((!g3122) & (g3128)) + ((g3122) & (!g3128)));
	assign g4142 = (((!g3047) & (!g3570) & (!g3053) & (g3074) & (g3088) & (g4141)) + ((!g3047) & (!g3570) & (g3053) & (!g3074) & (g3088) & (g4141)) + ((!g3047) & (!g3570) & (g3053) & (g3074) & (!g3088) & (g4141)) + ((!g3047) & (!g3570) & (g3053) & (g3074) & (g3088) & (g4141)) + ((!g3047) & (g3570) & (!g3053) & (g3074) & (g3088) & (g4141)) + ((!g3047) & (g3570) & (g3053) & (g3074) & (g3088) & (g4141)) + ((g3047) & (!g3570) & (!g3053) & (!g3074) & (g3088) & (g4141)) + ((g3047) & (!g3570) & (!g3053) & (g3074) & (!g3088) & (g4141)) + ((g3047) & (!g3570) & (!g3053) & (g3074) & (g3088) & (g4141)) + ((g3047) & (!g3570) & (g3053) & (!g3074) & (g3088) & (g4141)) + ((g3047) & (!g3570) & (g3053) & (g3074) & (!g3088) & (g4141)) + ((g3047) & (!g3570) & (g3053) & (g3074) & (g3088) & (g4141)) + ((g3047) & (g3570) & (!g3053) & (g3074) & (g3088) & (g4141)) + ((g3047) & (g3570) & (g3053) & (!g3074) & (g3088) & (g4141)) + ((g3047) & (g3570) & (g3053) & (g3074) & (!g3088) & (g4141)) + ((g3047) & (g3570) & (g3053) & (g3074) & (g3088) & (g4141)));
	assign g4143 = (((g3122) & (g3128)));
	assign g4144 = (((!g3163) & (!g4142) & (!g4143) & (g3149)) + ((!g3163) & (!g4142) & (g4143) & (!g3149)) + ((!g3163) & (g4142) & (!g4143) & (!g3149)) + ((!g3163) & (g4142) & (g4143) & (!g3149)) + ((g3163) & (!g4142) & (!g4143) & (!g3149)) + ((g3163) & (!g4142) & (g4143) & (g3149)) + ((g3163) & (g4142) & (!g4143) & (g3149)) + ((g3163) & (g4142) & (g4143) & (g3149)));
	assign g4145 = (((!g2210) & (!g2256) & (!g2868) & (g2889) & (!g3585)) + ((!g2210) & (!g2256) & (!g2868) & (g2889) & (g3585)) + ((!g2210) & (!g2256) & (g2868) & (!g2889) & (g3585)) + ((!g2210) & (!g2256) & (g2868) & (g2889) & (!g3585)) + ((!g2210) & (g2256) & (!g2868) & (!g2889) & (!g3585)) + ((!g2210) & (g2256) & (!g2868) & (!g2889) & (g3585)) + ((!g2210) & (g2256) & (g2868) & (!g2889) & (!g3585)) + ((!g2210) & (g2256) & (g2868) & (g2889) & (g3585)) + ((g2210) & (!g2256) & (!g2868) & (!g2889) & (g3585)) + ((g2210) & (!g2256) & (!g2868) & (g2889) & (!g3585)) + ((g2210) & (!g2256) & (g2868) & (!g2889) & (!g3585)) + ((g2210) & (!g2256) & (g2868) & (!g2889) & (g3585)) + ((g2210) & (g2256) & (!g2868) & (!g2889) & (!g3585)) + ((g2210) & (g2256) & (!g2868) & (g2889) & (g3585)) + ((g2210) & (g2256) & (g2868) & (g2889) & (!g3585)) + ((g2210) & (g2256) & (g2868) & (g2889) & (g3585)));
	assign g4146 = (((!g830) & (!g1914) & (!g2034) & (!g4144) & (!g4145) & (nonce[1])) + ((!g830) & (!g1914) & (!g2034) & (!g4144) & (g4145) & (nonce[1])) + ((!g830) & (!g1914) & (!g2034) & (g4144) & (!g4145) & (nonce[1])) + ((!g830) & (!g1914) & (!g2034) & (g4144) & (g4145) & (nonce[1])) + ((!g830) & (!g1914) & (g2034) & (!g4144) & (!g4145) & (nonce[1])) + ((!g830) & (!g1914) & (g2034) & (!g4144) & (g4145) & (nonce[1])) + ((!g830) & (!g1914) & (g2034) & (g4144) & (!g4145) & (nonce[1])) + ((!g830) & (!g1914) & (g2034) & (g4144) & (g4145) & (nonce[1])) + ((!g830) & (g1914) & (!g2034) & (!g4144) & (!g4145) & (nonce[1])) + ((!g830) & (g1914) & (!g2034) & (!g4144) & (g4145) & (nonce[1])) + ((!g830) & (g1914) & (!g2034) & (g4144) & (!g4145) & (nonce[1])) + ((!g830) & (g1914) & (!g2034) & (g4144) & (g4145) & (nonce[1])) + ((!g830) & (g1914) & (g2034) & (!g4144) & (!g4145) & (nonce[1])) + ((!g830) & (g1914) & (g2034) & (!g4144) & (g4145) & (nonce[1])) + ((!g830) & (g1914) & (g2034) & (g4144) & (!g4145) & (nonce[1])) + ((!g830) & (g1914) & (g2034) & (g4144) & (g4145) & (nonce[1])) + ((g830) & (!g1914) & (!g2034) & (!g4144) & (g4145) & (!nonce[1])) + ((g830) & (!g1914) & (!g2034) & (!g4144) & (g4145) & (nonce[1])) + ((g830) & (!g1914) & (!g2034) & (g4144) & (g4145) & (!nonce[1])) + ((g830) & (!g1914) & (!g2034) & (g4144) & (g4145) & (nonce[1])) + ((g830) & (!g1914) & (g2034) & (!g4144) & (!g4145) & (!nonce[1])) + ((g830) & (!g1914) & (g2034) & (!g4144) & (!g4145) & (nonce[1])) + ((g830) & (!g1914) & (g2034) & (g4144) & (!g4145) & (!nonce[1])) + ((g830) & (!g1914) & (g2034) & (g4144) & (!g4145) & (nonce[1])) + ((g830) & (g1914) & (!g2034) & (g4144) & (!g4145) & (!nonce[1])) + ((g830) & (g1914) & (!g2034) & (g4144) & (!g4145) & (nonce[1])) + ((g830) & (g1914) & (!g2034) & (g4144) & (g4145) & (!nonce[1])) + ((g830) & (g1914) & (!g2034) & (g4144) & (g4145) & (nonce[1])) + ((g830) & (g1914) & (g2034) & (!g4144) & (!g4145) & (!nonce[1])) + ((g830) & (g1914) & (g2034) & (!g4144) & (!g4145) & (nonce[1])) + ((g830) & (g1914) & (g2034) & (!g4144) & (g4145) & (!nonce[1])) + ((g830) & (g1914) & (g2034) & (!g4144) & (g4145) & (nonce[1])));
	assign g4147 = (((!g2607) & (!g2663) & (!g2640) & (g2669) & (!g3698)) + ((!g2607) & (!g2663) & (!g2640) & (g2669) & (g3698)) + ((!g2607) & (!g2663) & (g2640) & (!g2669) & (g3698)) + ((!g2607) & (!g2663) & (g2640) & (g2669) & (!g3698)) + ((!g2607) & (g2663) & (!g2640) & (!g2669) & (!g3698)) + ((!g2607) & (g2663) & (!g2640) & (!g2669) & (g3698)) + ((!g2607) & (g2663) & (g2640) & (!g2669) & (!g3698)) + ((!g2607) & (g2663) & (g2640) & (g2669) & (g3698)) + ((g2607) & (!g2663) & (!g2640) & (!g2669) & (g3698)) + ((g2607) & (!g2663) & (!g2640) & (g2669) & (!g3698)) + ((g2607) & (!g2663) & (g2640) & (!g2669) & (!g3698)) + ((g2607) & (!g2663) & (g2640) & (!g2669) & (g3698)) + ((g2607) & (g2663) & (!g2640) & (!g2669) & (!g3698)) + ((g2607) & (g2663) & (!g2640) & (g2669) & (g3698)) + ((g2607) & (g2663) & (g2640) & (g2669) & (!g3698)) + ((g2607) & (g2663) & (g2640) & (g2669) & (g3698)));
	assign g4148 = (((!g2559) & (!g2623) & (g2592) & (g2632) & (!g3706) & (g3707)) + ((!g2559) & (!g2623) & (g2592) & (g2632) & (g3706) & (!g3707)) + ((!g2559) & (!g2623) & (g2592) & (g2632) & (g3706) & (g3707)) + ((!g2559) & (g2623) & (!g2592) & (g2632) & (!g3706) & (!g3707)) + ((!g2559) & (g2623) & (!g2592) & (g2632) & (!g3706) & (g3707)) + ((!g2559) & (g2623) & (!g2592) & (g2632) & (g3706) & (!g3707)) + ((!g2559) & (g2623) & (!g2592) & (g2632) & (g3706) & (g3707)) + ((!g2559) & (g2623) & (g2592) & (!g2632) & (!g3706) & (g3707)) + ((!g2559) & (g2623) & (g2592) & (!g2632) & (g3706) & (!g3707)) + ((!g2559) & (g2623) & (g2592) & (!g2632) & (g3706) & (g3707)) + ((!g2559) & (g2623) & (g2592) & (g2632) & (!g3706) & (!g3707)) + ((!g2559) & (g2623) & (g2592) & (g2632) & (!g3706) & (g3707)) + ((!g2559) & (g2623) & (g2592) & (g2632) & (g3706) & (!g3707)) + ((!g2559) & (g2623) & (g2592) & (g2632) & (g3706) & (g3707)) + ((g2559) & (!g2623) & (!g2592) & (g2632) & (!g3706) & (g3707)) + ((g2559) & (!g2623) & (!g2592) & (g2632) & (g3706) & (!g3707)) + ((g2559) & (!g2623) & (!g2592) & (g2632) & (g3706) & (g3707)) + ((g2559) & (!g2623) & (g2592) & (g2632) & (!g3706) & (!g3707)) + ((g2559) & (!g2623) & (g2592) & (g2632) & (!g3706) & (g3707)) + ((g2559) & (!g2623) & (g2592) & (g2632) & (g3706) & (!g3707)) + ((g2559) & (!g2623) & (g2592) & (g2632) & (g3706) & (g3707)) + ((g2559) & (g2623) & (!g2592) & (!g2632) & (!g3706) & (g3707)) + ((g2559) & (g2623) & (!g2592) & (!g2632) & (g3706) & (!g3707)) + ((g2559) & (g2623) & (!g2592) & (!g2632) & (g3706) & (g3707)) + ((g2559) & (g2623) & (!g2592) & (g2632) & (!g3706) & (!g3707)) + ((g2559) & (g2623) & (!g2592) & (g2632) & (!g3706) & (g3707)) + ((g2559) & (g2623) & (!g2592) & (g2632) & (g3706) & (!g3707)) + ((g2559) & (g2623) & (!g2592) & (g2632) & (g3706) & (g3707)) + ((g2559) & (g2623) & (g2592) & (!g2632) & (!g3706) & (!g3707)) + ((g2559) & (g2623) & (g2592) & (!g2632) & (!g3706) & (g3707)) + ((g2559) & (g2623) & (g2592) & (!g2632) & (g3706) & (!g3707)) + ((g2559) & (g2623) & (g2592) & (!g2632) & (g3706) & (g3707)) + ((g2559) & (g2623) & (g2592) & (g2632) & (!g3706) & (!g3707)) + ((g2559) & (g2623) & (g2592) & (g2632) & (!g3706) & (g3707)) + ((g2559) & (g2623) & (g2592) & (g2632) & (g3706) & (!g3707)) + ((g2559) & (g2623) & (g2592) & (g2632) & (g3706) & (g3707)));
	assign g4149 = (((!g3053) & (g3050) & (!g3826)) + ((g3053) & (!g3050) & (!g3826)) + ((g3053) & (g3050) & (!g3826)) + ((g3053) & (g3050) & (g3826)));
	assign g4150 = (((g1914) & (!g3088) & (!g3080) & (g4149)) + ((g1914) & (!g3088) & (g3080) & (!g4149)) + ((g1914) & (g3088) & (!g3080) & (!g4149)) + ((g1914) & (g3088) & (g3080) & (g4149)));
	assign g4151 = (((!g2377) & (g3067) & (!g3843)) + ((g2377) & (!g3067) & (!g3843)) + ((g2377) & (g3067) & (!g3843)) + ((g2377) & (g3067) & (g3843)));
	assign g4152 = (((!g1914) & (!g2424) & (!g3097) & (g4151)) + ((!g1914) & (!g2424) & (g3097) & (!g4151)) + ((!g1914) & (g2424) & (!g3097) & (!g4151)) + ((!g1914) & (g2424) & (g3097) & (g4151)));
	assign g4153 = (((!g830) & (!g2038) & (!g4150) & (!g4152) & (nonce[33])) + ((!g830) & (!g2038) & (!g4150) & (g4152) & (nonce[33])) + ((!g830) & (!g2038) & (g4150) & (!g4152) & (nonce[33])) + ((!g830) & (!g2038) & (g4150) & (g4152) & (nonce[33])) + ((!g830) & (g2038) & (!g4150) & (!g4152) & (nonce[33])) + ((!g830) & (g2038) & (!g4150) & (g4152) & (nonce[33])) + ((!g830) & (g2038) & (g4150) & (!g4152) & (nonce[33])) + ((!g830) & (g2038) & (g4150) & (g4152) & (nonce[33])) + ((g830) & (!g2038) & (!g4150) & (g4152) & (!nonce[33])) + ((g830) & (!g2038) & (!g4150) & (g4152) & (nonce[33])) + ((g830) & (!g2038) & (g4150) & (!g4152) & (!nonce[33])) + ((g830) & (!g2038) & (g4150) & (!g4152) & (nonce[33])) + ((g830) & (!g2038) & (g4150) & (g4152) & (!nonce[33])) + ((g830) & (!g2038) & (g4150) & (g4152) & (nonce[33])) + ((g830) & (g2038) & (!g4150) & (!g4152) & (!nonce[33])) + ((g830) & (g2038) & (!g4150) & (!g4152) & (nonce[33])));
	assign g4154 = (((!g2213) & (!g2263) & (!g3601) & (!g2871) & (g2897)) + ((!g2213) & (!g2263) & (!g3601) & (g2871) & (g2897)) + ((!g2213) & (!g2263) & (g3601) & (!g2871) & (g2897)) + ((!g2213) & (!g2263) & (g3601) & (g2871) & (!g2897)) + ((!g2213) & (g2263) & (!g3601) & (!g2871) & (!g2897)) + ((!g2213) & (g2263) & (!g3601) & (g2871) & (!g2897)) + ((!g2213) & (g2263) & (g3601) & (!g2871) & (!g2897)) + ((!g2213) & (g2263) & (g3601) & (g2871) & (g2897)) + ((g2213) & (!g2263) & (!g3601) & (!g2871) & (g2897)) + ((g2213) & (!g2263) & (!g3601) & (g2871) & (!g2897)) + ((g2213) & (!g2263) & (g3601) & (!g2871) & (!g2897)) + ((g2213) & (!g2263) & (g3601) & (g2871) & (!g2897)) + ((g2213) & (g2263) & (!g3601) & (!g2871) & (!g2897)) + ((g2213) & (g2263) & (!g3601) & (g2871) & (g2897)) + ((g2213) & (g2263) & (g3601) & (!g2871) & (g2897)) + ((g2213) & (g2263) & (g3601) & (g2871) & (g2897)));
	assign g4155 = (((!g3113) & (g3125)) + ((g3113) & (!g3125)));
	assign g4156 = (((!g3038) & (!g3617) & (!g3050) & (g3078) & (g3080) & (g4155)) + ((!g3038) & (!g3617) & (g3050) & (!g3078) & (g3080) & (g4155)) + ((!g3038) & (!g3617) & (g3050) & (g3078) & (!g3080) & (g4155)) + ((!g3038) & (!g3617) & (g3050) & (g3078) & (g3080) & (g4155)) + ((!g3038) & (g3617) & (!g3050) & (g3078) & (g3080) & (g4155)) + ((!g3038) & (g3617) & (g3050) & (g3078) & (g3080) & (g4155)) + ((g3038) & (!g3617) & (!g3050) & (!g3078) & (g3080) & (g4155)) + ((g3038) & (!g3617) & (!g3050) & (g3078) & (!g3080) & (g4155)) + ((g3038) & (!g3617) & (!g3050) & (g3078) & (g3080) & (g4155)) + ((g3038) & (!g3617) & (g3050) & (!g3078) & (g3080) & (g4155)) + ((g3038) & (!g3617) & (g3050) & (g3078) & (!g3080) & (g4155)) + ((g3038) & (!g3617) & (g3050) & (g3078) & (g3080) & (g4155)) + ((g3038) & (g3617) & (!g3050) & (g3078) & (g3080) & (g4155)) + ((g3038) & (g3617) & (g3050) & (!g3078) & (g3080) & (g4155)) + ((g3038) & (g3617) & (g3050) & (g3078) & (!g3080) & (g4155)) + ((g3038) & (g3617) & (g3050) & (g3078) & (g3080) & (g4155)));
	assign g4157 = (((g3113) & (g3125)));
	assign g4158 = (((!g3153) & (!g4156) & (!g4157) & (g3155)) + ((!g3153) & (!g4156) & (g4157) & (!g3155)) + ((!g3153) & (g4156) & (!g4157) & (!g3155)) + ((!g3153) & (g4156) & (g4157) & (!g3155)) + ((g3153) & (!g4156) & (!g4157) & (!g3155)) + ((g3153) & (!g4156) & (g4157) & (g3155)) + ((g3153) & (g4156) & (!g4157) & (g3155)) + ((g3153) & (g4156) & (g4157) & (g3155)));
	assign g4159 = (((!g830) & (!g1914) & (!g2041) & (!g4154) & (!g4158) & (key[225])) + ((!g830) & (!g1914) & (!g2041) & (!g4154) & (g4158) & (key[225])) + ((!g830) & (!g1914) & (!g2041) & (g4154) & (!g4158) & (key[225])) + ((!g830) & (!g1914) & (!g2041) & (g4154) & (g4158) & (key[225])) + ((!g830) & (!g1914) & (g2041) & (!g4154) & (!g4158) & (key[225])) + ((!g830) & (!g1914) & (g2041) & (!g4154) & (g4158) & (key[225])) + ((!g830) & (!g1914) & (g2041) & (g4154) & (!g4158) & (key[225])) + ((!g830) & (!g1914) & (g2041) & (g4154) & (g4158) & (key[225])) + ((!g830) & (g1914) & (!g2041) & (!g4154) & (!g4158) & (key[225])) + ((!g830) & (g1914) & (!g2041) & (!g4154) & (g4158) & (key[225])) + ((!g830) & (g1914) & (!g2041) & (g4154) & (!g4158) & (key[225])) + ((!g830) & (g1914) & (!g2041) & (g4154) & (g4158) & (key[225])) + ((!g830) & (g1914) & (g2041) & (!g4154) & (!g4158) & (key[225])) + ((!g830) & (g1914) & (g2041) & (!g4154) & (g4158) & (key[225])) + ((!g830) & (g1914) & (g2041) & (g4154) & (!g4158) & (key[225])) + ((!g830) & (g1914) & (g2041) & (g4154) & (g4158) & (key[225])) + ((g830) & (!g1914) & (!g2041) & (!g4154) & (g4158) & (!key[225])) + ((g830) & (!g1914) & (!g2041) & (!g4154) & (g4158) & (key[225])) + ((g830) & (!g1914) & (!g2041) & (g4154) & (g4158) & (!key[225])) + ((g830) & (!g1914) & (!g2041) & (g4154) & (g4158) & (key[225])) + ((g830) & (!g1914) & (g2041) & (!g4154) & (!g4158) & (!key[225])) + ((g830) & (!g1914) & (g2041) & (!g4154) & (!g4158) & (key[225])) + ((g830) & (!g1914) & (g2041) & (g4154) & (!g4158) & (!key[225])) + ((g830) & (!g1914) & (g2041) & (g4154) & (!g4158) & (key[225])) + ((g830) & (g1914) & (!g2041) & (g4154) & (!g4158) & (!key[225])) + ((g830) & (g1914) & (!g2041) & (g4154) & (!g4158) & (key[225])) + ((g830) & (g1914) & (!g2041) & (g4154) & (g4158) & (!key[225])) + ((g830) & (g1914) & (!g2041) & (g4154) & (g4158) & (key[225])) + ((g830) & (g1914) & (g2041) & (!g4154) & (!g4158) & (!key[225])) + ((g830) & (g1914) & (g2041) & (!g4154) & (!g4158) & (key[225])) + ((g830) & (g1914) & (g2041) & (!g4154) & (g4158) & (!key[225])) + ((g830) & (g1914) & (g2041) & (!g4154) & (g4158) & (key[225])));
	assign g4160 = (((!g2379) & (g3067) & (!g3725)) + ((g2379) & (!g3067) & (!g3725)) + ((g2379) & (g3067) & (!g3725)) + ((g2379) & (g3067) & (g3725)));
	assign g4161 = (((g1914) & (!g2427) & (!g3097) & (g4160)) + ((g1914) & (!g2427) & (g3097) & (!g4160)) + ((g1914) & (g2427) & (!g3097) & (!g4160)) + ((g1914) & (g2427) & (g3097) & (g4160)));
	assign g4162 = (((!g3053) & (!g3742) & (g3041)) + ((g3053) & (!g3742) & (!g3041)) + ((g3053) & (!g3742) & (g3041)) + ((g3053) & (g3742) & (g3041)));
	assign g4163 = (((!g1914) & (!g3088) & (!g3086) & (g4162)) + ((!g1914) & (!g3088) & (g3086) & (!g4162)) + ((!g1914) & (g3088) & (!g3086) & (!g4162)) + ((!g1914) & (g3088) & (g3086) & (g4162)));
	assign g4164 = (((!g830) & (!g2043) & (!g4161) & (!g4163) & (key[193])) + ((!g830) & (!g2043) & (!g4161) & (g4163) & (key[193])) + ((!g830) & (!g2043) & (g4161) & (!g4163) & (key[193])) + ((!g830) & (!g2043) & (g4161) & (g4163) & (key[193])) + ((!g830) & (g2043) & (!g4161) & (!g4163) & (key[193])) + ((!g830) & (g2043) & (!g4161) & (g4163) & (key[193])) + ((!g830) & (g2043) & (g4161) & (!g4163) & (key[193])) + ((!g830) & (g2043) & (g4161) & (g4163) & (key[193])) + ((g830) & (!g2043) & (!g4161) & (g4163) & (!key[193])) + ((g830) & (!g2043) & (!g4161) & (g4163) & (key[193])) + ((g830) & (!g2043) & (g4161) & (!g4163) & (!key[193])) + ((g830) & (!g2043) & (g4161) & (!g4163) & (key[193])) + ((g830) & (!g2043) & (g4161) & (g4163) & (!key[193])) + ((g830) & (!g2043) & (g4161) & (g4163) & (key[193])) + ((g830) & (g2043) & (!g4161) & (!g4163) & (!key[193])) + ((g830) & (g2043) & (!g4161) & (!g4163) & (key[193])));
	assign g4165 = (((!g2620) & (!g2672) & (!g2632) & (g2674) & (!g3855)) + ((!g2620) & (!g2672) & (!g2632) & (g2674) & (g3855)) + ((!g2620) & (!g2672) & (g2632) & (!g2674) & (g3855)) + ((!g2620) & (!g2672) & (g2632) & (g2674) & (!g3855)) + ((!g2620) & (g2672) & (!g2632) & (!g2674) & (!g3855)) + ((!g2620) & (g2672) & (!g2632) & (!g2674) & (g3855)) + ((!g2620) & (g2672) & (g2632) & (!g2674) & (!g3855)) + ((!g2620) & (g2672) & (g2632) & (g2674) & (g3855)) + ((g2620) & (!g2672) & (!g2632) & (!g2674) & (g3855)) + ((g2620) & (!g2672) & (!g2632) & (g2674) & (!g3855)) + ((g2620) & (!g2672) & (g2632) & (!g2674) & (!g3855)) + ((g2620) & (!g2672) & (g2632) & (!g2674) & (g3855)) + ((g2620) & (g2672) & (!g2632) & (!g2674) & (!g3855)) + ((g2620) & (g2672) & (!g2632) & (g2674) & (g3855)) + ((g2620) & (g2672) & (g2632) & (g2674) & (!g3855)) + ((g2620) & (g2672) & (g2632) & (g2674) & (g3855)));
	assign g4166 = (((!g2572) & (!g2637) & (g2584) & (g2640) & (!g3863) & (g3864)) + ((!g2572) & (!g2637) & (g2584) & (g2640) & (g3863) & (!g3864)) + ((!g2572) & (!g2637) & (g2584) & (g2640) & (g3863) & (g3864)) + ((!g2572) & (g2637) & (!g2584) & (g2640) & (!g3863) & (!g3864)) + ((!g2572) & (g2637) & (!g2584) & (g2640) & (!g3863) & (g3864)) + ((!g2572) & (g2637) & (!g2584) & (g2640) & (g3863) & (!g3864)) + ((!g2572) & (g2637) & (!g2584) & (g2640) & (g3863) & (g3864)) + ((!g2572) & (g2637) & (g2584) & (!g2640) & (!g3863) & (g3864)) + ((!g2572) & (g2637) & (g2584) & (!g2640) & (g3863) & (!g3864)) + ((!g2572) & (g2637) & (g2584) & (!g2640) & (g3863) & (g3864)) + ((!g2572) & (g2637) & (g2584) & (g2640) & (!g3863) & (!g3864)) + ((!g2572) & (g2637) & (g2584) & (g2640) & (!g3863) & (g3864)) + ((!g2572) & (g2637) & (g2584) & (g2640) & (g3863) & (!g3864)) + ((!g2572) & (g2637) & (g2584) & (g2640) & (g3863) & (g3864)) + ((g2572) & (!g2637) & (!g2584) & (g2640) & (!g3863) & (g3864)) + ((g2572) & (!g2637) & (!g2584) & (g2640) & (g3863) & (!g3864)) + ((g2572) & (!g2637) & (!g2584) & (g2640) & (g3863) & (g3864)) + ((g2572) & (!g2637) & (g2584) & (g2640) & (!g3863) & (!g3864)) + ((g2572) & (!g2637) & (g2584) & (g2640) & (!g3863) & (g3864)) + ((g2572) & (!g2637) & (g2584) & (g2640) & (g3863) & (!g3864)) + ((g2572) & (!g2637) & (g2584) & (g2640) & (g3863) & (g3864)) + ((g2572) & (g2637) & (!g2584) & (!g2640) & (!g3863) & (g3864)) + ((g2572) & (g2637) & (!g2584) & (!g2640) & (g3863) & (!g3864)) + ((g2572) & (g2637) & (!g2584) & (!g2640) & (g3863) & (g3864)) + ((g2572) & (g2637) & (!g2584) & (g2640) & (!g3863) & (!g3864)) + ((g2572) & (g2637) & (!g2584) & (g2640) & (!g3863) & (g3864)) + ((g2572) & (g2637) & (!g2584) & (g2640) & (g3863) & (!g3864)) + ((g2572) & (g2637) & (!g2584) & (g2640) & (g3863) & (g3864)) + ((g2572) & (g2637) & (g2584) & (!g2640) & (!g3863) & (!g3864)) + ((g2572) & (g2637) & (g2584) & (!g2640) & (!g3863) & (g3864)) + ((g2572) & (g2637) & (g2584) & (!g2640) & (g3863) & (!g3864)) + ((g2572) & (g2637) & (g2584) & (!g2640) & (g3863) & (g3864)) + ((g2572) & (g2637) & (g2584) & (g2640) & (!g3863) & (!g3864)) + ((g2572) & (g2637) & (g2584) & (g2640) & (!g3863) & (g3864)) + ((g2572) & (g2637) & (g2584) & (g2640) & (g3863) & (!g3864)) + ((g2572) & (g2637) & (g2584) & (g2640) & (g3863) & (g3864)));
	assign g4167 = (((!g3502) & (!g3503)));
	assign g4168 = (((g1914) & (!g1031) & (!g4167) & (!g2233)) + ((g1914) & (!g1031) & (g4167) & (g2233)) + ((g1914) & (g1031) & (!g4167) & (g2233)) + ((g1914) & (g1031) & (g4167) & (!g2233)));
	assign g4169 = (((!g3519) & (!g3520)));
	assign g4170 = (((!g1914) & (!g2224) & (!g2230) & (!g4169)) + ((!g1914) & (!g2224) & (g2230) & (g4169)) + ((!g1914) & (g2224) & (!g2230) & (g4169)) + ((!g1914) & (g2224) & (g2230) & (!g4169)));
	assign g4171 = (((!g830) & (!g2047) & (!g4168) & (!g4170) & (key[47])) + ((!g830) & (!g2047) & (!g4168) & (g4170) & (key[47])) + ((!g830) & (!g2047) & (g4168) & (!g4170) & (key[47])) + ((!g830) & (!g2047) & (g4168) & (g4170) & (key[47])) + ((!g830) & (g2047) & (!g4168) & (!g4170) & (key[47])) + ((!g830) & (g2047) & (!g4168) & (g4170) & (key[47])) + ((!g830) & (g2047) & (g4168) & (!g4170) & (key[47])) + ((!g830) & (g2047) & (g4168) & (g4170) & (key[47])) + ((g830) & (!g2047) & (!g4168) & (g4170) & (!key[47])) + ((g830) & (!g2047) & (!g4168) & (g4170) & (key[47])) + ((g830) & (!g2047) & (g4168) & (!g4170) & (!key[47])) + ((g830) & (!g2047) & (g4168) & (!g4170) & (key[47])) + ((g830) & (!g2047) & (g4168) & (g4170) & (!key[47])) + ((g830) & (!g2047) & (g4168) & (g4170) & (key[47])) + ((g830) & (g2047) & (!g4168) & (!g4170) & (!key[47])) + ((g830) & (g2047) & (!g4168) & (!g4170) & (key[47])));
	assign g4172 = (((!g1890) & (!g1939) & (!g1941) & (!g1898) & (!g2022) & (g2071)) + ((!g1890) & (!g1939) & (!g1941) & (!g1898) & (g2022) & (g2071)) + ((!g1890) & (!g1939) & (!g1941) & (g1898) & (!g2022) & (g2071)) + ((!g1890) & (!g1939) & (!g1941) & (g1898) & (g2022) & (g2071)) + ((!g1890) & (!g1939) & (g1941) & (!g1898) & (!g2022) & (!g2071)) + ((!g1890) & (!g1939) & (g1941) & (!g1898) & (g2022) & (!g2071)) + ((!g1890) & (!g1939) & (g1941) & (g1898) & (!g2022) & (!g2071)) + ((!g1890) & (!g1939) & (g1941) & (g1898) & (g2022) & (!g2071)) + ((!g1890) & (g1939) & (!g1941) & (!g1898) & (!g2022) & (g2071)) + ((!g1890) & (g1939) & (!g1941) & (!g1898) & (g2022) & (!g2071)) + ((!g1890) & (g1939) & (!g1941) & (g1898) & (!g2022) & (g2071)) + ((!g1890) & (g1939) & (!g1941) & (g1898) & (g2022) & (!g2071)) + ((!g1890) & (g1939) & (g1941) & (!g1898) & (!g2022) & (!g2071)) + ((!g1890) & (g1939) & (g1941) & (!g1898) & (g2022) & (g2071)) + ((!g1890) & (g1939) & (g1941) & (g1898) & (!g2022) & (!g2071)) + ((!g1890) & (g1939) & (g1941) & (g1898) & (g2022) & (g2071)) + ((g1890) & (!g1939) & (!g1941) & (!g1898) & (!g2022) & (g2071)) + ((g1890) & (!g1939) & (!g1941) & (!g1898) & (g2022) & (g2071)) + ((g1890) & (!g1939) & (!g1941) & (g1898) & (!g2022) & (g2071)) + ((g1890) & (!g1939) & (!g1941) & (g1898) & (g2022) & (!g2071)) + ((g1890) & (!g1939) & (g1941) & (!g1898) & (!g2022) & (!g2071)) + ((g1890) & (!g1939) & (g1941) & (!g1898) & (g2022) & (!g2071)) + ((g1890) & (!g1939) & (g1941) & (g1898) & (!g2022) & (!g2071)) + ((g1890) & (!g1939) & (g1941) & (g1898) & (g2022) & (g2071)) + ((g1890) & (g1939) & (!g1941) & (!g1898) & (!g2022) & (g2071)) + ((g1890) & (g1939) & (!g1941) & (!g1898) & (g2022) & (!g2071)) + ((g1890) & (g1939) & (!g1941) & (g1898) & (!g2022) & (!g2071)) + ((g1890) & (g1939) & (!g1941) & (g1898) & (g2022) & (!g2071)) + ((g1890) & (g1939) & (g1941) & (!g1898) & (!g2022) & (!g2071)) + ((g1890) & (g1939) & (g1941) & (!g1898) & (g2022) & (g2071)) + ((g1890) & (g1939) & (g1941) & (g1898) & (!g2022) & (g2071)) + ((g1890) & (g1939) & (g1941) & (g1898) & (g2022) & (g2071)));
	assign g4173 = (((!g2334) & (!g2340) & (!g3763)) + ((!g2334) & (g2340) & (g3763)) + ((g2334) & (!g2340) & (g3763)) + ((g2334) & (g2340) & (!g3763)));
	assign g4174 = (((!g830) & (!g1914) & (!g2048) & (!g4172) & (!g4173) & (key[79])) + ((!g830) & (!g1914) & (!g2048) & (!g4172) & (g4173) & (key[79])) + ((!g830) & (!g1914) & (!g2048) & (g4172) & (!g4173) & (key[79])) + ((!g830) & (!g1914) & (!g2048) & (g4172) & (g4173) & (key[79])) + ((!g830) & (!g1914) & (g2048) & (!g4172) & (!g4173) & (key[79])) + ((!g830) & (!g1914) & (g2048) & (!g4172) & (g4173) & (key[79])) + ((!g830) & (!g1914) & (g2048) & (g4172) & (!g4173) & (key[79])) + ((!g830) & (!g1914) & (g2048) & (g4172) & (g4173) & (key[79])) + ((!g830) & (g1914) & (!g2048) & (!g4172) & (!g4173) & (key[79])) + ((!g830) & (g1914) & (!g2048) & (!g4172) & (g4173) & (key[79])) + ((!g830) & (g1914) & (!g2048) & (g4172) & (!g4173) & (key[79])) + ((!g830) & (g1914) & (!g2048) & (g4172) & (g4173) & (key[79])) + ((!g830) & (g1914) & (g2048) & (!g4172) & (!g4173) & (key[79])) + ((!g830) & (g1914) & (g2048) & (!g4172) & (g4173) & (key[79])) + ((!g830) & (g1914) & (g2048) & (g4172) & (!g4173) & (key[79])) + ((!g830) & (g1914) & (g2048) & (g4172) & (g4173) & (key[79])) + ((g830) & (!g1914) & (!g2048) & (!g4172) & (g4173) & (!key[79])) + ((g830) & (!g1914) & (!g2048) & (!g4172) & (g4173) & (key[79])) + ((g830) & (!g1914) & (!g2048) & (g4172) & (g4173) & (!key[79])) + ((g830) & (!g1914) & (!g2048) & (g4172) & (g4173) & (key[79])) + ((g830) & (!g1914) & (g2048) & (!g4172) & (!g4173) & (!key[79])) + ((g830) & (!g1914) & (g2048) & (!g4172) & (!g4173) & (key[79])) + ((g830) & (!g1914) & (g2048) & (g4172) & (!g4173) & (!key[79])) + ((g830) & (!g1914) & (g2048) & (g4172) & (!g4173) & (key[79])) + ((g830) & (g1914) & (!g2048) & (g4172) & (!g4173) & (!key[79])) + ((g830) & (g1914) & (!g2048) & (g4172) & (!g4173) & (key[79])) + ((g830) & (g1914) & (!g2048) & (g4172) & (g4173) & (!key[79])) + ((g830) & (g1914) & (!g2048) & (g4172) & (g4173) & (key[79])) + ((g830) & (g1914) & (g2048) & (!g4172) & (!g4173) & (!key[79])) + ((g830) & (g1914) & (g2048) & (!g4172) & (!g4173) & (key[79])) + ((g830) & (g1914) & (g2048) & (!g4172) & (g4173) & (!key[79])) + ((g830) & (g1914) & (g2048) & (!g4172) & (g4173) & (key[79])));
	assign g4175 = (((!g3412) & (g3413)) + ((g3412) & (!g3413)) + ((g3412) & (g3413)));
	assign g4176 = (((!g3394) & (g3395)) + ((g3394) & (!g3395)) + ((g3394) & (g3395)));
	assign g8293 = (((!g5560) & (g5586) & (!g4177)) + ((!g5560) & (g5586) & (g4177)) + ((g5560) & (!g5586) & (g4177)) + ((g5560) & (g5586) & (g4177)));
	assign g4178 = (((!g830) & (!g2051) & (!g6861) & (g4177)) + ((!g830) & (!g2051) & (g6861) & (g4177)) + ((!g830) & (g2051) & (!g6861) & (g4177)) + ((!g830) & (g2051) & (g6861) & (g4177)) + ((g830) & (!g2051) & (g6861) & (!g4177)) + ((g830) & (!g2051) & (g6861) & (g4177)) + ((g830) & (g2051) & (!g6861) & (!g4177)) + ((g830) & (g2051) & (!g6861) & (g4177)));
	assign g4179 = (((!g3469) & (!g2317) & (!g2340)) + ((!g3469) & (g2317) & (g2340)) + ((g3469) & (!g2317) & (g2340)) + ((g3469) & (g2317) & (!g2340)));
	assign g4180 = (((!g1884) & (!g1977) & (!g1979) & (!g1886) & (!g2032) & (g2055)) + ((!g1884) & (!g1977) & (!g1979) & (!g1886) & (g2032) & (g2055)) + ((!g1884) & (!g1977) & (!g1979) & (g1886) & (!g2032) & (g2055)) + ((!g1884) & (!g1977) & (!g1979) & (g1886) & (g2032) & (g2055)) + ((!g1884) & (!g1977) & (g1979) & (!g1886) & (!g2032) & (!g2055)) + ((!g1884) & (!g1977) & (g1979) & (!g1886) & (g2032) & (!g2055)) + ((!g1884) & (!g1977) & (g1979) & (g1886) & (!g2032) & (!g2055)) + ((!g1884) & (!g1977) & (g1979) & (g1886) & (g2032) & (!g2055)) + ((!g1884) & (g1977) & (!g1979) & (!g1886) & (!g2032) & (g2055)) + ((!g1884) & (g1977) & (!g1979) & (!g1886) & (g2032) & (!g2055)) + ((!g1884) & (g1977) & (!g1979) & (g1886) & (!g2032) & (g2055)) + ((!g1884) & (g1977) & (!g1979) & (g1886) & (g2032) & (!g2055)) + ((!g1884) & (g1977) & (g1979) & (!g1886) & (!g2032) & (!g2055)) + ((!g1884) & (g1977) & (g1979) & (!g1886) & (g2032) & (g2055)) + ((!g1884) & (g1977) & (g1979) & (g1886) & (!g2032) & (!g2055)) + ((!g1884) & (g1977) & (g1979) & (g1886) & (g2032) & (g2055)) + ((g1884) & (!g1977) & (!g1979) & (!g1886) & (!g2032) & (g2055)) + ((g1884) & (!g1977) & (!g1979) & (!g1886) & (g2032) & (g2055)) + ((g1884) & (!g1977) & (!g1979) & (g1886) & (!g2032) & (g2055)) + ((g1884) & (!g1977) & (!g1979) & (g1886) & (g2032) & (!g2055)) + ((g1884) & (!g1977) & (g1979) & (!g1886) & (!g2032) & (!g2055)) + ((g1884) & (!g1977) & (g1979) & (!g1886) & (g2032) & (!g2055)) + ((g1884) & (!g1977) & (g1979) & (g1886) & (!g2032) & (!g2055)) + ((g1884) & (!g1977) & (g1979) & (g1886) & (g2032) & (g2055)) + ((g1884) & (g1977) & (!g1979) & (!g1886) & (!g2032) & (g2055)) + ((g1884) & (g1977) & (!g1979) & (!g1886) & (g2032) & (!g2055)) + ((g1884) & (g1977) & (!g1979) & (g1886) & (!g2032) & (!g2055)) + ((g1884) & (g1977) & (!g1979) & (g1886) & (g2032) & (!g2055)) + ((g1884) & (g1977) & (g1979) & (!g1886) & (!g2032) & (!g2055)) + ((g1884) & (g1977) & (g1979) & (!g1886) & (g2032) & (g2055)) + ((g1884) & (g1977) & (g1979) & (g1886) & (!g2032) & (g2055)) + ((g1884) & (g1977) & (g1979) & (g1886) & (g2032) & (g2055)));
	assign g4181 = (((!g830) & (!g1914) & (!g2052) & (!g4179) & (!g4180) & (key[175])) + ((!g830) & (!g1914) & (!g2052) & (!g4179) & (g4180) & (key[175])) + ((!g830) & (!g1914) & (!g2052) & (g4179) & (!g4180) & (key[175])) + ((!g830) & (!g1914) & (!g2052) & (g4179) & (g4180) & (key[175])) + ((!g830) & (!g1914) & (g2052) & (!g4179) & (!g4180) & (key[175])) + ((!g830) & (!g1914) & (g2052) & (!g4179) & (g4180) & (key[175])) + ((!g830) & (!g1914) & (g2052) & (g4179) & (!g4180) & (key[175])) + ((!g830) & (!g1914) & (g2052) & (g4179) & (g4180) & (key[175])) + ((!g830) & (g1914) & (!g2052) & (!g4179) & (!g4180) & (key[175])) + ((!g830) & (g1914) & (!g2052) & (!g4179) & (g4180) & (key[175])) + ((!g830) & (g1914) & (!g2052) & (g4179) & (!g4180) & (key[175])) + ((!g830) & (g1914) & (!g2052) & (g4179) & (g4180) & (key[175])) + ((!g830) & (g1914) & (g2052) & (!g4179) & (!g4180) & (key[175])) + ((!g830) & (g1914) & (g2052) & (!g4179) & (g4180) & (key[175])) + ((!g830) & (g1914) & (g2052) & (g4179) & (!g4180) & (key[175])) + ((!g830) & (g1914) & (g2052) & (g4179) & (g4180) & (key[175])) + ((g830) & (!g1914) & (!g2052) & (!g4179) & (g4180) & (!key[175])) + ((g830) & (!g1914) & (!g2052) & (!g4179) & (g4180) & (key[175])) + ((g830) & (!g1914) & (!g2052) & (g4179) & (g4180) & (!key[175])) + ((g830) & (!g1914) & (!g2052) & (g4179) & (g4180) & (key[175])) + ((g830) & (!g1914) & (g2052) & (!g4179) & (!g4180) & (!key[175])) + ((g830) & (!g1914) & (g2052) & (!g4179) & (!g4180) & (key[175])) + ((g830) & (!g1914) & (g2052) & (g4179) & (!g4180) & (!key[175])) + ((g830) & (!g1914) & (g2052) & (g4179) & (!g4180) & (key[175])) + ((g830) & (g1914) & (!g2052) & (g4179) & (!g4180) & (!key[175])) + ((g830) & (g1914) & (!g2052) & (g4179) & (!g4180) & (key[175])) + ((g830) & (g1914) & (!g2052) & (g4179) & (g4180) & (!key[175])) + ((g830) & (g1914) & (!g2052) & (g4179) & (g4180) & (key[175])) + ((g830) & (g1914) & (g2052) & (!g4179) & (!g4180) & (!key[175])) + ((g830) & (g1914) & (g2052) & (!g4179) & (!g4180) & (key[175])) + ((g830) & (g1914) & (g2052) & (!g4179) & (g4180) & (!key[175])) + ((g830) & (g1914) & (g2052) & (!g4179) & (g4180) & (key[175])));
	assign g4182 = (((!g2887) & (g2902)) + ((g2887) & (!g2902)));
	assign g4183 = (((!g3442) & (!g2807) & (!g2830) & (g2857) & (g2863) & (g4182)) + ((!g3442) & (!g2807) & (g2830) & (!g2857) & (g2863) & (g4182)) + ((!g3442) & (!g2807) & (g2830) & (g2857) & (!g2863) & (g4182)) + ((!g3442) & (!g2807) & (g2830) & (g2857) & (g2863) & (g4182)) + ((!g3442) & (g2807) & (!g2830) & (!g2857) & (g2863) & (g4182)) + ((!g3442) & (g2807) & (!g2830) & (g2857) & (!g2863) & (g4182)) + ((!g3442) & (g2807) & (!g2830) & (g2857) & (g2863) & (g4182)) + ((!g3442) & (g2807) & (g2830) & (!g2857) & (g2863) & (g4182)) + ((!g3442) & (g2807) & (g2830) & (g2857) & (!g2863) & (g4182)) + ((!g3442) & (g2807) & (g2830) & (g2857) & (g2863) & (g4182)) + ((g3442) & (!g2807) & (!g2830) & (g2857) & (g2863) & (g4182)) + ((g3442) & (!g2807) & (g2830) & (g2857) & (g2863) & (g4182)) + ((g3442) & (g2807) & (!g2830) & (g2857) & (g2863) & (g4182)) + ((g3442) & (g2807) & (g2830) & (!g2857) & (g2863) & (g4182)) + ((g3442) & (g2807) & (g2830) & (g2857) & (!g2863) & (g4182)) + ((g3442) & (g2807) & (g2830) & (g2857) & (g2863) & (g4182)));
	assign g4184 = (((g2887) & (g2902)));
	assign g4185 = (((!g2956) & (!g4183) & (!g4184) & (g2968)) + ((!g2956) & (!g4183) & (g4184) & (!g2968)) + ((!g2956) & (g4183) & (!g4184) & (!g2968)) + ((!g2956) & (g4183) & (g4184) & (!g2968)) + ((g2956) & (!g4183) & (!g4184) & (!g2968)) + ((g2956) & (!g4183) & (g4184) & (g2968)) + ((g2956) & (g4183) & (!g4184) & (g2968)) + ((g2956) & (g4183) & (g4184) & (g2968)));
	assign g4186 = (((!g2556) & (!g1711) & (!g4137) & (!g4138)) + ((!g2556) & (!g1711) & (!g4137) & (g4138)) + ((!g2556) & (!g1711) & (g4137) & (!g4138)) + ((!g2556) & (!g1711) & (g4137) & (g4138)) + ((!g2556) & (g1711) & (!g4137) & (!g4138)) + ((g2556) & (!g1711) & (!g4137) & (!g4138)));
	assign g4187 = (((!g1914) & (!g2602) & (!g1744) & (!g4185) & (!g4186)) + ((!g1914) & (!g2602) & (!g1744) & (g4185) & (!g4186)) + ((!g1914) & (!g2602) & (g1744) & (!g4185) & (g4186)) + ((!g1914) & (!g2602) & (g1744) & (g4185) & (g4186)) + ((!g1914) & (g2602) & (!g1744) & (!g4185) & (g4186)) + ((!g1914) & (g2602) & (!g1744) & (g4185) & (g4186)) + ((!g1914) & (g2602) & (g1744) & (!g4185) & (!g4186)) + ((!g1914) & (g2602) & (g1744) & (g4185) & (!g4186)) + ((g1914) & (!g2602) & (!g1744) & (g4185) & (!g4186)) + ((g1914) & (!g2602) & (!g1744) & (g4185) & (g4186)) + ((g1914) & (!g2602) & (g1744) & (g4185) & (!g4186)) + ((g1914) & (!g2602) & (g1744) & (g4185) & (g4186)) + ((g1914) & (g2602) & (!g1744) & (g4185) & (!g4186)) + ((g1914) & (g2602) & (!g1744) & (g4185) & (g4186)) + ((g1914) & (g2602) & (g1744) & (g4185) & (!g4186)) + ((g1914) & (g2602) & (g1744) & (g4185) & (g4186)));
	assign g4188 = (((!g830) & (!g2055) & (!g4187) & (key[98])) + ((!g830) & (!g2055) & (g4187) & (key[98])) + ((!g830) & (g2055) & (!g4187) & (key[98])) + ((!g830) & (g2055) & (g4187) & (key[98])) + ((g830) & (!g2055) & (g4187) & (!key[98])) + ((g830) & (!g2055) & (g4187) & (key[98])) + ((g830) & (g2055) & (!g4187) & (!key[98])) + ((g830) & (g2055) & (!g4187) & (key[98])));
	assign g4189 = (((!g2051) & (g2659)) + ((g2051) & (!g2659)));
	assign g4190 = (((!g2011) & (!g2013) & (g3542) & (g2569) & (g2626) & (g4189)) + ((!g2011) & (g2013) & (!g3542) & (!g2569) & (g2626) & (g4189)) + ((!g2011) & (g2013) & (!g3542) & (g2569) & (g2626) & (g4189)) + ((!g2011) & (g2013) & (g3542) & (!g2569) & (g2626) & (g4189)) + ((!g2011) & (g2013) & (g3542) & (g2569) & (!g2626) & (g4189)) + ((!g2011) & (g2013) & (g3542) & (g2569) & (g2626) & (g4189)) + ((g2011) & (!g2013) & (!g3542) & (g2569) & (g2626) & (g4189)) + ((g2011) & (!g2013) & (g3542) & (!g2569) & (g2626) & (g4189)) + ((g2011) & (!g2013) & (g3542) & (g2569) & (g2626) & (g4189)) + ((g2011) & (g2013) & (!g3542) & (!g2569) & (g2626) & (g4189)) + ((g2011) & (g2013) & (!g3542) & (g2569) & (!g2626) & (g4189)) + ((g2011) & (g2013) & (!g3542) & (g2569) & (g2626) & (g4189)) + ((g2011) & (g2013) & (g3542) & (!g2569) & (!g2626) & (g4189)) + ((g2011) & (g2013) & (g3542) & (!g2569) & (g2626) & (g4189)) + ((g2011) & (g2013) & (g3542) & (g2569) & (!g2626) & (g4189)) + ((g2011) & (g2013) & (g3542) & (g2569) & (g2626) & (g4189)));
	assign g4191 = (((g2051) & (g2659)));
	assign g4192 = (((!g4190) & (g4191)) + ((g4190) & (!g4191)) + ((g4190) & (g4191)));
	assign g4193 = (((!g2047) & (!g2098) & (!g2665) & (g2708) & (!g4121)) + ((!g2047) & (!g2098) & (!g2665) & (g2708) & (g4121)) + ((!g2047) & (!g2098) & (g2665) & (!g2708) & (g4121)) + ((!g2047) & (!g2098) & (g2665) & (g2708) & (!g4121)) + ((!g2047) & (g2098) & (!g2665) & (!g2708) & (!g4121)) + ((!g2047) & (g2098) & (!g2665) & (!g2708) & (g4121)) + ((!g2047) & (g2098) & (g2665) & (!g2708) & (!g4121)) + ((!g2047) & (g2098) & (g2665) & (g2708) & (g4121)) + ((g2047) & (!g2098) & (!g2665) & (!g2708) & (g4121)) + ((g2047) & (!g2098) & (!g2665) & (g2708) & (!g4121)) + ((g2047) & (!g2098) & (g2665) & (!g2708) & (!g4121)) + ((g2047) & (!g2098) & (g2665) & (!g2708) & (g4121)) + ((g2047) & (g2098) & (!g2665) & (!g2708) & (!g4121)) + ((g2047) & (g2098) & (!g2665) & (g2708) & (g4121)) + ((g2047) & (g2098) & (g2665) & (g2708) & (!g4121)) + ((g2047) & (g2098) & (g2665) & (g2708) & (g4121)));
	assign g4194 = (((!g3163) & (!g4142) & (!g4143) & (!g3149)) + ((!g3163) & (!g4142) & (!g4143) & (g3149)) + ((!g3163) & (!g4142) & (g4143) & (!g3149)) + ((!g3163) & (g4142) & (!g4143) & (!g3149)) + ((!g3163) & (g4142) & (g4143) & (!g3149)) + ((g3163) & (!g4142) & (!g4143) & (!g3149)));
	assign g4195 = (((!g2256) & (g2889)) + ((g2256) & (!g2889)));
	assign g4196 = (((!g2177) & (!g2210) & (g2810) & (g2868) & (!g3584) & (g4195)) + ((!g2177) & (g2210) & (!g2810) & (g2868) & (!g3584) & (g4195)) + ((!g2177) & (g2210) & (!g2810) & (g2868) & (g3584) & (g4195)) + ((!g2177) & (g2210) & (g2810) & (!g2868) & (!g3584) & (g4195)) + ((!g2177) & (g2210) & (g2810) & (g2868) & (!g3584) & (g4195)) + ((!g2177) & (g2210) & (g2810) & (g2868) & (g3584) & (g4195)) + ((g2177) & (!g2210) & (!g2810) & (g2868) & (!g3584) & (g4195)) + ((g2177) & (!g2210) & (g2810) & (g2868) & (!g3584) & (g4195)) + ((g2177) & (!g2210) & (g2810) & (g2868) & (g3584) & (g4195)) + ((g2177) & (g2210) & (!g2810) & (!g2868) & (!g3584) & (g4195)) + ((g2177) & (g2210) & (!g2810) & (g2868) & (!g3584) & (g4195)) + ((g2177) & (g2210) & (!g2810) & (g2868) & (g3584) & (g4195)) + ((g2177) & (g2210) & (g2810) & (!g2868) & (!g3584) & (g4195)) + ((g2177) & (g2210) & (g2810) & (!g2868) & (g3584) & (g4195)) + ((g2177) & (g2210) & (g2810) & (g2868) & (!g3584) & (g4195)) + ((g2177) & (g2210) & (g2810) & (g2868) & (g3584) & (g4195)));
	assign g4197 = (((g2256) & (g2889)));
	assign g4198 = (((!g2295) & (!g2979) & (!g4196) & (g4197)) + ((!g2295) & (!g2979) & (g4196) & (!g4197)) + ((!g2295) & (!g2979) & (g4196) & (g4197)) + ((!g2295) & (g2979) & (!g4196) & (!g4197)) + ((g2295) & (!g2979) & (!g4196) & (!g4197)) + ((g2295) & (g2979) & (!g4196) & (g4197)) + ((g2295) & (g2979) & (g4196) & (!g4197)) + ((g2295) & (g2979) & (g4196) & (g4197)));
	assign g4199 = (((!g1914) & (!g4194) & (!g3193) & (!g3199) & (g4198)) + ((!g1914) & (!g4194) & (!g3193) & (g3199) & (g4198)) + ((!g1914) & (!g4194) & (g3193) & (!g3199) & (g4198)) + ((!g1914) & (!g4194) & (g3193) & (g3199) & (g4198)) + ((!g1914) & (g4194) & (!g3193) & (!g3199) & (g4198)) + ((!g1914) & (g4194) & (!g3193) & (g3199) & (g4198)) + ((!g1914) & (g4194) & (g3193) & (!g3199) & (g4198)) + ((!g1914) & (g4194) & (g3193) & (g3199) & (g4198)) + ((g1914) & (!g4194) & (!g3193) & (!g3199) & (!g4198)) + ((g1914) & (!g4194) & (!g3193) & (!g3199) & (g4198)) + ((g1914) & (!g4194) & (g3193) & (g3199) & (!g4198)) + ((g1914) & (!g4194) & (g3193) & (g3199) & (g4198)) + ((g1914) & (g4194) & (!g3193) & (g3199) & (!g4198)) + ((g1914) & (g4194) & (!g3193) & (g3199) & (g4198)) + ((g1914) & (g4194) & (g3193) & (!g3199) & (!g4198)) + ((g1914) & (g4194) & (g3193) & (!g3199) & (g4198)));
	assign g4200 = (((!g830) & (!g2065) & (!g4199) & (nonce[2])) + ((!g830) & (!g2065) & (g4199) & (nonce[2])) + ((!g830) & (g2065) & (!g4199) & (nonce[2])) + ((!g830) & (g2065) & (g4199) & (nonce[2])) + ((g830) & (!g2065) & (g4199) & (!nonce[2])) + ((g830) & (!g2065) & (g4199) & (nonce[2])) + ((g830) & (g2065) & (!g4199) & (!nonce[2])) + ((g830) & (g2065) & (!g4199) & (nonce[2])));
	assign g4201 = (((!g2263) & (g2897)) + ((g2263) & (!g2897)));
	assign g4202 = (((!g2181) & (!g2213) & (!g3600) & (g2822) & (g2871) & (g4201)) + ((!g2181) & (g2213) & (!g3600) & (!g2822) & (g2871) & (g4201)) + ((!g2181) & (g2213) & (!g3600) & (g2822) & (!g2871) & (g4201)) + ((!g2181) & (g2213) & (!g3600) & (g2822) & (g2871) & (g4201)) + ((!g2181) & (g2213) & (g3600) & (!g2822) & (g2871) & (g4201)) + ((!g2181) & (g2213) & (g3600) & (g2822) & (g2871) & (g4201)) + ((g2181) & (!g2213) & (!g3600) & (!g2822) & (g2871) & (g4201)) + ((g2181) & (!g2213) & (!g3600) & (g2822) & (g2871) & (g4201)) + ((g2181) & (!g2213) & (g3600) & (g2822) & (g2871) & (g4201)) + ((g2181) & (g2213) & (!g3600) & (!g2822) & (!g2871) & (g4201)) + ((g2181) & (g2213) & (!g3600) & (!g2822) & (g2871) & (g4201)) + ((g2181) & (g2213) & (!g3600) & (g2822) & (!g2871) & (g4201)) + ((g2181) & (g2213) & (!g3600) & (g2822) & (g2871) & (g4201)) + ((g2181) & (g2213) & (g3600) & (!g2822) & (g2871) & (g4201)) + ((g2181) & (g2213) & (g3600) & (g2822) & (!g2871) & (g4201)) + ((g2181) & (g2213) & (g3600) & (g2822) & (g2871) & (g4201)));
	assign g4203 = (((g2263) & (g2897)));
	assign g4204 = (((!g2299) & (!g4202) & (!g4203) & (g2985)) + ((!g2299) & (!g4202) & (g4203) & (!g2985)) + ((!g2299) & (g4202) & (!g4203) & (!g2985)) + ((!g2299) & (g4202) & (g4203) & (!g2985)) + ((g2299) & (!g4202) & (!g4203) & (!g2985)) + ((g2299) & (!g4202) & (g4203) & (g2985)) + ((g2299) & (g4202) & (!g4203) & (g2985)) + ((g2299) & (g4202) & (g4203) & (g2985)));
	assign g4205 = (((!g3153) & (!g4156) & (!g4157) & (!g3155)) + ((!g3153) & (!g4156) & (!g4157) & (g3155)) + ((!g3153) & (!g4156) & (g4157) & (!g3155)) + ((!g3153) & (g4156) & (!g4157) & (!g3155)) + ((!g3153) & (g4156) & (g4157) & (!g3155)) + ((g3153) & (!g4156) & (!g4157) & (!g3155)));
	assign g4206 = (((!g1914) & (!g4204) & (!g4205) & (!g3184) & (!g3196)) + ((!g1914) & (!g4204) & (!g4205) & (g3184) & (g3196)) + ((!g1914) & (!g4204) & (g4205) & (!g3184) & (g3196)) + ((!g1914) & (!g4204) & (g4205) & (g3184) & (!g3196)) + ((!g1914) & (g4204) & (!g4205) & (!g3184) & (!g3196)) + ((!g1914) & (g4204) & (!g4205) & (g3184) & (g3196)) + ((!g1914) & (g4204) & (g4205) & (!g3184) & (g3196)) + ((!g1914) & (g4204) & (g4205) & (g3184) & (!g3196)) + ((g1914) & (g4204) & (!g4205) & (!g3184) & (!g3196)) + ((g1914) & (g4204) & (!g4205) & (!g3184) & (g3196)) + ((g1914) & (g4204) & (!g4205) & (g3184) & (!g3196)) + ((g1914) & (g4204) & (!g4205) & (g3184) & (g3196)) + ((g1914) & (g4204) & (g4205) & (!g3184) & (!g3196)) + ((g1914) & (g4204) & (g4205) & (!g3184) & (g3196)) + ((g1914) & (g4204) & (g4205) & (g3184) & (!g3196)) + ((g1914) & (g4204) & (g4205) & (g3184) & (g3196)));
	assign g4207 = (((!g830) & (!g2068) & (!g4206) & (key[226])) + ((!g830) & (!g2068) & (g4206) & (key[226])) + ((!g830) & (g2068) & (!g4206) & (key[226])) + ((!g830) & (g2068) & (g4206) & (key[226])) + ((g830) & (!g2068) & (g4206) & (!key[226])) + ((g830) & (!g2068) & (g4206) & (key[226])) + ((g830) & (g2068) & (!g4206) & (!key[226])) + ((g830) & (g2068) & (!g4206) & (key[226])));
	assign g4208 = (((!g2552) & (!g1711) & (!g4115) & (!g4116)) + ((!g2552) & (!g1711) & (!g4115) & (g4116)) + ((!g2552) & (!g1711) & (g4115) & (!g4116)) + ((!g2552) & (!g1711) & (g4115) & (g4116)) + ((!g2552) & (g1711) & (!g4115) & (!g4116)) + ((g2552) & (!g1711) & (!g4115) & (!g4116)));
	assign g4209 = (((!g2893) & (g2897)) + ((g2893) & (!g2897)));
	assign g4210 = (((!g2822) & (!g2871) & (!g3650) & (g2816) & (g2848) & (g4209)) + ((!g2822) & (g2871) & (!g3650) & (!g2816) & (g2848) & (g4209)) + ((!g2822) & (g2871) & (!g3650) & (g2816) & (!g2848) & (g4209)) + ((!g2822) & (g2871) & (!g3650) & (g2816) & (g2848) & (g4209)) + ((!g2822) & (g2871) & (g3650) & (!g2816) & (g2848) & (g4209)) + ((!g2822) & (g2871) & (g3650) & (g2816) & (g2848) & (g4209)) + ((g2822) & (!g2871) & (!g3650) & (!g2816) & (g2848) & (g4209)) + ((g2822) & (!g2871) & (!g3650) & (g2816) & (g2848) & (g4209)) + ((g2822) & (!g2871) & (g3650) & (g2816) & (g2848) & (g4209)) + ((g2822) & (g2871) & (!g3650) & (!g2816) & (!g2848) & (g4209)) + ((g2822) & (g2871) & (!g3650) & (!g2816) & (g2848) & (g4209)) + ((g2822) & (g2871) & (!g3650) & (g2816) & (!g2848) & (g4209)) + ((g2822) & (g2871) & (!g3650) & (g2816) & (g2848) & (g4209)) + ((g2822) & (g2871) & (g3650) & (!g2816) & (g2848) & (g4209)) + ((g2822) & (g2871) & (g3650) & (g2816) & (!g2848) & (g4209)) + ((g2822) & (g2871) & (g3650) & (g2816) & (g2848) & (g4209)));
	assign g4211 = (((g2893) & (g2897)));
	assign g4212 = (((!g2938) & (!g2985) & (!g4210) & (g4211)) + ((!g2938) & (!g2985) & (g4210) & (!g4211)) + ((!g2938) & (!g2985) & (g4210) & (g4211)) + ((!g2938) & (g2985) & (!g4210) & (!g4211)) + ((g2938) & (!g2985) & (!g4210) & (!g4211)) + ((g2938) & (g2985) & (!g4210) & (g4211)) + ((g2938) & (g2985) & (g4210) & (!g4211)) + ((g2938) & (g2985) & (g4210) & (g4211)));
	assign g4213 = (((!g1914) & (!g2599) & (!g1744) & (!g4208) & (g4212)) + ((!g1914) & (!g2599) & (!g1744) & (g4208) & (g4212)) + ((!g1914) & (!g2599) & (g1744) & (!g4208) & (g4212)) + ((!g1914) & (!g2599) & (g1744) & (g4208) & (g4212)) + ((!g1914) & (g2599) & (!g1744) & (!g4208) & (g4212)) + ((!g1914) & (g2599) & (!g1744) & (g4208) & (g4212)) + ((!g1914) & (g2599) & (g1744) & (!g4208) & (g4212)) + ((!g1914) & (g2599) & (g1744) & (g4208) & (g4212)) + ((g1914) & (!g2599) & (!g1744) & (!g4208) & (!g4212)) + ((g1914) & (!g2599) & (!g1744) & (!g4208) & (g4212)) + ((g1914) & (!g2599) & (g1744) & (g4208) & (!g4212)) + ((g1914) & (!g2599) & (g1744) & (g4208) & (g4212)) + ((g1914) & (g2599) & (!g1744) & (g4208) & (!g4212)) + ((g1914) & (g2599) & (!g1744) & (g4208) & (g4212)) + ((g1914) & (g2599) & (g1744) & (!g4208) & (!g4212)) + ((g1914) & (g2599) & (g1744) & (!g4208) & (g4212)));
	assign g4214 = (((!g830) & (!g2071) & (!g4213) & (key[2])) + ((!g830) & (!g2071) & (g4213) & (key[2])) + ((!g830) & (g2071) & (!g4213) & (key[2])) + ((!g830) & (g2071) & (g4213) & (key[2])) + ((g830) & (!g2071) & (g4213) & (!key[2])) + ((g830) & (!g2071) & (g4213) & (key[2])) + ((g830) & (g2071) & (!g4213) & (!key[2])) + ((g830) & (g2071) & (!g4213) & (key[2])));
	assign g4215 = (((!g2262) & (g2900)) + ((g2262) & (!g2900)));
	assign g4216 = (((!g2180) & (!g2212) & (g2827) & (g2851) & (!g3666) & (g4215)) + ((!g2180) & (g2212) & (!g2827) & (g2851) & (!g3666) & (g4215)) + ((!g2180) & (g2212) & (!g2827) & (g2851) & (g3666) & (g4215)) + ((!g2180) & (g2212) & (g2827) & (!g2851) & (!g3666) & (g4215)) + ((!g2180) & (g2212) & (g2827) & (g2851) & (!g3666) & (g4215)) + ((!g2180) & (g2212) & (g2827) & (g2851) & (g3666) & (g4215)) + ((g2180) & (!g2212) & (!g2827) & (g2851) & (!g3666) & (g4215)) + ((g2180) & (!g2212) & (g2827) & (g2851) & (!g3666) & (g4215)) + ((g2180) & (!g2212) & (g2827) & (g2851) & (g3666) & (g4215)) + ((g2180) & (g2212) & (!g2827) & (!g2851) & (!g3666) & (g4215)) + ((g2180) & (g2212) & (!g2827) & (g2851) & (!g3666) & (g4215)) + ((g2180) & (g2212) & (!g2827) & (g2851) & (g3666) & (g4215)) + ((g2180) & (g2212) & (g2827) & (!g2851) & (!g3666) & (g4215)) + ((g2180) & (g2212) & (g2827) & (!g2851) & (g3666) & (g4215)) + ((g2180) & (g2212) & (g2827) & (g2851) & (!g3666) & (g4215)) + ((g2180) & (g2212) & (g2827) & (g2851) & (g3666) & (g4215)));
	assign g4217 = (((g2262) & (g2900)));
	assign g4218 = (((!g2298) & (!g2944) & (!g4216) & (g4217)) + ((!g2298) & (!g2944) & (g4216) & (!g4217)) + ((!g2298) & (!g2944) & (g4216) & (g4217)) + ((!g2298) & (g2944) & (!g4216) & (!g4217)) + ((g2298) & (!g2944) & (!g4216) & (!g4217)) + ((g2298) & (g2944) & (!g4216) & (g4217)) + ((g2298) & (g2944) & (g4216) & (!g4217)) + ((g2298) & (g2944) & (g4216) & (g4217)));
	assign g4219 = (((!g4124) & (!g4125) & (!g3159) & (!g3163)) + ((!g4124) & (!g4125) & (!g3159) & (g3163)) + ((!g4124) & (!g4125) & (g3159) & (!g3163)) + ((!g4124) & (g4125) & (!g3159) & (!g3163)) + ((g4124) & (!g4125) & (!g3159) & (!g3163)) + ((g4124) & (g4125) & (!g3159) & (!g3163)));
	assign g4220 = (((!g1914) & (!g3199) & (!g4218) & (!g4219) & (!g3177)) + ((!g1914) & (!g3199) & (!g4218) & (g4219) & (g3177)) + ((!g1914) & (!g3199) & (g4218) & (!g4219) & (!g3177)) + ((!g1914) & (!g3199) & (g4218) & (g4219) & (g3177)) + ((!g1914) & (g3199) & (!g4218) & (!g4219) & (g3177)) + ((!g1914) & (g3199) & (!g4218) & (g4219) & (!g3177)) + ((!g1914) & (g3199) & (g4218) & (!g4219) & (g3177)) + ((!g1914) & (g3199) & (g4218) & (g4219) & (!g3177)) + ((g1914) & (!g3199) & (g4218) & (!g4219) & (!g3177)) + ((g1914) & (!g3199) & (g4218) & (!g4219) & (g3177)) + ((g1914) & (!g3199) & (g4218) & (g4219) & (!g3177)) + ((g1914) & (!g3199) & (g4218) & (g4219) & (g3177)) + ((g1914) & (g3199) & (g4218) & (!g4219) & (!g3177)) + ((g1914) & (g3199) & (g4218) & (!g4219) & (g3177)) + ((g1914) & (g3199) & (g4218) & (g4219) & (!g3177)) + ((g1914) & (g3199) & (g4218) & (g4219) & (g3177)));
	assign g8294 = (((!g5560) & (g5587) & (!g4221)) + ((!g5560) & (g5587) & (g4221)) + ((g5560) & (!g5587) & (g4221)) + ((g5560) & (g5587) & (g4221)));
	assign g4222 = (((!g830) & (!g2074) & (!g4220) & (g4221)) + ((!g830) & (!g2074) & (g4220) & (g4221)) + ((!g830) & (g2074) & (!g4220) & (g4221)) + ((!g830) & (g2074) & (g4220) & (g4221)) + ((g830) & (!g2074) & (g4220) & (!g4221)) + ((g830) & (!g2074) & (g4220) & (g4221)) + ((g830) & (g2074) & (!g4220) & (!g4221)) + ((g830) & (g2074) & (!g4220) & (g4221)));
	assign g4223 = (((!g2468) & (!g2486) & (!g3695) & (!g3696) & (!g5771) & (g5772)) + ((!g2468) & (!g2486) & (!g3695) & (g3696) & (!g5771) & (g5772)) + ((!g2468) & (!g2486) & (g3695) & (!g3696) & (!g5771) & (g5772)) + ((!g2468) & (!g2486) & (g3695) & (g3696) & (!g5771) & (g5772)) + ((!g2468) & (g2486) & (!g3695) & (!g3696) & (!g5771) & (g5772)) + ((!g2468) & (g2486) & (!g3695) & (g3696) & (!g5771) & (g5772)) + ((!g2468) & (g2486) & (!g3695) & (g3696) & (g5771) & (g5772)) + ((!g2468) & (g2486) & (g3695) & (!g3696) & (!g5771) & (g5772)) + ((!g2468) & (g2486) & (g3695) & (!g3696) & (g5771) & (g5772)) + ((!g2468) & (g2486) & (g3695) & (g3696) & (!g5771) & (g5772)) + ((!g2468) & (g2486) & (g3695) & (g3696) & (g5771) & (g5772)) + ((g2468) & (!g2486) & (!g3695) & (!g3696) & (!g5771) & (g5772)) + ((g2468) & (!g2486) & (!g3695) & (g3696) & (!g5771) & (g5772)) + ((g2468) & (!g2486) & (!g3695) & (g3696) & (g5771) & (g5772)) + ((g2468) & (!g2486) & (g3695) & (!g3696) & (!g5771) & (g5772)) + ((g2468) & (!g2486) & (g3695) & (!g3696) & (g5771) & (g5772)) + ((g2468) & (!g2486) & (g3695) & (g3696) & (!g5771) & (g5772)) + ((g2468) & (!g2486) & (g3695) & (g3696) & (g5771) & (g5772)) + ((g2468) & (g2486) & (!g3695) & (!g3696) & (!g5771) & (g5772)) + ((g2468) & (g2486) & (!g3695) & (!g3696) & (g5771) & (g5772)) + ((g2468) & (g2486) & (!g3695) & (g3696) & (!g5771) & (g5772)) + ((g2468) & (g2486) & (!g3695) & (g3696) & (g5771) & (g5772)) + ((g2468) & (g2486) & (g3695) & (!g3696) & (!g5771) & (g5772)) + ((g2468) & (g2486) & (g3695) & (!g3696) & (g5771) & (g5772)) + ((g2468) & (g2486) & (g3695) & (g3696) & (!g5771) & (g5772)) + ((g2468) & (g2486) & (g3695) & (g3696) & (g5771) & (g5772)));
	assign g4224 = (((g2663) & (g2669)));
	assign g4225 = (((!g4223) & (g4224)) + ((g4223) & (!g4224)) + ((g4223) & (g4224)));
	assign g4226 = (((!g2653) & (!g2718) & (!g2674) & (g2733) & (!g4148)) + ((!g2653) & (!g2718) & (!g2674) & (g2733) & (g4148)) + ((!g2653) & (!g2718) & (g2674) & (!g2733) & (g4148)) + ((!g2653) & (!g2718) & (g2674) & (g2733) & (!g4148)) + ((!g2653) & (g2718) & (!g2674) & (!g2733) & (!g4148)) + ((!g2653) & (g2718) & (!g2674) & (!g2733) & (g4148)) + ((!g2653) & (g2718) & (g2674) & (!g2733) & (!g4148)) + ((!g2653) & (g2718) & (g2674) & (g2733) & (g4148)) + ((g2653) & (!g2718) & (!g2674) & (!g2733) & (g4148)) + ((g2653) & (!g2718) & (!g2674) & (g2733) & (!g4148)) + ((g2653) & (!g2718) & (g2674) & (!g2733) & (!g4148)) + ((g2653) & (!g2718) & (g2674) & (!g2733) & (g4148)) + ((g2653) & (g2718) & (!g2674) & (!g2733) & (!g4148)) + ((g2653) & (g2718) & (!g2674) & (g2733) & (g4148)) + ((g2653) & (g2718) & (g2674) & (g2733) & (!g4148)) + ((g2653) & (g2718) & (g2674) & (g2733) & (g4148)));
	assign g4227 = (((!g2427) & (!g2519) & (!g3097) & (g3142) & (!g4160)) + ((!g2427) & (!g2519) & (!g3097) & (g3142) & (g4160)) + ((!g2427) & (!g2519) & (g3097) & (!g3142) & (g4160)) + ((!g2427) & (!g2519) & (g3097) & (g3142) & (!g4160)) + ((!g2427) & (g2519) & (!g3097) & (!g3142) & (!g4160)) + ((!g2427) & (g2519) & (!g3097) & (!g3142) & (g4160)) + ((!g2427) & (g2519) & (g3097) & (!g3142) & (!g4160)) + ((!g2427) & (g2519) & (g3097) & (g3142) & (g4160)) + ((g2427) & (!g2519) & (!g3097) & (!g3142) & (g4160)) + ((g2427) & (!g2519) & (!g3097) & (g3142) & (!g4160)) + ((g2427) & (!g2519) & (g3097) & (!g3142) & (!g4160)) + ((g2427) & (!g2519) & (g3097) & (!g3142) & (g4160)) + ((g2427) & (g2519) & (!g3097) & (!g3142) & (!g4160)) + ((g2427) & (g2519) & (!g3097) & (g3142) & (g4160)) + ((g2427) & (g2519) & (g3097) & (g3142) & (!g4160)) + ((g2427) & (g2519) & (g3097) & (g3142) & (g4160)));
	assign g4228 = (((!g3088) & (!g3128) & (!g3086) & (g3116) & (!g4162)) + ((!g3088) & (!g3128) & (!g3086) & (g3116) & (g4162)) + ((!g3088) & (!g3128) & (g3086) & (!g3116) & (g4162)) + ((!g3088) & (!g3128) & (g3086) & (g3116) & (!g4162)) + ((!g3088) & (g3128) & (!g3086) & (!g3116) & (!g4162)) + ((!g3088) & (g3128) & (!g3086) & (!g3116) & (g4162)) + ((!g3088) & (g3128) & (g3086) & (!g3116) & (!g4162)) + ((!g3088) & (g3128) & (g3086) & (g3116) & (g4162)) + ((g3088) & (!g3128) & (!g3086) & (!g3116) & (g4162)) + ((g3088) & (!g3128) & (!g3086) & (g3116) & (!g4162)) + ((g3088) & (!g3128) & (g3086) & (!g3116) & (!g4162)) + ((g3088) & (!g3128) & (g3086) & (!g3116) & (g4162)) + ((g3088) & (g3128) & (!g3086) & (!g3116) & (!g4162)) + ((g3088) & (g3128) & (!g3086) & (g3116) & (g4162)) + ((g3088) & (g3128) & (g3086) & (g3116) & (!g4162)) + ((g3088) & (g3128) & (g3086) & (g3116) & (g4162)));
	assign g4229 = (((!g830) & (!g1914) & (!g2080) & (!g4227) & (!g4228) & (key[194])) + ((!g830) & (!g1914) & (!g2080) & (!g4227) & (g4228) & (key[194])) + ((!g830) & (!g1914) & (!g2080) & (g4227) & (!g4228) & (key[194])) + ((!g830) & (!g1914) & (!g2080) & (g4227) & (g4228) & (key[194])) + ((!g830) & (!g1914) & (g2080) & (!g4227) & (!g4228) & (key[194])) + ((!g830) & (!g1914) & (g2080) & (!g4227) & (g4228) & (key[194])) + ((!g830) & (!g1914) & (g2080) & (g4227) & (!g4228) & (key[194])) + ((!g830) & (!g1914) & (g2080) & (g4227) & (g4228) & (key[194])) + ((!g830) & (g1914) & (!g2080) & (!g4227) & (!g4228) & (key[194])) + ((!g830) & (g1914) & (!g2080) & (!g4227) & (g4228) & (key[194])) + ((!g830) & (g1914) & (!g2080) & (g4227) & (!g4228) & (key[194])) + ((!g830) & (g1914) & (!g2080) & (g4227) & (g4228) & (key[194])) + ((!g830) & (g1914) & (g2080) & (!g4227) & (!g4228) & (key[194])) + ((!g830) & (g1914) & (g2080) & (!g4227) & (g4228) & (key[194])) + ((!g830) & (g1914) & (g2080) & (g4227) & (!g4228) & (key[194])) + ((!g830) & (g1914) & (g2080) & (g4227) & (g4228) & (key[194])) + ((g830) & (!g1914) & (!g2080) & (!g4227) & (g4228) & (!key[194])) + ((g830) & (!g1914) & (!g2080) & (!g4227) & (g4228) & (key[194])) + ((g830) & (!g1914) & (!g2080) & (g4227) & (g4228) & (!key[194])) + ((g830) & (!g1914) & (!g2080) & (g4227) & (g4228) & (key[194])) + ((g830) & (!g1914) & (g2080) & (!g4227) & (!g4228) & (!key[194])) + ((g830) & (!g1914) & (g2080) & (!g4227) & (!g4228) & (key[194])) + ((g830) & (!g1914) & (g2080) & (g4227) & (!g4228) & (!key[194])) + ((g830) & (!g1914) & (g2080) & (g4227) & (!g4228) & (key[194])) + ((g830) & (g1914) & (!g2080) & (g4227) & (!g4228) & (!key[194])) + ((g830) & (g1914) & (!g2080) & (g4227) & (!g4228) & (key[194])) + ((g830) & (g1914) & (!g2080) & (g4227) & (g4228) & (!key[194])) + ((g830) & (g1914) & (!g2080) & (g4227) & (g4228) & (key[194])) + ((g830) & (g1914) & (g2080) & (!g4227) & (!g4228) & (!key[194])) + ((g830) & (g1914) & (g2080) & (!g4227) & (!g4228) & (key[194])) + ((g830) & (g1914) & (g2080) & (!g4227) & (g4228) & (!key[194])) + ((g830) & (g1914) & (g2080) & (!g4227) & (g4228) & (key[194])));
	assign g4230 = (((!g4130) & (!g4131) & (!g3153) & (!g3161)) + ((!g4130) & (!g4131) & (!g3153) & (g3161)) + ((!g4130) & (!g4131) & (g3153) & (!g3161)) + ((!g4130) & (g4131) & (!g3153) & (!g3161)) + ((g4130) & (!g4131) & (!g3153) & (!g3161)) + ((g4130) & (g4131) & (!g3153) & (!g3161)));
	assign g4231 = (((!g2257) & (g2902)) + ((g2257) & (!g2902)));
	assign g4232 = (((!g2178) & (!g2211) & (g2830) & (g2863) & (!g3807) & (g4231)) + ((!g2178) & (g2211) & (!g2830) & (g2863) & (!g3807) & (g4231)) + ((!g2178) & (g2211) & (!g2830) & (g2863) & (g3807) & (g4231)) + ((!g2178) & (g2211) & (g2830) & (!g2863) & (!g3807) & (g4231)) + ((!g2178) & (g2211) & (g2830) & (g2863) & (!g3807) & (g4231)) + ((!g2178) & (g2211) & (g2830) & (g2863) & (g3807) & (g4231)) + ((g2178) & (!g2211) & (!g2830) & (g2863) & (!g3807) & (g4231)) + ((g2178) & (!g2211) & (g2830) & (g2863) & (!g3807) & (g4231)) + ((g2178) & (!g2211) & (g2830) & (g2863) & (g3807) & (g4231)) + ((g2178) & (g2211) & (!g2830) & (!g2863) & (!g3807) & (g4231)) + ((g2178) & (g2211) & (!g2830) & (g2863) & (!g3807) & (g4231)) + ((g2178) & (g2211) & (!g2830) & (g2863) & (g3807) & (g4231)) + ((g2178) & (g2211) & (g2830) & (!g2863) & (!g3807) & (g4231)) + ((g2178) & (g2211) & (g2830) & (!g2863) & (g3807) & (g4231)) + ((g2178) & (g2211) & (g2830) & (g2863) & (!g3807) & (g4231)) + ((g2178) & (g2211) & (g2830) & (g2863) & (g3807) & (g4231)));
	assign g4233 = (((g2257) & (g2902)));
	assign g4234 = (((!g2296) & (!g2968) & (!g4232) & (g4233)) + ((!g2296) & (!g2968) & (g4232) & (!g4233)) + ((!g2296) & (!g2968) & (g4232) & (g4233)) + ((!g2296) & (g2968) & (!g4232) & (!g4233)) + ((g2296) & (!g2968) & (!g4232) & (!g4233)) + ((g2296) & (g2968) & (!g4232) & (g4233)) + ((g2296) & (g2968) & (g4232) & (!g4233)) + ((g2296) & (g2968) & (g4232) & (g4233)));
	assign g4235 = (((!g1914) & (!g3184) & (!g4230) & (!g3187) & (g4234)) + ((!g1914) & (!g3184) & (!g4230) & (g3187) & (g4234)) + ((!g1914) & (!g3184) & (g4230) & (!g3187) & (g4234)) + ((!g1914) & (!g3184) & (g4230) & (g3187) & (g4234)) + ((!g1914) & (g3184) & (!g4230) & (!g3187) & (g4234)) + ((!g1914) & (g3184) & (!g4230) & (g3187) & (g4234)) + ((!g1914) & (g3184) & (g4230) & (!g3187) & (g4234)) + ((!g1914) & (g3184) & (g4230) & (g3187) & (g4234)) + ((g1914) & (!g3184) & (!g4230) & (!g3187) & (!g4234)) + ((g1914) & (!g3184) & (!g4230) & (!g3187) & (g4234)) + ((g1914) & (!g3184) & (g4230) & (g3187) & (!g4234)) + ((g1914) & (!g3184) & (g4230) & (g3187) & (g4234)) + ((g1914) & (g3184) & (!g4230) & (g3187) & (!g4234)) + ((g1914) & (g3184) & (!g4230) & (g3187) & (g4234)) + ((g1914) & (g3184) & (g4230) & (!g3187) & (!g4234)) + ((g1914) & (g3184) & (g4230) & (!g3187) & (g4234)));
	assign g4236 = (((!g830) & (!g2085) & (!g4235) & (key[130])) + ((!g830) & (!g2085) & (g4235) & (key[130])) + ((!g830) & (g2085) & (!g4235) & (key[130])) + ((!g830) & (g2085) & (g4235) & (key[130])) + ((g830) & (!g2085) & (g4235) & (!key[130])) + ((g830) & (!g2085) & (g4235) & (key[130])) + ((g830) & (g2085) & (!g4235) & (!key[130])) + ((g830) & (g2085) & (!g4235) & (key[130])));
	assign g4237 = (((!g3088) & (!g3128) & (!g3080) & (g3125) & (!g4149)) + ((!g3088) & (!g3128) & (!g3080) & (g3125) & (g4149)) + ((!g3088) & (!g3128) & (g3080) & (!g3125) & (g4149)) + ((!g3088) & (!g3128) & (g3080) & (g3125) & (!g4149)) + ((!g3088) & (g3128) & (!g3080) & (!g3125) & (!g4149)) + ((!g3088) & (g3128) & (!g3080) & (!g3125) & (g4149)) + ((!g3088) & (g3128) & (g3080) & (!g3125) & (!g4149)) + ((!g3088) & (g3128) & (g3080) & (g3125) & (g4149)) + ((g3088) & (!g3128) & (!g3080) & (!g3125) & (g4149)) + ((g3088) & (!g3128) & (!g3080) & (g3125) & (!g4149)) + ((g3088) & (!g3128) & (g3080) & (!g3125) & (!g4149)) + ((g3088) & (!g3128) & (g3080) & (!g3125) & (g4149)) + ((g3088) & (g3128) & (!g3080) & (!g3125) & (!g4149)) + ((g3088) & (g3128) & (!g3080) & (g3125) & (g4149)) + ((g3088) & (g3128) & (g3080) & (g3125) & (!g4149)) + ((g3088) & (g3128) & (g3080) & (g3125) & (g4149)));
	assign g4238 = (((!g2424) & (!g2516) & (!g3097) & (g3142) & (!g4151)) + ((!g2424) & (!g2516) & (!g3097) & (g3142) & (g4151)) + ((!g2424) & (!g2516) & (g3097) & (!g3142) & (g4151)) + ((!g2424) & (!g2516) & (g3097) & (g3142) & (!g4151)) + ((!g2424) & (g2516) & (!g3097) & (!g3142) & (!g4151)) + ((!g2424) & (g2516) & (!g3097) & (!g3142) & (g4151)) + ((!g2424) & (g2516) & (g3097) & (!g3142) & (!g4151)) + ((!g2424) & (g2516) & (g3097) & (g3142) & (g4151)) + ((g2424) & (!g2516) & (!g3097) & (!g3142) & (g4151)) + ((g2424) & (!g2516) & (!g3097) & (g3142) & (!g4151)) + ((g2424) & (!g2516) & (g3097) & (!g3142) & (!g4151)) + ((g2424) & (!g2516) & (g3097) & (!g3142) & (g4151)) + ((g2424) & (g2516) & (!g3097) & (!g3142) & (!g4151)) + ((g2424) & (g2516) & (!g3097) & (g3142) & (g4151)) + ((g2424) & (g2516) & (g3097) & (g3142) & (!g4151)) + ((g2424) & (g2516) & (g3097) & (g3142) & (g4151)));
	assign g4239 = (((!g830) & (!g1914) & (!g2088) & (!g4237) & (!g4238) & (nonce[34])) + ((!g830) & (!g1914) & (!g2088) & (!g4237) & (g4238) & (nonce[34])) + ((!g830) & (!g1914) & (!g2088) & (g4237) & (!g4238) & (nonce[34])) + ((!g830) & (!g1914) & (!g2088) & (g4237) & (g4238) & (nonce[34])) + ((!g830) & (!g1914) & (g2088) & (!g4237) & (!g4238) & (nonce[34])) + ((!g830) & (!g1914) & (g2088) & (!g4237) & (g4238) & (nonce[34])) + ((!g830) & (!g1914) & (g2088) & (g4237) & (!g4238) & (nonce[34])) + ((!g830) & (!g1914) & (g2088) & (g4237) & (g4238) & (nonce[34])) + ((!g830) & (g1914) & (!g2088) & (!g4237) & (!g4238) & (nonce[34])) + ((!g830) & (g1914) & (!g2088) & (!g4237) & (g4238) & (nonce[34])) + ((!g830) & (g1914) & (!g2088) & (g4237) & (!g4238) & (nonce[34])) + ((!g830) & (g1914) & (!g2088) & (g4237) & (g4238) & (nonce[34])) + ((!g830) & (g1914) & (g2088) & (!g4237) & (!g4238) & (nonce[34])) + ((!g830) & (g1914) & (g2088) & (!g4237) & (g4238) & (nonce[34])) + ((!g830) & (g1914) & (g2088) & (g4237) & (!g4238) & (nonce[34])) + ((!g830) & (g1914) & (g2088) & (g4237) & (g4238) & (nonce[34])) + ((g830) & (!g1914) & (!g2088) & (!g4237) & (g4238) & (!nonce[34])) + ((g830) & (!g1914) & (!g2088) & (!g4237) & (g4238) & (nonce[34])) + ((g830) & (!g1914) & (!g2088) & (g4237) & (g4238) & (!nonce[34])) + ((g830) & (!g1914) & (!g2088) & (g4237) & (g4238) & (nonce[34])) + ((g830) & (!g1914) & (g2088) & (!g4237) & (!g4238) & (!nonce[34])) + ((g830) & (!g1914) & (g2088) & (!g4237) & (!g4238) & (nonce[34])) + ((g830) & (!g1914) & (g2088) & (g4237) & (!g4238) & (!nonce[34])) + ((g830) & (!g1914) & (g2088) & (g4237) & (!g4238) & (nonce[34])) + ((g830) & (g1914) & (!g2088) & (g4237) & (!g4238) & (!nonce[34])) + ((g830) & (g1914) & (!g2088) & (g4237) & (!g4238) & (nonce[34])) + ((g830) & (g1914) & (!g2088) & (g4237) & (g4238) & (!nonce[34])) + ((g830) & (g1914) & (!g2088) & (g4237) & (g4238) & (nonce[34])) + ((g830) & (g1914) & (g2088) & (!g4237) & (!g4238) & (!nonce[34])) + ((g830) & (g1914) & (g2088) & (!g4237) & (!g4238) & (nonce[34])) + ((g830) & (g1914) & (g2088) & (!g4237) & (g4238) & (!nonce[34])) + ((g830) & (g1914) & (g2088) & (!g4237) & (g4238) & (nonce[34])));
	assign g4240 = (((!g2497) & (!g2503) & (!g3852) & (!g3853) & (!g5774) & (g5775)) + ((!g2497) & (!g2503) & (!g3852) & (g3853) & (!g5774) & (g5775)) + ((!g2497) & (!g2503) & (g3852) & (!g3853) & (!g5774) & (g5775)) + ((!g2497) & (!g2503) & (g3852) & (g3853) & (!g5774) & (g5775)) + ((!g2497) & (g2503) & (!g3852) & (!g3853) & (!g5774) & (g5775)) + ((!g2497) & (g2503) & (!g3852) & (g3853) & (!g5774) & (g5775)) + ((!g2497) & (g2503) & (!g3852) & (g3853) & (g5774) & (g5775)) + ((!g2497) & (g2503) & (g3852) & (!g3853) & (!g5774) & (g5775)) + ((!g2497) & (g2503) & (g3852) & (!g3853) & (g5774) & (g5775)) + ((!g2497) & (g2503) & (g3852) & (g3853) & (!g5774) & (g5775)) + ((!g2497) & (g2503) & (g3852) & (g3853) & (g5774) & (g5775)) + ((g2497) & (!g2503) & (!g3852) & (!g3853) & (!g5774) & (g5775)) + ((g2497) & (!g2503) & (!g3852) & (g3853) & (!g5774) & (g5775)) + ((g2497) & (!g2503) & (!g3852) & (g3853) & (g5774) & (g5775)) + ((g2497) & (!g2503) & (g3852) & (!g3853) & (!g5774) & (g5775)) + ((g2497) & (!g2503) & (g3852) & (!g3853) & (g5774) & (g5775)) + ((g2497) & (!g2503) & (g3852) & (g3853) & (!g5774) & (g5775)) + ((g2497) & (!g2503) & (g3852) & (g3853) & (g5774) & (g5775)) + ((g2497) & (g2503) & (!g3852) & (!g3853) & (!g5774) & (g5775)) + ((g2497) & (g2503) & (!g3852) & (!g3853) & (g5774) & (g5775)) + ((g2497) & (g2503) & (!g3852) & (g3853) & (!g5774) & (g5775)) + ((g2497) & (g2503) & (!g3852) & (g3853) & (g5774) & (g5775)) + ((g2497) & (g2503) & (g3852) & (!g3853) & (!g5774) & (g5775)) + ((g2497) & (g2503) & (g3852) & (!g3853) & (g5774) & (g5775)) + ((g2497) & (g2503) & (g3852) & (g3853) & (!g5774) & (g5775)) + ((g2497) & (g2503) & (g3852) & (g3853) & (g5774) & (g5775)));
	assign g4241 = (((g2672) & (g2674)));
	assign g4242 = (((!g4240) & (g4241)) + ((g4240) & (!g4241)) + ((g4240) & (g4241)));
	assign g4243 = (((!g2661) & (!g2742) & (!g2669) & (g2747) & (!g4166)) + ((!g2661) & (!g2742) & (!g2669) & (g2747) & (g4166)) + ((!g2661) & (!g2742) & (g2669) & (!g2747) & (g4166)) + ((!g2661) & (!g2742) & (g2669) & (g2747) & (!g4166)) + ((!g2661) & (g2742) & (!g2669) & (!g2747) & (!g4166)) + ((!g2661) & (g2742) & (!g2669) & (!g2747) & (g4166)) + ((!g2661) & (g2742) & (g2669) & (!g2747) & (!g4166)) + ((!g2661) & (g2742) & (g2669) & (g2747) & (g4166)) + ((g2661) & (!g2742) & (!g2669) & (!g2747) & (g4166)) + ((g2661) & (!g2742) & (!g2669) & (g2747) & (!g4166)) + ((g2661) & (!g2742) & (g2669) & (!g2747) & (!g4166)) + ((g2661) & (!g2742) & (g2669) & (!g2747) & (g4166)) + ((g2661) & (g2742) & (!g2669) & (!g2747) & (!g4166)) + ((g2661) & (g2742) & (!g2669) & (g2747) & (g4166)) + ((g2661) & (g2742) & (g2669) & (g2747) & (!g4166)) + ((g2661) & (g2742) & (g2669) & (g2747) & (g4166)));
	assign g4244 = (((!g1031) & (!g1065) & (!g4167) & (!g2233) & (g2267)) + ((!g1031) & (!g1065) & (!g4167) & (g2233) & (!g2267)) + ((!g1031) & (!g1065) & (g4167) & (!g2233) & (g2267)) + ((!g1031) & (!g1065) & (g4167) & (g2233) & (g2267)) + ((!g1031) & (g1065) & (!g4167) & (!g2233) & (!g2267)) + ((!g1031) & (g1065) & (!g4167) & (g2233) & (g2267)) + ((!g1031) & (g1065) & (g4167) & (!g2233) & (!g2267)) + ((!g1031) & (g1065) & (g4167) & (g2233) & (!g2267)) + ((g1031) & (!g1065) & (!g4167) & (!g2233) & (!g2267)) + ((g1031) & (!g1065) & (!g4167) & (g2233) & (!g2267)) + ((g1031) & (!g1065) & (g4167) & (!g2233) & (g2267)) + ((g1031) & (!g1065) & (g4167) & (g2233) & (!g2267)) + ((g1031) & (g1065) & (!g4167) & (!g2233) & (g2267)) + ((g1031) & (g1065) & (!g4167) & (g2233) & (g2267)) + ((g1031) & (g1065) & (g4167) & (!g2233) & (!g2267)) + ((g1031) & (g1065) & (g4167) & (g2233) & (g2267)));
	assign g4245 = (((!g2224) & (!g2271) & (!g2230) & (g2286) & (!g4169)) + ((!g2224) & (!g2271) & (!g2230) & (g2286) & (g4169)) + ((!g2224) & (!g2271) & (g2230) & (!g2286) & (!g4169)) + ((!g2224) & (!g2271) & (g2230) & (g2286) & (g4169)) + ((!g2224) & (g2271) & (!g2230) & (!g2286) & (!g4169)) + ((!g2224) & (g2271) & (!g2230) & (!g2286) & (g4169)) + ((!g2224) & (g2271) & (g2230) & (!g2286) & (g4169)) + ((!g2224) & (g2271) & (g2230) & (g2286) & (!g4169)) + ((g2224) & (!g2271) & (!g2230) & (!g2286) & (!g4169)) + ((g2224) & (!g2271) & (!g2230) & (g2286) & (g4169)) + ((g2224) & (!g2271) & (g2230) & (!g2286) & (!g4169)) + ((g2224) & (!g2271) & (g2230) & (!g2286) & (g4169)) + ((g2224) & (g2271) & (!g2230) & (!g2286) & (g4169)) + ((g2224) & (g2271) & (!g2230) & (g2286) & (!g4169)) + ((g2224) & (g2271) & (g2230) & (g2286) & (!g4169)) + ((g2224) & (g2271) & (g2230) & (g2286) & (g4169)));
	assign g4246 = (((!g830) & (!g1914) & (!g2098) & (!g4244) & (!g4245) & (key[48])) + ((!g830) & (!g1914) & (!g2098) & (!g4244) & (g4245) & (key[48])) + ((!g830) & (!g1914) & (!g2098) & (g4244) & (!g4245) & (key[48])) + ((!g830) & (!g1914) & (!g2098) & (g4244) & (g4245) & (key[48])) + ((!g830) & (!g1914) & (g2098) & (!g4244) & (!g4245) & (key[48])) + ((!g830) & (!g1914) & (g2098) & (!g4244) & (g4245) & (key[48])) + ((!g830) & (!g1914) & (g2098) & (g4244) & (!g4245) & (key[48])) + ((!g830) & (!g1914) & (g2098) & (g4244) & (g4245) & (key[48])) + ((!g830) & (g1914) & (!g2098) & (!g4244) & (!g4245) & (key[48])) + ((!g830) & (g1914) & (!g2098) & (!g4244) & (g4245) & (key[48])) + ((!g830) & (g1914) & (!g2098) & (g4244) & (!g4245) & (key[48])) + ((!g830) & (g1914) & (!g2098) & (g4244) & (g4245) & (key[48])) + ((!g830) & (g1914) & (g2098) & (!g4244) & (!g4245) & (key[48])) + ((!g830) & (g1914) & (g2098) & (!g4244) & (g4245) & (key[48])) + ((!g830) & (g1914) & (g2098) & (g4244) & (!g4245) & (key[48])) + ((!g830) & (g1914) & (g2098) & (g4244) & (g4245) & (key[48])) + ((g830) & (!g1914) & (!g2098) & (!g4244) & (g4245) & (!key[48])) + ((g830) & (!g1914) & (!g2098) & (!g4244) & (g4245) & (key[48])) + ((g830) & (!g1914) & (!g2098) & (g4244) & (g4245) & (!key[48])) + ((g830) & (!g1914) & (!g2098) & (g4244) & (g4245) & (key[48])) + ((g830) & (!g1914) & (g2098) & (!g4244) & (!g4245) & (!key[48])) + ((g830) & (!g1914) & (g2098) & (!g4244) & (!g4245) & (key[48])) + ((g830) & (!g1914) & (g2098) & (g4244) & (!g4245) & (!key[48])) + ((g830) & (!g1914) & (g2098) & (g4244) & (!g4245) & (key[48])) + ((g830) & (g1914) & (!g2098) & (g4244) & (!g4245) & (!key[48])) + ((g830) & (g1914) & (!g2098) & (g4244) & (!g4245) & (key[48])) + ((g830) & (g1914) & (!g2098) & (g4244) & (g4245) & (!key[48])) + ((g830) & (g1914) & (!g2098) & (g4244) & (g4245) & (key[48])) + ((g830) & (g1914) & (g2098) & (!g4244) & (!g4245) & (!key[48])) + ((g830) & (g1914) & (g2098) & (!g4244) & (!g4245) & (key[48])) + ((g830) & (g1914) & (g2098) & (!g4244) & (g4245) & (!key[48])) + ((g830) & (g1914) & (g2098) & (!g4244) & (g4245) & (key[48])));
	assign g4247 = (((!g2334) & (g2340) & (!g3763)) + ((g2334) & (!g2340) & (!g3763)) + ((g2334) & (g2340) & (!g3763)) + ((g2334) & (g2340) & (g3763)));
	assign g4248 = (((!g1944) & (!g2104) & (g3745)) + ((!g1944) & (g2104) & (!g3745)) + ((g1944) & (!g2104) & (!g3745)) + ((g1944) & (g2104) & (g3745)));
	assign g4249 = (((!g1914) & (!g2358) & (!g2373) & (g4247) & (!g4248)) + ((!g1914) & (!g2358) & (!g2373) & (g4247) & (g4248)) + ((!g1914) & (!g2358) & (g2373) & (!g4247) & (!g4248)) + ((!g1914) & (!g2358) & (g2373) & (!g4247) & (g4248)) + ((!g1914) & (g2358) & (!g2373) & (!g4247) & (!g4248)) + ((!g1914) & (g2358) & (!g2373) & (!g4247) & (g4248)) + ((!g1914) & (g2358) & (g2373) & (g4247) & (!g4248)) + ((!g1914) & (g2358) & (g2373) & (g4247) & (g4248)) + ((g1914) & (!g2358) & (!g2373) & (!g4247) & (g4248)) + ((g1914) & (!g2358) & (!g2373) & (g4247) & (g4248)) + ((g1914) & (!g2358) & (g2373) & (!g4247) & (g4248)) + ((g1914) & (!g2358) & (g2373) & (g4247) & (g4248)) + ((g1914) & (g2358) & (!g2373) & (!g4247) & (g4248)) + ((g1914) & (g2358) & (!g2373) & (g4247) & (g4248)) + ((g1914) & (g2358) & (g2373) & (!g4247) & (g4248)) + ((g1914) & (g2358) & (g2373) & (g4247) & (g4248)));
	assign g4250 = (((!g830) & (!g2099) & (!g4249) & (key[80])) + ((!g830) & (!g2099) & (g4249) & (key[80])) + ((!g830) & (g2099) & (!g4249) & (key[80])) + ((!g830) & (g2099) & (g4249) & (key[80])) + ((g830) & (!g2099) & (g4249) & (!key[80])) + ((g830) & (!g2099) & (g4249) & (key[80])) + ((g830) & (g2099) & (!g4249) & (!key[80])) + ((g830) & (g2099) & (!g4249) & (key[80])));
	assign g4251 = (((!g4176) & (!g2224) & (!g2247) & (!g2271) & (g2275)) + ((!g4176) & (!g2224) & (!g2247) & (g2271) & (!g2275)) + ((!g4176) & (!g2224) & (g2247) & (!g2271) & (g2275)) + ((!g4176) & (!g2224) & (g2247) & (g2271) & (!g2275)) + ((!g4176) & (g2224) & (!g2247) & (!g2271) & (g2275)) + ((!g4176) & (g2224) & (!g2247) & (g2271) & (!g2275)) + ((!g4176) & (g2224) & (g2247) & (!g2271) & (!g2275)) + ((!g4176) & (g2224) & (g2247) & (g2271) & (g2275)) + ((g4176) & (!g2224) & (!g2247) & (!g2271) & (g2275)) + ((g4176) & (!g2224) & (!g2247) & (g2271) & (!g2275)) + ((g4176) & (!g2224) & (g2247) & (!g2271) & (!g2275)) + ((g4176) & (!g2224) & (g2247) & (g2271) & (g2275)) + ((g4176) & (g2224) & (!g2247) & (!g2271) & (!g2275)) + ((g4176) & (g2224) & (!g2247) & (g2271) & (g2275)) + ((g4176) & (g2224) & (g2247) & (!g2271) & (!g2275)) + ((g4176) & (g2224) & (g2247) & (g2271) & (g2275)));
	assign g8295 = (((!g5560) & (g5588) & (!g4252)) + ((!g5560) & (g5588) & (g4252)) + ((g5560) & (!g5588) & (g4252)) + ((g5560) & (g5588) & (g4252)));
	assign g4253 = (((!g830) & (!g2100) & (!g6830) & (g4252)) + ((!g830) & (!g2100) & (g6830) & (g4252)) + ((!g830) & (g2100) & (!g6830) & (g4252)) + ((!g830) & (g2100) & (g6830) & (g4252)) + ((g830) & (!g2100) & (g6830) & (!g4252)) + ((g830) & (!g2100) & (g6830) & (g4252)) + ((g830) & (g2100) & (!g6830) & (!g4252)) + ((g830) & (g2100) & (!g6830) & (g4252)));
	assign g4254 = (((!g3469) & (!g2317) & (g2340)) + ((!g3469) & (g2317) & (!g2340)) + ((!g3469) & (g2317) & (g2340)) + ((g3469) & (g2317) & (g2340)));
	assign g4255 = (((!g1982) & (!g2114) & (g3483)) + ((!g1982) & (g2114) & (!g3483)) + ((g1982) & (!g2114) & (!g3483)) + ((g1982) & (g2114) & (g3483)));
	assign g4256 = (((!g1914) & (!g4254) & (!g2369) & (!g2373) & (g4255)) + ((!g1914) & (!g4254) & (!g2369) & (g2373) & (g4255)) + ((!g1914) & (!g4254) & (g2369) & (!g2373) & (g4255)) + ((!g1914) & (!g4254) & (g2369) & (g2373) & (g4255)) + ((!g1914) & (g4254) & (!g2369) & (!g2373) & (g4255)) + ((!g1914) & (g4254) & (!g2369) & (g2373) & (g4255)) + ((!g1914) & (g4254) & (g2369) & (!g2373) & (g4255)) + ((!g1914) & (g4254) & (g2369) & (g2373) & (g4255)) + ((g1914) & (!g4254) & (!g2369) & (g2373) & (!g4255)) + ((g1914) & (!g4254) & (!g2369) & (g2373) & (g4255)) + ((g1914) & (!g4254) & (g2369) & (!g2373) & (!g4255)) + ((g1914) & (!g4254) & (g2369) & (!g2373) & (g4255)) + ((g1914) & (g4254) & (!g2369) & (!g2373) & (!g4255)) + ((g1914) & (g4254) & (!g2369) & (!g2373) & (g4255)) + ((g1914) & (g4254) & (g2369) & (g2373) & (!g4255)) + ((g1914) & (g4254) & (g2369) & (g2373) & (g4255)));
	assign g4257 = (((!g830) & (!g2101) & (!g4256) & (key[176])) + ((!g830) & (!g2101) & (g4256) & (key[176])) + ((!g830) & (g2101) & (!g4256) & (key[176])) + ((!g830) & (g2101) & (g4256) & (key[176])) + ((g830) & (!g2101) & (g4256) & (!key[176])) + ((g830) & (!g2101) & (g4256) & (key[176])) + ((g830) & (g2101) & (!g4256) & (!key[176])) + ((g830) & (g2101) & (!g4256) & (key[176])));
	assign g4258 = (((!g2552) & (!g2599) & (!g1711) & (!g1744) & (!g4115) & (!g4116)) + ((!g2552) & (!g2599) & (!g1711) & (!g1744) & (!g4115) & (g4116)) + ((!g2552) & (!g2599) & (!g1711) & (!g1744) & (g4115) & (!g4116)) + ((!g2552) & (!g2599) & (!g1711) & (!g1744) & (g4115) & (g4116)) + ((!g2552) & (!g2599) & (!g1711) & (g1744) & (!g4115) & (!g4116)) + ((!g2552) & (!g2599) & (!g1711) & (g1744) & (!g4115) & (g4116)) + ((!g2552) & (!g2599) & (!g1711) & (g1744) & (g4115) & (!g4116)) + ((!g2552) & (!g2599) & (!g1711) & (g1744) & (g4115) & (g4116)) + ((!g2552) & (!g2599) & (g1711) & (!g1744) & (!g4115) & (!g4116)) + ((!g2552) & (!g2599) & (g1711) & (!g1744) & (!g4115) & (g4116)) + ((!g2552) & (!g2599) & (g1711) & (!g1744) & (g4115) & (!g4116)) + ((!g2552) & (!g2599) & (g1711) & (!g1744) & (g4115) & (g4116)) + ((!g2552) & (!g2599) & (g1711) & (g1744) & (!g4115) & (!g4116)) + ((!g2552) & (g2599) & (!g1711) & (!g1744) & (!g4115) & (!g4116)) + ((!g2552) & (g2599) & (!g1711) & (!g1744) & (!g4115) & (g4116)) + ((!g2552) & (g2599) & (!g1711) & (!g1744) & (g4115) & (!g4116)) + ((!g2552) & (g2599) & (!g1711) & (!g1744) & (g4115) & (g4116)) + ((!g2552) & (g2599) & (g1711) & (!g1744) & (!g4115) & (!g4116)) + ((g2552) & (!g2599) & (!g1711) & (!g1744) & (!g4115) & (!g4116)) + ((g2552) & (!g2599) & (!g1711) & (!g1744) & (!g4115) & (g4116)) + ((g2552) & (!g2599) & (!g1711) & (!g1744) & (g4115) & (!g4116)) + ((g2552) & (!g2599) & (!g1711) & (!g1744) & (g4115) & (g4116)) + ((g2552) & (!g2599) & (!g1711) & (g1744) & (!g4115) & (!g4116)) + ((g2552) & (!g2599) & (g1711) & (!g1744) & (!g4115) & (!g4116)) + ((g2552) & (!g2599) & (g1711) & (!g1744) & (!g4115) & (g4116)) + ((g2552) & (!g2599) & (g1711) & (!g1744) & (g4115) & (!g4116)) + ((g2552) & (!g2599) & (g1711) & (!g1744) & (g4115) & (g4116)) + ((g2552) & (g2599) & (!g1711) & (!g1744) & (!g4115) & (!g4116)));
	assign g4259 = (((!g2938) & (!g3011) & (!g2985) & (!g4210) & (!g4211) & (g3015)) + ((!g2938) & (!g3011) & (!g2985) & (!g4210) & (g4211) & (g3015)) + ((!g2938) & (!g3011) & (!g2985) & (g4210) & (!g4211) & (g3015)) + ((!g2938) & (!g3011) & (!g2985) & (g4210) & (g4211) & (g3015)) + ((!g2938) & (!g3011) & (g2985) & (!g4210) & (!g4211) & (g3015)) + ((!g2938) & (!g3011) & (g2985) & (!g4210) & (g4211) & (!g3015)) + ((!g2938) & (!g3011) & (g2985) & (g4210) & (!g4211) & (!g3015)) + ((!g2938) & (!g3011) & (g2985) & (g4210) & (g4211) & (!g3015)) + ((!g2938) & (g3011) & (!g2985) & (!g4210) & (!g4211) & (!g3015)) + ((!g2938) & (g3011) & (!g2985) & (!g4210) & (g4211) & (!g3015)) + ((!g2938) & (g3011) & (!g2985) & (g4210) & (!g4211) & (!g3015)) + ((!g2938) & (g3011) & (!g2985) & (g4210) & (g4211) & (!g3015)) + ((!g2938) & (g3011) & (g2985) & (!g4210) & (!g4211) & (!g3015)) + ((!g2938) & (g3011) & (g2985) & (!g4210) & (g4211) & (g3015)) + ((!g2938) & (g3011) & (g2985) & (g4210) & (!g4211) & (g3015)) + ((!g2938) & (g3011) & (g2985) & (g4210) & (g4211) & (g3015)) + ((g2938) & (!g3011) & (!g2985) & (!g4210) & (!g4211) & (g3015)) + ((g2938) & (!g3011) & (!g2985) & (!g4210) & (g4211) & (!g3015)) + ((g2938) & (!g3011) & (!g2985) & (g4210) & (!g4211) & (!g3015)) + ((g2938) & (!g3011) & (!g2985) & (g4210) & (g4211) & (!g3015)) + ((g2938) & (!g3011) & (g2985) & (!g4210) & (!g4211) & (!g3015)) + ((g2938) & (!g3011) & (g2985) & (!g4210) & (g4211) & (!g3015)) + ((g2938) & (!g3011) & (g2985) & (g4210) & (!g4211) & (!g3015)) + ((g2938) & (!g3011) & (g2985) & (g4210) & (g4211) & (!g3015)) + ((g2938) & (g3011) & (!g2985) & (!g4210) & (!g4211) & (!g3015)) + ((g2938) & (g3011) & (!g2985) & (!g4210) & (g4211) & (g3015)) + ((g2938) & (g3011) & (!g2985) & (g4210) & (!g4211) & (g3015)) + ((g2938) & (g3011) & (!g2985) & (g4210) & (g4211) & (g3015)) + ((g2938) & (g3011) & (g2985) & (!g4210) & (!g4211) & (g3015)) + ((g2938) & (g3011) & (g2985) & (!g4210) & (g4211) & (g3015)) + ((g2938) & (g3011) & (g2985) & (g4210) & (!g4211) & (g3015)) + ((g2938) & (g3011) & (g2985) & (g4210) & (g4211) & (g3015)));
	assign g4260 = (((!g1914) & (!g2648) & (!g1778) & (!g4258) & (g4259)) + ((!g1914) & (!g2648) & (!g1778) & (g4258) & (g4259)) + ((!g1914) & (!g2648) & (g1778) & (!g4258) & (g4259)) + ((!g1914) & (!g2648) & (g1778) & (g4258) & (g4259)) + ((!g1914) & (g2648) & (!g1778) & (!g4258) & (g4259)) + ((!g1914) & (g2648) & (!g1778) & (g4258) & (g4259)) + ((!g1914) & (g2648) & (g1778) & (!g4258) & (g4259)) + ((!g1914) & (g2648) & (g1778) & (g4258) & (g4259)) + ((g1914) & (!g2648) & (!g1778) & (!g4258) & (!g4259)) + ((g1914) & (!g2648) & (!g1778) & (!g4258) & (g4259)) + ((g1914) & (!g2648) & (g1778) & (g4258) & (!g4259)) + ((g1914) & (!g2648) & (g1778) & (g4258) & (g4259)) + ((g1914) & (g2648) & (!g1778) & (g4258) & (!g4259)) + ((g1914) & (g2648) & (!g1778) & (g4258) & (g4259)) + ((g1914) & (g2648) & (g1778) & (!g4258) & (!g4259)) + ((g1914) & (g2648) & (g1778) & (!g4258) & (g4259)));
	assign g4261 = (((!g830) & (!g2104) & (!g4260) & (key[3])) + ((!g830) & (!g2104) & (g4260) & (key[3])) + ((!g830) & (g2104) & (!g4260) & (key[3])) + ((!g830) & (g2104) & (g4260) & (key[3])) + ((g830) & (!g2104) & (g4260) & (!key[3])) + ((g830) & (!g2104) & (g4260) & (key[3])) + ((g830) & (g2104) & (!g4260) & (!key[3])) + ((g830) & (g2104) & (!g4260) & (key[3])));
	assign g4262 = (((!g2100) & (!g2133) & (!g2723) & (g2770) & (!g4192)) + ((!g2100) & (!g2133) & (!g2723) & (g2770) & (g4192)) + ((!g2100) & (!g2133) & (g2723) & (!g2770) & (g4192)) + ((!g2100) & (!g2133) & (g2723) & (g2770) & (!g4192)) + ((!g2100) & (g2133) & (!g2723) & (!g2770) & (!g4192)) + ((!g2100) & (g2133) & (!g2723) & (!g2770) & (g4192)) + ((!g2100) & (g2133) & (g2723) & (!g2770) & (!g4192)) + ((!g2100) & (g2133) & (g2723) & (g2770) & (g4192)) + ((g2100) & (!g2133) & (!g2723) & (!g2770) & (g4192)) + ((g2100) & (!g2133) & (!g2723) & (g2770) & (!g4192)) + ((g2100) & (!g2133) & (g2723) & (!g2770) & (!g4192)) + ((g2100) & (!g2133) & (g2723) & (!g2770) & (g4192)) + ((g2100) & (g2133) & (!g2723) & (!g2770) & (!g4192)) + ((g2100) & (g2133) & (!g2723) & (g2770) & (g4192)) + ((g2100) & (g2133) & (g2723) & (g2770) & (!g4192)) + ((g2100) & (g2133) & (g2723) & (g2770) & (g4192)));
	assign g4263 = (((!g2047) & (!g2098) & (g2665) & (g2708) & (g4121)) + ((!g2047) & (g2098) & (!g2665) & (g2708) & (!g4121)) + ((!g2047) & (g2098) & (!g2665) & (g2708) & (g4121)) + ((!g2047) & (g2098) & (g2665) & (!g2708) & (g4121)) + ((!g2047) & (g2098) & (g2665) & (g2708) & (!g4121)) + ((!g2047) & (g2098) & (g2665) & (g2708) & (g4121)) + ((g2047) & (!g2098) & (!g2665) & (g2708) & (g4121)) + ((g2047) & (!g2098) & (g2665) & (g2708) & (!g4121)) + ((g2047) & (!g2098) & (g2665) & (g2708) & (g4121)) + ((g2047) & (g2098) & (!g2665) & (!g2708) & (g4121)) + ((g2047) & (g2098) & (!g2665) & (g2708) & (!g4121)) + ((g2047) & (g2098) & (!g2665) & (g2708) & (g4121)) + ((g2047) & (g2098) & (g2665) & (!g2708) & (!g4121)) + ((g2047) & (g2098) & (g2665) & (!g2708) & (g4121)) + ((g2047) & (g2098) & (g2665) & (g2708) & (!g4121)) + ((g2047) & (g2098) & (g2665) & (g2708) & (g4121)));
	assign g4264 = (((!g2298) & (!g2347) & (!g2944) & (g3018) & (!g4216) & (!g4217)) + ((!g2298) & (!g2347) & (!g2944) & (g3018) & (!g4216) & (g4217)) + ((!g2298) & (!g2347) & (!g2944) & (g3018) & (g4216) & (!g4217)) + ((!g2298) & (!g2347) & (!g2944) & (g3018) & (g4216) & (g4217)) + ((!g2298) & (!g2347) & (g2944) & (!g3018) & (!g4216) & (g4217)) + ((!g2298) & (!g2347) & (g2944) & (!g3018) & (g4216) & (!g4217)) + ((!g2298) & (!g2347) & (g2944) & (!g3018) & (g4216) & (g4217)) + ((!g2298) & (!g2347) & (g2944) & (g3018) & (!g4216) & (!g4217)) + ((!g2298) & (g2347) & (!g2944) & (!g3018) & (!g4216) & (!g4217)) + ((!g2298) & (g2347) & (!g2944) & (!g3018) & (!g4216) & (g4217)) + ((!g2298) & (g2347) & (!g2944) & (!g3018) & (g4216) & (!g4217)) + ((!g2298) & (g2347) & (!g2944) & (!g3018) & (g4216) & (g4217)) + ((!g2298) & (g2347) & (g2944) & (!g3018) & (!g4216) & (!g4217)) + ((!g2298) & (g2347) & (g2944) & (g3018) & (!g4216) & (g4217)) + ((!g2298) & (g2347) & (g2944) & (g3018) & (g4216) & (!g4217)) + ((!g2298) & (g2347) & (g2944) & (g3018) & (g4216) & (g4217)) + ((g2298) & (!g2347) & (!g2944) & (!g3018) & (!g4216) & (g4217)) + ((g2298) & (!g2347) & (!g2944) & (!g3018) & (g4216) & (!g4217)) + ((g2298) & (!g2347) & (!g2944) & (!g3018) & (g4216) & (g4217)) + ((g2298) & (!g2347) & (!g2944) & (g3018) & (!g4216) & (!g4217)) + ((g2298) & (!g2347) & (g2944) & (!g3018) & (!g4216) & (!g4217)) + ((g2298) & (!g2347) & (g2944) & (!g3018) & (!g4216) & (g4217)) + ((g2298) & (!g2347) & (g2944) & (!g3018) & (g4216) & (!g4217)) + ((g2298) & (!g2347) & (g2944) & (!g3018) & (g4216) & (g4217)) + ((g2298) & (g2347) & (!g2944) & (!g3018) & (!g4216) & (!g4217)) + ((g2298) & (g2347) & (!g2944) & (g3018) & (!g4216) & (g4217)) + ((g2298) & (g2347) & (!g2944) & (g3018) & (g4216) & (!g4217)) + ((g2298) & (g2347) & (!g2944) & (g3018) & (g4216) & (g4217)) + ((g2298) & (g2347) & (g2944) & (g3018) & (!g4216) & (!g4217)) + ((g2298) & (g2347) & (g2944) & (g3018) & (!g4216) & (g4217)) + ((g2298) & (g2347) & (g2944) & (g3018) & (g4216) & (!g4217)) + ((g2298) & (g2347) & (g2944) & (g3018) & (g4216) & (g4217)));
	assign g4265 = (((!g4124) & (!g4125) & (!g3159) & (!g3163) & (!g3199) & (!g3177)) + ((!g4124) & (!g4125) & (!g3159) & (!g3163) & (!g3199) & (g3177)) + ((!g4124) & (!g4125) & (!g3159) & (!g3163) & (g3199) & (!g3177)) + ((!g4124) & (!g4125) & (!g3159) & (g3163) & (!g3199) & (!g3177)) + ((!g4124) & (!g4125) & (!g3159) & (g3163) & (!g3199) & (g3177)) + ((!g4124) & (!g4125) & (!g3159) & (g3163) & (g3199) & (!g3177)) + ((!g4124) & (!g4125) & (g3159) & (!g3163) & (!g3199) & (!g3177)) + ((!g4124) & (!g4125) & (g3159) & (!g3163) & (!g3199) & (g3177)) + ((!g4124) & (!g4125) & (g3159) & (!g3163) & (g3199) & (!g3177)) + ((!g4124) & (!g4125) & (g3159) & (g3163) & (!g3199) & (!g3177)) + ((!g4124) & (g4125) & (!g3159) & (!g3163) & (!g3199) & (!g3177)) + ((!g4124) & (g4125) & (!g3159) & (!g3163) & (!g3199) & (g3177)) + ((!g4124) & (g4125) & (!g3159) & (!g3163) & (g3199) & (!g3177)) + ((!g4124) & (g4125) & (!g3159) & (g3163) & (!g3199) & (!g3177)) + ((!g4124) & (g4125) & (g3159) & (!g3163) & (!g3199) & (!g3177)) + ((!g4124) & (g4125) & (g3159) & (g3163) & (!g3199) & (!g3177)) + ((g4124) & (!g4125) & (!g3159) & (!g3163) & (!g3199) & (!g3177)) + ((g4124) & (!g4125) & (!g3159) & (!g3163) & (!g3199) & (g3177)) + ((g4124) & (!g4125) & (!g3159) & (!g3163) & (g3199) & (!g3177)) + ((g4124) & (!g4125) & (!g3159) & (g3163) & (!g3199) & (!g3177)) + ((g4124) & (!g4125) & (g3159) & (!g3163) & (!g3199) & (!g3177)) + ((g4124) & (!g4125) & (g3159) & (g3163) & (!g3199) & (!g3177)) + ((g4124) & (g4125) & (!g3159) & (!g3163) & (!g3199) & (!g3177)) + ((g4124) & (g4125) & (!g3159) & (!g3163) & (!g3199) & (g3177)) + ((g4124) & (g4125) & (!g3159) & (!g3163) & (g3199) & (!g3177)) + ((g4124) & (g4125) & (!g3159) & (g3163) & (!g3199) & (!g3177)) + ((g4124) & (g4125) & (g3159) & (!g3163) & (!g3199) & (!g3177)) + ((g4124) & (g4125) & (g3159) & (g3163) & (!g3199) & (!g3177)));
	assign g4266 = (((!g1914) & (!g4264) & (!g4265) & (!g3250) & (!g3260)) + ((!g1914) & (!g4264) & (!g4265) & (g3250) & (g3260)) + ((!g1914) & (!g4264) & (g4265) & (!g3250) & (g3260)) + ((!g1914) & (!g4264) & (g4265) & (g3250) & (!g3260)) + ((!g1914) & (g4264) & (!g4265) & (!g3250) & (!g3260)) + ((!g1914) & (g4264) & (!g4265) & (g3250) & (g3260)) + ((!g1914) & (g4264) & (g4265) & (!g3250) & (g3260)) + ((!g1914) & (g4264) & (g4265) & (g3250) & (!g3260)) + ((g1914) & (g4264) & (!g4265) & (!g3250) & (!g3260)) + ((g1914) & (g4264) & (!g4265) & (!g3250) & (g3260)) + ((g1914) & (g4264) & (!g4265) & (g3250) & (!g3260)) + ((g1914) & (g4264) & (!g4265) & (g3250) & (g3260)) + ((g1914) & (g4264) & (g4265) & (!g3250) & (!g3260)) + ((g1914) & (g4264) & (g4265) & (!g3250) & (g3260)) + ((g1914) & (g4264) & (g4265) & (g3250) & (!g3260)) + ((g1914) & (g4264) & (g4265) & (g3250) & (g3260)));
	assign g8296 = (((!g5560) & (g5589) & (!g4267)) + ((!g5560) & (g5589) & (g4267)) + ((g5560) & (!g5589) & (g4267)) + ((g5560) & (g5589) & (g4267)));
	assign g4268 = (((!g830) & (!g2110) & (!g4266) & (g4267)) + ((!g830) & (!g2110) & (g4266) & (g4267)) + ((!g830) & (g2110) & (!g4266) & (g4267)) + ((!g830) & (g2110) & (g4266) & (g4267)) + ((g830) & (!g2110) & (g4266) & (!g4267)) + ((g830) & (!g2110) & (g4266) & (g4267)) + ((g830) & (g2110) & (!g4266) & (!g4267)) + ((g830) & (g2110) & (!g4266) & (g4267)));
	assign g4269 = (((!g4130) & (!g4131) & (!g3153) & (!g3161) & (!g3184) & (!g3187)) + ((!g4130) & (!g4131) & (!g3153) & (!g3161) & (!g3184) & (g3187)) + ((!g4130) & (!g4131) & (!g3153) & (!g3161) & (g3184) & (!g3187)) + ((!g4130) & (!g4131) & (!g3153) & (g3161) & (!g3184) & (!g3187)) + ((!g4130) & (!g4131) & (!g3153) & (g3161) & (!g3184) & (g3187)) + ((!g4130) & (!g4131) & (!g3153) & (g3161) & (g3184) & (!g3187)) + ((!g4130) & (!g4131) & (g3153) & (!g3161) & (!g3184) & (!g3187)) + ((!g4130) & (!g4131) & (g3153) & (!g3161) & (!g3184) & (g3187)) + ((!g4130) & (!g4131) & (g3153) & (!g3161) & (g3184) & (!g3187)) + ((!g4130) & (!g4131) & (g3153) & (g3161) & (!g3184) & (!g3187)) + ((!g4130) & (g4131) & (!g3153) & (!g3161) & (!g3184) & (!g3187)) + ((!g4130) & (g4131) & (!g3153) & (!g3161) & (!g3184) & (g3187)) + ((!g4130) & (g4131) & (!g3153) & (!g3161) & (g3184) & (!g3187)) + ((!g4130) & (g4131) & (!g3153) & (g3161) & (!g3184) & (!g3187)) + ((!g4130) & (g4131) & (g3153) & (!g3161) & (!g3184) & (!g3187)) + ((!g4130) & (g4131) & (g3153) & (g3161) & (!g3184) & (!g3187)) + ((g4130) & (!g4131) & (!g3153) & (!g3161) & (!g3184) & (!g3187)) + ((g4130) & (!g4131) & (!g3153) & (!g3161) & (!g3184) & (g3187)) + ((g4130) & (!g4131) & (!g3153) & (!g3161) & (g3184) & (!g3187)) + ((g4130) & (!g4131) & (!g3153) & (g3161) & (!g3184) & (!g3187)) + ((g4130) & (!g4131) & (g3153) & (!g3161) & (!g3184) & (!g3187)) + ((g4130) & (!g4131) & (g3153) & (g3161) & (!g3184) & (!g3187)) + ((g4130) & (g4131) & (!g3153) & (!g3161) & (!g3184) & (!g3187)) + ((g4130) & (g4131) & (!g3153) & (!g3161) & (!g3184) & (g3187)) + ((g4130) & (g4131) & (!g3153) & (!g3161) & (g3184) & (!g3187)) + ((g4130) & (g4131) & (!g3153) & (g3161) & (!g3184) & (!g3187)) + ((g4130) & (g4131) & (g3153) & (!g3161) & (!g3184) & (!g3187)) + ((g4130) & (g4131) & (g3153) & (g3161) & (!g3184) & (!g3187)));
	assign g4270 = (((!g2296) & (!g2344) & (!g2968) & (!g4232) & (!g4233) & (g3020)) + ((!g2296) & (!g2344) & (!g2968) & (!g4232) & (g4233) & (g3020)) + ((!g2296) & (!g2344) & (!g2968) & (g4232) & (!g4233) & (g3020)) + ((!g2296) & (!g2344) & (!g2968) & (g4232) & (g4233) & (g3020)) + ((!g2296) & (!g2344) & (g2968) & (!g4232) & (!g4233) & (g3020)) + ((!g2296) & (!g2344) & (g2968) & (!g4232) & (g4233) & (!g3020)) + ((!g2296) & (!g2344) & (g2968) & (g4232) & (!g4233) & (!g3020)) + ((!g2296) & (!g2344) & (g2968) & (g4232) & (g4233) & (!g3020)) + ((!g2296) & (g2344) & (!g2968) & (!g4232) & (!g4233) & (!g3020)) + ((!g2296) & (g2344) & (!g2968) & (!g4232) & (g4233) & (!g3020)) + ((!g2296) & (g2344) & (!g2968) & (g4232) & (!g4233) & (!g3020)) + ((!g2296) & (g2344) & (!g2968) & (g4232) & (g4233) & (!g3020)) + ((!g2296) & (g2344) & (g2968) & (!g4232) & (!g4233) & (!g3020)) + ((!g2296) & (g2344) & (g2968) & (!g4232) & (g4233) & (g3020)) + ((!g2296) & (g2344) & (g2968) & (g4232) & (!g4233) & (g3020)) + ((!g2296) & (g2344) & (g2968) & (g4232) & (g4233) & (g3020)) + ((g2296) & (!g2344) & (!g2968) & (!g4232) & (!g4233) & (g3020)) + ((g2296) & (!g2344) & (!g2968) & (!g4232) & (g4233) & (!g3020)) + ((g2296) & (!g2344) & (!g2968) & (g4232) & (!g4233) & (!g3020)) + ((g2296) & (!g2344) & (!g2968) & (g4232) & (g4233) & (!g3020)) + ((g2296) & (!g2344) & (g2968) & (!g4232) & (!g4233) & (!g3020)) + ((g2296) & (!g2344) & (g2968) & (!g4232) & (g4233) & (!g3020)) + ((g2296) & (!g2344) & (g2968) & (g4232) & (!g4233) & (!g3020)) + ((g2296) & (!g2344) & (g2968) & (g4232) & (g4233) & (!g3020)) + ((g2296) & (g2344) & (!g2968) & (!g4232) & (!g4233) & (!g3020)) + ((g2296) & (g2344) & (!g2968) & (!g4232) & (g4233) & (g3020)) + ((g2296) & (g2344) & (!g2968) & (g4232) & (!g4233) & (g3020)) + ((g2296) & (g2344) & (!g2968) & (g4232) & (g4233) & (g3020)) + ((g2296) & (g2344) & (g2968) & (!g4232) & (!g4233) & (g3020)) + ((g2296) & (g2344) & (g2968) & (!g4232) & (g4233) & (g3020)) + ((g2296) & (g2344) & (g2968) & (g4232) & (!g4233) & (g3020)) + ((g2296) & (g2344) & (g2968) & (g4232) & (g4233) & (g3020)));
	assign g4271 = (((!g1914) & (!g4269) & (!g3235) & (!g3255) & (g4270)) + ((!g1914) & (!g4269) & (!g3235) & (g3255) & (g4270)) + ((!g1914) & (!g4269) & (g3235) & (!g3255) & (g4270)) + ((!g1914) & (!g4269) & (g3235) & (g3255) & (g4270)) + ((!g1914) & (g4269) & (!g3235) & (!g3255) & (g4270)) + ((!g1914) & (g4269) & (!g3235) & (g3255) & (g4270)) + ((!g1914) & (g4269) & (g3235) & (!g3255) & (g4270)) + ((!g1914) & (g4269) & (g3235) & (g3255) & (g4270)) + ((g1914) & (!g4269) & (!g3235) & (!g3255) & (!g4270)) + ((g1914) & (!g4269) & (!g3235) & (!g3255) & (g4270)) + ((g1914) & (!g4269) & (g3235) & (g3255) & (!g4270)) + ((g1914) & (!g4269) & (g3235) & (g3255) & (g4270)) + ((g1914) & (g4269) & (!g3235) & (g3255) & (!g4270)) + ((g1914) & (g4269) & (!g3235) & (g3255) & (g4270)) + ((g1914) & (g4269) & (g3235) & (!g3255) & (!g4270)) + ((g1914) & (g4269) & (g3235) & (!g3255) & (g4270)));
	assign g4272 = (((!g830) & (!g2112) & (!g4271) & (key[131])) + ((!g830) & (!g2112) & (g4271) & (key[131])) + ((!g830) & (g2112) & (!g4271) & (key[131])) + ((!g830) & (g2112) & (g4271) & (key[131])) + ((g830) & (!g2112) & (g4271) & (!key[131])) + ((g830) & (!g2112) & (g4271) & (key[131])) + ((g830) & (g2112) & (!g4271) & (!key[131])) + ((g830) & (g2112) & (!g4271) & (key[131])));
	assign g4273 = (((!g2956) & (!g3005) & (!g4183) & (!g4184) & (!g2968) & (g3020)) + ((!g2956) & (!g3005) & (!g4183) & (!g4184) & (g2968) & (g3020)) + ((!g2956) & (!g3005) & (!g4183) & (g4184) & (!g2968) & (g3020)) + ((!g2956) & (!g3005) & (!g4183) & (g4184) & (g2968) & (!g3020)) + ((!g2956) & (!g3005) & (g4183) & (!g4184) & (!g2968) & (g3020)) + ((!g2956) & (!g3005) & (g4183) & (!g4184) & (g2968) & (!g3020)) + ((!g2956) & (!g3005) & (g4183) & (g4184) & (!g2968) & (g3020)) + ((!g2956) & (!g3005) & (g4183) & (g4184) & (g2968) & (!g3020)) + ((!g2956) & (g3005) & (!g4183) & (!g4184) & (!g2968) & (!g3020)) + ((!g2956) & (g3005) & (!g4183) & (!g4184) & (g2968) & (!g3020)) + ((!g2956) & (g3005) & (!g4183) & (g4184) & (!g2968) & (!g3020)) + ((!g2956) & (g3005) & (!g4183) & (g4184) & (g2968) & (g3020)) + ((!g2956) & (g3005) & (g4183) & (!g4184) & (!g2968) & (!g3020)) + ((!g2956) & (g3005) & (g4183) & (!g4184) & (g2968) & (g3020)) + ((!g2956) & (g3005) & (g4183) & (g4184) & (!g2968) & (!g3020)) + ((!g2956) & (g3005) & (g4183) & (g4184) & (g2968) & (g3020)) + ((g2956) & (!g3005) & (!g4183) & (!g4184) & (!g2968) & (g3020)) + ((g2956) & (!g3005) & (!g4183) & (!g4184) & (g2968) & (!g3020)) + ((g2956) & (!g3005) & (!g4183) & (g4184) & (!g2968) & (!g3020)) + ((g2956) & (!g3005) & (!g4183) & (g4184) & (g2968) & (!g3020)) + ((g2956) & (!g3005) & (g4183) & (!g4184) & (!g2968) & (!g3020)) + ((g2956) & (!g3005) & (g4183) & (!g4184) & (g2968) & (!g3020)) + ((g2956) & (!g3005) & (g4183) & (g4184) & (!g2968) & (!g3020)) + ((g2956) & (!g3005) & (g4183) & (g4184) & (g2968) & (!g3020)) + ((g2956) & (g3005) & (!g4183) & (!g4184) & (!g2968) & (!g3020)) + ((g2956) & (g3005) & (!g4183) & (!g4184) & (g2968) & (g3020)) + ((g2956) & (g3005) & (!g4183) & (g4184) & (!g2968) & (g3020)) + ((g2956) & (g3005) & (!g4183) & (g4184) & (g2968) & (g3020)) + ((g2956) & (g3005) & (g4183) & (!g4184) & (!g2968) & (g3020)) + ((g2956) & (g3005) & (g4183) & (!g4184) & (g2968) & (g3020)) + ((g2956) & (g3005) & (g4183) & (g4184) & (!g2968) & (g3020)) + ((g2956) & (g3005) & (g4183) & (g4184) & (g2968) & (g3020)));
	assign g4274 = (((!g2556) & (!g2602) & (!g1711) & (!g1744) & (!g4137) & (!g4138)) + ((!g2556) & (!g2602) & (!g1711) & (!g1744) & (!g4137) & (g4138)) + ((!g2556) & (!g2602) & (!g1711) & (!g1744) & (g4137) & (!g4138)) + ((!g2556) & (!g2602) & (!g1711) & (!g1744) & (g4137) & (g4138)) + ((!g2556) & (!g2602) & (!g1711) & (g1744) & (!g4137) & (!g4138)) + ((!g2556) & (!g2602) & (!g1711) & (g1744) & (!g4137) & (g4138)) + ((!g2556) & (!g2602) & (!g1711) & (g1744) & (g4137) & (!g4138)) + ((!g2556) & (!g2602) & (!g1711) & (g1744) & (g4137) & (g4138)) + ((!g2556) & (!g2602) & (g1711) & (!g1744) & (!g4137) & (!g4138)) + ((!g2556) & (!g2602) & (g1711) & (!g1744) & (!g4137) & (g4138)) + ((!g2556) & (!g2602) & (g1711) & (!g1744) & (g4137) & (!g4138)) + ((!g2556) & (!g2602) & (g1711) & (!g1744) & (g4137) & (g4138)) + ((!g2556) & (!g2602) & (g1711) & (g1744) & (!g4137) & (!g4138)) + ((!g2556) & (g2602) & (!g1711) & (!g1744) & (!g4137) & (!g4138)) + ((!g2556) & (g2602) & (!g1711) & (!g1744) & (!g4137) & (g4138)) + ((!g2556) & (g2602) & (!g1711) & (!g1744) & (g4137) & (!g4138)) + ((!g2556) & (g2602) & (!g1711) & (!g1744) & (g4137) & (g4138)) + ((!g2556) & (g2602) & (g1711) & (!g1744) & (!g4137) & (!g4138)) + ((g2556) & (!g2602) & (!g1711) & (!g1744) & (!g4137) & (!g4138)) + ((g2556) & (!g2602) & (!g1711) & (!g1744) & (!g4137) & (g4138)) + ((g2556) & (!g2602) & (!g1711) & (!g1744) & (g4137) & (!g4138)) + ((g2556) & (!g2602) & (!g1711) & (!g1744) & (g4137) & (g4138)) + ((g2556) & (!g2602) & (!g1711) & (g1744) & (!g4137) & (!g4138)) + ((g2556) & (!g2602) & (g1711) & (!g1744) & (!g4137) & (!g4138)) + ((g2556) & (!g2602) & (g1711) & (!g1744) & (!g4137) & (g4138)) + ((g2556) & (!g2602) & (g1711) & (!g1744) & (g4137) & (!g4138)) + ((g2556) & (!g2602) & (g1711) & (!g1744) & (g4137) & (g4138)) + ((g2556) & (g2602) & (!g1711) & (!g1744) & (!g4137) & (!g4138)));
	assign g4275 = (((!g1914) & (!g2650) & (!g1778) & (!g4273) & (!g4274)) + ((!g1914) & (!g2650) & (!g1778) & (g4273) & (!g4274)) + ((!g1914) & (!g2650) & (g1778) & (!g4273) & (g4274)) + ((!g1914) & (!g2650) & (g1778) & (g4273) & (g4274)) + ((!g1914) & (g2650) & (!g1778) & (!g4273) & (g4274)) + ((!g1914) & (g2650) & (!g1778) & (g4273) & (g4274)) + ((!g1914) & (g2650) & (g1778) & (!g4273) & (!g4274)) + ((!g1914) & (g2650) & (g1778) & (g4273) & (!g4274)) + ((g1914) & (!g2650) & (!g1778) & (g4273) & (!g4274)) + ((g1914) & (!g2650) & (!g1778) & (g4273) & (g4274)) + ((g1914) & (!g2650) & (g1778) & (g4273) & (!g4274)) + ((g1914) & (!g2650) & (g1778) & (g4273) & (g4274)) + ((g1914) & (g2650) & (!g1778) & (g4273) & (!g4274)) + ((g1914) & (g2650) & (!g1778) & (g4273) & (g4274)) + ((g1914) & (g2650) & (g1778) & (g4273) & (!g4274)) + ((g1914) & (g2650) & (g1778) & (g4273) & (g4274)));
	assign g4276 = (((!g830) & (!g2114) & (!g4275) & (key[99])) + ((!g830) & (!g2114) & (g4275) & (key[99])) + ((!g830) & (g2114) & (!g4275) & (key[99])) + ((!g830) & (g2114) & (g4275) & (key[99])) + ((g830) & (!g2114) & (g4275) & (!key[99])) + ((g830) & (!g2114) & (g4275) & (key[99])) + ((g830) & (g2114) & (!g4275) & (!key[99])) + ((g830) & (g2114) & (!g4275) & (key[99])));
	assign g4277 = (((!g3163) & (!g4142) & (!g4143) & (!g3149) & (!g3193) & (!g3199)) + ((!g3163) & (!g4142) & (!g4143) & (!g3149) & (!g3193) & (g3199)) + ((!g3163) & (!g4142) & (!g4143) & (!g3149) & (g3193) & (!g3199)) + ((!g3163) & (!g4142) & (!g4143) & (g3149) & (!g3193) & (!g3199)) + ((!g3163) & (!g4142) & (!g4143) & (g3149) & (!g3193) & (g3199)) + ((!g3163) & (!g4142) & (!g4143) & (g3149) & (g3193) & (!g3199)) + ((!g3163) & (!g4142) & (g4143) & (!g3149) & (!g3193) & (!g3199)) + ((!g3163) & (!g4142) & (g4143) & (!g3149) & (!g3193) & (g3199)) + ((!g3163) & (!g4142) & (g4143) & (!g3149) & (g3193) & (!g3199)) + ((!g3163) & (!g4142) & (g4143) & (g3149) & (!g3193) & (!g3199)) + ((!g3163) & (g4142) & (!g4143) & (!g3149) & (!g3193) & (!g3199)) + ((!g3163) & (g4142) & (!g4143) & (!g3149) & (!g3193) & (g3199)) + ((!g3163) & (g4142) & (!g4143) & (!g3149) & (g3193) & (!g3199)) + ((!g3163) & (g4142) & (!g4143) & (g3149) & (!g3193) & (!g3199)) + ((!g3163) & (g4142) & (g4143) & (!g3149) & (!g3193) & (!g3199)) + ((!g3163) & (g4142) & (g4143) & (!g3149) & (!g3193) & (g3199)) + ((!g3163) & (g4142) & (g4143) & (!g3149) & (g3193) & (!g3199)) + ((!g3163) & (g4142) & (g4143) & (g3149) & (!g3193) & (!g3199)) + ((g3163) & (!g4142) & (!g4143) & (!g3149) & (!g3193) & (!g3199)) + ((g3163) & (!g4142) & (!g4143) & (!g3149) & (!g3193) & (g3199)) + ((g3163) & (!g4142) & (!g4143) & (!g3149) & (g3193) & (!g3199)) + ((g3163) & (!g4142) & (!g4143) & (g3149) & (!g3193) & (!g3199)) + ((g3163) & (!g4142) & (g4143) & (!g3149) & (!g3193) & (!g3199)) + ((g3163) & (!g4142) & (g4143) & (g3149) & (!g3193) & (!g3199)) + ((g3163) & (g4142) & (!g4143) & (!g3149) & (!g3193) & (!g3199)) + ((g3163) & (g4142) & (!g4143) & (g3149) & (!g3193) & (!g3199)) + ((g3163) & (g4142) & (g4143) & (!g3149) & (!g3193) & (!g3199)) + ((g3163) & (g4142) & (g4143) & (g3149) & (!g3193) & (!g3199)));
	assign g4278 = (((!g2295) & (!g2343) & (!g2979) & (g3007) & (!g4196) & (!g4197)) + ((!g2295) & (!g2343) & (!g2979) & (g3007) & (!g4196) & (g4197)) + ((!g2295) & (!g2343) & (!g2979) & (g3007) & (g4196) & (!g4197)) + ((!g2295) & (!g2343) & (!g2979) & (g3007) & (g4196) & (g4197)) + ((!g2295) & (!g2343) & (g2979) & (!g3007) & (!g4196) & (g4197)) + ((!g2295) & (!g2343) & (g2979) & (!g3007) & (g4196) & (!g4197)) + ((!g2295) & (!g2343) & (g2979) & (!g3007) & (g4196) & (g4197)) + ((!g2295) & (!g2343) & (g2979) & (g3007) & (!g4196) & (!g4197)) + ((!g2295) & (g2343) & (!g2979) & (!g3007) & (!g4196) & (!g4197)) + ((!g2295) & (g2343) & (!g2979) & (!g3007) & (!g4196) & (g4197)) + ((!g2295) & (g2343) & (!g2979) & (!g3007) & (g4196) & (!g4197)) + ((!g2295) & (g2343) & (!g2979) & (!g3007) & (g4196) & (g4197)) + ((!g2295) & (g2343) & (g2979) & (!g3007) & (!g4196) & (!g4197)) + ((!g2295) & (g2343) & (g2979) & (g3007) & (!g4196) & (g4197)) + ((!g2295) & (g2343) & (g2979) & (g3007) & (g4196) & (!g4197)) + ((!g2295) & (g2343) & (g2979) & (g3007) & (g4196) & (g4197)) + ((g2295) & (!g2343) & (!g2979) & (!g3007) & (!g4196) & (g4197)) + ((g2295) & (!g2343) & (!g2979) & (!g3007) & (g4196) & (!g4197)) + ((g2295) & (!g2343) & (!g2979) & (!g3007) & (g4196) & (g4197)) + ((g2295) & (!g2343) & (!g2979) & (g3007) & (!g4196) & (!g4197)) + ((g2295) & (!g2343) & (g2979) & (!g3007) & (!g4196) & (!g4197)) + ((g2295) & (!g2343) & (g2979) & (!g3007) & (!g4196) & (g4197)) + ((g2295) & (!g2343) & (g2979) & (!g3007) & (g4196) & (!g4197)) + ((g2295) & (!g2343) & (g2979) & (!g3007) & (g4196) & (g4197)) + ((g2295) & (g2343) & (!g2979) & (!g3007) & (!g4196) & (!g4197)) + ((g2295) & (g2343) & (!g2979) & (g3007) & (!g4196) & (g4197)) + ((g2295) & (g2343) & (!g2979) & (g3007) & (g4196) & (!g4197)) + ((g2295) & (g2343) & (!g2979) & (g3007) & (g4196) & (g4197)) + ((g2295) & (g2343) & (g2979) & (g3007) & (!g4196) & (!g4197)) + ((g2295) & (g2343) & (g2979) & (g3007) & (!g4196) & (g4197)) + ((g2295) & (g2343) & (g2979) & (g3007) & (g4196) & (!g4197)) + ((g2295) & (g2343) & (g2979) & (g3007) & (g4196) & (g4197)));
	assign g4279 = (((!g1914) & (!g3260) & (!g4277) & (!g3222) & (g4278)) + ((!g1914) & (!g3260) & (!g4277) & (g3222) & (g4278)) + ((!g1914) & (!g3260) & (g4277) & (!g3222) & (g4278)) + ((!g1914) & (!g3260) & (g4277) & (g3222) & (g4278)) + ((!g1914) & (g3260) & (!g4277) & (!g3222) & (g4278)) + ((!g1914) & (g3260) & (!g4277) & (g3222) & (g4278)) + ((!g1914) & (g3260) & (g4277) & (!g3222) & (g4278)) + ((!g1914) & (g3260) & (g4277) & (g3222) & (g4278)) + ((g1914) & (!g3260) & (!g4277) & (!g3222) & (!g4278)) + ((g1914) & (!g3260) & (!g4277) & (!g3222) & (g4278)) + ((g1914) & (!g3260) & (g4277) & (g3222) & (!g4278)) + ((g1914) & (!g3260) & (g4277) & (g3222) & (g4278)) + ((g1914) & (g3260) & (!g4277) & (g3222) & (!g4278)) + ((g1914) & (g3260) & (!g4277) & (g3222) & (g4278)) + ((g1914) & (g3260) & (g4277) & (!g3222) & (!g4278)) + ((g1914) & (g3260) & (g4277) & (!g3222) & (g4278)));
	assign g4280 = (((!g830) & (!g2116) & (!g4279) & (nonce[3])) + ((!g830) & (!g2116) & (g4279) & (nonce[3])) + ((!g830) & (g2116) & (!g4279) & (nonce[3])) + ((!g830) & (g2116) & (g4279) & (nonce[3])) + ((g830) & (!g2116) & (g4279) & (!nonce[3])) + ((g830) & (!g2116) & (g4279) & (nonce[3])) + ((g830) & (g2116) & (!g4279) & (!nonce[3])) + ((g830) & (g2116) & (!g4279) & (nonce[3])));
	assign g4281 = (((!g2690) & (!g2774) & (!g2747) & (g2780) & (!g4225)) + ((!g2690) & (!g2774) & (!g2747) & (g2780) & (g4225)) + ((!g2690) & (!g2774) & (g2747) & (!g2780) & (g4225)) + ((!g2690) & (!g2774) & (g2747) & (g2780) & (!g4225)) + ((!g2690) & (g2774) & (!g2747) & (!g2780) & (!g4225)) + ((!g2690) & (g2774) & (!g2747) & (!g2780) & (g4225)) + ((!g2690) & (g2774) & (g2747) & (!g2780) & (!g4225)) + ((!g2690) & (g2774) & (g2747) & (g2780) & (g4225)) + ((g2690) & (!g2774) & (!g2747) & (!g2780) & (g4225)) + ((g2690) & (!g2774) & (!g2747) & (g2780) & (!g4225)) + ((g2690) & (!g2774) & (g2747) & (!g2780) & (!g4225)) + ((g2690) & (!g2774) & (g2747) & (!g2780) & (g4225)) + ((g2690) & (g2774) & (!g2747) & (!g2780) & (!g4225)) + ((g2690) & (g2774) & (!g2747) & (g2780) & (g4225)) + ((g2690) & (g2774) & (g2747) & (g2780) & (!g4225)) + ((g2690) & (g2774) & (g2747) & (g2780) & (g4225)));
	assign g4282 = (((!g2653) & (!g2718) & (g2674) & (g2733) & (g4148)) + ((!g2653) & (g2718) & (!g2674) & (g2733) & (!g4148)) + ((!g2653) & (g2718) & (!g2674) & (g2733) & (g4148)) + ((!g2653) & (g2718) & (g2674) & (!g2733) & (g4148)) + ((!g2653) & (g2718) & (g2674) & (g2733) & (!g4148)) + ((!g2653) & (g2718) & (g2674) & (g2733) & (g4148)) + ((g2653) & (!g2718) & (!g2674) & (g2733) & (g4148)) + ((g2653) & (!g2718) & (g2674) & (g2733) & (!g4148)) + ((g2653) & (!g2718) & (g2674) & (g2733) & (g4148)) + ((g2653) & (g2718) & (!g2674) & (!g2733) & (g4148)) + ((g2653) & (g2718) & (!g2674) & (g2733) & (!g4148)) + ((g2653) & (g2718) & (!g2674) & (g2733) & (g4148)) + ((g2653) & (g2718) & (g2674) & (!g2733) & (!g4148)) + ((g2653) & (g2718) & (g2674) & (!g2733) & (g4148)) + ((g2653) & (g2718) & (g2674) & (g2733) & (!g4148)) + ((g2653) & (g2718) & (g2674) & (g2733) & (g4148)));
	assign g4283 = (((!g3128) & (g3125)) + ((g3128) & (!g3125)));
	assign g4284 = (((!g3053) & (!g3088) & (g3050) & (g3080) & (!g3826) & (g4283)) + ((!g3053) & (g3088) & (!g3050) & (g3080) & (!g3826) & (g4283)) + ((!g3053) & (g3088) & (!g3050) & (g3080) & (g3826) & (g4283)) + ((!g3053) & (g3088) & (g3050) & (!g3080) & (!g3826) & (g4283)) + ((!g3053) & (g3088) & (g3050) & (g3080) & (!g3826) & (g4283)) + ((!g3053) & (g3088) & (g3050) & (g3080) & (g3826) & (g4283)) + ((g3053) & (!g3088) & (!g3050) & (g3080) & (!g3826) & (g4283)) + ((g3053) & (!g3088) & (g3050) & (g3080) & (!g3826) & (g4283)) + ((g3053) & (!g3088) & (g3050) & (g3080) & (g3826) & (g4283)) + ((g3053) & (g3088) & (!g3050) & (!g3080) & (!g3826) & (g4283)) + ((g3053) & (g3088) & (!g3050) & (g3080) & (!g3826) & (g4283)) + ((g3053) & (g3088) & (!g3050) & (g3080) & (g3826) & (g4283)) + ((g3053) & (g3088) & (g3050) & (!g3080) & (!g3826) & (g4283)) + ((g3053) & (g3088) & (g3050) & (!g3080) & (g3826) & (g4283)) + ((g3053) & (g3088) & (g3050) & (g3080) & (!g3826) & (g4283)) + ((g3053) & (g3088) & (g3050) & (g3080) & (g3826) & (g4283)));
	assign g4285 = (((g3128) & (g3125)));
	assign g4286 = (((!g3163) & (!g3155) & (!g4284) & (g4285)) + ((!g3163) & (!g3155) & (g4284) & (!g4285)) + ((!g3163) & (!g3155) & (g4284) & (g4285)) + ((!g3163) & (g3155) & (!g4284) & (!g4285)) + ((g3163) & (!g3155) & (!g4284) & (!g4285)) + ((g3163) & (g3155) & (!g4284) & (g4285)) + ((g3163) & (g3155) & (g4284) & (!g4285)) + ((g3163) & (g3155) & (g4284) & (g4285)));
	assign g4287 = (((!g2516) & (g3142)) + ((g2516) & (!g3142)));
	assign g4288 = (((!g2377) & (!g2424) & (g3067) & (g3097) & (!g3843) & (g4287)) + ((!g2377) & (g2424) & (!g3067) & (g3097) & (!g3843) & (g4287)) + ((!g2377) & (g2424) & (!g3067) & (g3097) & (g3843) & (g4287)) + ((!g2377) & (g2424) & (g3067) & (!g3097) & (!g3843) & (g4287)) + ((!g2377) & (g2424) & (g3067) & (g3097) & (!g3843) & (g4287)) + ((!g2377) & (g2424) & (g3067) & (g3097) & (g3843) & (g4287)) + ((g2377) & (!g2424) & (!g3067) & (g3097) & (!g3843) & (g4287)) + ((g2377) & (!g2424) & (g3067) & (g3097) & (!g3843) & (g4287)) + ((g2377) & (!g2424) & (g3067) & (g3097) & (g3843) & (g4287)) + ((g2377) & (g2424) & (!g3067) & (!g3097) & (!g3843) & (g4287)) + ((g2377) & (g2424) & (!g3067) & (g3097) & (!g3843) & (g4287)) + ((g2377) & (g2424) & (!g3067) & (g3097) & (g3843) & (g4287)) + ((g2377) & (g2424) & (g3067) & (!g3097) & (!g3843) & (g4287)) + ((g2377) & (g2424) & (g3067) & (!g3097) & (g3843) & (g4287)) + ((g2377) & (g2424) & (g3067) & (g3097) & (!g3843) & (g4287)) + ((g2377) & (g2424) & (g3067) & (g3097) & (g3843) & (g4287)));
	assign g4289 = (((g2516) & (g3142)));
	assign g4290 = (((!g2552) & (!g3172) & (!g4288) & (g4289)) + ((!g2552) & (!g3172) & (g4288) & (!g4289)) + ((!g2552) & (!g3172) & (g4288) & (g4289)) + ((!g2552) & (g3172) & (!g4288) & (!g4289)) + ((g2552) & (!g3172) & (!g4288) & (!g4289)) + ((g2552) & (g3172) & (!g4288) & (g4289)) + ((g2552) & (g3172) & (g4288) & (!g4289)) + ((g2552) & (g3172) & (g4288) & (g4289)));
	assign g4291 = (((!g830) & (!g1914) & (!g2120) & (!g4286) & (!g4290) & (nonce[35])) + ((!g830) & (!g1914) & (!g2120) & (!g4286) & (g4290) & (nonce[35])) + ((!g830) & (!g1914) & (!g2120) & (g4286) & (!g4290) & (nonce[35])) + ((!g830) & (!g1914) & (!g2120) & (g4286) & (g4290) & (nonce[35])) + ((!g830) & (!g1914) & (g2120) & (!g4286) & (!g4290) & (nonce[35])) + ((!g830) & (!g1914) & (g2120) & (!g4286) & (g4290) & (nonce[35])) + ((!g830) & (!g1914) & (g2120) & (g4286) & (!g4290) & (nonce[35])) + ((!g830) & (!g1914) & (g2120) & (g4286) & (g4290) & (nonce[35])) + ((!g830) & (g1914) & (!g2120) & (!g4286) & (!g4290) & (nonce[35])) + ((!g830) & (g1914) & (!g2120) & (!g4286) & (g4290) & (nonce[35])) + ((!g830) & (g1914) & (!g2120) & (g4286) & (!g4290) & (nonce[35])) + ((!g830) & (g1914) & (!g2120) & (g4286) & (g4290) & (nonce[35])) + ((!g830) & (g1914) & (g2120) & (!g4286) & (!g4290) & (nonce[35])) + ((!g830) & (g1914) & (g2120) & (!g4286) & (g4290) & (nonce[35])) + ((!g830) & (g1914) & (g2120) & (g4286) & (!g4290) & (nonce[35])) + ((!g830) & (g1914) & (g2120) & (g4286) & (g4290) & (nonce[35])) + ((g830) & (!g1914) & (!g2120) & (!g4286) & (g4290) & (!nonce[35])) + ((g830) & (!g1914) & (!g2120) & (!g4286) & (g4290) & (nonce[35])) + ((g830) & (!g1914) & (!g2120) & (g4286) & (g4290) & (!nonce[35])) + ((g830) & (!g1914) & (!g2120) & (g4286) & (g4290) & (nonce[35])) + ((g830) & (!g1914) & (g2120) & (!g4286) & (!g4290) & (!nonce[35])) + ((g830) & (!g1914) & (g2120) & (!g4286) & (!g4290) & (nonce[35])) + ((g830) & (!g1914) & (g2120) & (g4286) & (!g4290) & (!nonce[35])) + ((g830) & (!g1914) & (g2120) & (g4286) & (!g4290) & (nonce[35])) + ((g830) & (g1914) & (!g2120) & (g4286) & (!g4290) & (!nonce[35])) + ((g830) & (g1914) & (!g2120) & (g4286) & (!g4290) & (nonce[35])) + ((g830) & (g1914) & (!g2120) & (g4286) & (g4290) & (!nonce[35])) + ((g830) & (g1914) & (!g2120) & (g4286) & (g4290) & (nonce[35])) + ((g830) & (g1914) & (g2120) & (!g4286) & (!g4290) & (!nonce[35])) + ((g830) & (g1914) & (g2120) & (!g4286) & (!g4290) & (nonce[35])) + ((g830) & (g1914) & (g2120) & (!g4286) & (g4290) & (!nonce[35])) + ((g830) & (g1914) & (g2120) & (!g4286) & (g4290) & (nonce[35])));
	assign g4292 = (((!g2299) & (!g2348) & (!g4202) & (!g4203) & (!g2985) & (g3015)) + ((!g2299) & (!g2348) & (!g4202) & (!g4203) & (g2985) & (g3015)) + ((!g2299) & (!g2348) & (!g4202) & (g4203) & (!g2985) & (g3015)) + ((!g2299) & (!g2348) & (!g4202) & (g4203) & (g2985) & (!g3015)) + ((!g2299) & (!g2348) & (g4202) & (!g4203) & (!g2985) & (g3015)) + ((!g2299) & (!g2348) & (g4202) & (!g4203) & (g2985) & (!g3015)) + ((!g2299) & (!g2348) & (g4202) & (g4203) & (!g2985) & (g3015)) + ((!g2299) & (!g2348) & (g4202) & (g4203) & (g2985) & (!g3015)) + ((!g2299) & (g2348) & (!g4202) & (!g4203) & (!g2985) & (!g3015)) + ((!g2299) & (g2348) & (!g4202) & (!g4203) & (g2985) & (!g3015)) + ((!g2299) & (g2348) & (!g4202) & (g4203) & (!g2985) & (!g3015)) + ((!g2299) & (g2348) & (!g4202) & (g4203) & (g2985) & (g3015)) + ((!g2299) & (g2348) & (g4202) & (!g4203) & (!g2985) & (!g3015)) + ((!g2299) & (g2348) & (g4202) & (!g4203) & (g2985) & (g3015)) + ((!g2299) & (g2348) & (g4202) & (g4203) & (!g2985) & (!g3015)) + ((!g2299) & (g2348) & (g4202) & (g4203) & (g2985) & (g3015)) + ((g2299) & (!g2348) & (!g4202) & (!g4203) & (!g2985) & (g3015)) + ((g2299) & (!g2348) & (!g4202) & (!g4203) & (g2985) & (!g3015)) + ((g2299) & (!g2348) & (!g4202) & (g4203) & (!g2985) & (!g3015)) + ((g2299) & (!g2348) & (!g4202) & (g4203) & (g2985) & (!g3015)) + ((g2299) & (!g2348) & (g4202) & (!g4203) & (!g2985) & (!g3015)) + ((g2299) & (!g2348) & (g4202) & (!g4203) & (g2985) & (!g3015)) + ((g2299) & (!g2348) & (g4202) & (g4203) & (!g2985) & (!g3015)) + ((g2299) & (!g2348) & (g4202) & (g4203) & (g2985) & (!g3015)) + ((g2299) & (g2348) & (!g4202) & (!g4203) & (!g2985) & (!g3015)) + ((g2299) & (g2348) & (!g4202) & (!g4203) & (g2985) & (g3015)) + ((g2299) & (g2348) & (!g4202) & (g4203) & (!g2985) & (g3015)) + ((g2299) & (g2348) & (!g4202) & (g4203) & (g2985) & (g3015)) + ((g2299) & (g2348) & (g4202) & (!g4203) & (!g2985) & (g3015)) + ((g2299) & (g2348) & (g4202) & (!g4203) & (g2985) & (g3015)) + ((g2299) & (g2348) & (g4202) & (g4203) & (!g2985) & (g3015)) + ((g2299) & (g2348) & (g4202) & (g4203) & (g2985) & (g3015)));
	assign g4293 = (((!g3153) & (!g4156) & (!g4157) & (!g3155) & (!g3184) & (!g3196)) + ((!g3153) & (!g4156) & (!g4157) & (!g3155) & (!g3184) & (g3196)) + ((!g3153) & (!g4156) & (!g4157) & (!g3155) & (g3184) & (!g3196)) + ((!g3153) & (!g4156) & (!g4157) & (g3155) & (!g3184) & (!g3196)) + ((!g3153) & (!g4156) & (!g4157) & (g3155) & (!g3184) & (g3196)) + ((!g3153) & (!g4156) & (!g4157) & (g3155) & (g3184) & (!g3196)) + ((!g3153) & (!g4156) & (g4157) & (!g3155) & (!g3184) & (!g3196)) + ((!g3153) & (!g4156) & (g4157) & (!g3155) & (!g3184) & (g3196)) + ((!g3153) & (!g4156) & (g4157) & (!g3155) & (g3184) & (!g3196)) + ((!g3153) & (!g4156) & (g4157) & (g3155) & (!g3184) & (!g3196)) + ((!g3153) & (g4156) & (!g4157) & (!g3155) & (!g3184) & (!g3196)) + ((!g3153) & (g4156) & (!g4157) & (!g3155) & (!g3184) & (g3196)) + ((!g3153) & (g4156) & (!g4157) & (!g3155) & (g3184) & (!g3196)) + ((!g3153) & (g4156) & (!g4157) & (g3155) & (!g3184) & (!g3196)) + ((!g3153) & (g4156) & (g4157) & (!g3155) & (!g3184) & (!g3196)) + ((!g3153) & (g4156) & (g4157) & (!g3155) & (!g3184) & (g3196)) + ((!g3153) & (g4156) & (g4157) & (!g3155) & (g3184) & (!g3196)) + ((!g3153) & (g4156) & (g4157) & (g3155) & (!g3184) & (!g3196)) + ((g3153) & (!g4156) & (!g4157) & (!g3155) & (!g3184) & (!g3196)) + ((g3153) & (!g4156) & (!g4157) & (!g3155) & (!g3184) & (g3196)) + ((g3153) & (!g4156) & (!g4157) & (!g3155) & (g3184) & (!g3196)) + ((g3153) & (!g4156) & (!g4157) & (g3155) & (!g3184) & (!g3196)) + ((g3153) & (!g4156) & (g4157) & (!g3155) & (!g3184) & (!g3196)) + ((g3153) & (!g4156) & (g4157) & (g3155) & (!g3184) & (!g3196)) + ((g3153) & (g4156) & (!g4157) & (!g3155) & (!g3184) & (!g3196)) + ((g3153) & (g4156) & (!g4157) & (g3155) & (!g3184) & (!g3196)) + ((g3153) & (g4156) & (g4157) & (!g3155) & (!g3184) & (!g3196)) + ((g3153) & (g4156) & (g4157) & (g3155) & (!g3184) & (!g3196)));
	assign g4294 = (((!g1914) & (!g3235) & (!g4292) & (!g4293) & (!g3240)) + ((!g1914) & (!g3235) & (!g4292) & (g4293) & (g3240)) + ((!g1914) & (!g3235) & (g4292) & (!g4293) & (!g3240)) + ((!g1914) & (!g3235) & (g4292) & (g4293) & (g3240)) + ((!g1914) & (g3235) & (!g4292) & (!g4293) & (g3240)) + ((!g1914) & (g3235) & (!g4292) & (g4293) & (!g3240)) + ((!g1914) & (g3235) & (g4292) & (!g4293) & (g3240)) + ((!g1914) & (g3235) & (g4292) & (g4293) & (!g3240)) + ((g1914) & (!g3235) & (g4292) & (!g4293) & (!g3240)) + ((g1914) & (!g3235) & (g4292) & (!g4293) & (g3240)) + ((g1914) & (!g3235) & (g4292) & (g4293) & (!g3240)) + ((g1914) & (!g3235) & (g4292) & (g4293) & (g3240)) + ((g1914) & (g3235) & (g4292) & (!g4293) & (!g3240)) + ((g1914) & (g3235) & (g4292) & (!g4293) & (g3240)) + ((g1914) & (g3235) & (g4292) & (g4293) & (!g3240)) + ((g1914) & (g3235) & (g4292) & (g4293) & (g3240)));
	assign g4295 = (((!g830) & (!g2123) & (!g4294) & (key[227])) + ((!g830) & (!g2123) & (g4294) & (key[227])) + ((!g830) & (g2123) & (!g4294) & (key[227])) + ((!g830) & (g2123) & (g4294) & (key[227])) + ((g830) & (!g2123) & (g4294) & (!key[227])) + ((g830) & (!g2123) & (g4294) & (key[227])) + ((g830) & (g2123) & (!g4294) & (!key[227])) + ((g830) & (g2123) & (!g4294) & (key[227])));
	assign g4296 = (((!g2519) & (g3142)) + ((g2519) & (!g3142)));
	assign g4297 = (((!g2379) & (!g2427) & (g3067) & (g3097) & (!g3725) & (g4296)) + ((!g2379) & (g2427) & (!g3067) & (g3097) & (!g3725) & (g4296)) + ((!g2379) & (g2427) & (!g3067) & (g3097) & (g3725) & (g4296)) + ((!g2379) & (g2427) & (g3067) & (!g3097) & (!g3725) & (g4296)) + ((!g2379) & (g2427) & (g3067) & (g3097) & (!g3725) & (g4296)) + ((!g2379) & (g2427) & (g3067) & (g3097) & (g3725) & (g4296)) + ((g2379) & (!g2427) & (!g3067) & (g3097) & (!g3725) & (g4296)) + ((g2379) & (!g2427) & (g3067) & (g3097) & (!g3725) & (g4296)) + ((g2379) & (!g2427) & (g3067) & (g3097) & (g3725) & (g4296)) + ((g2379) & (g2427) & (!g3067) & (!g3097) & (!g3725) & (g4296)) + ((g2379) & (g2427) & (!g3067) & (g3097) & (!g3725) & (g4296)) + ((g2379) & (g2427) & (!g3067) & (g3097) & (g3725) & (g4296)) + ((g2379) & (g2427) & (g3067) & (!g3097) & (!g3725) & (g4296)) + ((g2379) & (g2427) & (g3067) & (!g3097) & (g3725) & (g4296)) + ((g2379) & (g2427) & (g3067) & (g3097) & (!g3725) & (g4296)) + ((g2379) & (g2427) & (g3067) & (g3097) & (g3725) & (g4296)));
	assign g4298 = (((g2519) & (g3142)));
	assign g4299 = (((!g2556) & (!g3172) & (!g4297) & (g4298)) + ((!g2556) & (!g3172) & (g4297) & (!g4298)) + ((!g2556) & (!g3172) & (g4297) & (g4298)) + ((!g2556) & (g3172) & (!g4297) & (!g4298)) + ((g2556) & (!g3172) & (!g4297) & (!g4298)) + ((g2556) & (g3172) & (!g4297) & (g4298)) + ((g2556) & (g3172) & (g4297) & (!g4298)) + ((g2556) & (g3172) & (g4297) & (g4298)));
	assign g4300 = (((!g3128) & (g3116)) + ((g3128) & (!g3116)));
	assign g4301 = (((!g3053) & (!g3088) & (!g3742) & (g3041) & (g3086) & (g4300)) + ((!g3053) & (g3088) & (!g3742) & (!g3041) & (g3086) & (g4300)) + ((!g3053) & (g3088) & (!g3742) & (g3041) & (!g3086) & (g4300)) + ((!g3053) & (g3088) & (!g3742) & (g3041) & (g3086) & (g4300)) + ((!g3053) & (g3088) & (g3742) & (!g3041) & (g3086) & (g4300)) + ((!g3053) & (g3088) & (g3742) & (g3041) & (g3086) & (g4300)) + ((g3053) & (!g3088) & (!g3742) & (!g3041) & (g3086) & (g4300)) + ((g3053) & (!g3088) & (!g3742) & (g3041) & (g3086) & (g4300)) + ((g3053) & (!g3088) & (g3742) & (g3041) & (g3086) & (g4300)) + ((g3053) & (g3088) & (!g3742) & (!g3041) & (!g3086) & (g4300)) + ((g3053) & (g3088) & (!g3742) & (!g3041) & (g3086) & (g4300)) + ((g3053) & (g3088) & (!g3742) & (g3041) & (!g3086) & (g4300)) + ((g3053) & (g3088) & (!g3742) & (g3041) & (g3086) & (g4300)) + ((g3053) & (g3088) & (g3742) & (!g3041) & (g3086) & (g4300)) + ((g3053) & (g3088) & (g3742) & (g3041) & (!g3086) & (g4300)) + ((g3053) & (g3088) & (g3742) & (g3041) & (g3086) & (g4300)));
	assign g4302 = (((g3128) & (g3116)));
	assign g4303 = (((!g3163) & (!g3161) & (!g4301) & (g4302)) + ((!g3163) & (!g3161) & (g4301) & (!g4302)) + ((!g3163) & (!g3161) & (g4301) & (g4302)) + ((!g3163) & (g3161) & (!g4301) & (!g4302)) + ((g3163) & (!g3161) & (!g4301) & (!g4302)) + ((g3163) & (g3161) & (!g4301) & (g4302)) + ((g3163) & (g3161) & (g4301) & (!g4302)) + ((g3163) & (g3161) & (g4301) & (g4302)));
	assign g4304 = (((!g830) & (!g1914) & (!g2125) & (!g4299) & (!g4303) & (key[195])) + ((!g830) & (!g1914) & (!g2125) & (!g4299) & (g4303) & (key[195])) + ((!g830) & (!g1914) & (!g2125) & (g4299) & (!g4303) & (key[195])) + ((!g830) & (!g1914) & (!g2125) & (g4299) & (g4303) & (key[195])) + ((!g830) & (!g1914) & (g2125) & (!g4299) & (!g4303) & (key[195])) + ((!g830) & (!g1914) & (g2125) & (!g4299) & (g4303) & (key[195])) + ((!g830) & (!g1914) & (g2125) & (g4299) & (!g4303) & (key[195])) + ((!g830) & (!g1914) & (g2125) & (g4299) & (g4303) & (key[195])) + ((!g830) & (g1914) & (!g2125) & (!g4299) & (!g4303) & (key[195])) + ((!g830) & (g1914) & (!g2125) & (!g4299) & (g4303) & (key[195])) + ((!g830) & (g1914) & (!g2125) & (g4299) & (!g4303) & (key[195])) + ((!g830) & (g1914) & (!g2125) & (g4299) & (g4303) & (key[195])) + ((!g830) & (g1914) & (g2125) & (!g4299) & (!g4303) & (key[195])) + ((!g830) & (g1914) & (g2125) & (!g4299) & (g4303) & (key[195])) + ((!g830) & (g1914) & (g2125) & (g4299) & (!g4303) & (key[195])) + ((!g830) & (g1914) & (g2125) & (g4299) & (g4303) & (key[195])) + ((g830) & (!g1914) & (!g2125) & (!g4299) & (g4303) & (!key[195])) + ((g830) & (!g1914) & (!g2125) & (!g4299) & (g4303) & (key[195])) + ((g830) & (!g1914) & (!g2125) & (g4299) & (g4303) & (!key[195])) + ((g830) & (!g1914) & (!g2125) & (g4299) & (g4303) & (key[195])) + ((g830) & (!g1914) & (g2125) & (!g4299) & (!g4303) & (!key[195])) + ((g830) & (!g1914) & (g2125) & (!g4299) & (!g4303) & (key[195])) + ((g830) & (!g1914) & (g2125) & (g4299) & (!g4303) & (!key[195])) + ((g830) & (!g1914) & (g2125) & (g4299) & (!g4303) & (key[195])) + ((g830) & (g1914) & (!g2125) & (g4299) & (!g4303) & (!key[195])) + ((g830) & (g1914) & (!g2125) & (g4299) & (!g4303) & (key[195])) + ((g830) & (g1914) & (!g2125) & (g4299) & (g4303) & (!key[195])) + ((g830) & (g1914) & (!g2125) & (g4299) & (g4303) & (key[195])) + ((g830) & (g1914) & (g2125) & (!g4299) & (!g4303) & (!key[195])) + ((g830) & (g1914) & (g2125) & (!g4299) & (!g4303) & (key[195])) + ((g830) & (g1914) & (g2125) & (!g4299) & (g4303) & (!key[195])) + ((g830) & (g1914) & (g2125) & (!g4299) & (g4303) & (key[195])));
	assign g4305 = (((!g2713) & (!g2783) & (!g2733) & (g2785) & (!g4242)) + ((!g2713) & (!g2783) & (!g2733) & (g2785) & (g4242)) + ((!g2713) & (!g2783) & (g2733) & (!g2785) & (g4242)) + ((!g2713) & (!g2783) & (g2733) & (g2785) & (!g4242)) + ((!g2713) & (g2783) & (!g2733) & (!g2785) & (!g4242)) + ((!g2713) & (g2783) & (!g2733) & (!g2785) & (g4242)) + ((!g2713) & (g2783) & (g2733) & (!g2785) & (!g4242)) + ((!g2713) & (g2783) & (g2733) & (g2785) & (g4242)) + ((g2713) & (!g2783) & (!g2733) & (!g2785) & (g4242)) + ((g2713) & (!g2783) & (!g2733) & (g2785) & (!g4242)) + ((g2713) & (!g2783) & (g2733) & (!g2785) & (!g4242)) + ((g2713) & (!g2783) & (g2733) & (!g2785) & (g4242)) + ((g2713) & (g2783) & (!g2733) & (!g2785) & (!g4242)) + ((g2713) & (g2783) & (!g2733) & (g2785) & (g4242)) + ((g2713) & (g2783) & (g2733) & (g2785) & (!g4242)) + ((g2713) & (g2783) & (g2733) & (g2785) & (g4242)));
	assign g4306 = (((!g2661) & (!g2742) & (g2669) & (g2747) & (g4166)) + ((!g2661) & (g2742) & (!g2669) & (g2747) & (!g4166)) + ((!g2661) & (g2742) & (!g2669) & (g2747) & (g4166)) + ((!g2661) & (g2742) & (g2669) & (!g2747) & (g4166)) + ((!g2661) & (g2742) & (g2669) & (g2747) & (!g4166)) + ((!g2661) & (g2742) & (g2669) & (g2747) & (g4166)) + ((g2661) & (!g2742) & (!g2669) & (g2747) & (g4166)) + ((g2661) & (!g2742) & (g2669) & (g2747) & (!g4166)) + ((g2661) & (!g2742) & (g2669) & (g2747) & (g4166)) + ((g2661) & (g2742) & (!g2669) & (!g2747) & (g4166)) + ((g2661) & (g2742) & (!g2669) & (g2747) & (!g4166)) + ((g2661) & (g2742) & (!g2669) & (g2747) & (g4166)) + ((g2661) & (g2742) & (g2669) & (!g2747) & (!g4166)) + ((g2661) & (g2742) & (g2669) & (!g2747) & (g4166)) + ((g2661) & (g2742) & (g2669) & (g2747) & (!g4166)) + ((g2661) & (g2742) & (g2669) & (g2747) & (g4166)));
	assign g4307 = (((!g1098) & (!g3504) & (!g2320)) + ((!g1098) & (g3504) & (g2320)) + ((g1098) & (!g3504) & (g2320)) + ((g1098) & (g3504) & (!g2320)));
	assign g4308 = (((!g2311) & (!g2317) & (!g3521)) + ((!g2311) & (g2317) & (g3521)) + ((g2311) & (!g2317) & (g3521)) + ((g2311) & (g2317) & (!g3521)));
	assign g4309 = (((!g830) & (!g1914) & (!g2129) & (!g4307) & (!g4308) & (key[49])) + ((!g830) & (!g1914) & (!g2129) & (!g4307) & (g4308) & (key[49])) + ((!g830) & (!g1914) & (!g2129) & (g4307) & (!g4308) & (key[49])) + ((!g830) & (!g1914) & (!g2129) & (g4307) & (g4308) & (key[49])) + ((!g830) & (!g1914) & (g2129) & (!g4307) & (!g4308) & (key[49])) + ((!g830) & (!g1914) & (g2129) & (!g4307) & (g4308) & (key[49])) + ((!g830) & (!g1914) & (g2129) & (g4307) & (!g4308) & (key[49])) + ((!g830) & (!g1914) & (g2129) & (g4307) & (g4308) & (key[49])) + ((!g830) & (g1914) & (!g2129) & (!g4307) & (!g4308) & (key[49])) + ((!g830) & (g1914) & (!g2129) & (!g4307) & (g4308) & (key[49])) + ((!g830) & (g1914) & (!g2129) & (g4307) & (!g4308) & (key[49])) + ((!g830) & (g1914) & (!g2129) & (g4307) & (g4308) & (key[49])) + ((!g830) & (g1914) & (g2129) & (!g4307) & (!g4308) & (key[49])) + ((!g830) & (g1914) & (g2129) & (!g4307) & (g4308) & (key[49])) + ((!g830) & (g1914) & (g2129) & (g4307) & (!g4308) & (key[49])) + ((!g830) & (g1914) & (g2129) & (g4307) & (g4308) & (key[49])) + ((g830) & (!g1914) & (!g2129) & (!g4307) & (g4308) & (!key[49])) + ((g830) & (!g1914) & (!g2129) & (!g4307) & (g4308) & (key[49])) + ((g830) & (!g1914) & (!g2129) & (g4307) & (g4308) & (!key[49])) + ((g830) & (!g1914) & (!g2129) & (g4307) & (g4308) & (key[49])) + ((g830) & (!g1914) & (g2129) & (!g4307) & (!g4308) & (!key[49])) + ((g830) & (!g1914) & (g2129) & (!g4307) & (!g4308) & (key[49])) + ((g830) & (!g1914) & (g2129) & (g4307) & (!g4308) & (!key[49])) + ((g830) & (!g1914) & (g2129) & (g4307) & (!g4308) & (key[49])) + ((g830) & (g1914) & (!g2129) & (g4307) & (!g4308) & (!key[49])) + ((g830) & (g1914) & (!g2129) & (g4307) & (!g4308) & (key[49])) + ((g830) & (g1914) & (!g2129) & (g4307) & (g4308) & (!key[49])) + ((g830) & (g1914) & (!g2129) & (g4307) & (g4308) & (key[49])) + ((g830) & (g1914) & (g2129) & (!g4307) & (!g4308) & (!key[49])) + ((g830) & (g1914) & (g2129) & (!g4307) & (!g4308) & (key[49])) + ((g830) & (g1914) & (g2129) & (!g4307) & (g4308) & (!key[49])) + ((g830) & (g1914) & (g2129) & (!g4307) & (g4308) & (key[49])));
	assign g4310 = (((!g1944) & (g2104) & (g3745)) + ((g1944) & (!g2104) & (g3745)) + ((g1944) & (g2104) & (!g3745)) + ((g1944) & (g2104) & (g3745)));
	assign g4311 = (((!g1946) & (!g2153) & (g4310)) + ((!g1946) & (g2153) & (!g4310)) + ((g1946) & (!g2153) & (!g4310)) + ((g1946) & (g2153) & (g4310)));
	assign g4312 = (((!g830) & (!g2130) & (!g6800) & (key[81])) + ((!g830) & (!g2130) & (g6800) & (key[81])) + ((!g830) & (g2130) & (!g6800) & (key[81])) + ((!g830) & (g2130) & (g6800) & (key[81])) + ((g830) & (!g2130) & (g6800) & (!key[81])) + ((g830) & (!g2130) & (g6800) & (key[81])) + ((g830) & (g2130) & (!g6800) & (!key[81])) + ((g830) & (g2130) & (!g6800) & (key[81])));
	assign g4313 = (((!g3396) & (!g2311) & (!g2334)) + ((!g3396) & (g2311) & (g2334)) + ((g3396) & (!g2311) & (g2334)) + ((g3396) & (g2311) & (!g2334)));
	assign g4314 = (((!g1098) & (!g3414) & (!g2304)) + ((!g1098) & (g3414) & (g2304)) + ((g1098) & (!g3414) & (g2304)) + ((g1098) & (g3414) & (!g2304)));
	assign g8297 = (((!g5560) & (g5591) & (!g4315)) + ((!g5560) & (g5591) & (g4315)) + ((g5560) & (!g5591) & (g4315)) + ((g5560) & (g5591) & (g4315)));
	assign g4316 = (((!g830) & (!g1914) & (!g2133) & (!g4313) & (!g4314) & (g4315)) + ((!g830) & (!g1914) & (!g2133) & (!g4313) & (g4314) & (g4315)) + ((!g830) & (!g1914) & (!g2133) & (g4313) & (!g4314) & (g4315)) + ((!g830) & (!g1914) & (!g2133) & (g4313) & (g4314) & (g4315)) + ((!g830) & (!g1914) & (g2133) & (!g4313) & (!g4314) & (g4315)) + ((!g830) & (!g1914) & (g2133) & (!g4313) & (g4314) & (g4315)) + ((!g830) & (!g1914) & (g2133) & (g4313) & (!g4314) & (g4315)) + ((!g830) & (!g1914) & (g2133) & (g4313) & (g4314) & (g4315)) + ((!g830) & (g1914) & (!g2133) & (!g4313) & (!g4314) & (g4315)) + ((!g830) & (g1914) & (!g2133) & (!g4313) & (g4314) & (g4315)) + ((!g830) & (g1914) & (!g2133) & (g4313) & (!g4314) & (g4315)) + ((!g830) & (g1914) & (!g2133) & (g4313) & (g4314) & (g4315)) + ((!g830) & (g1914) & (g2133) & (!g4313) & (!g4314) & (g4315)) + ((!g830) & (g1914) & (g2133) & (!g4313) & (g4314) & (g4315)) + ((!g830) & (g1914) & (g2133) & (g4313) & (!g4314) & (g4315)) + ((!g830) & (g1914) & (g2133) & (g4313) & (g4314) & (g4315)) + ((g830) & (!g1914) & (!g2133) & (!g4313) & (g4314) & (!g4315)) + ((g830) & (!g1914) & (!g2133) & (!g4313) & (g4314) & (g4315)) + ((g830) & (!g1914) & (!g2133) & (g4313) & (g4314) & (!g4315)) + ((g830) & (!g1914) & (!g2133) & (g4313) & (g4314) & (g4315)) + ((g830) & (!g1914) & (g2133) & (!g4313) & (!g4314) & (!g4315)) + ((g830) & (!g1914) & (g2133) & (!g4313) & (!g4314) & (g4315)) + ((g830) & (!g1914) & (g2133) & (g4313) & (!g4314) & (!g4315)) + ((g830) & (!g1914) & (g2133) & (g4313) & (!g4314) & (g4315)) + ((g830) & (g1914) & (!g2133) & (g4313) & (!g4314) & (!g4315)) + ((g830) & (g1914) & (!g2133) & (g4313) & (!g4314) & (g4315)) + ((g830) & (g1914) & (!g2133) & (g4313) & (g4314) & (!g4315)) + ((g830) & (g1914) & (!g2133) & (g4313) & (g4314) & (g4315)) + ((g830) & (g1914) & (g2133) & (!g4313) & (!g4314) & (!g4315)) + ((g830) & (g1914) & (g2133) & (!g4313) & (!g4314) & (g4315)) + ((g830) & (g1914) & (g2133) & (!g4313) & (g4314) & (!g4315)) + ((g830) & (g1914) & (g2133) & (!g4313) & (g4314) & (g4315)));
	assign g4317 = (((!g1982) & (g2114) & (g3483)) + ((g1982) & (!g2114) & (g3483)) + ((g1982) & (g2114) & (!g3483)) + ((g1982) & (g2114) & (g3483)));
	assign g4318 = (((!g1984) & (!g2137) & (g4317)) + ((!g1984) & (g2137) & (!g4317)) + ((g1984) & (!g2137) & (!g4317)) + ((g1984) & (g2137) & (g4317)));
	assign g4319 = (((!g830) & (!g2134) & (!g6789) & (key[177])) + ((!g830) & (!g2134) & (g6789) & (key[177])) + ((!g830) & (g2134) & (!g6789) & (key[177])) + ((!g830) & (g2134) & (g6789) & (key[177])) + ((g830) & (!g2134) & (g6789) & (!key[177])) + ((g830) & (!g2134) & (g6789) & (key[177])) + ((g830) & (g2134) & (!g6789) & (!key[177])) + ((g830) & (g2134) & (!g6789) & (key[177])));
	assign g4320 = (((!g2956) & (!g3005) & (!g4183) & (!g4184) & (!g2968) & (!g3020)) + ((!g2956) & (!g3005) & (!g4183) & (!g4184) & (!g2968) & (g3020)) + ((!g2956) & (!g3005) & (!g4183) & (!g4184) & (g2968) & (!g3020)) + ((!g2956) & (!g3005) & (!g4183) & (!g4184) & (g2968) & (g3020)) + ((!g2956) & (!g3005) & (!g4183) & (g4184) & (!g2968) & (!g3020)) + ((!g2956) & (!g3005) & (!g4183) & (g4184) & (!g2968) & (g3020)) + ((!g2956) & (!g3005) & (!g4183) & (g4184) & (g2968) & (!g3020)) + ((!g2956) & (!g3005) & (g4183) & (!g4184) & (!g2968) & (!g3020)) + ((!g2956) & (!g3005) & (g4183) & (!g4184) & (!g2968) & (g3020)) + ((!g2956) & (!g3005) & (g4183) & (!g4184) & (g2968) & (!g3020)) + ((!g2956) & (!g3005) & (g4183) & (g4184) & (!g2968) & (!g3020)) + ((!g2956) & (!g3005) & (g4183) & (g4184) & (!g2968) & (g3020)) + ((!g2956) & (!g3005) & (g4183) & (g4184) & (g2968) & (!g3020)) + ((!g2956) & (g3005) & (!g4183) & (!g4184) & (!g2968) & (!g3020)) + ((!g2956) & (g3005) & (!g4183) & (!g4184) & (g2968) & (!g3020)) + ((!g2956) & (g3005) & (!g4183) & (g4184) & (!g2968) & (!g3020)) + ((!g2956) & (g3005) & (g4183) & (!g4184) & (!g2968) & (!g3020)) + ((!g2956) & (g3005) & (g4183) & (g4184) & (!g2968) & (!g3020)) + ((g2956) & (!g3005) & (!g4183) & (!g4184) & (!g2968) & (!g3020)) + ((g2956) & (!g3005) & (!g4183) & (!g4184) & (!g2968) & (g3020)) + ((g2956) & (!g3005) & (!g4183) & (!g4184) & (g2968) & (!g3020)) + ((g2956) & (!g3005) & (!g4183) & (g4184) & (!g2968) & (!g3020)) + ((g2956) & (!g3005) & (!g4183) & (g4184) & (g2968) & (!g3020)) + ((g2956) & (!g3005) & (g4183) & (!g4184) & (!g2968) & (!g3020)) + ((g2956) & (!g3005) & (g4183) & (!g4184) & (g2968) & (!g3020)) + ((g2956) & (!g3005) & (g4183) & (g4184) & (!g2968) & (!g3020)) + ((g2956) & (!g3005) & (g4183) & (g4184) & (g2968) & (!g3020)) + ((g2956) & (g3005) & (!g4183) & (!g4184) & (!g2968) & (!g3020)));
	assign g4321 = (((!g3050) & (!g4320) & (!g3056)) + ((!g3050) & (g4320) & (g3056)) + ((g3050) & (!g4320) & (g3056)) + ((g3050) & (g4320) & (!g3056)));
	assign g4322 = (((!g2650) & (!g2684) & (!g1778) & (g1814) & (!g4274)) + ((!g2650) & (!g2684) & (!g1778) & (g1814) & (g4274)) + ((!g2650) & (!g2684) & (g1778) & (!g1814) & (!g4274)) + ((!g2650) & (!g2684) & (g1778) & (g1814) & (g4274)) + ((!g2650) & (g2684) & (!g1778) & (!g1814) & (!g4274)) + ((!g2650) & (g2684) & (!g1778) & (!g1814) & (g4274)) + ((!g2650) & (g2684) & (g1778) & (!g1814) & (g4274)) + ((!g2650) & (g2684) & (g1778) & (g1814) & (!g4274)) + ((g2650) & (!g2684) & (!g1778) & (!g1814) & (!g4274)) + ((g2650) & (!g2684) & (!g1778) & (g1814) & (g4274)) + ((g2650) & (!g2684) & (g1778) & (!g1814) & (!g4274)) + ((g2650) & (!g2684) & (g1778) & (!g1814) & (g4274)) + ((g2650) & (g2684) & (!g1778) & (!g1814) & (g4274)) + ((g2650) & (g2684) & (!g1778) & (g1814) & (!g4274)) + ((g2650) & (g2684) & (g1778) & (g1814) & (!g4274)) + ((g2650) & (g2684) & (g1778) & (g1814) & (g4274)));
	assign g4323 = (((!g830) & (!g1914) & (!g2137) & (!g4321) & (!g4322) & (key[100])) + ((!g830) & (!g1914) & (!g2137) & (!g4321) & (g4322) & (key[100])) + ((!g830) & (!g1914) & (!g2137) & (g4321) & (!g4322) & (key[100])) + ((!g830) & (!g1914) & (!g2137) & (g4321) & (g4322) & (key[100])) + ((!g830) & (!g1914) & (g2137) & (!g4321) & (!g4322) & (key[100])) + ((!g830) & (!g1914) & (g2137) & (!g4321) & (g4322) & (key[100])) + ((!g830) & (!g1914) & (g2137) & (g4321) & (!g4322) & (key[100])) + ((!g830) & (!g1914) & (g2137) & (g4321) & (g4322) & (key[100])) + ((!g830) & (g1914) & (!g2137) & (!g4321) & (!g4322) & (key[100])) + ((!g830) & (g1914) & (!g2137) & (!g4321) & (g4322) & (key[100])) + ((!g830) & (g1914) & (!g2137) & (g4321) & (!g4322) & (key[100])) + ((!g830) & (g1914) & (!g2137) & (g4321) & (g4322) & (key[100])) + ((!g830) & (g1914) & (g2137) & (!g4321) & (!g4322) & (key[100])) + ((!g830) & (g1914) & (g2137) & (!g4321) & (g4322) & (key[100])) + ((!g830) & (g1914) & (g2137) & (g4321) & (!g4322) & (key[100])) + ((!g830) & (g1914) & (g2137) & (g4321) & (g4322) & (key[100])) + ((g830) & (!g1914) & (!g2137) & (!g4321) & (g4322) & (!key[100])) + ((g830) & (!g1914) & (!g2137) & (!g4321) & (g4322) & (key[100])) + ((g830) & (!g1914) & (!g2137) & (g4321) & (g4322) & (!key[100])) + ((g830) & (!g1914) & (!g2137) & (g4321) & (g4322) & (key[100])) + ((g830) & (!g1914) & (g2137) & (!g4321) & (!g4322) & (!key[100])) + ((g830) & (!g1914) & (g2137) & (!g4321) & (!g4322) & (key[100])) + ((g830) & (!g1914) & (g2137) & (g4321) & (!g4322) & (!key[100])) + ((g830) & (!g1914) & (g2137) & (g4321) & (!g4322) & (key[100])) + ((g830) & (g1914) & (!g2137) & (g4321) & (!g4322) & (!key[100])) + ((g830) & (g1914) & (!g2137) & (g4321) & (!g4322) & (key[100])) + ((g830) & (g1914) & (!g2137) & (g4321) & (g4322) & (!key[100])) + ((g830) & (g1914) & (!g2137) & (g4321) & (g4322) & (key[100])) + ((g830) & (g1914) & (g2137) & (!g4321) & (!g4322) & (!key[100])) + ((g830) & (g1914) & (g2137) & (!g4321) & (!g4322) & (key[100])) + ((g830) & (g1914) & (g2137) & (!g4321) & (g4322) & (!key[100])) + ((g830) & (g1914) & (g2137) & (!g4321) & (g4322) & (key[100])));
	assign g4324 = (((!g2100) & (!g2133) & (g2723) & (g2770) & (!g4190) & (g4191)) + ((!g2100) & (!g2133) & (g2723) & (g2770) & (g4190) & (!g4191)) + ((!g2100) & (!g2133) & (g2723) & (g2770) & (g4190) & (g4191)) + ((!g2100) & (g2133) & (!g2723) & (g2770) & (!g4190) & (!g4191)) + ((!g2100) & (g2133) & (!g2723) & (g2770) & (!g4190) & (g4191)) + ((!g2100) & (g2133) & (!g2723) & (g2770) & (g4190) & (!g4191)) + ((!g2100) & (g2133) & (!g2723) & (g2770) & (g4190) & (g4191)) + ((!g2100) & (g2133) & (g2723) & (!g2770) & (!g4190) & (g4191)) + ((!g2100) & (g2133) & (g2723) & (!g2770) & (g4190) & (!g4191)) + ((!g2100) & (g2133) & (g2723) & (!g2770) & (g4190) & (g4191)) + ((!g2100) & (g2133) & (g2723) & (g2770) & (!g4190) & (!g4191)) + ((!g2100) & (g2133) & (g2723) & (g2770) & (!g4190) & (g4191)) + ((!g2100) & (g2133) & (g2723) & (g2770) & (g4190) & (!g4191)) + ((!g2100) & (g2133) & (g2723) & (g2770) & (g4190) & (g4191)) + ((g2100) & (!g2133) & (!g2723) & (g2770) & (!g4190) & (g4191)) + ((g2100) & (!g2133) & (!g2723) & (g2770) & (g4190) & (!g4191)) + ((g2100) & (!g2133) & (!g2723) & (g2770) & (g4190) & (g4191)) + ((g2100) & (!g2133) & (g2723) & (g2770) & (!g4190) & (!g4191)) + ((g2100) & (!g2133) & (g2723) & (g2770) & (!g4190) & (g4191)) + ((g2100) & (!g2133) & (g2723) & (g2770) & (g4190) & (!g4191)) + ((g2100) & (!g2133) & (g2723) & (g2770) & (g4190) & (g4191)) + ((g2100) & (g2133) & (!g2723) & (!g2770) & (!g4190) & (g4191)) + ((g2100) & (g2133) & (!g2723) & (!g2770) & (g4190) & (!g4191)) + ((g2100) & (g2133) & (!g2723) & (!g2770) & (g4190) & (g4191)) + ((g2100) & (g2133) & (!g2723) & (g2770) & (!g4190) & (!g4191)) + ((g2100) & (g2133) & (!g2723) & (g2770) & (!g4190) & (g4191)) + ((g2100) & (g2133) & (!g2723) & (g2770) & (g4190) & (!g4191)) + ((g2100) & (g2133) & (!g2723) & (g2770) & (g4190) & (g4191)) + ((g2100) & (g2133) & (g2723) & (!g2770) & (!g4190) & (!g4191)) + ((g2100) & (g2133) & (g2723) & (!g2770) & (!g4190) & (g4191)) + ((g2100) & (g2133) & (g2723) & (!g2770) & (g4190) & (!g4191)) + ((g2100) & (g2133) & (g2723) & (!g2770) & (g4190) & (g4191)) + ((g2100) & (g2133) & (g2723) & (g2770) & (!g4190) & (!g4191)) + ((g2100) & (g2133) & (g2723) & (g2770) & (!g4190) & (g4191)) + ((g2100) & (g2133) & (g2723) & (g2770) & (g4190) & (!g4191)) + ((g2100) & (g2133) & (g2723) & (g2770) & (g4190) & (g4191)));
	assign g4325 = (((!g2129) & (g2776) & (g4263)) + ((g2129) & (!g2776) & (g4263)) + ((g2129) & (g2776) & (!g4263)) + ((g2129) & (g2776) & (g4263)));
	assign g4326 = (((!g2177) & (!g2807) & (g4325)) + ((!g2177) & (g2807) & (!g4325)) + ((g2177) & (!g2807) & (!g4325)) + ((g2177) & (g2807) & (g4325)));
	assign g4327 = (((!g3260) & (!g4277) & (!g3222) & (!g3301) & (g3305)) + ((!g3260) & (!g4277) & (!g3222) & (g3301) & (!g3305)) + ((!g3260) & (!g4277) & (g3222) & (!g3301) & (!g3305)) + ((!g3260) & (!g4277) & (g3222) & (g3301) & (g3305)) + ((!g3260) & (g4277) & (!g3222) & (!g3301) & (g3305)) + ((!g3260) & (g4277) & (!g3222) & (g3301) & (!g3305)) + ((!g3260) & (g4277) & (g3222) & (!g3301) & (g3305)) + ((!g3260) & (g4277) & (g3222) & (g3301) & (!g3305)) + ((g3260) & (!g4277) & (!g3222) & (!g3301) & (!g3305)) + ((g3260) & (!g4277) & (!g3222) & (g3301) & (g3305)) + ((g3260) & (!g4277) & (g3222) & (!g3301) & (!g3305)) + ((g3260) & (!g4277) & (g3222) & (g3301) & (g3305)) + ((g3260) & (g4277) & (!g3222) & (!g3301) & (g3305)) + ((g3260) & (g4277) & (!g3222) & (g3301) & (!g3305)) + ((g3260) & (g4277) & (g3222) & (!g3301) & (!g3305)) + ((g3260) & (g4277) & (g3222) & (g3301) & (g3305)));
	assign g4328 = (((!g2295) & (!g2343) & (!g2979) & (!g3007) & (!g4196) & (!g4197)) + ((!g2295) & (!g2343) & (!g2979) & (!g3007) & (!g4196) & (g4197)) + ((!g2295) & (!g2343) & (!g2979) & (!g3007) & (g4196) & (!g4197)) + ((!g2295) & (!g2343) & (!g2979) & (!g3007) & (g4196) & (g4197)) + ((!g2295) & (!g2343) & (!g2979) & (g3007) & (!g4196) & (!g4197)) + ((!g2295) & (!g2343) & (!g2979) & (g3007) & (!g4196) & (g4197)) + ((!g2295) & (!g2343) & (!g2979) & (g3007) & (g4196) & (!g4197)) + ((!g2295) & (!g2343) & (!g2979) & (g3007) & (g4196) & (g4197)) + ((!g2295) & (!g2343) & (g2979) & (!g3007) & (!g4196) & (!g4197)) + ((!g2295) & (!g2343) & (g2979) & (!g3007) & (!g4196) & (g4197)) + ((!g2295) & (!g2343) & (g2979) & (!g3007) & (g4196) & (!g4197)) + ((!g2295) & (!g2343) & (g2979) & (!g3007) & (g4196) & (g4197)) + ((!g2295) & (!g2343) & (g2979) & (g3007) & (!g4196) & (!g4197)) + ((!g2295) & (g2343) & (!g2979) & (!g3007) & (!g4196) & (!g4197)) + ((!g2295) & (g2343) & (!g2979) & (!g3007) & (!g4196) & (g4197)) + ((!g2295) & (g2343) & (!g2979) & (!g3007) & (g4196) & (!g4197)) + ((!g2295) & (g2343) & (!g2979) & (!g3007) & (g4196) & (g4197)) + ((!g2295) & (g2343) & (g2979) & (!g3007) & (!g4196) & (!g4197)) + ((g2295) & (!g2343) & (!g2979) & (!g3007) & (!g4196) & (!g4197)) + ((g2295) & (!g2343) & (!g2979) & (!g3007) & (!g4196) & (g4197)) + ((g2295) & (!g2343) & (!g2979) & (!g3007) & (g4196) & (!g4197)) + ((g2295) & (!g2343) & (!g2979) & (!g3007) & (g4196) & (g4197)) + ((g2295) & (!g2343) & (!g2979) & (g3007) & (!g4196) & (!g4197)) + ((g2295) & (!g2343) & (g2979) & (!g3007) & (!g4196) & (!g4197)) + ((g2295) & (!g2343) & (g2979) & (!g3007) & (!g4196) & (g4197)) + ((g2295) & (!g2343) & (g2979) & (!g3007) & (g4196) & (!g4197)) + ((g2295) & (!g2343) & (g2979) & (!g3007) & (g4196) & (g4197)) + ((g2295) & (g2343) & (!g2979) & (!g3007) & (!g4196) & (!g4197)));
	assign g4329 = (((!g2376) & (!g3061) & (!g4328)) + ((!g2376) & (g3061) & (g4328)) + ((g2376) & (!g3061) & (g4328)) + ((g2376) & (g3061) & (!g4328)));
	assign g4330 = (((!g830) & (!g1914) & (!g2147) & (!g4327) & (!g4329) & (nonce[4])) + ((!g830) & (!g1914) & (!g2147) & (!g4327) & (g4329) & (nonce[4])) + ((!g830) & (!g1914) & (!g2147) & (g4327) & (!g4329) & (nonce[4])) + ((!g830) & (!g1914) & (!g2147) & (g4327) & (g4329) & (nonce[4])) + ((!g830) & (!g1914) & (g2147) & (!g4327) & (!g4329) & (nonce[4])) + ((!g830) & (!g1914) & (g2147) & (!g4327) & (g4329) & (nonce[4])) + ((!g830) & (!g1914) & (g2147) & (g4327) & (!g4329) & (nonce[4])) + ((!g830) & (!g1914) & (g2147) & (g4327) & (g4329) & (nonce[4])) + ((!g830) & (g1914) & (!g2147) & (!g4327) & (!g4329) & (nonce[4])) + ((!g830) & (g1914) & (!g2147) & (!g4327) & (g4329) & (nonce[4])) + ((!g830) & (g1914) & (!g2147) & (g4327) & (!g4329) & (nonce[4])) + ((!g830) & (g1914) & (!g2147) & (g4327) & (g4329) & (nonce[4])) + ((!g830) & (g1914) & (g2147) & (!g4327) & (!g4329) & (nonce[4])) + ((!g830) & (g1914) & (g2147) & (!g4327) & (g4329) & (nonce[4])) + ((!g830) & (g1914) & (g2147) & (g4327) & (!g4329) & (nonce[4])) + ((!g830) & (g1914) & (g2147) & (g4327) & (g4329) & (nonce[4])) + ((g830) & (!g1914) & (!g2147) & (!g4327) & (g4329) & (!nonce[4])) + ((g830) & (!g1914) & (!g2147) & (!g4327) & (g4329) & (nonce[4])) + ((g830) & (!g1914) & (!g2147) & (g4327) & (g4329) & (!nonce[4])) + ((g830) & (!g1914) & (!g2147) & (g4327) & (g4329) & (nonce[4])) + ((g830) & (!g1914) & (g2147) & (!g4327) & (!g4329) & (!nonce[4])) + ((g830) & (!g1914) & (g2147) & (!g4327) & (!g4329) & (nonce[4])) + ((g830) & (!g1914) & (g2147) & (g4327) & (!g4329) & (!nonce[4])) + ((g830) & (!g1914) & (g2147) & (g4327) & (!g4329) & (nonce[4])) + ((g830) & (g1914) & (!g2147) & (g4327) & (!g4329) & (!nonce[4])) + ((g830) & (g1914) & (!g2147) & (g4327) & (!g4329) & (nonce[4])) + ((g830) & (g1914) & (!g2147) & (g4327) & (g4329) & (!nonce[4])) + ((g830) & (g1914) & (!g2147) & (g4327) & (g4329) & (nonce[4])) + ((g830) & (g1914) & (g2147) & (!g4327) & (!g4329) & (!nonce[4])) + ((g830) & (g1914) & (g2147) & (!g4327) & (!g4329) & (nonce[4])) + ((g830) & (g1914) & (g2147) & (!g4327) & (g4329) & (!nonce[4])) + ((g830) & (g1914) & (g2147) & (!g4327) & (g4329) & (nonce[4])));
	assign g4331 = (((!g2299) & (!g2348) & (!g4202) & (!g4203) & (!g2985) & (!g3015)) + ((!g2299) & (!g2348) & (!g4202) & (!g4203) & (!g2985) & (g3015)) + ((!g2299) & (!g2348) & (!g4202) & (!g4203) & (g2985) & (!g3015)) + ((!g2299) & (!g2348) & (!g4202) & (!g4203) & (g2985) & (g3015)) + ((!g2299) & (!g2348) & (!g4202) & (g4203) & (!g2985) & (!g3015)) + ((!g2299) & (!g2348) & (!g4202) & (g4203) & (!g2985) & (g3015)) + ((!g2299) & (!g2348) & (!g4202) & (g4203) & (g2985) & (!g3015)) + ((!g2299) & (!g2348) & (g4202) & (!g4203) & (!g2985) & (!g3015)) + ((!g2299) & (!g2348) & (g4202) & (!g4203) & (!g2985) & (g3015)) + ((!g2299) & (!g2348) & (g4202) & (!g4203) & (g2985) & (!g3015)) + ((!g2299) & (!g2348) & (g4202) & (g4203) & (!g2985) & (!g3015)) + ((!g2299) & (!g2348) & (g4202) & (g4203) & (!g2985) & (g3015)) + ((!g2299) & (!g2348) & (g4202) & (g4203) & (g2985) & (!g3015)) + ((!g2299) & (g2348) & (!g4202) & (!g4203) & (!g2985) & (!g3015)) + ((!g2299) & (g2348) & (!g4202) & (!g4203) & (g2985) & (!g3015)) + ((!g2299) & (g2348) & (!g4202) & (g4203) & (!g2985) & (!g3015)) + ((!g2299) & (g2348) & (g4202) & (!g4203) & (!g2985) & (!g3015)) + ((!g2299) & (g2348) & (g4202) & (g4203) & (!g2985) & (!g3015)) + ((g2299) & (!g2348) & (!g4202) & (!g4203) & (!g2985) & (!g3015)) + ((g2299) & (!g2348) & (!g4202) & (!g4203) & (!g2985) & (g3015)) + ((g2299) & (!g2348) & (!g4202) & (!g4203) & (g2985) & (!g3015)) + ((g2299) & (!g2348) & (!g4202) & (g4203) & (!g2985) & (!g3015)) + ((g2299) & (!g2348) & (!g4202) & (g4203) & (g2985) & (!g3015)) + ((g2299) & (!g2348) & (g4202) & (!g4203) & (!g2985) & (!g3015)) + ((g2299) & (!g2348) & (g4202) & (!g4203) & (g2985) & (!g3015)) + ((g2299) & (!g2348) & (g4202) & (g4203) & (!g2985) & (!g3015)) + ((g2299) & (!g2348) & (g4202) & (g4203) & (g2985) & (!g3015)) + ((g2299) & (g2348) & (!g4202) & (!g4203) & (!g2985) & (!g3015)));
	assign g4332 = (((!g2379) & (!g4331) & (!g3064)) + ((!g2379) & (g4331) & (g3064)) + ((g2379) & (!g4331) & (g3064)) + ((g2379) & (g4331) & (!g3064)));
	assign g4333 = (((!g3235) & (!g4293) & (!g3240) & (!g3295) & (g3303)) + ((!g3235) & (!g4293) & (!g3240) & (g3295) & (!g3303)) + ((!g3235) & (!g4293) & (g3240) & (!g3295) & (!g3303)) + ((!g3235) & (!g4293) & (g3240) & (g3295) & (g3303)) + ((!g3235) & (g4293) & (!g3240) & (!g3295) & (g3303)) + ((!g3235) & (g4293) & (!g3240) & (g3295) & (!g3303)) + ((!g3235) & (g4293) & (g3240) & (!g3295) & (g3303)) + ((!g3235) & (g4293) & (g3240) & (g3295) & (!g3303)) + ((g3235) & (!g4293) & (!g3240) & (!g3295) & (!g3303)) + ((g3235) & (!g4293) & (!g3240) & (g3295) & (g3303)) + ((g3235) & (!g4293) & (g3240) & (!g3295) & (!g3303)) + ((g3235) & (!g4293) & (g3240) & (g3295) & (g3303)) + ((g3235) & (g4293) & (!g3240) & (!g3295) & (g3303)) + ((g3235) & (g4293) & (!g3240) & (g3295) & (!g3303)) + ((g3235) & (g4293) & (g3240) & (!g3295) & (!g3303)) + ((g3235) & (g4293) & (g3240) & (g3295) & (g3303)));
	assign g4334 = (((!g830) & (!g1914) & (!g2150) & (!g4332) & (!g4333) & (key[228])) + ((!g830) & (!g1914) & (!g2150) & (!g4332) & (g4333) & (key[228])) + ((!g830) & (!g1914) & (!g2150) & (g4332) & (!g4333) & (key[228])) + ((!g830) & (!g1914) & (!g2150) & (g4332) & (g4333) & (key[228])) + ((!g830) & (!g1914) & (g2150) & (!g4332) & (!g4333) & (key[228])) + ((!g830) & (!g1914) & (g2150) & (!g4332) & (g4333) & (key[228])) + ((!g830) & (!g1914) & (g2150) & (g4332) & (!g4333) & (key[228])) + ((!g830) & (!g1914) & (g2150) & (g4332) & (g4333) & (key[228])) + ((!g830) & (g1914) & (!g2150) & (!g4332) & (!g4333) & (key[228])) + ((!g830) & (g1914) & (!g2150) & (!g4332) & (g4333) & (key[228])) + ((!g830) & (g1914) & (!g2150) & (g4332) & (!g4333) & (key[228])) + ((!g830) & (g1914) & (!g2150) & (g4332) & (g4333) & (key[228])) + ((!g830) & (g1914) & (g2150) & (!g4332) & (!g4333) & (key[228])) + ((!g830) & (g1914) & (g2150) & (!g4332) & (g4333) & (key[228])) + ((!g830) & (g1914) & (g2150) & (g4332) & (!g4333) & (key[228])) + ((!g830) & (g1914) & (g2150) & (g4332) & (g4333) & (key[228])) + ((g830) & (!g1914) & (!g2150) & (!g4332) & (g4333) & (!key[228])) + ((g830) & (!g1914) & (!g2150) & (!g4332) & (g4333) & (key[228])) + ((g830) & (!g1914) & (!g2150) & (g4332) & (g4333) & (!key[228])) + ((g830) & (!g1914) & (!g2150) & (g4332) & (g4333) & (key[228])) + ((g830) & (!g1914) & (g2150) & (!g4332) & (!g4333) & (!key[228])) + ((g830) & (!g1914) & (g2150) & (!g4332) & (!g4333) & (key[228])) + ((g830) & (!g1914) & (g2150) & (g4332) & (!g4333) & (!key[228])) + ((g830) & (!g1914) & (g2150) & (g4332) & (!g4333) & (key[228])) + ((g830) & (g1914) & (!g2150) & (g4332) & (!g4333) & (!key[228])) + ((g830) & (g1914) & (!g2150) & (g4332) & (!g4333) & (key[228])) + ((g830) & (g1914) & (!g2150) & (g4332) & (g4333) & (!key[228])) + ((g830) & (g1914) & (!g2150) & (g4332) & (g4333) & (key[228])) + ((g830) & (g1914) & (g2150) & (!g4332) & (!g4333) & (!key[228])) + ((g830) & (g1914) & (g2150) & (!g4332) & (!g4333) & (key[228])) + ((g830) & (g1914) & (g2150) & (!g4332) & (g4333) & (!key[228])) + ((g830) & (g1914) & (g2150) & (!g4332) & (g4333) & (key[228])));
	assign g4335 = (((!g2648) & (!g2679) & (!g1778) & (g1814) & (!g4258)) + ((!g2648) & (!g2679) & (!g1778) & (g1814) & (g4258)) + ((!g2648) & (!g2679) & (g1778) & (!g1814) & (!g4258)) + ((!g2648) & (!g2679) & (g1778) & (g1814) & (g4258)) + ((!g2648) & (g2679) & (!g1778) & (!g1814) & (!g4258)) + ((!g2648) & (g2679) & (!g1778) & (!g1814) & (g4258)) + ((!g2648) & (g2679) & (g1778) & (!g1814) & (g4258)) + ((!g2648) & (g2679) & (g1778) & (g1814) & (!g4258)) + ((g2648) & (!g2679) & (!g1778) & (!g1814) & (!g4258)) + ((g2648) & (!g2679) & (!g1778) & (g1814) & (g4258)) + ((g2648) & (!g2679) & (g1778) & (!g1814) & (!g4258)) + ((g2648) & (!g2679) & (g1778) & (!g1814) & (g4258)) + ((g2648) & (g2679) & (!g1778) & (!g1814) & (g4258)) + ((g2648) & (g2679) & (!g1778) & (g1814) & (!g4258)) + ((g2648) & (g2679) & (g1778) & (g1814) & (!g4258)) + ((g2648) & (g2679) & (g1778) & (g1814) & (g4258)));
	assign g4336 = (((!g2938) & (!g3011) & (!g2985) & (!g4210) & (!g4211) & (!g3015)) + ((!g2938) & (!g3011) & (!g2985) & (!g4210) & (!g4211) & (g3015)) + ((!g2938) & (!g3011) & (!g2985) & (!g4210) & (g4211) & (!g3015)) + ((!g2938) & (!g3011) & (!g2985) & (!g4210) & (g4211) & (g3015)) + ((!g2938) & (!g3011) & (!g2985) & (g4210) & (!g4211) & (!g3015)) + ((!g2938) & (!g3011) & (!g2985) & (g4210) & (!g4211) & (g3015)) + ((!g2938) & (!g3011) & (!g2985) & (g4210) & (g4211) & (!g3015)) + ((!g2938) & (!g3011) & (!g2985) & (g4210) & (g4211) & (g3015)) + ((!g2938) & (!g3011) & (g2985) & (!g4210) & (!g4211) & (!g3015)) + ((!g2938) & (!g3011) & (g2985) & (!g4210) & (!g4211) & (g3015)) + ((!g2938) & (!g3011) & (g2985) & (!g4210) & (g4211) & (!g3015)) + ((!g2938) & (!g3011) & (g2985) & (g4210) & (!g4211) & (!g3015)) + ((!g2938) & (!g3011) & (g2985) & (g4210) & (g4211) & (!g3015)) + ((!g2938) & (g3011) & (!g2985) & (!g4210) & (!g4211) & (!g3015)) + ((!g2938) & (g3011) & (!g2985) & (!g4210) & (g4211) & (!g3015)) + ((!g2938) & (g3011) & (!g2985) & (g4210) & (!g4211) & (!g3015)) + ((!g2938) & (g3011) & (!g2985) & (g4210) & (g4211) & (!g3015)) + ((!g2938) & (g3011) & (g2985) & (!g4210) & (!g4211) & (!g3015)) + ((g2938) & (!g3011) & (!g2985) & (!g4210) & (!g4211) & (!g3015)) + ((g2938) & (!g3011) & (!g2985) & (!g4210) & (!g4211) & (g3015)) + ((g2938) & (!g3011) & (!g2985) & (!g4210) & (g4211) & (!g3015)) + ((g2938) & (!g3011) & (!g2985) & (g4210) & (!g4211) & (!g3015)) + ((g2938) & (!g3011) & (!g2985) & (g4210) & (g4211) & (!g3015)) + ((g2938) & (!g3011) & (g2985) & (!g4210) & (!g4211) & (!g3015)) + ((g2938) & (!g3011) & (g2985) & (!g4210) & (g4211) & (!g3015)) + ((g2938) & (!g3011) & (g2985) & (g4210) & (!g4211) & (!g3015)) + ((g2938) & (!g3011) & (g2985) & (g4210) & (g4211) & (!g3015)) + ((g2938) & (g3011) & (!g2985) & (!g4210) & (!g4211) & (!g3015)));
	assign g4337 = (((!g3041) & (!g3064) & (!g4336)) + ((!g3041) & (g3064) & (g4336)) + ((g3041) & (!g3064) & (g4336)) + ((g3041) & (g3064) & (!g4336)));
	assign g4338 = (((!g830) & (!g1914) & (!g2153) & (!g4335) & (!g4337) & (key[4])) + ((!g830) & (!g1914) & (!g2153) & (!g4335) & (g4337) & (key[4])) + ((!g830) & (!g1914) & (!g2153) & (g4335) & (!g4337) & (key[4])) + ((!g830) & (!g1914) & (!g2153) & (g4335) & (g4337) & (key[4])) + ((!g830) & (!g1914) & (g2153) & (!g4335) & (!g4337) & (key[4])) + ((!g830) & (!g1914) & (g2153) & (!g4335) & (g4337) & (key[4])) + ((!g830) & (!g1914) & (g2153) & (g4335) & (!g4337) & (key[4])) + ((!g830) & (!g1914) & (g2153) & (g4335) & (g4337) & (key[4])) + ((!g830) & (g1914) & (!g2153) & (!g4335) & (!g4337) & (key[4])) + ((!g830) & (g1914) & (!g2153) & (!g4335) & (g4337) & (key[4])) + ((!g830) & (g1914) & (!g2153) & (g4335) & (!g4337) & (key[4])) + ((!g830) & (g1914) & (!g2153) & (g4335) & (g4337) & (key[4])) + ((!g830) & (g1914) & (g2153) & (!g4335) & (!g4337) & (key[4])) + ((!g830) & (g1914) & (g2153) & (!g4335) & (g4337) & (key[4])) + ((!g830) & (g1914) & (g2153) & (g4335) & (!g4337) & (key[4])) + ((!g830) & (g1914) & (g2153) & (g4335) & (g4337) & (key[4])) + ((g830) & (!g1914) & (!g2153) & (!g4335) & (g4337) & (!key[4])) + ((g830) & (!g1914) & (!g2153) & (!g4335) & (g4337) & (key[4])) + ((g830) & (!g1914) & (!g2153) & (g4335) & (g4337) & (!key[4])) + ((g830) & (!g1914) & (!g2153) & (g4335) & (g4337) & (key[4])) + ((g830) & (!g1914) & (g2153) & (!g4335) & (!g4337) & (!key[4])) + ((g830) & (!g1914) & (g2153) & (!g4335) & (!g4337) & (key[4])) + ((g830) & (!g1914) & (g2153) & (g4335) & (!g4337) & (!key[4])) + ((g830) & (!g1914) & (g2153) & (g4335) & (!g4337) & (key[4])) + ((g830) & (g1914) & (!g2153) & (g4335) & (!g4337) & (!key[4])) + ((g830) & (g1914) & (!g2153) & (g4335) & (!g4337) & (key[4])) + ((g830) & (g1914) & (!g2153) & (g4335) & (g4337) & (!key[4])) + ((g830) & (g1914) & (!g2153) & (g4335) & (g4337) & (key[4])) + ((g830) & (g1914) & (g2153) & (!g4335) & (!g4337) & (!key[4])) + ((g830) & (g1914) & (g2153) & (!g4335) & (!g4337) & (key[4])) + ((g830) & (g1914) & (g2153) & (!g4335) & (g4337) & (!key[4])) + ((g830) & (g1914) & (g2153) & (!g4335) & (g4337) & (key[4])));
	assign g4339 = (((!g2298) & (!g2347) & (!g2944) & (!g3018) & (!g4216) & (!g4217)) + ((!g2298) & (!g2347) & (!g2944) & (!g3018) & (!g4216) & (g4217)) + ((!g2298) & (!g2347) & (!g2944) & (!g3018) & (g4216) & (!g4217)) + ((!g2298) & (!g2347) & (!g2944) & (!g3018) & (g4216) & (g4217)) + ((!g2298) & (!g2347) & (!g2944) & (g3018) & (!g4216) & (!g4217)) + ((!g2298) & (!g2347) & (!g2944) & (g3018) & (!g4216) & (g4217)) + ((!g2298) & (!g2347) & (!g2944) & (g3018) & (g4216) & (!g4217)) + ((!g2298) & (!g2347) & (!g2944) & (g3018) & (g4216) & (g4217)) + ((!g2298) & (!g2347) & (g2944) & (!g3018) & (!g4216) & (!g4217)) + ((!g2298) & (!g2347) & (g2944) & (!g3018) & (!g4216) & (g4217)) + ((!g2298) & (!g2347) & (g2944) & (!g3018) & (g4216) & (!g4217)) + ((!g2298) & (!g2347) & (g2944) & (!g3018) & (g4216) & (g4217)) + ((!g2298) & (!g2347) & (g2944) & (g3018) & (!g4216) & (!g4217)) + ((!g2298) & (g2347) & (!g2944) & (!g3018) & (!g4216) & (!g4217)) + ((!g2298) & (g2347) & (!g2944) & (!g3018) & (!g4216) & (g4217)) + ((!g2298) & (g2347) & (!g2944) & (!g3018) & (g4216) & (!g4217)) + ((!g2298) & (g2347) & (!g2944) & (!g3018) & (g4216) & (g4217)) + ((!g2298) & (g2347) & (g2944) & (!g3018) & (!g4216) & (!g4217)) + ((g2298) & (!g2347) & (!g2944) & (!g3018) & (!g4216) & (!g4217)) + ((g2298) & (!g2347) & (!g2944) & (!g3018) & (!g4216) & (g4217)) + ((g2298) & (!g2347) & (!g2944) & (!g3018) & (g4216) & (!g4217)) + ((g2298) & (!g2347) & (!g2944) & (!g3018) & (g4216) & (g4217)) + ((g2298) & (!g2347) & (!g2944) & (g3018) & (!g4216) & (!g4217)) + ((g2298) & (!g2347) & (g2944) & (!g3018) & (!g4216) & (!g4217)) + ((g2298) & (!g2347) & (g2944) & (!g3018) & (!g4216) & (g4217)) + ((g2298) & (!g2347) & (g2944) & (!g3018) & (g4216) & (!g4217)) + ((g2298) & (!g2347) & (g2944) & (!g3018) & (g4216) & (g4217)) + ((g2298) & (g2347) & (!g2944) & (!g3018) & (!g4216) & (!g4217)));
	assign g4340 = (((!g2378) & (!g3044) & (!g4339)) + ((!g2378) & (g3044) & (g4339)) + ((g2378) & (!g3044) & (g4339)) + ((g2378) & (g3044) & (!g4339)));
	assign g4341 = (((!g4265) & (!g3250) & (!g3260) & (!g3305) & (g3291)) + ((!g4265) & (!g3250) & (!g3260) & (g3305) & (!g3291)) + ((!g4265) & (!g3250) & (g3260) & (!g3305) & (!g3291)) + ((!g4265) & (!g3250) & (g3260) & (g3305) & (g3291)) + ((!g4265) & (g3250) & (!g3260) & (!g3305) & (!g3291)) + ((!g4265) & (g3250) & (!g3260) & (g3305) & (g3291)) + ((!g4265) & (g3250) & (g3260) & (!g3305) & (!g3291)) + ((!g4265) & (g3250) & (g3260) & (g3305) & (g3291)) + ((g4265) & (!g3250) & (!g3260) & (!g3305) & (g3291)) + ((g4265) & (!g3250) & (!g3260) & (g3305) & (!g3291)) + ((g4265) & (!g3250) & (g3260) & (!g3305) & (g3291)) + ((g4265) & (!g3250) & (g3260) & (g3305) & (!g3291)) + ((g4265) & (g3250) & (!g3260) & (!g3305) & (g3291)) + ((g4265) & (g3250) & (!g3260) & (g3305) & (!g3291)) + ((g4265) & (g3250) & (g3260) & (!g3305) & (!g3291)) + ((g4265) & (g3250) & (g3260) & (g3305) & (g3291)));
	assign g8298 = (((!g5560) & (g5593) & (!g4342)) + ((!g5560) & (g5593) & (g4342)) + ((g5560) & (!g5593) & (g4342)) + ((g5560) & (g5593) & (g4342)));
	assign g4343 = (((!g830) & (!g1914) & (!g2156) & (!g4340) & (!g4341) & (g4342)) + ((!g830) & (!g1914) & (!g2156) & (!g4340) & (g4341) & (g4342)) + ((!g830) & (!g1914) & (!g2156) & (g4340) & (!g4341) & (g4342)) + ((!g830) & (!g1914) & (!g2156) & (g4340) & (g4341) & (g4342)) + ((!g830) & (!g1914) & (g2156) & (!g4340) & (!g4341) & (g4342)) + ((!g830) & (!g1914) & (g2156) & (!g4340) & (g4341) & (g4342)) + ((!g830) & (!g1914) & (g2156) & (g4340) & (!g4341) & (g4342)) + ((!g830) & (!g1914) & (g2156) & (g4340) & (g4341) & (g4342)) + ((!g830) & (g1914) & (!g2156) & (!g4340) & (!g4341) & (g4342)) + ((!g830) & (g1914) & (!g2156) & (!g4340) & (g4341) & (g4342)) + ((!g830) & (g1914) & (!g2156) & (g4340) & (!g4341) & (g4342)) + ((!g830) & (g1914) & (!g2156) & (g4340) & (g4341) & (g4342)) + ((!g830) & (g1914) & (g2156) & (!g4340) & (!g4341) & (g4342)) + ((!g830) & (g1914) & (g2156) & (!g4340) & (g4341) & (g4342)) + ((!g830) & (g1914) & (g2156) & (g4340) & (!g4341) & (g4342)) + ((!g830) & (g1914) & (g2156) & (g4340) & (g4341) & (g4342)) + ((g830) & (!g1914) & (!g2156) & (!g4340) & (g4341) & (!g4342)) + ((g830) & (!g1914) & (!g2156) & (!g4340) & (g4341) & (g4342)) + ((g830) & (!g1914) & (!g2156) & (g4340) & (g4341) & (!g4342)) + ((g830) & (!g1914) & (!g2156) & (g4340) & (g4341) & (g4342)) + ((g830) & (!g1914) & (g2156) & (!g4340) & (!g4341) & (!g4342)) + ((g830) & (!g1914) & (g2156) & (!g4340) & (!g4341) & (g4342)) + ((g830) & (!g1914) & (g2156) & (g4340) & (!g4341) & (!g4342)) + ((g830) & (!g1914) & (g2156) & (g4340) & (!g4341) & (g4342)) + ((g830) & (g1914) & (!g2156) & (g4340) & (!g4341) & (!g4342)) + ((g830) & (g1914) & (!g2156) & (g4340) & (!g4341) & (g4342)) + ((g830) & (g1914) & (!g2156) & (g4340) & (g4341) & (!g4342)) + ((g830) & (g1914) & (!g2156) & (g4340) & (g4341) & (g4342)) + ((g830) & (g1914) & (g2156) & (!g4340) & (!g4341) & (!g4342)) + ((g830) & (g1914) & (g2156) & (!g4340) & (!g4341) & (g4342)) + ((g830) & (g1914) & (g2156) & (!g4340) & (g4341) & (!g4342)) + ((g830) & (g1914) & (g2156) & (!g4340) & (g4341) & (g4342)));
	assign g4344 = (((!g2690) & (!g2774) & (g2747) & (g2780) & (!g4223) & (g4224)) + ((!g2690) & (!g2774) & (g2747) & (g2780) & (g4223) & (!g4224)) + ((!g2690) & (!g2774) & (g2747) & (g2780) & (g4223) & (g4224)) + ((!g2690) & (g2774) & (!g2747) & (g2780) & (!g4223) & (!g4224)) + ((!g2690) & (g2774) & (!g2747) & (g2780) & (!g4223) & (g4224)) + ((!g2690) & (g2774) & (!g2747) & (g2780) & (g4223) & (!g4224)) + ((!g2690) & (g2774) & (!g2747) & (g2780) & (g4223) & (g4224)) + ((!g2690) & (g2774) & (g2747) & (!g2780) & (!g4223) & (g4224)) + ((!g2690) & (g2774) & (g2747) & (!g2780) & (g4223) & (!g4224)) + ((!g2690) & (g2774) & (g2747) & (!g2780) & (g4223) & (g4224)) + ((!g2690) & (g2774) & (g2747) & (g2780) & (!g4223) & (!g4224)) + ((!g2690) & (g2774) & (g2747) & (g2780) & (!g4223) & (g4224)) + ((!g2690) & (g2774) & (g2747) & (g2780) & (g4223) & (!g4224)) + ((!g2690) & (g2774) & (g2747) & (g2780) & (g4223) & (g4224)) + ((g2690) & (!g2774) & (!g2747) & (g2780) & (!g4223) & (g4224)) + ((g2690) & (!g2774) & (!g2747) & (g2780) & (g4223) & (!g4224)) + ((g2690) & (!g2774) & (!g2747) & (g2780) & (g4223) & (g4224)) + ((g2690) & (!g2774) & (g2747) & (g2780) & (!g4223) & (!g4224)) + ((g2690) & (!g2774) & (g2747) & (g2780) & (!g4223) & (g4224)) + ((g2690) & (!g2774) & (g2747) & (g2780) & (g4223) & (!g4224)) + ((g2690) & (!g2774) & (g2747) & (g2780) & (g4223) & (g4224)) + ((g2690) & (g2774) & (!g2747) & (!g2780) & (!g4223) & (g4224)) + ((g2690) & (g2774) & (!g2747) & (!g2780) & (g4223) & (!g4224)) + ((g2690) & (g2774) & (!g2747) & (!g2780) & (g4223) & (g4224)) + ((g2690) & (g2774) & (!g2747) & (g2780) & (!g4223) & (!g4224)) + ((g2690) & (g2774) & (!g2747) & (g2780) & (!g4223) & (g4224)) + ((g2690) & (g2774) & (!g2747) & (g2780) & (g4223) & (!g4224)) + ((g2690) & (g2774) & (!g2747) & (g2780) & (g4223) & (g4224)) + ((g2690) & (g2774) & (g2747) & (!g2780) & (!g4223) & (!g4224)) + ((g2690) & (g2774) & (g2747) & (!g2780) & (!g4223) & (g4224)) + ((g2690) & (g2774) & (g2747) & (!g2780) & (g4223) & (!g4224)) + ((g2690) & (g2774) & (g2747) & (!g2780) & (g4223) & (g4224)) + ((g2690) & (g2774) & (g2747) & (g2780) & (!g4223) & (!g4224)) + ((g2690) & (g2774) & (g2747) & (g2780) & (!g4223) & (g4224)) + ((g2690) & (g2774) & (g2747) & (g2780) & (g4223) & (!g4224)) + ((g2690) & (g2774) & (g2747) & (g2780) & (g4223) & (g4224)));
	assign g4345 = (((!g2764) & (g2785) & (g4282)) + ((g2764) & (!g2785) & (g4282)) + ((g2764) & (g2785) & (!g4282)) + ((g2764) & (g2785) & (g4282)));
	assign g4346 = (((!g2813) & (!g2822) & (g4345)) + ((!g2813) & (g2822) & (!g4345)) + ((g2813) & (!g2822) & (!g4345)) + ((g2813) & (g2822) & (g4345)));
	assign g4347 = (((!g2556) & (!g3172) & (!g4297) & (!g4298)) + ((!g2556) & (!g3172) & (!g4297) & (g4298)) + ((!g2556) & (!g3172) & (g4297) & (!g4298)) + ((!g2556) & (!g3172) & (g4297) & (g4298)) + ((!g2556) & (g3172) & (!g4297) & (!g4298)) + ((g2556) & (!g3172) & (!g4297) & (!g4298)));
	assign g4348 = (((g1914) & (!g2602) & (!g3213) & (!g4347)) + ((g1914) & (!g2602) & (g3213) & (g4347)) + ((g1914) & (g2602) & (!g3213) & (g4347)) + ((g1914) & (g2602) & (g3213) & (!g4347)));
	assign g4349 = (((!g3163) & (!g3161) & (!g4301) & (!g4302)) + ((!g3163) & (!g3161) & (!g4301) & (g4302)) + ((!g3163) & (!g3161) & (g4301) & (!g4302)) + ((!g3163) & (!g3161) & (g4301) & (g4302)) + ((!g3163) & (g3161) & (!g4301) & (!g4302)) + ((g3163) & (!g3161) & (!g4301) & (!g4302)));
	assign g4350 = (((!g1914) & (!g3199) & (!g3187) & (!g4349)) + ((!g1914) & (!g3199) & (g3187) & (g4349)) + ((!g1914) & (g3199) & (!g3187) & (g4349)) + ((!g1914) & (g3199) & (g3187) & (!g4349)));
	assign g4351 = (((!g830) & (!g2162) & (!g4348) & (!g4350) & (key[196])) + ((!g830) & (!g2162) & (!g4348) & (g4350) & (key[196])) + ((!g830) & (!g2162) & (g4348) & (!g4350) & (key[196])) + ((!g830) & (!g2162) & (g4348) & (g4350) & (key[196])) + ((!g830) & (g2162) & (!g4348) & (!g4350) & (key[196])) + ((!g830) & (g2162) & (!g4348) & (g4350) & (key[196])) + ((!g830) & (g2162) & (g4348) & (!g4350) & (key[196])) + ((!g830) & (g2162) & (g4348) & (g4350) & (key[196])) + ((g830) & (!g2162) & (!g4348) & (g4350) & (!key[196])) + ((g830) & (!g2162) & (!g4348) & (g4350) & (key[196])) + ((g830) & (!g2162) & (g4348) & (!g4350) & (!key[196])) + ((g830) & (!g2162) & (g4348) & (!g4350) & (key[196])) + ((g830) & (!g2162) & (g4348) & (g4350) & (!key[196])) + ((g830) & (!g2162) & (g4348) & (g4350) & (key[196])) + ((g830) & (g2162) & (!g4348) & (!g4350) & (!key[196])) + ((g830) & (g2162) & (!g4348) & (!g4350) & (key[196])));
	assign g4352 = (((!g4269) & (!g3235) & (!g3255) & (!g3295) & (g3297)) + ((!g4269) & (!g3235) & (!g3255) & (g3295) & (!g3297)) + ((!g4269) & (!g3235) & (g3255) & (!g3295) & (!g3297)) + ((!g4269) & (!g3235) & (g3255) & (g3295) & (g3297)) + ((!g4269) & (g3235) & (!g3255) & (!g3295) & (!g3297)) + ((!g4269) & (g3235) & (!g3255) & (g3295) & (g3297)) + ((!g4269) & (g3235) & (g3255) & (!g3295) & (!g3297)) + ((!g4269) & (g3235) & (g3255) & (g3295) & (g3297)) + ((g4269) & (!g3235) & (!g3255) & (!g3295) & (g3297)) + ((g4269) & (!g3235) & (!g3255) & (g3295) & (!g3297)) + ((g4269) & (!g3235) & (g3255) & (!g3295) & (g3297)) + ((g4269) & (!g3235) & (g3255) & (g3295) & (!g3297)) + ((g4269) & (g3235) & (!g3255) & (!g3295) & (g3297)) + ((g4269) & (g3235) & (!g3255) & (g3295) & (!g3297)) + ((g4269) & (g3235) & (g3255) & (!g3295) & (!g3297)) + ((g4269) & (g3235) & (g3255) & (g3295) & (g3297)));
	assign g4353 = (((!g2296) & (!g2344) & (!g2968) & (!g4232) & (!g4233) & (!g3020)) + ((!g2296) & (!g2344) & (!g2968) & (!g4232) & (!g4233) & (g3020)) + ((!g2296) & (!g2344) & (!g2968) & (!g4232) & (g4233) & (!g3020)) + ((!g2296) & (!g2344) & (!g2968) & (!g4232) & (g4233) & (g3020)) + ((!g2296) & (!g2344) & (!g2968) & (g4232) & (!g4233) & (!g3020)) + ((!g2296) & (!g2344) & (!g2968) & (g4232) & (!g4233) & (g3020)) + ((!g2296) & (!g2344) & (!g2968) & (g4232) & (g4233) & (!g3020)) + ((!g2296) & (!g2344) & (!g2968) & (g4232) & (g4233) & (g3020)) + ((!g2296) & (!g2344) & (g2968) & (!g4232) & (!g4233) & (!g3020)) + ((!g2296) & (!g2344) & (g2968) & (!g4232) & (!g4233) & (g3020)) + ((!g2296) & (!g2344) & (g2968) & (!g4232) & (g4233) & (!g3020)) + ((!g2296) & (!g2344) & (g2968) & (g4232) & (!g4233) & (!g3020)) + ((!g2296) & (!g2344) & (g2968) & (g4232) & (g4233) & (!g3020)) + ((!g2296) & (g2344) & (!g2968) & (!g4232) & (!g4233) & (!g3020)) + ((!g2296) & (g2344) & (!g2968) & (!g4232) & (g4233) & (!g3020)) + ((!g2296) & (g2344) & (!g2968) & (g4232) & (!g4233) & (!g3020)) + ((!g2296) & (g2344) & (!g2968) & (g4232) & (g4233) & (!g3020)) + ((!g2296) & (g2344) & (g2968) & (!g4232) & (!g4233) & (!g3020)) + ((g2296) & (!g2344) & (!g2968) & (!g4232) & (!g4233) & (!g3020)) + ((g2296) & (!g2344) & (!g2968) & (!g4232) & (!g4233) & (g3020)) + ((g2296) & (!g2344) & (!g2968) & (!g4232) & (g4233) & (!g3020)) + ((g2296) & (!g2344) & (!g2968) & (g4232) & (!g4233) & (!g3020)) + ((g2296) & (!g2344) & (!g2968) & (g4232) & (g4233) & (!g3020)) + ((g2296) & (!g2344) & (g2968) & (!g4232) & (!g4233) & (!g3020)) + ((g2296) & (!g2344) & (g2968) & (!g4232) & (g4233) & (!g3020)) + ((g2296) & (!g2344) & (g2968) & (g4232) & (!g4233) & (!g3020)) + ((g2296) & (!g2344) & (g2968) & (g4232) & (g4233) & (!g3020)) + ((g2296) & (g2344) & (!g2968) & (!g4232) & (!g4233) & (!g3020)));
	assign g4354 = (((!g2377) & (!g3056) & (!g4353)) + ((!g2377) & (g3056) & (g4353)) + ((g2377) & (!g3056) & (g4353)) + ((g2377) & (g3056) & (!g4353)));
	assign g4355 = (((!g830) & (!g1914) & (!g2167) & (!g4352) & (!g4354) & (key[132])) + ((!g830) & (!g1914) & (!g2167) & (!g4352) & (g4354) & (key[132])) + ((!g830) & (!g1914) & (!g2167) & (g4352) & (!g4354) & (key[132])) + ((!g830) & (!g1914) & (!g2167) & (g4352) & (g4354) & (key[132])) + ((!g830) & (!g1914) & (g2167) & (!g4352) & (!g4354) & (key[132])) + ((!g830) & (!g1914) & (g2167) & (!g4352) & (g4354) & (key[132])) + ((!g830) & (!g1914) & (g2167) & (g4352) & (!g4354) & (key[132])) + ((!g830) & (!g1914) & (g2167) & (g4352) & (g4354) & (key[132])) + ((!g830) & (g1914) & (!g2167) & (!g4352) & (!g4354) & (key[132])) + ((!g830) & (g1914) & (!g2167) & (!g4352) & (g4354) & (key[132])) + ((!g830) & (g1914) & (!g2167) & (g4352) & (!g4354) & (key[132])) + ((!g830) & (g1914) & (!g2167) & (g4352) & (g4354) & (key[132])) + ((!g830) & (g1914) & (g2167) & (!g4352) & (!g4354) & (key[132])) + ((!g830) & (g1914) & (g2167) & (!g4352) & (g4354) & (key[132])) + ((!g830) & (g1914) & (g2167) & (g4352) & (!g4354) & (key[132])) + ((!g830) & (g1914) & (g2167) & (g4352) & (g4354) & (key[132])) + ((g830) & (!g1914) & (!g2167) & (!g4352) & (g4354) & (!key[132])) + ((g830) & (!g1914) & (!g2167) & (!g4352) & (g4354) & (key[132])) + ((g830) & (!g1914) & (!g2167) & (g4352) & (g4354) & (!key[132])) + ((g830) & (!g1914) & (!g2167) & (g4352) & (g4354) & (key[132])) + ((g830) & (!g1914) & (g2167) & (!g4352) & (!g4354) & (!key[132])) + ((g830) & (!g1914) & (g2167) & (!g4352) & (!g4354) & (key[132])) + ((g830) & (!g1914) & (g2167) & (g4352) & (!g4354) & (!key[132])) + ((g830) & (!g1914) & (g2167) & (g4352) & (!g4354) & (key[132])) + ((g830) & (g1914) & (!g2167) & (g4352) & (!g4354) & (!key[132])) + ((g830) & (g1914) & (!g2167) & (g4352) & (!g4354) & (key[132])) + ((g830) & (g1914) & (!g2167) & (g4352) & (g4354) & (!key[132])) + ((g830) & (g1914) & (!g2167) & (g4352) & (g4354) & (key[132])) + ((g830) & (g1914) & (g2167) & (!g4352) & (!g4354) & (!key[132])) + ((g830) & (g1914) & (g2167) & (!g4352) & (!g4354) & (key[132])) + ((g830) & (g1914) & (g2167) & (!g4352) & (g4354) & (!key[132])) + ((g830) & (g1914) & (g2167) & (!g4352) & (g4354) & (key[132])));
	assign g4356 = (((!g3163) & (!g3155) & (!g4284) & (!g4285)) + ((!g3163) & (!g3155) & (!g4284) & (g4285)) + ((!g3163) & (!g3155) & (g4284) & (!g4285)) + ((!g3163) & (!g3155) & (g4284) & (g4285)) + ((!g3163) & (g3155) & (!g4284) & (!g4285)) + ((g3163) & (!g3155) & (!g4284) & (!g4285)));
	assign g4357 = (((g1914) & (!g3199) & (!g3196) & (!g4356)) + ((g1914) & (!g3199) & (g3196) & (g4356)) + ((g1914) & (g3199) & (!g3196) & (g4356)) + ((g1914) & (g3199) & (g3196) & (!g4356)));
	assign g4358 = (((!g2552) & (!g3172) & (!g4288) & (!g4289)) + ((!g2552) & (!g3172) & (!g4288) & (g4289)) + ((!g2552) & (!g3172) & (g4288) & (!g4289)) + ((!g2552) & (!g3172) & (g4288) & (g4289)) + ((!g2552) & (g3172) & (!g4288) & (!g4289)) + ((g2552) & (!g3172) & (!g4288) & (!g4289)));
	assign g4359 = (((!g1914) & (!g2599) & (!g3213) & (!g4358)) + ((!g1914) & (!g2599) & (g3213) & (g4358)) + ((!g1914) & (g2599) & (!g3213) & (g4358)) + ((!g1914) & (g2599) & (g3213) & (!g4358)));
	assign g4360 = (((!g830) & (!g2170) & (!g4357) & (!g4359) & (nonce[36])) + ((!g830) & (!g2170) & (!g4357) & (g4359) & (nonce[36])) + ((!g830) & (!g2170) & (g4357) & (!g4359) & (nonce[36])) + ((!g830) & (!g2170) & (g4357) & (g4359) & (nonce[36])) + ((!g830) & (g2170) & (!g4357) & (!g4359) & (nonce[36])) + ((!g830) & (g2170) & (!g4357) & (g4359) & (nonce[36])) + ((!g830) & (g2170) & (g4357) & (!g4359) & (nonce[36])) + ((!g830) & (g2170) & (g4357) & (g4359) & (nonce[36])) + ((g830) & (!g2170) & (!g4357) & (g4359) & (!nonce[36])) + ((g830) & (!g2170) & (!g4357) & (g4359) & (nonce[36])) + ((g830) & (!g2170) & (g4357) & (!g4359) & (!nonce[36])) + ((g830) & (!g2170) & (g4357) & (!g4359) & (nonce[36])) + ((g830) & (!g2170) & (g4357) & (g4359) & (!nonce[36])) + ((g830) & (!g2170) & (g4357) & (g4359) & (nonce[36])) + ((g830) & (g2170) & (!g4357) & (!g4359) & (!nonce[36])) + ((g830) & (g2170) & (!g4357) & (!g4359) & (nonce[36])));
	assign g4361 = (((!g2713) & (!g2783) & (g2733) & (g2785) & (!g4240) & (g4241)) + ((!g2713) & (!g2783) & (g2733) & (g2785) & (g4240) & (!g4241)) + ((!g2713) & (!g2783) & (g2733) & (g2785) & (g4240) & (g4241)) + ((!g2713) & (g2783) & (!g2733) & (g2785) & (!g4240) & (!g4241)) + ((!g2713) & (g2783) & (!g2733) & (g2785) & (!g4240) & (g4241)) + ((!g2713) & (g2783) & (!g2733) & (g2785) & (g4240) & (!g4241)) + ((!g2713) & (g2783) & (!g2733) & (g2785) & (g4240) & (g4241)) + ((!g2713) & (g2783) & (g2733) & (!g2785) & (!g4240) & (g4241)) + ((!g2713) & (g2783) & (g2733) & (!g2785) & (g4240) & (!g4241)) + ((!g2713) & (g2783) & (g2733) & (!g2785) & (g4240) & (g4241)) + ((!g2713) & (g2783) & (g2733) & (g2785) & (!g4240) & (!g4241)) + ((!g2713) & (g2783) & (g2733) & (g2785) & (!g4240) & (g4241)) + ((!g2713) & (g2783) & (g2733) & (g2785) & (g4240) & (!g4241)) + ((!g2713) & (g2783) & (g2733) & (g2785) & (g4240) & (g4241)) + ((g2713) & (!g2783) & (!g2733) & (g2785) & (!g4240) & (g4241)) + ((g2713) & (!g2783) & (!g2733) & (g2785) & (g4240) & (!g4241)) + ((g2713) & (!g2783) & (!g2733) & (g2785) & (g4240) & (g4241)) + ((g2713) & (!g2783) & (g2733) & (g2785) & (!g4240) & (!g4241)) + ((g2713) & (!g2783) & (g2733) & (g2785) & (!g4240) & (g4241)) + ((g2713) & (!g2783) & (g2733) & (g2785) & (g4240) & (!g4241)) + ((g2713) & (!g2783) & (g2733) & (g2785) & (g4240) & (g4241)) + ((g2713) & (g2783) & (!g2733) & (!g2785) & (!g4240) & (g4241)) + ((g2713) & (g2783) & (!g2733) & (!g2785) & (g4240) & (!g4241)) + ((g2713) & (g2783) & (!g2733) & (!g2785) & (g4240) & (g4241)) + ((g2713) & (g2783) & (!g2733) & (g2785) & (!g4240) & (!g4241)) + ((g2713) & (g2783) & (!g2733) & (g2785) & (!g4240) & (g4241)) + ((g2713) & (g2783) & (!g2733) & (g2785) & (g4240) & (!g4241)) + ((g2713) & (g2783) & (!g2733) & (g2785) & (g4240) & (g4241)) + ((g2713) & (g2783) & (g2733) & (!g2785) & (!g4240) & (!g4241)) + ((g2713) & (g2783) & (g2733) & (!g2785) & (!g4240) & (g4241)) + ((g2713) & (g2783) & (g2733) & (!g2785) & (g4240) & (!g4241)) + ((g2713) & (g2783) & (g2733) & (!g2785) & (g4240) & (g4241)) + ((g2713) & (g2783) & (g2733) & (g2785) & (!g4240) & (!g4241)) + ((g2713) & (g2783) & (g2733) & (g2785) & (!g4240) & (g4241)) + ((g2713) & (g2783) & (g2733) & (g2785) & (g4240) & (!g4241)) + ((g2713) & (g2783) & (g2733) & (g2785) & (g4240) & (g4241)));
	assign g4362 = (((!g2772) & (g2780) & (g4306)) + ((g2772) & (!g2780) & (g4306)) + ((g2772) & (g2780) & (!g4306)) + ((g2772) & (g2780) & (g4306)));
	assign g4363 = (((!g2827) & (!g2830) & (g4362)) + ((!g2827) & (g2830) & (!g4362)) + ((g2827) & (!g2830) & (!g4362)) + ((g2827) & (g2830) & (g4362)));
	assign g4364 = (((!g1098) & (!g3504) & (g2320)) + ((g1098) & (!g3504) & (!g2320)) + ((g1098) & (!g3504) & (g2320)) + ((g1098) & (g3504) & (g2320)));
	assign g4365 = (((g1914) & (!g1132) & (!g4364) & (g2350)) + ((g1914) & (!g1132) & (g4364) & (!g2350)) + ((g1914) & (g1132) & (!g4364) & (!g2350)) + ((g1914) & (g1132) & (g4364) & (g2350)));
	assign g4366 = (((!g2311) & (g2317) & (!g3521)) + ((g2311) & (!g2317) & (!g3521)) + ((g2311) & (g2317) & (!g3521)) + ((g2311) & (g2317) & (g3521)));
	assign g4367 = (((!g1914) & (!g2354) & (!g2369) & (g4366)) + ((!g1914) & (!g2354) & (g2369) & (!g4366)) + ((!g1914) & (g2354) & (!g2369) & (!g4366)) + ((!g1914) & (g2354) & (g2369) & (g4366)));
	assign g4368 = (((!g830) & (!g2177) & (!g4365) & (!g4367) & (key[50])) + ((!g830) & (!g2177) & (!g4365) & (g4367) & (key[50])) + ((!g830) & (!g2177) & (g4365) & (!g4367) & (key[50])) + ((!g830) & (!g2177) & (g4365) & (g4367) & (key[50])) + ((!g830) & (g2177) & (!g4365) & (!g4367) & (key[50])) + ((!g830) & (g2177) & (!g4365) & (g4367) & (key[50])) + ((!g830) & (g2177) & (g4365) & (!g4367) & (key[50])) + ((!g830) & (g2177) & (g4365) & (g4367) & (key[50])) + ((g830) & (!g2177) & (!g4365) & (g4367) & (!key[50])) + ((g830) & (!g2177) & (!g4365) & (g4367) & (key[50])) + ((g830) & (!g2177) & (g4365) & (!g4367) & (!key[50])) + ((g830) & (!g2177) & (g4365) & (!g4367) & (key[50])) + ((g830) & (!g2177) & (g4365) & (g4367) & (!key[50])) + ((g830) & (!g2177) & (g4365) & (g4367) & (key[50])) + ((g830) & (g2177) & (!g4365) & (!g4367) & (!key[50])) + ((g830) & (g2177) & (!g4365) & (!g4367) & (key[50])));
	assign g4369 = (((!g3765) & (!g3766)));
	assign g4370 = (((!g1946) & (!g1948) & (!g2153) & (g2184) & (!g4310)) + ((!g1946) & (!g1948) & (!g2153) & (g2184) & (g4310)) + ((!g1946) & (!g1948) & (g2153) & (!g2184) & (g4310)) + ((!g1946) & (!g1948) & (g2153) & (g2184) & (!g4310)) + ((!g1946) & (g1948) & (!g2153) & (!g2184) & (!g4310)) + ((!g1946) & (g1948) & (!g2153) & (!g2184) & (g4310)) + ((!g1946) & (g1948) & (g2153) & (!g2184) & (!g4310)) + ((!g1946) & (g1948) & (g2153) & (g2184) & (g4310)) + ((g1946) & (!g1948) & (!g2153) & (!g2184) & (g4310)) + ((g1946) & (!g1948) & (!g2153) & (g2184) & (!g4310)) + ((g1946) & (!g1948) & (g2153) & (!g2184) & (!g4310)) + ((g1946) & (!g1948) & (g2153) & (!g2184) & (g4310)) + ((g1946) & (g1948) & (!g2153) & (!g2184) & (!g4310)) + ((g1946) & (g1948) & (!g2153) & (g2184) & (g4310)) + ((g1946) & (g1948) & (g2153) & (g2184) & (!g4310)) + ((g1946) & (g1948) & (g2153) & (g2184) & (g4310)));
	assign g4371 = (((!g1914) & (!g2462) & (!g2509) & (!g4369) & (!g4370)) + ((!g1914) & (!g2462) & (!g2509) & (!g4369) & (g4370)) + ((!g1914) & (!g2462) & (g2509) & (g4369) & (!g4370)) + ((!g1914) & (!g2462) & (g2509) & (g4369) & (g4370)) + ((!g1914) & (g2462) & (!g2509) & (g4369) & (!g4370)) + ((!g1914) & (g2462) & (!g2509) & (g4369) & (g4370)) + ((!g1914) & (g2462) & (g2509) & (!g4369) & (!g4370)) + ((!g1914) & (g2462) & (g2509) & (!g4369) & (g4370)) + ((g1914) & (!g2462) & (!g2509) & (!g4369) & (g4370)) + ((g1914) & (!g2462) & (!g2509) & (g4369) & (g4370)) + ((g1914) & (!g2462) & (g2509) & (!g4369) & (g4370)) + ((g1914) & (!g2462) & (g2509) & (g4369) & (g4370)) + ((g1914) & (g2462) & (!g2509) & (!g4369) & (g4370)) + ((g1914) & (g2462) & (!g2509) & (g4369) & (g4370)) + ((g1914) & (g2462) & (g2509) & (!g4369) & (g4370)) + ((g1914) & (g2462) & (g2509) & (g4369) & (g4370)));
	assign g4372 = (((!g830) & (!g2178) & (!g4371) & (key[82])) + ((!g830) & (!g2178) & (g4371) & (key[82])) + ((!g830) & (g2178) & (!g4371) & (key[82])) + ((!g830) & (g2178) & (g4371) & (key[82])) + ((g830) & (!g2178) & (g4371) & (!key[82])) + ((g830) & (!g2178) & (g4371) & (key[82])) + ((g830) & (g2178) & (!g4371) & (!key[82])) + ((g830) & (g2178) & (!g4371) & (key[82])));
	assign g4373 = (((!g1098) & (!g3414) & (g2304)) + ((g1098) & (!g3414) & (!g2304)) + ((g1098) & (!g3414) & (g2304)) + ((g1098) & (g3414) & (g2304)));
	assign g4374 = (((!g3396) & (!g2311) & (g2334)) + ((!g3396) & (g2311) & (!g2334)) + ((!g3396) & (g2311) & (g2334)) + ((g3396) & (g2311) & (g2334)));
	assign g4375 = (((!g4374) & (!g2354) & (g2358)) + ((!g4374) & (g2354) & (!g2358)) + ((g4374) & (!g2354) & (!g2358)) + ((g4374) & (g2354) & (g2358)));
	assign g4376 = (((!g1914) & (!g1132) & (!g4373) & (g2360) & (!g4375)) + ((!g1914) & (!g1132) & (!g4373) & (g2360) & (g4375)) + ((!g1914) & (!g1132) & (g4373) & (!g2360) & (!g4375)) + ((!g1914) & (!g1132) & (g4373) & (!g2360) & (g4375)) + ((!g1914) & (g1132) & (!g4373) & (!g2360) & (!g4375)) + ((!g1914) & (g1132) & (!g4373) & (!g2360) & (g4375)) + ((!g1914) & (g1132) & (g4373) & (g2360) & (!g4375)) + ((!g1914) & (g1132) & (g4373) & (g2360) & (g4375)) + ((g1914) & (!g1132) & (!g4373) & (!g2360) & (g4375)) + ((g1914) & (!g1132) & (!g4373) & (g2360) & (g4375)) + ((g1914) & (!g1132) & (g4373) & (!g2360) & (g4375)) + ((g1914) & (!g1132) & (g4373) & (g2360) & (g4375)) + ((g1914) & (g1132) & (!g4373) & (!g2360) & (g4375)) + ((g1914) & (g1132) & (!g4373) & (g2360) & (g4375)) + ((g1914) & (g1132) & (g4373) & (!g2360) & (g4375)) + ((g1914) & (g1132) & (g4373) & (g2360) & (g4375)));
	assign g8299 = (((!g5560) & (g5594) & (!g4377)) + ((!g5560) & (g5594) & (g4377)) + ((g5560) & (!g5594) & (g4377)) + ((g5560) & (g5594) & (g4377)));
	assign g4378 = (((!g830) & (!g2180) & (!g4376) & (g4377)) + ((!g830) & (!g2180) & (g4376) & (g4377)) + ((!g830) & (g2180) & (!g4376) & (g4377)) + ((!g830) & (g2180) & (g4376) & (g4377)) + ((g830) & (!g2180) & (g4376) & (!g4377)) + ((g830) & (!g2180) & (g4376) & (g4377)) + ((g830) & (g2180) & (!g4376) & (!g4377)) + ((g830) & (g2180) & (!g4376) & (g4377)));
	assign g4379 = (((!g3471) & (!g3472)));
	assign g4380 = (((!g1984) & (!g1986) & (!g2137) & (g2194) & (!g4317)) + ((!g1984) & (!g1986) & (!g2137) & (g2194) & (g4317)) + ((!g1984) & (!g1986) & (g2137) & (!g2194) & (g4317)) + ((!g1984) & (!g1986) & (g2137) & (g2194) & (!g4317)) + ((!g1984) & (g1986) & (!g2137) & (!g2194) & (!g4317)) + ((!g1984) & (g1986) & (!g2137) & (!g2194) & (g4317)) + ((!g1984) & (g1986) & (g2137) & (!g2194) & (!g4317)) + ((!g1984) & (g1986) & (g2137) & (g2194) & (g4317)) + ((g1984) & (!g1986) & (!g2137) & (!g2194) & (g4317)) + ((g1984) & (!g1986) & (!g2137) & (g2194) & (!g4317)) + ((g1984) & (!g1986) & (g2137) & (!g2194) & (!g4317)) + ((g1984) & (!g1986) & (g2137) & (!g2194) & (g4317)) + ((g1984) & (g1986) & (!g2137) & (!g2194) & (!g4317)) + ((g1984) & (g1986) & (!g2137) & (g2194) & (g4317)) + ((g1984) & (g1986) & (g2137) & (g2194) & (!g4317)) + ((g1984) & (g1986) & (g2137) & (g2194) & (g4317)));
	assign g4381 = (((!g1914) & (!g4379) & (!g2497) & (!g2509) & (g4380)) + ((!g1914) & (!g4379) & (!g2497) & (g2509) & (g4380)) + ((!g1914) & (!g4379) & (g2497) & (!g2509) & (g4380)) + ((!g1914) & (!g4379) & (g2497) & (g2509) & (g4380)) + ((!g1914) & (g4379) & (!g2497) & (!g2509) & (g4380)) + ((!g1914) & (g4379) & (!g2497) & (g2509) & (g4380)) + ((!g1914) & (g4379) & (g2497) & (!g2509) & (g4380)) + ((!g1914) & (g4379) & (g2497) & (g2509) & (g4380)) + ((g1914) & (!g4379) & (!g2497) & (!g2509) & (!g4380)) + ((g1914) & (!g4379) & (!g2497) & (!g2509) & (g4380)) + ((g1914) & (!g4379) & (g2497) & (g2509) & (!g4380)) + ((g1914) & (!g4379) & (g2497) & (g2509) & (g4380)) + ((g1914) & (g4379) & (!g2497) & (g2509) & (!g4380)) + ((g1914) & (g4379) & (!g2497) & (g2509) & (g4380)) + ((g1914) & (g4379) & (g2497) & (!g2509) & (!g4380)) + ((g1914) & (g4379) & (g2497) & (!g2509) & (g4380)));
	assign g4382 = (((!g830) & (!g2181) & (!g4381) & (key[178])) + ((!g830) & (!g2181) & (g4381) & (key[178])) + ((!g830) & (g2181) & (!g4381) & (key[178])) + ((!g830) & (g2181) & (g4381) & (key[178])) + ((g830) & (!g2181) & (g4381) & (!key[178])) + ((g830) & (!g2181) & (g4381) & (key[178])) + ((g830) & (g2181) & (!g4381) & (!key[178])) + ((g830) & (g2181) & (!g4381) & (key[178])));
	assign g4383 = (((!g2648) & (!g2679) & (g1778) & (g1814) & (!g4258)) + ((!g2648) & (g2679) & (!g1778) & (g1814) & (!g4258)) + ((!g2648) & (g2679) & (!g1778) & (g1814) & (g4258)) + ((!g2648) & (g2679) & (g1778) & (!g1814) & (!g4258)) + ((!g2648) & (g2679) & (g1778) & (g1814) & (!g4258)) + ((!g2648) & (g2679) & (g1778) & (g1814) & (g4258)) + ((g2648) & (!g2679) & (!g1778) & (g1814) & (!g4258)) + ((g2648) & (!g2679) & (g1778) & (g1814) & (!g4258)) + ((g2648) & (!g2679) & (g1778) & (g1814) & (g4258)) + ((g2648) & (g2679) & (!g1778) & (!g1814) & (!g4258)) + ((g2648) & (g2679) & (!g1778) & (g1814) & (!g4258)) + ((g2648) & (g2679) & (!g1778) & (g1814) & (g4258)) + ((g2648) & (g2679) & (g1778) & (!g1814) & (!g4258)) + ((g2648) & (g2679) & (g1778) & (!g1814) & (g4258)) + ((g2648) & (g2679) & (g1778) & (g1814) & (!g4258)) + ((g2648) & (g2679) & (g1778) & (g1814) & (g4258)));
	assign g4384 = (((!g3041) & (g3064) & (!g4336)) + ((g3041) & (!g3064) & (!g4336)) + ((g3041) & (g3064) & (!g4336)) + ((g3041) & (g3064) & (g4336)));
	assign g4385 = (((!g830) & (key[5]) & (!g1914) & (!g4383) & (!g4384) & (!g5664)) + ((!g830) & (key[5]) & (!g1914) & (!g4383) & (!g4384) & (g5664)) + ((!g830) & (key[5]) & (!g1914) & (!g4383) & (g4384) & (!g5664)) + ((!g830) & (key[5]) & (!g1914) & (!g4383) & (g4384) & (g5664)) + ((!g830) & (key[5]) & (!g1914) & (g4383) & (!g4384) & (!g5664)) + ((!g830) & (key[5]) & (!g1914) & (g4383) & (!g4384) & (g5664)) + ((!g830) & (key[5]) & (!g1914) & (g4383) & (g4384) & (!g5664)) + ((!g830) & (key[5]) & (!g1914) & (g4383) & (g4384) & (g5664)) + ((!g830) & (key[5]) & (g1914) & (!g4383) & (!g4384) & (!g5664)) + ((!g830) & (key[5]) & (g1914) & (!g4383) & (!g4384) & (g5664)) + ((!g830) & (key[5]) & (g1914) & (!g4383) & (g4384) & (!g5664)) + ((!g830) & (key[5]) & (g1914) & (!g4383) & (g4384) & (g5664)) + ((!g830) & (key[5]) & (g1914) & (g4383) & (!g4384) & (!g5664)) + ((!g830) & (key[5]) & (g1914) & (g4383) & (!g4384) & (g5664)) + ((!g830) & (key[5]) & (g1914) & (g4383) & (g4384) & (!g5664)) + ((!g830) & (key[5]) & (g1914) & (g4383) & (g4384) & (g5664)) + ((g830) & (!key[5]) & (!g1914) & (!g4383) & (!g4384) & (!g5664)) + ((g830) & (!key[5]) & (!g1914) & (!g4383) & (g4384) & (g5664)) + ((g830) & (!key[5]) & (!g1914) & (g4383) & (!g4384) & (!g5664)) + ((g830) & (!key[5]) & (!g1914) & (g4383) & (g4384) & (g5664)) + ((g830) & (!key[5]) & (g1914) & (!g4383) & (!g4384) & (!g5664)) + ((g830) & (!key[5]) & (g1914) & (!g4383) & (g4384) & (!g5664)) + ((g830) & (!key[5]) & (g1914) & (g4383) & (!g4384) & (g5664)) + ((g830) & (!key[5]) & (g1914) & (g4383) & (g4384) & (g5664)) + ((g830) & (key[5]) & (!g1914) & (!g4383) & (!g4384) & (!g5664)) + ((g830) & (key[5]) & (!g1914) & (!g4383) & (g4384) & (g5664)) + ((g830) & (key[5]) & (!g1914) & (g4383) & (!g4384) & (!g5664)) + ((g830) & (key[5]) & (!g1914) & (g4383) & (g4384) & (g5664)) + ((g830) & (key[5]) & (g1914) & (!g4383) & (!g4384) & (!g5664)) + ((g830) & (key[5]) & (g1914) & (!g4383) & (g4384) & (!g5664)) + ((g830) & (key[5]) & (g1914) & (g4383) & (!g4384) & (g5664)) + ((g830) & (key[5]) & (g1914) & (g4383) & (g4384) & (g5664)));
	assign g4386 = (((!g2180) & (g2816) & (g4324)) + ((g2180) & (!g2816) & (g4324)) + ((g2180) & (g2816) & (!g4324)) + ((g2180) & (g2816) & (g4324)));
	assign g4387 = (((!g2177) & (!g2210) & (!g2807) & (g2857) & (!g4325)) + ((!g2177) & (!g2210) & (!g2807) & (g2857) & (g4325)) + ((!g2177) & (!g2210) & (g2807) & (!g2857) & (g4325)) + ((!g2177) & (!g2210) & (g2807) & (g2857) & (!g4325)) + ((!g2177) & (g2210) & (!g2807) & (!g2857) & (!g4325)) + ((!g2177) & (g2210) & (!g2807) & (!g2857) & (g4325)) + ((!g2177) & (g2210) & (g2807) & (!g2857) & (!g4325)) + ((!g2177) & (g2210) & (g2807) & (g2857) & (g4325)) + ((g2177) & (!g2210) & (!g2807) & (!g2857) & (g4325)) + ((g2177) & (!g2210) & (!g2807) & (g2857) & (!g4325)) + ((g2177) & (!g2210) & (g2807) & (!g2857) & (!g4325)) + ((g2177) & (!g2210) & (g2807) & (!g2857) & (g4325)) + ((g2177) & (g2210) & (!g2807) & (!g2857) & (!g4325)) + ((g2177) & (g2210) & (!g2807) & (g2857) & (g4325)) + ((g2177) & (g2210) & (g2807) & (g2857) & (!g4325)) + ((g2177) & (g2210) & (g2807) & (g2857) & (g4325)));
	assign g4388 = (((!g2378) & (g3044) & (!g4339)) + ((g2378) & (!g3044) & (!g4339)) + ((g2378) & (g3044) & (!g4339)) + ((g2378) & (g3044) & (g4339)));
	assign g4389 = (((!g4265) & (!g3250) & (!g3260) & (g3305) & (g3291)) + ((!g4265) & (!g3250) & (g3260) & (!g3305) & (g3291)) + ((!g4265) & (!g3250) & (g3260) & (g3305) & (!g3291)) + ((!g4265) & (!g3250) & (g3260) & (g3305) & (g3291)) + ((!g4265) & (g3250) & (!g3260) & (!g3305) & (g3291)) + ((!g4265) & (g3250) & (!g3260) & (g3305) & (!g3291)) + ((!g4265) & (g3250) & (!g3260) & (g3305) & (g3291)) + ((!g4265) & (g3250) & (g3260) & (!g3305) & (g3291)) + ((!g4265) & (g3250) & (g3260) & (g3305) & (!g3291)) + ((!g4265) & (g3250) & (g3260) & (g3305) & (g3291)) + ((g4265) & (!g3250) & (!g3260) & (g3305) & (g3291)) + ((g4265) & (!g3250) & (g3260) & (g3305) & (g3291)) + ((g4265) & (g3250) & (!g3260) & (g3305) & (g3291)) + ((g4265) & (g3250) & (g3260) & (!g3305) & (g3291)) + ((g4265) & (g3250) & (g3260) & (g3305) & (!g3291)) + ((g4265) & (g3250) & (g3260) & (g3305) & (g3291)));
	assign g8300 = (((!g5560) & (g5595) & (!g4390)) + ((!g5560) & (g5595) & (g4390)) + ((g5560) & (!g5595) & (g4390)) + ((g5560) & (g5595) & (g4390)));
	assign g4391 = (((!g830) & (g4390) & (!g1914) & (!g4389) & (!g4388) & (!g5666)) + ((!g830) & (g4390) & (!g1914) & (!g4389) & (!g4388) & (g5666)) + ((!g830) & (g4390) & (!g1914) & (!g4389) & (g4388) & (!g5666)) + ((!g830) & (g4390) & (!g1914) & (!g4389) & (g4388) & (g5666)) + ((!g830) & (g4390) & (!g1914) & (g4389) & (!g4388) & (!g5666)) + ((!g830) & (g4390) & (!g1914) & (g4389) & (!g4388) & (g5666)) + ((!g830) & (g4390) & (!g1914) & (g4389) & (g4388) & (!g5666)) + ((!g830) & (g4390) & (!g1914) & (g4389) & (g4388) & (g5666)) + ((!g830) & (g4390) & (g1914) & (!g4389) & (!g4388) & (!g5666)) + ((!g830) & (g4390) & (g1914) & (!g4389) & (!g4388) & (g5666)) + ((!g830) & (g4390) & (g1914) & (!g4389) & (g4388) & (!g5666)) + ((!g830) & (g4390) & (g1914) & (!g4389) & (g4388) & (g5666)) + ((!g830) & (g4390) & (g1914) & (g4389) & (!g4388) & (!g5666)) + ((!g830) & (g4390) & (g1914) & (g4389) & (!g4388) & (g5666)) + ((!g830) & (g4390) & (g1914) & (g4389) & (g4388) & (!g5666)) + ((!g830) & (g4390) & (g1914) & (g4389) & (g4388) & (g5666)) + ((g830) & (!g4390) & (!g1914) & (!g4389) & (!g4388) & (!g5666)) + ((g830) & (!g4390) & (!g1914) & (!g4389) & (g4388) & (!g5666)) + ((g830) & (!g4390) & (!g1914) & (g4389) & (!g4388) & (g5666)) + ((g830) & (!g4390) & (!g1914) & (g4389) & (g4388) & (g5666)) + ((g830) & (!g4390) & (g1914) & (!g4389) & (!g4388) & (!g5666)) + ((g830) & (!g4390) & (g1914) & (!g4389) & (g4388) & (g5666)) + ((g830) & (!g4390) & (g1914) & (g4389) & (!g4388) & (!g5666)) + ((g830) & (!g4390) & (g1914) & (g4389) & (g4388) & (g5666)) + ((g830) & (g4390) & (!g1914) & (!g4389) & (!g4388) & (!g5666)) + ((g830) & (g4390) & (!g1914) & (!g4389) & (g4388) & (!g5666)) + ((g830) & (g4390) & (!g1914) & (g4389) & (!g4388) & (g5666)) + ((g830) & (g4390) & (!g1914) & (g4389) & (g4388) & (g5666)) + ((g830) & (g4390) & (g1914) & (!g4389) & (!g4388) & (!g5666)) + ((g830) & (g4390) & (g1914) & (!g4389) & (g4388) & (g5666)) + ((g830) & (g4390) & (g1914) & (g4389) & (!g4388) & (!g5666)) + ((g830) & (g4390) & (g1914) & (g4389) & (g4388) & (g5666)));
	assign g4392 = (((!g4269) & (!g3235) & (!g3255) & (g3295) & (g3297)) + ((!g4269) & (!g3235) & (g3255) & (!g3295) & (g3297)) + ((!g4269) & (!g3235) & (g3255) & (g3295) & (!g3297)) + ((!g4269) & (!g3235) & (g3255) & (g3295) & (g3297)) + ((!g4269) & (g3235) & (!g3255) & (!g3295) & (g3297)) + ((!g4269) & (g3235) & (!g3255) & (g3295) & (!g3297)) + ((!g4269) & (g3235) & (!g3255) & (g3295) & (g3297)) + ((!g4269) & (g3235) & (g3255) & (!g3295) & (g3297)) + ((!g4269) & (g3235) & (g3255) & (g3295) & (!g3297)) + ((!g4269) & (g3235) & (g3255) & (g3295) & (g3297)) + ((g4269) & (!g3235) & (!g3255) & (g3295) & (g3297)) + ((g4269) & (!g3235) & (g3255) & (g3295) & (g3297)) + ((g4269) & (g3235) & (!g3255) & (g3295) & (g3297)) + ((g4269) & (g3235) & (g3255) & (!g3295) & (g3297)) + ((g4269) & (g3235) & (g3255) & (g3295) & (!g3297)) + ((g4269) & (g3235) & (g3255) & (g3295) & (g3297)));
	assign g4393 = (((!g2377) & (g3056) & (!g4353)) + ((g2377) & (!g3056) & (!g4353)) + ((g2377) & (g3056) & (!g4353)) + ((g2377) & (g3056) & (g4353)));
	assign g4394 = (((!g830) & (key[133]) & (!g1914) & (!g4392) & (!g4393) & (!g5667)) + ((!g830) & (key[133]) & (!g1914) & (!g4392) & (!g4393) & (g5667)) + ((!g830) & (key[133]) & (!g1914) & (!g4392) & (g4393) & (!g5667)) + ((!g830) & (key[133]) & (!g1914) & (!g4392) & (g4393) & (g5667)) + ((!g830) & (key[133]) & (!g1914) & (g4392) & (!g4393) & (!g5667)) + ((!g830) & (key[133]) & (!g1914) & (g4392) & (!g4393) & (g5667)) + ((!g830) & (key[133]) & (!g1914) & (g4392) & (g4393) & (!g5667)) + ((!g830) & (key[133]) & (!g1914) & (g4392) & (g4393) & (g5667)) + ((!g830) & (key[133]) & (g1914) & (!g4392) & (!g4393) & (!g5667)) + ((!g830) & (key[133]) & (g1914) & (!g4392) & (!g4393) & (g5667)) + ((!g830) & (key[133]) & (g1914) & (!g4392) & (g4393) & (!g5667)) + ((!g830) & (key[133]) & (g1914) & (!g4392) & (g4393) & (g5667)) + ((!g830) & (key[133]) & (g1914) & (g4392) & (!g4393) & (!g5667)) + ((!g830) & (key[133]) & (g1914) & (g4392) & (!g4393) & (g5667)) + ((!g830) & (key[133]) & (g1914) & (g4392) & (g4393) & (!g5667)) + ((!g830) & (key[133]) & (g1914) & (g4392) & (g4393) & (g5667)) + ((g830) & (!key[133]) & (!g1914) & (!g4392) & (!g4393) & (!g5667)) + ((g830) & (!key[133]) & (!g1914) & (!g4392) & (g4393) & (g5667)) + ((g830) & (!key[133]) & (!g1914) & (g4392) & (!g4393) & (!g5667)) + ((g830) & (!key[133]) & (!g1914) & (g4392) & (g4393) & (g5667)) + ((g830) & (!key[133]) & (g1914) & (!g4392) & (!g4393) & (!g5667)) + ((g830) & (!key[133]) & (g1914) & (!g4392) & (g4393) & (!g5667)) + ((g830) & (!key[133]) & (g1914) & (g4392) & (!g4393) & (g5667)) + ((g830) & (!key[133]) & (g1914) & (g4392) & (g4393) & (g5667)) + ((g830) & (key[133]) & (!g1914) & (!g4392) & (!g4393) & (!g5667)) + ((g830) & (key[133]) & (!g1914) & (!g4392) & (g4393) & (g5667)) + ((g830) & (key[133]) & (!g1914) & (g4392) & (!g4393) & (!g5667)) + ((g830) & (key[133]) & (!g1914) & (g4392) & (g4393) & (g5667)) + ((g830) & (key[133]) & (g1914) & (!g4392) & (!g4393) & (!g5667)) + ((g830) & (key[133]) & (g1914) & (!g4392) & (g4393) & (!g5667)) + ((g830) & (key[133]) & (g1914) & (g4392) & (!g4393) & (g5667)) + ((g830) & (key[133]) & (g1914) & (g4392) & (g4393) & (g5667)));
	assign g4395 = (((!g3050) & (!g4320) & (g3056)) + ((g3050) & (!g4320) & (!g3056)) + ((g3050) & (!g4320) & (g3056)) + ((g3050) & (g4320) & (g3056)));
	assign g4396 = (((!g2650) & (!g2684) & (g1778) & (g1814) & (!g4274)) + ((!g2650) & (g2684) & (!g1778) & (g1814) & (!g4274)) + ((!g2650) & (g2684) & (!g1778) & (g1814) & (g4274)) + ((!g2650) & (g2684) & (g1778) & (!g1814) & (!g4274)) + ((!g2650) & (g2684) & (g1778) & (g1814) & (!g4274)) + ((!g2650) & (g2684) & (g1778) & (g1814) & (g4274)) + ((g2650) & (!g2684) & (!g1778) & (g1814) & (!g4274)) + ((g2650) & (!g2684) & (g1778) & (g1814) & (!g4274)) + ((g2650) & (!g2684) & (g1778) & (g1814) & (g4274)) + ((g2650) & (g2684) & (!g1778) & (!g1814) & (!g4274)) + ((g2650) & (g2684) & (!g1778) & (g1814) & (!g4274)) + ((g2650) & (g2684) & (!g1778) & (g1814) & (g4274)) + ((g2650) & (g2684) & (g1778) & (!g1814) & (!g4274)) + ((g2650) & (g2684) & (g1778) & (!g1814) & (g4274)) + ((g2650) & (g2684) & (g1778) & (g1814) & (!g4274)) + ((g2650) & (g2684) & (g1778) & (g1814) & (g4274)));
	assign g4397 = (((!g830) & (key[101]) & (!g1914) & (!g4396) & (!g4395) & (!g5668)) + ((!g830) & (key[101]) & (!g1914) & (!g4396) & (!g4395) & (g5668)) + ((!g830) & (key[101]) & (!g1914) & (!g4396) & (g4395) & (!g5668)) + ((!g830) & (key[101]) & (!g1914) & (!g4396) & (g4395) & (g5668)) + ((!g830) & (key[101]) & (!g1914) & (g4396) & (!g4395) & (!g5668)) + ((!g830) & (key[101]) & (!g1914) & (g4396) & (!g4395) & (g5668)) + ((!g830) & (key[101]) & (!g1914) & (g4396) & (g4395) & (!g5668)) + ((!g830) & (key[101]) & (!g1914) & (g4396) & (g4395) & (g5668)) + ((!g830) & (key[101]) & (g1914) & (!g4396) & (!g4395) & (!g5668)) + ((!g830) & (key[101]) & (g1914) & (!g4396) & (!g4395) & (g5668)) + ((!g830) & (key[101]) & (g1914) & (!g4396) & (g4395) & (!g5668)) + ((!g830) & (key[101]) & (g1914) & (!g4396) & (g4395) & (g5668)) + ((!g830) & (key[101]) & (g1914) & (g4396) & (!g4395) & (!g5668)) + ((!g830) & (key[101]) & (g1914) & (g4396) & (!g4395) & (g5668)) + ((!g830) & (key[101]) & (g1914) & (g4396) & (g4395) & (!g5668)) + ((!g830) & (key[101]) & (g1914) & (g4396) & (g4395) & (g5668)) + ((g830) & (!key[101]) & (!g1914) & (!g4396) & (!g4395) & (!g5668)) + ((g830) & (!key[101]) & (!g1914) & (!g4396) & (g4395) & (!g5668)) + ((g830) & (!key[101]) & (!g1914) & (g4396) & (!g4395) & (g5668)) + ((g830) & (!key[101]) & (!g1914) & (g4396) & (g4395) & (g5668)) + ((g830) & (!key[101]) & (g1914) & (!g4396) & (!g4395) & (!g5668)) + ((g830) & (!key[101]) & (g1914) & (!g4396) & (g4395) & (g5668)) + ((g830) & (!key[101]) & (g1914) & (g4396) & (!g4395) & (!g5668)) + ((g830) & (!key[101]) & (g1914) & (g4396) & (g4395) & (g5668)) + ((g830) & (key[101]) & (!g1914) & (!g4396) & (!g4395) & (!g5668)) + ((g830) & (key[101]) & (!g1914) & (!g4396) & (g4395) & (!g5668)) + ((g830) & (key[101]) & (!g1914) & (g4396) & (!g4395) & (g5668)) + ((g830) & (key[101]) & (!g1914) & (g4396) & (g4395) & (g5668)) + ((g830) & (key[101]) & (g1914) & (!g4396) & (!g4395) & (!g5668)) + ((g830) & (key[101]) & (g1914) & (!g4396) & (g4395) & (g5668)) + ((g830) & (key[101]) & (g1914) & (g4396) & (!g4395) & (!g5668)) + ((g830) & (key[101]) & (g1914) & (g4396) & (g4395) & (g5668)));
	assign g4398 = (((!g3260) & (!g4277) & (!g3222) & (g3301) & (g3305)) + ((!g3260) & (!g4277) & (g3222) & (!g3301) & (g3305)) + ((!g3260) & (!g4277) & (g3222) & (g3301) & (!g3305)) + ((!g3260) & (!g4277) & (g3222) & (g3301) & (g3305)) + ((!g3260) & (g4277) & (!g3222) & (g3301) & (g3305)) + ((!g3260) & (g4277) & (g3222) & (g3301) & (g3305)) + ((g3260) & (!g4277) & (!g3222) & (!g3301) & (g3305)) + ((g3260) & (!g4277) & (!g3222) & (g3301) & (!g3305)) + ((g3260) & (!g4277) & (!g3222) & (g3301) & (g3305)) + ((g3260) & (!g4277) & (g3222) & (!g3301) & (g3305)) + ((g3260) & (!g4277) & (g3222) & (g3301) & (!g3305)) + ((g3260) & (!g4277) & (g3222) & (g3301) & (g3305)) + ((g3260) & (g4277) & (!g3222) & (g3301) & (g3305)) + ((g3260) & (g4277) & (g3222) & (!g3301) & (g3305)) + ((g3260) & (g4277) & (g3222) & (g3301) & (!g3305)) + ((g3260) & (g4277) & (g3222) & (g3301) & (g3305)));
	assign g4399 = (((!g2376) & (g3061) & (!g4328)) + ((g2376) & (!g3061) & (!g4328)) + ((g2376) & (g3061) & (!g4328)) + ((g2376) & (g3061) & (g4328)));
	assign g4400 = (((!g830) & (nonce[5]) & (!g1914) & (!g4398) & (!g4399) & (!g5669)) + ((!g830) & (nonce[5]) & (!g1914) & (!g4398) & (!g4399) & (g5669)) + ((!g830) & (nonce[5]) & (!g1914) & (!g4398) & (g4399) & (!g5669)) + ((!g830) & (nonce[5]) & (!g1914) & (!g4398) & (g4399) & (g5669)) + ((!g830) & (nonce[5]) & (!g1914) & (g4398) & (!g4399) & (!g5669)) + ((!g830) & (nonce[5]) & (!g1914) & (g4398) & (!g4399) & (g5669)) + ((!g830) & (nonce[5]) & (!g1914) & (g4398) & (g4399) & (!g5669)) + ((!g830) & (nonce[5]) & (!g1914) & (g4398) & (g4399) & (g5669)) + ((!g830) & (nonce[5]) & (g1914) & (!g4398) & (!g4399) & (!g5669)) + ((!g830) & (nonce[5]) & (g1914) & (!g4398) & (!g4399) & (g5669)) + ((!g830) & (nonce[5]) & (g1914) & (!g4398) & (g4399) & (!g5669)) + ((!g830) & (nonce[5]) & (g1914) & (!g4398) & (g4399) & (g5669)) + ((!g830) & (nonce[5]) & (g1914) & (g4398) & (!g4399) & (!g5669)) + ((!g830) & (nonce[5]) & (g1914) & (g4398) & (!g4399) & (g5669)) + ((!g830) & (nonce[5]) & (g1914) & (g4398) & (g4399) & (!g5669)) + ((!g830) & (nonce[5]) & (g1914) & (g4398) & (g4399) & (g5669)) + ((g830) & (!nonce[5]) & (!g1914) & (!g4398) & (!g4399) & (!g5669)) + ((g830) & (!nonce[5]) & (!g1914) & (!g4398) & (g4399) & (g5669)) + ((g830) & (!nonce[5]) & (!g1914) & (g4398) & (!g4399) & (!g5669)) + ((g830) & (!nonce[5]) & (!g1914) & (g4398) & (g4399) & (g5669)) + ((g830) & (!nonce[5]) & (g1914) & (!g4398) & (!g4399) & (!g5669)) + ((g830) & (!nonce[5]) & (g1914) & (!g4398) & (g4399) & (!g5669)) + ((g830) & (!nonce[5]) & (g1914) & (g4398) & (!g4399) & (g5669)) + ((g830) & (!nonce[5]) & (g1914) & (g4398) & (g4399) & (g5669)) + ((g830) & (nonce[5]) & (!g1914) & (!g4398) & (!g4399) & (!g5669)) + ((g830) & (nonce[5]) & (!g1914) & (!g4398) & (g4399) & (g5669)) + ((g830) & (nonce[5]) & (!g1914) & (g4398) & (!g4399) & (!g5669)) + ((g830) & (nonce[5]) & (!g1914) & (g4398) & (g4399) & (g5669)) + ((g830) & (nonce[5]) & (g1914) & (!g4398) & (!g4399) & (!g5669)) + ((g830) & (nonce[5]) & (g1914) & (!g4398) & (g4399) & (!g5669)) + ((g830) & (nonce[5]) & (g1914) & (g4398) & (!g4399) & (g5669)) + ((g830) & (nonce[5]) & (g1914) & (g4398) & (g4399) & (g5669)));
	assign g4401 = (((!g2797) & (g2830) & (g4344)) + ((g2797) & (!g2830) & (g4344)) + ((g2797) & (g2830) & (!g4344)) + ((g2797) & (g2830) & (g4344)));
	assign g4402 = (((!g2813) & (!g2838) & (!g2822) & (g2871) & (!g4345)) + ((!g2813) & (!g2838) & (!g2822) & (g2871) & (g4345)) + ((!g2813) & (!g2838) & (g2822) & (!g2871) & (g4345)) + ((!g2813) & (!g2838) & (g2822) & (g2871) & (!g4345)) + ((!g2813) & (g2838) & (!g2822) & (!g2871) & (!g4345)) + ((!g2813) & (g2838) & (!g2822) & (!g2871) & (g4345)) + ((!g2813) & (g2838) & (g2822) & (!g2871) & (!g4345)) + ((!g2813) & (g2838) & (g2822) & (g2871) & (g4345)) + ((g2813) & (!g2838) & (!g2822) & (!g2871) & (g4345)) + ((g2813) & (!g2838) & (!g2822) & (g2871) & (!g4345)) + ((g2813) & (!g2838) & (g2822) & (!g2871) & (!g4345)) + ((g2813) & (!g2838) & (g2822) & (!g2871) & (g4345)) + ((g2813) & (g2838) & (!g2822) & (!g2871) & (!g4345)) + ((g2813) & (g2838) & (!g2822) & (g2871) & (g4345)) + ((g2813) & (g2838) & (g2822) & (g2871) & (!g4345)) + ((g2813) & (g2838) & (g2822) & (g2871) & (g4345)));
	assign g4403 = (((!g3163) & (!g3155) & (!g3199) & (!g3196) & (!g4284) & (!g4285)) + ((!g3163) & (!g3155) & (!g3199) & (!g3196) & (!g4284) & (g4285)) + ((!g3163) & (!g3155) & (!g3199) & (!g3196) & (g4284) & (!g4285)) + ((!g3163) & (!g3155) & (!g3199) & (!g3196) & (g4284) & (g4285)) + ((!g3163) & (!g3155) & (!g3199) & (g3196) & (!g4284) & (!g4285)) + ((!g3163) & (!g3155) & (!g3199) & (g3196) & (!g4284) & (g4285)) + ((!g3163) & (!g3155) & (!g3199) & (g3196) & (g4284) & (!g4285)) + ((!g3163) & (!g3155) & (!g3199) & (g3196) & (g4284) & (g4285)) + ((!g3163) & (!g3155) & (g3199) & (!g3196) & (!g4284) & (!g4285)) + ((!g3163) & (!g3155) & (g3199) & (!g3196) & (!g4284) & (g4285)) + ((!g3163) & (!g3155) & (g3199) & (!g3196) & (g4284) & (!g4285)) + ((!g3163) & (!g3155) & (g3199) & (!g3196) & (g4284) & (g4285)) + ((!g3163) & (g3155) & (!g3199) & (!g3196) & (!g4284) & (!g4285)) + ((!g3163) & (g3155) & (!g3199) & (!g3196) & (!g4284) & (g4285)) + ((!g3163) & (g3155) & (!g3199) & (!g3196) & (g4284) & (!g4285)) + ((!g3163) & (g3155) & (!g3199) & (!g3196) & (g4284) & (g4285)) + ((!g3163) & (g3155) & (!g3199) & (g3196) & (!g4284) & (!g4285)) + ((!g3163) & (g3155) & (g3199) & (!g3196) & (!g4284) & (!g4285)) + ((g3163) & (!g3155) & (!g3199) & (!g3196) & (!g4284) & (!g4285)) + ((g3163) & (!g3155) & (!g3199) & (!g3196) & (!g4284) & (g4285)) + ((g3163) & (!g3155) & (!g3199) & (!g3196) & (g4284) & (!g4285)) + ((g3163) & (!g3155) & (!g3199) & (!g3196) & (g4284) & (g4285)) + ((g3163) & (!g3155) & (!g3199) & (g3196) & (!g4284) & (!g4285)) + ((g3163) & (!g3155) & (g3199) & (!g3196) & (!g4284) & (!g4285)) + ((g3163) & (g3155) & (!g3199) & (!g3196) & (!g4284) & (!g4285)) + ((g3163) & (g3155) & (!g3199) & (!g3196) & (!g4284) & (g4285)) + ((g3163) & (g3155) & (!g3199) & (!g3196) & (g4284) & (!g4285)) + ((g3163) & (g3155) & (!g3199) & (!g3196) & (g4284) & (g4285)));
	assign g4404 = (((g1914) & (!g3260) & (!g3240) & (!g4403)) + ((g1914) & (!g3260) & (g3240) & (g4403)) + ((g1914) & (g3260) & (!g3240) & (g4403)) + ((g1914) & (g3260) & (g3240) & (!g4403)));
	assign g4405 = (((!g2552) & (!g2599) & (!g3172) & (!g3213) & (!g4288) & (!g4289)) + ((!g2552) & (!g2599) & (!g3172) & (!g3213) & (!g4288) & (g4289)) + ((!g2552) & (!g2599) & (!g3172) & (!g3213) & (g4288) & (!g4289)) + ((!g2552) & (!g2599) & (!g3172) & (!g3213) & (g4288) & (g4289)) + ((!g2552) & (!g2599) & (!g3172) & (g3213) & (!g4288) & (!g4289)) + ((!g2552) & (!g2599) & (!g3172) & (g3213) & (!g4288) & (g4289)) + ((!g2552) & (!g2599) & (!g3172) & (g3213) & (g4288) & (!g4289)) + ((!g2552) & (!g2599) & (!g3172) & (g3213) & (g4288) & (g4289)) + ((!g2552) & (!g2599) & (g3172) & (!g3213) & (!g4288) & (!g4289)) + ((!g2552) & (!g2599) & (g3172) & (!g3213) & (!g4288) & (g4289)) + ((!g2552) & (!g2599) & (g3172) & (!g3213) & (g4288) & (!g4289)) + ((!g2552) & (!g2599) & (g3172) & (!g3213) & (g4288) & (g4289)) + ((!g2552) & (!g2599) & (g3172) & (g3213) & (!g4288) & (!g4289)) + ((!g2552) & (g2599) & (!g3172) & (!g3213) & (!g4288) & (!g4289)) + ((!g2552) & (g2599) & (!g3172) & (!g3213) & (!g4288) & (g4289)) + ((!g2552) & (g2599) & (!g3172) & (!g3213) & (g4288) & (!g4289)) + ((!g2552) & (g2599) & (!g3172) & (!g3213) & (g4288) & (g4289)) + ((!g2552) & (g2599) & (g3172) & (!g3213) & (!g4288) & (!g4289)) + ((g2552) & (!g2599) & (!g3172) & (!g3213) & (!g4288) & (!g4289)) + ((g2552) & (!g2599) & (!g3172) & (!g3213) & (!g4288) & (g4289)) + ((g2552) & (!g2599) & (!g3172) & (!g3213) & (g4288) & (!g4289)) + ((g2552) & (!g2599) & (!g3172) & (!g3213) & (g4288) & (g4289)) + ((g2552) & (!g2599) & (!g3172) & (g3213) & (!g4288) & (!g4289)) + ((g2552) & (!g2599) & (g3172) & (!g3213) & (!g4288) & (!g4289)) + ((g2552) & (!g2599) & (g3172) & (!g3213) & (!g4288) & (g4289)) + ((g2552) & (!g2599) & (g3172) & (!g3213) & (g4288) & (!g4289)) + ((g2552) & (!g2599) & (g3172) & (!g3213) & (g4288) & (g4289)) + ((g2552) & (g2599) & (!g3172) & (!g3213) & (!g4288) & (!g4289)));
	assign g4406 = (((!g1914) & (!g2648) & (!g3284) & (!g4405)) + ((!g1914) & (!g2648) & (g3284) & (g4405)) + ((!g1914) & (g2648) & (!g3284) & (g4405)) + ((!g1914) & (g2648) & (g3284) & (!g4405)));
	assign g4407 = (((!g830) & (!g2200) & (!g4404) & (!g4406) & (nonce[37])) + ((!g830) & (!g2200) & (!g4404) & (g4406) & (nonce[37])) + ((!g830) & (!g2200) & (g4404) & (!g4406) & (nonce[37])) + ((!g830) & (!g2200) & (g4404) & (g4406) & (nonce[37])) + ((!g830) & (g2200) & (!g4404) & (!g4406) & (nonce[37])) + ((!g830) & (g2200) & (!g4404) & (g4406) & (nonce[37])) + ((!g830) & (g2200) & (g4404) & (!g4406) & (nonce[37])) + ((!g830) & (g2200) & (g4404) & (g4406) & (nonce[37])) + ((g830) & (!g2200) & (!g4404) & (g4406) & (!nonce[37])) + ((g830) & (!g2200) & (!g4404) & (g4406) & (nonce[37])) + ((g830) & (!g2200) & (g4404) & (!g4406) & (!nonce[37])) + ((g830) & (!g2200) & (g4404) & (!g4406) & (nonce[37])) + ((g830) & (!g2200) & (g4404) & (g4406) & (!nonce[37])) + ((g830) & (!g2200) & (g4404) & (g4406) & (nonce[37])) + ((g830) & (g2200) & (!g4404) & (!g4406) & (!nonce[37])) + ((g830) & (g2200) & (!g4404) & (!g4406) & (nonce[37])));
	assign g4408 = (((!g2379) & (!g4331) & (g3064)) + ((g2379) & (!g4331) & (!g3064)) + ((g2379) & (!g4331) & (g3064)) + ((g2379) & (g4331) & (g3064)));
	assign g4409 = (((!g3235) & (!g4293) & (!g3240) & (g3295) & (g3303)) + ((!g3235) & (!g4293) & (g3240) & (!g3295) & (g3303)) + ((!g3235) & (!g4293) & (g3240) & (g3295) & (!g3303)) + ((!g3235) & (!g4293) & (g3240) & (g3295) & (g3303)) + ((!g3235) & (g4293) & (!g3240) & (g3295) & (g3303)) + ((!g3235) & (g4293) & (g3240) & (g3295) & (g3303)) + ((g3235) & (!g4293) & (!g3240) & (!g3295) & (g3303)) + ((g3235) & (!g4293) & (!g3240) & (g3295) & (!g3303)) + ((g3235) & (!g4293) & (!g3240) & (g3295) & (g3303)) + ((g3235) & (!g4293) & (g3240) & (!g3295) & (g3303)) + ((g3235) & (!g4293) & (g3240) & (g3295) & (!g3303)) + ((g3235) & (!g4293) & (g3240) & (g3295) & (g3303)) + ((g3235) & (g4293) & (!g3240) & (g3295) & (g3303)) + ((g3235) & (g4293) & (g3240) & (!g3295) & (g3303)) + ((g3235) & (g4293) & (g3240) & (g3295) & (!g3303)) + ((g3235) & (g4293) & (g3240) & (g3295) & (g3303)));
	assign g4410 = (((!g830) & (key[229]) & (!g1914) & (!g4409) & (!g4408) & (!g5671)) + ((!g830) & (key[229]) & (!g1914) & (!g4409) & (!g4408) & (g5671)) + ((!g830) & (key[229]) & (!g1914) & (!g4409) & (g4408) & (!g5671)) + ((!g830) & (key[229]) & (!g1914) & (!g4409) & (g4408) & (g5671)) + ((!g830) & (key[229]) & (!g1914) & (g4409) & (!g4408) & (!g5671)) + ((!g830) & (key[229]) & (!g1914) & (g4409) & (!g4408) & (g5671)) + ((!g830) & (key[229]) & (!g1914) & (g4409) & (g4408) & (!g5671)) + ((!g830) & (key[229]) & (!g1914) & (g4409) & (g4408) & (g5671)) + ((!g830) & (key[229]) & (g1914) & (!g4409) & (!g4408) & (!g5671)) + ((!g830) & (key[229]) & (g1914) & (!g4409) & (!g4408) & (g5671)) + ((!g830) & (key[229]) & (g1914) & (!g4409) & (g4408) & (!g5671)) + ((!g830) & (key[229]) & (g1914) & (!g4409) & (g4408) & (g5671)) + ((!g830) & (key[229]) & (g1914) & (g4409) & (!g4408) & (!g5671)) + ((!g830) & (key[229]) & (g1914) & (g4409) & (!g4408) & (g5671)) + ((!g830) & (key[229]) & (g1914) & (g4409) & (g4408) & (!g5671)) + ((!g830) & (key[229]) & (g1914) & (g4409) & (g4408) & (g5671)) + ((g830) & (!key[229]) & (!g1914) & (!g4409) & (!g4408) & (!g5671)) + ((g830) & (!key[229]) & (!g1914) & (!g4409) & (g4408) & (!g5671)) + ((g830) & (!key[229]) & (!g1914) & (g4409) & (!g4408) & (g5671)) + ((g830) & (!key[229]) & (!g1914) & (g4409) & (g4408) & (g5671)) + ((g830) & (!key[229]) & (g1914) & (!g4409) & (!g4408) & (!g5671)) + ((g830) & (!key[229]) & (g1914) & (!g4409) & (g4408) & (g5671)) + ((g830) & (!key[229]) & (g1914) & (g4409) & (!g4408) & (!g5671)) + ((g830) & (!key[229]) & (g1914) & (g4409) & (g4408) & (g5671)) + ((g830) & (key[229]) & (!g1914) & (!g4409) & (!g4408) & (!g5671)) + ((g830) & (key[229]) & (!g1914) & (!g4409) & (g4408) & (!g5671)) + ((g830) & (key[229]) & (!g1914) & (g4409) & (!g4408) & (g5671)) + ((g830) & (key[229]) & (!g1914) & (g4409) & (g4408) & (g5671)) + ((g830) & (key[229]) & (g1914) & (!g4409) & (!g4408) & (!g5671)) + ((g830) & (key[229]) & (g1914) & (!g4409) & (g4408) & (g5671)) + ((g830) & (key[229]) & (g1914) & (g4409) & (!g4408) & (!g5671)) + ((g830) & (key[229]) & (g1914) & (g4409) & (g4408) & (g5671)));
	assign g4411 = (((!g2556) & (!g2602) & (!g3172) & (!g3213) & (!g4297) & (!g4298)) + ((!g2556) & (!g2602) & (!g3172) & (!g3213) & (!g4297) & (g4298)) + ((!g2556) & (!g2602) & (!g3172) & (!g3213) & (g4297) & (!g4298)) + ((!g2556) & (!g2602) & (!g3172) & (!g3213) & (g4297) & (g4298)) + ((!g2556) & (!g2602) & (!g3172) & (g3213) & (!g4297) & (!g4298)) + ((!g2556) & (!g2602) & (!g3172) & (g3213) & (!g4297) & (g4298)) + ((!g2556) & (!g2602) & (!g3172) & (g3213) & (g4297) & (!g4298)) + ((!g2556) & (!g2602) & (!g3172) & (g3213) & (g4297) & (g4298)) + ((!g2556) & (!g2602) & (g3172) & (!g3213) & (!g4297) & (!g4298)) + ((!g2556) & (!g2602) & (g3172) & (!g3213) & (!g4297) & (g4298)) + ((!g2556) & (!g2602) & (g3172) & (!g3213) & (g4297) & (!g4298)) + ((!g2556) & (!g2602) & (g3172) & (!g3213) & (g4297) & (g4298)) + ((!g2556) & (!g2602) & (g3172) & (g3213) & (!g4297) & (!g4298)) + ((!g2556) & (g2602) & (!g3172) & (!g3213) & (!g4297) & (!g4298)) + ((!g2556) & (g2602) & (!g3172) & (!g3213) & (!g4297) & (g4298)) + ((!g2556) & (g2602) & (!g3172) & (!g3213) & (g4297) & (!g4298)) + ((!g2556) & (g2602) & (!g3172) & (!g3213) & (g4297) & (g4298)) + ((!g2556) & (g2602) & (g3172) & (!g3213) & (!g4297) & (!g4298)) + ((g2556) & (!g2602) & (!g3172) & (!g3213) & (!g4297) & (!g4298)) + ((g2556) & (!g2602) & (!g3172) & (!g3213) & (!g4297) & (g4298)) + ((g2556) & (!g2602) & (!g3172) & (!g3213) & (g4297) & (!g4298)) + ((g2556) & (!g2602) & (!g3172) & (!g3213) & (g4297) & (g4298)) + ((g2556) & (!g2602) & (!g3172) & (g3213) & (!g4297) & (!g4298)) + ((g2556) & (!g2602) & (g3172) & (!g3213) & (!g4297) & (!g4298)) + ((g2556) & (!g2602) & (g3172) & (!g3213) & (!g4297) & (g4298)) + ((g2556) & (!g2602) & (g3172) & (!g3213) & (g4297) & (!g4298)) + ((g2556) & (!g2602) & (g3172) & (!g3213) & (g4297) & (g4298)) + ((g2556) & (g2602) & (!g3172) & (!g3213) & (!g4297) & (!g4298)));
	assign g4412 = (((g1914) & (!g2650) & (!g3284) & (!g4411)) + ((g1914) & (!g2650) & (g3284) & (g4411)) + ((g1914) & (g2650) & (!g3284) & (g4411)) + ((g1914) & (g2650) & (g3284) & (!g4411)));
	assign g4413 = (((!g3163) & (!g3161) & (!g3199) & (!g3187) & (!g4301) & (!g4302)) + ((!g3163) & (!g3161) & (!g3199) & (!g3187) & (!g4301) & (g4302)) + ((!g3163) & (!g3161) & (!g3199) & (!g3187) & (g4301) & (!g4302)) + ((!g3163) & (!g3161) & (!g3199) & (!g3187) & (g4301) & (g4302)) + ((!g3163) & (!g3161) & (!g3199) & (g3187) & (!g4301) & (!g4302)) + ((!g3163) & (!g3161) & (!g3199) & (g3187) & (!g4301) & (g4302)) + ((!g3163) & (!g3161) & (!g3199) & (g3187) & (g4301) & (!g4302)) + ((!g3163) & (!g3161) & (!g3199) & (g3187) & (g4301) & (g4302)) + ((!g3163) & (!g3161) & (g3199) & (!g3187) & (!g4301) & (!g4302)) + ((!g3163) & (!g3161) & (g3199) & (!g3187) & (!g4301) & (g4302)) + ((!g3163) & (!g3161) & (g3199) & (!g3187) & (g4301) & (!g4302)) + ((!g3163) & (!g3161) & (g3199) & (!g3187) & (g4301) & (g4302)) + ((!g3163) & (g3161) & (!g3199) & (!g3187) & (!g4301) & (!g4302)) + ((!g3163) & (g3161) & (!g3199) & (!g3187) & (!g4301) & (g4302)) + ((!g3163) & (g3161) & (!g3199) & (!g3187) & (g4301) & (!g4302)) + ((!g3163) & (g3161) & (!g3199) & (!g3187) & (g4301) & (g4302)) + ((!g3163) & (g3161) & (!g3199) & (g3187) & (!g4301) & (!g4302)) + ((!g3163) & (g3161) & (g3199) & (!g3187) & (!g4301) & (!g4302)) + ((g3163) & (!g3161) & (!g3199) & (!g3187) & (!g4301) & (!g4302)) + ((g3163) & (!g3161) & (!g3199) & (!g3187) & (!g4301) & (g4302)) + ((g3163) & (!g3161) & (!g3199) & (!g3187) & (g4301) & (!g4302)) + ((g3163) & (!g3161) & (!g3199) & (!g3187) & (g4301) & (g4302)) + ((g3163) & (!g3161) & (!g3199) & (g3187) & (!g4301) & (!g4302)) + ((g3163) & (!g3161) & (g3199) & (!g3187) & (!g4301) & (!g4302)) + ((g3163) & (g3161) & (!g3199) & (!g3187) & (!g4301) & (!g4302)) + ((g3163) & (g3161) & (!g3199) & (!g3187) & (!g4301) & (g4302)) + ((g3163) & (g3161) & (!g3199) & (!g3187) & (g4301) & (!g4302)) + ((g3163) & (g3161) & (!g3199) & (!g3187) & (g4301) & (g4302)));
	assign g4414 = (((!g1914) & (!g3260) & (!g3255) & (!g4413)) + ((!g1914) & (!g3260) & (g3255) & (g4413)) + ((!g1914) & (g3260) & (!g3255) & (g4413)) + ((!g1914) & (g3260) & (g3255) & (!g4413)));
	assign g4415 = (((!g830) & (!g2205) & (!g4412) & (!g4414) & (key[197])) + ((!g830) & (!g2205) & (!g4412) & (g4414) & (key[197])) + ((!g830) & (!g2205) & (g4412) & (!g4414) & (key[197])) + ((!g830) & (!g2205) & (g4412) & (g4414) & (key[197])) + ((!g830) & (g2205) & (!g4412) & (!g4414) & (key[197])) + ((!g830) & (g2205) & (!g4412) & (g4414) & (key[197])) + ((!g830) & (g2205) & (g4412) & (!g4414) & (key[197])) + ((!g830) & (g2205) & (g4412) & (g4414) & (key[197])) + ((g830) & (!g2205) & (!g4412) & (g4414) & (!key[197])) + ((g830) & (!g2205) & (!g4412) & (g4414) & (key[197])) + ((g830) & (!g2205) & (g4412) & (!g4414) & (!key[197])) + ((g830) & (!g2205) & (g4412) & (!g4414) & (key[197])) + ((g830) & (!g2205) & (g4412) & (g4414) & (!key[197])) + ((g830) & (!g2205) & (g4412) & (g4414) & (key[197])) + ((g830) & (g2205) & (!g4412) & (!g4414) & (!key[197])) + ((g830) & (g2205) & (!g4412) & (!g4414) & (key[197])));
	assign g4416 = (((!g2810) & (g2822) & (g4361)) + ((g2810) & (!g2822) & (g4361)) + ((g2810) & (g2822) & (!g4361)) + ((g2810) & (g2822) & (g4361)));
	assign g4417 = (((!g2827) & (!g2851) & (!g2830) & (g2863) & (!g4362)) + ((!g2827) & (!g2851) & (!g2830) & (g2863) & (g4362)) + ((!g2827) & (!g2851) & (g2830) & (!g2863) & (g4362)) + ((!g2827) & (!g2851) & (g2830) & (g2863) & (!g4362)) + ((!g2827) & (g2851) & (!g2830) & (!g2863) & (!g4362)) + ((!g2827) & (g2851) & (!g2830) & (!g2863) & (g4362)) + ((!g2827) & (g2851) & (g2830) & (!g2863) & (!g4362)) + ((!g2827) & (g2851) & (g2830) & (g2863) & (g4362)) + ((g2827) & (!g2851) & (!g2830) & (!g2863) & (g4362)) + ((g2827) & (!g2851) & (!g2830) & (g2863) & (!g4362)) + ((g2827) & (!g2851) & (g2830) & (!g2863) & (!g4362)) + ((g2827) & (!g2851) & (g2830) & (!g2863) & (g4362)) + ((g2827) & (g2851) & (!g2830) & (!g2863) & (!g4362)) + ((g2827) & (g2851) & (!g2830) & (g2863) & (g4362)) + ((g2827) & (g2851) & (g2830) & (g2863) & (!g4362)) + ((g2827) & (g2851) & (g2830) & (g2863) & (g4362)));
	assign g4418 = (((!g1132) & (!g1165) & (!g4364) & (!g2350) & (g2399)) + ((!g1132) & (!g1165) & (!g4364) & (g2350) & (g2399)) + ((!g1132) & (!g1165) & (g4364) & (!g2350) & (g2399)) + ((!g1132) & (!g1165) & (g4364) & (g2350) & (!g2399)) + ((!g1132) & (g1165) & (!g4364) & (!g2350) & (!g2399)) + ((!g1132) & (g1165) & (!g4364) & (g2350) & (!g2399)) + ((!g1132) & (g1165) & (g4364) & (!g2350) & (!g2399)) + ((!g1132) & (g1165) & (g4364) & (g2350) & (g2399)) + ((g1132) & (!g1165) & (!g4364) & (!g2350) & (g2399)) + ((g1132) & (!g1165) & (!g4364) & (g2350) & (!g2399)) + ((g1132) & (!g1165) & (g4364) & (!g2350) & (!g2399)) + ((g1132) & (!g1165) & (g4364) & (g2350) & (!g2399)) + ((g1132) & (g1165) & (!g4364) & (!g2350) & (!g2399)) + ((g1132) & (g1165) & (!g4364) & (g2350) & (g2399)) + ((g1132) & (g1165) & (g4364) & (!g2350) & (g2399)) + ((g1132) & (g1165) & (g4364) & (g2350) & (g2399)));
	assign g4419 = (((!g2354) & (!g2390) & (!g2369) & (g2396) & (!g4366)) + ((!g2354) & (!g2390) & (!g2369) & (g2396) & (g4366)) + ((!g2354) & (!g2390) & (g2369) & (!g2396) & (g4366)) + ((!g2354) & (!g2390) & (g2369) & (g2396) & (!g4366)) + ((!g2354) & (g2390) & (!g2369) & (!g2396) & (!g4366)) + ((!g2354) & (g2390) & (!g2369) & (!g2396) & (g4366)) + ((!g2354) & (g2390) & (g2369) & (!g2396) & (!g4366)) + ((!g2354) & (g2390) & (g2369) & (g2396) & (g4366)) + ((g2354) & (!g2390) & (!g2369) & (!g2396) & (g4366)) + ((g2354) & (!g2390) & (!g2369) & (g2396) & (!g4366)) + ((g2354) & (!g2390) & (g2369) & (!g2396) & (!g4366)) + ((g2354) & (!g2390) & (g2369) & (!g2396) & (g4366)) + ((g2354) & (g2390) & (!g2369) & (!g2396) & (!g4366)) + ((g2354) & (g2390) & (!g2369) & (g2396) & (g4366)) + ((g2354) & (g2390) & (g2369) & (g2396) & (!g4366)) + ((g2354) & (g2390) & (g2369) & (g2396) & (g4366)));
	assign g4420 = (((!g830) & (!g1914) & (!g2210) & (!g4418) & (!g4419) & (key[51])) + ((!g830) & (!g1914) & (!g2210) & (!g4418) & (g4419) & (key[51])) + ((!g830) & (!g1914) & (!g2210) & (g4418) & (!g4419) & (key[51])) + ((!g830) & (!g1914) & (!g2210) & (g4418) & (g4419) & (key[51])) + ((!g830) & (!g1914) & (g2210) & (!g4418) & (!g4419) & (key[51])) + ((!g830) & (!g1914) & (g2210) & (!g4418) & (g4419) & (key[51])) + ((!g830) & (!g1914) & (g2210) & (g4418) & (!g4419) & (key[51])) + ((!g830) & (!g1914) & (g2210) & (g4418) & (g4419) & (key[51])) + ((!g830) & (g1914) & (!g2210) & (!g4418) & (!g4419) & (key[51])) + ((!g830) & (g1914) & (!g2210) & (!g4418) & (g4419) & (key[51])) + ((!g830) & (g1914) & (!g2210) & (g4418) & (!g4419) & (key[51])) + ((!g830) & (g1914) & (!g2210) & (g4418) & (g4419) & (key[51])) + ((!g830) & (g1914) & (g2210) & (!g4418) & (!g4419) & (key[51])) + ((!g830) & (g1914) & (g2210) & (!g4418) & (g4419) & (key[51])) + ((!g830) & (g1914) & (g2210) & (g4418) & (!g4419) & (key[51])) + ((!g830) & (g1914) & (g2210) & (g4418) & (g4419) & (key[51])) + ((g830) & (!g1914) & (!g2210) & (!g4418) & (g4419) & (!key[51])) + ((g830) & (!g1914) & (!g2210) & (!g4418) & (g4419) & (key[51])) + ((g830) & (!g1914) & (!g2210) & (g4418) & (g4419) & (!key[51])) + ((g830) & (!g1914) & (!g2210) & (g4418) & (g4419) & (key[51])) + ((g830) & (!g1914) & (g2210) & (!g4418) & (!g4419) & (!key[51])) + ((g830) & (!g1914) & (g2210) & (!g4418) & (!g4419) & (key[51])) + ((g830) & (!g1914) & (g2210) & (g4418) & (!g4419) & (!key[51])) + ((g830) & (!g1914) & (g2210) & (g4418) & (!g4419) & (key[51])) + ((g830) & (g1914) & (!g2210) & (g4418) & (!g4419) & (!key[51])) + ((g830) & (g1914) & (!g2210) & (g4418) & (!g4419) & (key[51])) + ((g830) & (g1914) & (!g2210) & (g4418) & (g4419) & (!key[51])) + ((g830) & (g1914) & (!g2210) & (g4418) & (g4419) & (key[51])) + ((g830) & (g1914) & (g2210) & (!g4418) & (!g4419) & (!key[51])) + ((g830) & (g1914) & (g2210) & (!g4418) & (!g4419) & (key[51])) + ((g830) & (g1914) & (g2210) & (!g4418) & (g4419) & (!key[51])) + ((g830) & (g1914) & (g2210) & (!g4418) & (g4419) & (key[51])));
	assign g4421 = (((!g3747) & (!g3748)));
	assign g4422 = (((!g1953) & (!g2233) & (!g4421)) + ((!g1953) & (g2233) & (g4421)) + ((g1953) & (!g2233) & (g4421)) + ((g1953) & (g2233) & (!g4421)));
	assign g4423 = (((!g2462) & (!g2542) & (!g2509) & (g2546) & (!g4369)) + ((!g2462) & (!g2542) & (!g2509) & (g2546) & (g4369)) + ((!g2462) & (!g2542) & (g2509) & (!g2546) & (!g4369)) + ((!g2462) & (!g2542) & (g2509) & (g2546) & (g4369)) + ((!g2462) & (g2542) & (!g2509) & (!g2546) & (!g4369)) + ((!g2462) & (g2542) & (!g2509) & (!g2546) & (g4369)) + ((!g2462) & (g2542) & (g2509) & (!g2546) & (g4369)) + ((!g2462) & (g2542) & (g2509) & (g2546) & (!g4369)) + ((g2462) & (!g2542) & (!g2509) & (!g2546) & (!g4369)) + ((g2462) & (!g2542) & (!g2509) & (g2546) & (g4369)) + ((g2462) & (!g2542) & (g2509) & (!g2546) & (!g4369)) + ((g2462) & (!g2542) & (g2509) & (!g2546) & (g4369)) + ((g2462) & (g2542) & (!g2509) & (!g2546) & (g4369)) + ((g2462) & (g2542) & (!g2509) & (g2546) & (!g4369)) + ((g2462) & (g2542) & (g2509) & (g2546) & (!g4369)) + ((g2462) & (g2542) & (g2509) & (g2546) & (g4369)));
	assign g4424 = (((!g830) & (!g1914) & (!g2211) & (!g4422) & (!g4423) & (key[83])) + ((!g830) & (!g1914) & (!g2211) & (!g4422) & (g4423) & (key[83])) + ((!g830) & (!g1914) & (!g2211) & (g4422) & (!g4423) & (key[83])) + ((!g830) & (!g1914) & (!g2211) & (g4422) & (g4423) & (key[83])) + ((!g830) & (!g1914) & (g2211) & (!g4422) & (!g4423) & (key[83])) + ((!g830) & (!g1914) & (g2211) & (!g4422) & (g4423) & (key[83])) + ((!g830) & (!g1914) & (g2211) & (g4422) & (!g4423) & (key[83])) + ((!g830) & (!g1914) & (g2211) & (g4422) & (g4423) & (key[83])) + ((!g830) & (g1914) & (!g2211) & (!g4422) & (!g4423) & (key[83])) + ((!g830) & (g1914) & (!g2211) & (!g4422) & (g4423) & (key[83])) + ((!g830) & (g1914) & (!g2211) & (g4422) & (!g4423) & (key[83])) + ((!g830) & (g1914) & (!g2211) & (g4422) & (g4423) & (key[83])) + ((!g830) & (g1914) & (g2211) & (!g4422) & (!g4423) & (key[83])) + ((!g830) & (g1914) & (g2211) & (!g4422) & (g4423) & (key[83])) + ((!g830) & (g1914) & (g2211) & (g4422) & (!g4423) & (key[83])) + ((!g830) & (g1914) & (g2211) & (g4422) & (g4423) & (key[83])) + ((g830) & (!g1914) & (!g2211) & (!g4422) & (g4423) & (!key[83])) + ((g830) & (!g1914) & (!g2211) & (!g4422) & (g4423) & (key[83])) + ((g830) & (!g1914) & (!g2211) & (g4422) & (g4423) & (!key[83])) + ((g830) & (!g1914) & (!g2211) & (g4422) & (g4423) & (key[83])) + ((g830) & (!g1914) & (g2211) & (!g4422) & (!g4423) & (!key[83])) + ((g830) & (!g1914) & (g2211) & (!g4422) & (!g4423) & (key[83])) + ((g830) & (!g1914) & (g2211) & (g4422) & (!g4423) & (!key[83])) + ((g830) & (!g1914) & (g2211) & (g4422) & (!g4423) & (key[83])) + ((g830) & (g1914) & (!g2211) & (g4422) & (!g4423) & (!key[83])) + ((g830) & (g1914) & (!g2211) & (g4422) & (!g4423) & (key[83])) + ((g830) & (g1914) & (!g2211) & (g4422) & (g4423) & (!key[83])) + ((g830) & (g1914) & (!g2211) & (g4422) & (g4423) & (key[83])) + ((g830) & (g1914) & (g2211) & (!g4422) & (!g4423) & (!key[83])) + ((g830) & (g1914) & (g2211) & (!g4422) & (!g4423) & (key[83])) + ((g830) & (g1914) & (g2211) & (!g4422) & (g4423) & (!key[83])) + ((g830) & (g1914) & (g2211) & (!g4422) & (g4423) & (key[83])));
	assign g4425 = (((!g4374) & (!g2354) & (!g2358) & (!g2390) & (g2413)) + ((!g4374) & (!g2354) & (!g2358) & (g2390) & (!g2413)) + ((!g4374) & (!g2354) & (g2358) & (!g2390) & (g2413)) + ((!g4374) & (!g2354) & (g2358) & (g2390) & (!g2413)) + ((!g4374) & (g2354) & (!g2358) & (!g2390) & (g2413)) + ((!g4374) & (g2354) & (!g2358) & (g2390) & (!g2413)) + ((!g4374) & (g2354) & (g2358) & (!g2390) & (!g2413)) + ((!g4374) & (g2354) & (g2358) & (g2390) & (g2413)) + ((g4374) & (!g2354) & (!g2358) & (!g2390) & (g2413)) + ((g4374) & (!g2354) & (!g2358) & (g2390) & (!g2413)) + ((g4374) & (!g2354) & (g2358) & (!g2390) & (!g2413)) + ((g4374) & (!g2354) & (g2358) & (g2390) & (g2413)) + ((g4374) & (g2354) & (!g2358) & (!g2390) & (!g2413)) + ((g4374) & (g2354) & (!g2358) & (g2390) & (g2413)) + ((g4374) & (g2354) & (g2358) & (!g2390) & (!g2413)) + ((g4374) & (g2354) & (g2358) & (g2390) & (g2413)));
	assign g8301 = (((!g5560) & (g5596) & (!g4426)) + ((!g5560) & (g5596) & (g4426)) + ((g5560) & (!g5596) & (g4426)) + ((g5560) & (g5596) & (g4426)));
	assign g4427 = (((!g830) & (!g2212) & (!g6737) & (g4426)) + ((!g830) & (!g2212) & (g6737) & (g4426)) + ((!g830) & (g2212) & (!g6737) & (g4426)) + ((!g830) & (g2212) & (g6737) & (g4426)) + ((g830) & (!g2212) & (g6737) & (!g4426)) + ((g830) & (!g2212) & (g6737) & (g4426)) + ((g830) & (g2212) & (!g6737) & (!g4426)) + ((g830) & (g2212) & (!g6737) & (g4426)));
	assign g4428 = (((!g4379) & (!g2497) & (!g2509) & (!g2531) & (g2546)) + ((!g4379) & (!g2497) & (!g2509) & (g2531) & (!g2546)) + ((!g4379) & (!g2497) & (g2509) & (!g2531) & (!g2546)) + ((!g4379) & (!g2497) & (g2509) & (g2531) & (g2546)) + ((!g4379) & (g2497) & (!g2509) & (!g2531) & (!g2546)) + ((!g4379) & (g2497) & (!g2509) & (g2531) & (g2546)) + ((!g4379) & (g2497) & (g2509) & (!g2531) & (!g2546)) + ((!g4379) & (g2497) & (g2509) & (g2531) & (g2546)) + ((g4379) & (!g2497) & (!g2509) & (!g2531) & (g2546)) + ((g4379) & (!g2497) & (!g2509) & (g2531) & (!g2546)) + ((g4379) & (!g2497) & (g2509) & (!g2531) & (g2546)) + ((g4379) & (!g2497) & (g2509) & (g2531) & (!g2546)) + ((g4379) & (g2497) & (!g2509) & (!g2531) & (g2546)) + ((g4379) & (g2497) & (!g2509) & (g2531) & (!g2546)) + ((g4379) & (g2497) & (g2509) & (!g2531) & (!g2546)) + ((g4379) & (g2497) & (g2509) & (g2531) & (g2546)));
	assign g4429 = (((!g3485) & (!g3486)));
	assign g4430 = (((!g1991) & (!g2217) & (!g4429)) + ((!g1991) & (g2217) & (g4429)) + ((g1991) & (!g2217) & (g4429)) + ((g1991) & (g2217) & (!g4429)));
	assign g4431 = (((!g830) & (!g1914) & (!g2213) & (!g4428) & (!g4430) & (key[179])) + ((!g830) & (!g1914) & (!g2213) & (!g4428) & (g4430) & (key[179])) + ((!g830) & (!g1914) & (!g2213) & (g4428) & (!g4430) & (key[179])) + ((!g830) & (!g1914) & (!g2213) & (g4428) & (g4430) & (key[179])) + ((!g830) & (!g1914) & (g2213) & (!g4428) & (!g4430) & (key[179])) + ((!g830) & (!g1914) & (g2213) & (!g4428) & (g4430) & (key[179])) + ((!g830) & (!g1914) & (g2213) & (g4428) & (!g4430) & (key[179])) + ((!g830) & (!g1914) & (g2213) & (g4428) & (g4430) & (key[179])) + ((!g830) & (g1914) & (!g2213) & (!g4428) & (!g4430) & (key[179])) + ((!g830) & (g1914) & (!g2213) & (!g4428) & (g4430) & (key[179])) + ((!g830) & (g1914) & (!g2213) & (g4428) & (!g4430) & (key[179])) + ((!g830) & (g1914) & (!g2213) & (g4428) & (g4430) & (key[179])) + ((!g830) & (g1914) & (g2213) & (!g4428) & (!g4430) & (key[179])) + ((!g830) & (g1914) & (g2213) & (!g4428) & (g4430) & (key[179])) + ((!g830) & (g1914) & (g2213) & (g4428) & (!g4430) & (key[179])) + ((!g830) & (g1914) & (g2213) & (g4428) & (g4430) & (key[179])) + ((g830) & (!g1914) & (!g2213) & (!g4428) & (g4430) & (!key[179])) + ((g830) & (!g1914) & (!g2213) & (!g4428) & (g4430) & (key[179])) + ((g830) & (!g1914) & (!g2213) & (g4428) & (g4430) & (!key[179])) + ((g830) & (!g1914) & (!g2213) & (g4428) & (g4430) & (key[179])) + ((g830) & (!g1914) & (g2213) & (!g4428) & (!g4430) & (!key[179])) + ((g830) & (!g1914) & (g2213) & (!g4428) & (!g4430) & (key[179])) + ((g830) & (!g1914) & (g2213) & (g4428) & (!g4430) & (!key[179])) + ((g830) & (!g1914) & (g2213) & (g4428) & (!g4430) & (key[179])) + ((g830) & (g1914) & (!g2213) & (g4428) & (!g4430) & (!key[179])) + ((g830) & (g1914) & (!g2213) & (g4428) & (!g4430) & (key[179])) + ((g830) & (g1914) & (!g2213) & (g4428) & (g4430) & (!key[179])) + ((g830) & (g1914) & (!g2213) & (g4428) & (g4430) & (key[179])) + ((g830) & (g1914) & (g2213) & (!g4428) & (!g4430) & (!key[179])) + ((g830) & (g1914) & (g2213) & (!g4428) & (!g4430) & (key[179])) + ((g830) & (g1914) & (g2213) & (!g4428) & (g4430) & (!key[179])) + ((g830) & (g1914) & (g2213) & (!g4428) & (g4430) & (key[179])));
	assign g4432 = (((!g3080) & (!g3125) & (!g3095) & (!g4395) & (g3131)) + ((!g3080) & (!g3125) & (!g3095) & (g4395) & (g3131)) + ((!g3080) & (!g3125) & (g3095) & (!g4395) & (g3131)) + ((!g3080) & (!g3125) & (g3095) & (g4395) & (!g3131)) + ((!g3080) & (g3125) & (!g3095) & (!g4395) & (!g3131)) + ((!g3080) & (g3125) & (!g3095) & (g4395) & (!g3131)) + ((!g3080) & (g3125) & (g3095) & (!g4395) & (!g3131)) + ((!g3080) & (g3125) & (g3095) & (g4395) & (g3131)) + ((g3080) & (!g3125) & (!g3095) & (!g4395) & (g3131)) + ((g3080) & (!g3125) & (!g3095) & (g4395) & (!g3131)) + ((g3080) & (!g3125) & (g3095) & (!g4395) & (!g3131)) + ((g3080) & (!g3125) & (g3095) & (g4395) & (!g3131)) + ((g3080) & (g3125) & (!g3095) & (!g4395) & (!g3131)) + ((g3080) & (g3125) & (!g3095) & (g4395) & (g3131)) + ((g3080) & (g3125) & (g3095) & (!g4395) & (g3131)) + ((g3080) & (g3125) & (g3095) & (g4395) & (g3131)));
	assign g4433 = (((!g2761) & (!g2794) & (!g1847) & (g1881) & (!g4396)) + ((!g2761) & (!g2794) & (!g1847) & (g1881) & (g4396)) + ((!g2761) & (!g2794) & (g1847) & (!g1881) & (g4396)) + ((!g2761) & (!g2794) & (g1847) & (g1881) & (!g4396)) + ((!g2761) & (g2794) & (!g1847) & (!g1881) & (!g4396)) + ((!g2761) & (g2794) & (!g1847) & (!g1881) & (g4396)) + ((!g2761) & (g2794) & (g1847) & (!g1881) & (!g4396)) + ((!g2761) & (g2794) & (g1847) & (g1881) & (g4396)) + ((g2761) & (!g2794) & (!g1847) & (!g1881) & (g4396)) + ((g2761) & (!g2794) & (!g1847) & (g1881) & (!g4396)) + ((g2761) & (!g2794) & (g1847) & (!g1881) & (!g4396)) + ((g2761) & (!g2794) & (g1847) & (!g1881) & (g4396)) + ((g2761) & (g2794) & (!g1847) & (!g1881) & (!g4396)) + ((g2761) & (g2794) & (!g1847) & (g1881) & (g4396)) + ((g2761) & (g2794) & (g1847) & (g1881) & (!g4396)) + ((g2761) & (g2794) & (g1847) & (g1881) & (g4396)));
	assign g4434 = (((!g830) & (!g1914) & (!g2217) & (!g4432) & (!g4433) & (key[102])) + ((!g830) & (!g1914) & (!g2217) & (!g4432) & (g4433) & (key[102])) + ((!g830) & (!g1914) & (!g2217) & (g4432) & (!g4433) & (key[102])) + ((!g830) & (!g1914) & (!g2217) & (g4432) & (g4433) & (key[102])) + ((!g830) & (!g1914) & (g2217) & (!g4432) & (!g4433) & (key[102])) + ((!g830) & (!g1914) & (g2217) & (!g4432) & (g4433) & (key[102])) + ((!g830) & (!g1914) & (g2217) & (g4432) & (!g4433) & (key[102])) + ((!g830) & (!g1914) & (g2217) & (g4432) & (g4433) & (key[102])) + ((!g830) & (g1914) & (!g2217) & (!g4432) & (!g4433) & (key[102])) + ((!g830) & (g1914) & (!g2217) & (!g4432) & (g4433) & (key[102])) + ((!g830) & (g1914) & (!g2217) & (g4432) & (!g4433) & (key[102])) + ((!g830) & (g1914) & (!g2217) & (g4432) & (g4433) & (key[102])) + ((!g830) & (g1914) & (g2217) & (!g4432) & (!g4433) & (key[102])) + ((!g830) & (g1914) & (g2217) & (!g4432) & (g4433) & (key[102])) + ((!g830) & (g1914) & (g2217) & (g4432) & (!g4433) & (key[102])) + ((!g830) & (g1914) & (g2217) & (g4432) & (g4433) & (key[102])) + ((g830) & (!g1914) & (!g2217) & (!g4432) & (g4433) & (!key[102])) + ((g830) & (!g1914) & (!g2217) & (!g4432) & (g4433) & (key[102])) + ((g830) & (!g1914) & (!g2217) & (g4432) & (g4433) & (!key[102])) + ((g830) & (!g1914) & (!g2217) & (g4432) & (g4433) & (key[102])) + ((g830) & (!g1914) & (g2217) & (!g4432) & (!g4433) & (!key[102])) + ((g830) & (!g1914) & (g2217) & (!g4432) & (!g4433) & (key[102])) + ((g830) & (!g1914) & (g2217) & (g4432) & (!g4433) & (!key[102])) + ((g830) & (!g1914) & (g2217) & (g4432) & (!g4433) & (key[102])) + ((g830) & (g1914) & (!g2217) & (g4432) & (!g4433) & (!key[102])) + ((g830) & (g1914) & (!g2217) & (g4432) & (!g4433) & (key[102])) + ((g830) & (g1914) & (!g2217) & (g4432) & (g4433) & (!key[102])) + ((g830) & (g1914) & (!g2217) & (g4432) & (g4433) & (key[102])) + ((g830) & (g1914) & (g2217) & (!g4432) & (!g4433) & (!key[102])) + ((g830) & (g1914) & (g2217) & (!g4432) & (!g4433) & (key[102])) + ((g830) & (g1914) & (g2217) & (!g4432) & (g4433) & (!key[102])) + ((g830) & (g1914) & (g2217) & (!g4432) & (g4433) & (key[102])));
	assign g4435 = (((!g2212) & (!g2262) & (!g2848) & (g2893) & (!g4386)) + ((!g2212) & (!g2262) & (!g2848) & (g2893) & (g4386)) + ((!g2212) & (!g2262) & (g2848) & (!g2893) & (g4386)) + ((!g2212) & (!g2262) & (g2848) & (g2893) & (!g4386)) + ((!g2212) & (g2262) & (!g2848) & (!g2893) & (!g4386)) + ((!g2212) & (g2262) & (!g2848) & (!g2893) & (g4386)) + ((!g2212) & (g2262) & (g2848) & (!g2893) & (!g4386)) + ((!g2212) & (g2262) & (g2848) & (g2893) & (g4386)) + ((g2212) & (!g2262) & (!g2848) & (!g2893) & (g4386)) + ((g2212) & (!g2262) & (!g2848) & (g2893) & (!g4386)) + ((g2212) & (!g2262) & (g2848) & (!g2893) & (!g4386)) + ((g2212) & (!g2262) & (g2848) & (!g2893) & (g4386)) + ((g2212) & (g2262) & (!g2848) & (!g2893) & (!g4386)) + ((g2212) & (g2262) & (!g2848) & (g2893) & (g4386)) + ((g2212) & (g2262) & (g2848) & (g2893) & (!g4386)) + ((g2212) & (g2262) & (g2848) & (g2893) & (g4386)));
	assign g4436 = (((!g2047) & (!g2665) & (!g4121) & (g5778) & (!g5779) & (!g5780)) + ((!g2047) & (!g2665) & (!g4121) & (g5778) & (!g5779) & (g5780)) + ((!g2047) & (!g2665) & (g4121) & (g5778) & (!g5779) & (!g5780)) + ((!g2047) & (!g2665) & (g4121) & (g5778) & (!g5779) & (g5780)) + ((!g2047) & (g2665) & (!g4121) & (g5778) & (!g5779) & (!g5780)) + ((!g2047) & (g2665) & (!g4121) & (g5778) & (!g5779) & (g5780)) + ((!g2047) & (g2665) & (g4121) & (g5778) & (!g5779) & (!g5780)) + ((!g2047) & (g2665) & (g4121) & (g5778) & (!g5779) & (g5780)) + ((!g2047) & (g2665) & (g4121) & (g5778) & (g5779) & (!g5780)) + ((g2047) & (!g2665) & (!g4121) & (g5778) & (!g5779) & (!g5780)) + ((g2047) & (!g2665) & (!g4121) & (g5778) & (!g5779) & (g5780)) + ((g2047) & (!g2665) & (g4121) & (g5778) & (!g5779) & (!g5780)) + ((g2047) & (!g2665) & (g4121) & (g5778) & (!g5779) & (g5780)) + ((g2047) & (!g2665) & (g4121) & (g5778) & (g5779) & (!g5780)) + ((g2047) & (g2665) & (!g4121) & (g5778) & (!g5779) & (!g5780)) + ((g2047) & (g2665) & (!g4121) & (g5778) & (!g5779) & (g5780)) + ((g2047) & (g2665) & (!g4121) & (g5778) & (g5779) & (!g5780)) + ((g2047) & (g2665) & (g4121) & (g5778) & (!g5779) & (!g5780)) + ((g2047) & (g2665) & (g4121) & (g5778) & (!g5779) & (g5780)) + ((g2047) & (g2665) & (g4121) & (g5778) & (g5779) & (!g5780)));
	assign g4437 = (((g2210) & (g2857)));
	assign g4438 = (((!g2256) & (!g2887) & (!g4436) & (g4437)) + ((!g2256) & (!g2887) & (g4436) & (!g4437)) + ((!g2256) & (!g2887) & (g4436) & (g4437)) + ((!g2256) & (g2887) & (!g4436) & (!g4437)) + ((g2256) & (!g2887) & (!g4436) & (!g4437)) + ((g2256) & (g2887) & (!g4436) & (g4437)) + ((g2256) & (g2887) & (g4436) & (!g4437)) + ((g2256) & (g2887) & (g4436) & (g4437)));
	assign g4439 = (((g830) & (!g1914) & (!g2224) & (!g4435) & (g4438)) + ((g830) & (!g1914) & (!g2224) & (g4435) & (g4438)) + ((g830) & (!g1914) & (g2224) & (!g4435) & (!g4438)) + ((g830) & (!g1914) & (g2224) & (g4435) & (!g4438)) + ((g830) & (g1914) & (!g2224) & (g4435) & (!g4438)) + ((g830) & (g1914) & (!g2224) & (g4435) & (g4438)) + ((g830) & (g1914) & (g2224) & (!g4435) & (!g4438)) + ((g830) & (g1914) & (g2224) & (!g4435) & (g4438)));
	assign g4440 = (((!g3345) & (!g4398) & (!g3323) & (!g3376) & (g3380)) + ((!g3345) & (!g4398) & (!g3323) & (g3376) & (!g3380)) + ((!g3345) & (!g4398) & (g3323) & (!g3376) & (g3380)) + ((!g3345) & (!g4398) & (g3323) & (g3376) & (!g3380)) + ((!g3345) & (g4398) & (!g3323) & (!g3376) & (g3380)) + ((!g3345) & (g4398) & (!g3323) & (g3376) & (!g3380)) + ((!g3345) & (g4398) & (g3323) & (!g3376) & (!g3380)) + ((!g3345) & (g4398) & (g3323) & (g3376) & (g3380)) + ((g3345) & (!g4398) & (!g3323) & (!g3376) & (g3380)) + ((g3345) & (!g4398) & (!g3323) & (g3376) & (!g3380)) + ((g3345) & (!g4398) & (g3323) & (!g3376) & (!g3380)) + ((g3345) & (!g4398) & (g3323) & (g3376) & (g3380)) + ((g3345) & (g4398) & (!g3323) & (!g3376) & (!g3380)) + ((g3345) & (g4398) & (!g3323) & (g3376) & (g3380)) + ((g3345) & (g4398) & (g3323) & (!g3376) & (!g3380)) + ((g3345) & (g4398) & (g3323) & (g3376) & (g3380)));
	assign g4441 = (((!g2423) & (!g2515) & (!g3082) & (g3136) & (!g4399)) + ((!g2423) & (!g2515) & (!g3082) & (g3136) & (g4399)) + ((!g2423) & (!g2515) & (g3082) & (!g3136) & (g4399)) + ((!g2423) & (!g2515) & (g3082) & (g3136) & (!g4399)) + ((!g2423) & (g2515) & (!g3082) & (!g3136) & (!g4399)) + ((!g2423) & (g2515) & (!g3082) & (!g3136) & (g4399)) + ((!g2423) & (g2515) & (g3082) & (!g3136) & (!g4399)) + ((!g2423) & (g2515) & (g3082) & (g3136) & (g4399)) + ((g2423) & (!g2515) & (!g3082) & (!g3136) & (g4399)) + ((g2423) & (!g2515) & (!g3082) & (g3136) & (!g4399)) + ((g2423) & (!g2515) & (g3082) & (!g3136) & (!g4399)) + ((g2423) & (!g2515) & (g3082) & (!g3136) & (g4399)) + ((g2423) & (g2515) & (!g3082) & (!g3136) & (!g4399)) + ((g2423) & (g2515) & (!g3082) & (g3136) & (g4399)) + ((g2423) & (g2515) & (g3082) & (g3136) & (!g4399)) + ((g2423) & (g2515) & (g3082) & (g3136) & (g4399)));
	assign g4442 = (((!g830) & (!g1914) & (!g2227) & (!g4440) & (!g4441) & (nonce[6])) + ((!g830) & (!g1914) & (!g2227) & (!g4440) & (g4441) & (nonce[6])) + ((!g830) & (!g1914) & (!g2227) & (g4440) & (!g4441) & (nonce[6])) + ((!g830) & (!g1914) & (!g2227) & (g4440) & (g4441) & (nonce[6])) + ((!g830) & (!g1914) & (g2227) & (!g4440) & (!g4441) & (nonce[6])) + ((!g830) & (!g1914) & (g2227) & (!g4440) & (g4441) & (nonce[6])) + ((!g830) & (!g1914) & (g2227) & (g4440) & (!g4441) & (nonce[6])) + ((!g830) & (!g1914) & (g2227) & (g4440) & (g4441) & (nonce[6])) + ((!g830) & (g1914) & (!g2227) & (!g4440) & (!g4441) & (nonce[6])) + ((!g830) & (g1914) & (!g2227) & (!g4440) & (g4441) & (nonce[6])) + ((!g830) & (g1914) & (!g2227) & (g4440) & (!g4441) & (nonce[6])) + ((!g830) & (g1914) & (!g2227) & (g4440) & (g4441) & (nonce[6])) + ((!g830) & (g1914) & (g2227) & (!g4440) & (!g4441) & (nonce[6])) + ((!g830) & (g1914) & (g2227) & (!g4440) & (g4441) & (nonce[6])) + ((!g830) & (g1914) & (g2227) & (g4440) & (!g4441) & (nonce[6])) + ((!g830) & (g1914) & (g2227) & (g4440) & (g4441) & (nonce[6])) + ((g830) & (!g1914) & (!g2227) & (!g4440) & (g4441) & (!nonce[6])) + ((g830) & (!g1914) & (!g2227) & (!g4440) & (g4441) & (nonce[6])) + ((g830) & (!g1914) & (!g2227) & (g4440) & (g4441) & (!nonce[6])) + ((g830) & (!g1914) & (!g2227) & (g4440) & (g4441) & (nonce[6])) + ((g830) & (!g1914) & (g2227) & (!g4440) & (!g4441) & (!nonce[6])) + ((g830) & (!g1914) & (g2227) & (!g4440) & (!g4441) & (nonce[6])) + ((g830) & (!g1914) & (g2227) & (g4440) & (!g4441) & (!nonce[6])) + ((g830) & (!g1914) & (g2227) & (g4440) & (!g4441) & (nonce[6])) + ((g830) & (g1914) & (!g2227) & (g4440) & (!g4441) & (!nonce[6])) + ((g830) & (g1914) & (!g2227) & (g4440) & (!g4441) & (nonce[6])) + ((g830) & (g1914) & (!g2227) & (g4440) & (g4441) & (!nonce[6])) + ((g830) & (g1914) & (!g2227) & (g4440) & (g4441) & (nonce[6])) + ((g830) & (g1914) & (g2227) & (!g4440) & (!g4441) & (!nonce[6])) + ((g830) & (g1914) & (g2227) & (!g4440) & (!g4441) & (nonce[6])) + ((g830) & (g1914) & (g2227) & (!g4440) & (g4441) & (!nonce[6])) + ((g830) & (g1914) & (g2227) & (!g4440) & (g4441) & (nonce[6])));
	assign g4443 = (((!g2427) & (!g2519) & (!g3090) & (!g4408) & (g3139)) + ((!g2427) & (!g2519) & (!g3090) & (g4408) & (g3139)) + ((!g2427) & (!g2519) & (g3090) & (!g4408) & (g3139)) + ((!g2427) & (!g2519) & (g3090) & (g4408) & (!g3139)) + ((!g2427) & (g2519) & (!g3090) & (!g4408) & (!g3139)) + ((!g2427) & (g2519) & (!g3090) & (g4408) & (!g3139)) + ((!g2427) & (g2519) & (g3090) & (!g4408) & (!g3139)) + ((!g2427) & (g2519) & (g3090) & (g4408) & (g3139)) + ((g2427) & (!g2519) & (!g3090) & (!g4408) & (g3139)) + ((g2427) & (!g2519) & (!g3090) & (g4408) & (!g3139)) + ((g2427) & (!g2519) & (g3090) & (!g4408) & (!g3139)) + ((g2427) & (!g2519) & (g3090) & (g4408) & (!g3139)) + ((g2427) & (g2519) & (!g3090) & (!g4408) & (!g3139)) + ((g2427) & (g2519) & (!g3090) & (g4408) & (g3139)) + ((g2427) & (g2519) & (g3090) & (!g4408) & (g3139)) + ((g2427) & (g2519) & (g3090) & (g4408) & (g3139)));
	assign g4444 = (((!g3330) & (!g4409) & (!g3333) & (!g3370) & (g3378)) + ((!g3330) & (!g4409) & (!g3333) & (g3370) & (!g3378)) + ((!g3330) & (!g4409) & (g3333) & (!g3370) & (g3378)) + ((!g3330) & (!g4409) & (g3333) & (g3370) & (!g3378)) + ((!g3330) & (g4409) & (!g3333) & (!g3370) & (g3378)) + ((!g3330) & (g4409) & (!g3333) & (g3370) & (!g3378)) + ((!g3330) & (g4409) & (g3333) & (!g3370) & (!g3378)) + ((!g3330) & (g4409) & (g3333) & (g3370) & (g3378)) + ((g3330) & (!g4409) & (!g3333) & (!g3370) & (g3378)) + ((g3330) & (!g4409) & (!g3333) & (g3370) & (!g3378)) + ((g3330) & (!g4409) & (g3333) & (!g3370) & (!g3378)) + ((g3330) & (!g4409) & (g3333) & (g3370) & (g3378)) + ((g3330) & (g4409) & (!g3333) & (!g3370) & (!g3378)) + ((g3330) & (g4409) & (!g3333) & (g3370) & (g3378)) + ((g3330) & (g4409) & (g3333) & (!g3370) & (!g3378)) + ((g3330) & (g4409) & (g3333) & (g3370) & (g3378)));
	assign g4445 = (((!g830) & (!g1914) & (!g2230) & (!g4443) & (!g4444) & (key[230])) + ((!g830) & (!g1914) & (!g2230) & (!g4443) & (g4444) & (key[230])) + ((!g830) & (!g1914) & (!g2230) & (g4443) & (!g4444) & (key[230])) + ((!g830) & (!g1914) & (!g2230) & (g4443) & (g4444) & (key[230])) + ((!g830) & (!g1914) & (g2230) & (!g4443) & (!g4444) & (key[230])) + ((!g830) & (!g1914) & (g2230) & (!g4443) & (g4444) & (key[230])) + ((!g830) & (!g1914) & (g2230) & (g4443) & (!g4444) & (key[230])) + ((!g830) & (!g1914) & (g2230) & (g4443) & (g4444) & (key[230])) + ((!g830) & (g1914) & (!g2230) & (!g4443) & (!g4444) & (key[230])) + ((!g830) & (g1914) & (!g2230) & (!g4443) & (g4444) & (key[230])) + ((!g830) & (g1914) & (!g2230) & (g4443) & (!g4444) & (key[230])) + ((!g830) & (g1914) & (!g2230) & (g4443) & (g4444) & (key[230])) + ((!g830) & (g1914) & (g2230) & (!g4443) & (!g4444) & (key[230])) + ((!g830) & (g1914) & (g2230) & (!g4443) & (g4444) & (key[230])) + ((!g830) & (g1914) & (g2230) & (g4443) & (!g4444) & (key[230])) + ((!g830) & (g1914) & (g2230) & (g4443) & (g4444) & (key[230])) + ((g830) & (!g1914) & (!g2230) & (!g4443) & (g4444) & (!key[230])) + ((g830) & (!g1914) & (!g2230) & (!g4443) & (g4444) & (key[230])) + ((g830) & (!g1914) & (!g2230) & (g4443) & (g4444) & (!key[230])) + ((g830) & (!g1914) & (!g2230) & (g4443) & (g4444) & (key[230])) + ((g830) & (!g1914) & (g2230) & (!g4443) & (!g4444) & (!key[230])) + ((g830) & (!g1914) & (g2230) & (!g4443) & (!g4444) & (key[230])) + ((g830) & (!g1914) & (g2230) & (g4443) & (!g4444) & (!key[230])) + ((g830) & (!g1914) & (g2230) & (g4443) & (!g4444) & (key[230])) + ((g830) & (g1914) & (!g2230) & (g4443) & (!g4444) & (!key[230])) + ((g830) & (g1914) & (!g2230) & (g4443) & (!g4444) & (key[230])) + ((g830) & (g1914) & (!g2230) & (g4443) & (g4444) & (!key[230])) + ((g830) & (g1914) & (!g2230) & (g4443) & (g4444) & (key[230])) + ((g830) & (g1914) & (g2230) & (!g4443) & (!g4444) & (!key[230])) + ((g830) & (g1914) & (g2230) & (!g4443) & (!g4444) & (key[230])) + ((g830) & (g1914) & (g2230) & (!g4443) & (g4444) & (!key[230])) + ((g830) & (g1914) & (g2230) & (!g4443) & (g4444) & (key[230])));
	assign g4446 = (((!g2759) & (!g2790) & (!g1847) & (g1881) & (!g4383)) + ((!g2759) & (!g2790) & (!g1847) & (g1881) & (g4383)) + ((!g2759) & (!g2790) & (g1847) & (!g1881) & (g4383)) + ((!g2759) & (!g2790) & (g1847) & (g1881) & (!g4383)) + ((!g2759) & (g2790) & (!g1847) & (!g1881) & (!g4383)) + ((!g2759) & (g2790) & (!g1847) & (!g1881) & (g4383)) + ((!g2759) & (g2790) & (g1847) & (!g1881) & (!g4383)) + ((!g2759) & (g2790) & (g1847) & (g1881) & (g4383)) + ((g2759) & (!g2790) & (!g1847) & (!g1881) & (g4383)) + ((g2759) & (!g2790) & (!g1847) & (g1881) & (!g4383)) + ((g2759) & (!g2790) & (g1847) & (!g1881) & (!g4383)) + ((g2759) & (!g2790) & (g1847) & (!g1881) & (g4383)) + ((g2759) & (g2790) & (!g1847) & (!g1881) & (!g4383)) + ((g2759) & (g2790) & (!g1847) & (g1881) & (g4383)) + ((g2759) & (g2790) & (g1847) & (g1881) & (!g4383)) + ((g2759) & (g2790) & (g1847) & (g1881) & (g4383)));
	assign g4447 = (((!g3086) & (!g3116) & (!g4384) & (!g3090) & (g3139)) + ((!g3086) & (!g3116) & (!g4384) & (g3090) & (g3139)) + ((!g3086) & (!g3116) & (g4384) & (!g3090) & (g3139)) + ((!g3086) & (!g3116) & (g4384) & (g3090) & (!g3139)) + ((!g3086) & (g3116) & (!g4384) & (!g3090) & (!g3139)) + ((!g3086) & (g3116) & (!g4384) & (g3090) & (!g3139)) + ((!g3086) & (g3116) & (g4384) & (!g3090) & (!g3139)) + ((!g3086) & (g3116) & (g4384) & (g3090) & (g3139)) + ((g3086) & (!g3116) & (!g4384) & (!g3090) & (g3139)) + ((g3086) & (!g3116) & (!g4384) & (g3090) & (!g3139)) + ((g3086) & (!g3116) & (g4384) & (!g3090) & (!g3139)) + ((g3086) & (!g3116) & (g4384) & (g3090) & (!g3139)) + ((g3086) & (g3116) & (!g4384) & (!g3090) & (!g3139)) + ((g3086) & (g3116) & (!g4384) & (g3090) & (g3139)) + ((g3086) & (g3116) & (g4384) & (!g3090) & (g3139)) + ((g3086) & (g3116) & (g4384) & (g3090) & (g3139)));
	assign g4448 = (((!g830) & (!g1914) & (!g2233) & (!g4446) & (!g4447) & (key[6])) + ((!g830) & (!g1914) & (!g2233) & (!g4446) & (g4447) & (key[6])) + ((!g830) & (!g1914) & (!g2233) & (g4446) & (!g4447) & (key[6])) + ((!g830) & (!g1914) & (!g2233) & (g4446) & (g4447) & (key[6])) + ((!g830) & (!g1914) & (g2233) & (!g4446) & (!g4447) & (key[6])) + ((!g830) & (!g1914) & (g2233) & (!g4446) & (g4447) & (key[6])) + ((!g830) & (!g1914) & (g2233) & (g4446) & (!g4447) & (key[6])) + ((!g830) & (!g1914) & (g2233) & (g4446) & (g4447) & (key[6])) + ((!g830) & (g1914) & (!g2233) & (!g4446) & (!g4447) & (key[6])) + ((!g830) & (g1914) & (!g2233) & (!g4446) & (g4447) & (key[6])) + ((!g830) & (g1914) & (!g2233) & (g4446) & (!g4447) & (key[6])) + ((!g830) & (g1914) & (!g2233) & (g4446) & (g4447) & (key[6])) + ((!g830) & (g1914) & (g2233) & (!g4446) & (!g4447) & (key[6])) + ((!g830) & (g1914) & (g2233) & (!g4446) & (g4447) & (key[6])) + ((!g830) & (g1914) & (g2233) & (g4446) & (!g4447) & (key[6])) + ((!g830) & (g1914) & (g2233) & (g4446) & (g4447) & (key[6])) + ((g830) & (!g1914) & (!g2233) & (!g4446) & (g4447) & (!key[6])) + ((g830) & (!g1914) & (!g2233) & (!g4446) & (g4447) & (key[6])) + ((g830) & (!g1914) & (!g2233) & (g4446) & (g4447) & (!key[6])) + ((g830) & (!g1914) & (!g2233) & (g4446) & (g4447) & (key[6])) + ((g830) & (!g1914) & (g2233) & (!g4446) & (!g4447) & (!key[6])) + ((g830) & (!g1914) & (g2233) & (!g4446) & (!g4447) & (key[6])) + ((g830) & (!g1914) & (g2233) & (g4446) & (!g4447) & (!key[6])) + ((g830) & (!g1914) & (g2233) & (g4446) & (!g4447) & (key[6])) + ((g830) & (g1914) & (!g2233) & (g4446) & (!g4447) & (!key[6])) + ((g830) & (g1914) & (!g2233) & (g4446) & (!g4447) & (key[6])) + ((g830) & (g1914) & (!g2233) & (g4446) & (g4447) & (!key[6])) + ((g830) & (g1914) & (!g2233) & (g4446) & (g4447) & (key[6])) + ((g830) & (g1914) & (g2233) & (!g4446) & (!g4447) & (!key[6])) + ((g830) & (g1914) & (g2233) & (!g4446) & (!g4447) & (key[6])) + ((g830) & (g1914) & (g2233) & (!g4446) & (g4447) & (!key[6])) + ((g830) & (g1914) & (g2233) & (!g4446) & (g4447) & (key[6])));
	assign g4449 = (((!g2426) & (!g2518) & (!g3093) & (g3119) & (!g4388)) + ((!g2426) & (!g2518) & (!g3093) & (g3119) & (g4388)) + ((!g2426) & (!g2518) & (g3093) & (!g3119) & (g4388)) + ((!g2426) & (!g2518) & (g3093) & (g3119) & (!g4388)) + ((!g2426) & (g2518) & (!g3093) & (!g3119) & (!g4388)) + ((!g2426) & (g2518) & (!g3093) & (!g3119) & (g4388)) + ((!g2426) & (g2518) & (g3093) & (!g3119) & (!g4388)) + ((!g2426) & (g2518) & (g3093) & (g3119) & (g4388)) + ((g2426) & (!g2518) & (!g3093) & (!g3119) & (g4388)) + ((g2426) & (!g2518) & (!g3093) & (g3119) & (!g4388)) + ((g2426) & (!g2518) & (g3093) & (!g3119) & (!g4388)) + ((g2426) & (!g2518) & (g3093) & (!g3119) & (g4388)) + ((g2426) & (g2518) & (!g3093) & (!g3119) & (!g4388)) + ((g2426) & (g2518) & (!g3093) & (g3119) & (g4388)) + ((g2426) & (g2518) & (g3093) & (g3119) & (!g4388)) + ((g2426) & (g2518) & (g3093) & (g3119) & (g4388)));
	assign g4450 = (((!g4389) & (!g3339) & (!g3345) & (!g3380) & (g3366)) + ((!g4389) & (!g3339) & (!g3345) & (g3380) & (!g3366)) + ((!g4389) & (!g3339) & (g3345) & (!g3380) & (g3366)) + ((!g4389) & (!g3339) & (g3345) & (g3380) & (!g3366)) + ((!g4389) & (g3339) & (!g3345) & (!g3380) & (g3366)) + ((!g4389) & (g3339) & (!g3345) & (g3380) & (!g3366)) + ((!g4389) & (g3339) & (g3345) & (!g3380) & (!g3366)) + ((!g4389) & (g3339) & (g3345) & (g3380) & (g3366)) + ((g4389) & (!g3339) & (!g3345) & (!g3380) & (g3366)) + ((g4389) & (!g3339) & (!g3345) & (g3380) & (!g3366)) + ((g4389) & (!g3339) & (g3345) & (!g3380) & (!g3366)) + ((g4389) & (!g3339) & (g3345) & (g3380) & (g3366)) + ((g4389) & (g3339) & (!g3345) & (!g3380) & (!g3366)) + ((g4389) & (g3339) & (!g3345) & (g3380) & (g3366)) + ((g4389) & (g3339) & (g3345) & (!g3380) & (!g3366)) + ((g4389) & (g3339) & (g3345) & (g3380) & (g3366)));
	assign g8302 = (((!g5560) & (g5598) & (!g4451)) + ((!g5560) & (g5598) & (g4451)) + ((g5560) & (!g5598) & (g4451)) + ((g5560) & (g5598) & (g4451)));
	assign g4452 = (((!g830) & (!g1914) & (!g2236) & (!g4449) & (!g4450) & (g4451)) + ((!g830) & (!g1914) & (!g2236) & (!g4449) & (g4450) & (g4451)) + ((!g830) & (!g1914) & (!g2236) & (g4449) & (!g4450) & (g4451)) + ((!g830) & (!g1914) & (!g2236) & (g4449) & (g4450) & (g4451)) + ((!g830) & (!g1914) & (g2236) & (!g4449) & (!g4450) & (g4451)) + ((!g830) & (!g1914) & (g2236) & (!g4449) & (g4450) & (g4451)) + ((!g830) & (!g1914) & (g2236) & (g4449) & (!g4450) & (g4451)) + ((!g830) & (!g1914) & (g2236) & (g4449) & (g4450) & (g4451)) + ((!g830) & (g1914) & (!g2236) & (!g4449) & (!g4450) & (g4451)) + ((!g830) & (g1914) & (!g2236) & (!g4449) & (g4450) & (g4451)) + ((!g830) & (g1914) & (!g2236) & (g4449) & (!g4450) & (g4451)) + ((!g830) & (g1914) & (!g2236) & (g4449) & (g4450) & (g4451)) + ((!g830) & (g1914) & (g2236) & (!g4449) & (!g4450) & (g4451)) + ((!g830) & (g1914) & (g2236) & (!g4449) & (g4450) & (g4451)) + ((!g830) & (g1914) & (g2236) & (g4449) & (!g4450) & (g4451)) + ((!g830) & (g1914) & (g2236) & (g4449) & (g4450) & (g4451)) + ((g830) & (!g1914) & (!g2236) & (!g4449) & (g4450) & (!g4451)) + ((g830) & (!g1914) & (!g2236) & (!g4449) & (g4450) & (g4451)) + ((g830) & (!g1914) & (!g2236) & (g4449) & (g4450) & (!g4451)) + ((g830) & (!g1914) & (!g2236) & (g4449) & (g4450) & (g4451)) + ((g830) & (!g1914) & (g2236) & (!g4449) & (!g4450) & (!g4451)) + ((g830) & (!g1914) & (g2236) & (!g4449) & (!g4450) & (g4451)) + ((g830) & (!g1914) & (g2236) & (g4449) & (!g4450) & (!g4451)) + ((g830) & (!g1914) & (g2236) & (g4449) & (!g4450) & (g4451)) + ((g830) & (g1914) & (!g2236) & (g4449) & (!g4450) & (!g4451)) + ((g830) & (g1914) & (!g2236) & (g4449) & (!g4450) & (g4451)) + ((g830) & (g1914) & (!g2236) & (g4449) & (g4450) & (!g4451)) + ((g830) & (g1914) & (!g2236) & (g4449) & (g4450) & (g4451)) + ((g830) & (g1914) & (g2236) & (!g4449) & (!g4450) & (!g4451)) + ((g830) & (g1914) & (g2236) & (!g4449) & (!g4450) & (g4451)) + ((g830) & (g1914) & (g2236) & (!g4449) & (g4450) & (!g4451)) + ((g830) & (g1914) & (g2236) & (!g4449) & (g4450) & (g4451)));
	assign g4453 = (((!g2854) & (!g2881) & (!g2863) & (g2902) & (!g4401)) + ((!g2854) & (!g2881) & (!g2863) & (g2902) & (g4401)) + ((!g2854) & (!g2881) & (g2863) & (!g2902) & (g4401)) + ((!g2854) & (!g2881) & (g2863) & (g2902) & (!g4401)) + ((!g2854) & (g2881) & (!g2863) & (!g2902) & (!g4401)) + ((!g2854) & (g2881) & (!g2863) & (!g2902) & (g4401)) + ((!g2854) & (g2881) & (g2863) & (!g2902) & (!g4401)) + ((!g2854) & (g2881) & (g2863) & (g2902) & (g4401)) + ((g2854) & (!g2881) & (!g2863) & (!g2902) & (g4401)) + ((g2854) & (!g2881) & (!g2863) & (g2902) & (!g4401)) + ((g2854) & (!g2881) & (g2863) & (!g2902) & (!g4401)) + ((g2854) & (!g2881) & (g2863) & (!g2902) & (g4401)) + ((g2854) & (g2881) & (!g2863) & (!g2902) & (!g4401)) + ((g2854) & (g2881) & (!g2863) & (g2902) & (g4401)) + ((g2854) & (g2881) & (g2863) & (g2902) & (!g4401)) + ((g2854) & (g2881) & (g2863) & (g2902) & (g4401)));
	assign g4454 = (((!g2653) & (!g2674) & (!g4148) & (g5781) & (!g5782) & (!g5783)) + ((!g2653) & (!g2674) & (!g4148) & (g5781) & (!g5782) & (g5783)) + ((!g2653) & (!g2674) & (g4148) & (g5781) & (!g5782) & (!g5783)) + ((!g2653) & (!g2674) & (g4148) & (g5781) & (!g5782) & (g5783)) + ((!g2653) & (g2674) & (!g4148) & (g5781) & (!g5782) & (!g5783)) + ((!g2653) & (g2674) & (!g4148) & (g5781) & (!g5782) & (g5783)) + ((!g2653) & (g2674) & (g4148) & (g5781) & (!g5782) & (!g5783)) + ((!g2653) & (g2674) & (g4148) & (g5781) & (!g5782) & (g5783)) + ((!g2653) & (g2674) & (g4148) & (g5781) & (g5782) & (!g5783)) + ((g2653) & (!g2674) & (!g4148) & (g5781) & (!g5782) & (!g5783)) + ((g2653) & (!g2674) & (!g4148) & (g5781) & (!g5782) & (g5783)) + ((g2653) & (!g2674) & (g4148) & (g5781) & (!g5782) & (!g5783)) + ((g2653) & (!g2674) & (g4148) & (g5781) & (!g5782) & (g5783)) + ((g2653) & (!g2674) & (g4148) & (g5781) & (g5782) & (!g5783)) + ((g2653) & (g2674) & (!g4148) & (g5781) & (!g5782) & (!g5783)) + ((g2653) & (g2674) & (!g4148) & (g5781) & (!g5782) & (g5783)) + ((g2653) & (g2674) & (!g4148) & (g5781) & (g5782) & (!g5783)) + ((g2653) & (g2674) & (g4148) & (g5781) & (!g5782) & (!g5783)) + ((g2653) & (g2674) & (g4148) & (g5781) & (!g5782) & (g5783)) + ((g2653) & (g2674) & (g4148) & (g5781) & (g5782) & (!g5783)));
	assign g4455 = (((g2838) & (g2871)));
	assign g4456 = (((!g2891) & (!g2897) & (!g4454) & (g4455)) + ((!g2891) & (!g2897) & (g4454) & (!g4455)) + ((!g2891) & (!g2897) & (g4454) & (g4455)) + ((!g2891) & (g2897) & (!g4454) & (!g4455)) + ((g2891) & (!g2897) & (!g4454) & (!g4455)) + ((g2891) & (g2897) & (!g4454) & (g4455)) + ((g2891) & (g2897) & (g4454) & (!g4455)) + ((g2891) & (g2897) & (g4454) & (g4455)));
	assign g4457 = (((!g830) & (!g1914) & (!g2239) & (!g4453) & (!g4456)) + ((!g830) & (!g1914) & (!g2239) & (!g4453) & (g4456)) + ((!g830) & (!g1914) & (!g2239) & (g4453) & (!g4456)) + ((!g830) & (!g1914) & (!g2239) & (g4453) & (g4456)) + ((!g830) & (!g1914) & (g2239) & (!g4453) & (!g4456)) + ((!g830) & (!g1914) & (g2239) & (!g4453) & (g4456)) + ((!g830) & (!g1914) & (g2239) & (g4453) & (!g4456)) + ((!g830) & (!g1914) & (g2239) & (g4453) & (g4456)) + ((!g830) & (g1914) & (!g2239) & (!g4453) & (!g4456)) + ((!g830) & (g1914) & (!g2239) & (!g4453) & (g4456)) + ((!g830) & (g1914) & (!g2239) & (g4453) & (!g4456)) + ((!g830) & (g1914) & (!g2239) & (g4453) & (g4456)) + ((!g830) & (g1914) & (g2239) & (!g4453) & (!g4456)) + ((!g830) & (g1914) & (g2239) & (!g4453) & (g4456)) + ((!g830) & (g1914) & (g2239) & (g4453) & (!g4456)) + ((!g830) & (g1914) & (g2239) & (g4453) & (g4456)) + ((g830) & (!g1914) & (!g2239) & (!g4453) & (g4456)) + ((g830) & (!g1914) & (!g2239) & (g4453) & (g4456)) + ((g830) & (!g1914) & (g2239) & (!g4453) & (!g4456)) + ((g830) & (!g1914) & (g2239) & (g4453) & (!g4456)) + ((g830) & (g1914) & (!g2239) & (g4453) & (!g4456)) + ((g830) & (g1914) & (!g2239) & (g4453) & (g4456)) + ((g830) & (g1914) & (g2239) & (!g4453) & (!g4456)) + ((g830) & (g1914) & (g2239) & (!g4453) & (g4456)));
	assign g4458 = (((!g2650) & (!g2684) & (!g3284) & (g3314) & (!g4411)) + ((!g2650) & (!g2684) & (!g3284) & (g3314) & (g4411)) + ((!g2650) & (!g2684) & (g3284) & (!g3314) & (!g4411)) + ((!g2650) & (!g2684) & (g3284) & (g3314) & (g4411)) + ((!g2650) & (g2684) & (!g3284) & (!g3314) & (!g4411)) + ((!g2650) & (g2684) & (!g3284) & (!g3314) & (g4411)) + ((!g2650) & (g2684) & (g3284) & (!g3314) & (g4411)) + ((!g2650) & (g2684) & (g3284) & (g3314) & (!g4411)) + ((g2650) & (!g2684) & (!g3284) & (!g3314) & (!g4411)) + ((g2650) & (!g2684) & (!g3284) & (g3314) & (g4411)) + ((g2650) & (!g2684) & (g3284) & (!g3314) & (!g4411)) + ((g2650) & (!g2684) & (g3284) & (!g3314) & (g4411)) + ((g2650) & (g2684) & (!g3284) & (!g3314) & (g4411)) + ((g2650) & (g2684) & (!g3284) & (g3314) & (!g4411)) + ((g2650) & (g2684) & (g3284) & (g3314) & (!g4411)) + ((g2650) & (g2684) & (g3284) & (g3314) & (g4411)));
	assign g4459 = (((!g3260) & (!g3255) & (!g3305) & (g3297) & (!g4413)) + ((!g3260) & (!g3255) & (!g3305) & (g3297) & (g4413)) + ((!g3260) & (!g3255) & (g3305) & (!g3297) & (!g4413)) + ((!g3260) & (!g3255) & (g3305) & (!g3297) & (g4413)) + ((!g3260) & (g3255) & (!g3305) & (!g3297) & (!g4413)) + ((!g3260) & (g3255) & (!g3305) & (g3297) & (g4413)) + ((!g3260) & (g3255) & (g3305) & (!g3297) & (g4413)) + ((!g3260) & (g3255) & (g3305) & (g3297) & (!g4413)) + ((g3260) & (!g3255) & (!g3305) & (!g3297) & (!g4413)) + ((g3260) & (!g3255) & (!g3305) & (g3297) & (g4413)) + ((g3260) & (!g3255) & (g3305) & (!g3297) & (g4413)) + ((g3260) & (!g3255) & (g3305) & (g3297) & (!g4413)) + ((g3260) & (g3255) & (!g3305) & (!g3297) & (!g4413)) + ((g3260) & (g3255) & (!g3305) & (!g3297) & (g4413)) + ((g3260) & (g3255) & (g3305) & (g3297) & (!g4413)) + ((g3260) & (g3255) & (g3305) & (g3297) & (g4413)));
	assign g4460 = (((!g830) & (!g1914) & (!g2242) & (!g4458) & (!g4459) & (key[198])) + ((!g830) & (!g1914) & (!g2242) & (!g4458) & (g4459) & (key[198])) + ((!g830) & (!g1914) & (!g2242) & (g4458) & (!g4459) & (key[198])) + ((!g830) & (!g1914) & (!g2242) & (g4458) & (g4459) & (key[198])) + ((!g830) & (!g1914) & (g2242) & (!g4458) & (!g4459) & (key[198])) + ((!g830) & (!g1914) & (g2242) & (!g4458) & (g4459) & (key[198])) + ((!g830) & (!g1914) & (g2242) & (g4458) & (!g4459) & (key[198])) + ((!g830) & (!g1914) & (g2242) & (g4458) & (g4459) & (key[198])) + ((!g830) & (g1914) & (!g2242) & (!g4458) & (!g4459) & (key[198])) + ((!g830) & (g1914) & (!g2242) & (!g4458) & (g4459) & (key[198])) + ((!g830) & (g1914) & (!g2242) & (g4458) & (!g4459) & (key[198])) + ((!g830) & (g1914) & (!g2242) & (g4458) & (g4459) & (key[198])) + ((!g830) & (g1914) & (g2242) & (!g4458) & (!g4459) & (key[198])) + ((!g830) & (g1914) & (g2242) & (!g4458) & (g4459) & (key[198])) + ((!g830) & (g1914) & (g2242) & (g4458) & (!g4459) & (key[198])) + ((!g830) & (g1914) & (g2242) & (g4458) & (g4459) & (key[198])) + ((g830) & (!g1914) & (!g2242) & (!g4458) & (g4459) & (!key[198])) + ((g830) & (!g1914) & (!g2242) & (!g4458) & (g4459) & (key[198])) + ((g830) & (!g1914) & (!g2242) & (g4458) & (g4459) & (!key[198])) + ((g830) & (!g1914) & (!g2242) & (g4458) & (g4459) & (key[198])) + ((g830) & (!g1914) & (g2242) & (!g4458) & (!g4459) & (!key[198])) + ((g830) & (!g1914) & (g2242) & (!g4458) & (!g4459) & (key[198])) + ((g830) & (!g1914) & (g2242) & (g4458) & (!g4459) & (!key[198])) + ((g830) & (!g1914) & (g2242) & (g4458) & (!g4459) & (key[198])) + ((g830) & (g1914) & (!g2242) & (g4458) & (!g4459) & (!key[198])) + ((g830) & (g1914) & (!g2242) & (g4458) & (!g4459) & (key[198])) + ((g830) & (g1914) & (!g2242) & (g4458) & (g4459) & (!key[198])) + ((g830) & (g1914) & (!g2242) & (g4458) & (g4459) & (key[198])) + ((g830) & (g1914) & (g2242) & (!g4458) & (!g4459) & (!key[198])) + ((g830) & (g1914) & (g2242) & (!g4458) & (!g4459) & (key[198])) + ((g830) & (g1914) & (g2242) & (!g4458) & (g4459) & (!key[198])) + ((g830) & (g1914) & (g2242) & (!g4458) & (g4459) & (key[198])));
	assign g4461 = (((!g4392) & (!g3330) & (!g3342) & (!g3370) & (g3372)) + ((!g4392) & (!g3330) & (!g3342) & (g3370) & (!g3372)) + ((!g4392) & (!g3330) & (g3342) & (!g3370) & (g3372)) + ((!g4392) & (!g3330) & (g3342) & (g3370) & (!g3372)) + ((!g4392) & (g3330) & (!g3342) & (!g3370) & (g3372)) + ((!g4392) & (g3330) & (!g3342) & (g3370) & (!g3372)) + ((!g4392) & (g3330) & (g3342) & (!g3370) & (!g3372)) + ((!g4392) & (g3330) & (g3342) & (g3370) & (g3372)) + ((g4392) & (!g3330) & (!g3342) & (!g3370) & (g3372)) + ((g4392) & (!g3330) & (!g3342) & (g3370) & (!g3372)) + ((g4392) & (!g3330) & (g3342) & (!g3370) & (!g3372)) + ((g4392) & (!g3330) & (g3342) & (g3370) & (g3372)) + ((g4392) & (g3330) & (!g3342) & (!g3370) & (!g3372)) + ((g4392) & (g3330) & (!g3342) & (g3370) & (g3372)) + ((g4392) & (g3330) & (g3342) & (!g3370) & (!g3372)) + ((g4392) & (g3330) & (g3342) & (g3370) & (g3372)));
	assign g4462 = (((!g2424) & (!g2516) & (!g4393) & (!g3095) & (g3131)) + ((!g2424) & (!g2516) & (!g4393) & (g3095) & (g3131)) + ((!g2424) & (!g2516) & (g4393) & (!g3095) & (g3131)) + ((!g2424) & (!g2516) & (g4393) & (g3095) & (!g3131)) + ((!g2424) & (g2516) & (!g4393) & (!g3095) & (!g3131)) + ((!g2424) & (g2516) & (!g4393) & (g3095) & (!g3131)) + ((!g2424) & (g2516) & (g4393) & (!g3095) & (!g3131)) + ((!g2424) & (g2516) & (g4393) & (g3095) & (g3131)) + ((g2424) & (!g2516) & (!g4393) & (!g3095) & (g3131)) + ((g2424) & (!g2516) & (!g4393) & (g3095) & (!g3131)) + ((g2424) & (!g2516) & (g4393) & (!g3095) & (!g3131)) + ((g2424) & (!g2516) & (g4393) & (g3095) & (!g3131)) + ((g2424) & (g2516) & (!g4393) & (!g3095) & (!g3131)) + ((g2424) & (g2516) & (!g4393) & (g3095) & (g3131)) + ((g2424) & (g2516) & (g4393) & (!g3095) & (g3131)) + ((g2424) & (g2516) & (g4393) & (g3095) & (g3131)));
	assign g4463 = (((!g830) & (!g1914) & (!g2247) & (!g4461) & (!g4462) & (key[134])) + ((!g830) & (!g1914) & (!g2247) & (!g4461) & (g4462) & (key[134])) + ((!g830) & (!g1914) & (!g2247) & (g4461) & (!g4462) & (key[134])) + ((!g830) & (!g1914) & (!g2247) & (g4461) & (g4462) & (key[134])) + ((!g830) & (!g1914) & (g2247) & (!g4461) & (!g4462) & (key[134])) + ((!g830) & (!g1914) & (g2247) & (!g4461) & (g4462) & (key[134])) + ((!g830) & (!g1914) & (g2247) & (g4461) & (!g4462) & (key[134])) + ((!g830) & (!g1914) & (g2247) & (g4461) & (g4462) & (key[134])) + ((!g830) & (g1914) & (!g2247) & (!g4461) & (!g4462) & (key[134])) + ((!g830) & (g1914) & (!g2247) & (!g4461) & (g4462) & (key[134])) + ((!g830) & (g1914) & (!g2247) & (g4461) & (!g4462) & (key[134])) + ((!g830) & (g1914) & (!g2247) & (g4461) & (g4462) & (key[134])) + ((!g830) & (g1914) & (g2247) & (!g4461) & (!g4462) & (key[134])) + ((!g830) & (g1914) & (g2247) & (!g4461) & (g4462) & (key[134])) + ((!g830) & (g1914) & (g2247) & (g4461) & (!g4462) & (key[134])) + ((!g830) & (g1914) & (g2247) & (g4461) & (g4462) & (key[134])) + ((g830) & (!g1914) & (!g2247) & (!g4461) & (g4462) & (!key[134])) + ((g830) & (!g1914) & (!g2247) & (!g4461) & (g4462) & (key[134])) + ((g830) & (!g1914) & (!g2247) & (g4461) & (g4462) & (!key[134])) + ((g830) & (!g1914) & (!g2247) & (g4461) & (g4462) & (key[134])) + ((g830) & (!g1914) & (g2247) & (!g4461) & (!g4462) & (!key[134])) + ((g830) & (!g1914) & (g2247) & (!g4461) & (!g4462) & (key[134])) + ((g830) & (!g1914) & (g2247) & (g4461) & (!g4462) & (!key[134])) + ((g830) & (!g1914) & (g2247) & (g4461) & (!g4462) & (key[134])) + ((g830) & (g1914) & (!g2247) & (g4461) & (!g4462) & (!key[134])) + ((g830) & (g1914) & (!g2247) & (g4461) & (!g4462) & (key[134])) + ((g830) & (g1914) & (!g2247) & (g4461) & (g4462) & (!key[134])) + ((g830) & (g1914) & (!g2247) & (g4461) & (g4462) & (key[134])) + ((g830) & (g1914) & (g2247) & (!g4461) & (!g4462) & (!key[134])) + ((g830) & (g1914) & (g2247) & (!g4461) & (!g4462) & (key[134])) + ((g830) & (g1914) & (g2247) & (!g4461) & (g4462) & (!key[134])) + ((g830) & (g1914) & (g2247) & (!g4461) & (g4462) & (key[134])));
	assign g4464 = (((!g3260) & (!g3240) & (!g3305) & (g3303) & (!g4403)) + ((!g3260) & (!g3240) & (!g3305) & (g3303) & (g4403)) + ((!g3260) & (!g3240) & (g3305) & (!g3303) & (!g4403)) + ((!g3260) & (!g3240) & (g3305) & (!g3303) & (g4403)) + ((!g3260) & (g3240) & (!g3305) & (!g3303) & (!g4403)) + ((!g3260) & (g3240) & (!g3305) & (g3303) & (g4403)) + ((!g3260) & (g3240) & (g3305) & (!g3303) & (g4403)) + ((!g3260) & (g3240) & (g3305) & (g3303) & (!g4403)) + ((g3260) & (!g3240) & (!g3305) & (!g3303) & (!g4403)) + ((g3260) & (!g3240) & (!g3305) & (g3303) & (g4403)) + ((g3260) & (!g3240) & (g3305) & (!g3303) & (g4403)) + ((g3260) & (!g3240) & (g3305) & (g3303) & (!g4403)) + ((g3260) & (g3240) & (!g3305) & (!g3303) & (!g4403)) + ((g3260) & (g3240) & (!g3305) & (!g3303) & (g4403)) + ((g3260) & (g3240) & (g3305) & (g3303) & (!g4403)) + ((g3260) & (g3240) & (g3305) & (g3303) & (g4403)));
	assign g4465 = (((!g2648) & (!g2679) & (!g3284) & (g3314) & (!g4405)) + ((!g2648) & (!g2679) & (!g3284) & (g3314) & (g4405)) + ((!g2648) & (!g2679) & (g3284) & (!g3314) & (!g4405)) + ((!g2648) & (!g2679) & (g3284) & (g3314) & (g4405)) + ((!g2648) & (g2679) & (!g3284) & (!g3314) & (!g4405)) + ((!g2648) & (g2679) & (!g3284) & (!g3314) & (g4405)) + ((!g2648) & (g2679) & (g3284) & (!g3314) & (g4405)) + ((!g2648) & (g2679) & (g3284) & (g3314) & (!g4405)) + ((g2648) & (!g2679) & (!g3284) & (!g3314) & (!g4405)) + ((g2648) & (!g2679) & (!g3284) & (g3314) & (g4405)) + ((g2648) & (!g2679) & (g3284) & (!g3314) & (!g4405)) + ((g2648) & (!g2679) & (g3284) & (!g3314) & (g4405)) + ((g2648) & (g2679) & (!g3284) & (!g3314) & (g4405)) + ((g2648) & (g2679) & (!g3284) & (g3314) & (!g4405)) + ((g2648) & (g2679) & (g3284) & (g3314) & (!g4405)) + ((g2648) & (g2679) & (g3284) & (g3314) & (g4405)));
	assign g4466 = (((!g830) & (!g1914) & (!g2250) & (!g4464) & (!g4465) & (nonce[38])) + ((!g830) & (!g1914) & (!g2250) & (!g4464) & (g4465) & (nonce[38])) + ((!g830) & (!g1914) & (!g2250) & (g4464) & (!g4465) & (nonce[38])) + ((!g830) & (!g1914) & (!g2250) & (g4464) & (g4465) & (nonce[38])) + ((!g830) & (!g1914) & (g2250) & (!g4464) & (!g4465) & (nonce[38])) + ((!g830) & (!g1914) & (g2250) & (!g4464) & (g4465) & (nonce[38])) + ((!g830) & (!g1914) & (g2250) & (g4464) & (!g4465) & (nonce[38])) + ((!g830) & (!g1914) & (g2250) & (g4464) & (g4465) & (nonce[38])) + ((!g830) & (g1914) & (!g2250) & (!g4464) & (!g4465) & (nonce[38])) + ((!g830) & (g1914) & (!g2250) & (!g4464) & (g4465) & (nonce[38])) + ((!g830) & (g1914) & (!g2250) & (g4464) & (!g4465) & (nonce[38])) + ((!g830) & (g1914) & (!g2250) & (g4464) & (g4465) & (nonce[38])) + ((!g830) & (g1914) & (g2250) & (!g4464) & (!g4465) & (nonce[38])) + ((!g830) & (g1914) & (g2250) & (!g4464) & (g4465) & (nonce[38])) + ((!g830) & (g1914) & (g2250) & (g4464) & (!g4465) & (nonce[38])) + ((!g830) & (g1914) & (g2250) & (g4464) & (g4465) & (nonce[38])) + ((g830) & (!g1914) & (!g2250) & (!g4464) & (g4465) & (!nonce[38])) + ((g830) & (!g1914) & (!g2250) & (!g4464) & (g4465) & (nonce[38])) + ((g830) & (!g1914) & (!g2250) & (g4464) & (g4465) & (!nonce[38])) + ((g830) & (!g1914) & (!g2250) & (g4464) & (g4465) & (nonce[38])) + ((g830) & (!g1914) & (g2250) & (!g4464) & (!g4465) & (!nonce[38])) + ((g830) & (!g1914) & (g2250) & (!g4464) & (!g4465) & (nonce[38])) + ((g830) & (!g1914) & (g2250) & (g4464) & (!g4465) & (!nonce[38])) + ((g830) & (!g1914) & (g2250) & (g4464) & (!g4465) & (nonce[38])) + ((g830) & (g1914) & (!g2250) & (g4464) & (!g4465) & (!nonce[38])) + ((g830) & (g1914) & (!g2250) & (g4464) & (!g4465) & (nonce[38])) + ((g830) & (g1914) & (!g2250) & (g4464) & (g4465) & (!nonce[38])) + ((g830) & (g1914) & (!g2250) & (g4464) & (g4465) & (nonce[38])) + ((g830) & (g1914) & (g2250) & (!g4464) & (!g4465) & (!nonce[38])) + ((g830) & (g1914) & (g2250) & (!g4464) & (!g4465) & (nonce[38])) + ((g830) & (g1914) & (g2250) & (!g4464) & (g4465) & (!nonce[38])) + ((g830) & (g1914) & (g2250) & (!g4464) & (g4465) & (nonce[38])));
	assign g4467 = (((!g2868) & (!g2889) & (!g2871) & (g2897) & (!g4416)) + ((!g2868) & (!g2889) & (!g2871) & (g2897) & (g4416)) + ((!g2868) & (!g2889) & (g2871) & (!g2897) & (g4416)) + ((!g2868) & (!g2889) & (g2871) & (g2897) & (!g4416)) + ((!g2868) & (g2889) & (!g2871) & (!g2897) & (!g4416)) + ((!g2868) & (g2889) & (!g2871) & (!g2897) & (g4416)) + ((!g2868) & (g2889) & (g2871) & (!g2897) & (!g4416)) + ((!g2868) & (g2889) & (g2871) & (g2897) & (g4416)) + ((g2868) & (!g2889) & (!g2871) & (!g2897) & (g4416)) + ((g2868) & (!g2889) & (!g2871) & (g2897) & (!g4416)) + ((g2868) & (!g2889) & (g2871) & (!g2897) & (!g4416)) + ((g2868) & (!g2889) & (g2871) & (!g2897) & (g4416)) + ((g2868) & (g2889) & (!g2871) & (!g2897) & (!g4416)) + ((g2868) & (g2889) & (!g2871) & (g2897) & (g4416)) + ((g2868) & (g2889) & (g2871) & (g2897) & (!g4416)) + ((g2868) & (g2889) & (g2871) & (g2897) & (g4416)));
	assign g4468 = (((!g2661) & (!g2669) & (!g4166) & (g5784) & (!g5785) & (!g5786)) + ((!g2661) & (!g2669) & (!g4166) & (g5784) & (!g5785) & (g5786)) + ((!g2661) & (!g2669) & (g4166) & (g5784) & (!g5785) & (!g5786)) + ((!g2661) & (!g2669) & (g4166) & (g5784) & (!g5785) & (g5786)) + ((!g2661) & (g2669) & (!g4166) & (g5784) & (!g5785) & (!g5786)) + ((!g2661) & (g2669) & (!g4166) & (g5784) & (!g5785) & (g5786)) + ((!g2661) & (g2669) & (g4166) & (g5784) & (!g5785) & (!g5786)) + ((!g2661) & (g2669) & (g4166) & (g5784) & (!g5785) & (g5786)) + ((!g2661) & (g2669) & (g4166) & (g5784) & (g5785) & (!g5786)) + ((g2661) & (!g2669) & (!g4166) & (g5784) & (!g5785) & (!g5786)) + ((g2661) & (!g2669) & (!g4166) & (g5784) & (!g5785) & (g5786)) + ((g2661) & (!g2669) & (g4166) & (g5784) & (!g5785) & (!g5786)) + ((g2661) & (!g2669) & (g4166) & (g5784) & (!g5785) & (g5786)) + ((g2661) & (!g2669) & (g4166) & (g5784) & (g5785) & (!g5786)) + ((g2661) & (g2669) & (!g4166) & (g5784) & (!g5785) & (!g5786)) + ((g2661) & (g2669) & (!g4166) & (g5784) & (!g5785) & (g5786)) + ((g2661) & (g2669) & (!g4166) & (g5784) & (g5785) & (!g5786)) + ((g2661) & (g2669) & (g4166) & (g5784) & (!g5785) & (!g5786)) + ((g2661) & (g2669) & (g4166) & (g5784) & (!g5785) & (g5786)) + ((g2661) & (g2669) & (g4166) & (g5784) & (g5785) & (!g5786)));
	assign g4469 = (((g2851) & (g2863)));
	assign g4470 = (((!g2900) & (!g2902) & (!g4468) & (g4469)) + ((!g2900) & (!g2902) & (g4468) & (!g4469)) + ((!g2900) & (!g2902) & (g4468) & (g4469)) + ((!g2900) & (g2902) & (!g4468) & (!g4469)) + ((g2900) & (!g2902) & (!g4468) & (!g4469)) + ((g2900) & (g2902) & (!g4468) & (g4469)) + ((g2900) & (g2902) & (g4468) & (!g4469)) + ((g2900) & (g2902) & (g4468) & (g4469)));
	assign g4471 = (((!g830) & (!g1914) & (!g2253) & (!g4467) & (!g4470)) + ((!g830) & (!g1914) & (!g2253) & (!g4467) & (g4470)) + ((!g830) & (!g1914) & (!g2253) & (g4467) & (!g4470)) + ((!g830) & (!g1914) & (!g2253) & (g4467) & (g4470)) + ((!g830) & (!g1914) & (g2253) & (!g4467) & (!g4470)) + ((!g830) & (!g1914) & (g2253) & (!g4467) & (g4470)) + ((!g830) & (!g1914) & (g2253) & (g4467) & (!g4470)) + ((!g830) & (!g1914) & (g2253) & (g4467) & (g4470)) + ((!g830) & (g1914) & (!g2253) & (!g4467) & (!g4470)) + ((!g830) & (g1914) & (!g2253) & (!g4467) & (g4470)) + ((!g830) & (g1914) & (!g2253) & (g4467) & (!g4470)) + ((!g830) & (g1914) & (!g2253) & (g4467) & (g4470)) + ((!g830) & (g1914) & (g2253) & (!g4467) & (!g4470)) + ((!g830) & (g1914) & (g2253) & (!g4467) & (g4470)) + ((!g830) & (g1914) & (g2253) & (g4467) & (!g4470)) + ((!g830) & (g1914) & (g2253) & (g4467) & (g4470)) + ((g830) & (!g1914) & (!g2253) & (!g4467) & (g4470)) + ((g830) & (!g1914) & (!g2253) & (g4467) & (g4470)) + ((g830) & (!g1914) & (g2253) & (!g4467) & (!g4470)) + ((g830) & (!g1914) & (g2253) & (g4467) & (!g4470)) + ((g830) & (g1914) & (!g2253) & (g4467) & (!g4470)) + ((g830) & (g1914) & (!g2253) & (g4467) & (g4470)) + ((g830) & (g1914) & (g2253) & (!g4467) & (!g4470)) + ((g830) & (g1914) & (g2253) & (!g4467) & (g4470)));
	assign g4472 = (((!g3505) & (!g3506)));
	assign g4473 = (((g1914) & (!g1199) & (!g4472) & (!g2434)) + ((g1914) & (!g1199) & (g4472) & (g2434)) + ((g1914) & (g1199) & (!g4472) & (g2434)) + ((g1914) & (g1199) & (g4472) & (!g2434)));
	assign g4474 = (((!g3523) & (!g3524)));
	assign g4475 = (((!g1914) & (!g2450) & (!g2497) & (!g4474)) + ((!g1914) & (!g2450) & (g2497) & (g4474)) + ((!g1914) & (g2450) & (!g2497) & (g4474)) + ((!g1914) & (g2450) & (g2497) & (!g4474)));
	assign g4476 = (((!g830) & (!g2256) & (!g4473) & (!g4475) & (key[52])) + ((!g830) & (!g2256) & (!g4473) & (g4475) & (key[52])) + ((!g830) & (!g2256) & (g4473) & (!g4475) & (key[52])) + ((!g830) & (!g2256) & (g4473) & (g4475) & (key[52])) + ((!g830) & (g2256) & (!g4473) & (!g4475) & (key[52])) + ((!g830) & (g2256) & (!g4473) & (g4475) & (key[52])) + ((!g830) & (g2256) & (g4473) & (!g4475) & (key[52])) + ((!g830) & (g2256) & (g4473) & (g4475) & (key[52])) + ((g830) & (!g2256) & (!g4473) & (g4475) & (!key[52])) + ((g830) & (!g2256) & (!g4473) & (g4475) & (key[52])) + ((g830) & (!g2256) & (g4473) & (!g4475) & (!key[52])) + ((g830) & (!g2256) & (g4473) & (!g4475) & (key[52])) + ((g830) & (!g2256) & (g4473) & (g4475) & (!key[52])) + ((g830) & (!g2256) & (g4473) & (g4475) & (key[52])) + ((g830) & (g2256) & (!g4473) & (!g4475) & (!key[52])) + ((g830) & (g2256) & (!g4473) & (!g4475) & (key[52])));
	assign g4477 = (((!g1953) & (!g1955) & (!g2233) & (g2267) & (!g4421)) + ((!g1953) & (!g1955) & (!g2233) & (g2267) & (g4421)) + ((!g1953) & (!g1955) & (g2233) & (!g2267) & (!g4421)) + ((!g1953) & (!g1955) & (g2233) & (g2267) & (g4421)) + ((!g1953) & (g1955) & (!g2233) & (!g2267) & (!g4421)) + ((!g1953) & (g1955) & (!g2233) & (!g2267) & (g4421)) + ((!g1953) & (g1955) & (g2233) & (!g2267) & (g4421)) + ((!g1953) & (g1955) & (g2233) & (g2267) & (!g4421)) + ((g1953) & (!g1955) & (!g2233) & (!g2267) & (!g4421)) + ((g1953) & (!g1955) & (!g2233) & (g2267) & (g4421)) + ((g1953) & (!g1955) & (g2233) & (!g2267) & (!g4421)) + ((g1953) & (!g1955) & (g2233) & (!g2267) & (g4421)) + ((g1953) & (g1955) & (!g2233) & (!g2267) & (g4421)) + ((g1953) & (g1955) & (!g2233) & (g2267) & (!g4421)) + ((g1953) & (g1955) & (g2233) & (g2267) & (!g4421)) + ((g1953) & (g1955) & (g2233) & (g2267) & (g4421)));
	assign g4478 = (((!g2572) & (!g2595) & (!g3767)) + ((!g2572) & (g2595) & (g3767)) + ((g2572) & (!g2595) & (g3767)) + ((g2572) & (g2595) & (!g3767)));
	assign g4479 = (((!g830) & (!g1914) & (!g2257) & (!g4477) & (!g4478) & (key[84])) + ((!g830) & (!g1914) & (!g2257) & (!g4477) & (g4478) & (key[84])) + ((!g830) & (!g1914) & (!g2257) & (g4477) & (!g4478) & (key[84])) + ((!g830) & (!g1914) & (!g2257) & (g4477) & (g4478) & (key[84])) + ((!g830) & (!g1914) & (g2257) & (!g4477) & (!g4478) & (key[84])) + ((!g830) & (!g1914) & (g2257) & (!g4477) & (g4478) & (key[84])) + ((!g830) & (!g1914) & (g2257) & (g4477) & (!g4478) & (key[84])) + ((!g830) & (!g1914) & (g2257) & (g4477) & (g4478) & (key[84])) + ((!g830) & (g1914) & (!g2257) & (!g4477) & (!g4478) & (key[84])) + ((!g830) & (g1914) & (!g2257) & (!g4477) & (g4478) & (key[84])) + ((!g830) & (g1914) & (!g2257) & (g4477) & (!g4478) & (key[84])) + ((!g830) & (g1914) & (!g2257) & (g4477) & (g4478) & (key[84])) + ((!g830) & (g1914) & (g2257) & (!g4477) & (!g4478) & (key[84])) + ((!g830) & (g1914) & (g2257) & (!g4477) & (g4478) & (key[84])) + ((!g830) & (g1914) & (g2257) & (g4477) & (!g4478) & (key[84])) + ((!g830) & (g1914) & (g2257) & (g4477) & (g4478) & (key[84])) + ((g830) & (!g1914) & (!g2257) & (!g4477) & (g4478) & (!key[84])) + ((g830) & (!g1914) & (!g2257) & (!g4477) & (g4478) & (key[84])) + ((g830) & (!g1914) & (!g2257) & (g4477) & (g4478) & (!key[84])) + ((g830) & (!g1914) & (!g2257) & (g4477) & (g4478) & (key[84])) + ((g830) & (!g1914) & (g2257) & (!g4477) & (!g4478) & (!key[84])) + ((g830) & (!g1914) & (g2257) & (!g4477) & (!g4478) & (key[84])) + ((g830) & (!g1914) & (g2257) & (g4477) & (!g4478) & (!key[84])) + ((g830) & (!g1914) & (g2257) & (g4477) & (!g4478) & (key[84])) + ((g830) & (g1914) & (!g2257) & (g4477) & (!g4478) & (!key[84])) + ((g830) & (g1914) & (!g2257) & (g4477) & (!g4478) & (key[84])) + ((g830) & (g1914) & (!g2257) & (g4477) & (g4478) & (!key[84])) + ((g830) & (g1914) & (!g2257) & (g4477) & (g4478) & (key[84])) + ((g830) & (g1914) & (g2257) & (!g4477) & (!g4478) & (!key[84])) + ((g830) & (g1914) & (g2257) & (!g4477) & (!g4478) & (key[84])) + ((g830) & (g1914) & (g2257) & (!g4477) & (g4478) & (!key[84])) + ((g830) & (g1914) & (g2257) & (!g4477) & (g4478) & (key[84])));
	assign g4480 = (((!g3415) & (g3416)) + ((g3415) & (!g3416)) + ((g3415) & (g3416)));
	assign g4481 = (((!g3398) & (g3399)) + ((g3398) & (!g3399)) + ((g3398) & (g3399)));
	assign g8303 = (((!g5560) & (g5599) & (!g4482)) + ((!g5560) & (g5599) & (g4482)) + ((g5560) & (!g5599) & (g4482)) + ((g5560) & (g5599) & (g4482)));
	assign g4483 = (((!g830) & (!g2262) & (!g6724) & (g4482)) + ((!g830) & (!g2262) & (g6724) & (g4482)) + ((!g830) & (g2262) & (!g6724) & (g4482)) + ((!g830) & (g2262) & (g6724) & (g4482)) + ((g830) & (!g2262) & (g6724) & (!g4482)) + ((g830) & (!g2262) & (g6724) & (g4482)) + ((g830) & (g2262) & (!g6724) & (!g4482)) + ((g830) & (g2262) & (!g6724) & (g4482)));
	assign g4484 = (((!g3473) & (!g2589) & (!g2595)) + ((!g3473) & (g2589) & (g2595)) + ((g3473) & (!g2589) & (g2595)) + ((g3473) & (g2589) & (!g2595)));
	assign g4485 = (((!g1991) & (!g1993) & (!g2217) & (g2277) & (!g4429)) + ((!g1991) & (!g1993) & (!g2217) & (g2277) & (g4429)) + ((!g1991) & (!g1993) & (g2217) & (!g2277) & (!g4429)) + ((!g1991) & (!g1993) & (g2217) & (g2277) & (g4429)) + ((!g1991) & (g1993) & (!g2217) & (!g2277) & (!g4429)) + ((!g1991) & (g1993) & (!g2217) & (!g2277) & (g4429)) + ((!g1991) & (g1993) & (g2217) & (!g2277) & (g4429)) + ((!g1991) & (g1993) & (g2217) & (g2277) & (!g4429)) + ((g1991) & (!g1993) & (!g2217) & (!g2277) & (!g4429)) + ((g1991) & (!g1993) & (!g2217) & (g2277) & (g4429)) + ((g1991) & (!g1993) & (g2217) & (!g2277) & (!g4429)) + ((g1991) & (!g1993) & (g2217) & (!g2277) & (g4429)) + ((g1991) & (g1993) & (!g2217) & (!g2277) & (g4429)) + ((g1991) & (g1993) & (!g2217) & (g2277) & (!g4429)) + ((g1991) & (g1993) & (g2217) & (g2277) & (!g4429)) + ((g1991) & (g1993) & (g2217) & (g2277) & (g4429)));
	assign g4486 = (((!g830) & (!g1914) & (!g2263) & (!g4484) & (!g4485) & (key[180])) + ((!g830) & (!g1914) & (!g2263) & (!g4484) & (g4485) & (key[180])) + ((!g830) & (!g1914) & (!g2263) & (g4484) & (!g4485) & (key[180])) + ((!g830) & (!g1914) & (!g2263) & (g4484) & (g4485) & (key[180])) + ((!g830) & (!g1914) & (g2263) & (!g4484) & (!g4485) & (key[180])) + ((!g830) & (!g1914) & (g2263) & (!g4484) & (g4485) & (key[180])) + ((!g830) & (!g1914) & (g2263) & (g4484) & (!g4485) & (key[180])) + ((!g830) & (!g1914) & (g2263) & (g4484) & (g4485) & (key[180])) + ((!g830) & (g1914) & (!g2263) & (!g4484) & (!g4485) & (key[180])) + ((!g830) & (g1914) & (!g2263) & (!g4484) & (g4485) & (key[180])) + ((!g830) & (g1914) & (!g2263) & (g4484) & (!g4485) & (key[180])) + ((!g830) & (g1914) & (!g2263) & (g4484) & (g4485) & (key[180])) + ((!g830) & (g1914) & (g2263) & (!g4484) & (!g4485) & (key[180])) + ((!g830) & (g1914) & (g2263) & (!g4484) & (g4485) & (key[180])) + ((!g830) & (g1914) & (g2263) & (g4484) & (!g4485) & (key[180])) + ((!g830) & (g1914) & (g2263) & (g4484) & (g4485) & (key[180])) + ((g830) & (!g1914) & (!g2263) & (!g4484) & (g4485) & (!key[180])) + ((g830) & (!g1914) & (!g2263) & (!g4484) & (g4485) & (key[180])) + ((g830) & (!g1914) & (!g2263) & (g4484) & (g4485) & (!key[180])) + ((g830) & (!g1914) & (!g2263) & (g4484) & (g4485) & (key[180])) + ((g830) & (!g1914) & (g2263) & (!g4484) & (!g4485) & (!key[180])) + ((g830) & (!g1914) & (g2263) & (!g4484) & (!g4485) & (key[180])) + ((g830) & (!g1914) & (g2263) & (g4484) & (!g4485) & (!key[180])) + ((g830) & (!g1914) & (g2263) & (g4484) & (!g4485) & (key[180])) + ((g830) & (g1914) & (!g2263) & (g4484) & (!g4485) & (!key[180])) + ((g830) & (g1914) & (!g2263) & (g4484) & (!g4485) & (key[180])) + ((g830) & (g1914) & (!g2263) & (g4484) & (g4485) & (!key[180])) + ((g830) & (g1914) & (!g2263) & (g4484) & (g4485) & (key[180])) + ((g830) & (g1914) & (g2263) & (!g4484) & (!g4485) & (!key[180])) + ((g830) & (g1914) & (g2263) & (!g4484) & (!g4485) & (key[180])) + ((g830) & (g1914) & (g2263) & (!g4484) & (g4485) & (!key[180])) + ((g830) & (g1914) & (g2263) & (!g4484) & (g4485) & (key[180])));
	assign g4487 = (((!g3116) & (g3139)) + ((g3116) & (!g3139)));
	assign g4488 = (((!g3041) & (!g3086) & (g3064) & (!g4336) & (g3090) & (g4487)) + ((!g3041) & (g3086) & (!g3064) & (!g4336) & (g3090) & (g4487)) + ((!g3041) & (g3086) & (!g3064) & (g4336) & (g3090) & (g4487)) + ((!g3041) & (g3086) & (g3064) & (!g4336) & (!g3090) & (g4487)) + ((!g3041) & (g3086) & (g3064) & (!g4336) & (g3090) & (g4487)) + ((!g3041) & (g3086) & (g3064) & (g4336) & (g3090) & (g4487)) + ((g3041) & (!g3086) & (!g3064) & (!g4336) & (g3090) & (g4487)) + ((g3041) & (!g3086) & (g3064) & (!g4336) & (g3090) & (g4487)) + ((g3041) & (!g3086) & (g3064) & (g4336) & (g3090) & (g4487)) + ((g3041) & (g3086) & (!g3064) & (!g4336) & (!g3090) & (g4487)) + ((g3041) & (g3086) & (!g3064) & (!g4336) & (g3090) & (g4487)) + ((g3041) & (g3086) & (!g3064) & (g4336) & (g3090) & (g4487)) + ((g3041) & (g3086) & (g3064) & (!g4336) & (!g3090) & (g4487)) + ((g3041) & (g3086) & (g3064) & (!g4336) & (g3090) & (g4487)) + ((g3041) & (g3086) & (g3064) & (g4336) & (!g3090) & (g4487)) + ((g3041) & (g3086) & (g3064) & (g4336) & (g3090) & (g4487)));
	assign g4489 = (((g3116) & (g3139)));
	assign g4490 = (((!g3161) & (!g4488) & (!g4489) & (g3165)) + ((!g3161) & (!g4488) & (g4489) & (!g3165)) + ((!g3161) & (g4488) & (!g4489) & (!g3165)) + ((!g3161) & (g4488) & (g4489) & (!g3165)) + ((g3161) & (!g4488) & (!g4489) & (!g3165)) + ((g3161) & (!g4488) & (g4489) & (g3165)) + ((g3161) & (g4488) & (!g4489) & (g3165)) + ((g3161) & (g4488) & (g4489) & (g3165)));
	assign g4491 = (((!g2262) & (g2893)) + ((g2262) & (!g2893)));
	assign g4492 = (((!g2180) & (!g2212) & (g2816) & (g2848) & (g4324) & (g4491)) + ((!g2180) & (g2212) & (!g2816) & (g2848) & (!g4324) & (g4491)) + ((!g2180) & (g2212) & (!g2816) & (g2848) & (g4324) & (g4491)) + ((!g2180) & (g2212) & (g2816) & (!g2848) & (g4324) & (g4491)) + ((!g2180) & (g2212) & (g2816) & (g2848) & (!g4324) & (g4491)) + ((!g2180) & (g2212) & (g2816) & (g2848) & (g4324) & (g4491)) + ((g2180) & (!g2212) & (!g2816) & (g2848) & (g4324) & (g4491)) + ((g2180) & (!g2212) & (g2816) & (g2848) & (!g4324) & (g4491)) + ((g2180) & (!g2212) & (g2816) & (g2848) & (g4324) & (g4491)) + ((g2180) & (g2212) & (!g2816) & (!g2848) & (g4324) & (g4491)) + ((g2180) & (g2212) & (!g2816) & (g2848) & (!g4324) & (g4491)) + ((g2180) & (g2212) & (!g2816) & (g2848) & (g4324) & (g4491)) + ((g2180) & (g2212) & (g2816) & (!g2848) & (!g4324) & (g4491)) + ((g2180) & (g2212) & (g2816) & (!g2848) & (g4324) & (g4491)) + ((g2180) & (g2212) & (g2816) & (g2848) & (!g4324) & (g4491)) + ((g2180) & (g2212) & (g2816) & (g2848) & (g4324) & (g4491)));
	assign g4493 = (((g2262) & (g2893)));
	assign g4494 = (((!g2298) & (!g2938) & (!g4492) & (g4493)) + ((!g2298) & (!g2938) & (g4492) & (!g4493)) + ((!g2298) & (!g2938) & (g4492) & (g4493)) + ((!g2298) & (g2938) & (!g4492) & (!g4493)) + ((g2298) & (!g2938) & (!g4492) & (!g4493)) + ((g2298) & (g2938) & (!g4492) & (g4493)) + ((g2298) & (g2938) & (g4492) & (!g4493)) + ((g2298) & (g2938) & (g4492) & (g4493)));
	assign g4495 = (((!g2256) & (!g2295) & (!g2887) & (g2956) & (!g4436) & (!g4437)) + ((!g2256) & (!g2295) & (!g2887) & (g2956) & (!g4436) & (g4437)) + ((!g2256) & (!g2295) & (!g2887) & (g2956) & (g4436) & (!g4437)) + ((!g2256) & (!g2295) & (!g2887) & (g2956) & (g4436) & (g4437)) + ((!g2256) & (!g2295) & (g2887) & (!g2956) & (!g4436) & (g4437)) + ((!g2256) & (!g2295) & (g2887) & (!g2956) & (g4436) & (!g4437)) + ((!g2256) & (!g2295) & (g2887) & (!g2956) & (g4436) & (g4437)) + ((!g2256) & (!g2295) & (g2887) & (g2956) & (!g4436) & (!g4437)) + ((!g2256) & (g2295) & (!g2887) & (!g2956) & (!g4436) & (!g4437)) + ((!g2256) & (g2295) & (!g2887) & (!g2956) & (!g4436) & (g4437)) + ((!g2256) & (g2295) & (!g2887) & (!g2956) & (g4436) & (!g4437)) + ((!g2256) & (g2295) & (!g2887) & (!g2956) & (g4436) & (g4437)) + ((!g2256) & (g2295) & (g2887) & (!g2956) & (!g4436) & (!g4437)) + ((!g2256) & (g2295) & (g2887) & (g2956) & (!g4436) & (g4437)) + ((!g2256) & (g2295) & (g2887) & (g2956) & (g4436) & (!g4437)) + ((!g2256) & (g2295) & (g2887) & (g2956) & (g4436) & (g4437)) + ((g2256) & (!g2295) & (!g2887) & (!g2956) & (!g4436) & (g4437)) + ((g2256) & (!g2295) & (!g2887) & (!g2956) & (g4436) & (!g4437)) + ((g2256) & (!g2295) & (!g2887) & (!g2956) & (g4436) & (g4437)) + ((g2256) & (!g2295) & (!g2887) & (g2956) & (!g4436) & (!g4437)) + ((g2256) & (!g2295) & (g2887) & (!g2956) & (!g4436) & (!g4437)) + ((g2256) & (!g2295) & (g2887) & (!g2956) & (!g4436) & (g4437)) + ((g2256) & (!g2295) & (g2887) & (!g2956) & (g4436) & (!g4437)) + ((g2256) & (!g2295) & (g2887) & (!g2956) & (g4436) & (g4437)) + ((g2256) & (g2295) & (!g2887) & (!g2956) & (!g4436) & (!g4437)) + ((g2256) & (g2295) & (!g2887) & (g2956) & (!g4436) & (g4437)) + ((g2256) & (g2295) & (!g2887) & (g2956) & (g4436) & (!g4437)) + ((g2256) & (g2295) & (!g2887) & (g2956) & (g4436) & (g4437)) + ((g2256) & (g2295) & (g2887) & (g2956) & (!g4436) & (!g4437)) + ((g2256) & (g2295) & (g2887) & (g2956) & (!g4436) & (g4437)) + ((g2256) & (g2295) & (g2887) & (g2956) & (g4436) & (!g4437)) + ((g2256) & (g2295) & (g2887) & (g2956) & (g4436) & (g4437)));
	assign g4496 = (((g830) & (!g1914) & (!g2271) & (!g4494) & (g4495)) + ((g830) & (!g1914) & (!g2271) & (g4494) & (g4495)) + ((g830) & (!g1914) & (g2271) & (!g4494) & (!g4495)) + ((g830) & (!g1914) & (g2271) & (g4494) & (!g4495)) + ((g830) & (g1914) & (!g2271) & (g4494) & (!g4495)) + ((g830) & (g1914) & (!g2271) & (g4494) & (g4495)) + ((g830) & (g1914) & (g2271) & (!g4494) & (!g4495)) + ((g830) & (g1914) & (g2271) & (!g4494) & (g4495)));
	assign g4497 = (((!g2518) & (g3119)) + ((g2518) & (!g3119)));
	assign g4498 = (((!g2378) & (!g2426) & (g3044) & (g3093) & (!g4339) & (g4497)) + ((!g2378) & (g2426) & (!g3044) & (g3093) & (!g4339) & (g4497)) + ((!g2378) & (g2426) & (!g3044) & (g3093) & (g4339) & (g4497)) + ((!g2378) & (g2426) & (g3044) & (!g3093) & (!g4339) & (g4497)) + ((!g2378) & (g2426) & (g3044) & (g3093) & (!g4339) & (g4497)) + ((!g2378) & (g2426) & (g3044) & (g3093) & (g4339) & (g4497)) + ((g2378) & (!g2426) & (!g3044) & (g3093) & (!g4339) & (g4497)) + ((g2378) & (!g2426) & (g3044) & (g3093) & (!g4339) & (g4497)) + ((g2378) & (!g2426) & (g3044) & (g3093) & (g4339) & (g4497)) + ((g2378) & (g2426) & (!g3044) & (!g3093) & (!g4339) & (g4497)) + ((g2378) & (g2426) & (!g3044) & (g3093) & (!g4339) & (g4497)) + ((g2378) & (g2426) & (!g3044) & (g3093) & (g4339) & (g4497)) + ((g2378) & (g2426) & (g3044) & (!g3093) & (!g4339) & (g4497)) + ((g2378) & (g2426) & (g3044) & (!g3093) & (g4339) & (g4497)) + ((g2378) & (g2426) & (g3044) & (g3093) & (!g4339) & (g4497)) + ((g2378) & (g2426) & (g3044) & (g3093) & (g4339) & (g4497)));
	assign g4499 = (((g2518) & (g3119)));
	assign g4500 = (((!g2555) & (!g3168) & (!g4498) & (g4499)) + ((!g2555) & (!g3168) & (g4498) & (!g4499)) + ((!g2555) & (!g3168) & (g4498) & (g4499)) + ((!g2555) & (g3168) & (!g4498) & (!g4499)) + ((g2555) & (!g3168) & (!g4498) & (!g4499)) + ((g2555) & (g3168) & (!g4498) & (g4499)) + ((g2555) & (g3168) & (g4498) & (!g4499)) + ((g2555) & (g3168) & (g4498) & (g4499)));
	assign g8304 = (((!g5560) & (g5600) & (!g4501)) + ((!g5560) & (g5600) & (g4501)) + ((g5560) & (!g5600) & (g4501)) + ((g5560) & (g5600) & (g4501)));
	assign g4502 = (((!g2516) & (g3131)) + ((g2516) & (!g3131)));
	assign g4503 = (((!g2377) & (!g2424) & (g3056) & (!g4353) & (g3095) & (g4502)) + ((!g2377) & (g2424) & (!g3056) & (!g4353) & (g3095) & (g4502)) + ((!g2377) & (g2424) & (!g3056) & (g4353) & (g3095) & (g4502)) + ((!g2377) & (g2424) & (g3056) & (!g4353) & (!g3095) & (g4502)) + ((!g2377) & (g2424) & (g3056) & (!g4353) & (g3095) & (g4502)) + ((!g2377) & (g2424) & (g3056) & (g4353) & (g3095) & (g4502)) + ((g2377) & (!g2424) & (!g3056) & (!g4353) & (g3095) & (g4502)) + ((g2377) & (!g2424) & (g3056) & (!g4353) & (g3095) & (g4502)) + ((g2377) & (!g2424) & (g3056) & (g4353) & (g3095) & (g4502)) + ((g2377) & (g2424) & (!g3056) & (!g4353) & (!g3095) & (g4502)) + ((g2377) & (g2424) & (!g3056) & (!g4353) & (g3095) & (g4502)) + ((g2377) & (g2424) & (!g3056) & (g4353) & (g3095) & (g4502)) + ((g2377) & (g2424) & (g3056) & (!g4353) & (!g3095) & (g4502)) + ((g2377) & (g2424) & (g3056) & (!g4353) & (g3095) & (g4502)) + ((g2377) & (g2424) & (g3056) & (g4353) & (!g3095) & (g4502)) + ((g2377) & (g2424) & (g3056) & (g4353) & (g3095) & (g4502)));
	assign g4504 = (((g2516) & (g3131)));
	assign g4505 = (((!g2552) & (!g4503) & (!g4504) & (g3170)) + ((!g2552) & (!g4503) & (g4504) & (!g3170)) + ((!g2552) & (g4503) & (!g4504) & (!g3170)) + ((!g2552) & (g4503) & (g4504) & (!g3170)) + ((g2552) & (!g4503) & (!g4504) & (!g3170)) + ((g2552) & (!g4503) & (g4504) & (g3170)) + ((g2552) & (g4503) & (!g4504) & (g3170)) + ((g2552) & (g4503) & (g4504) & (g3170)));
	assign g4506 = (((!g3125) & (g3131)) + ((g3125) & (!g3131)));
	assign g4507 = (((!g3050) & (!g3080) & (!g4320) & (g3056) & (g3095) & (g4506)) + ((!g3050) & (g3080) & (!g4320) & (!g3056) & (g3095) & (g4506)) + ((!g3050) & (g3080) & (!g4320) & (g3056) & (!g3095) & (g4506)) + ((!g3050) & (g3080) & (!g4320) & (g3056) & (g3095) & (g4506)) + ((!g3050) & (g3080) & (g4320) & (!g3056) & (g3095) & (g4506)) + ((!g3050) & (g3080) & (g4320) & (g3056) & (g3095) & (g4506)) + ((g3050) & (!g3080) & (!g4320) & (!g3056) & (g3095) & (g4506)) + ((g3050) & (!g3080) & (!g4320) & (g3056) & (g3095) & (g4506)) + ((g3050) & (!g3080) & (g4320) & (g3056) & (g3095) & (g4506)) + ((g3050) & (g3080) & (!g4320) & (!g3056) & (!g3095) & (g4506)) + ((g3050) & (g3080) & (!g4320) & (!g3056) & (g3095) & (g4506)) + ((g3050) & (g3080) & (!g4320) & (g3056) & (!g3095) & (g4506)) + ((g3050) & (g3080) & (!g4320) & (g3056) & (g3095) & (g4506)) + ((g3050) & (g3080) & (g4320) & (!g3056) & (g3095) & (g4506)) + ((g3050) & (g3080) & (g4320) & (g3056) & (!g3095) & (g4506)) + ((g3050) & (g3080) & (g4320) & (g3056) & (g3095) & (g4506)));
	assign g4508 = (((g3125) & (g3131)));
	assign g4509 = (((!g3155) & (!g3170) & (!g4507) & (g4508)) + ((!g3155) & (!g3170) & (g4507) & (!g4508)) + ((!g3155) & (!g3170) & (g4507) & (g4508)) + ((!g3155) & (g3170) & (!g4507) & (!g4508)) + ((g3155) & (!g3170) & (!g4507) & (!g4508)) + ((g3155) & (g3170) & (!g4507) & (g4508)) + ((g3155) & (g3170) & (g4507) & (!g4508)) + ((g3155) & (g3170) & (g4507) & (g4508)));
	assign g4510 = (((!g2515) & (g3136)) + ((g2515) & (!g3136)));
	assign g4511 = (((!g2376) & (!g2423) & (g3061) & (g3082) & (!g4328) & (g4510)) + ((!g2376) & (g2423) & (!g3061) & (g3082) & (!g4328) & (g4510)) + ((!g2376) & (g2423) & (!g3061) & (g3082) & (g4328) & (g4510)) + ((!g2376) & (g2423) & (g3061) & (!g3082) & (!g4328) & (g4510)) + ((!g2376) & (g2423) & (g3061) & (g3082) & (!g4328) & (g4510)) + ((!g2376) & (g2423) & (g3061) & (g3082) & (g4328) & (g4510)) + ((g2376) & (!g2423) & (!g3061) & (g3082) & (!g4328) & (g4510)) + ((g2376) & (!g2423) & (g3061) & (g3082) & (!g4328) & (g4510)) + ((g2376) & (!g2423) & (g3061) & (g3082) & (g4328) & (g4510)) + ((g2376) & (g2423) & (!g3061) & (!g3082) & (!g4328) & (g4510)) + ((g2376) & (g2423) & (!g3061) & (g3082) & (!g4328) & (g4510)) + ((g2376) & (g2423) & (!g3061) & (g3082) & (g4328) & (g4510)) + ((g2376) & (g2423) & (g3061) & (!g3082) & (!g4328) & (g4510)) + ((g2376) & (g2423) & (g3061) & (!g3082) & (g4328) & (g4510)) + ((g2376) & (g2423) & (g3061) & (g3082) & (!g4328) & (g4510)) + ((g2376) & (g2423) & (g3061) & (g3082) & (g4328) & (g4510)));
	assign g4512 = (((g2515) & (g3136)));
	assign g4513 = (((!g2551) & (!g3157) & (!g4511) & (g4512)) + ((!g2551) & (!g3157) & (g4511) & (!g4512)) + ((!g2551) & (!g3157) & (g4511) & (g4512)) + ((!g2551) & (g3157) & (!g4511) & (!g4512)) + ((g2551) & (!g3157) & (!g4511) & (!g4512)) + ((g2551) & (g3157) & (!g4511) & (g4512)) + ((g2551) & (g3157) & (g4511) & (!g4512)) + ((g2551) & (g3157) & (g4511) & (g4512)));
	assign g4514 = (((!g2881) & (g2902)) + ((g2881) & (!g2902)));
	assign g4515 = (((!g2797) & (!g2854) & (g2830) & (g2863) & (g4344) & (g4514)) + ((!g2797) & (g2854) & (!g2830) & (g2863) & (!g4344) & (g4514)) + ((!g2797) & (g2854) & (!g2830) & (g2863) & (g4344) & (g4514)) + ((!g2797) & (g2854) & (g2830) & (!g2863) & (g4344) & (g4514)) + ((!g2797) & (g2854) & (g2830) & (g2863) & (!g4344) & (g4514)) + ((!g2797) & (g2854) & (g2830) & (g2863) & (g4344) & (g4514)) + ((g2797) & (!g2854) & (!g2830) & (g2863) & (g4344) & (g4514)) + ((g2797) & (!g2854) & (g2830) & (g2863) & (!g4344) & (g4514)) + ((g2797) & (!g2854) & (g2830) & (g2863) & (g4344) & (g4514)) + ((g2797) & (g2854) & (!g2830) & (!g2863) & (g4344) & (g4514)) + ((g2797) & (g2854) & (!g2830) & (g2863) & (!g4344) & (g4514)) + ((g2797) & (g2854) & (!g2830) & (g2863) & (g4344) & (g4514)) + ((g2797) & (g2854) & (g2830) & (!g2863) & (!g4344) & (g4514)) + ((g2797) & (g2854) & (g2830) & (!g2863) & (g4344) & (g4514)) + ((g2797) & (g2854) & (g2830) & (g2863) & (!g4344) & (g4514)) + ((g2797) & (g2854) & (g2830) & (g2863) & (g4344) & (g4514)));
	assign g4516 = (((g2881) & (g2902)));
	assign g4517 = (((!g2950) & (!g2968) & (!g4515) & (g4516)) + ((!g2950) & (!g2968) & (g4515) & (!g4516)) + ((!g2950) & (!g2968) & (g4515) & (g4516)) + ((!g2950) & (g2968) & (!g4515) & (!g4516)) + ((g2950) & (!g2968) & (!g4515) & (!g4516)) + ((g2950) & (g2968) & (!g4515) & (g4516)) + ((g2950) & (g2968) & (g4515) & (!g4516)) + ((g2950) & (g2968) & (g4515) & (g4516)));
	assign g4518 = (((!g2891) & (!g2916) & (!g2897) & (g2985) & (!g4454) & (!g4455)) + ((!g2891) & (!g2916) & (!g2897) & (g2985) & (!g4454) & (g4455)) + ((!g2891) & (!g2916) & (!g2897) & (g2985) & (g4454) & (!g4455)) + ((!g2891) & (!g2916) & (!g2897) & (g2985) & (g4454) & (g4455)) + ((!g2891) & (!g2916) & (g2897) & (!g2985) & (!g4454) & (g4455)) + ((!g2891) & (!g2916) & (g2897) & (!g2985) & (g4454) & (!g4455)) + ((!g2891) & (!g2916) & (g2897) & (!g2985) & (g4454) & (g4455)) + ((!g2891) & (!g2916) & (g2897) & (g2985) & (!g4454) & (!g4455)) + ((!g2891) & (g2916) & (!g2897) & (!g2985) & (!g4454) & (!g4455)) + ((!g2891) & (g2916) & (!g2897) & (!g2985) & (!g4454) & (g4455)) + ((!g2891) & (g2916) & (!g2897) & (!g2985) & (g4454) & (!g4455)) + ((!g2891) & (g2916) & (!g2897) & (!g2985) & (g4454) & (g4455)) + ((!g2891) & (g2916) & (g2897) & (!g2985) & (!g4454) & (!g4455)) + ((!g2891) & (g2916) & (g2897) & (g2985) & (!g4454) & (g4455)) + ((!g2891) & (g2916) & (g2897) & (g2985) & (g4454) & (!g4455)) + ((!g2891) & (g2916) & (g2897) & (g2985) & (g4454) & (g4455)) + ((g2891) & (!g2916) & (!g2897) & (!g2985) & (!g4454) & (g4455)) + ((g2891) & (!g2916) & (!g2897) & (!g2985) & (g4454) & (!g4455)) + ((g2891) & (!g2916) & (!g2897) & (!g2985) & (g4454) & (g4455)) + ((g2891) & (!g2916) & (!g2897) & (g2985) & (!g4454) & (!g4455)) + ((g2891) & (!g2916) & (g2897) & (!g2985) & (!g4454) & (!g4455)) + ((g2891) & (!g2916) & (g2897) & (!g2985) & (!g4454) & (g4455)) + ((g2891) & (!g2916) & (g2897) & (!g2985) & (g4454) & (!g4455)) + ((g2891) & (!g2916) & (g2897) & (!g2985) & (g4454) & (g4455)) + ((g2891) & (g2916) & (!g2897) & (!g2985) & (!g4454) & (!g4455)) + ((g2891) & (g2916) & (!g2897) & (g2985) & (!g4454) & (g4455)) + ((g2891) & (g2916) & (!g2897) & (g2985) & (g4454) & (!g4455)) + ((g2891) & (g2916) & (!g2897) & (g2985) & (g4454) & (g4455)) + ((g2891) & (g2916) & (g2897) & (g2985) & (!g4454) & (!g4455)) + ((g2891) & (g2916) & (g2897) & (g2985) & (!g4454) & (g4455)) + ((g2891) & (g2916) & (g2897) & (g2985) & (g4454) & (!g4455)) + ((g2891) & (g2916) & (g2897) & (g2985) & (g4454) & (g4455)));
	assign g4519 = (((g830) & (!g1914) & (!g2281) & (!g4517) & (g4518)) + ((g830) & (!g1914) & (!g2281) & (g4517) & (g4518)) + ((g830) & (!g1914) & (g2281) & (!g4517) & (!g4518)) + ((g830) & (!g1914) & (g2281) & (g4517) & (!g4518)) + ((g830) & (g1914) & (!g2281) & (g4517) & (!g4518)) + ((g830) & (g1914) & (!g2281) & (g4517) & (g4518)) + ((g830) & (g1914) & (g2281) & (!g4517) & (!g4518)) + ((g830) & (g1914) & (g2281) & (!g4517) & (g4518)));
	assign g4520 = (((!g3260) & (!g3240) & (g3305) & (g3303) & (!g4403)) + ((!g3260) & (!g3240) & (g3305) & (g3303) & (g4403)) + ((!g3260) & (g3240) & (!g3305) & (g3303) & (!g4403)) + ((!g3260) & (g3240) & (g3305) & (!g3303) & (!g4403)) + ((!g3260) & (g3240) & (g3305) & (g3303) & (!g4403)) + ((!g3260) & (g3240) & (g3305) & (g3303) & (g4403)) + ((g3260) & (!g3240) & (!g3305) & (g3303) & (!g4403)) + ((g3260) & (!g3240) & (g3305) & (!g3303) & (!g4403)) + ((g3260) & (!g3240) & (g3305) & (g3303) & (!g4403)) + ((g3260) & (!g3240) & (g3305) & (g3303) & (g4403)) + ((g3260) & (g3240) & (!g3305) & (g3303) & (!g4403)) + ((g3260) & (g3240) & (!g3305) & (g3303) & (g4403)) + ((g3260) & (g3240) & (g3305) & (!g3303) & (!g4403)) + ((g3260) & (g3240) & (g3305) & (!g3303) & (g4403)) + ((g3260) & (g3240) & (g3305) & (g3303) & (!g4403)) + ((g3260) & (g3240) & (g3305) & (g3303) & (g4403)));
	assign g4521 = (((!g2648) & (!g2679) & (g3284) & (g3314) & (!g4405)) + ((!g2648) & (g2679) & (!g3284) & (g3314) & (!g4405)) + ((!g2648) & (g2679) & (!g3284) & (g3314) & (g4405)) + ((!g2648) & (g2679) & (g3284) & (!g3314) & (!g4405)) + ((!g2648) & (g2679) & (g3284) & (g3314) & (!g4405)) + ((!g2648) & (g2679) & (g3284) & (g3314) & (g4405)) + ((g2648) & (!g2679) & (!g3284) & (g3314) & (!g4405)) + ((g2648) & (!g2679) & (g3284) & (g3314) & (!g4405)) + ((g2648) & (!g2679) & (g3284) & (g3314) & (g4405)) + ((g2648) & (g2679) & (!g3284) & (!g3314) & (!g4405)) + ((g2648) & (g2679) & (!g3284) & (g3314) & (!g4405)) + ((g2648) & (g2679) & (!g3284) & (g3314) & (g4405)) + ((g2648) & (g2679) & (g3284) & (!g3314) & (!g4405)) + ((g2648) & (g2679) & (g3284) & (!g3314) & (g4405)) + ((g2648) & (g2679) & (g3284) & (g3314) & (!g4405)) + ((g2648) & (g2679) & (g3284) & (g3314) & (g4405)));
	assign g4522 = (((!g830) & (nonce[39]) & (!g1914) & (!g4520) & (!g4521) & (!g5674)) + ((!g830) & (nonce[39]) & (!g1914) & (!g4520) & (!g4521) & (g5674)) + ((!g830) & (nonce[39]) & (!g1914) & (!g4520) & (g4521) & (!g5674)) + ((!g830) & (nonce[39]) & (!g1914) & (!g4520) & (g4521) & (g5674)) + ((!g830) & (nonce[39]) & (!g1914) & (g4520) & (!g4521) & (!g5674)) + ((!g830) & (nonce[39]) & (!g1914) & (g4520) & (!g4521) & (g5674)) + ((!g830) & (nonce[39]) & (!g1914) & (g4520) & (g4521) & (!g5674)) + ((!g830) & (nonce[39]) & (!g1914) & (g4520) & (g4521) & (g5674)) + ((!g830) & (nonce[39]) & (g1914) & (!g4520) & (!g4521) & (!g5674)) + ((!g830) & (nonce[39]) & (g1914) & (!g4520) & (!g4521) & (g5674)) + ((!g830) & (nonce[39]) & (g1914) & (!g4520) & (g4521) & (!g5674)) + ((!g830) & (nonce[39]) & (g1914) & (!g4520) & (g4521) & (g5674)) + ((!g830) & (nonce[39]) & (g1914) & (g4520) & (!g4521) & (!g5674)) + ((!g830) & (nonce[39]) & (g1914) & (g4520) & (!g4521) & (g5674)) + ((!g830) & (nonce[39]) & (g1914) & (g4520) & (g4521) & (!g5674)) + ((!g830) & (nonce[39]) & (g1914) & (g4520) & (g4521) & (g5674)) + ((g830) & (!nonce[39]) & (!g1914) & (!g4520) & (!g4521) & (!g5674)) + ((g830) & (!nonce[39]) & (!g1914) & (!g4520) & (g4521) & (g5674)) + ((g830) & (!nonce[39]) & (!g1914) & (g4520) & (!g4521) & (!g5674)) + ((g830) & (!nonce[39]) & (!g1914) & (g4520) & (g4521) & (g5674)) + ((g830) & (!nonce[39]) & (g1914) & (!g4520) & (!g4521) & (!g5674)) + ((g830) & (!nonce[39]) & (g1914) & (!g4520) & (g4521) & (!g5674)) + ((g830) & (!nonce[39]) & (g1914) & (g4520) & (!g4521) & (g5674)) + ((g830) & (!nonce[39]) & (g1914) & (g4520) & (g4521) & (g5674)) + ((g830) & (nonce[39]) & (!g1914) & (!g4520) & (!g4521) & (!g5674)) + ((g830) & (nonce[39]) & (!g1914) & (!g4520) & (g4521) & (g5674)) + ((g830) & (nonce[39]) & (!g1914) & (g4520) & (!g4521) & (!g5674)) + ((g830) & (nonce[39]) & (!g1914) & (g4520) & (g4521) & (g5674)) + ((g830) & (nonce[39]) & (g1914) & (!g4520) & (!g4521) & (!g5674)) + ((g830) & (nonce[39]) & (g1914) & (!g4520) & (g4521) & (!g5674)) + ((g830) & (nonce[39]) & (g1914) & (g4520) & (!g4521) & (g5674)) + ((g830) & (nonce[39]) & (g1914) & (g4520) & (g4521) & (g5674)));
	assign g4523 = (((!g2519) & (g3139)) + ((g2519) & (!g3139)));
	assign g4524 = (((!g2379) & (!g2427) & (!g4331) & (g3064) & (g3090) & (g4523)) + ((!g2379) & (g2427) & (!g4331) & (!g3064) & (g3090) & (g4523)) + ((!g2379) & (g2427) & (!g4331) & (g3064) & (!g3090) & (g4523)) + ((!g2379) & (g2427) & (!g4331) & (g3064) & (g3090) & (g4523)) + ((!g2379) & (g2427) & (g4331) & (!g3064) & (g3090) & (g4523)) + ((!g2379) & (g2427) & (g4331) & (g3064) & (g3090) & (g4523)) + ((g2379) & (!g2427) & (!g4331) & (!g3064) & (g3090) & (g4523)) + ((g2379) & (!g2427) & (!g4331) & (g3064) & (g3090) & (g4523)) + ((g2379) & (!g2427) & (g4331) & (g3064) & (g3090) & (g4523)) + ((g2379) & (g2427) & (!g4331) & (!g3064) & (!g3090) & (g4523)) + ((g2379) & (g2427) & (!g4331) & (!g3064) & (g3090) & (g4523)) + ((g2379) & (g2427) & (!g4331) & (g3064) & (!g3090) & (g4523)) + ((g2379) & (g2427) & (!g4331) & (g3064) & (g3090) & (g4523)) + ((g2379) & (g2427) & (g4331) & (!g3064) & (g3090) & (g4523)) + ((g2379) & (g2427) & (g4331) & (g3064) & (!g3090) & (g4523)) + ((g2379) & (g2427) & (g4331) & (g3064) & (g3090) & (g4523)));
	assign g4525 = (((g2519) & (g3139)));
	assign g4526 = (((!g2556) & (!g3165) & (!g4524) & (g4525)) + ((!g2556) & (!g3165) & (g4524) & (!g4525)) + ((!g2556) & (!g3165) & (g4524) & (g4525)) + ((!g2556) & (g3165) & (!g4524) & (!g4525)) + ((g2556) & (!g3165) & (!g4524) & (!g4525)) + ((g2556) & (g3165) & (!g4524) & (g4525)) + ((g2556) & (g3165) & (g4524) & (!g4525)) + ((g2556) & (g3165) & (g4524) & (g4525)));
	assign g4527 = (((!g2650) & (!g2684) & (g3284) & (g3314) & (!g4411)) + ((!g2650) & (g2684) & (!g3284) & (g3314) & (!g4411)) + ((!g2650) & (g2684) & (!g3284) & (g3314) & (g4411)) + ((!g2650) & (g2684) & (g3284) & (!g3314) & (!g4411)) + ((!g2650) & (g2684) & (g3284) & (g3314) & (!g4411)) + ((!g2650) & (g2684) & (g3284) & (g3314) & (g4411)) + ((g2650) & (!g2684) & (!g3284) & (g3314) & (!g4411)) + ((g2650) & (!g2684) & (g3284) & (g3314) & (!g4411)) + ((g2650) & (!g2684) & (g3284) & (g3314) & (g4411)) + ((g2650) & (g2684) & (!g3284) & (!g3314) & (!g4411)) + ((g2650) & (g2684) & (!g3284) & (g3314) & (!g4411)) + ((g2650) & (g2684) & (!g3284) & (g3314) & (g4411)) + ((g2650) & (g2684) & (g3284) & (!g3314) & (!g4411)) + ((g2650) & (g2684) & (g3284) & (!g3314) & (g4411)) + ((g2650) & (g2684) & (g3284) & (g3314) & (!g4411)) + ((g2650) & (g2684) & (g3284) & (g3314) & (g4411)));
	assign g4528 = (((!g3260) & (!g3255) & (g3305) & (g3297) & (!g4413)) + ((!g3260) & (!g3255) & (g3305) & (g3297) & (g4413)) + ((!g3260) & (g3255) & (!g3305) & (g3297) & (!g4413)) + ((!g3260) & (g3255) & (g3305) & (!g3297) & (!g4413)) + ((!g3260) & (g3255) & (g3305) & (g3297) & (!g4413)) + ((!g3260) & (g3255) & (g3305) & (g3297) & (g4413)) + ((g3260) & (!g3255) & (!g3305) & (g3297) & (!g4413)) + ((g3260) & (!g3255) & (g3305) & (!g3297) & (!g4413)) + ((g3260) & (!g3255) & (g3305) & (g3297) & (!g4413)) + ((g3260) & (!g3255) & (g3305) & (g3297) & (g4413)) + ((g3260) & (g3255) & (!g3305) & (g3297) & (!g4413)) + ((g3260) & (g3255) & (!g3305) & (g3297) & (g4413)) + ((g3260) & (g3255) & (g3305) & (!g3297) & (!g4413)) + ((g3260) & (g3255) & (g3305) & (!g3297) & (g4413)) + ((g3260) & (g3255) & (g3305) & (g3297) & (!g4413)) + ((g3260) & (g3255) & (g3305) & (g3297) & (g4413)));
	assign g4529 = (((!g830) & (key[199]) & (!g1914) & (!g4527) & (!g4528) & (!g5675)) + ((!g830) & (key[199]) & (!g1914) & (!g4527) & (!g4528) & (g5675)) + ((!g830) & (key[199]) & (!g1914) & (!g4527) & (g4528) & (!g5675)) + ((!g830) & (key[199]) & (!g1914) & (!g4527) & (g4528) & (g5675)) + ((!g830) & (key[199]) & (!g1914) & (g4527) & (!g4528) & (!g5675)) + ((!g830) & (key[199]) & (!g1914) & (g4527) & (!g4528) & (g5675)) + ((!g830) & (key[199]) & (!g1914) & (g4527) & (g4528) & (!g5675)) + ((!g830) & (key[199]) & (!g1914) & (g4527) & (g4528) & (g5675)) + ((!g830) & (key[199]) & (g1914) & (!g4527) & (!g4528) & (!g5675)) + ((!g830) & (key[199]) & (g1914) & (!g4527) & (!g4528) & (g5675)) + ((!g830) & (key[199]) & (g1914) & (!g4527) & (g4528) & (!g5675)) + ((!g830) & (key[199]) & (g1914) & (!g4527) & (g4528) & (g5675)) + ((!g830) & (key[199]) & (g1914) & (g4527) & (!g4528) & (!g5675)) + ((!g830) & (key[199]) & (g1914) & (g4527) & (!g4528) & (g5675)) + ((!g830) & (key[199]) & (g1914) & (g4527) & (g4528) & (!g5675)) + ((!g830) & (key[199]) & (g1914) & (g4527) & (g4528) & (g5675)) + ((g830) & (!key[199]) & (!g1914) & (!g4527) & (!g4528) & (!g5675)) + ((g830) & (!key[199]) & (!g1914) & (!g4527) & (g4528) & (g5675)) + ((g830) & (!key[199]) & (!g1914) & (g4527) & (!g4528) & (!g5675)) + ((g830) & (!key[199]) & (!g1914) & (g4527) & (g4528) & (g5675)) + ((g830) & (!key[199]) & (g1914) & (!g4527) & (!g4528) & (!g5675)) + ((g830) & (!key[199]) & (g1914) & (!g4527) & (g4528) & (!g5675)) + ((g830) & (!key[199]) & (g1914) & (g4527) & (!g4528) & (g5675)) + ((g830) & (!key[199]) & (g1914) & (g4527) & (g4528) & (g5675)) + ((g830) & (key[199]) & (!g1914) & (!g4527) & (!g4528) & (!g5675)) + ((g830) & (key[199]) & (!g1914) & (!g4527) & (g4528) & (g5675)) + ((g830) & (key[199]) & (!g1914) & (g4527) & (!g4528) & (!g5675)) + ((g830) & (key[199]) & (!g1914) & (g4527) & (g4528) & (g5675)) + ((g830) & (key[199]) & (g1914) & (!g4527) & (!g4528) & (!g5675)) + ((g830) & (key[199]) & (g1914) & (!g4527) & (g4528) & (!g5675)) + ((g830) & (key[199]) & (g1914) & (g4527) & (!g4528) & (g5675)) + ((g830) & (key[199]) & (g1914) & (g4527) & (g4528) & (g5675)));
	assign g4530 = (((!g2889) & (g2897)) + ((g2889) & (!g2897)));
	assign g4531 = (((!g2810) & (!g2868) & (g2822) & (g2871) & (g4361) & (g4530)) + ((!g2810) & (g2868) & (!g2822) & (g2871) & (!g4361) & (g4530)) + ((!g2810) & (g2868) & (!g2822) & (g2871) & (g4361) & (g4530)) + ((!g2810) & (g2868) & (g2822) & (!g2871) & (g4361) & (g4530)) + ((!g2810) & (g2868) & (g2822) & (g2871) & (!g4361) & (g4530)) + ((!g2810) & (g2868) & (g2822) & (g2871) & (g4361) & (g4530)) + ((g2810) & (!g2868) & (!g2822) & (g2871) & (g4361) & (g4530)) + ((g2810) & (!g2868) & (g2822) & (g2871) & (!g4361) & (g4530)) + ((g2810) & (!g2868) & (g2822) & (g2871) & (g4361) & (g4530)) + ((g2810) & (g2868) & (!g2822) & (!g2871) & (g4361) & (g4530)) + ((g2810) & (g2868) & (!g2822) & (g2871) & (!g4361) & (g4530)) + ((g2810) & (g2868) & (!g2822) & (g2871) & (g4361) & (g4530)) + ((g2810) & (g2868) & (g2822) & (!g2871) & (!g4361) & (g4530)) + ((g2810) & (g2868) & (g2822) & (!g2871) & (g4361) & (g4530)) + ((g2810) & (g2868) & (g2822) & (g2871) & (!g4361) & (g4530)) + ((g2810) & (g2868) & (g2822) & (g2871) & (g4361) & (g4530)));
	assign g4532 = (((g2889) & (g2897)));
	assign g4533 = (((!g2979) & (!g2985) & (!g4531) & (g4532)) + ((!g2979) & (!g2985) & (g4531) & (!g4532)) + ((!g2979) & (!g2985) & (g4531) & (g4532)) + ((!g2979) & (g2985) & (!g4531) & (!g4532)) + ((g2979) & (!g2985) & (!g4531) & (!g4532)) + ((g2979) & (g2985) & (!g4531) & (g4532)) + ((g2979) & (g2985) & (g4531) & (!g4532)) + ((g2979) & (g2985) & (g4531) & (g4532)));
	assign g4534 = (((!g2900) & (!g2944) & (!g2902) & (g2968) & (!g4468) & (!g4469)) + ((!g2900) & (!g2944) & (!g2902) & (g2968) & (!g4468) & (g4469)) + ((!g2900) & (!g2944) & (!g2902) & (g2968) & (g4468) & (!g4469)) + ((!g2900) & (!g2944) & (!g2902) & (g2968) & (g4468) & (g4469)) + ((!g2900) & (!g2944) & (g2902) & (!g2968) & (!g4468) & (g4469)) + ((!g2900) & (!g2944) & (g2902) & (!g2968) & (g4468) & (!g4469)) + ((!g2900) & (!g2944) & (g2902) & (!g2968) & (g4468) & (g4469)) + ((!g2900) & (!g2944) & (g2902) & (g2968) & (!g4468) & (!g4469)) + ((!g2900) & (g2944) & (!g2902) & (!g2968) & (!g4468) & (!g4469)) + ((!g2900) & (g2944) & (!g2902) & (!g2968) & (!g4468) & (g4469)) + ((!g2900) & (g2944) & (!g2902) & (!g2968) & (g4468) & (!g4469)) + ((!g2900) & (g2944) & (!g2902) & (!g2968) & (g4468) & (g4469)) + ((!g2900) & (g2944) & (g2902) & (!g2968) & (!g4468) & (!g4469)) + ((!g2900) & (g2944) & (g2902) & (g2968) & (!g4468) & (g4469)) + ((!g2900) & (g2944) & (g2902) & (g2968) & (g4468) & (!g4469)) + ((!g2900) & (g2944) & (g2902) & (g2968) & (g4468) & (g4469)) + ((g2900) & (!g2944) & (!g2902) & (!g2968) & (!g4468) & (g4469)) + ((g2900) & (!g2944) & (!g2902) & (!g2968) & (g4468) & (!g4469)) + ((g2900) & (!g2944) & (!g2902) & (!g2968) & (g4468) & (g4469)) + ((g2900) & (!g2944) & (!g2902) & (g2968) & (!g4468) & (!g4469)) + ((g2900) & (!g2944) & (g2902) & (!g2968) & (!g4468) & (!g4469)) + ((g2900) & (!g2944) & (g2902) & (!g2968) & (!g4468) & (g4469)) + ((g2900) & (!g2944) & (g2902) & (!g2968) & (g4468) & (!g4469)) + ((g2900) & (!g2944) & (g2902) & (!g2968) & (g4468) & (g4469)) + ((g2900) & (g2944) & (!g2902) & (!g2968) & (!g4468) & (!g4469)) + ((g2900) & (g2944) & (!g2902) & (g2968) & (!g4468) & (g4469)) + ((g2900) & (g2944) & (!g2902) & (g2968) & (g4468) & (!g4469)) + ((g2900) & (g2944) & (!g2902) & (g2968) & (g4468) & (g4469)) + ((g2900) & (g2944) & (g2902) & (g2968) & (!g4468) & (!g4469)) + ((g2900) & (g2944) & (g2902) & (g2968) & (!g4468) & (g4469)) + ((g2900) & (g2944) & (g2902) & (g2968) & (g4468) & (!g4469)) + ((g2900) & (g2944) & (g2902) & (g2968) & (g4468) & (g4469)));
	assign g4535 = (((g830) & (!g1914) & (!g2290) & (!g4533) & (g4534)) + ((g830) & (!g1914) & (!g2290) & (g4533) & (g4534)) + ((g830) & (!g1914) & (g2290) & (!g4533) & (!g4534)) + ((g830) & (!g1914) & (g2290) & (g4533) & (!g4534)) + ((g830) & (g1914) & (!g2290) & (g4533) & (!g4534)) + ((g830) & (g1914) & (!g2290) & (g4533) & (g4534)) + ((g830) & (g1914) & (g2290) & (!g4533) & (!g4534)) + ((g830) & (g1914) & (g2290) & (!g4533) & (g4534)));
	assign g4536 = (((!g1199) & (!g1236) & (!g4472) & (!g2434) & (g2533)) + ((!g1199) & (!g1236) & (!g4472) & (g2434) & (!g2533)) + ((!g1199) & (!g1236) & (g4472) & (!g2434) & (g2533)) + ((!g1199) & (!g1236) & (g4472) & (g2434) & (g2533)) + ((!g1199) & (g1236) & (!g4472) & (!g2434) & (!g2533)) + ((!g1199) & (g1236) & (!g4472) & (g2434) & (g2533)) + ((!g1199) & (g1236) & (g4472) & (!g2434) & (!g2533)) + ((!g1199) & (g1236) & (g4472) & (g2434) & (!g2533)) + ((g1199) & (!g1236) & (!g4472) & (!g2434) & (!g2533)) + ((g1199) & (!g1236) & (!g4472) & (g2434) & (!g2533)) + ((g1199) & (!g1236) & (g4472) & (!g2434) & (g2533)) + ((g1199) & (!g1236) & (g4472) & (g2434) & (!g2533)) + ((g1199) & (g1236) & (!g4472) & (!g2434) & (g2533)) + ((g1199) & (g1236) & (!g4472) & (g2434) & (g2533)) + ((g1199) & (g1236) & (g4472) & (!g2434) & (!g2533)) + ((g1199) & (g1236) & (g4472) & (g2434) & (g2533)));
	assign g4537 = (((!g2450) & (!g2527) & (!g2497) & (g2531) & (!g4474)) + ((!g2450) & (!g2527) & (!g2497) & (g2531) & (g4474)) + ((!g2450) & (!g2527) & (g2497) & (!g2531) & (!g4474)) + ((!g2450) & (!g2527) & (g2497) & (g2531) & (g4474)) + ((!g2450) & (g2527) & (!g2497) & (!g2531) & (!g4474)) + ((!g2450) & (g2527) & (!g2497) & (!g2531) & (g4474)) + ((!g2450) & (g2527) & (g2497) & (!g2531) & (g4474)) + ((!g2450) & (g2527) & (g2497) & (g2531) & (!g4474)) + ((g2450) & (!g2527) & (!g2497) & (!g2531) & (!g4474)) + ((g2450) & (!g2527) & (!g2497) & (g2531) & (g4474)) + ((g2450) & (!g2527) & (g2497) & (!g2531) & (!g4474)) + ((g2450) & (!g2527) & (g2497) & (!g2531) & (g4474)) + ((g2450) & (g2527) & (!g2497) & (!g2531) & (g4474)) + ((g2450) & (g2527) & (!g2497) & (g2531) & (!g4474)) + ((g2450) & (g2527) & (g2497) & (g2531) & (!g4474)) + ((g2450) & (g2527) & (g2497) & (g2531) & (g4474)));
	assign g4538 = (((!g830) & (!g1914) & (!g2295) & (!g4536) & (!g4537) & (key[53])) + ((!g830) & (!g1914) & (!g2295) & (!g4536) & (g4537) & (key[53])) + ((!g830) & (!g1914) & (!g2295) & (g4536) & (!g4537) & (key[53])) + ((!g830) & (!g1914) & (!g2295) & (g4536) & (g4537) & (key[53])) + ((!g830) & (!g1914) & (g2295) & (!g4536) & (!g4537) & (key[53])) + ((!g830) & (!g1914) & (g2295) & (!g4536) & (g4537) & (key[53])) + ((!g830) & (!g1914) & (g2295) & (g4536) & (!g4537) & (key[53])) + ((!g830) & (!g1914) & (g2295) & (g4536) & (g4537) & (key[53])) + ((!g830) & (g1914) & (!g2295) & (!g4536) & (!g4537) & (key[53])) + ((!g830) & (g1914) & (!g2295) & (!g4536) & (g4537) & (key[53])) + ((!g830) & (g1914) & (!g2295) & (g4536) & (!g4537) & (key[53])) + ((!g830) & (g1914) & (!g2295) & (g4536) & (g4537) & (key[53])) + ((!g830) & (g1914) & (g2295) & (!g4536) & (!g4537) & (key[53])) + ((!g830) & (g1914) & (g2295) & (!g4536) & (g4537) & (key[53])) + ((!g830) & (g1914) & (g2295) & (g4536) & (!g4537) & (key[53])) + ((!g830) & (g1914) & (g2295) & (g4536) & (g4537) & (key[53])) + ((g830) & (!g1914) & (!g2295) & (!g4536) & (g4537) & (!key[53])) + ((g830) & (!g1914) & (!g2295) & (!g4536) & (g4537) & (key[53])) + ((g830) & (!g1914) & (!g2295) & (g4536) & (g4537) & (!key[53])) + ((g830) & (!g1914) & (!g2295) & (g4536) & (g4537) & (key[53])) + ((g830) & (!g1914) & (g2295) & (!g4536) & (!g4537) & (!key[53])) + ((g830) & (!g1914) & (g2295) & (!g4536) & (!g4537) & (key[53])) + ((g830) & (!g1914) & (g2295) & (g4536) & (!g4537) & (!key[53])) + ((g830) & (!g1914) & (g2295) & (g4536) & (!g4537) & (key[53])) + ((g830) & (g1914) & (!g2295) & (g4536) & (!g4537) & (!key[53])) + ((g830) & (g1914) & (!g2295) & (g4536) & (!g4537) & (key[53])) + ((g830) & (g1914) & (!g2295) & (g4536) & (g4537) & (!key[53])) + ((g830) & (g1914) & (!g2295) & (g4536) & (g4537) & (key[53])) + ((g830) & (g1914) & (g2295) & (!g4536) & (!g4537) & (!key[53])) + ((g830) & (g1914) & (g2295) & (!g4536) & (!g4537) & (key[53])) + ((g830) & (g1914) & (g2295) & (!g4536) & (g4537) & (!key[53])) + ((g830) & (g1914) & (g2295) & (!g4536) & (g4537) & (key[53])));
	assign g4539 = (((!g2572) & (g2595) & (!g3767)) + ((g2572) & (!g2595) & (!g3767)) + ((g2572) & (g2595) & (!g3767)) + ((g2572) & (g2595) & (g3767)));
	assign g4540 = (((!g1958) & (!g2320) & (!g3749)) + ((!g1958) & (g2320) & (g3749)) + ((g1958) & (!g2320) & (g3749)) + ((g1958) & (g2320) & (!g3749)));
	assign g4541 = (((!g1914) & (!g2637) & (!g2643) & (g4539) & (!g4540)) + ((!g1914) & (!g2637) & (!g2643) & (g4539) & (g4540)) + ((!g1914) & (!g2637) & (g2643) & (!g4539) & (!g4540)) + ((!g1914) & (!g2637) & (g2643) & (!g4539) & (g4540)) + ((!g1914) & (g2637) & (!g2643) & (!g4539) & (!g4540)) + ((!g1914) & (g2637) & (!g2643) & (!g4539) & (g4540)) + ((!g1914) & (g2637) & (g2643) & (g4539) & (!g4540)) + ((!g1914) & (g2637) & (g2643) & (g4539) & (g4540)) + ((g1914) & (!g2637) & (!g2643) & (!g4539) & (g4540)) + ((g1914) & (!g2637) & (!g2643) & (g4539) & (g4540)) + ((g1914) & (!g2637) & (g2643) & (!g4539) & (g4540)) + ((g1914) & (!g2637) & (g2643) & (g4539) & (g4540)) + ((g1914) & (g2637) & (!g2643) & (!g4539) & (g4540)) + ((g1914) & (g2637) & (!g2643) & (g4539) & (g4540)) + ((g1914) & (g2637) & (g2643) & (!g4539) & (g4540)) + ((g1914) & (g2637) & (g2643) & (g4539) & (g4540)));
	assign g4542 = (((!g830) & (!g2296) & (!g4541) & (key[85])) + ((!g830) & (!g2296) & (g4541) & (key[85])) + ((!g830) & (g2296) & (!g4541) & (key[85])) + ((!g830) & (g2296) & (g4541) & (key[85])) + ((g830) & (!g2296) & (g4541) & (!key[85])) + ((g830) & (!g2296) & (g4541) & (key[85])) + ((g830) & (g2296) & (!g4541) & (!key[85])) + ((g830) & (g2296) & (!g4541) & (key[85])));
	assign g4543 = (((!g4481) & (!g2450) & (!g2462) & (!g2527) & (g2542)) + ((!g4481) & (!g2450) & (!g2462) & (g2527) & (!g2542)) + ((!g4481) & (!g2450) & (g2462) & (!g2527) & (g2542)) + ((!g4481) & (!g2450) & (g2462) & (g2527) & (!g2542)) + ((!g4481) & (g2450) & (!g2462) & (!g2527) & (g2542)) + ((!g4481) & (g2450) & (!g2462) & (g2527) & (!g2542)) + ((!g4481) & (g2450) & (g2462) & (!g2527) & (!g2542)) + ((!g4481) & (g2450) & (g2462) & (g2527) & (g2542)) + ((g4481) & (!g2450) & (!g2462) & (!g2527) & (g2542)) + ((g4481) & (!g2450) & (!g2462) & (g2527) & (!g2542)) + ((g4481) & (!g2450) & (g2462) & (!g2527) & (!g2542)) + ((g4481) & (!g2450) & (g2462) & (g2527) & (g2542)) + ((g4481) & (g2450) & (!g2462) & (!g2527) & (!g2542)) + ((g4481) & (g2450) & (!g2462) & (g2527) & (g2542)) + ((g4481) & (g2450) & (g2462) & (!g2527) & (!g2542)) + ((g4481) & (g2450) & (g2462) & (g2527) & (g2542)));
	assign g4544 = (((!g1199) & (!g1236) & (!g4480) & (!g2468) & (g2523)) + ((!g1199) & (!g1236) & (!g4480) & (g2468) & (g2523)) + ((!g1199) & (!g1236) & (g4480) & (!g2468) & (g2523)) + ((!g1199) & (!g1236) & (g4480) & (g2468) & (!g2523)) + ((!g1199) & (g1236) & (!g4480) & (!g2468) & (!g2523)) + ((!g1199) & (g1236) & (!g4480) & (g2468) & (!g2523)) + ((!g1199) & (g1236) & (g4480) & (!g2468) & (!g2523)) + ((!g1199) & (g1236) & (g4480) & (g2468) & (g2523)) + ((g1199) & (!g1236) & (!g4480) & (!g2468) & (g2523)) + ((g1199) & (!g1236) & (!g4480) & (g2468) & (!g2523)) + ((g1199) & (!g1236) & (g4480) & (!g2468) & (!g2523)) + ((g1199) & (!g1236) & (g4480) & (g2468) & (!g2523)) + ((g1199) & (g1236) & (!g4480) & (!g2468) & (!g2523)) + ((g1199) & (g1236) & (!g4480) & (g2468) & (g2523)) + ((g1199) & (g1236) & (g4480) & (!g2468) & (g2523)) + ((g1199) & (g1236) & (g4480) & (g2468) & (g2523)));
	assign g8305 = (((!g5560) & (g5601) & (!g4545)) + ((!g5560) & (g5601) & (g4545)) + ((g5560) & (!g5601) & (g4545)) + ((g5560) & (g5601) & (g4545)));
	assign g4546 = (((!g830) & (!g1914) & (!g2298) & (!g4543) & (!g4544) & (g4545)) + ((!g830) & (!g1914) & (!g2298) & (!g4543) & (g4544) & (g4545)) + ((!g830) & (!g1914) & (!g2298) & (g4543) & (!g4544) & (g4545)) + ((!g830) & (!g1914) & (!g2298) & (g4543) & (g4544) & (g4545)) + ((!g830) & (!g1914) & (g2298) & (!g4543) & (!g4544) & (g4545)) + ((!g830) & (!g1914) & (g2298) & (!g4543) & (g4544) & (g4545)) + ((!g830) & (!g1914) & (g2298) & (g4543) & (!g4544) & (g4545)) + ((!g830) & (!g1914) & (g2298) & (g4543) & (g4544) & (g4545)) + ((!g830) & (g1914) & (!g2298) & (!g4543) & (!g4544) & (g4545)) + ((!g830) & (g1914) & (!g2298) & (!g4543) & (g4544) & (g4545)) + ((!g830) & (g1914) & (!g2298) & (g4543) & (!g4544) & (g4545)) + ((!g830) & (g1914) & (!g2298) & (g4543) & (g4544) & (g4545)) + ((!g830) & (g1914) & (g2298) & (!g4543) & (!g4544) & (g4545)) + ((!g830) & (g1914) & (g2298) & (!g4543) & (g4544) & (g4545)) + ((!g830) & (g1914) & (g2298) & (g4543) & (!g4544) & (g4545)) + ((!g830) & (g1914) & (g2298) & (g4543) & (g4544) & (g4545)) + ((g830) & (!g1914) & (!g2298) & (!g4543) & (g4544) & (!g4545)) + ((g830) & (!g1914) & (!g2298) & (!g4543) & (g4544) & (g4545)) + ((g830) & (!g1914) & (!g2298) & (g4543) & (g4544) & (!g4545)) + ((g830) & (!g1914) & (!g2298) & (g4543) & (g4544) & (g4545)) + ((g830) & (!g1914) & (g2298) & (!g4543) & (!g4544) & (!g4545)) + ((g830) & (!g1914) & (g2298) & (!g4543) & (!g4544) & (g4545)) + ((g830) & (!g1914) & (g2298) & (g4543) & (!g4544) & (!g4545)) + ((g830) & (!g1914) & (g2298) & (g4543) & (!g4544) & (g4545)) + ((g830) & (g1914) & (!g2298) & (g4543) & (!g4544) & (!g4545)) + ((g830) & (g1914) & (!g2298) & (g4543) & (!g4544) & (g4545)) + ((g830) & (g1914) & (!g2298) & (g4543) & (g4544) & (!g4545)) + ((g830) & (g1914) & (!g2298) & (g4543) & (g4544) & (g4545)) + ((g830) & (g1914) & (g2298) & (!g4543) & (!g4544) & (!g4545)) + ((g830) & (g1914) & (g2298) & (!g4543) & (!g4544) & (g4545)) + ((g830) & (g1914) & (g2298) & (!g4543) & (g4544) & (!g4545)) + ((g830) & (g1914) & (g2298) & (!g4543) & (g4544) & (g4545)));
	assign g4547 = (((!g3473) & (!g2589) & (g2595)) + ((!g3473) & (g2589) & (!g2595)) + ((!g3473) & (g2589) & (g2595)) + ((g3473) & (g2589) & (g2595)));
	assign g4548 = (((!g1996) & (!g2304) & (!g3487)) + ((!g1996) & (g2304) & (g3487)) + ((g1996) & (!g2304) & (g3487)) + ((g1996) & (g2304) & (!g3487)));
	assign g4549 = (((!g1914) & (!g4547) & (!g2620) & (!g2643) & (g4548)) + ((!g1914) & (!g4547) & (!g2620) & (g2643) & (g4548)) + ((!g1914) & (!g4547) & (g2620) & (!g2643) & (g4548)) + ((!g1914) & (!g4547) & (g2620) & (g2643) & (g4548)) + ((!g1914) & (g4547) & (!g2620) & (!g2643) & (g4548)) + ((!g1914) & (g4547) & (!g2620) & (g2643) & (g4548)) + ((!g1914) & (g4547) & (g2620) & (!g2643) & (g4548)) + ((!g1914) & (g4547) & (g2620) & (g2643) & (g4548)) + ((g1914) & (!g4547) & (!g2620) & (g2643) & (!g4548)) + ((g1914) & (!g4547) & (!g2620) & (g2643) & (g4548)) + ((g1914) & (!g4547) & (g2620) & (!g2643) & (!g4548)) + ((g1914) & (!g4547) & (g2620) & (!g2643) & (g4548)) + ((g1914) & (g4547) & (!g2620) & (!g2643) & (!g4548)) + ((g1914) & (g4547) & (!g2620) & (!g2643) & (g4548)) + ((g1914) & (g4547) & (g2620) & (g2643) & (!g4548)) + ((g1914) & (g4547) & (g2620) & (g2643) & (g4548)));
	assign g4550 = (((!g830) & (!g2299) & (!g4549) & (key[181])) + ((!g830) & (!g2299) & (g4549) & (key[181])) + ((!g830) & (g2299) & (!g4549) & (key[181])) + ((!g830) & (g2299) & (g4549) & (key[181])) + ((g830) & (!g2299) & (g4549) & (!key[181])) + ((g830) & (!g2299) & (g4549) & (key[181])) + ((g830) & (g2299) & (!g4549) & (!key[181])) + ((g830) & (g2299) & (!g4549) & (key[181])));
	assign g4551 = (((!g3155) & (!g3170) & (!g4507) & (!g4508)) + ((!g3155) & (!g3170) & (!g4507) & (g4508)) + ((!g3155) & (!g3170) & (g4507) & (!g4508)) + ((!g3155) & (!g3170) & (g4507) & (g4508)) + ((!g3155) & (g3170) & (!g4507) & (!g4508)) + ((g3155) & (!g3170) & (!g4507) & (!g4508)));
	assign g4552 = (((!g1888) & (!g1978) & (!g828) & (g864)) + ((!g1888) & (!g1978) & (g828) & (g864)) + ((!g1888) & (g1978) & (!g828) & (!g864)) + ((!g1888) & (g1978) & (g828) & (!g864)) + ((g1888) & (!g1978) & (!g828) & (g864)) + ((g1888) & (!g1978) & (g828) & (!g864)) + ((g1888) & (g1978) & (!g828) & (!g864)) + ((g1888) & (g1978) & (g828) & (g864)));
	assign g4553 = (((!g1914) & (!g3196) & (!g4551) & (!g3202) & (g4552)) + ((!g1914) & (!g3196) & (!g4551) & (g3202) & (g4552)) + ((!g1914) & (!g3196) & (g4551) & (!g3202) & (g4552)) + ((!g1914) & (!g3196) & (g4551) & (g3202) & (g4552)) + ((!g1914) & (g3196) & (!g4551) & (!g3202) & (g4552)) + ((!g1914) & (g3196) & (!g4551) & (g3202) & (g4552)) + ((!g1914) & (g3196) & (g4551) & (!g3202) & (g4552)) + ((!g1914) & (g3196) & (g4551) & (g3202) & (g4552)) + ((g1914) & (!g3196) & (!g4551) & (!g3202) & (!g4552)) + ((g1914) & (!g3196) & (!g4551) & (!g3202) & (g4552)) + ((g1914) & (!g3196) & (g4551) & (g3202) & (!g4552)) + ((g1914) & (!g3196) & (g4551) & (g3202) & (g4552)) + ((g1914) & (g3196) & (!g4551) & (g3202) & (!g4552)) + ((g1914) & (g3196) & (!g4551) & (g3202) & (g4552)) + ((g1914) & (g3196) & (g4551) & (!g3202) & (!g4552)) + ((g1914) & (g3196) & (g4551) & (!g3202) & (g4552)));
	assign g4554 = (((!g830) & (!g2304) & (!g4553) & (key[104])) + ((!g830) & (!g2304) & (g4553) & (key[104])) + ((!g830) & (g2304) & (!g4553) & (key[104])) + ((!g830) & (g2304) & (g4553) & (key[104])) + ((g830) & (!g2304) & (g4553) & (!key[104])) + ((g830) & (!g2304) & (g4553) & (key[104])) + ((g830) & (g2304) & (!g4553) & (!key[104])) + ((g830) & (g2304) & (!g4553) & (key[104])));
	assign g4555 = (((!g2298) & (!g2347) & (!g2938) & (g3011) & (!g4492) & (!g4493)) + ((!g2298) & (!g2347) & (!g2938) & (g3011) & (!g4492) & (g4493)) + ((!g2298) & (!g2347) & (!g2938) & (g3011) & (g4492) & (!g4493)) + ((!g2298) & (!g2347) & (!g2938) & (g3011) & (g4492) & (g4493)) + ((!g2298) & (!g2347) & (g2938) & (!g3011) & (!g4492) & (g4493)) + ((!g2298) & (!g2347) & (g2938) & (!g3011) & (g4492) & (!g4493)) + ((!g2298) & (!g2347) & (g2938) & (!g3011) & (g4492) & (g4493)) + ((!g2298) & (!g2347) & (g2938) & (g3011) & (!g4492) & (!g4493)) + ((!g2298) & (g2347) & (!g2938) & (!g3011) & (!g4492) & (!g4493)) + ((!g2298) & (g2347) & (!g2938) & (!g3011) & (!g4492) & (g4493)) + ((!g2298) & (g2347) & (!g2938) & (!g3011) & (g4492) & (!g4493)) + ((!g2298) & (g2347) & (!g2938) & (!g3011) & (g4492) & (g4493)) + ((!g2298) & (g2347) & (g2938) & (!g3011) & (!g4492) & (!g4493)) + ((!g2298) & (g2347) & (g2938) & (g3011) & (!g4492) & (g4493)) + ((!g2298) & (g2347) & (g2938) & (g3011) & (g4492) & (!g4493)) + ((!g2298) & (g2347) & (g2938) & (g3011) & (g4492) & (g4493)) + ((g2298) & (!g2347) & (!g2938) & (!g3011) & (!g4492) & (g4493)) + ((g2298) & (!g2347) & (!g2938) & (!g3011) & (g4492) & (!g4493)) + ((g2298) & (!g2347) & (!g2938) & (!g3011) & (g4492) & (g4493)) + ((g2298) & (!g2347) & (!g2938) & (g3011) & (!g4492) & (!g4493)) + ((g2298) & (!g2347) & (g2938) & (!g3011) & (!g4492) & (!g4493)) + ((g2298) & (!g2347) & (g2938) & (!g3011) & (!g4492) & (g4493)) + ((g2298) & (!g2347) & (g2938) & (!g3011) & (g4492) & (!g4493)) + ((g2298) & (!g2347) & (g2938) & (!g3011) & (g4492) & (g4493)) + ((g2298) & (g2347) & (!g2938) & (!g3011) & (!g4492) & (!g4493)) + ((g2298) & (g2347) & (!g2938) & (g3011) & (!g4492) & (g4493)) + ((g2298) & (g2347) & (!g2938) & (g3011) & (g4492) & (!g4493)) + ((g2298) & (g2347) & (!g2938) & (g3011) & (g4492) & (g4493)) + ((g2298) & (g2347) & (g2938) & (g3011) & (!g4492) & (!g4493)) + ((g2298) & (g2347) & (g2938) & (g3011) & (!g4492) & (g4493)) + ((g2298) & (g2347) & (g2938) & (g3011) & (g4492) & (!g4493)) + ((g2298) & (g2347) & (g2938) & (g3011) & (g4492) & (g4493)));
	assign g4556 = (((!g2256) & (!g2295) & (g2887) & (g2956) & (!g4436) & (g4437)) + ((!g2256) & (!g2295) & (g2887) & (g2956) & (g4436) & (!g4437)) + ((!g2256) & (!g2295) & (g2887) & (g2956) & (g4436) & (g4437)) + ((!g2256) & (g2295) & (!g2887) & (g2956) & (!g4436) & (!g4437)) + ((!g2256) & (g2295) & (!g2887) & (g2956) & (!g4436) & (g4437)) + ((!g2256) & (g2295) & (!g2887) & (g2956) & (g4436) & (!g4437)) + ((!g2256) & (g2295) & (!g2887) & (g2956) & (g4436) & (g4437)) + ((!g2256) & (g2295) & (g2887) & (!g2956) & (!g4436) & (g4437)) + ((!g2256) & (g2295) & (g2887) & (!g2956) & (g4436) & (!g4437)) + ((!g2256) & (g2295) & (g2887) & (!g2956) & (g4436) & (g4437)) + ((!g2256) & (g2295) & (g2887) & (g2956) & (!g4436) & (!g4437)) + ((!g2256) & (g2295) & (g2887) & (g2956) & (!g4436) & (g4437)) + ((!g2256) & (g2295) & (g2887) & (g2956) & (g4436) & (!g4437)) + ((!g2256) & (g2295) & (g2887) & (g2956) & (g4436) & (g4437)) + ((g2256) & (!g2295) & (!g2887) & (g2956) & (!g4436) & (g4437)) + ((g2256) & (!g2295) & (!g2887) & (g2956) & (g4436) & (!g4437)) + ((g2256) & (!g2295) & (!g2887) & (g2956) & (g4436) & (g4437)) + ((g2256) & (!g2295) & (g2887) & (g2956) & (!g4436) & (!g4437)) + ((g2256) & (!g2295) & (g2887) & (g2956) & (!g4436) & (g4437)) + ((g2256) & (!g2295) & (g2887) & (g2956) & (g4436) & (!g4437)) + ((g2256) & (!g2295) & (g2887) & (g2956) & (g4436) & (g4437)) + ((g2256) & (g2295) & (!g2887) & (!g2956) & (!g4436) & (g4437)) + ((g2256) & (g2295) & (!g2887) & (!g2956) & (g4436) & (!g4437)) + ((g2256) & (g2295) & (!g2887) & (!g2956) & (g4436) & (g4437)) + ((g2256) & (g2295) & (!g2887) & (g2956) & (!g4436) & (!g4437)) + ((g2256) & (g2295) & (!g2887) & (g2956) & (!g4436) & (g4437)) + ((g2256) & (g2295) & (!g2887) & (g2956) & (g4436) & (!g4437)) + ((g2256) & (g2295) & (!g2887) & (g2956) & (g4436) & (g4437)) + ((g2256) & (g2295) & (g2887) & (!g2956) & (!g4436) & (!g4437)) + ((g2256) & (g2295) & (g2887) & (!g2956) & (!g4436) & (g4437)) + ((g2256) & (g2295) & (g2887) & (!g2956) & (g4436) & (!g4437)) + ((g2256) & (g2295) & (g2887) & (!g2956) & (g4436) & (g4437)) + ((g2256) & (g2295) & (g2887) & (g2956) & (!g4436) & (!g4437)) + ((g2256) & (g2295) & (g2887) & (g2956) & (!g4436) & (g4437)) + ((g2256) & (g2295) & (g2887) & (g2956) & (g4436) & (!g4437)) + ((g2256) & (g2295) & (g2887) & (g2956) & (g4436) & (g4437)));
	assign g4557 = (((!g1886) & (!g2032) & (!g1902) & (g2036)) + ((!g1886) & (!g2032) & (g1902) & (g2036)) + ((!g1886) & (g2032) & (!g1902) & (!g2036)) + ((!g1886) & (g2032) & (g1902) & (!g2036)) + ((g1886) & (!g2032) & (!g1902) & (g2036)) + ((g1886) & (!g2032) & (g1902) & (!g2036)) + ((g1886) & (g2032) & (!g1902) & (!g2036)) + ((g1886) & (g2032) & (g1902) & (g2036)));
	assign g4558 = (((!g2551) & (!g3157) & (!g4511) & (!g4512)) + ((!g2551) & (!g3157) & (!g4511) & (g4512)) + ((!g2551) & (!g3157) & (g4511) & (!g4512)) + ((!g2551) & (!g3157) & (g4511) & (g4512)) + ((!g2551) & (g3157) & (!g4511) & (!g4512)) + ((g2551) & (!g3157) & (!g4511) & (!g4512)));
	assign g4559 = (((!g1914) & (!g2598) & (!g3207) & (!g4557) & (!g4558)) + ((!g1914) & (!g2598) & (!g3207) & (g4557) & (!g4558)) + ((!g1914) & (!g2598) & (g3207) & (!g4557) & (g4558)) + ((!g1914) & (!g2598) & (g3207) & (g4557) & (g4558)) + ((!g1914) & (g2598) & (!g3207) & (!g4557) & (g4558)) + ((!g1914) & (g2598) & (!g3207) & (g4557) & (g4558)) + ((!g1914) & (g2598) & (g3207) & (!g4557) & (!g4558)) + ((!g1914) & (g2598) & (g3207) & (g4557) & (!g4558)) + ((g1914) & (!g2598) & (!g3207) & (g4557) & (!g4558)) + ((g1914) & (!g2598) & (!g3207) & (g4557) & (g4558)) + ((g1914) & (!g2598) & (g3207) & (g4557) & (!g4558)) + ((g1914) & (!g2598) & (g3207) & (g4557) & (g4558)) + ((g1914) & (g2598) & (!g3207) & (g4557) & (!g4558)) + ((g1914) & (g2598) & (!g3207) & (g4557) & (g4558)) + ((g1914) & (g2598) & (g3207) & (g4557) & (!g4558)) + ((g1914) & (g2598) & (g3207) & (g4557) & (g4558)));
	assign g4560 = (((!g830) & (!g2314) & (!g4559) & (nonce[8])) + ((!g830) & (!g2314) & (g4559) & (nonce[8])) + ((!g830) & (g2314) & (!g4559) & (nonce[8])) + ((!g830) & (g2314) & (g4559) & (nonce[8])) + ((g830) & (!g2314) & (g4559) & (!nonce[8])) + ((g830) & (!g2314) & (g4559) & (nonce[8])) + ((g830) & (g2314) & (!g4559) & (!nonce[8])) + ((g830) & (g2314) & (!g4559) & (nonce[8])));
	assign g4561 = (((!g2556) & (!g3165) & (!g4524) & (!g4525)) + ((!g2556) & (!g3165) & (!g4524) & (g4525)) + ((!g2556) & (!g3165) & (g4524) & (!g4525)) + ((!g2556) & (!g3165) & (g4524) & (g4525)) + ((!g2556) & (g3165) & (!g4524) & (!g4525)) + ((g2556) & (!g3165) & (!g4524) & (!g4525)));
	assign g4562 = (((!g1892) & (!g2026) & (!g1894) & (g2034)) + ((!g1892) & (!g2026) & (g1894) & (g2034)) + ((!g1892) & (g2026) & (!g1894) & (!g2034)) + ((!g1892) & (g2026) & (g1894) & (!g2034)) + ((g1892) & (!g2026) & (!g1894) & (g2034)) + ((g1892) & (!g2026) & (g1894) & (!g2034)) + ((g1892) & (g2026) & (!g1894) & (!g2034)) + ((g1892) & (g2026) & (g1894) & (g2034)));
	assign g4563 = (((!g1914) & (!g2602) & (!g4561) & (!g3210) & (g4562)) + ((!g1914) & (!g2602) & (!g4561) & (g3210) & (g4562)) + ((!g1914) & (!g2602) & (g4561) & (!g3210) & (g4562)) + ((!g1914) & (!g2602) & (g4561) & (g3210) & (g4562)) + ((!g1914) & (g2602) & (!g4561) & (!g3210) & (g4562)) + ((!g1914) & (g2602) & (!g4561) & (g3210) & (g4562)) + ((!g1914) & (g2602) & (g4561) & (!g3210) & (g4562)) + ((!g1914) & (g2602) & (g4561) & (g3210) & (g4562)) + ((g1914) & (!g2602) & (!g4561) & (!g3210) & (!g4562)) + ((g1914) & (!g2602) & (!g4561) & (!g3210) & (g4562)) + ((g1914) & (!g2602) & (g4561) & (g3210) & (!g4562)) + ((g1914) & (!g2602) & (g4561) & (g3210) & (g4562)) + ((g1914) & (g2602) & (!g4561) & (g3210) & (!g4562)) + ((g1914) & (g2602) & (!g4561) & (g3210) & (g4562)) + ((g1914) & (g2602) & (g4561) & (!g3210) & (!g4562)) + ((g1914) & (g2602) & (g4561) & (!g3210) & (g4562)));
	assign g4564 = (((!g830) & (!g2317) & (!g4563) & (key[232])) + ((!g830) & (!g2317) & (g4563) & (key[232])) + ((!g830) & (g2317) & (!g4563) & (key[232])) + ((!g830) & (g2317) & (g4563) & (key[232])) + ((g830) & (!g2317) & (g4563) & (!key[232])) + ((g830) & (!g2317) & (g4563) & (key[232])) + ((g830) & (g2317) & (!g4563) & (!key[232])) + ((g830) & (g2317) & (!g4563) & (key[232])));
	assign g4565 = (((!g1906) & (!g1940) & (!g828) & (g864)) + ((!g1906) & (!g1940) & (g828) & (g864)) + ((!g1906) & (g1940) & (!g828) & (!g864)) + ((!g1906) & (g1940) & (g828) & (!g864)) + ((g1906) & (!g1940) & (!g828) & (g864)) + ((g1906) & (!g1940) & (g828) & (!g864)) + ((g1906) & (g1940) & (!g828) & (!g864)) + ((g1906) & (g1940) & (g828) & (g864)));
	assign g4566 = (((!g3161) & (!g4488) & (!g4489) & (!g3165)) + ((!g3161) & (!g4488) & (!g4489) & (g3165)) + ((!g3161) & (!g4488) & (g4489) & (!g3165)) + ((!g3161) & (g4488) & (!g4489) & (!g3165)) + ((!g3161) & (g4488) & (g4489) & (!g3165)) + ((g3161) & (!g4488) & (!g4489) & (!g3165)));
	assign g4567 = (((!g1914) & (!g3187) & (!g3210) & (!g4565) & (!g4566)) + ((!g1914) & (!g3187) & (!g3210) & (g4565) & (!g4566)) + ((!g1914) & (!g3187) & (g3210) & (!g4565) & (g4566)) + ((!g1914) & (!g3187) & (g3210) & (g4565) & (g4566)) + ((!g1914) & (g3187) & (!g3210) & (!g4565) & (g4566)) + ((!g1914) & (g3187) & (!g3210) & (g4565) & (g4566)) + ((!g1914) & (g3187) & (g3210) & (!g4565) & (!g4566)) + ((!g1914) & (g3187) & (g3210) & (g4565) & (!g4566)) + ((g1914) & (!g3187) & (!g3210) & (g4565) & (!g4566)) + ((g1914) & (!g3187) & (!g3210) & (g4565) & (g4566)) + ((g1914) & (!g3187) & (g3210) & (g4565) & (!g4566)) + ((g1914) & (!g3187) & (g3210) & (g4565) & (g4566)) + ((g1914) & (g3187) & (!g3210) & (g4565) & (!g4566)) + ((g1914) & (g3187) & (!g3210) & (g4565) & (g4566)) + ((g1914) & (g3187) & (g3210) & (g4565) & (!g4566)) + ((g1914) & (g3187) & (g3210) & (g4565) & (g4566)));
	assign g4568 = (((!g830) & (!g2320) & (!g4567) & (key[8])) + ((!g830) & (!g2320) & (g4567) & (key[8])) + ((!g830) & (g2320) & (!g4567) & (key[8])) + ((!g830) & (g2320) & (g4567) & (key[8])) + ((g830) & (!g2320) & (g4567) & (!key[8])) + ((g830) & (!g2320) & (g4567) & (key[8])) + ((g830) & (g2320) & (!g4567) & (!key[8])) + ((g830) & (g2320) & (!g4567) & (key[8])));
	assign g4569 = (((!g2555) & (!g3168) & (!g4498) & (!g4499)) + ((!g2555) & (!g3168) & (!g4498) & (g4499)) + ((!g2555) & (!g3168) & (g4498) & (!g4499)) + ((!g2555) & (!g3168) & (g4498) & (g4499)) + ((!g2555) & (g3168) & (!g4498) & (!g4499)) + ((g2555) & (!g3168) & (!g4498) & (!g4499)));
	assign g4570 = (((!g1898) & (!g2022) & (!g1902) & (g2036)) + ((!g1898) & (!g2022) & (g1902) & (g2036)) + ((!g1898) & (g2022) & (!g1902) & (!g2036)) + ((!g1898) & (g2022) & (g1902) & (!g2036)) + ((g1898) & (!g2022) & (!g1902) & (g2036)) + ((g1898) & (!g2022) & (g1902) & (!g2036)) + ((g1898) & (g2022) & (!g1902) & (!g2036)) + ((g1898) & (g2022) & (g1902) & (g2036)));
	assign g4571 = (((!g1914) & (!g2601) & (!g3190) & (!g4569) & (g4570)) + ((!g1914) & (!g2601) & (!g3190) & (g4569) & (g4570)) + ((!g1914) & (!g2601) & (g3190) & (!g4569) & (g4570)) + ((!g1914) & (!g2601) & (g3190) & (g4569) & (g4570)) + ((!g1914) & (g2601) & (!g3190) & (!g4569) & (g4570)) + ((!g1914) & (g2601) & (!g3190) & (g4569) & (g4570)) + ((!g1914) & (g2601) & (g3190) & (!g4569) & (g4570)) + ((!g1914) & (g2601) & (g3190) & (g4569) & (g4570)) + ((g1914) & (!g2601) & (!g3190) & (!g4569) & (!g4570)) + ((g1914) & (!g2601) & (!g3190) & (!g4569) & (g4570)) + ((g1914) & (!g2601) & (g3190) & (g4569) & (!g4570)) + ((g1914) & (!g2601) & (g3190) & (g4569) & (g4570)) + ((g1914) & (g2601) & (!g3190) & (g4569) & (!g4570)) + ((g1914) & (g2601) & (!g3190) & (g4569) & (g4570)) + ((g1914) & (g2601) & (g3190) & (!g4569) & (!g4570)) + ((g1914) & (g2601) & (g3190) & (!g4569) & (g4570)));
	assign g8306 = (((!g5560) & (g5602) & (!g4572)) + ((!g5560) & (g5602) & (g4572)) + ((g5560) & (!g5602) & (g4572)) + ((g5560) & (g5602) & (g4572)));
	assign g4573 = (((!g830) & (!g2323) & (!g4571) & (g4572)) + ((!g830) & (!g2323) & (g4571) & (g4572)) + ((!g830) & (g2323) & (!g4571) & (g4572)) + ((!g830) & (g2323) & (g4571) & (g4572)) + ((g830) & (!g2323) & (g4571) & (!g4572)) + ((g830) & (!g2323) & (g4571) & (g4572)) + ((g830) & (g2323) & (!g4571) & (!g4572)) + ((g830) & (g2323) & (!g4571) & (g4572)));
	assign g4574 = (((!g2950) & (!g2999) & (!g2968) & (g3020) & (!g4515) & (!g4516)) + ((!g2950) & (!g2999) & (!g2968) & (g3020) & (!g4515) & (g4516)) + ((!g2950) & (!g2999) & (!g2968) & (g3020) & (g4515) & (!g4516)) + ((!g2950) & (!g2999) & (!g2968) & (g3020) & (g4515) & (g4516)) + ((!g2950) & (!g2999) & (g2968) & (!g3020) & (!g4515) & (g4516)) + ((!g2950) & (!g2999) & (g2968) & (!g3020) & (g4515) & (!g4516)) + ((!g2950) & (!g2999) & (g2968) & (!g3020) & (g4515) & (g4516)) + ((!g2950) & (!g2999) & (g2968) & (g3020) & (!g4515) & (!g4516)) + ((!g2950) & (g2999) & (!g2968) & (!g3020) & (!g4515) & (!g4516)) + ((!g2950) & (g2999) & (!g2968) & (!g3020) & (!g4515) & (g4516)) + ((!g2950) & (g2999) & (!g2968) & (!g3020) & (g4515) & (!g4516)) + ((!g2950) & (g2999) & (!g2968) & (!g3020) & (g4515) & (g4516)) + ((!g2950) & (g2999) & (g2968) & (!g3020) & (!g4515) & (!g4516)) + ((!g2950) & (g2999) & (g2968) & (g3020) & (!g4515) & (g4516)) + ((!g2950) & (g2999) & (g2968) & (g3020) & (g4515) & (!g4516)) + ((!g2950) & (g2999) & (g2968) & (g3020) & (g4515) & (g4516)) + ((g2950) & (!g2999) & (!g2968) & (!g3020) & (!g4515) & (g4516)) + ((g2950) & (!g2999) & (!g2968) & (!g3020) & (g4515) & (!g4516)) + ((g2950) & (!g2999) & (!g2968) & (!g3020) & (g4515) & (g4516)) + ((g2950) & (!g2999) & (!g2968) & (g3020) & (!g4515) & (!g4516)) + ((g2950) & (!g2999) & (g2968) & (!g3020) & (!g4515) & (!g4516)) + ((g2950) & (!g2999) & (g2968) & (!g3020) & (!g4515) & (g4516)) + ((g2950) & (!g2999) & (g2968) & (!g3020) & (g4515) & (!g4516)) + ((g2950) & (!g2999) & (g2968) & (!g3020) & (g4515) & (g4516)) + ((g2950) & (g2999) & (!g2968) & (!g3020) & (!g4515) & (!g4516)) + ((g2950) & (g2999) & (!g2968) & (g3020) & (!g4515) & (g4516)) + ((g2950) & (g2999) & (!g2968) & (g3020) & (g4515) & (!g4516)) + ((g2950) & (g2999) & (!g2968) & (g3020) & (g4515) & (g4516)) + ((g2950) & (g2999) & (g2968) & (g3020) & (!g4515) & (!g4516)) + ((g2950) & (g2999) & (g2968) & (g3020) & (!g4515) & (g4516)) + ((g2950) & (g2999) & (g2968) & (g3020) & (g4515) & (!g4516)) + ((g2950) & (g2999) & (g2968) & (g3020) & (g4515) & (g4516)));
	assign g4575 = (((!g2891) & (!g2916) & (g2897) & (g2985) & (!g4454) & (g4455)) + ((!g2891) & (!g2916) & (g2897) & (g2985) & (g4454) & (!g4455)) + ((!g2891) & (!g2916) & (g2897) & (g2985) & (g4454) & (g4455)) + ((!g2891) & (g2916) & (!g2897) & (g2985) & (!g4454) & (!g4455)) + ((!g2891) & (g2916) & (!g2897) & (g2985) & (!g4454) & (g4455)) + ((!g2891) & (g2916) & (!g2897) & (g2985) & (g4454) & (!g4455)) + ((!g2891) & (g2916) & (!g2897) & (g2985) & (g4454) & (g4455)) + ((!g2891) & (g2916) & (g2897) & (!g2985) & (!g4454) & (g4455)) + ((!g2891) & (g2916) & (g2897) & (!g2985) & (g4454) & (!g4455)) + ((!g2891) & (g2916) & (g2897) & (!g2985) & (g4454) & (g4455)) + ((!g2891) & (g2916) & (g2897) & (g2985) & (!g4454) & (!g4455)) + ((!g2891) & (g2916) & (g2897) & (g2985) & (!g4454) & (g4455)) + ((!g2891) & (g2916) & (g2897) & (g2985) & (g4454) & (!g4455)) + ((!g2891) & (g2916) & (g2897) & (g2985) & (g4454) & (g4455)) + ((g2891) & (!g2916) & (!g2897) & (g2985) & (!g4454) & (g4455)) + ((g2891) & (!g2916) & (!g2897) & (g2985) & (g4454) & (!g4455)) + ((g2891) & (!g2916) & (!g2897) & (g2985) & (g4454) & (g4455)) + ((g2891) & (!g2916) & (g2897) & (g2985) & (!g4454) & (!g4455)) + ((g2891) & (!g2916) & (g2897) & (g2985) & (!g4454) & (g4455)) + ((g2891) & (!g2916) & (g2897) & (g2985) & (g4454) & (!g4455)) + ((g2891) & (!g2916) & (g2897) & (g2985) & (g4454) & (g4455)) + ((g2891) & (g2916) & (!g2897) & (!g2985) & (!g4454) & (g4455)) + ((g2891) & (g2916) & (!g2897) & (!g2985) & (g4454) & (!g4455)) + ((g2891) & (g2916) & (!g2897) & (!g2985) & (g4454) & (g4455)) + ((g2891) & (g2916) & (!g2897) & (g2985) & (!g4454) & (!g4455)) + ((g2891) & (g2916) & (!g2897) & (g2985) & (!g4454) & (g4455)) + ((g2891) & (g2916) & (!g2897) & (g2985) & (g4454) & (!g4455)) + ((g2891) & (g2916) & (!g2897) & (g2985) & (g4454) & (g4455)) + ((g2891) & (g2916) & (g2897) & (!g2985) & (!g4454) & (!g4455)) + ((g2891) & (g2916) & (g2897) & (!g2985) & (!g4454) & (g4455)) + ((g2891) & (g2916) & (g2897) & (!g2985) & (g4454) & (!g4455)) + ((g2891) & (g2916) & (g2897) & (!g2985) & (g4454) & (g4455)) + ((g2891) & (g2916) & (g2897) & (g2985) & (!g4454) & (!g4455)) + ((g2891) & (g2916) & (g2897) & (g2985) & (!g4454) & (g4455)) + ((g2891) & (g2916) & (g2897) & (g2985) & (g4454) & (!g4455)) + ((g2891) & (g2916) & (g2897) & (g2985) & (g4454) & (g4455)));
	assign g4576 = (((!g2761) & (!g2794) & (!g3359) & (g3389) & (!g4527)) + ((!g2761) & (!g2794) & (!g3359) & (g3389) & (g4527)) + ((!g2761) & (!g2794) & (g3359) & (!g3389) & (g4527)) + ((!g2761) & (!g2794) & (g3359) & (g3389) & (!g4527)) + ((!g2761) & (g2794) & (!g3359) & (!g3389) & (!g4527)) + ((!g2761) & (g2794) & (!g3359) & (!g3389) & (g4527)) + ((!g2761) & (g2794) & (g3359) & (!g3389) & (!g4527)) + ((!g2761) & (g2794) & (g3359) & (g3389) & (g4527)) + ((g2761) & (!g2794) & (!g3359) & (!g3389) & (g4527)) + ((g2761) & (!g2794) & (!g3359) & (g3389) & (!g4527)) + ((g2761) & (!g2794) & (g3359) & (!g3389) & (!g4527)) + ((g2761) & (!g2794) & (g3359) & (!g3389) & (g4527)) + ((g2761) & (g2794) & (!g3359) & (!g3389) & (!g4527)) + ((g2761) & (g2794) & (!g3359) & (g3389) & (g4527)) + ((g2761) & (g2794) & (g3359) & (g3389) & (!g4527)) + ((g2761) & (g2794) & (g3359) & (g3389) & (g4527)));
	assign g4577 = (((!g3345) & (!g3342) & (!g3380) & (g3372) & (!g4528)) + ((!g3345) & (!g3342) & (!g3380) & (g3372) & (g4528)) + ((!g3345) & (!g3342) & (g3380) & (!g3372) & (!g4528)) + ((!g3345) & (!g3342) & (g3380) & (!g3372) & (g4528)) + ((!g3345) & (g3342) & (!g3380) & (!g3372) & (g4528)) + ((!g3345) & (g3342) & (!g3380) & (g3372) & (!g4528)) + ((!g3345) & (g3342) & (g3380) & (!g3372) & (!g4528)) + ((!g3345) & (g3342) & (g3380) & (g3372) & (g4528)) + ((g3345) & (!g3342) & (!g3380) & (!g3372) & (g4528)) + ((g3345) & (!g3342) & (!g3380) & (g3372) & (!g4528)) + ((g3345) & (!g3342) & (g3380) & (!g3372) & (!g4528)) + ((g3345) & (!g3342) & (g3380) & (g3372) & (g4528)) + ((g3345) & (g3342) & (!g3380) & (!g3372) & (!g4528)) + ((g3345) & (g3342) & (!g3380) & (!g3372) & (g4528)) + ((g3345) & (g3342) & (g3380) & (g3372) & (!g4528)) + ((g3345) & (g3342) & (g3380) & (g3372) & (g4528)));
	assign g4578 = (((!g830) & (!g1914) & (!g2329) & (!g4576) & (!g4577) & (key[200])) + ((!g830) & (!g1914) & (!g2329) & (!g4576) & (g4577) & (key[200])) + ((!g830) & (!g1914) & (!g2329) & (g4576) & (!g4577) & (key[200])) + ((!g830) & (!g1914) & (!g2329) & (g4576) & (g4577) & (key[200])) + ((!g830) & (!g1914) & (g2329) & (!g4576) & (!g4577) & (key[200])) + ((!g830) & (!g1914) & (g2329) & (!g4576) & (g4577) & (key[200])) + ((!g830) & (!g1914) & (g2329) & (g4576) & (!g4577) & (key[200])) + ((!g830) & (!g1914) & (g2329) & (g4576) & (g4577) & (key[200])) + ((!g830) & (g1914) & (!g2329) & (!g4576) & (!g4577) & (key[200])) + ((!g830) & (g1914) & (!g2329) & (!g4576) & (g4577) & (key[200])) + ((!g830) & (g1914) & (!g2329) & (g4576) & (!g4577) & (key[200])) + ((!g830) & (g1914) & (!g2329) & (g4576) & (g4577) & (key[200])) + ((!g830) & (g1914) & (g2329) & (!g4576) & (!g4577) & (key[200])) + ((!g830) & (g1914) & (g2329) & (!g4576) & (g4577) & (key[200])) + ((!g830) & (g1914) & (g2329) & (g4576) & (!g4577) & (key[200])) + ((!g830) & (g1914) & (g2329) & (g4576) & (g4577) & (key[200])) + ((g830) & (!g1914) & (!g2329) & (!g4576) & (g4577) & (!key[200])) + ((g830) & (!g1914) & (!g2329) & (!g4576) & (g4577) & (key[200])) + ((g830) & (!g1914) & (!g2329) & (g4576) & (g4577) & (!key[200])) + ((g830) & (!g1914) & (!g2329) & (g4576) & (g4577) & (key[200])) + ((g830) & (!g1914) & (g2329) & (!g4576) & (!g4577) & (!key[200])) + ((g830) & (!g1914) & (g2329) & (!g4576) & (!g4577) & (key[200])) + ((g830) & (!g1914) & (g2329) & (g4576) & (!g4577) & (!key[200])) + ((g830) & (!g1914) & (g2329) & (g4576) & (!g4577) & (key[200])) + ((g830) & (g1914) & (!g2329) & (g4576) & (!g4577) & (!key[200])) + ((g830) & (g1914) & (!g2329) & (g4576) & (!g4577) & (key[200])) + ((g830) & (g1914) & (!g2329) & (g4576) & (g4577) & (!key[200])) + ((g830) & (g1914) & (!g2329) & (g4576) & (g4577) & (key[200])) + ((g830) & (g1914) & (g2329) & (!g4576) & (!g4577) & (!key[200])) + ((g830) & (g1914) & (g2329) & (!g4576) & (!g4577) & (key[200])) + ((g830) & (g1914) & (g2329) & (!g4576) & (g4577) & (!key[200])) + ((g830) & (g1914) & (g2329) & (!g4576) & (g4577) & (key[200])));
	assign g4579 = (((!g1892) & (!g2026) & (!g1900) & (g2028)) + ((!g1892) & (!g2026) & (g1900) & (g2028)) + ((!g1892) & (g2026) & (!g1900) & (!g2028)) + ((!g1892) & (g2026) & (g1900) & (!g2028)) + ((g1892) & (!g2026) & (!g1900) & (g2028)) + ((g1892) & (!g2026) & (g1900) & (!g2028)) + ((g1892) & (g2026) & (!g1900) & (!g2028)) + ((g1892) & (g2026) & (g1900) & (g2028)));
	assign g4580 = (((!g2552) & (!g4503) & (!g4504) & (!g3170)) + ((!g2552) & (!g4503) & (!g4504) & (g3170)) + ((!g2552) & (!g4503) & (g4504) & (!g3170)) + ((!g2552) & (g4503) & (!g4504) & (!g3170)) + ((!g2552) & (g4503) & (g4504) & (!g3170)) + ((g2552) & (!g4503) & (!g4504) & (!g3170)));
	assign g4581 = (((!g1914) & (!g2599) & (!g3202) & (!g4579) & (!g4580)) + ((!g1914) & (!g2599) & (!g3202) & (g4579) & (!g4580)) + ((!g1914) & (!g2599) & (g3202) & (!g4579) & (g4580)) + ((!g1914) & (!g2599) & (g3202) & (g4579) & (g4580)) + ((!g1914) & (g2599) & (!g3202) & (!g4579) & (g4580)) + ((!g1914) & (g2599) & (!g3202) & (g4579) & (g4580)) + ((!g1914) & (g2599) & (g3202) & (!g4579) & (!g4580)) + ((!g1914) & (g2599) & (g3202) & (g4579) & (!g4580)) + ((g1914) & (!g2599) & (!g3202) & (g4579) & (!g4580)) + ((g1914) & (!g2599) & (!g3202) & (g4579) & (g4580)) + ((g1914) & (!g2599) & (g3202) & (g4579) & (!g4580)) + ((g1914) & (!g2599) & (g3202) & (g4579) & (g4580)) + ((g1914) & (g2599) & (!g3202) & (g4579) & (!g4580)) + ((g1914) & (g2599) & (!g3202) & (g4579) & (g4580)) + ((g1914) & (g2599) & (g3202) & (g4579) & (!g4580)) + ((g1914) & (g2599) & (g3202) & (g4579) & (g4580)));
	assign g4582 = (((!g830) & (!g2334) & (!g4581) & (key[136])) + ((!g830) & (!g2334) & (g4581) & (key[136])) + ((!g830) & (g2334) & (!g4581) & (key[136])) + ((!g830) & (g2334) & (g4581) & (key[136])) + ((g830) & (!g2334) & (g4581) & (!key[136])) + ((g830) & (!g2334) & (g4581) & (key[136])) + ((g830) & (g2334) & (!g4581) & (!key[136])) + ((g830) & (g2334) & (!g4581) & (key[136])));
	assign g4583 = (((!g3345) & (!g3333) & (!g3380) & (g3378) & (!g4520)) + ((!g3345) & (!g3333) & (!g3380) & (g3378) & (g4520)) + ((!g3345) & (!g3333) & (g3380) & (!g3378) & (!g4520)) + ((!g3345) & (!g3333) & (g3380) & (!g3378) & (g4520)) + ((!g3345) & (g3333) & (!g3380) & (!g3378) & (g4520)) + ((!g3345) & (g3333) & (!g3380) & (g3378) & (!g4520)) + ((!g3345) & (g3333) & (g3380) & (!g3378) & (!g4520)) + ((!g3345) & (g3333) & (g3380) & (g3378) & (g4520)) + ((g3345) & (!g3333) & (!g3380) & (!g3378) & (g4520)) + ((g3345) & (!g3333) & (!g3380) & (g3378) & (!g4520)) + ((g3345) & (!g3333) & (g3380) & (!g3378) & (!g4520)) + ((g3345) & (!g3333) & (g3380) & (g3378) & (g4520)) + ((g3345) & (g3333) & (!g3380) & (!g3378) & (!g4520)) + ((g3345) & (g3333) & (!g3380) & (!g3378) & (g4520)) + ((g3345) & (g3333) & (g3380) & (g3378) & (!g4520)) + ((g3345) & (g3333) & (g3380) & (g3378) & (g4520)));
	assign g4584 = (((!g2759) & (!g2790) & (!g3359) & (g3389) & (!g4521)) + ((!g2759) & (!g2790) & (!g3359) & (g3389) & (g4521)) + ((!g2759) & (!g2790) & (g3359) & (!g3389) & (g4521)) + ((!g2759) & (!g2790) & (g3359) & (g3389) & (!g4521)) + ((!g2759) & (g2790) & (!g3359) & (!g3389) & (!g4521)) + ((!g2759) & (g2790) & (!g3359) & (!g3389) & (g4521)) + ((!g2759) & (g2790) & (g3359) & (!g3389) & (!g4521)) + ((!g2759) & (g2790) & (g3359) & (g3389) & (g4521)) + ((g2759) & (!g2790) & (!g3359) & (!g3389) & (g4521)) + ((g2759) & (!g2790) & (!g3359) & (g3389) & (!g4521)) + ((g2759) & (!g2790) & (g3359) & (!g3389) & (!g4521)) + ((g2759) & (!g2790) & (g3359) & (!g3389) & (g4521)) + ((g2759) & (g2790) & (!g3359) & (!g3389) & (!g4521)) + ((g2759) & (g2790) & (!g3359) & (g3389) & (g4521)) + ((g2759) & (g2790) & (g3359) & (g3389) & (!g4521)) + ((g2759) & (g2790) & (g3359) & (g3389) & (g4521)));
	assign g4585 = (((!g830) & (!g1914) & (!g2337) & (!g4583) & (!g4584) & (nonce[40])) + ((!g830) & (!g1914) & (!g2337) & (!g4583) & (g4584) & (nonce[40])) + ((!g830) & (!g1914) & (!g2337) & (g4583) & (!g4584) & (nonce[40])) + ((!g830) & (!g1914) & (!g2337) & (g4583) & (g4584) & (nonce[40])) + ((!g830) & (!g1914) & (g2337) & (!g4583) & (!g4584) & (nonce[40])) + ((!g830) & (!g1914) & (g2337) & (!g4583) & (g4584) & (nonce[40])) + ((!g830) & (!g1914) & (g2337) & (g4583) & (!g4584) & (nonce[40])) + ((!g830) & (!g1914) & (g2337) & (g4583) & (g4584) & (nonce[40])) + ((!g830) & (g1914) & (!g2337) & (!g4583) & (!g4584) & (nonce[40])) + ((!g830) & (g1914) & (!g2337) & (!g4583) & (g4584) & (nonce[40])) + ((!g830) & (g1914) & (!g2337) & (g4583) & (!g4584) & (nonce[40])) + ((!g830) & (g1914) & (!g2337) & (g4583) & (g4584) & (nonce[40])) + ((!g830) & (g1914) & (g2337) & (!g4583) & (!g4584) & (nonce[40])) + ((!g830) & (g1914) & (g2337) & (!g4583) & (g4584) & (nonce[40])) + ((!g830) & (g1914) & (g2337) & (g4583) & (!g4584) & (nonce[40])) + ((!g830) & (g1914) & (g2337) & (g4583) & (g4584) & (nonce[40])) + ((g830) & (!g1914) & (!g2337) & (!g4583) & (g4584) & (!nonce[40])) + ((g830) & (!g1914) & (!g2337) & (!g4583) & (g4584) & (nonce[40])) + ((g830) & (!g1914) & (!g2337) & (g4583) & (g4584) & (!nonce[40])) + ((g830) & (!g1914) & (!g2337) & (g4583) & (g4584) & (nonce[40])) + ((g830) & (!g1914) & (g2337) & (!g4583) & (!g4584) & (!nonce[40])) + ((g830) & (!g1914) & (g2337) & (!g4583) & (!g4584) & (nonce[40])) + ((g830) & (!g1914) & (g2337) & (g4583) & (!g4584) & (!nonce[40])) + ((g830) & (!g1914) & (g2337) & (g4583) & (!g4584) & (nonce[40])) + ((g830) & (g1914) & (!g2337) & (g4583) & (!g4584) & (!nonce[40])) + ((g830) & (g1914) & (!g2337) & (g4583) & (!g4584) & (nonce[40])) + ((g830) & (g1914) & (!g2337) & (g4583) & (g4584) & (!nonce[40])) + ((g830) & (g1914) & (!g2337) & (g4583) & (g4584) & (nonce[40])) + ((g830) & (g1914) & (g2337) & (!g4583) & (!g4584) & (!nonce[40])) + ((g830) & (g1914) & (g2337) & (!g4583) & (!g4584) & (nonce[40])) + ((g830) & (g1914) & (g2337) & (!g4583) & (g4584) & (!nonce[40])) + ((g830) & (g1914) & (g2337) & (!g4583) & (g4584) & (nonce[40])));
	assign g4586 = (((!g2979) & (!g3007) & (!g2985) & (g3015) & (!g4531) & (!g4532)) + ((!g2979) & (!g3007) & (!g2985) & (g3015) & (!g4531) & (g4532)) + ((!g2979) & (!g3007) & (!g2985) & (g3015) & (g4531) & (!g4532)) + ((!g2979) & (!g3007) & (!g2985) & (g3015) & (g4531) & (g4532)) + ((!g2979) & (!g3007) & (g2985) & (!g3015) & (!g4531) & (g4532)) + ((!g2979) & (!g3007) & (g2985) & (!g3015) & (g4531) & (!g4532)) + ((!g2979) & (!g3007) & (g2985) & (!g3015) & (g4531) & (g4532)) + ((!g2979) & (!g3007) & (g2985) & (g3015) & (!g4531) & (!g4532)) + ((!g2979) & (g3007) & (!g2985) & (!g3015) & (!g4531) & (!g4532)) + ((!g2979) & (g3007) & (!g2985) & (!g3015) & (!g4531) & (g4532)) + ((!g2979) & (g3007) & (!g2985) & (!g3015) & (g4531) & (!g4532)) + ((!g2979) & (g3007) & (!g2985) & (!g3015) & (g4531) & (g4532)) + ((!g2979) & (g3007) & (g2985) & (!g3015) & (!g4531) & (!g4532)) + ((!g2979) & (g3007) & (g2985) & (g3015) & (!g4531) & (g4532)) + ((!g2979) & (g3007) & (g2985) & (g3015) & (g4531) & (!g4532)) + ((!g2979) & (g3007) & (g2985) & (g3015) & (g4531) & (g4532)) + ((g2979) & (!g3007) & (!g2985) & (!g3015) & (!g4531) & (g4532)) + ((g2979) & (!g3007) & (!g2985) & (!g3015) & (g4531) & (!g4532)) + ((g2979) & (!g3007) & (!g2985) & (!g3015) & (g4531) & (g4532)) + ((g2979) & (!g3007) & (!g2985) & (g3015) & (!g4531) & (!g4532)) + ((g2979) & (!g3007) & (g2985) & (!g3015) & (!g4531) & (!g4532)) + ((g2979) & (!g3007) & (g2985) & (!g3015) & (!g4531) & (g4532)) + ((g2979) & (!g3007) & (g2985) & (!g3015) & (g4531) & (!g4532)) + ((g2979) & (!g3007) & (g2985) & (!g3015) & (g4531) & (g4532)) + ((g2979) & (g3007) & (!g2985) & (!g3015) & (!g4531) & (!g4532)) + ((g2979) & (g3007) & (!g2985) & (g3015) & (!g4531) & (g4532)) + ((g2979) & (g3007) & (!g2985) & (g3015) & (g4531) & (!g4532)) + ((g2979) & (g3007) & (!g2985) & (g3015) & (g4531) & (g4532)) + ((g2979) & (g3007) & (g2985) & (g3015) & (!g4531) & (!g4532)) + ((g2979) & (g3007) & (g2985) & (g3015) & (!g4531) & (g4532)) + ((g2979) & (g3007) & (g2985) & (g3015) & (g4531) & (!g4532)) + ((g2979) & (g3007) & (g2985) & (g3015) & (g4531) & (g4532)));
	assign g4587 = (((!g2900) & (!g2944) & (g2902) & (g2968) & (!g4468) & (g4469)) + ((!g2900) & (!g2944) & (g2902) & (g2968) & (g4468) & (!g4469)) + ((!g2900) & (!g2944) & (g2902) & (g2968) & (g4468) & (g4469)) + ((!g2900) & (g2944) & (!g2902) & (g2968) & (!g4468) & (!g4469)) + ((!g2900) & (g2944) & (!g2902) & (g2968) & (!g4468) & (g4469)) + ((!g2900) & (g2944) & (!g2902) & (g2968) & (g4468) & (!g4469)) + ((!g2900) & (g2944) & (!g2902) & (g2968) & (g4468) & (g4469)) + ((!g2900) & (g2944) & (g2902) & (!g2968) & (!g4468) & (g4469)) + ((!g2900) & (g2944) & (g2902) & (!g2968) & (g4468) & (!g4469)) + ((!g2900) & (g2944) & (g2902) & (!g2968) & (g4468) & (g4469)) + ((!g2900) & (g2944) & (g2902) & (g2968) & (!g4468) & (!g4469)) + ((!g2900) & (g2944) & (g2902) & (g2968) & (!g4468) & (g4469)) + ((!g2900) & (g2944) & (g2902) & (g2968) & (g4468) & (!g4469)) + ((!g2900) & (g2944) & (g2902) & (g2968) & (g4468) & (g4469)) + ((g2900) & (!g2944) & (!g2902) & (g2968) & (!g4468) & (g4469)) + ((g2900) & (!g2944) & (!g2902) & (g2968) & (g4468) & (!g4469)) + ((g2900) & (!g2944) & (!g2902) & (g2968) & (g4468) & (g4469)) + ((g2900) & (!g2944) & (g2902) & (g2968) & (!g4468) & (!g4469)) + ((g2900) & (!g2944) & (g2902) & (g2968) & (!g4468) & (g4469)) + ((g2900) & (!g2944) & (g2902) & (g2968) & (g4468) & (!g4469)) + ((g2900) & (!g2944) & (g2902) & (g2968) & (g4468) & (g4469)) + ((g2900) & (g2944) & (!g2902) & (!g2968) & (!g4468) & (g4469)) + ((g2900) & (g2944) & (!g2902) & (!g2968) & (g4468) & (!g4469)) + ((g2900) & (g2944) & (!g2902) & (!g2968) & (g4468) & (g4469)) + ((g2900) & (g2944) & (!g2902) & (g2968) & (!g4468) & (!g4469)) + ((g2900) & (g2944) & (!g2902) & (g2968) & (!g4468) & (g4469)) + ((g2900) & (g2944) & (!g2902) & (g2968) & (g4468) & (!g4469)) + ((g2900) & (g2944) & (!g2902) & (g2968) & (g4468) & (g4469)) + ((g2900) & (g2944) & (g2902) & (!g2968) & (!g4468) & (!g4469)) + ((g2900) & (g2944) & (g2902) & (!g2968) & (!g4468) & (g4469)) + ((g2900) & (g2944) & (g2902) & (!g2968) & (g4468) & (!g4469)) + ((g2900) & (g2944) & (g2902) & (!g2968) & (g4468) & (g4469)) + ((g2900) & (g2944) & (g2902) & (g2968) & (!g4468) & (!g4469)) + ((g2900) & (g2944) & (g2902) & (g2968) & (!g4468) & (g4469)) + ((g2900) & (g2944) & (g2902) & (g2968) & (g4468) & (!g4469)) + ((g2900) & (g2944) & (g2902) & (g2968) & (g4468) & (g4469)));
	assign g4588 = (((!g1269) & (!g3507) & (!g2559)) + ((!g1269) & (g3507) & (g2559)) + ((g1269) & (!g3507) & (g2559)) + ((g1269) & (g3507) & (!g2559)));
	assign g4589 = (((!g2566) & (!g2589) & (!g3525)) + ((!g2566) & (g2589) & (g3525)) + ((g2566) & (!g2589) & (g3525)) + ((g2566) & (g2589) & (!g3525)));
	assign g4590 = (((!g830) & (!g1914) & (!g2343) & (!g4588) & (!g4589) & (key[54])) + ((!g830) & (!g1914) & (!g2343) & (!g4588) & (g4589) & (key[54])) + ((!g830) & (!g1914) & (!g2343) & (g4588) & (!g4589) & (key[54])) + ((!g830) & (!g1914) & (!g2343) & (g4588) & (g4589) & (key[54])) + ((!g830) & (!g1914) & (g2343) & (!g4588) & (!g4589) & (key[54])) + ((!g830) & (!g1914) & (g2343) & (!g4588) & (g4589) & (key[54])) + ((!g830) & (!g1914) & (g2343) & (g4588) & (!g4589) & (key[54])) + ((!g830) & (!g1914) & (g2343) & (g4588) & (g4589) & (key[54])) + ((!g830) & (g1914) & (!g2343) & (!g4588) & (!g4589) & (key[54])) + ((!g830) & (g1914) & (!g2343) & (!g4588) & (g4589) & (key[54])) + ((!g830) & (g1914) & (!g2343) & (g4588) & (!g4589) & (key[54])) + ((!g830) & (g1914) & (!g2343) & (g4588) & (g4589) & (key[54])) + ((!g830) & (g1914) & (g2343) & (!g4588) & (!g4589) & (key[54])) + ((!g830) & (g1914) & (g2343) & (!g4588) & (g4589) & (key[54])) + ((!g830) & (g1914) & (g2343) & (g4588) & (!g4589) & (key[54])) + ((!g830) & (g1914) & (g2343) & (g4588) & (g4589) & (key[54])) + ((g830) & (!g1914) & (!g2343) & (!g4588) & (g4589) & (!key[54])) + ((g830) & (!g1914) & (!g2343) & (!g4588) & (g4589) & (key[54])) + ((g830) & (!g1914) & (!g2343) & (g4588) & (g4589) & (!key[54])) + ((g830) & (!g1914) & (!g2343) & (g4588) & (g4589) & (key[54])) + ((g830) & (!g1914) & (g2343) & (!g4588) & (!g4589) & (!key[54])) + ((g830) & (!g1914) & (g2343) & (!g4588) & (!g4589) & (key[54])) + ((g830) & (!g1914) & (g2343) & (g4588) & (!g4589) & (!key[54])) + ((g830) & (!g1914) & (g2343) & (g4588) & (!g4589) & (key[54])) + ((g830) & (g1914) & (!g2343) & (g4588) & (!g4589) & (!key[54])) + ((g830) & (g1914) & (!g2343) & (g4588) & (!g4589) & (key[54])) + ((g830) & (g1914) & (!g2343) & (g4588) & (g4589) & (!key[54])) + ((g830) & (g1914) & (!g2343) & (g4588) & (g4589) & (key[54])) + ((g830) & (g1914) & (g2343) & (!g4588) & (!g4589) & (!key[54])) + ((g830) & (g1914) & (g2343) & (!g4588) & (!g4589) & (key[54])) + ((g830) & (g1914) & (g2343) & (!g4588) & (g4589) & (!key[54])) + ((g830) & (g1914) & (g2343) & (!g4588) & (g4589) & (key[54])));
	assign g4591 = (((!g1958) & (g2320) & (!g3749)) + ((g1958) & (!g2320) & (!g3749)) + ((g1958) & (g2320) & (!g3749)) + ((g1958) & (g2320) & (g3749)));
	assign g4592 = (((!g1960) & (!g2350) & (g4591)) + ((!g1960) & (g2350) & (!g4591)) + ((g1960) & (!g2350) & (!g4591)) + ((g1960) & (g2350) & (g4591)));
	assign g4593 = (((!g830) & (!g2344) & (!g6627) & (key[86])) + ((!g830) & (!g2344) & (g6627) & (key[86])) + ((!g830) & (g2344) & (!g6627) & (key[86])) + ((!g830) & (g2344) & (g6627) & (key[86])) + ((g830) & (!g2344) & (g6627) & (!key[86])) + ((g830) & (!g2344) & (g6627) & (key[86])) + ((g830) & (g2344) & (!g6627) & (!key[86])) + ((g830) & (g2344) & (!g6627) & (key[86])));
	assign g4594 = (((!g3400) & (!g2566) & (!g2572)) + ((!g3400) & (g2566) & (g2572)) + ((g3400) & (!g2566) & (g2572)) + ((g3400) & (g2566) & (!g2572)));
	assign g4595 = (((!g1269) & (!g3417) & (!g2575)) + ((!g1269) & (g3417) & (g2575)) + ((g1269) & (!g3417) & (g2575)) + ((g1269) & (g3417) & (!g2575)));
	assign g8307 = (((!g5560) & (g5603) & (!g4596)) + ((!g5560) & (g5603) & (g4596)) + ((g5560) & (!g5603) & (g4596)) + ((g5560) & (g5603) & (g4596)));
	assign g4597 = (((!g830) & (!g1914) & (!g2347) & (!g4594) & (!g4595) & (g4596)) + ((!g830) & (!g1914) & (!g2347) & (!g4594) & (g4595) & (g4596)) + ((!g830) & (!g1914) & (!g2347) & (g4594) & (!g4595) & (g4596)) + ((!g830) & (!g1914) & (!g2347) & (g4594) & (g4595) & (g4596)) + ((!g830) & (!g1914) & (g2347) & (!g4594) & (!g4595) & (g4596)) + ((!g830) & (!g1914) & (g2347) & (!g4594) & (g4595) & (g4596)) + ((!g830) & (!g1914) & (g2347) & (g4594) & (!g4595) & (g4596)) + ((!g830) & (!g1914) & (g2347) & (g4594) & (g4595) & (g4596)) + ((!g830) & (g1914) & (!g2347) & (!g4594) & (!g4595) & (g4596)) + ((!g830) & (g1914) & (!g2347) & (!g4594) & (g4595) & (g4596)) + ((!g830) & (g1914) & (!g2347) & (g4594) & (!g4595) & (g4596)) + ((!g830) & (g1914) & (!g2347) & (g4594) & (g4595) & (g4596)) + ((!g830) & (g1914) & (g2347) & (!g4594) & (!g4595) & (g4596)) + ((!g830) & (g1914) & (g2347) & (!g4594) & (g4595) & (g4596)) + ((!g830) & (g1914) & (g2347) & (g4594) & (!g4595) & (g4596)) + ((!g830) & (g1914) & (g2347) & (g4594) & (g4595) & (g4596)) + ((g830) & (!g1914) & (!g2347) & (!g4594) & (g4595) & (!g4596)) + ((g830) & (!g1914) & (!g2347) & (!g4594) & (g4595) & (g4596)) + ((g830) & (!g1914) & (!g2347) & (g4594) & (g4595) & (!g4596)) + ((g830) & (!g1914) & (!g2347) & (g4594) & (g4595) & (g4596)) + ((g830) & (!g1914) & (g2347) & (!g4594) & (!g4595) & (!g4596)) + ((g830) & (!g1914) & (g2347) & (!g4594) & (!g4595) & (g4596)) + ((g830) & (!g1914) & (g2347) & (g4594) & (!g4595) & (!g4596)) + ((g830) & (!g1914) & (g2347) & (g4594) & (!g4595) & (g4596)) + ((g830) & (g1914) & (!g2347) & (g4594) & (!g4595) & (!g4596)) + ((g830) & (g1914) & (!g2347) & (g4594) & (!g4595) & (g4596)) + ((g830) & (g1914) & (!g2347) & (g4594) & (g4595) & (!g4596)) + ((g830) & (g1914) & (!g2347) & (g4594) & (g4595) & (g4596)) + ((g830) & (g1914) & (g2347) & (!g4594) & (!g4595) & (!g4596)) + ((g830) & (g1914) & (g2347) & (!g4594) & (!g4595) & (g4596)) + ((g830) & (g1914) & (g2347) & (!g4594) & (g4595) & (!g4596)) + ((g830) & (g1914) & (g2347) & (!g4594) & (g4595) & (g4596)));
	assign g4598 = (((!g1996) & (g2304) & (!g3487)) + ((g1996) & (!g2304) & (!g3487)) + ((g1996) & (g2304) & (!g3487)) + ((g1996) & (g2304) & (g3487)));
	assign g4599 = (((!g1998) & (!g2360) & (g4598)) + ((!g1998) & (g2360) & (!g4598)) + ((g1998) & (!g2360) & (!g4598)) + ((g1998) & (g2360) & (g4598)));
	assign g4600 = (((!g830) & (!g2348) & (!g6616) & (key[182])) + ((!g830) & (!g2348) & (g6616) & (key[182])) + ((!g830) & (g2348) & (!g6616) & (key[182])) + ((!g830) & (g2348) & (g6616) & (key[182])) + ((g830) & (!g2348) & (g6616) & (!key[182])) + ((g830) & (!g2348) & (g6616) & (key[182])) + ((g830) & (g2348) & (!g6616) & (!key[182])) + ((g830) & (g2348) & (!g6616) & (key[182])));
	assign g4601 = (((!g1906) & (!g1940) & (!g1942) & (!g828) & (!g864) & (g897)) + ((!g1906) & (!g1940) & (!g1942) & (!g828) & (g864) & (g897)) + ((!g1906) & (!g1940) & (!g1942) & (g828) & (!g864) & (g897)) + ((!g1906) & (!g1940) & (!g1942) & (g828) & (g864) & (g897)) + ((!g1906) & (!g1940) & (g1942) & (!g828) & (!g864) & (!g897)) + ((!g1906) & (!g1940) & (g1942) & (!g828) & (g864) & (!g897)) + ((!g1906) & (!g1940) & (g1942) & (g828) & (!g864) & (!g897)) + ((!g1906) & (!g1940) & (g1942) & (g828) & (g864) & (!g897)) + ((!g1906) & (g1940) & (!g1942) & (!g828) & (!g864) & (g897)) + ((!g1906) & (g1940) & (!g1942) & (!g828) & (g864) & (!g897)) + ((!g1906) & (g1940) & (!g1942) & (g828) & (!g864) & (g897)) + ((!g1906) & (g1940) & (!g1942) & (g828) & (g864) & (!g897)) + ((!g1906) & (g1940) & (g1942) & (!g828) & (!g864) & (!g897)) + ((!g1906) & (g1940) & (g1942) & (!g828) & (g864) & (g897)) + ((!g1906) & (g1940) & (g1942) & (g828) & (!g864) & (!g897)) + ((!g1906) & (g1940) & (g1942) & (g828) & (g864) & (g897)) + ((g1906) & (!g1940) & (!g1942) & (!g828) & (!g864) & (g897)) + ((g1906) & (!g1940) & (!g1942) & (!g828) & (g864) & (g897)) + ((g1906) & (!g1940) & (!g1942) & (g828) & (!g864) & (g897)) + ((g1906) & (!g1940) & (!g1942) & (g828) & (g864) & (!g897)) + ((g1906) & (!g1940) & (g1942) & (!g828) & (!g864) & (!g897)) + ((g1906) & (!g1940) & (g1942) & (!g828) & (g864) & (!g897)) + ((g1906) & (!g1940) & (g1942) & (g828) & (!g864) & (!g897)) + ((g1906) & (!g1940) & (g1942) & (g828) & (g864) & (g897)) + ((g1906) & (g1940) & (!g1942) & (!g828) & (!g864) & (g897)) + ((g1906) & (g1940) & (!g1942) & (!g828) & (g864) & (!g897)) + ((g1906) & (g1940) & (!g1942) & (g828) & (!g864) & (!g897)) + ((g1906) & (g1940) & (!g1942) & (g828) & (g864) & (!g897)) + ((g1906) & (g1940) & (g1942) & (!g828) & (!g864) & (!g897)) + ((g1906) & (g1940) & (g1942) & (!g828) & (g864) & (g897)) + ((g1906) & (g1940) & (g1942) & (g828) & (!g864) & (g897)) + ((g1906) & (g1940) & (g1942) & (g828) & (g864) & (g897)));
	assign g4602 = (((!g3161) & (!g3187) & (!g4488) & (!g4489) & (!g3165) & (!g3210)) + ((!g3161) & (!g3187) & (!g4488) & (!g4489) & (!g3165) & (g3210)) + ((!g3161) & (!g3187) & (!g4488) & (!g4489) & (g3165) & (!g3210)) + ((!g3161) & (!g3187) & (!g4488) & (!g4489) & (g3165) & (g3210)) + ((!g3161) & (!g3187) & (!g4488) & (g4489) & (!g3165) & (!g3210)) + ((!g3161) & (!g3187) & (!g4488) & (g4489) & (!g3165) & (g3210)) + ((!g3161) & (!g3187) & (!g4488) & (g4489) & (g3165) & (!g3210)) + ((!g3161) & (!g3187) & (g4488) & (!g4489) & (!g3165) & (!g3210)) + ((!g3161) & (!g3187) & (g4488) & (!g4489) & (!g3165) & (g3210)) + ((!g3161) & (!g3187) & (g4488) & (!g4489) & (g3165) & (!g3210)) + ((!g3161) & (!g3187) & (g4488) & (g4489) & (!g3165) & (!g3210)) + ((!g3161) & (!g3187) & (g4488) & (g4489) & (!g3165) & (g3210)) + ((!g3161) & (!g3187) & (g4488) & (g4489) & (g3165) & (!g3210)) + ((!g3161) & (g3187) & (!g4488) & (!g4489) & (!g3165) & (!g3210)) + ((!g3161) & (g3187) & (!g4488) & (!g4489) & (g3165) & (!g3210)) + ((!g3161) & (g3187) & (!g4488) & (g4489) & (!g3165) & (!g3210)) + ((!g3161) & (g3187) & (g4488) & (!g4489) & (!g3165) & (!g3210)) + ((!g3161) & (g3187) & (g4488) & (g4489) & (!g3165) & (!g3210)) + ((g3161) & (!g3187) & (!g4488) & (!g4489) & (!g3165) & (!g3210)) + ((g3161) & (!g3187) & (!g4488) & (!g4489) & (!g3165) & (g3210)) + ((g3161) & (!g3187) & (!g4488) & (!g4489) & (g3165) & (!g3210)) + ((g3161) & (!g3187) & (!g4488) & (g4489) & (!g3165) & (!g3210)) + ((g3161) & (!g3187) & (!g4488) & (g4489) & (g3165) & (!g3210)) + ((g3161) & (!g3187) & (g4488) & (!g4489) & (!g3165) & (!g3210)) + ((g3161) & (!g3187) & (g4488) & (!g4489) & (g3165) & (!g3210)) + ((g3161) & (!g3187) & (g4488) & (g4489) & (!g3165) & (!g3210)) + ((g3161) & (!g3187) & (g4488) & (g4489) & (g3165) & (!g3210)) + ((g3161) & (g3187) & (!g4488) & (!g4489) & (!g3165) & (!g3210)));
	assign g4603 = (((!g1914) & (!g3255) & (!g4601) & (!g4602) & (!g3265)) + ((!g1914) & (!g3255) & (!g4601) & (g4602) & (g3265)) + ((!g1914) & (!g3255) & (g4601) & (!g4602) & (!g3265)) + ((!g1914) & (!g3255) & (g4601) & (g4602) & (g3265)) + ((!g1914) & (g3255) & (!g4601) & (!g4602) & (g3265)) + ((!g1914) & (g3255) & (!g4601) & (g4602) & (!g3265)) + ((!g1914) & (g3255) & (g4601) & (!g4602) & (g3265)) + ((!g1914) & (g3255) & (g4601) & (g4602) & (!g3265)) + ((g1914) & (!g3255) & (g4601) & (!g4602) & (!g3265)) + ((g1914) & (!g3255) & (g4601) & (!g4602) & (g3265)) + ((g1914) & (!g3255) & (g4601) & (g4602) & (!g3265)) + ((g1914) & (!g3255) & (g4601) & (g4602) & (g3265)) + ((g1914) & (g3255) & (g4601) & (!g4602) & (!g3265)) + ((g1914) & (g3255) & (g4601) & (!g4602) & (g3265)) + ((g1914) & (g3255) & (g4601) & (g4602) & (!g3265)) + ((g1914) & (g3255) & (g4601) & (g4602) & (g3265)));
	assign g4604 = (((!g830) & (!g2350) & (!g4603) & (key[9])) + ((!g830) & (!g2350) & (g4603) & (key[9])) + ((!g830) & (g2350) & (!g4603) & (key[9])) + ((!g830) & (g2350) & (g4603) & (key[9])) + ((g830) & (!g2350) & (g4603) & (!key[9])) + ((g830) & (!g2350) & (g4603) & (key[9])) + ((g830) & (g2350) & (!g4603) & (!key[9])) + ((g830) & (g2350) & (!g4603) & (key[9])));
	assign g4605 = (((!g2298) & (!g2347) & (g2938) & (g3011) & (!g4492) & (g4493)) + ((!g2298) & (!g2347) & (g2938) & (g3011) & (g4492) & (!g4493)) + ((!g2298) & (!g2347) & (g2938) & (g3011) & (g4492) & (g4493)) + ((!g2298) & (g2347) & (!g2938) & (g3011) & (!g4492) & (!g4493)) + ((!g2298) & (g2347) & (!g2938) & (g3011) & (!g4492) & (g4493)) + ((!g2298) & (g2347) & (!g2938) & (g3011) & (g4492) & (!g4493)) + ((!g2298) & (g2347) & (!g2938) & (g3011) & (g4492) & (g4493)) + ((!g2298) & (g2347) & (g2938) & (!g3011) & (!g4492) & (g4493)) + ((!g2298) & (g2347) & (g2938) & (!g3011) & (g4492) & (!g4493)) + ((!g2298) & (g2347) & (g2938) & (!g3011) & (g4492) & (g4493)) + ((!g2298) & (g2347) & (g2938) & (g3011) & (!g4492) & (!g4493)) + ((!g2298) & (g2347) & (g2938) & (g3011) & (!g4492) & (g4493)) + ((!g2298) & (g2347) & (g2938) & (g3011) & (g4492) & (!g4493)) + ((!g2298) & (g2347) & (g2938) & (g3011) & (g4492) & (g4493)) + ((g2298) & (!g2347) & (!g2938) & (g3011) & (!g4492) & (g4493)) + ((g2298) & (!g2347) & (!g2938) & (g3011) & (g4492) & (!g4493)) + ((g2298) & (!g2347) & (!g2938) & (g3011) & (g4492) & (g4493)) + ((g2298) & (!g2347) & (g2938) & (g3011) & (!g4492) & (!g4493)) + ((g2298) & (!g2347) & (g2938) & (g3011) & (!g4492) & (g4493)) + ((g2298) & (!g2347) & (g2938) & (g3011) & (g4492) & (!g4493)) + ((g2298) & (!g2347) & (g2938) & (g3011) & (g4492) & (g4493)) + ((g2298) & (g2347) & (!g2938) & (!g3011) & (!g4492) & (g4493)) + ((g2298) & (g2347) & (!g2938) & (!g3011) & (g4492) & (!g4493)) + ((g2298) & (g2347) & (!g2938) & (!g3011) & (g4492) & (g4493)) + ((g2298) & (g2347) & (!g2938) & (g3011) & (!g4492) & (!g4493)) + ((g2298) & (g2347) & (!g2938) & (g3011) & (!g4492) & (g4493)) + ((g2298) & (g2347) & (!g2938) & (g3011) & (g4492) & (!g4493)) + ((g2298) & (g2347) & (!g2938) & (g3011) & (g4492) & (g4493)) + ((g2298) & (g2347) & (g2938) & (!g3011) & (!g4492) & (!g4493)) + ((g2298) & (g2347) & (g2938) & (!g3011) & (!g4492) & (g4493)) + ((g2298) & (g2347) & (g2938) & (!g3011) & (g4492) & (!g4493)) + ((g2298) & (g2347) & (g2938) & (!g3011) & (g4492) & (g4493)) + ((g2298) & (g2347) & (g2938) & (g3011) & (!g4492) & (!g4493)) + ((g2298) & (g2347) & (g2938) & (g3011) & (!g4492) & (g4493)) + ((g2298) & (g2347) & (g2938) & (g3011) & (g4492) & (!g4493)) + ((g2298) & (g2347) & (g2938) & (g3011) & (g4492) & (g4493)));
	assign g4606 = (((!g2343) & (!g2376) & (!g3005) & (g3050) & (!g4556)) + ((!g2343) & (!g2376) & (!g3005) & (g3050) & (g4556)) + ((!g2343) & (!g2376) & (g3005) & (!g3050) & (g4556)) + ((!g2343) & (!g2376) & (g3005) & (g3050) & (!g4556)) + ((!g2343) & (g2376) & (!g3005) & (!g3050) & (!g4556)) + ((!g2343) & (g2376) & (!g3005) & (!g3050) & (g4556)) + ((!g2343) & (g2376) & (g3005) & (!g3050) & (!g4556)) + ((!g2343) & (g2376) & (g3005) & (g3050) & (g4556)) + ((g2343) & (!g2376) & (!g3005) & (!g3050) & (g4556)) + ((g2343) & (!g2376) & (!g3005) & (g3050) & (!g4556)) + ((g2343) & (!g2376) & (g3005) & (!g3050) & (!g4556)) + ((g2343) & (!g2376) & (g3005) & (!g3050) & (g4556)) + ((g2343) & (g2376) & (!g3005) & (!g3050) & (!g4556)) + ((g2343) & (g2376) & (!g3005) & (g3050) & (g4556)) + ((g2343) & (g2376) & (g3005) & (g3050) & (!g4556)) + ((g2343) & (g2376) & (g3005) & (g3050) & (g4556)));
	assign g4607 = (((!g2555) & (!g2601) & (!g3168) & (!g3190) & (!g4498) & (!g4499)) + ((!g2555) & (!g2601) & (!g3168) & (!g3190) & (!g4498) & (g4499)) + ((!g2555) & (!g2601) & (!g3168) & (!g3190) & (g4498) & (!g4499)) + ((!g2555) & (!g2601) & (!g3168) & (!g3190) & (g4498) & (g4499)) + ((!g2555) & (!g2601) & (!g3168) & (g3190) & (!g4498) & (!g4499)) + ((!g2555) & (!g2601) & (!g3168) & (g3190) & (!g4498) & (g4499)) + ((!g2555) & (!g2601) & (!g3168) & (g3190) & (g4498) & (!g4499)) + ((!g2555) & (!g2601) & (!g3168) & (g3190) & (g4498) & (g4499)) + ((!g2555) & (!g2601) & (g3168) & (!g3190) & (!g4498) & (!g4499)) + ((!g2555) & (!g2601) & (g3168) & (!g3190) & (!g4498) & (g4499)) + ((!g2555) & (!g2601) & (g3168) & (!g3190) & (g4498) & (!g4499)) + ((!g2555) & (!g2601) & (g3168) & (!g3190) & (g4498) & (g4499)) + ((!g2555) & (!g2601) & (g3168) & (g3190) & (!g4498) & (!g4499)) + ((!g2555) & (g2601) & (!g3168) & (!g3190) & (!g4498) & (!g4499)) + ((!g2555) & (g2601) & (!g3168) & (!g3190) & (!g4498) & (g4499)) + ((!g2555) & (g2601) & (!g3168) & (!g3190) & (g4498) & (!g4499)) + ((!g2555) & (g2601) & (!g3168) & (!g3190) & (g4498) & (g4499)) + ((!g2555) & (g2601) & (g3168) & (!g3190) & (!g4498) & (!g4499)) + ((g2555) & (!g2601) & (!g3168) & (!g3190) & (!g4498) & (!g4499)) + ((g2555) & (!g2601) & (!g3168) & (!g3190) & (!g4498) & (g4499)) + ((g2555) & (!g2601) & (!g3168) & (!g3190) & (g4498) & (!g4499)) + ((g2555) & (!g2601) & (!g3168) & (!g3190) & (g4498) & (g4499)) + ((g2555) & (!g2601) & (!g3168) & (g3190) & (!g4498) & (!g4499)) + ((g2555) & (!g2601) & (g3168) & (!g3190) & (!g4498) & (!g4499)) + ((g2555) & (!g2601) & (g3168) & (!g3190) & (!g4498) & (g4499)) + ((g2555) & (!g2601) & (g3168) & (!g3190) & (g4498) & (!g4499)) + ((g2555) & (!g2601) & (g3168) & (!g3190) & (g4498) & (g4499)) + ((g2555) & (g2601) & (!g3168) & (!g3190) & (!g4498) & (!g4499)));
	assign g4608 = (((!g1898) & (!g2022) & (!g2071) & (!g1902) & (!g2036) & (g2077)) + ((!g1898) & (!g2022) & (!g2071) & (!g1902) & (g2036) & (g2077)) + ((!g1898) & (!g2022) & (!g2071) & (g1902) & (!g2036) & (g2077)) + ((!g1898) & (!g2022) & (!g2071) & (g1902) & (g2036) & (g2077)) + ((!g1898) & (!g2022) & (g2071) & (!g1902) & (!g2036) & (!g2077)) + ((!g1898) & (!g2022) & (g2071) & (!g1902) & (g2036) & (!g2077)) + ((!g1898) & (!g2022) & (g2071) & (g1902) & (!g2036) & (!g2077)) + ((!g1898) & (!g2022) & (g2071) & (g1902) & (g2036) & (!g2077)) + ((!g1898) & (g2022) & (!g2071) & (!g1902) & (!g2036) & (g2077)) + ((!g1898) & (g2022) & (!g2071) & (!g1902) & (g2036) & (!g2077)) + ((!g1898) & (g2022) & (!g2071) & (g1902) & (!g2036) & (g2077)) + ((!g1898) & (g2022) & (!g2071) & (g1902) & (g2036) & (!g2077)) + ((!g1898) & (g2022) & (g2071) & (!g1902) & (!g2036) & (!g2077)) + ((!g1898) & (g2022) & (g2071) & (!g1902) & (g2036) & (g2077)) + ((!g1898) & (g2022) & (g2071) & (g1902) & (!g2036) & (!g2077)) + ((!g1898) & (g2022) & (g2071) & (g1902) & (g2036) & (g2077)) + ((g1898) & (!g2022) & (!g2071) & (!g1902) & (!g2036) & (g2077)) + ((g1898) & (!g2022) & (!g2071) & (!g1902) & (g2036) & (g2077)) + ((g1898) & (!g2022) & (!g2071) & (g1902) & (!g2036) & (g2077)) + ((g1898) & (!g2022) & (!g2071) & (g1902) & (g2036) & (!g2077)) + ((g1898) & (!g2022) & (g2071) & (!g1902) & (!g2036) & (!g2077)) + ((g1898) & (!g2022) & (g2071) & (!g1902) & (g2036) & (!g2077)) + ((g1898) & (!g2022) & (g2071) & (g1902) & (!g2036) & (!g2077)) + ((g1898) & (!g2022) & (g2071) & (g1902) & (g2036) & (g2077)) + ((g1898) & (g2022) & (!g2071) & (!g1902) & (!g2036) & (g2077)) + ((g1898) & (g2022) & (!g2071) & (!g1902) & (g2036) & (!g2077)) + ((g1898) & (g2022) & (!g2071) & (g1902) & (!g2036) & (!g2077)) + ((g1898) & (g2022) & (!g2071) & (g1902) & (g2036) & (!g2077)) + ((g1898) & (g2022) & (g2071) & (!g1902) & (!g2036) & (!g2077)) + ((g1898) & (g2022) & (g2071) & (!g1902) & (g2036) & (g2077)) + ((g1898) & (g2022) & (g2071) & (g1902) & (!g2036) & (g2077)) + ((g1898) & (g2022) & (g2071) & (g1902) & (g2036) & (g2077)));
	assign g4609 = (((!g1914) & (!g2649) & (!g3274) & (!g4607) & (g4608)) + ((!g1914) & (!g2649) & (!g3274) & (g4607) & (g4608)) + ((!g1914) & (!g2649) & (g3274) & (!g4607) & (g4608)) + ((!g1914) & (!g2649) & (g3274) & (g4607) & (g4608)) + ((!g1914) & (g2649) & (!g3274) & (!g4607) & (g4608)) + ((!g1914) & (g2649) & (!g3274) & (g4607) & (g4608)) + ((!g1914) & (g2649) & (g3274) & (!g4607) & (g4608)) + ((!g1914) & (g2649) & (g3274) & (g4607) & (g4608)) + ((g1914) & (!g2649) & (!g3274) & (!g4607) & (!g4608)) + ((g1914) & (!g2649) & (!g3274) & (!g4607) & (g4608)) + ((g1914) & (!g2649) & (g3274) & (g4607) & (!g4608)) + ((g1914) & (!g2649) & (g3274) & (g4607) & (g4608)) + ((g1914) & (g2649) & (!g3274) & (g4607) & (!g4608)) + ((g1914) & (g2649) & (!g3274) & (g4607) & (g4608)) + ((g1914) & (g2649) & (g3274) & (!g4607) & (!g4608)) + ((g1914) & (g2649) & (g3274) & (!g4607) & (g4608)));
	assign g8308 = (((!g5560) & (g5605) & (!g4610)) + ((!g5560) & (g5605) & (g4610)) + ((g5560) & (!g5605) & (g4610)) + ((g5560) & (g5605) & (g4610)));
	assign g4611 = (((!g830) & (!g2356) & (!g4609) & (g4610)) + ((!g830) & (!g2356) & (g4609) & (g4610)) + ((!g830) & (g2356) & (!g4609) & (g4610)) + ((!g830) & (g2356) & (g4609) & (g4610)) + ((g830) & (!g2356) & (g4609) & (!g4610)) + ((g830) & (!g2356) & (g4609) & (g4610)) + ((g830) & (g2356) & (!g4609) & (!g4610)) + ((g830) & (g2356) & (!g4609) & (g4610)));
	assign g4612 = (((!g1892) & (!g2026) & (!g2062) & (!g1900) & (!g2028) & (g2074)) + ((!g1892) & (!g2026) & (!g2062) & (!g1900) & (g2028) & (g2074)) + ((!g1892) & (!g2026) & (!g2062) & (g1900) & (!g2028) & (g2074)) + ((!g1892) & (!g2026) & (!g2062) & (g1900) & (g2028) & (g2074)) + ((!g1892) & (!g2026) & (g2062) & (!g1900) & (!g2028) & (!g2074)) + ((!g1892) & (!g2026) & (g2062) & (!g1900) & (g2028) & (!g2074)) + ((!g1892) & (!g2026) & (g2062) & (g1900) & (!g2028) & (!g2074)) + ((!g1892) & (!g2026) & (g2062) & (g1900) & (g2028) & (!g2074)) + ((!g1892) & (g2026) & (!g2062) & (!g1900) & (!g2028) & (g2074)) + ((!g1892) & (g2026) & (!g2062) & (!g1900) & (g2028) & (!g2074)) + ((!g1892) & (g2026) & (!g2062) & (g1900) & (!g2028) & (g2074)) + ((!g1892) & (g2026) & (!g2062) & (g1900) & (g2028) & (!g2074)) + ((!g1892) & (g2026) & (g2062) & (!g1900) & (!g2028) & (!g2074)) + ((!g1892) & (g2026) & (g2062) & (!g1900) & (g2028) & (g2074)) + ((!g1892) & (g2026) & (g2062) & (g1900) & (!g2028) & (!g2074)) + ((!g1892) & (g2026) & (g2062) & (g1900) & (g2028) & (g2074)) + ((g1892) & (!g2026) & (!g2062) & (!g1900) & (!g2028) & (g2074)) + ((g1892) & (!g2026) & (!g2062) & (!g1900) & (g2028) & (g2074)) + ((g1892) & (!g2026) & (!g2062) & (g1900) & (!g2028) & (g2074)) + ((g1892) & (!g2026) & (!g2062) & (g1900) & (g2028) & (!g2074)) + ((g1892) & (!g2026) & (g2062) & (!g1900) & (!g2028) & (!g2074)) + ((g1892) & (!g2026) & (g2062) & (!g1900) & (g2028) & (!g2074)) + ((g1892) & (!g2026) & (g2062) & (g1900) & (!g2028) & (!g2074)) + ((g1892) & (!g2026) & (g2062) & (g1900) & (g2028) & (g2074)) + ((g1892) & (g2026) & (!g2062) & (!g1900) & (!g2028) & (g2074)) + ((g1892) & (g2026) & (!g2062) & (!g1900) & (g2028) & (!g2074)) + ((g1892) & (g2026) & (!g2062) & (g1900) & (!g2028) & (!g2074)) + ((g1892) & (g2026) & (!g2062) & (g1900) & (g2028) & (!g2074)) + ((g1892) & (g2026) & (g2062) & (!g1900) & (!g2028) & (!g2074)) + ((g1892) & (g2026) & (g2062) & (!g1900) & (g2028) & (g2074)) + ((g1892) & (g2026) & (g2062) & (g1900) & (!g2028) & (g2074)) + ((g1892) & (g2026) & (g2062) & (g1900) & (g2028) & (g2074)));
	assign g4613 = (((!g2552) & (!g2599) & (!g4503) & (!g4504) & (!g3170) & (!g3202)) + ((!g2552) & (!g2599) & (!g4503) & (!g4504) & (!g3170) & (g3202)) + ((!g2552) & (!g2599) & (!g4503) & (!g4504) & (g3170) & (!g3202)) + ((!g2552) & (!g2599) & (!g4503) & (!g4504) & (g3170) & (g3202)) + ((!g2552) & (!g2599) & (!g4503) & (g4504) & (!g3170) & (!g3202)) + ((!g2552) & (!g2599) & (!g4503) & (g4504) & (!g3170) & (g3202)) + ((!g2552) & (!g2599) & (!g4503) & (g4504) & (g3170) & (!g3202)) + ((!g2552) & (!g2599) & (g4503) & (!g4504) & (!g3170) & (!g3202)) + ((!g2552) & (!g2599) & (g4503) & (!g4504) & (!g3170) & (g3202)) + ((!g2552) & (!g2599) & (g4503) & (!g4504) & (g3170) & (!g3202)) + ((!g2552) & (!g2599) & (g4503) & (g4504) & (!g3170) & (!g3202)) + ((!g2552) & (!g2599) & (g4503) & (g4504) & (!g3170) & (g3202)) + ((!g2552) & (!g2599) & (g4503) & (g4504) & (g3170) & (!g3202)) + ((!g2552) & (g2599) & (!g4503) & (!g4504) & (!g3170) & (!g3202)) + ((!g2552) & (g2599) & (!g4503) & (!g4504) & (g3170) & (!g3202)) + ((!g2552) & (g2599) & (!g4503) & (g4504) & (!g3170) & (!g3202)) + ((!g2552) & (g2599) & (g4503) & (!g4504) & (!g3170) & (!g3202)) + ((!g2552) & (g2599) & (g4503) & (g4504) & (!g3170) & (!g3202)) + ((g2552) & (!g2599) & (!g4503) & (!g4504) & (!g3170) & (!g3202)) + ((g2552) & (!g2599) & (!g4503) & (!g4504) & (!g3170) & (g3202)) + ((g2552) & (!g2599) & (!g4503) & (!g4504) & (g3170) & (!g3202)) + ((g2552) & (!g2599) & (!g4503) & (g4504) & (!g3170) & (!g3202)) + ((g2552) & (!g2599) & (!g4503) & (g4504) & (g3170) & (!g3202)) + ((g2552) & (!g2599) & (g4503) & (!g4504) & (!g3170) & (!g3202)) + ((g2552) & (!g2599) & (g4503) & (!g4504) & (g3170) & (!g3202)) + ((g2552) & (!g2599) & (g4503) & (g4504) & (!g3170) & (!g3202)) + ((g2552) & (!g2599) & (g4503) & (g4504) & (g3170) & (!g3202)) + ((g2552) & (g2599) & (!g4503) & (!g4504) & (!g3170) & (!g3202)));
	assign g4614 = (((!g1914) & (!g2648) & (!g4612) & (!g4613) & (!g3279)) + ((!g1914) & (!g2648) & (!g4612) & (g4613) & (g3279)) + ((!g1914) & (!g2648) & (g4612) & (!g4613) & (!g3279)) + ((!g1914) & (!g2648) & (g4612) & (g4613) & (g3279)) + ((!g1914) & (g2648) & (!g4612) & (!g4613) & (g3279)) + ((!g1914) & (g2648) & (!g4612) & (g4613) & (!g3279)) + ((!g1914) & (g2648) & (g4612) & (!g4613) & (g3279)) + ((!g1914) & (g2648) & (g4612) & (g4613) & (!g3279)) + ((g1914) & (!g2648) & (g4612) & (!g4613) & (!g3279)) + ((g1914) & (!g2648) & (g4612) & (!g4613) & (g3279)) + ((g1914) & (!g2648) & (g4612) & (g4613) & (!g3279)) + ((g1914) & (!g2648) & (g4612) & (g4613) & (g3279)) + ((g1914) & (g2648) & (g4612) & (!g4613) & (!g3279)) + ((g1914) & (g2648) & (g4612) & (!g4613) & (g3279)) + ((g1914) & (g2648) & (g4612) & (g4613) & (!g3279)) + ((g1914) & (g2648) & (g4612) & (g4613) & (g3279)));
	assign g4615 = (((!g830) & (!g2358) & (!g4614) & (key[137])) + ((!g830) & (!g2358) & (g4614) & (key[137])) + ((!g830) & (g2358) & (!g4614) & (key[137])) + ((!g830) & (g2358) & (g4614) & (key[137])) + ((g830) & (!g2358) & (g4614) & (!key[137])) + ((g830) & (!g2358) & (g4614) & (key[137])) + ((g830) & (g2358) & (!g4614) & (!key[137])) + ((g830) & (g2358) & (!g4614) & (key[137])));
	assign g4616 = (((!g3155) & (!g3196) & (!g3170) & (!g4507) & (!g4508) & (!g3202)) + ((!g3155) & (!g3196) & (!g3170) & (!g4507) & (!g4508) & (g3202)) + ((!g3155) & (!g3196) & (!g3170) & (!g4507) & (g4508) & (!g3202)) + ((!g3155) & (!g3196) & (!g3170) & (!g4507) & (g4508) & (g3202)) + ((!g3155) & (!g3196) & (!g3170) & (g4507) & (!g4508) & (!g3202)) + ((!g3155) & (!g3196) & (!g3170) & (g4507) & (!g4508) & (g3202)) + ((!g3155) & (!g3196) & (!g3170) & (g4507) & (g4508) & (!g3202)) + ((!g3155) & (!g3196) & (!g3170) & (g4507) & (g4508) & (g3202)) + ((!g3155) & (!g3196) & (g3170) & (!g4507) & (!g4508) & (!g3202)) + ((!g3155) & (!g3196) & (g3170) & (!g4507) & (!g4508) & (g3202)) + ((!g3155) & (!g3196) & (g3170) & (!g4507) & (g4508) & (!g3202)) + ((!g3155) & (!g3196) & (g3170) & (g4507) & (!g4508) & (!g3202)) + ((!g3155) & (!g3196) & (g3170) & (g4507) & (g4508) & (!g3202)) + ((!g3155) & (g3196) & (!g3170) & (!g4507) & (!g4508) & (!g3202)) + ((!g3155) & (g3196) & (!g3170) & (!g4507) & (g4508) & (!g3202)) + ((!g3155) & (g3196) & (!g3170) & (g4507) & (!g4508) & (!g3202)) + ((!g3155) & (g3196) & (!g3170) & (g4507) & (g4508) & (!g3202)) + ((!g3155) & (g3196) & (g3170) & (!g4507) & (!g4508) & (!g3202)) + ((g3155) & (!g3196) & (!g3170) & (!g4507) & (!g4508) & (!g3202)) + ((g3155) & (!g3196) & (!g3170) & (!g4507) & (!g4508) & (g3202)) + ((g3155) & (!g3196) & (!g3170) & (!g4507) & (g4508) & (!g3202)) + ((g3155) & (!g3196) & (!g3170) & (g4507) & (!g4508) & (!g3202)) + ((g3155) & (!g3196) & (!g3170) & (g4507) & (g4508) & (!g3202)) + ((g3155) & (!g3196) & (g3170) & (!g4507) & (!g4508) & (!g3202)) + ((g3155) & (!g3196) & (g3170) & (!g4507) & (g4508) & (!g3202)) + ((g3155) & (!g3196) & (g3170) & (g4507) & (!g4508) & (!g3202)) + ((g3155) & (!g3196) & (g3170) & (g4507) & (g4508) & (!g3202)) + ((g3155) & (g3196) & (!g3170) & (!g4507) & (!g4508) & (!g3202)));
	assign g4617 = (((!g1888) & (!g1978) & (!g1980) & (!g828) & (!g864) & (g897)) + ((!g1888) & (!g1978) & (!g1980) & (!g828) & (g864) & (g897)) + ((!g1888) & (!g1978) & (!g1980) & (g828) & (!g864) & (g897)) + ((!g1888) & (!g1978) & (!g1980) & (g828) & (g864) & (g897)) + ((!g1888) & (!g1978) & (g1980) & (!g828) & (!g864) & (!g897)) + ((!g1888) & (!g1978) & (g1980) & (!g828) & (g864) & (!g897)) + ((!g1888) & (!g1978) & (g1980) & (g828) & (!g864) & (!g897)) + ((!g1888) & (!g1978) & (g1980) & (g828) & (g864) & (!g897)) + ((!g1888) & (g1978) & (!g1980) & (!g828) & (!g864) & (g897)) + ((!g1888) & (g1978) & (!g1980) & (!g828) & (g864) & (!g897)) + ((!g1888) & (g1978) & (!g1980) & (g828) & (!g864) & (g897)) + ((!g1888) & (g1978) & (!g1980) & (g828) & (g864) & (!g897)) + ((!g1888) & (g1978) & (g1980) & (!g828) & (!g864) & (!g897)) + ((!g1888) & (g1978) & (g1980) & (!g828) & (g864) & (g897)) + ((!g1888) & (g1978) & (g1980) & (g828) & (!g864) & (!g897)) + ((!g1888) & (g1978) & (g1980) & (g828) & (g864) & (g897)) + ((g1888) & (!g1978) & (!g1980) & (!g828) & (!g864) & (g897)) + ((g1888) & (!g1978) & (!g1980) & (!g828) & (g864) & (g897)) + ((g1888) & (!g1978) & (!g1980) & (g828) & (!g864) & (g897)) + ((g1888) & (!g1978) & (!g1980) & (g828) & (g864) & (!g897)) + ((g1888) & (!g1978) & (g1980) & (!g828) & (!g864) & (!g897)) + ((g1888) & (!g1978) & (g1980) & (!g828) & (g864) & (!g897)) + ((g1888) & (!g1978) & (g1980) & (g828) & (!g864) & (!g897)) + ((g1888) & (!g1978) & (g1980) & (g828) & (g864) & (g897)) + ((g1888) & (g1978) & (!g1980) & (!g828) & (!g864) & (g897)) + ((g1888) & (g1978) & (!g1980) & (!g828) & (g864) & (!g897)) + ((g1888) & (g1978) & (!g1980) & (g828) & (!g864) & (!g897)) + ((g1888) & (g1978) & (!g1980) & (g828) & (g864) & (!g897)) + ((g1888) & (g1978) & (g1980) & (!g828) & (!g864) & (!g897)) + ((g1888) & (g1978) & (g1980) & (!g828) & (g864) & (g897)) + ((g1888) & (g1978) & (g1980) & (g828) & (!g864) & (g897)) + ((g1888) & (g1978) & (g1980) & (g828) & (g864) & (g897)));
	assign g4618 = (((!g1914) & (!g3240) & (!g3279) & (!g4616) & (g4617)) + ((!g1914) & (!g3240) & (!g3279) & (g4616) & (g4617)) + ((!g1914) & (!g3240) & (g3279) & (!g4616) & (g4617)) + ((!g1914) & (!g3240) & (g3279) & (g4616) & (g4617)) + ((!g1914) & (g3240) & (!g3279) & (!g4616) & (g4617)) + ((!g1914) & (g3240) & (!g3279) & (g4616) & (g4617)) + ((!g1914) & (g3240) & (g3279) & (!g4616) & (g4617)) + ((!g1914) & (g3240) & (g3279) & (g4616) & (g4617)) + ((g1914) & (!g3240) & (!g3279) & (!g4616) & (!g4617)) + ((g1914) & (!g3240) & (!g3279) & (!g4616) & (g4617)) + ((g1914) & (!g3240) & (g3279) & (g4616) & (!g4617)) + ((g1914) & (!g3240) & (g3279) & (g4616) & (g4617)) + ((g1914) & (g3240) & (!g3279) & (g4616) & (!g4617)) + ((g1914) & (g3240) & (!g3279) & (g4616) & (g4617)) + ((g1914) & (g3240) & (g3279) & (!g4616) & (!g4617)) + ((g1914) & (g3240) & (g3279) & (!g4616) & (g4617)));
	assign g4619 = (((!g830) & (!g2360) & (!g4618) & (key[105])) + ((!g830) & (!g2360) & (g4618) & (key[105])) + ((!g830) & (g2360) & (!g4618) & (key[105])) + ((!g830) & (g2360) & (g4618) & (key[105])) + ((g830) & (!g2360) & (g4618) & (!key[105])) + ((g830) & (!g2360) & (g4618) & (key[105])) + ((g830) & (g2360) & (!g4618) & (!key[105])) + ((g830) & (g2360) & (!g4618) & (key[105])));
	assign g4620 = (((!g1886) & (!g2032) & (!g2055) & (!g1902) & (!g2036) & (g2077)) + ((!g1886) & (!g2032) & (!g2055) & (!g1902) & (g2036) & (g2077)) + ((!g1886) & (!g2032) & (!g2055) & (g1902) & (!g2036) & (g2077)) + ((!g1886) & (!g2032) & (!g2055) & (g1902) & (g2036) & (g2077)) + ((!g1886) & (!g2032) & (g2055) & (!g1902) & (!g2036) & (!g2077)) + ((!g1886) & (!g2032) & (g2055) & (!g1902) & (g2036) & (!g2077)) + ((!g1886) & (!g2032) & (g2055) & (g1902) & (!g2036) & (!g2077)) + ((!g1886) & (!g2032) & (g2055) & (g1902) & (g2036) & (!g2077)) + ((!g1886) & (g2032) & (!g2055) & (!g1902) & (!g2036) & (g2077)) + ((!g1886) & (g2032) & (!g2055) & (!g1902) & (g2036) & (!g2077)) + ((!g1886) & (g2032) & (!g2055) & (g1902) & (!g2036) & (g2077)) + ((!g1886) & (g2032) & (!g2055) & (g1902) & (g2036) & (!g2077)) + ((!g1886) & (g2032) & (g2055) & (!g1902) & (!g2036) & (!g2077)) + ((!g1886) & (g2032) & (g2055) & (!g1902) & (g2036) & (g2077)) + ((!g1886) & (g2032) & (g2055) & (g1902) & (!g2036) & (!g2077)) + ((!g1886) & (g2032) & (g2055) & (g1902) & (g2036) & (g2077)) + ((g1886) & (!g2032) & (!g2055) & (!g1902) & (!g2036) & (g2077)) + ((g1886) & (!g2032) & (!g2055) & (!g1902) & (g2036) & (g2077)) + ((g1886) & (!g2032) & (!g2055) & (g1902) & (!g2036) & (g2077)) + ((g1886) & (!g2032) & (!g2055) & (g1902) & (g2036) & (!g2077)) + ((g1886) & (!g2032) & (g2055) & (!g1902) & (!g2036) & (!g2077)) + ((g1886) & (!g2032) & (g2055) & (!g1902) & (g2036) & (!g2077)) + ((g1886) & (!g2032) & (g2055) & (g1902) & (!g2036) & (!g2077)) + ((g1886) & (!g2032) & (g2055) & (g1902) & (g2036) & (g2077)) + ((g1886) & (g2032) & (!g2055) & (!g1902) & (!g2036) & (g2077)) + ((g1886) & (g2032) & (!g2055) & (!g1902) & (g2036) & (!g2077)) + ((g1886) & (g2032) & (!g2055) & (g1902) & (!g2036) & (!g2077)) + ((g1886) & (g2032) & (!g2055) & (g1902) & (g2036) & (!g2077)) + ((g1886) & (g2032) & (g2055) & (!g1902) & (!g2036) & (!g2077)) + ((g1886) & (g2032) & (g2055) & (!g1902) & (g2036) & (g2077)) + ((g1886) & (g2032) & (g2055) & (g1902) & (!g2036) & (g2077)) + ((g1886) & (g2032) & (g2055) & (g1902) & (g2036) & (g2077)));
	assign g4621 = (((!g2551) & (!g2598) & (!g3157) & (!g3207) & (!g4511) & (!g4512)) + ((!g2551) & (!g2598) & (!g3157) & (!g3207) & (!g4511) & (g4512)) + ((!g2551) & (!g2598) & (!g3157) & (!g3207) & (g4511) & (!g4512)) + ((!g2551) & (!g2598) & (!g3157) & (!g3207) & (g4511) & (g4512)) + ((!g2551) & (!g2598) & (!g3157) & (g3207) & (!g4511) & (!g4512)) + ((!g2551) & (!g2598) & (!g3157) & (g3207) & (!g4511) & (g4512)) + ((!g2551) & (!g2598) & (!g3157) & (g3207) & (g4511) & (!g4512)) + ((!g2551) & (!g2598) & (!g3157) & (g3207) & (g4511) & (g4512)) + ((!g2551) & (!g2598) & (g3157) & (!g3207) & (!g4511) & (!g4512)) + ((!g2551) & (!g2598) & (g3157) & (!g3207) & (!g4511) & (g4512)) + ((!g2551) & (!g2598) & (g3157) & (!g3207) & (g4511) & (!g4512)) + ((!g2551) & (!g2598) & (g3157) & (!g3207) & (g4511) & (g4512)) + ((!g2551) & (!g2598) & (g3157) & (g3207) & (!g4511) & (!g4512)) + ((!g2551) & (g2598) & (!g3157) & (!g3207) & (!g4511) & (!g4512)) + ((!g2551) & (g2598) & (!g3157) & (!g3207) & (!g4511) & (g4512)) + ((!g2551) & (g2598) & (!g3157) & (!g3207) & (g4511) & (!g4512)) + ((!g2551) & (g2598) & (!g3157) & (!g3207) & (g4511) & (g4512)) + ((!g2551) & (g2598) & (g3157) & (!g3207) & (!g4511) & (!g4512)) + ((g2551) & (!g2598) & (!g3157) & (!g3207) & (!g4511) & (!g4512)) + ((g2551) & (!g2598) & (!g3157) & (!g3207) & (!g4511) & (g4512)) + ((g2551) & (!g2598) & (!g3157) & (!g3207) & (g4511) & (!g4512)) + ((g2551) & (!g2598) & (!g3157) & (!g3207) & (g4511) & (g4512)) + ((g2551) & (!g2598) & (!g3157) & (g3207) & (!g4511) & (!g4512)) + ((g2551) & (!g2598) & (g3157) & (!g3207) & (!g4511) & (!g4512)) + ((g2551) & (!g2598) & (g3157) & (!g3207) & (!g4511) & (g4512)) + ((g2551) & (!g2598) & (g3157) & (!g3207) & (g4511) & (!g4512)) + ((g2551) & (!g2598) & (g3157) & (!g3207) & (g4511) & (g4512)) + ((g2551) & (g2598) & (!g3157) & (!g3207) & (!g4511) & (!g4512)));
	assign g4622 = (((!g1914) & (!g2647) & (!g3245) & (!g4620) & (!g4621)) + ((!g1914) & (!g2647) & (!g3245) & (g4620) & (!g4621)) + ((!g1914) & (!g2647) & (g3245) & (!g4620) & (g4621)) + ((!g1914) & (!g2647) & (g3245) & (g4620) & (g4621)) + ((!g1914) & (g2647) & (!g3245) & (!g4620) & (g4621)) + ((!g1914) & (g2647) & (!g3245) & (g4620) & (g4621)) + ((!g1914) & (g2647) & (g3245) & (!g4620) & (!g4621)) + ((!g1914) & (g2647) & (g3245) & (g4620) & (!g4621)) + ((g1914) & (!g2647) & (!g3245) & (g4620) & (!g4621)) + ((g1914) & (!g2647) & (!g3245) & (g4620) & (g4621)) + ((g1914) & (!g2647) & (g3245) & (g4620) & (!g4621)) + ((g1914) & (!g2647) & (g3245) & (g4620) & (g4621)) + ((g1914) & (g2647) & (!g3245) & (g4620) & (!g4621)) + ((g1914) & (g2647) & (!g3245) & (g4620) & (g4621)) + ((g1914) & (g2647) & (g3245) & (g4620) & (!g4621)) + ((g1914) & (g2647) & (g3245) & (g4620) & (g4621)));
	assign g4623 = (((!g830) & (!g2362) & (!g4622) & (nonce[9])) + ((!g830) & (!g2362) & (g4622) & (nonce[9])) + ((!g830) & (g2362) & (!g4622) & (nonce[9])) + ((!g830) & (g2362) & (g4622) & (nonce[9])) + ((g830) & (!g2362) & (g4622) & (!nonce[9])) + ((g830) & (!g2362) & (g4622) & (nonce[9])) + ((g830) & (g2362) & (!g4622) & (!nonce[9])) + ((g830) & (g2362) & (!g4622) & (nonce[9])));
	assign g4624 = (((!g2950) & (!g2999) & (g2968) & (g3020) & (!g4515) & (g4516)) + ((!g2950) & (!g2999) & (g2968) & (g3020) & (g4515) & (!g4516)) + ((!g2950) & (!g2999) & (g2968) & (g3020) & (g4515) & (g4516)) + ((!g2950) & (g2999) & (!g2968) & (g3020) & (!g4515) & (!g4516)) + ((!g2950) & (g2999) & (!g2968) & (g3020) & (!g4515) & (g4516)) + ((!g2950) & (g2999) & (!g2968) & (g3020) & (g4515) & (!g4516)) + ((!g2950) & (g2999) & (!g2968) & (g3020) & (g4515) & (g4516)) + ((!g2950) & (g2999) & (g2968) & (!g3020) & (!g4515) & (g4516)) + ((!g2950) & (g2999) & (g2968) & (!g3020) & (g4515) & (!g4516)) + ((!g2950) & (g2999) & (g2968) & (!g3020) & (g4515) & (g4516)) + ((!g2950) & (g2999) & (g2968) & (g3020) & (!g4515) & (!g4516)) + ((!g2950) & (g2999) & (g2968) & (g3020) & (!g4515) & (g4516)) + ((!g2950) & (g2999) & (g2968) & (g3020) & (g4515) & (!g4516)) + ((!g2950) & (g2999) & (g2968) & (g3020) & (g4515) & (g4516)) + ((g2950) & (!g2999) & (!g2968) & (g3020) & (!g4515) & (g4516)) + ((g2950) & (!g2999) & (!g2968) & (g3020) & (g4515) & (!g4516)) + ((g2950) & (!g2999) & (!g2968) & (g3020) & (g4515) & (g4516)) + ((g2950) & (!g2999) & (g2968) & (g3020) & (!g4515) & (!g4516)) + ((g2950) & (!g2999) & (g2968) & (g3020) & (!g4515) & (g4516)) + ((g2950) & (!g2999) & (g2968) & (g3020) & (g4515) & (!g4516)) + ((g2950) & (!g2999) & (g2968) & (g3020) & (g4515) & (g4516)) + ((g2950) & (g2999) & (!g2968) & (!g3020) & (!g4515) & (g4516)) + ((g2950) & (g2999) & (!g2968) & (!g3020) & (g4515) & (!g4516)) + ((g2950) & (g2999) & (!g2968) & (!g3020) & (g4515) & (g4516)) + ((g2950) & (g2999) & (!g2968) & (g3020) & (!g4515) & (!g4516)) + ((g2950) & (g2999) & (!g2968) & (g3020) & (!g4515) & (g4516)) + ((g2950) & (g2999) & (!g2968) & (g3020) & (g4515) & (!g4516)) + ((g2950) & (g2999) & (!g2968) & (g3020) & (g4515) & (g4516)) + ((g2950) & (g2999) & (g2968) & (!g3020) & (!g4515) & (!g4516)) + ((g2950) & (g2999) & (g2968) & (!g3020) & (!g4515) & (g4516)) + ((g2950) & (g2999) & (g2968) & (!g3020) & (g4515) & (!g4516)) + ((g2950) & (g2999) & (g2968) & (!g3020) & (g4515) & (g4516)) + ((g2950) & (g2999) & (g2968) & (g3020) & (!g4515) & (!g4516)) + ((g2950) & (g2999) & (g2968) & (g3020) & (!g4515) & (g4516)) + ((g2950) & (g2999) & (g2968) & (g3020) & (g4515) & (!g4516)) + ((g2950) & (g2999) & (g2968) & (g3020) & (g4515) & (g4516)));
	assign g4625 = (((!g3009) & (!g3031) & (!g3015) & (g3064) & (!g4575)) + ((!g3009) & (!g3031) & (!g3015) & (g3064) & (g4575)) + ((!g3009) & (!g3031) & (g3015) & (!g3064) & (g4575)) + ((!g3009) & (!g3031) & (g3015) & (g3064) & (!g4575)) + ((!g3009) & (g3031) & (!g3015) & (!g3064) & (!g4575)) + ((!g3009) & (g3031) & (!g3015) & (!g3064) & (g4575)) + ((!g3009) & (g3031) & (g3015) & (!g3064) & (!g4575)) + ((!g3009) & (g3031) & (g3015) & (g3064) & (g4575)) + ((g3009) & (!g3031) & (!g3015) & (!g3064) & (g4575)) + ((g3009) & (!g3031) & (!g3015) & (g3064) & (!g4575)) + ((g3009) & (!g3031) & (g3015) & (!g3064) & (!g4575)) + ((g3009) & (!g3031) & (g3015) & (!g3064) & (g4575)) + ((g3009) & (g3031) & (!g3015) & (!g3064) & (!g4575)) + ((g3009) & (g3031) & (!g3015) & (g3064) & (g4575)) + ((g3009) & (g3031) & (g3015) & (g3064) & (!g4575)) + ((g3009) & (g3031) & (g3015) & (g3064) & (g4575)));
	assign g4626 = (((!g1914) & (!g1906) & (!g1894) & (g1912) & (!g1902)) + ((!g1914) & (!g1906) & (!g1894) & (g1912) & (g1902)) + ((!g1914) & (!g1906) & (g1894) & (g1912) & (!g1902)) + ((!g1914) & (!g1906) & (g1894) & (g1912) & (g1902)) + ((!g1914) & (g1906) & (!g1894) & (!g1912) & (!g1902)) + ((!g1914) & (g1906) & (!g1894) & (!g1912) & (g1902)) + ((!g1914) & (g1906) & (g1894) & (!g1912) & (!g1902)) + ((!g1914) & (g1906) & (g1894) & (!g1912) & (g1902)) + ((g1914) & (!g1906) & (!g1894) & (!g1912) & (g1902)) + ((g1914) & (!g1906) & (!g1894) & (g1912) & (g1902)) + ((g1914) & (!g1906) & (g1894) & (!g1912) & (!g1902)) + ((g1914) & (!g1906) & (g1894) & (g1912) & (!g1902)) + ((g1914) & (g1906) & (!g1894) & (!g1912) & (g1902)) + ((g1914) & (g1906) & (!g1894) & (g1912) & (g1902)) + ((g1914) & (g1906) & (g1894) & (!g1912) & (!g1902)) + ((g1914) & (g1906) & (g1894) & (g1912) & (!g1902)));
	assign g4627 = (((!g830) & (!g2366) & (!g4626) & (nonce[41])) + ((!g830) & (!g2366) & (g4626) & (nonce[41])) + ((!g830) & (g2366) & (!g4626) & (nonce[41])) + ((!g830) & (g2366) & (g4626) & (nonce[41])) + ((g830) & (!g2366) & (g4626) & (!nonce[41])) + ((g830) & (!g2366) & (g4626) & (nonce[41])) + ((g830) & (g2366) & (!g4626) & (!nonce[41])) + ((g830) & (g2366) & (!g4626) & (nonce[41])));
	assign g4628 = (((!g2556) & (!g2602) & (!g3165) & (!g4524) & (!g4525) & (!g3210)) + ((!g2556) & (!g2602) & (!g3165) & (!g4524) & (!g4525) & (g3210)) + ((!g2556) & (!g2602) & (!g3165) & (!g4524) & (g4525) & (!g3210)) + ((!g2556) & (!g2602) & (!g3165) & (!g4524) & (g4525) & (g3210)) + ((!g2556) & (!g2602) & (!g3165) & (g4524) & (!g4525) & (!g3210)) + ((!g2556) & (!g2602) & (!g3165) & (g4524) & (!g4525) & (g3210)) + ((!g2556) & (!g2602) & (!g3165) & (g4524) & (g4525) & (!g3210)) + ((!g2556) & (!g2602) & (!g3165) & (g4524) & (g4525) & (g3210)) + ((!g2556) & (!g2602) & (g3165) & (!g4524) & (!g4525) & (!g3210)) + ((!g2556) & (!g2602) & (g3165) & (!g4524) & (!g4525) & (g3210)) + ((!g2556) & (!g2602) & (g3165) & (!g4524) & (g4525) & (!g3210)) + ((!g2556) & (!g2602) & (g3165) & (g4524) & (!g4525) & (!g3210)) + ((!g2556) & (!g2602) & (g3165) & (g4524) & (g4525) & (!g3210)) + ((!g2556) & (g2602) & (!g3165) & (!g4524) & (!g4525) & (!g3210)) + ((!g2556) & (g2602) & (!g3165) & (!g4524) & (g4525) & (!g3210)) + ((!g2556) & (g2602) & (!g3165) & (g4524) & (!g4525) & (!g3210)) + ((!g2556) & (g2602) & (!g3165) & (g4524) & (g4525) & (!g3210)) + ((!g2556) & (g2602) & (g3165) & (!g4524) & (!g4525) & (!g3210)) + ((g2556) & (!g2602) & (!g3165) & (!g4524) & (!g4525) & (!g3210)) + ((g2556) & (!g2602) & (!g3165) & (!g4524) & (!g4525) & (g3210)) + ((g2556) & (!g2602) & (!g3165) & (!g4524) & (g4525) & (!g3210)) + ((g2556) & (!g2602) & (!g3165) & (g4524) & (!g4525) & (!g3210)) + ((g2556) & (!g2602) & (!g3165) & (g4524) & (g4525) & (!g3210)) + ((g2556) & (!g2602) & (g3165) & (!g4524) & (!g4525) & (!g3210)) + ((g2556) & (!g2602) & (g3165) & (!g4524) & (g4525) & (!g3210)) + ((g2556) & (!g2602) & (g3165) & (g4524) & (!g4525) & (!g3210)) + ((g2556) & (!g2602) & (g3165) & (g4524) & (g4525) & (!g3210)) + ((g2556) & (g2602) & (!g3165) & (!g4524) & (!g4525) & (!g3210)));
	assign g4629 = (((!g1892) & (!g2026) & (!g2062) & (!g1894) & (!g2034) & (g2065)) + ((!g1892) & (!g2026) & (!g2062) & (!g1894) & (g2034) & (g2065)) + ((!g1892) & (!g2026) & (!g2062) & (g1894) & (!g2034) & (g2065)) + ((!g1892) & (!g2026) & (!g2062) & (g1894) & (g2034) & (g2065)) + ((!g1892) & (!g2026) & (g2062) & (!g1894) & (!g2034) & (!g2065)) + ((!g1892) & (!g2026) & (g2062) & (!g1894) & (g2034) & (!g2065)) + ((!g1892) & (!g2026) & (g2062) & (g1894) & (!g2034) & (!g2065)) + ((!g1892) & (!g2026) & (g2062) & (g1894) & (g2034) & (!g2065)) + ((!g1892) & (g2026) & (!g2062) & (!g1894) & (!g2034) & (g2065)) + ((!g1892) & (g2026) & (!g2062) & (!g1894) & (g2034) & (!g2065)) + ((!g1892) & (g2026) & (!g2062) & (g1894) & (!g2034) & (g2065)) + ((!g1892) & (g2026) & (!g2062) & (g1894) & (g2034) & (!g2065)) + ((!g1892) & (g2026) & (g2062) & (!g1894) & (!g2034) & (!g2065)) + ((!g1892) & (g2026) & (g2062) & (!g1894) & (g2034) & (g2065)) + ((!g1892) & (g2026) & (g2062) & (g1894) & (!g2034) & (!g2065)) + ((!g1892) & (g2026) & (g2062) & (g1894) & (g2034) & (g2065)) + ((g1892) & (!g2026) & (!g2062) & (!g1894) & (!g2034) & (g2065)) + ((g1892) & (!g2026) & (!g2062) & (!g1894) & (g2034) & (g2065)) + ((g1892) & (!g2026) & (!g2062) & (g1894) & (!g2034) & (g2065)) + ((g1892) & (!g2026) & (!g2062) & (g1894) & (g2034) & (!g2065)) + ((g1892) & (!g2026) & (g2062) & (!g1894) & (!g2034) & (!g2065)) + ((g1892) & (!g2026) & (g2062) & (!g1894) & (g2034) & (!g2065)) + ((g1892) & (!g2026) & (g2062) & (g1894) & (!g2034) & (!g2065)) + ((g1892) & (!g2026) & (g2062) & (g1894) & (g2034) & (g2065)) + ((g1892) & (g2026) & (!g2062) & (!g1894) & (!g2034) & (g2065)) + ((g1892) & (g2026) & (!g2062) & (!g1894) & (g2034) & (!g2065)) + ((g1892) & (g2026) & (!g2062) & (g1894) & (!g2034) & (!g2065)) + ((g1892) & (g2026) & (!g2062) & (g1894) & (g2034) & (!g2065)) + ((g1892) & (g2026) & (g2062) & (!g1894) & (!g2034) & (!g2065)) + ((g1892) & (g2026) & (g2062) & (!g1894) & (g2034) & (g2065)) + ((g1892) & (g2026) & (g2062) & (g1894) & (!g2034) & (g2065)) + ((g1892) & (g2026) & (g2062) & (g1894) & (g2034) & (g2065)));
	assign g4630 = (((!g1914) & (!g2650) & (!g3265) & (!g4628) & (g4629)) + ((!g1914) & (!g2650) & (!g3265) & (g4628) & (g4629)) + ((!g1914) & (!g2650) & (g3265) & (!g4628) & (g4629)) + ((!g1914) & (!g2650) & (g3265) & (g4628) & (g4629)) + ((!g1914) & (g2650) & (!g3265) & (!g4628) & (g4629)) + ((!g1914) & (g2650) & (!g3265) & (g4628) & (g4629)) + ((!g1914) & (g2650) & (g3265) & (!g4628) & (g4629)) + ((!g1914) & (g2650) & (g3265) & (g4628) & (g4629)) + ((g1914) & (!g2650) & (!g3265) & (!g4628) & (!g4629)) + ((g1914) & (!g2650) & (!g3265) & (!g4628) & (g4629)) + ((g1914) & (!g2650) & (g3265) & (g4628) & (!g4629)) + ((g1914) & (!g2650) & (g3265) & (g4628) & (g4629)) + ((g1914) & (g2650) & (!g3265) & (g4628) & (!g4629)) + ((g1914) & (g2650) & (!g3265) & (g4628) & (g4629)) + ((g1914) & (g2650) & (g3265) & (!g4628) & (!g4629)) + ((g1914) & (g2650) & (g3265) & (!g4628) & (g4629)));
	assign g4631 = (((!g830) & (!g2369) & (!g4630) & (key[233])) + ((!g830) & (!g2369) & (g4630) & (key[233])) + ((!g830) & (g2369) & (!g4630) & (key[233])) + ((!g830) & (g2369) & (g4630) & (key[233])) + ((g830) & (!g2369) & (g4630) & (!key[233])) + ((g830) & (!g2369) & (g4630) & (key[233])) + ((g830) & (g2369) & (!g4630) & (!key[233])) + ((g830) & (g2369) & (!g4630) & (key[233])));
	assign g4632 = (((!g1914) & (!g1888) & (!g1912) & (!g1900) & (g1902)) + ((!g1914) & (!g1888) & (!g1912) & (g1900) & (!g1902)) + ((!g1914) & (!g1888) & (g1912) & (!g1900) & (g1902)) + ((!g1914) & (!g1888) & (g1912) & (g1900) & (!g1902)) + ((!g1914) & (g1888) & (!g1912) & (!g1900) & (g1902)) + ((!g1914) & (g1888) & (!g1912) & (g1900) & (!g1902)) + ((!g1914) & (g1888) & (g1912) & (!g1900) & (g1902)) + ((!g1914) & (g1888) & (g1912) & (g1900) & (!g1902)) + ((g1914) & (!g1888) & (g1912) & (!g1900) & (!g1902)) + ((g1914) & (!g1888) & (g1912) & (!g1900) & (g1902)) + ((g1914) & (!g1888) & (g1912) & (g1900) & (!g1902)) + ((g1914) & (!g1888) & (g1912) & (g1900) & (g1902)) + ((g1914) & (g1888) & (!g1912) & (!g1900) & (!g1902)) + ((g1914) & (g1888) & (!g1912) & (!g1900) & (g1902)) + ((g1914) & (g1888) & (!g1912) & (g1900) & (!g1902)) + ((g1914) & (g1888) & (!g1912) & (g1900) & (g1902)));
	assign g4633 = (((!g830) & (!g2371) & (!g4632) & (key[201])) + ((!g830) & (!g2371) & (g4632) & (key[201])) + ((!g830) & (g2371) & (!g4632) & (key[201])) + ((!g830) & (g2371) & (g4632) & (key[201])) + ((g830) & (!g2371) & (g4632) & (!key[201])) + ((g830) & (!g2371) & (g4632) & (key[201])) + ((g830) & (g2371) & (!g4632) & (!key[201])) + ((g830) & (g2371) & (!g4632) & (key[201])));
	assign g4634 = (((!g2979) & (!g3007) & (g2985) & (g3015) & (!g4531) & (g4532)) + ((!g2979) & (!g3007) & (g2985) & (g3015) & (g4531) & (!g4532)) + ((!g2979) & (!g3007) & (g2985) & (g3015) & (g4531) & (g4532)) + ((!g2979) & (g3007) & (!g2985) & (g3015) & (!g4531) & (!g4532)) + ((!g2979) & (g3007) & (!g2985) & (g3015) & (!g4531) & (g4532)) + ((!g2979) & (g3007) & (!g2985) & (g3015) & (g4531) & (!g4532)) + ((!g2979) & (g3007) & (!g2985) & (g3015) & (g4531) & (g4532)) + ((!g2979) & (g3007) & (g2985) & (!g3015) & (!g4531) & (g4532)) + ((!g2979) & (g3007) & (g2985) & (!g3015) & (g4531) & (!g4532)) + ((!g2979) & (g3007) & (g2985) & (!g3015) & (g4531) & (g4532)) + ((!g2979) & (g3007) & (g2985) & (g3015) & (!g4531) & (!g4532)) + ((!g2979) & (g3007) & (g2985) & (g3015) & (!g4531) & (g4532)) + ((!g2979) & (g3007) & (g2985) & (g3015) & (g4531) & (!g4532)) + ((!g2979) & (g3007) & (g2985) & (g3015) & (g4531) & (g4532)) + ((g2979) & (!g3007) & (!g2985) & (g3015) & (!g4531) & (g4532)) + ((g2979) & (!g3007) & (!g2985) & (g3015) & (g4531) & (!g4532)) + ((g2979) & (!g3007) & (!g2985) & (g3015) & (g4531) & (g4532)) + ((g2979) & (!g3007) & (g2985) & (g3015) & (!g4531) & (!g4532)) + ((g2979) & (!g3007) & (g2985) & (g3015) & (!g4531) & (g4532)) + ((g2979) & (!g3007) & (g2985) & (g3015) & (g4531) & (!g4532)) + ((g2979) & (!g3007) & (g2985) & (g3015) & (g4531) & (g4532)) + ((g2979) & (g3007) & (!g2985) & (!g3015) & (!g4531) & (g4532)) + ((g2979) & (g3007) & (!g2985) & (!g3015) & (g4531) & (!g4532)) + ((g2979) & (g3007) & (!g2985) & (!g3015) & (g4531) & (g4532)) + ((g2979) & (g3007) & (!g2985) & (g3015) & (!g4531) & (!g4532)) + ((g2979) & (g3007) & (!g2985) & (g3015) & (!g4531) & (g4532)) + ((g2979) & (g3007) & (!g2985) & (g3015) & (g4531) & (!g4532)) + ((g2979) & (g3007) & (!g2985) & (g3015) & (g4531) & (g4532)) + ((g2979) & (g3007) & (g2985) & (!g3015) & (!g4531) & (!g4532)) + ((g2979) & (g3007) & (g2985) & (!g3015) & (!g4531) & (g4532)) + ((g2979) & (g3007) & (g2985) & (!g3015) & (g4531) & (!g4532)) + ((g2979) & (g3007) & (g2985) & (!g3015) & (g4531) & (g4532)) + ((g2979) & (g3007) & (g2985) & (g3015) & (!g4531) & (!g4532)) + ((g2979) & (g3007) & (g2985) & (g3015) & (!g4531) & (g4532)) + ((g2979) & (g3007) & (g2985) & (g3015) & (g4531) & (!g4532)) + ((g2979) & (g3007) & (g2985) & (g3015) & (g4531) & (g4532)));
	assign g4635 = (((!g3018) & (!g3044) & (!g3020) & (g3056) & (!g4587)) + ((!g3018) & (!g3044) & (!g3020) & (g3056) & (g4587)) + ((!g3018) & (!g3044) & (g3020) & (!g3056) & (g4587)) + ((!g3018) & (!g3044) & (g3020) & (g3056) & (!g4587)) + ((!g3018) & (g3044) & (!g3020) & (!g3056) & (!g4587)) + ((!g3018) & (g3044) & (!g3020) & (!g3056) & (g4587)) + ((!g3018) & (g3044) & (g3020) & (!g3056) & (!g4587)) + ((!g3018) & (g3044) & (g3020) & (g3056) & (g4587)) + ((g3018) & (!g3044) & (!g3020) & (!g3056) & (g4587)) + ((g3018) & (!g3044) & (!g3020) & (g3056) & (!g4587)) + ((g3018) & (!g3044) & (g3020) & (!g3056) & (!g4587)) + ((g3018) & (!g3044) & (g3020) & (!g3056) & (g4587)) + ((g3018) & (g3044) & (!g3020) & (!g3056) & (!g4587)) + ((g3018) & (g3044) & (!g3020) & (g3056) & (g4587)) + ((g3018) & (g3044) & (g3020) & (g3056) & (!g4587)) + ((g3018) & (g3044) & (g3020) & (g3056) & (g4587)));
	assign g4636 = (((!g1269) & (!g3507) & (g2559)) + ((g1269) & (!g3507) & (!g2559)) + ((g1269) & (!g3507) & (g2559)) + ((g1269) & (g3507) & (g2559)));
	assign g4637 = (((g1914) & (!g1303) & (!g4636) & (g2623)) + ((g1914) & (!g1303) & (g4636) & (!g2623)) + ((g1914) & (g1303) & (!g4636) & (!g2623)) + ((g1914) & (g1303) & (g4636) & (g2623)));
	assign g4638 = (((!g2566) & (g2589) & (!g3525)) + ((g2566) & (!g2589) & (!g3525)) + ((g2566) & (g2589) & (!g3525)) + ((g2566) & (g2589) & (g3525)));
	assign g4639 = (((!g1914) & (!g2614) & (!g2620) & (g4638)) + ((!g1914) & (!g2614) & (g2620) & (!g4638)) + ((!g1914) & (g2614) & (!g2620) & (!g4638)) + ((!g1914) & (g2614) & (g2620) & (g4638)));
	assign g4640 = (((!g830) & (!g2376) & (!g4637) & (!g4639) & (key[55])) + ((!g830) & (!g2376) & (!g4637) & (g4639) & (key[55])) + ((!g830) & (!g2376) & (g4637) & (!g4639) & (key[55])) + ((!g830) & (!g2376) & (g4637) & (g4639) & (key[55])) + ((!g830) & (g2376) & (!g4637) & (!g4639) & (key[55])) + ((!g830) & (g2376) & (!g4637) & (g4639) & (key[55])) + ((!g830) & (g2376) & (g4637) & (!g4639) & (key[55])) + ((!g830) & (g2376) & (g4637) & (g4639) & (key[55])) + ((g830) & (!g2376) & (!g4637) & (g4639) & (!key[55])) + ((g830) & (!g2376) & (!g4637) & (g4639) & (key[55])) + ((g830) & (!g2376) & (g4637) & (!g4639) & (!key[55])) + ((g830) & (!g2376) & (g4637) & (!g4639) & (key[55])) + ((g830) & (!g2376) & (g4637) & (g4639) & (!key[55])) + ((g830) & (!g2376) & (g4637) & (g4639) & (key[55])) + ((g830) & (g2376) & (!g4637) & (!g4639) & (!key[55])) + ((g830) & (g2376) & (!g4637) & (!g4639) & (key[55])));
	assign g4641 = (((!g3768) & (g3769)) + ((g3768) & (!g3769)) + ((g3768) & (g3769)));
	assign g4642 = (((!g1960) & (!g1962) & (!g2350) & (g2399) & (!g4591)) + ((!g1960) & (!g1962) & (!g2350) & (g2399) & (g4591)) + ((!g1960) & (!g1962) & (g2350) & (!g2399) & (g4591)) + ((!g1960) & (!g1962) & (g2350) & (g2399) & (!g4591)) + ((!g1960) & (g1962) & (!g2350) & (!g2399) & (!g4591)) + ((!g1960) & (g1962) & (!g2350) & (!g2399) & (g4591)) + ((!g1960) & (g1962) & (g2350) & (!g2399) & (!g4591)) + ((!g1960) & (g1962) & (g2350) & (g2399) & (g4591)) + ((g1960) & (!g1962) & (!g2350) & (!g2399) & (g4591)) + ((g1960) & (!g1962) & (!g2350) & (g2399) & (!g4591)) + ((g1960) & (!g1962) & (g2350) & (!g2399) & (!g4591)) + ((g1960) & (!g1962) & (g2350) & (!g2399) & (g4591)) + ((g1960) & (g1962) & (!g2350) & (!g2399) & (!g4591)) + ((g1960) & (g1962) & (!g2350) & (g2399) & (g4591)) + ((g1960) & (g1962) & (g2350) & (g2399) & (!g4591)) + ((g1960) & (g1962) & (g2350) & (g2399) & (g4591)));
	assign g4643 = (((!g1914) & (!g2742) & (!g2752) & (g4641) & (!g4642)) + ((!g1914) & (!g2742) & (!g2752) & (g4641) & (g4642)) + ((!g1914) & (!g2742) & (g2752) & (!g4641) & (!g4642)) + ((!g1914) & (!g2742) & (g2752) & (!g4641) & (g4642)) + ((!g1914) & (g2742) & (!g2752) & (!g4641) & (!g4642)) + ((!g1914) & (g2742) & (!g2752) & (!g4641) & (g4642)) + ((!g1914) & (g2742) & (g2752) & (g4641) & (!g4642)) + ((!g1914) & (g2742) & (g2752) & (g4641) & (g4642)) + ((g1914) & (!g2742) & (!g2752) & (!g4641) & (g4642)) + ((g1914) & (!g2742) & (!g2752) & (g4641) & (g4642)) + ((g1914) & (!g2742) & (g2752) & (!g4641) & (g4642)) + ((g1914) & (!g2742) & (g2752) & (g4641) & (g4642)) + ((g1914) & (g2742) & (!g2752) & (!g4641) & (g4642)) + ((g1914) & (g2742) & (!g2752) & (g4641) & (g4642)) + ((g1914) & (g2742) & (g2752) & (!g4641) & (g4642)) + ((g1914) & (g2742) & (g2752) & (g4641) & (g4642)));
	assign g4644 = (((!g830) & (!g2377) & (!g4643) & (key[87])) + ((!g830) & (!g2377) & (g4643) & (key[87])) + ((!g830) & (g2377) & (!g4643) & (key[87])) + ((!g830) & (g2377) & (g4643) & (key[87])) + ((g830) & (!g2377) & (g4643) & (!key[87])) + ((g830) & (!g2377) & (g4643) & (key[87])) + ((g830) & (g2377) & (!g4643) & (!key[87])) + ((g830) & (g2377) & (!g4643) & (key[87])));
	assign g4645 = (((!g1269) & (!g3417) & (g2575)) + ((g1269) & (!g3417) & (!g2575)) + ((g1269) & (!g3417) & (g2575)) + ((g1269) & (g3417) & (g2575)));
	assign g4646 = (((!g3400) & (!g2566) & (g2572)) + ((!g3400) & (g2566) & (!g2572)) + ((!g3400) & (g2566) & (g2572)) + ((g3400) & (g2566) & (g2572)));
	assign g4647 = (((!g4646) & (!g2614) & (g2637)) + ((!g4646) & (g2614) & (!g2637)) + ((g4646) & (!g2614) & (!g2637)) + ((g4646) & (g2614) & (g2637)));
	assign g4648 = (((!g1914) & (!g1303) & (!g4645) & (g2607) & (!g4647)) + ((!g1914) & (!g1303) & (!g4645) & (g2607) & (g4647)) + ((!g1914) & (!g1303) & (g4645) & (!g2607) & (!g4647)) + ((!g1914) & (!g1303) & (g4645) & (!g2607) & (g4647)) + ((!g1914) & (g1303) & (!g4645) & (!g2607) & (!g4647)) + ((!g1914) & (g1303) & (!g4645) & (!g2607) & (g4647)) + ((!g1914) & (g1303) & (g4645) & (g2607) & (!g4647)) + ((!g1914) & (g1303) & (g4645) & (g2607) & (g4647)) + ((g1914) & (!g1303) & (!g4645) & (!g2607) & (g4647)) + ((g1914) & (!g1303) & (!g4645) & (g2607) & (g4647)) + ((g1914) & (!g1303) & (g4645) & (!g2607) & (g4647)) + ((g1914) & (!g1303) & (g4645) & (g2607) & (g4647)) + ((g1914) & (g1303) & (!g4645) & (!g2607) & (g4647)) + ((g1914) & (g1303) & (!g4645) & (g2607) & (g4647)) + ((g1914) & (g1303) & (g4645) & (!g2607) & (g4647)) + ((g1914) & (g1303) & (g4645) & (g2607) & (g4647)));
	assign g8309 = (((!g5560) & (g5607) & (!g4649)) + ((!g5560) & (g5607) & (g4649)) + ((g5560) & (!g5607) & (g4649)) + ((g5560) & (g5607) & (g4649)));
	assign g4650 = (((!g830) & (!g2378) & (!g4648) & (g4649)) + ((!g830) & (!g2378) & (g4648) & (g4649)) + ((!g830) & (g2378) & (!g4648) & (g4649)) + ((!g830) & (g2378) & (g4648) & (g4649)) + ((g830) & (!g2378) & (g4648) & (!g4649)) + ((g830) & (!g2378) & (g4648) & (g4649)) + ((g830) & (g2378) & (!g4648) & (!g4649)) + ((g830) & (g2378) & (!g4648) & (g4649)));
	assign g4651 = (((!g3475) & (g3476)) + ((g3475) & (!g3476)) + ((g3475) & (g3476)));
	assign g4652 = (((!g1998) & (!g2001) & (!g2360) & (g2383) & (!g4598)) + ((!g1998) & (!g2001) & (!g2360) & (g2383) & (g4598)) + ((!g1998) & (!g2001) & (g2360) & (!g2383) & (g4598)) + ((!g1998) & (!g2001) & (g2360) & (g2383) & (!g4598)) + ((!g1998) & (g2001) & (!g2360) & (!g2383) & (!g4598)) + ((!g1998) & (g2001) & (!g2360) & (!g2383) & (g4598)) + ((!g1998) & (g2001) & (g2360) & (!g2383) & (!g4598)) + ((!g1998) & (g2001) & (g2360) & (g2383) & (g4598)) + ((g1998) & (!g2001) & (!g2360) & (!g2383) & (g4598)) + ((g1998) & (!g2001) & (!g2360) & (g2383) & (!g4598)) + ((g1998) & (!g2001) & (g2360) & (!g2383) & (!g4598)) + ((g1998) & (!g2001) & (g2360) & (!g2383) & (g4598)) + ((g1998) & (g2001) & (!g2360) & (!g2383) & (!g4598)) + ((g1998) & (g2001) & (!g2360) & (g2383) & (g4598)) + ((g1998) & (g2001) & (g2360) & (g2383) & (!g4598)) + ((g1998) & (g2001) & (g2360) & (g2383) & (g4598)));
	assign g4653 = (((!g1914) & (!g4651) & (!g2713) & (!g2752) & (g4652)) + ((!g1914) & (!g4651) & (!g2713) & (g2752) & (g4652)) + ((!g1914) & (!g4651) & (g2713) & (!g2752) & (g4652)) + ((!g1914) & (!g4651) & (g2713) & (g2752) & (g4652)) + ((!g1914) & (g4651) & (!g2713) & (!g2752) & (g4652)) + ((!g1914) & (g4651) & (!g2713) & (g2752) & (g4652)) + ((!g1914) & (g4651) & (g2713) & (!g2752) & (g4652)) + ((!g1914) & (g4651) & (g2713) & (g2752) & (g4652)) + ((g1914) & (!g4651) & (!g2713) & (g2752) & (!g4652)) + ((g1914) & (!g4651) & (!g2713) & (g2752) & (g4652)) + ((g1914) & (!g4651) & (g2713) & (!g2752) & (!g4652)) + ((g1914) & (!g4651) & (g2713) & (!g2752) & (g4652)) + ((g1914) & (g4651) & (!g2713) & (!g2752) & (!g4652)) + ((g1914) & (g4651) & (!g2713) & (!g2752) & (g4652)) + ((g1914) & (g4651) & (g2713) & (g2752) & (!g4652)) + ((g1914) & (g4651) & (g2713) & (g2752) & (g4652)));
	assign g4654 = (((!g830) & (!g2379) & (!g4653) & (key[183])) + ((!g830) & (!g2379) & (g4653) & (key[183])) + ((!g830) & (g2379) & (!g4653) & (key[183])) + ((!g830) & (g2379) & (g4653) & (key[183])) + ((g830) & (!g2379) & (g4653) & (!key[183])) + ((g830) & (!g2379) & (g4653) & (key[183])) + ((g830) & (g2379) & (!g4653) & (!key[183])) + ((g830) & (g2379) & (!g4653) & (key[183])));
	assign g4655 = (((!g3240) & (!g3303) & (!g3279) & (!g4616) & (g3307)) + ((!g3240) & (!g3303) & (!g3279) & (g4616) & (g3307)) + ((!g3240) & (!g3303) & (g3279) & (!g4616) & (!g3307)) + ((!g3240) & (!g3303) & (g3279) & (g4616) & (g3307)) + ((!g3240) & (g3303) & (!g3279) & (!g4616) & (!g3307)) + ((!g3240) & (g3303) & (!g3279) & (g4616) & (!g3307)) + ((!g3240) & (g3303) & (g3279) & (!g4616) & (g3307)) + ((!g3240) & (g3303) & (g3279) & (g4616) & (!g3307)) + ((g3240) & (!g3303) & (!g3279) & (!g4616) & (!g3307)) + ((g3240) & (!g3303) & (!g3279) & (g4616) & (g3307)) + ((g3240) & (!g3303) & (g3279) & (!g4616) & (!g3307)) + ((g3240) & (!g3303) & (g3279) & (g4616) & (!g3307)) + ((g3240) & (g3303) & (!g3279) & (!g4616) & (g3307)) + ((g3240) & (g3303) & (!g3279) & (g4616) & (!g3307)) + ((g3240) & (g3303) & (g3279) & (!g4616) & (g3307)) + ((g3240) & (g3303) & (g3279) & (g4616) & (g3307)));
	assign g4656 = (((!g1983) & (!g931) & (g3444)) + ((!g1983) & (g931) & (!g3444)) + ((g1983) & (!g931) & (!g3444)) + ((g1983) & (g931) & (g3444)));
	assign g4657 = (((!g830) & (!g1914) & (!g2383) & (!g4655) & (!g4656) & (key[106])) + ((!g830) & (!g1914) & (!g2383) & (!g4655) & (g4656) & (key[106])) + ((!g830) & (!g1914) & (!g2383) & (g4655) & (!g4656) & (key[106])) + ((!g830) & (!g1914) & (!g2383) & (g4655) & (g4656) & (key[106])) + ((!g830) & (!g1914) & (g2383) & (!g4655) & (!g4656) & (key[106])) + ((!g830) & (!g1914) & (g2383) & (!g4655) & (g4656) & (key[106])) + ((!g830) & (!g1914) & (g2383) & (g4655) & (!g4656) & (key[106])) + ((!g830) & (!g1914) & (g2383) & (g4655) & (g4656) & (key[106])) + ((!g830) & (g1914) & (!g2383) & (!g4655) & (!g4656) & (key[106])) + ((!g830) & (g1914) & (!g2383) & (!g4655) & (g4656) & (key[106])) + ((!g830) & (g1914) & (!g2383) & (g4655) & (!g4656) & (key[106])) + ((!g830) & (g1914) & (!g2383) & (g4655) & (g4656) & (key[106])) + ((!g830) & (g1914) & (g2383) & (!g4655) & (!g4656) & (key[106])) + ((!g830) & (g1914) & (g2383) & (!g4655) & (g4656) & (key[106])) + ((!g830) & (g1914) & (g2383) & (g4655) & (!g4656) & (key[106])) + ((!g830) & (g1914) & (g2383) & (g4655) & (g4656) & (key[106])) + ((g830) & (!g1914) & (!g2383) & (!g4655) & (g4656) & (!key[106])) + ((g830) & (!g1914) & (!g2383) & (!g4655) & (g4656) & (key[106])) + ((g830) & (!g1914) & (!g2383) & (g4655) & (g4656) & (!key[106])) + ((g830) & (!g1914) & (!g2383) & (g4655) & (g4656) & (key[106])) + ((g830) & (!g1914) & (g2383) & (!g4655) & (!g4656) & (!key[106])) + ((g830) & (!g1914) & (g2383) & (!g4655) & (!g4656) & (key[106])) + ((g830) & (!g1914) & (g2383) & (g4655) & (!g4656) & (!key[106])) + ((g830) & (!g1914) & (g2383) & (g4655) & (!g4656) & (key[106])) + ((g830) & (g1914) & (!g2383) & (g4655) & (!g4656) & (!key[106])) + ((g830) & (g1914) & (!g2383) & (g4655) & (!g4656) & (key[106])) + ((g830) & (g1914) & (!g2383) & (g4655) & (g4656) & (!key[106])) + ((g830) & (g1914) & (!g2383) & (g4655) & (g4656) & (key[106])) + ((g830) & (g1914) & (g2383) & (!g4655) & (!g4656) & (!key[106])) + ((g830) & (g1914) & (g2383) & (!g4655) & (!g4656) & (key[106])) + ((g830) & (g1914) & (g2383) & (!g4655) & (g4656) & (!key[106])) + ((g830) & (g1914) & (g2383) & (!g4655) & (g4656) & (key[106])));
	assign g4658 = (((!g2378) & (g3041) & (g4605)) + ((g2378) & (!g3041) & (g4605)) + ((g2378) & (g3041) & (!g4605)) + ((g2378) & (g3041) & (g4605)));
	assign g4659 = (((!g2343) & (!g2376) & (g3005) & (g3050) & (g4556)) + ((!g2343) & (g2376) & (!g3005) & (g3050) & (!g4556)) + ((!g2343) & (g2376) & (!g3005) & (g3050) & (g4556)) + ((!g2343) & (g2376) & (g3005) & (!g3050) & (g4556)) + ((!g2343) & (g2376) & (g3005) & (g3050) & (!g4556)) + ((!g2343) & (g2376) & (g3005) & (g3050) & (g4556)) + ((g2343) & (!g2376) & (!g3005) & (g3050) & (g4556)) + ((g2343) & (!g2376) & (g3005) & (g3050) & (!g4556)) + ((g2343) & (!g2376) & (g3005) & (g3050) & (g4556)) + ((g2343) & (g2376) & (!g3005) & (!g3050) & (g4556)) + ((g2343) & (g2376) & (!g3005) & (g3050) & (!g4556)) + ((g2343) & (g2376) & (!g3005) & (g3050) & (g4556)) + ((g2343) & (g2376) & (g3005) & (!g3050) & (!g4556)) + ((g2343) & (g2376) & (g3005) & (!g3050) & (g4556)) + ((g2343) & (g2376) & (g3005) & (g3050) & (!g4556)) + ((g2343) & (g2376) & (g3005) & (g3050) & (g4556)));
	assign g4660 = (((!g2423) & (!g3080) & (g4659)) + ((!g2423) & (g3080) & (!g4659)) + ((g2423) & (!g3080) & (!g4659)) + ((g2423) & (g3080) & (g4659)));
	assign g4661 = (((!g2114) & (!g3555) & (g2118)) + ((!g2114) & (g3555) & (!g2118)) + ((g2114) & (!g3555) & (!g2118)) + ((g2114) & (g3555) & (g2118)));
	assign g4662 = (((!g2647) & (!g2678) & (!g3245) & (g3310) & (!g4621)) + ((!g2647) & (!g2678) & (!g3245) & (g3310) & (g4621)) + ((!g2647) & (!g2678) & (g3245) & (!g3310) & (!g4621)) + ((!g2647) & (!g2678) & (g3245) & (g3310) & (g4621)) + ((!g2647) & (g2678) & (!g3245) & (!g3310) & (!g4621)) + ((!g2647) & (g2678) & (!g3245) & (!g3310) & (g4621)) + ((!g2647) & (g2678) & (g3245) & (!g3310) & (g4621)) + ((!g2647) & (g2678) & (g3245) & (g3310) & (!g4621)) + ((g2647) & (!g2678) & (!g3245) & (!g3310) & (!g4621)) + ((g2647) & (!g2678) & (!g3245) & (g3310) & (g4621)) + ((g2647) & (!g2678) & (g3245) & (!g3310) & (!g4621)) + ((g2647) & (!g2678) & (g3245) & (!g3310) & (g4621)) + ((g2647) & (g2678) & (!g3245) & (!g3310) & (g4621)) + ((g2647) & (g2678) & (!g3245) & (g3310) & (!g4621)) + ((g2647) & (g2678) & (g3245) & (g3310) & (!g4621)) + ((g2647) & (g2678) & (g3245) & (g3310) & (g4621)));
	assign g4663 = (((!g830) & (!g1914) & (!g2393) & (!g4661) & (!g4662) & (nonce[10])) + ((!g830) & (!g1914) & (!g2393) & (!g4661) & (g4662) & (nonce[10])) + ((!g830) & (!g1914) & (!g2393) & (g4661) & (!g4662) & (nonce[10])) + ((!g830) & (!g1914) & (!g2393) & (g4661) & (g4662) & (nonce[10])) + ((!g830) & (!g1914) & (g2393) & (!g4661) & (!g4662) & (nonce[10])) + ((!g830) & (!g1914) & (g2393) & (!g4661) & (g4662) & (nonce[10])) + ((!g830) & (!g1914) & (g2393) & (g4661) & (!g4662) & (nonce[10])) + ((!g830) & (!g1914) & (g2393) & (g4661) & (g4662) & (nonce[10])) + ((!g830) & (g1914) & (!g2393) & (!g4661) & (!g4662) & (nonce[10])) + ((!g830) & (g1914) & (!g2393) & (!g4661) & (g4662) & (nonce[10])) + ((!g830) & (g1914) & (!g2393) & (g4661) & (!g4662) & (nonce[10])) + ((!g830) & (g1914) & (!g2393) & (g4661) & (g4662) & (nonce[10])) + ((!g830) & (g1914) & (g2393) & (!g4661) & (!g4662) & (nonce[10])) + ((!g830) & (g1914) & (g2393) & (!g4661) & (g4662) & (nonce[10])) + ((!g830) & (g1914) & (g2393) & (g4661) & (!g4662) & (nonce[10])) + ((!g830) & (g1914) & (g2393) & (g4661) & (g4662) & (nonce[10])) + ((g830) & (!g1914) & (!g2393) & (!g4661) & (g4662) & (!nonce[10])) + ((g830) & (!g1914) & (!g2393) & (!g4661) & (g4662) & (nonce[10])) + ((g830) & (!g1914) & (!g2393) & (g4661) & (g4662) & (!nonce[10])) + ((g830) & (!g1914) & (!g2393) & (g4661) & (g4662) & (nonce[10])) + ((g830) & (!g1914) & (g2393) & (!g4661) & (!g4662) & (!nonce[10])) + ((g830) & (!g1914) & (g2393) & (!g4661) & (!g4662) & (nonce[10])) + ((g830) & (!g1914) & (g2393) & (g4661) & (!g4662) & (!nonce[10])) + ((g830) & (!g1914) & (g2393) & (g4661) & (!g4662) & (nonce[10])) + ((g830) & (g1914) & (!g2393) & (g4661) & (!g4662) & (!nonce[10])) + ((g830) & (g1914) & (!g2393) & (g4661) & (!g4662) & (nonce[10])) + ((g830) & (g1914) & (!g2393) & (g4661) & (g4662) & (!nonce[10])) + ((g830) & (g1914) & (!g2393) & (g4661) & (g4662) & (nonce[10])) + ((g830) & (g1914) & (g2393) & (!g4661) & (!g4662) & (!nonce[10])) + ((g830) & (g1914) & (g2393) & (!g4661) & (!g4662) & (nonce[10])) + ((g830) & (g1914) & (g2393) & (!g4661) & (g4662) & (!nonce[10])) + ((g830) & (g1914) & (g2393) & (!g4661) & (g4662) & (nonce[10])));
	assign g4664 = (((!g2650) & (!g2684) & (!g3265) & (!g4628) & (g3312)) + ((!g2650) & (!g2684) & (!g3265) & (g4628) & (g3312)) + ((!g2650) & (!g2684) & (g3265) & (!g4628) & (!g3312)) + ((!g2650) & (!g2684) & (g3265) & (g4628) & (g3312)) + ((!g2650) & (g2684) & (!g3265) & (!g4628) & (!g3312)) + ((!g2650) & (g2684) & (!g3265) & (g4628) & (!g3312)) + ((!g2650) & (g2684) & (g3265) & (!g4628) & (g3312)) + ((!g2650) & (g2684) & (g3265) & (g4628) & (!g3312)) + ((g2650) & (!g2684) & (!g3265) & (!g4628) & (!g3312)) + ((g2650) & (!g2684) & (!g3265) & (g4628) & (g3312)) + ((g2650) & (!g2684) & (g3265) & (!g4628) & (!g3312)) + ((g2650) & (!g2684) & (g3265) & (g4628) & (!g3312)) + ((g2650) & (g2684) & (!g3265) & (!g4628) & (g3312)) + ((g2650) & (g2684) & (!g3265) & (g4628) & (!g3312)) + ((g2650) & (g2684) & (g3265) & (!g4628) & (g3312)) + ((g2650) & (g2684) & (g3265) & (g4628) & (g3312)));
	assign g4665 = (((!g2108) & (!g2116) & (g3602)) + ((!g2108) & (g2116) & (!g3602)) + ((g2108) & (!g2116) & (!g3602)) + ((g2108) & (g2116) & (g3602)));
	assign g4666 = (((!g830) & (!g1914) & (!g2396) & (!g4664) & (!g4665) & (key[234])) + ((!g830) & (!g1914) & (!g2396) & (!g4664) & (g4665) & (key[234])) + ((!g830) & (!g1914) & (!g2396) & (g4664) & (!g4665) & (key[234])) + ((!g830) & (!g1914) & (!g2396) & (g4664) & (g4665) & (key[234])) + ((!g830) & (!g1914) & (g2396) & (!g4664) & (!g4665) & (key[234])) + ((!g830) & (!g1914) & (g2396) & (!g4664) & (g4665) & (key[234])) + ((!g830) & (!g1914) & (g2396) & (g4664) & (!g4665) & (key[234])) + ((!g830) & (!g1914) & (g2396) & (g4664) & (g4665) & (key[234])) + ((!g830) & (g1914) & (!g2396) & (!g4664) & (!g4665) & (key[234])) + ((!g830) & (g1914) & (!g2396) & (!g4664) & (g4665) & (key[234])) + ((!g830) & (g1914) & (!g2396) & (g4664) & (!g4665) & (key[234])) + ((!g830) & (g1914) & (!g2396) & (g4664) & (g4665) & (key[234])) + ((!g830) & (g1914) & (g2396) & (!g4664) & (!g4665) & (key[234])) + ((!g830) & (g1914) & (g2396) & (!g4664) & (g4665) & (key[234])) + ((!g830) & (g1914) & (g2396) & (g4664) & (!g4665) & (key[234])) + ((!g830) & (g1914) & (g2396) & (g4664) & (g4665) & (key[234])) + ((g830) & (!g1914) & (!g2396) & (!g4664) & (g4665) & (!key[234])) + ((g830) & (!g1914) & (!g2396) & (!g4664) & (g4665) & (key[234])) + ((g830) & (!g1914) & (!g2396) & (g4664) & (g4665) & (!key[234])) + ((g830) & (!g1914) & (!g2396) & (g4664) & (g4665) & (key[234])) + ((g830) & (!g1914) & (g2396) & (!g4664) & (!g4665) & (!key[234])) + ((g830) & (!g1914) & (g2396) & (!g4664) & (!g4665) & (key[234])) + ((g830) & (!g1914) & (g2396) & (g4664) & (!g4665) & (!key[234])) + ((g830) & (!g1914) & (g2396) & (g4664) & (!g4665) & (key[234])) + ((g830) & (g1914) & (!g2396) & (g4664) & (!g4665) & (!key[234])) + ((g830) & (g1914) & (!g2396) & (g4664) & (!g4665) & (key[234])) + ((g830) & (g1914) & (!g2396) & (g4664) & (g4665) & (!key[234])) + ((g830) & (g1914) & (!g2396) & (g4664) & (g4665) & (key[234])) + ((g830) & (g1914) & (g2396) & (!g4664) & (!g4665) & (!key[234])) + ((g830) & (g1914) & (g2396) & (!g4664) & (!g4665) & (key[234])) + ((g830) & (g1914) & (g2396) & (!g4664) & (g4665) & (!key[234])) + ((g830) & (g1914) & (g2396) & (!g4664) & (g4665) & (key[234])));
	assign g4667 = (((!g1945) & (!g931) & (g3621)) + ((!g1945) & (g931) & (!g3621)) + ((g1945) & (!g931) & (!g3621)) + ((g1945) & (g931) & (g3621)));
	assign g4668 = (((!g3255) & (!g3297) & (!g4602) & (!g3265) & (g3312)) + ((!g3255) & (!g3297) & (!g4602) & (g3265) & (!g3312)) + ((!g3255) & (!g3297) & (g4602) & (!g3265) & (g3312)) + ((!g3255) & (!g3297) & (g4602) & (g3265) & (g3312)) + ((!g3255) & (g3297) & (!g4602) & (!g3265) & (!g3312)) + ((!g3255) & (g3297) & (!g4602) & (g3265) & (g3312)) + ((!g3255) & (g3297) & (g4602) & (!g3265) & (!g3312)) + ((!g3255) & (g3297) & (g4602) & (g3265) & (!g3312)) + ((g3255) & (!g3297) & (!g4602) & (!g3265) & (!g3312)) + ((g3255) & (!g3297) & (!g4602) & (g3265) & (!g3312)) + ((g3255) & (!g3297) & (g4602) & (!g3265) & (g3312)) + ((g3255) & (!g3297) & (g4602) & (g3265) & (!g3312)) + ((g3255) & (g3297) & (!g4602) & (!g3265) & (g3312)) + ((g3255) & (g3297) & (!g4602) & (g3265) & (g3312)) + ((g3255) & (g3297) & (g4602) & (!g3265) & (!g3312)) + ((g3255) & (g3297) & (g4602) & (g3265) & (g3312)));
	assign g4669 = (((!g830) & (!g1914) & (!g2399) & (!g4667) & (!g4668) & (key[10])) + ((!g830) & (!g1914) & (!g2399) & (!g4667) & (g4668) & (key[10])) + ((!g830) & (!g1914) & (!g2399) & (g4667) & (!g4668) & (key[10])) + ((!g830) & (!g1914) & (!g2399) & (g4667) & (g4668) & (key[10])) + ((!g830) & (!g1914) & (g2399) & (!g4667) & (!g4668) & (key[10])) + ((!g830) & (!g1914) & (g2399) & (!g4667) & (g4668) & (key[10])) + ((!g830) & (!g1914) & (g2399) & (g4667) & (!g4668) & (key[10])) + ((!g830) & (!g1914) & (g2399) & (g4667) & (g4668) & (key[10])) + ((!g830) & (g1914) & (!g2399) & (!g4667) & (!g4668) & (key[10])) + ((!g830) & (g1914) & (!g2399) & (!g4667) & (g4668) & (key[10])) + ((!g830) & (g1914) & (!g2399) & (g4667) & (!g4668) & (key[10])) + ((!g830) & (g1914) & (!g2399) & (g4667) & (g4668) & (key[10])) + ((!g830) & (g1914) & (g2399) & (!g4667) & (!g4668) & (key[10])) + ((!g830) & (g1914) & (g2399) & (!g4667) & (g4668) & (key[10])) + ((!g830) & (g1914) & (g2399) & (g4667) & (!g4668) & (key[10])) + ((!g830) & (g1914) & (g2399) & (g4667) & (g4668) & (key[10])) + ((g830) & (!g1914) & (!g2399) & (!g4667) & (g4668) & (!key[10])) + ((g830) & (!g1914) & (!g2399) & (!g4667) & (g4668) & (key[10])) + ((g830) & (!g1914) & (!g2399) & (g4667) & (g4668) & (!key[10])) + ((g830) & (!g1914) & (!g2399) & (g4667) & (g4668) & (key[10])) + ((g830) & (!g1914) & (g2399) & (!g4667) & (!g4668) & (!key[10])) + ((g830) & (!g1914) & (g2399) & (!g4667) & (!g4668) & (key[10])) + ((g830) & (!g1914) & (g2399) & (g4667) & (!g4668) & (!key[10])) + ((g830) & (!g1914) & (g2399) & (g4667) & (!g4668) & (key[10])) + ((g830) & (g1914) & (!g2399) & (g4667) & (!g4668) & (!key[10])) + ((g830) & (g1914) & (!g2399) & (g4667) & (!g4668) & (key[10])) + ((g830) & (g1914) & (!g2399) & (g4667) & (g4668) & (!key[10])) + ((g830) & (g1914) & (!g2399) & (g4667) & (g4668) & (key[10])) + ((g830) & (g1914) & (g2399) & (!g4667) & (!g4668) & (!key[10])) + ((g830) & (g1914) & (g2399) & (!g4667) & (!g4668) & (key[10])) + ((g830) & (g1914) & (g2399) & (!g4667) & (g4668) & (!key[10])) + ((g830) & (g1914) & (g2399) & (!g4667) & (g4668) & (key[10])));
	assign g4670 = (((!g2649) & (!g2683) & (!g3274) & (g3299) & (!g4607)) + ((!g2649) & (!g2683) & (!g3274) & (g3299) & (g4607)) + ((!g2649) & (!g2683) & (g3274) & (!g3299) & (!g4607)) + ((!g2649) & (!g2683) & (g3274) & (g3299) & (g4607)) + ((!g2649) & (g2683) & (!g3274) & (!g3299) & (!g4607)) + ((!g2649) & (g2683) & (!g3274) & (!g3299) & (g4607)) + ((!g2649) & (g2683) & (g3274) & (!g3299) & (g4607)) + ((!g2649) & (g2683) & (g3274) & (g3299) & (!g4607)) + ((g2649) & (!g2683) & (!g3274) & (!g3299) & (!g4607)) + ((g2649) & (!g2683) & (!g3274) & (g3299) & (g4607)) + ((g2649) & (!g2683) & (g3274) & (!g3299) & (!g4607)) + ((g2649) & (!g2683) & (g3274) & (!g3299) & (g4607)) + ((g2649) & (g2683) & (!g3274) & (!g3299) & (g4607)) + ((g2649) & (g2683) & (!g3274) & (g3299) & (!g4607)) + ((g2649) & (g2683) & (g3274) & (g3299) & (!g4607)) + ((g2649) & (g2683) & (g3274) & (g3299) & (g4607)));
	assign g4671 = (((!g2104) & (!g2118) & (g3669)) + ((!g2104) & (g2118) & (!g3669)) + ((g2104) & (!g2118) & (!g3669)) + ((g2104) & (g2118) & (g3669)));
	assign g8310 = (((!g5560) & (g5608) & (!g4672)) + ((!g5560) & (g5608) & (g4672)) + ((g5560) & (!g5608) & (g4672)) + ((g5560) & (g5608) & (g4672)));
	assign g4673 = (((!g830) & (!g1914) & (!g2402) & (!g4670) & (!g4671) & (g4672)) + ((!g830) & (!g1914) & (!g2402) & (!g4670) & (g4671) & (g4672)) + ((!g830) & (!g1914) & (!g2402) & (g4670) & (!g4671) & (g4672)) + ((!g830) & (!g1914) & (!g2402) & (g4670) & (g4671) & (g4672)) + ((!g830) & (!g1914) & (g2402) & (!g4670) & (!g4671) & (g4672)) + ((!g830) & (!g1914) & (g2402) & (!g4670) & (g4671) & (g4672)) + ((!g830) & (!g1914) & (g2402) & (g4670) & (!g4671) & (g4672)) + ((!g830) & (!g1914) & (g2402) & (g4670) & (g4671) & (g4672)) + ((!g830) & (g1914) & (!g2402) & (!g4670) & (!g4671) & (g4672)) + ((!g830) & (g1914) & (!g2402) & (!g4670) & (g4671) & (g4672)) + ((!g830) & (g1914) & (!g2402) & (g4670) & (!g4671) & (g4672)) + ((!g830) & (g1914) & (!g2402) & (g4670) & (g4671) & (g4672)) + ((!g830) & (g1914) & (g2402) & (!g4670) & (!g4671) & (g4672)) + ((!g830) & (g1914) & (g2402) & (!g4670) & (g4671) & (g4672)) + ((!g830) & (g1914) & (g2402) & (g4670) & (!g4671) & (g4672)) + ((!g830) & (g1914) & (g2402) & (g4670) & (g4671) & (g4672)) + ((g830) & (!g1914) & (!g2402) & (!g4670) & (g4671) & (!g4672)) + ((g830) & (!g1914) & (!g2402) & (!g4670) & (g4671) & (g4672)) + ((g830) & (!g1914) & (!g2402) & (g4670) & (g4671) & (!g4672)) + ((g830) & (!g1914) & (!g2402) & (g4670) & (g4671) & (g4672)) + ((g830) & (!g1914) & (g2402) & (!g4670) & (!g4671) & (!g4672)) + ((g830) & (!g1914) & (g2402) & (!g4670) & (!g4671) & (g4672)) + ((g830) & (!g1914) & (g2402) & (g4670) & (!g4671) & (!g4672)) + ((g830) & (!g1914) & (g2402) & (g4670) & (!g4671) & (g4672)) + ((g830) & (g1914) & (!g2402) & (g4670) & (!g4671) & (!g4672)) + ((g830) & (g1914) & (!g2402) & (g4670) & (!g4671) & (g4672)) + ((g830) & (g1914) & (!g2402) & (g4670) & (g4671) & (!g4672)) + ((g830) & (g1914) & (!g2402) & (g4670) & (g4671) & (g4672)) + ((g830) & (g1914) & (g2402) & (!g4670) & (!g4671) & (!g4672)) + ((g830) & (g1914) & (g2402) & (!g4670) & (!g4671) & (g4672)) + ((g830) & (g1914) & (g2402) & (!g4670) & (g4671) & (!g4672)) + ((g830) & (g1914) & (g2402) & (!g4670) & (g4671) & (g4672)));
	assign g4674 = (((!g3047) & (g3056) & (g4624)) + ((g3047) & (!g3056) & (g4624)) + ((g3047) & (g3056) & (!g4624)) + ((g3047) & (g3056) & (g4624)));
	assign g4675 = (((!g3009) & (!g3031) & (g3015) & (g3064) & (g4575)) + ((!g3009) & (g3031) & (!g3015) & (g3064) & (!g4575)) + ((!g3009) & (g3031) & (!g3015) & (g3064) & (g4575)) + ((!g3009) & (g3031) & (g3015) & (!g3064) & (g4575)) + ((!g3009) & (g3031) & (g3015) & (g3064) & (!g4575)) + ((!g3009) & (g3031) & (g3015) & (g3064) & (g4575)) + ((g3009) & (!g3031) & (!g3015) & (g3064) & (g4575)) + ((g3009) & (!g3031) & (g3015) & (g3064) & (!g4575)) + ((g3009) & (!g3031) & (g3015) & (g3064) & (g4575)) + ((g3009) & (g3031) & (!g3015) & (!g3064) & (g4575)) + ((g3009) & (g3031) & (!g3015) & (g3064) & (!g4575)) + ((g3009) & (g3031) & (!g3015) & (g3064) & (g4575)) + ((g3009) & (g3031) & (g3015) & (!g3064) & (!g4575)) + ((g3009) & (g3031) & (g3015) & (!g3064) & (g4575)) + ((g3009) & (g3031) & (g3015) & (g3064) & (!g4575)) + ((g3009) & (g3031) & (g3015) & (g3064) & (g4575)));
	assign g4676 = (((!g3084) & (!g3090) & (g4675)) + ((!g3084) & (g3090) & (!g4675)) + ((g3084) & (!g3090) & (!g4675)) + ((g3084) & (g3090) & (g4675)));
	assign g4677 = (((g1914) & (!g1888) & (!g1978) & (!g1912) & (g2045)) + ((g1914) & (!g1888) & (!g1978) & (g1912) & (g2045)) + ((g1914) & (!g1888) & (g1978) & (!g1912) & (!g2045)) + ((g1914) & (!g1888) & (g1978) & (g1912) & (!g2045)) + ((g1914) & (g1888) & (!g1978) & (!g1912) & (g2045)) + ((g1914) & (g1888) & (!g1978) & (g1912) & (!g2045)) + ((g1914) & (g1888) & (g1978) & (!g1912) & (!g2045)) + ((g1914) & (g1888) & (g1978) & (g1912) & (g2045)));
	assign g4678 = (((!g1914) & (!g1900) & (!g2028) & (!g1902) & (g2036)) + ((!g1914) & (!g1900) & (!g2028) & (g1902) & (g2036)) + ((!g1914) & (!g1900) & (g2028) & (!g1902) & (!g2036)) + ((!g1914) & (!g1900) & (g2028) & (g1902) & (!g2036)) + ((!g1914) & (g1900) & (!g2028) & (!g1902) & (g2036)) + ((!g1914) & (g1900) & (!g2028) & (g1902) & (!g2036)) + ((!g1914) & (g1900) & (g2028) & (!g1902) & (!g2036)) + ((!g1914) & (g1900) & (g2028) & (g1902) & (g2036)));
	assign g4679 = (((!g830) & (!g2408) & (!g4677) & (!g4678) & (key[202])) + ((!g830) & (!g2408) & (!g4677) & (g4678) & (key[202])) + ((!g830) & (!g2408) & (g4677) & (!g4678) & (key[202])) + ((!g830) & (!g2408) & (g4677) & (g4678) & (key[202])) + ((!g830) & (g2408) & (!g4677) & (!g4678) & (key[202])) + ((!g830) & (g2408) & (!g4677) & (g4678) & (key[202])) + ((!g830) & (g2408) & (g4677) & (!g4678) & (key[202])) + ((!g830) & (g2408) & (g4677) & (g4678) & (key[202])) + ((g830) & (!g2408) & (!g4677) & (g4678) & (!key[202])) + ((g830) & (!g2408) & (!g4677) & (g4678) & (key[202])) + ((g830) & (!g2408) & (g4677) & (!g4678) & (!key[202])) + ((g830) & (!g2408) & (g4677) & (!g4678) & (key[202])) + ((g830) & (!g2408) & (g4677) & (g4678) & (!key[202])) + ((g830) & (!g2408) & (g4677) & (g4678) & (key[202])) + ((g830) & (g2408) & (!g4677) & (!g4678) & (!key[202])) + ((g830) & (g2408) & (!g4677) & (!g4678) & (key[202])));
	assign g4680 = (((!g2108) & (!g2110) & (g3778)) + ((!g2108) & (g2110) & (!g3778)) + ((g2108) & (!g2110) & (!g3778)) + ((g2108) & (g2110) & (g3778)));
	assign g4681 = (((!g2648) & (!g2679) & (!g4613) & (!g3279) & (g3307)) + ((!g2648) & (!g2679) & (!g4613) & (g3279) & (!g3307)) + ((!g2648) & (!g2679) & (g4613) & (!g3279) & (g3307)) + ((!g2648) & (!g2679) & (g4613) & (g3279) & (g3307)) + ((!g2648) & (g2679) & (!g4613) & (!g3279) & (!g3307)) + ((!g2648) & (g2679) & (!g4613) & (g3279) & (g3307)) + ((!g2648) & (g2679) & (g4613) & (!g3279) & (!g3307)) + ((!g2648) & (g2679) & (g4613) & (g3279) & (!g3307)) + ((g2648) & (!g2679) & (!g4613) & (!g3279) & (!g3307)) + ((g2648) & (!g2679) & (!g4613) & (g3279) & (!g3307)) + ((g2648) & (!g2679) & (g4613) & (!g3279) & (g3307)) + ((g2648) & (!g2679) & (g4613) & (g3279) & (!g3307)) + ((g2648) & (g2679) & (!g4613) & (!g3279) & (g3307)) + ((g2648) & (g2679) & (!g4613) & (g3279) & (g3307)) + ((g2648) & (g2679) & (g4613) & (!g3279) & (!g3307)) + ((g2648) & (g2679) & (g4613) & (g3279) & (g3307)));
	assign g4682 = (((!g830) & (!g1914) & (!g2413) & (!g4680) & (!g4681) & (key[138])) + ((!g830) & (!g1914) & (!g2413) & (!g4680) & (g4681) & (key[138])) + ((!g830) & (!g1914) & (!g2413) & (g4680) & (!g4681) & (key[138])) + ((!g830) & (!g1914) & (!g2413) & (g4680) & (g4681) & (key[138])) + ((!g830) & (!g1914) & (g2413) & (!g4680) & (!g4681) & (key[138])) + ((!g830) & (!g1914) & (g2413) & (!g4680) & (g4681) & (key[138])) + ((!g830) & (!g1914) & (g2413) & (g4680) & (!g4681) & (key[138])) + ((!g830) & (!g1914) & (g2413) & (g4680) & (g4681) & (key[138])) + ((!g830) & (g1914) & (!g2413) & (!g4680) & (!g4681) & (key[138])) + ((!g830) & (g1914) & (!g2413) & (!g4680) & (g4681) & (key[138])) + ((!g830) & (g1914) & (!g2413) & (g4680) & (!g4681) & (key[138])) + ((!g830) & (g1914) & (!g2413) & (g4680) & (g4681) & (key[138])) + ((!g830) & (g1914) & (g2413) & (!g4680) & (!g4681) & (key[138])) + ((!g830) & (g1914) & (g2413) & (!g4680) & (g4681) & (key[138])) + ((!g830) & (g1914) & (g2413) & (g4680) & (!g4681) & (key[138])) + ((!g830) & (g1914) & (g2413) & (g4680) & (g4681) & (key[138])) + ((g830) & (!g1914) & (!g2413) & (!g4680) & (g4681) & (!key[138])) + ((g830) & (!g1914) & (!g2413) & (!g4680) & (g4681) & (key[138])) + ((g830) & (!g1914) & (!g2413) & (g4680) & (g4681) & (!key[138])) + ((g830) & (!g1914) & (!g2413) & (g4680) & (g4681) & (key[138])) + ((g830) & (!g1914) & (g2413) & (!g4680) & (!g4681) & (!key[138])) + ((g830) & (!g1914) & (g2413) & (!g4680) & (!g4681) & (key[138])) + ((g830) & (!g1914) & (g2413) & (g4680) & (!g4681) & (!key[138])) + ((g830) & (!g1914) & (g2413) & (g4680) & (!g4681) & (key[138])) + ((g830) & (g1914) & (!g2413) & (g4680) & (!g4681) & (!key[138])) + ((g830) & (g1914) & (!g2413) & (g4680) & (!g4681) & (key[138])) + ((g830) & (g1914) & (!g2413) & (g4680) & (g4681) & (!key[138])) + ((g830) & (g1914) & (!g2413) & (g4680) & (g4681) & (key[138])) + ((g830) & (g1914) & (g2413) & (!g4680) & (!g4681) & (!key[138])) + ((g830) & (g1914) & (g2413) & (!g4680) & (!g4681) & (key[138])) + ((g830) & (g1914) & (g2413) & (!g4680) & (g4681) & (!key[138])) + ((g830) & (g1914) & (g2413) & (!g4680) & (g4681) & (key[138])));
	assign g4683 = (((g1914) & (!g1894) & (!g2034) & (!g1902) & (g2036)) + ((g1914) & (!g1894) & (!g2034) & (g1902) & (g2036)) + ((g1914) & (!g1894) & (g2034) & (!g1902) & (!g2036)) + ((g1914) & (!g1894) & (g2034) & (g1902) & (!g2036)) + ((g1914) & (g1894) & (!g2034) & (!g1902) & (g2036)) + ((g1914) & (g1894) & (!g2034) & (g1902) & (!g2036)) + ((g1914) & (g1894) & (g2034) & (!g1902) & (!g2036)) + ((g1914) & (g1894) & (g2034) & (g1902) & (g2036)));
	assign g4684 = (((!g1914) & (!g1906) & (!g1940) & (!g1912) & (g2045)) + ((!g1914) & (!g1906) & (!g1940) & (g1912) & (g2045)) + ((!g1914) & (!g1906) & (g1940) & (!g1912) & (!g2045)) + ((!g1914) & (!g1906) & (g1940) & (g1912) & (!g2045)) + ((!g1914) & (g1906) & (!g1940) & (!g1912) & (g2045)) + ((!g1914) & (g1906) & (!g1940) & (g1912) & (!g2045)) + ((!g1914) & (g1906) & (g1940) & (!g1912) & (!g2045)) + ((!g1914) & (g1906) & (g1940) & (g1912) & (g2045)));
	assign g4685 = (((!g830) & (!g2416) & (!g4683) & (!g4684) & (nonce[42])) + ((!g830) & (!g2416) & (!g4683) & (g4684) & (nonce[42])) + ((!g830) & (!g2416) & (g4683) & (!g4684) & (nonce[42])) + ((!g830) & (!g2416) & (g4683) & (g4684) & (nonce[42])) + ((!g830) & (g2416) & (!g4683) & (!g4684) & (nonce[42])) + ((!g830) & (g2416) & (!g4683) & (g4684) & (nonce[42])) + ((!g830) & (g2416) & (g4683) & (!g4684) & (nonce[42])) + ((!g830) & (g2416) & (g4683) & (g4684) & (nonce[42])) + ((g830) & (!g2416) & (!g4683) & (g4684) & (!nonce[42])) + ((g830) & (!g2416) & (!g4683) & (g4684) & (nonce[42])) + ((g830) & (!g2416) & (g4683) & (!g4684) & (!nonce[42])) + ((g830) & (!g2416) & (g4683) & (!g4684) & (nonce[42])) + ((g830) & (!g2416) & (g4683) & (g4684) & (!nonce[42])) + ((g830) & (!g2416) & (g4683) & (g4684) & (nonce[42])) + ((g830) & (g2416) & (!g4683) & (!g4684) & (!nonce[42])) + ((g830) & (g2416) & (!g4683) & (!g4684) & (nonce[42])));
	assign g4686 = (((!g3061) & (g3064) & (g4634)) + ((g3061) & (!g3064) & (g4634)) + ((g3061) & (g3064) & (!g4634)) + ((g3061) & (g3064) & (g4634)));
	assign g4687 = (((!g3018) & (!g3044) & (g3020) & (g3056) & (g4587)) + ((!g3018) & (g3044) & (!g3020) & (g3056) & (!g4587)) + ((!g3018) & (g3044) & (!g3020) & (g3056) & (g4587)) + ((!g3018) & (g3044) & (g3020) & (!g3056) & (g4587)) + ((!g3018) & (g3044) & (g3020) & (g3056) & (!g4587)) + ((!g3018) & (g3044) & (g3020) & (g3056) & (g4587)) + ((g3018) & (!g3044) & (!g3020) & (g3056) & (g4587)) + ((g3018) & (!g3044) & (g3020) & (g3056) & (!g4587)) + ((g3018) & (!g3044) & (g3020) & (g3056) & (g4587)) + ((g3018) & (g3044) & (!g3020) & (!g3056) & (g4587)) + ((g3018) & (g3044) & (!g3020) & (g3056) & (!g4587)) + ((g3018) & (g3044) & (!g3020) & (g3056) & (g4587)) + ((g3018) & (g3044) & (g3020) & (!g3056) & (!g4587)) + ((g3018) & (g3044) & (g3020) & (!g3056) & (g4587)) + ((g3018) & (g3044) & (g3020) & (g3056) & (!g4587)) + ((g3018) & (g3044) & (g3020) & (g3056) & (g4587)));
	assign g4688 = (((!g3093) & (!g3095) & (g4687)) + ((!g3093) & (g3095) & (!g4687)) + ((g3093) & (!g3095) & (!g4687)) + ((g3093) & (g3095) & (g4687)));
	assign g4689 = (((!g1303) & (!g1337) & (!g4636) & (!g2623) & (g2653)) + ((!g1303) & (!g1337) & (!g4636) & (g2623) & (g2653)) + ((!g1303) & (!g1337) & (g4636) & (!g2623) & (g2653)) + ((!g1303) & (!g1337) & (g4636) & (g2623) & (!g2653)) + ((!g1303) & (g1337) & (!g4636) & (!g2623) & (!g2653)) + ((!g1303) & (g1337) & (!g4636) & (g2623) & (!g2653)) + ((!g1303) & (g1337) & (g4636) & (!g2623) & (!g2653)) + ((!g1303) & (g1337) & (g4636) & (g2623) & (g2653)) + ((g1303) & (!g1337) & (!g4636) & (!g2623) & (g2653)) + ((g1303) & (!g1337) & (!g4636) & (g2623) & (!g2653)) + ((g1303) & (!g1337) & (g4636) & (!g2623) & (!g2653)) + ((g1303) & (!g1337) & (g4636) & (g2623) & (!g2653)) + ((g1303) & (g1337) & (!g4636) & (!g2623) & (!g2653)) + ((g1303) & (g1337) & (!g4636) & (g2623) & (g2653)) + ((g1303) & (g1337) & (g4636) & (!g2623) & (g2653)) + ((g1303) & (g1337) & (g4636) & (g2623) & (g2653)));
	assign g4690 = (((!g2614) & (!g2657) & (!g2620) & (g2672) & (!g4638)) + ((!g2614) & (!g2657) & (!g2620) & (g2672) & (g4638)) + ((!g2614) & (!g2657) & (g2620) & (!g2672) & (g4638)) + ((!g2614) & (!g2657) & (g2620) & (g2672) & (!g4638)) + ((!g2614) & (g2657) & (!g2620) & (!g2672) & (!g4638)) + ((!g2614) & (g2657) & (!g2620) & (!g2672) & (g4638)) + ((!g2614) & (g2657) & (g2620) & (!g2672) & (!g4638)) + ((!g2614) & (g2657) & (g2620) & (g2672) & (g4638)) + ((g2614) & (!g2657) & (!g2620) & (!g2672) & (g4638)) + ((g2614) & (!g2657) & (!g2620) & (g2672) & (!g4638)) + ((g2614) & (!g2657) & (g2620) & (!g2672) & (!g4638)) + ((g2614) & (!g2657) & (g2620) & (!g2672) & (g4638)) + ((g2614) & (g2657) & (!g2620) & (!g2672) & (!g4638)) + ((g2614) & (g2657) & (!g2620) & (g2672) & (g4638)) + ((g2614) & (g2657) & (g2620) & (g2672) & (!g4638)) + ((g2614) & (g2657) & (g2620) & (g2672) & (g4638)));
	assign g4691 = (((!g830) & (!g1914) & (!g2423) & (!g4689) & (!g4690) & (key[56])) + ((!g830) & (!g1914) & (!g2423) & (!g4689) & (g4690) & (key[56])) + ((!g830) & (!g1914) & (!g2423) & (g4689) & (!g4690) & (key[56])) + ((!g830) & (!g1914) & (!g2423) & (g4689) & (g4690) & (key[56])) + ((!g830) & (!g1914) & (g2423) & (!g4689) & (!g4690) & (key[56])) + ((!g830) & (!g1914) & (g2423) & (!g4689) & (g4690) & (key[56])) + ((!g830) & (!g1914) & (g2423) & (g4689) & (!g4690) & (key[56])) + ((!g830) & (!g1914) & (g2423) & (g4689) & (g4690) & (key[56])) + ((!g830) & (g1914) & (!g2423) & (!g4689) & (!g4690) & (key[56])) + ((!g830) & (g1914) & (!g2423) & (!g4689) & (g4690) & (key[56])) + ((!g830) & (g1914) & (!g2423) & (g4689) & (!g4690) & (key[56])) + ((!g830) & (g1914) & (!g2423) & (g4689) & (g4690) & (key[56])) + ((!g830) & (g1914) & (g2423) & (!g4689) & (!g4690) & (key[56])) + ((!g830) & (g1914) & (g2423) & (!g4689) & (g4690) & (key[56])) + ((!g830) & (g1914) & (g2423) & (g4689) & (!g4690) & (key[56])) + ((!g830) & (g1914) & (g2423) & (g4689) & (g4690) & (key[56])) + ((g830) & (!g1914) & (!g2423) & (!g4689) & (g4690) & (!key[56])) + ((g830) & (!g1914) & (!g2423) & (!g4689) & (g4690) & (key[56])) + ((g830) & (!g1914) & (!g2423) & (g4689) & (g4690) & (!key[56])) + ((g830) & (!g1914) & (!g2423) & (g4689) & (g4690) & (key[56])) + ((g830) & (!g1914) & (g2423) & (!g4689) & (!g4690) & (!key[56])) + ((g830) & (!g1914) & (g2423) & (!g4689) & (!g4690) & (key[56])) + ((g830) & (!g1914) & (g2423) & (g4689) & (!g4690) & (!key[56])) + ((g830) & (!g1914) & (g2423) & (g4689) & (!g4690) & (key[56])) + ((g830) & (g1914) & (!g2423) & (g4689) & (!g4690) & (!key[56])) + ((g830) & (g1914) & (!g2423) & (g4689) & (!g4690) & (key[56])) + ((g830) & (g1914) & (!g2423) & (g4689) & (g4690) & (!key[56])) + ((g830) & (g1914) & (!g2423) & (g4689) & (g4690) & (key[56])) + ((g830) & (g1914) & (g2423) & (!g4689) & (!g4690) & (!key[56])) + ((g830) & (g1914) & (g2423) & (!g4689) & (!g4690) & (key[56])) + ((g830) & (g1914) & (g2423) & (!g4689) & (g4690) & (!key[56])) + ((g830) & (g1914) & (g2423) & (!g4689) & (g4690) & (key[56])));
	assign g4692 = (((!g3751) & (!g3752)));
	assign g4693 = (((!g1967) & (!g2434) & (!g4692)) + ((!g1967) & (g2434) & (g4692)) + ((g1967) & (!g2434) & (g4692)) + ((g1967) & (g2434) & (!g4692)));
	assign g4694 = (((!g830) & (!g2424) & (!g6566) & (key[88])) + ((!g830) & (!g2424) & (g6566) & (key[88])) + ((!g830) & (g2424) & (!g6566) & (key[88])) + ((!g830) & (g2424) & (g6566) & (key[88])) + ((g830) & (!g2424) & (g6566) & (!key[88])) + ((g830) & (!g2424) & (g6566) & (key[88])) + ((g830) & (g2424) & (!g6566) & (!key[88])) + ((g830) & (g2424) & (!g6566) & (key[88])));
	assign g4695 = (((!g4646) & (!g2614) & (!g2637) & (!g2657) & (g2661)) + ((!g4646) & (!g2614) & (!g2637) & (g2657) & (!g2661)) + ((!g4646) & (!g2614) & (g2637) & (!g2657) & (g2661)) + ((!g4646) & (!g2614) & (g2637) & (g2657) & (!g2661)) + ((!g4646) & (g2614) & (!g2637) & (!g2657) & (g2661)) + ((!g4646) & (g2614) & (!g2637) & (g2657) & (!g2661)) + ((!g4646) & (g2614) & (g2637) & (!g2657) & (!g2661)) + ((!g4646) & (g2614) & (g2637) & (g2657) & (g2661)) + ((g4646) & (!g2614) & (!g2637) & (!g2657) & (g2661)) + ((g4646) & (!g2614) & (!g2637) & (g2657) & (!g2661)) + ((g4646) & (!g2614) & (g2637) & (!g2657) & (!g2661)) + ((g4646) & (!g2614) & (g2637) & (g2657) & (g2661)) + ((g4646) & (g2614) & (!g2637) & (!g2657) & (!g2661)) + ((g4646) & (g2614) & (!g2637) & (g2657) & (g2661)) + ((g4646) & (g2614) & (g2637) & (!g2657) & (!g2661)) + ((g4646) & (g2614) & (g2637) & (g2657) & (g2661)));
	assign g8311 = (((!g5560) & (g5609) & (!g4696)) + ((!g5560) & (g5609) & (g4696)) + ((g5560) & (!g5609) & (g4696)) + ((g5560) & (g5609) & (g4696)));
	assign g4697 = (((!g830) & (!g2426) & (!g6555) & (g4696)) + ((!g830) & (!g2426) & (g6555) & (g4696)) + ((!g830) & (g2426) & (!g6555) & (g4696)) + ((!g830) & (g2426) & (g6555) & (g4696)) + ((g830) & (!g2426) & (g6555) & (!g4696)) + ((g830) & (!g2426) & (g6555) & (g4696)) + ((g830) & (g2426) & (!g6555) & (!g4696)) + ((g830) & (g2426) & (!g6555) & (g4696)));
	assign g4698 = (((!g3489) & (!g3490)));
	assign g4699 = (((!g2003) & (!g2468) & (!g4698)) + ((!g2003) & (g2468) & (g4698)) + ((g2003) & (!g2468) & (g4698)) + ((g2003) & (g2468) & (!g4698)));
	assign g4700 = (((!g830) & (!g2427) & (!g6544) & (key[184])) + ((!g830) & (!g2427) & (g6544) & (key[184])) + ((!g830) & (g2427) & (!g6544) & (key[184])) + ((!g830) & (g2427) & (g6544) & (key[184])) + ((g830) & (!g2427) & (g6544) & (!key[184])) + ((g830) & (!g2427) & (g6544) & (key[184])) + ((g830) & (g2427) & (!g6544) & (!key[184])) + ((g830) & (g2427) & (!g6544) & (key[184])));
	assign g4701 = (((!g1945) & (g931) & (g3621)) + ((g1945) & (!g931) & (g3621)) + ((g1945) & (g931) & (!g3621)) + ((g1945) & (g931) & (g3621)));
	assign g4702 = (((!g3255) & (!g3297) & (!g4602) & (g3265) & (g3312)) + ((!g3255) & (g3297) & (!g4602) & (!g3265) & (g3312)) + ((!g3255) & (g3297) & (!g4602) & (g3265) & (!g3312)) + ((!g3255) & (g3297) & (!g4602) & (g3265) & (g3312)) + ((!g3255) & (g3297) & (g4602) & (!g3265) & (g3312)) + ((!g3255) & (g3297) & (g4602) & (g3265) & (g3312)) + ((g3255) & (!g3297) & (!g4602) & (!g3265) & (g3312)) + ((g3255) & (!g3297) & (!g4602) & (g3265) & (g3312)) + ((g3255) & (!g3297) & (g4602) & (g3265) & (g3312)) + ((g3255) & (g3297) & (!g4602) & (!g3265) & (!g3312)) + ((g3255) & (g3297) & (!g4602) & (!g3265) & (g3312)) + ((g3255) & (g3297) & (!g4602) & (g3265) & (!g3312)) + ((g3255) & (g3297) & (!g4602) & (g3265) & (g3312)) + ((g3255) & (g3297) & (g4602) & (!g3265) & (g3312)) + ((g3255) & (g3297) & (g4602) & (g3265) & (!g3312)) + ((g3255) & (g3297) & (g4602) & (g3265) & (g3312)));
	assign g4703 = (((!g830) & (key[11]) & (!g1914) & (!g4702) & (!g1947) & (!g5676)) + ((!g830) & (key[11]) & (!g1914) & (!g4702) & (!g1947) & (g5676)) + ((!g830) & (key[11]) & (!g1914) & (!g4702) & (g1947) & (!g5676)) + ((!g830) & (key[11]) & (!g1914) & (!g4702) & (g1947) & (g5676)) + ((!g830) & (key[11]) & (!g1914) & (g4702) & (!g1947) & (!g5676)) + ((!g830) & (key[11]) & (!g1914) & (g4702) & (!g1947) & (g5676)) + ((!g830) & (key[11]) & (!g1914) & (g4702) & (g1947) & (!g5676)) + ((!g830) & (key[11]) & (!g1914) & (g4702) & (g1947) & (g5676)) + ((!g830) & (key[11]) & (g1914) & (!g4702) & (!g1947) & (!g5676)) + ((!g830) & (key[11]) & (g1914) & (!g4702) & (!g1947) & (g5676)) + ((!g830) & (key[11]) & (g1914) & (!g4702) & (g1947) & (!g5676)) + ((!g830) & (key[11]) & (g1914) & (!g4702) & (g1947) & (g5676)) + ((!g830) & (key[11]) & (g1914) & (g4702) & (!g1947) & (!g5676)) + ((!g830) & (key[11]) & (g1914) & (g4702) & (!g1947) & (g5676)) + ((!g830) & (key[11]) & (g1914) & (g4702) & (g1947) & (!g5676)) + ((!g830) & (key[11]) & (g1914) & (g4702) & (g1947) & (g5676)) + ((g830) & (!key[11]) & (!g1914) & (!g4702) & (!g1947) & (!g5676)) + ((g830) & (!key[11]) & (!g1914) & (!g4702) & (g1947) & (!g5676)) + ((g830) & (!key[11]) & (!g1914) & (g4702) & (!g1947) & (g5676)) + ((g830) & (!key[11]) & (!g1914) & (g4702) & (g1947) & (g5676)) + ((g830) & (!key[11]) & (g1914) & (!g4702) & (!g1947) & (!g5676)) + ((g830) & (!key[11]) & (g1914) & (!g4702) & (g1947) & (g5676)) + ((g830) & (!key[11]) & (g1914) & (g4702) & (!g1947) & (!g5676)) + ((g830) & (!key[11]) & (g1914) & (g4702) & (g1947) & (g5676)) + ((g830) & (key[11]) & (!g1914) & (!g4702) & (!g1947) & (!g5676)) + ((g830) & (key[11]) & (!g1914) & (!g4702) & (g1947) & (!g5676)) + ((g830) & (key[11]) & (!g1914) & (g4702) & (!g1947) & (g5676)) + ((g830) & (key[11]) & (!g1914) & (g4702) & (g1947) & (g5676)) + ((g830) & (key[11]) & (g1914) & (!g4702) & (!g1947) & (!g5676)) + ((g830) & (key[11]) & (g1914) & (!g4702) & (g1947) & (g5676)) + ((g830) & (key[11]) & (g1914) & (g4702) & (!g1947) & (!g5676)) + ((g830) & (key[11]) & (g1914) & (g4702) & (g1947) & (g5676)));
	assign g4704 = (((!g2426) & (!g2518) & (!g3086) & (g3116) & (!g4658)) + ((!g2426) & (!g2518) & (!g3086) & (g3116) & (g4658)) + ((!g2426) & (!g2518) & (g3086) & (!g3116) & (g4658)) + ((!g2426) & (!g2518) & (g3086) & (g3116) & (!g4658)) + ((!g2426) & (g2518) & (!g3086) & (!g3116) & (!g4658)) + ((!g2426) & (g2518) & (!g3086) & (!g3116) & (g4658)) + ((!g2426) & (g2518) & (g3086) & (!g3116) & (!g4658)) + ((!g2426) & (g2518) & (g3086) & (g3116) & (g4658)) + ((g2426) & (!g2518) & (!g3086) & (!g3116) & (g4658)) + ((g2426) & (!g2518) & (!g3086) & (g3116) & (!g4658)) + ((g2426) & (!g2518) & (g3086) & (!g3116) & (!g4658)) + ((g2426) & (!g2518) & (g3086) & (!g3116) & (g4658)) + ((g2426) & (g2518) & (!g3086) & (!g3116) & (!g4658)) + ((g2426) & (g2518) & (!g3086) & (g3116) & (g4658)) + ((g2426) & (g2518) & (g3086) & (g3116) & (!g4658)) + ((g2426) & (g2518) & (g3086) & (g3116) & (g4658)));
	assign g4705 = (((!g2423) & (!g2515) & (!g3080) & (g3125) & (!g4659)) + ((!g2423) & (!g2515) & (!g3080) & (g3125) & (g4659)) + ((!g2423) & (!g2515) & (g3080) & (!g3125) & (g4659)) + ((!g2423) & (!g2515) & (g3080) & (g3125) & (!g4659)) + ((!g2423) & (g2515) & (!g3080) & (!g3125) & (!g4659)) + ((!g2423) & (g2515) & (!g3080) & (!g3125) & (g4659)) + ((!g2423) & (g2515) & (g3080) & (!g3125) & (!g4659)) + ((!g2423) & (g2515) & (g3080) & (g3125) & (g4659)) + ((g2423) & (!g2515) & (!g3080) & (!g3125) & (g4659)) + ((g2423) & (!g2515) & (!g3080) & (g3125) & (!g4659)) + ((g2423) & (!g2515) & (g3080) & (!g3125) & (!g4659)) + ((g2423) & (!g2515) & (g3080) & (!g3125) & (g4659)) + ((g2423) & (g2515) & (!g3080) & (!g3125) & (!g4659)) + ((g2423) & (g2515) & (!g3080) & (g3125) & (g4659)) + ((g2423) & (g2515) & (g3080) & (g3125) & (!g4659)) + ((g2423) & (g2515) & (g3080) & (g3125) & (g4659)));
	assign g4706 = (((!g830) & (!g1914) & (!g2450) & (!g4704) & (!g4705)) + ((!g830) & (!g1914) & (!g2450) & (!g4704) & (g4705)) + ((!g830) & (!g1914) & (!g2450) & (g4704) & (!g4705)) + ((!g830) & (!g1914) & (!g2450) & (g4704) & (g4705)) + ((!g830) & (!g1914) & (g2450) & (!g4704) & (!g4705)) + ((!g830) & (!g1914) & (g2450) & (!g4704) & (g4705)) + ((!g830) & (!g1914) & (g2450) & (g4704) & (!g4705)) + ((!g830) & (!g1914) & (g2450) & (g4704) & (g4705)) + ((!g830) & (g1914) & (!g2450) & (!g4704) & (!g4705)) + ((!g830) & (g1914) & (!g2450) & (!g4704) & (g4705)) + ((!g830) & (g1914) & (!g2450) & (g4704) & (!g4705)) + ((!g830) & (g1914) & (!g2450) & (g4704) & (g4705)) + ((!g830) & (g1914) & (g2450) & (!g4704) & (!g4705)) + ((!g830) & (g1914) & (g2450) & (!g4704) & (g4705)) + ((!g830) & (g1914) & (g2450) & (g4704) & (!g4705)) + ((!g830) & (g1914) & (g2450) & (g4704) & (g4705)) + ((g830) & (!g1914) & (!g2450) & (!g4704) & (g4705)) + ((g830) & (!g1914) & (!g2450) & (g4704) & (g4705)) + ((g830) & (!g1914) & (g2450) & (!g4704) & (!g4705)) + ((g830) & (!g1914) & (g2450) & (g4704) & (!g4705)) + ((g830) & (g1914) & (!g2450) & (g4704) & (!g4705)) + ((g830) & (g1914) & (!g2450) & (g4704) & (g4705)) + ((g830) & (g1914) & (g2450) & (!g4704) & (!g4705)) + ((g830) & (g1914) & (g2450) & (!g4704) & (g4705)));
	assign g4707 = (((!g2649) & (!g2683) & (g3274) & (g3299) & (!g4607)) + ((!g2649) & (g2683) & (!g3274) & (g3299) & (!g4607)) + ((!g2649) & (g2683) & (!g3274) & (g3299) & (g4607)) + ((!g2649) & (g2683) & (g3274) & (!g3299) & (!g4607)) + ((!g2649) & (g2683) & (g3274) & (g3299) & (!g4607)) + ((!g2649) & (g2683) & (g3274) & (g3299) & (g4607)) + ((g2649) & (!g2683) & (!g3274) & (g3299) & (!g4607)) + ((g2649) & (!g2683) & (g3274) & (g3299) & (!g4607)) + ((g2649) & (!g2683) & (g3274) & (g3299) & (g4607)) + ((g2649) & (g2683) & (!g3274) & (!g3299) & (!g4607)) + ((g2649) & (g2683) & (!g3274) & (g3299) & (!g4607)) + ((g2649) & (g2683) & (!g3274) & (g3299) & (g4607)) + ((g2649) & (g2683) & (g3274) & (!g3299) & (!g4607)) + ((g2649) & (g2683) & (g3274) & (!g3299) & (g4607)) + ((g2649) & (g2683) & (g3274) & (g3299) & (!g4607)) + ((g2649) & (g2683) & (g3274) & (g3299) & (g4607)));
	assign g4708 = (((!g2104) & (g2118) & (g3669)) + ((g2104) & (!g2118) & (g3669)) + ((g2104) & (g2118) & (!g3669)) + ((g2104) & (g2118) & (g3669)));
	assign g8312 = (((!g5560) & (g5610) & (!g4709)) + ((!g5560) & (g5610) & (g4709)) + ((g5560) & (!g5610) & (g4709)) + ((g5560) & (g5610) & (g4709)));
	assign g4710 = (((!g830) & (g4709) & (!g1914) & (!g4707) & (!g2153) & (!g5678)) + ((!g830) & (g4709) & (!g1914) & (!g4707) & (!g2153) & (g5678)) + ((!g830) & (g4709) & (!g1914) & (!g4707) & (g2153) & (!g5678)) + ((!g830) & (g4709) & (!g1914) & (!g4707) & (g2153) & (g5678)) + ((!g830) & (g4709) & (!g1914) & (g4707) & (!g2153) & (!g5678)) + ((!g830) & (g4709) & (!g1914) & (g4707) & (!g2153) & (g5678)) + ((!g830) & (g4709) & (!g1914) & (g4707) & (g2153) & (!g5678)) + ((!g830) & (g4709) & (!g1914) & (g4707) & (g2153) & (g5678)) + ((!g830) & (g4709) & (g1914) & (!g4707) & (!g2153) & (!g5678)) + ((!g830) & (g4709) & (g1914) & (!g4707) & (!g2153) & (g5678)) + ((!g830) & (g4709) & (g1914) & (!g4707) & (g2153) & (!g5678)) + ((!g830) & (g4709) & (g1914) & (!g4707) & (g2153) & (g5678)) + ((!g830) & (g4709) & (g1914) & (g4707) & (!g2153) & (!g5678)) + ((!g830) & (g4709) & (g1914) & (g4707) & (!g2153) & (g5678)) + ((!g830) & (g4709) & (g1914) & (g4707) & (g2153) & (!g5678)) + ((!g830) & (g4709) & (g1914) & (g4707) & (g2153) & (g5678)) + ((g830) & (!g4709) & (!g1914) & (!g4707) & (!g2153) & (!g5678)) + ((g830) & (!g4709) & (!g1914) & (!g4707) & (g2153) & (g5678)) + ((g830) & (!g4709) & (!g1914) & (g4707) & (!g2153) & (!g5678)) + ((g830) & (!g4709) & (!g1914) & (g4707) & (g2153) & (g5678)) + ((g830) & (!g4709) & (g1914) & (!g4707) & (!g2153) & (!g5678)) + ((g830) & (!g4709) & (g1914) & (!g4707) & (g2153) & (!g5678)) + ((g830) & (!g4709) & (g1914) & (g4707) & (!g2153) & (g5678)) + ((g830) & (!g4709) & (g1914) & (g4707) & (g2153) & (g5678)) + ((g830) & (g4709) & (!g1914) & (!g4707) & (!g2153) & (!g5678)) + ((g830) & (g4709) & (!g1914) & (!g4707) & (g2153) & (g5678)) + ((g830) & (g4709) & (!g1914) & (g4707) & (!g2153) & (!g5678)) + ((g830) & (g4709) & (!g1914) & (g4707) & (g2153) & (g5678)) + ((g830) & (g4709) & (g1914) & (!g4707) & (!g2153) & (!g5678)) + ((g830) & (g4709) & (g1914) & (!g4707) & (g2153) & (!g5678)) + ((g830) & (g4709) & (g1914) & (g4707) & (!g2153) & (g5678)) + ((g830) & (g4709) & (g1914) & (g4707) & (g2153) & (g5678)));
	assign g4711 = (((!g2108) & (g2110) & (g3778)) + ((g2108) & (!g2110) & (g3778)) + ((g2108) & (g2110) & (!g3778)) + ((g2108) & (g2110) & (g3778)));
	assign g4712 = (((!g2648) & (!g2679) & (!g4613) & (g3279) & (g3307)) + ((!g2648) & (g2679) & (!g4613) & (!g3279) & (g3307)) + ((!g2648) & (g2679) & (!g4613) & (g3279) & (!g3307)) + ((!g2648) & (g2679) & (!g4613) & (g3279) & (g3307)) + ((!g2648) & (g2679) & (g4613) & (!g3279) & (g3307)) + ((!g2648) & (g2679) & (g4613) & (g3279) & (g3307)) + ((g2648) & (!g2679) & (!g4613) & (!g3279) & (g3307)) + ((g2648) & (!g2679) & (!g4613) & (g3279) & (g3307)) + ((g2648) & (!g2679) & (g4613) & (g3279) & (g3307)) + ((g2648) & (g2679) & (!g4613) & (!g3279) & (!g3307)) + ((g2648) & (g2679) & (!g4613) & (!g3279) & (g3307)) + ((g2648) & (g2679) & (!g4613) & (g3279) & (!g3307)) + ((g2648) & (g2679) & (!g4613) & (g3279) & (g3307)) + ((g2648) & (g2679) & (g4613) & (!g3279) & (g3307)) + ((g2648) & (g2679) & (g4613) & (g3279) & (!g3307)) + ((g2648) & (g2679) & (g4613) & (g3279) & (g3307)));
	assign g4713 = (((!g830) & (key[139]) & (!g1914) & (!g4712) & (!g2144) & (!g5679)) + ((!g830) & (key[139]) & (!g1914) & (!g4712) & (!g2144) & (g5679)) + ((!g830) & (key[139]) & (!g1914) & (!g4712) & (g2144) & (!g5679)) + ((!g830) & (key[139]) & (!g1914) & (!g4712) & (g2144) & (g5679)) + ((!g830) & (key[139]) & (!g1914) & (g4712) & (!g2144) & (!g5679)) + ((!g830) & (key[139]) & (!g1914) & (g4712) & (!g2144) & (g5679)) + ((!g830) & (key[139]) & (!g1914) & (g4712) & (g2144) & (!g5679)) + ((!g830) & (key[139]) & (!g1914) & (g4712) & (g2144) & (g5679)) + ((!g830) & (key[139]) & (g1914) & (!g4712) & (!g2144) & (!g5679)) + ((!g830) & (key[139]) & (g1914) & (!g4712) & (!g2144) & (g5679)) + ((!g830) & (key[139]) & (g1914) & (!g4712) & (g2144) & (!g5679)) + ((!g830) & (key[139]) & (g1914) & (!g4712) & (g2144) & (g5679)) + ((!g830) & (key[139]) & (g1914) & (g4712) & (!g2144) & (!g5679)) + ((!g830) & (key[139]) & (g1914) & (g4712) & (!g2144) & (g5679)) + ((!g830) & (key[139]) & (g1914) & (g4712) & (g2144) & (!g5679)) + ((!g830) & (key[139]) & (g1914) & (g4712) & (g2144) & (g5679)) + ((g830) & (!key[139]) & (!g1914) & (!g4712) & (!g2144) & (!g5679)) + ((g830) & (!key[139]) & (!g1914) & (!g4712) & (g2144) & (!g5679)) + ((g830) & (!key[139]) & (!g1914) & (g4712) & (!g2144) & (g5679)) + ((g830) & (!key[139]) & (!g1914) & (g4712) & (g2144) & (g5679)) + ((g830) & (!key[139]) & (g1914) & (!g4712) & (!g2144) & (!g5679)) + ((g830) & (!key[139]) & (g1914) & (!g4712) & (g2144) & (g5679)) + ((g830) & (!key[139]) & (g1914) & (g4712) & (!g2144) & (!g5679)) + ((g830) & (!key[139]) & (g1914) & (g4712) & (g2144) & (g5679)) + ((g830) & (key[139]) & (!g1914) & (!g4712) & (!g2144) & (!g5679)) + ((g830) & (key[139]) & (!g1914) & (!g4712) & (g2144) & (!g5679)) + ((g830) & (key[139]) & (!g1914) & (g4712) & (!g2144) & (g5679)) + ((g830) & (key[139]) & (!g1914) & (g4712) & (g2144) & (g5679)) + ((g830) & (key[139]) & (g1914) & (!g4712) & (!g2144) & (!g5679)) + ((g830) & (key[139]) & (g1914) & (!g4712) & (g2144) & (g5679)) + ((g830) & (key[139]) & (g1914) & (g4712) & (!g2144) & (!g5679)) + ((g830) & (key[139]) & (g1914) & (g4712) & (g2144) & (g5679)));
	assign g4714 = (((!g3240) & (!g3303) & (g3279) & (!g4616) & (g3307)) + ((!g3240) & (g3303) & (!g3279) & (!g4616) & (g3307)) + ((!g3240) & (g3303) & (!g3279) & (g4616) & (g3307)) + ((!g3240) & (g3303) & (g3279) & (!g4616) & (!g3307)) + ((!g3240) & (g3303) & (g3279) & (!g4616) & (g3307)) + ((!g3240) & (g3303) & (g3279) & (g4616) & (g3307)) + ((g3240) & (!g3303) & (!g3279) & (!g4616) & (g3307)) + ((g3240) & (!g3303) & (g3279) & (!g4616) & (g3307)) + ((g3240) & (!g3303) & (g3279) & (g4616) & (g3307)) + ((g3240) & (g3303) & (!g3279) & (!g4616) & (!g3307)) + ((g3240) & (g3303) & (!g3279) & (!g4616) & (g3307)) + ((g3240) & (g3303) & (!g3279) & (g4616) & (g3307)) + ((g3240) & (g3303) & (g3279) & (!g4616) & (!g3307)) + ((g3240) & (g3303) & (g3279) & (!g4616) & (g3307)) + ((g3240) & (g3303) & (g3279) & (g4616) & (!g3307)) + ((g3240) & (g3303) & (g3279) & (g4616) & (g3307)));
	assign g4715 = (((!g1983) & (g931) & (g3444)) + ((g1983) & (!g931) & (g3444)) + ((g1983) & (g931) & (!g3444)) + ((g1983) & (g931) & (g3444)));
	assign g4716 = (((!g830) & (key[107]) & (!g1914) & (!g4714) & (!g1985) & (!g5680)) + ((!g830) & (key[107]) & (!g1914) & (!g4714) & (!g1985) & (g5680)) + ((!g830) & (key[107]) & (!g1914) & (!g4714) & (g1985) & (!g5680)) + ((!g830) & (key[107]) & (!g1914) & (!g4714) & (g1985) & (g5680)) + ((!g830) & (key[107]) & (!g1914) & (g4714) & (!g1985) & (!g5680)) + ((!g830) & (key[107]) & (!g1914) & (g4714) & (!g1985) & (g5680)) + ((!g830) & (key[107]) & (!g1914) & (g4714) & (g1985) & (!g5680)) + ((!g830) & (key[107]) & (!g1914) & (g4714) & (g1985) & (g5680)) + ((!g830) & (key[107]) & (g1914) & (!g4714) & (!g1985) & (!g5680)) + ((!g830) & (key[107]) & (g1914) & (!g4714) & (!g1985) & (g5680)) + ((!g830) & (key[107]) & (g1914) & (!g4714) & (g1985) & (!g5680)) + ((!g830) & (key[107]) & (g1914) & (!g4714) & (g1985) & (g5680)) + ((!g830) & (key[107]) & (g1914) & (g4714) & (!g1985) & (!g5680)) + ((!g830) & (key[107]) & (g1914) & (g4714) & (!g1985) & (g5680)) + ((!g830) & (key[107]) & (g1914) & (g4714) & (g1985) & (!g5680)) + ((!g830) & (key[107]) & (g1914) & (g4714) & (g1985) & (g5680)) + ((g830) & (!key[107]) & (!g1914) & (!g4714) & (!g1985) & (!g5680)) + ((g830) & (!key[107]) & (!g1914) & (!g4714) & (g1985) & (g5680)) + ((g830) & (!key[107]) & (!g1914) & (g4714) & (!g1985) & (!g5680)) + ((g830) & (!key[107]) & (!g1914) & (g4714) & (g1985) & (g5680)) + ((g830) & (!key[107]) & (g1914) & (!g4714) & (!g1985) & (!g5680)) + ((g830) & (!key[107]) & (g1914) & (!g4714) & (g1985) & (!g5680)) + ((g830) & (!key[107]) & (g1914) & (g4714) & (!g1985) & (g5680)) + ((g830) & (!key[107]) & (g1914) & (g4714) & (g1985) & (g5680)) + ((g830) & (key[107]) & (!g1914) & (!g4714) & (!g1985) & (!g5680)) + ((g830) & (key[107]) & (!g1914) & (!g4714) & (g1985) & (g5680)) + ((g830) & (key[107]) & (!g1914) & (g4714) & (!g1985) & (!g5680)) + ((g830) & (key[107]) & (!g1914) & (g4714) & (g1985) & (g5680)) + ((g830) & (key[107]) & (g1914) & (!g4714) & (!g1985) & (!g5680)) + ((g830) & (key[107]) & (g1914) & (!g4714) & (g1985) & (!g5680)) + ((g830) & (key[107]) & (g1914) & (g4714) & (!g1985) & (g5680)) + ((g830) & (key[107]) & (g1914) & (g4714) & (g1985) & (g5680)));
	assign g4717 = (((!g2114) & (g3555) & (g2118)) + ((g2114) & (!g3555) & (g2118)) + ((g2114) & (g3555) & (!g2118)) + ((g2114) & (g3555) & (g2118)));
	assign g4718 = (((!g2647) & (!g2678) & (g3245) & (g3310) & (!g4621)) + ((!g2647) & (g2678) & (!g3245) & (g3310) & (!g4621)) + ((!g2647) & (g2678) & (!g3245) & (g3310) & (g4621)) + ((!g2647) & (g2678) & (g3245) & (!g3310) & (!g4621)) + ((!g2647) & (g2678) & (g3245) & (g3310) & (!g4621)) + ((!g2647) & (g2678) & (g3245) & (g3310) & (g4621)) + ((g2647) & (!g2678) & (!g3245) & (g3310) & (!g4621)) + ((g2647) & (!g2678) & (g3245) & (g3310) & (!g4621)) + ((g2647) & (!g2678) & (g3245) & (g3310) & (g4621)) + ((g2647) & (g2678) & (!g3245) & (!g3310) & (!g4621)) + ((g2647) & (g2678) & (!g3245) & (g3310) & (!g4621)) + ((g2647) & (g2678) & (!g3245) & (g3310) & (g4621)) + ((g2647) & (g2678) & (g3245) & (!g3310) & (!g4621)) + ((g2647) & (g2678) & (g3245) & (!g3310) & (g4621)) + ((g2647) & (g2678) & (g3245) & (g3310) & (!g4621)) + ((g2647) & (g2678) & (g3245) & (g3310) & (g4621)));
	assign g4719 = (((!g830) & (nonce[11]) & (!g1914) & (!g4718) & (!g2137) & (!g5681)) + ((!g830) & (nonce[11]) & (!g1914) & (!g4718) & (!g2137) & (g5681)) + ((!g830) & (nonce[11]) & (!g1914) & (!g4718) & (g2137) & (!g5681)) + ((!g830) & (nonce[11]) & (!g1914) & (!g4718) & (g2137) & (g5681)) + ((!g830) & (nonce[11]) & (!g1914) & (g4718) & (!g2137) & (!g5681)) + ((!g830) & (nonce[11]) & (!g1914) & (g4718) & (!g2137) & (g5681)) + ((!g830) & (nonce[11]) & (!g1914) & (g4718) & (g2137) & (!g5681)) + ((!g830) & (nonce[11]) & (!g1914) & (g4718) & (g2137) & (g5681)) + ((!g830) & (nonce[11]) & (g1914) & (!g4718) & (!g2137) & (!g5681)) + ((!g830) & (nonce[11]) & (g1914) & (!g4718) & (!g2137) & (g5681)) + ((!g830) & (nonce[11]) & (g1914) & (!g4718) & (g2137) & (!g5681)) + ((!g830) & (nonce[11]) & (g1914) & (!g4718) & (g2137) & (g5681)) + ((!g830) & (nonce[11]) & (g1914) & (g4718) & (!g2137) & (!g5681)) + ((!g830) & (nonce[11]) & (g1914) & (g4718) & (!g2137) & (g5681)) + ((!g830) & (nonce[11]) & (g1914) & (g4718) & (g2137) & (!g5681)) + ((!g830) & (nonce[11]) & (g1914) & (g4718) & (g2137) & (g5681)) + ((g830) & (!nonce[11]) & (!g1914) & (!g4718) & (!g2137) & (!g5681)) + ((g830) & (!nonce[11]) & (!g1914) & (!g4718) & (g2137) & (!g5681)) + ((g830) & (!nonce[11]) & (!g1914) & (g4718) & (!g2137) & (g5681)) + ((g830) & (!nonce[11]) & (!g1914) & (g4718) & (g2137) & (g5681)) + ((g830) & (!nonce[11]) & (g1914) & (!g4718) & (!g2137) & (!g5681)) + ((g830) & (!nonce[11]) & (g1914) & (!g4718) & (g2137) & (g5681)) + ((g830) & (!nonce[11]) & (g1914) & (g4718) & (!g2137) & (!g5681)) + ((g830) & (!nonce[11]) & (g1914) & (g4718) & (g2137) & (g5681)) + ((g830) & (nonce[11]) & (!g1914) & (!g4718) & (!g2137) & (!g5681)) + ((g830) & (nonce[11]) & (!g1914) & (!g4718) & (g2137) & (!g5681)) + ((g830) & (nonce[11]) & (!g1914) & (g4718) & (!g2137) & (g5681)) + ((g830) & (nonce[11]) & (!g1914) & (g4718) & (g2137) & (g5681)) + ((g830) & (nonce[11]) & (g1914) & (!g4718) & (!g2137) & (!g5681)) + ((g830) & (nonce[11]) & (g1914) & (!g4718) & (g2137) & (g5681)) + ((g830) & (nonce[11]) & (g1914) & (g4718) & (!g2137) & (!g5681)) + ((g830) & (nonce[11]) & (g1914) & (g4718) & (g2137) & (g5681)));
	assign g4720 = (((!g3074) & (!g3122) & (!g3095) & (g3131) & (!g4674)) + ((!g3074) & (!g3122) & (!g3095) & (g3131) & (g4674)) + ((!g3074) & (!g3122) & (g3095) & (!g3131) & (g4674)) + ((!g3074) & (!g3122) & (g3095) & (g3131) & (!g4674)) + ((!g3074) & (g3122) & (!g3095) & (!g3131) & (!g4674)) + ((!g3074) & (g3122) & (!g3095) & (!g3131) & (g4674)) + ((!g3074) & (g3122) & (g3095) & (!g3131) & (!g4674)) + ((!g3074) & (g3122) & (g3095) & (g3131) & (g4674)) + ((g3074) & (!g3122) & (!g3095) & (!g3131) & (g4674)) + ((g3074) & (!g3122) & (!g3095) & (g3131) & (!g4674)) + ((g3074) & (!g3122) & (g3095) & (!g3131) & (!g4674)) + ((g3074) & (!g3122) & (g3095) & (!g3131) & (g4674)) + ((g3074) & (g3122) & (!g3095) & (!g3131) & (!g4674)) + ((g3074) & (g3122) & (!g3095) & (g3131) & (g4674)) + ((g3074) & (g3122) & (g3095) & (g3131) & (!g4674)) + ((g3074) & (g3122) & (g3095) & (g3131) & (g4674)));
	assign g4721 = (((!g3084) & (!g3106) & (!g3090) & (g3139) & (!g4675)) + ((!g3084) & (!g3106) & (!g3090) & (g3139) & (g4675)) + ((!g3084) & (!g3106) & (g3090) & (!g3139) & (g4675)) + ((!g3084) & (!g3106) & (g3090) & (g3139) & (!g4675)) + ((!g3084) & (g3106) & (!g3090) & (!g3139) & (!g4675)) + ((!g3084) & (g3106) & (!g3090) & (!g3139) & (g4675)) + ((!g3084) & (g3106) & (g3090) & (!g3139) & (!g4675)) + ((!g3084) & (g3106) & (g3090) & (g3139) & (g4675)) + ((g3084) & (!g3106) & (!g3090) & (!g3139) & (g4675)) + ((g3084) & (!g3106) & (!g3090) & (g3139) & (!g4675)) + ((g3084) & (!g3106) & (g3090) & (!g3139) & (!g4675)) + ((g3084) & (!g3106) & (g3090) & (!g3139) & (g4675)) + ((g3084) & (g3106) & (!g3090) & (!g3139) & (!g4675)) + ((g3084) & (g3106) & (!g3090) & (g3139) & (g4675)) + ((g3084) & (g3106) & (g3090) & (g3139) & (!g4675)) + ((g3084) & (g3106) & (g3090) & (g3139) & (g4675)));
	assign g4722 = (((g830) & (!g1914) & (!g2480) & (!g4720) & (g4721)) + ((g830) & (!g1914) & (!g2480) & (g4720) & (g4721)) + ((g830) & (!g1914) & (g2480) & (!g4720) & (!g4721)) + ((g830) & (!g1914) & (g2480) & (g4720) & (!g4721)) + ((g830) & (g1914) & (!g2480) & (g4720) & (!g4721)) + ((g830) & (g1914) & (!g2480) & (g4720) & (g4721)) + ((g830) & (g1914) & (g2480) & (!g4720) & (!g4721)) + ((g830) & (g1914) & (g2480) & (!g4720) & (g4721)));
	assign g4723 = (((!g1894) & (g2034) & (!g1902) & (g2036)) + ((!g1894) & (g2034) & (g1902) & (g2036)) + ((g1894) & (!g2034) & (g1902) & (g2036)) + ((g1894) & (g2034) & (!g1902) & (g2036)) + ((g1894) & (g2034) & (g1902) & (!g2036)) + ((g1894) & (g2034) & (g1902) & (g2036)));
	assign g4724 = (((g1914) & (!g2065) & (!g2077) & (g4723)) + ((g1914) & (!g2065) & (g2077) & (!g4723)) + ((g1914) & (g2065) & (!g2077) & (!g4723)) + ((g1914) & (g2065) & (g2077) & (g4723)));
	assign g4725 = (((!g1906) & (g1940) & (!g1912) & (g2045)) + ((!g1906) & (g1940) & (g1912) & (g2045)) + ((g1906) & (!g1940) & (g1912) & (g2045)) + ((g1906) & (g1940) & (!g1912) & (g2045)) + ((g1906) & (g1940) & (g1912) & (!g2045)) + ((g1906) & (g1940) & (g1912) & (g2045)));
	assign g4726 = (((!g1914) & (!g1942) & (!g2091) & (g4725)) + ((!g1914) & (!g1942) & (g2091) & (!g4725)) + ((!g1914) & (g1942) & (!g2091) & (!g4725)) + ((!g1914) & (g1942) & (g2091) & (g4725)));
	assign g4727 = (((!g830) & (!g2486) & (!g4724) & (!g4726) & (nonce[43])) + ((!g830) & (!g2486) & (!g4724) & (g4726) & (nonce[43])) + ((!g830) & (!g2486) & (g4724) & (!g4726) & (nonce[43])) + ((!g830) & (!g2486) & (g4724) & (g4726) & (nonce[43])) + ((!g830) & (g2486) & (!g4724) & (!g4726) & (nonce[43])) + ((!g830) & (g2486) & (!g4724) & (g4726) & (nonce[43])) + ((!g830) & (g2486) & (g4724) & (!g4726) & (nonce[43])) + ((!g830) & (g2486) & (g4724) & (g4726) & (nonce[43])) + ((g830) & (!g2486) & (!g4724) & (g4726) & (!nonce[43])) + ((g830) & (!g2486) & (!g4724) & (g4726) & (nonce[43])) + ((g830) & (!g2486) & (g4724) & (!g4726) & (!nonce[43])) + ((g830) & (!g2486) & (g4724) & (!g4726) & (nonce[43])) + ((g830) & (!g2486) & (g4724) & (g4726) & (!nonce[43])) + ((g830) & (!g2486) & (g4724) & (g4726) & (nonce[43])) + ((g830) & (g2486) & (!g4724) & (!g4726) & (!nonce[43])) + ((g830) & (g2486) & (!g4724) & (!g4726) & (nonce[43])));
	assign g4728 = (((!g2650) & (!g2684) & (g3265) & (!g4628) & (g3312)) + ((!g2650) & (g2684) & (!g3265) & (!g4628) & (g3312)) + ((!g2650) & (g2684) & (!g3265) & (g4628) & (g3312)) + ((!g2650) & (g2684) & (g3265) & (!g4628) & (!g3312)) + ((!g2650) & (g2684) & (g3265) & (!g4628) & (g3312)) + ((!g2650) & (g2684) & (g3265) & (g4628) & (g3312)) + ((g2650) & (!g2684) & (!g3265) & (!g4628) & (g3312)) + ((g2650) & (!g2684) & (g3265) & (!g4628) & (g3312)) + ((g2650) & (!g2684) & (g3265) & (g4628) & (g3312)) + ((g2650) & (g2684) & (!g3265) & (!g4628) & (!g3312)) + ((g2650) & (g2684) & (!g3265) & (!g4628) & (g3312)) + ((g2650) & (g2684) & (!g3265) & (g4628) & (g3312)) + ((g2650) & (g2684) & (g3265) & (!g4628) & (!g3312)) + ((g2650) & (g2684) & (g3265) & (!g4628) & (g3312)) + ((g2650) & (g2684) & (g3265) & (g4628) & (!g3312)) + ((g2650) & (g2684) & (g3265) & (g4628) & (g3312)));
	assign g4729 = (((!g2108) & (g2116) & (g3602)) + ((g2108) & (!g2116) & (g3602)) + ((g2108) & (g2116) & (!g3602)) + ((g2108) & (g2116) & (g3602)));
	assign g4730 = (((!g830) & (key[235]) & (!g1914) & (!g4728) & (!g2144) & (!g5683)) + ((!g830) & (key[235]) & (!g1914) & (!g4728) & (!g2144) & (g5683)) + ((!g830) & (key[235]) & (!g1914) & (!g4728) & (g2144) & (!g5683)) + ((!g830) & (key[235]) & (!g1914) & (!g4728) & (g2144) & (g5683)) + ((!g830) & (key[235]) & (!g1914) & (g4728) & (!g2144) & (!g5683)) + ((!g830) & (key[235]) & (!g1914) & (g4728) & (!g2144) & (g5683)) + ((!g830) & (key[235]) & (!g1914) & (g4728) & (g2144) & (!g5683)) + ((!g830) & (key[235]) & (!g1914) & (g4728) & (g2144) & (g5683)) + ((!g830) & (key[235]) & (g1914) & (!g4728) & (!g2144) & (!g5683)) + ((!g830) & (key[235]) & (g1914) & (!g4728) & (!g2144) & (g5683)) + ((!g830) & (key[235]) & (g1914) & (!g4728) & (g2144) & (!g5683)) + ((!g830) & (key[235]) & (g1914) & (!g4728) & (g2144) & (g5683)) + ((!g830) & (key[235]) & (g1914) & (g4728) & (!g2144) & (!g5683)) + ((!g830) & (key[235]) & (g1914) & (g4728) & (!g2144) & (g5683)) + ((!g830) & (key[235]) & (g1914) & (g4728) & (g2144) & (!g5683)) + ((!g830) & (key[235]) & (g1914) & (g4728) & (g2144) & (g5683)) + ((g830) & (!key[235]) & (!g1914) & (!g4728) & (!g2144) & (!g5683)) + ((g830) & (!key[235]) & (!g1914) & (!g4728) & (g2144) & (g5683)) + ((g830) & (!key[235]) & (!g1914) & (g4728) & (!g2144) & (!g5683)) + ((g830) & (!key[235]) & (!g1914) & (g4728) & (g2144) & (g5683)) + ((g830) & (!key[235]) & (g1914) & (!g4728) & (!g2144) & (!g5683)) + ((g830) & (!key[235]) & (g1914) & (!g4728) & (g2144) & (!g5683)) + ((g830) & (!key[235]) & (g1914) & (g4728) & (!g2144) & (g5683)) + ((g830) & (!key[235]) & (g1914) & (g4728) & (g2144) & (g5683)) + ((g830) & (key[235]) & (!g1914) & (!g4728) & (!g2144) & (!g5683)) + ((g830) & (key[235]) & (!g1914) & (!g4728) & (g2144) & (g5683)) + ((g830) & (key[235]) & (!g1914) & (g4728) & (!g2144) & (!g5683)) + ((g830) & (key[235]) & (!g1914) & (g4728) & (g2144) & (g5683)) + ((g830) & (key[235]) & (g1914) & (!g4728) & (!g2144) & (!g5683)) + ((g830) & (key[235]) & (g1914) & (!g4728) & (g2144) & (!g5683)) + ((g830) & (key[235]) & (g1914) & (g4728) & (!g2144) & (g5683)) + ((g830) & (key[235]) & (g1914) & (g4728) & (g2144) & (g5683)));
	assign g4731 = (((!g1888) & (g1978) & (!g1912) & (g2045)) + ((!g1888) & (g1978) & (g1912) & (g2045)) + ((g1888) & (!g1978) & (g1912) & (g2045)) + ((g1888) & (g1978) & (!g1912) & (g2045)) + ((g1888) & (g1978) & (g1912) & (!g2045)) + ((g1888) & (g1978) & (g1912) & (g2045)));
	assign g4732 = (((g1914) & (!g1980) & (!g2091) & (g4731)) + ((g1914) & (!g1980) & (g2091) & (!g4731)) + ((g1914) & (g1980) & (!g2091) & (!g4731)) + ((g1914) & (g1980) & (g2091) & (g4731)));
	assign g4733 = (((!g1900) & (g2028) & (!g1902) & (g2036)) + ((!g1900) & (g2028) & (g1902) & (g2036)) + ((g1900) & (!g2028) & (g1902) & (g2036)) + ((g1900) & (g2028) & (!g1902) & (g2036)) + ((g1900) & (g2028) & (g1902) & (!g2036)) + ((g1900) & (g2028) & (g1902) & (g2036)));
	assign g4734 = (((!g1914) & (!g2074) & (!g2077) & (g4733)) + ((!g1914) & (!g2074) & (g2077) & (!g4733)) + ((!g1914) & (g2074) & (!g2077) & (!g4733)) + ((!g1914) & (g2074) & (g2077) & (g4733)));
	assign g4735 = (((!g830) & (!g2503) & (!g4732) & (!g4734) & (key[203])) + ((!g830) & (!g2503) & (!g4732) & (g4734) & (key[203])) + ((!g830) & (!g2503) & (g4732) & (!g4734) & (key[203])) + ((!g830) & (!g2503) & (g4732) & (g4734) & (key[203])) + ((!g830) & (g2503) & (!g4732) & (!g4734) & (key[203])) + ((!g830) & (g2503) & (!g4732) & (g4734) & (key[203])) + ((!g830) & (g2503) & (g4732) & (!g4734) & (key[203])) + ((!g830) & (g2503) & (g4732) & (g4734) & (key[203])) + ((g830) & (!g2503) & (!g4732) & (g4734) & (!key[203])) + ((g830) & (!g2503) & (!g4732) & (g4734) & (key[203])) + ((g830) & (!g2503) & (g4732) & (!g4734) & (!key[203])) + ((g830) & (!g2503) & (g4732) & (!g4734) & (key[203])) + ((g830) & (!g2503) & (g4732) & (g4734) & (!key[203])) + ((g830) & (!g2503) & (g4732) & (g4734) & (key[203])) + ((g830) & (g2503) & (!g4732) & (!g4734) & (!key[203])) + ((g830) & (g2503) & (!g4732) & (!g4734) & (key[203])));
	assign g4736 = (((!g3082) & (!g3136) & (!g3090) & (g3139) & (!g4686)) + ((!g3082) & (!g3136) & (!g3090) & (g3139) & (g4686)) + ((!g3082) & (!g3136) & (g3090) & (!g3139) & (g4686)) + ((!g3082) & (!g3136) & (g3090) & (g3139) & (!g4686)) + ((!g3082) & (g3136) & (!g3090) & (!g3139) & (!g4686)) + ((!g3082) & (g3136) & (!g3090) & (!g3139) & (g4686)) + ((!g3082) & (g3136) & (g3090) & (!g3139) & (!g4686)) + ((!g3082) & (g3136) & (g3090) & (g3139) & (g4686)) + ((g3082) & (!g3136) & (!g3090) & (!g3139) & (g4686)) + ((g3082) & (!g3136) & (!g3090) & (g3139) & (!g4686)) + ((g3082) & (!g3136) & (g3090) & (!g3139) & (!g4686)) + ((g3082) & (!g3136) & (g3090) & (!g3139) & (g4686)) + ((g3082) & (g3136) & (!g3090) & (!g3139) & (!g4686)) + ((g3082) & (g3136) & (!g3090) & (g3139) & (g4686)) + ((g3082) & (g3136) & (g3090) & (g3139) & (!g4686)) + ((g3082) & (g3136) & (g3090) & (g3139) & (g4686)));
	assign g4737 = (((!g3093) & (!g3119) & (!g3095) & (g3131) & (!g4687)) + ((!g3093) & (!g3119) & (!g3095) & (g3131) & (g4687)) + ((!g3093) & (!g3119) & (g3095) & (!g3131) & (g4687)) + ((!g3093) & (!g3119) & (g3095) & (g3131) & (!g4687)) + ((!g3093) & (g3119) & (!g3095) & (!g3131) & (!g4687)) + ((!g3093) & (g3119) & (!g3095) & (!g3131) & (g4687)) + ((!g3093) & (g3119) & (g3095) & (!g3131) & (!g4687)) + ((!g3093) & (g3119) & (g3095) & (g3131) & (g4687)) + ((g3093) & (!g3119) & (!g3095) & (!g3131) & (g4687)) + ((g3093) & (!g3119) & (!g3095) & (g3131) & (!g4687)) + ((g3093) & (!g3119) & (g3095) & (!g3131) & (!g4687)) + ((g3093) & (!g3119) & (g3095) & (!g3131) & (g4687)) + ((g3093) & (g3119) & (!g3095) & (!g3131) & (!g4687)) + ((g3093) & (g3119) & (!g3095) & (g3131) & (g4687)) + ((g3093) & (g3119) & (g3095) & (g3131) & (!g4687)) + ((g3093) & (g3119) & (g3095) & (g3131) & (g4687)));
	assign g4738 = (((g830) & (!g1914) & (!g2509) & (!g4736) & (g4737)) + ((g830) & (!g1914) & (!g2509) & (g4736) & (g4737)) + ((g830) & (!g1914) & (g2509) & (!g4736) & (!g4737)) + ((g830) & (!g1914) & (g2509) & (g4736) & (!g4737)) + ((g830) & (g1914) & (!g2509) & (g4736) & (!g4737)) + ((g830) & (g1914) & (!g2509) & (g4736) & (g4737)) + ((g830) & (g1914) & (g2509) & (!g4736) & (!g4737)) + ((g830) & (g1914) & (g2509) & (!g4736) & (g4737)));
	assign g4739 = (((!g3509) & (!g3510)));
	assign g4740 = (((g1914) & (!g1370) & (!g4739) & (!g2718)) + ((g1914) & (!g1370) & (g4739) & (g2718)) + ((g1914) & (g1370) & (!g4739) & (g2718)) + ((g1914) & (g1370) & (g4739) & (!g2718)));
	assign g4741 = (((!g3526) & (!g3527)));
	assign g4742 = (((!g1914) & (!g2703) & (!g2713) & (!g4741)) + ((!g1914) & (!g2703) & (g2713) & (g4741)) + ((!g1914) & (g2703) & (!g2713) & (g4741)) + ((!g1914) & (g2703) & (g2713) & (!g4741)));
	assign g4743 = (((!g830) & (!g2515) & (!g4740) & (!g4742) & (key[57])) + ((!g830) & (!g2515) & (!g4740) & (g4742) & (key[57])) + ((!g830) & (!g2515) & (g4740) & (!g4742) & (key[57])) + ((!g830) & (!g2515) & (g4740) & (g4742) & (key[57])) + ((!g830) & (g2515) & (!g4740) & (!g4742) & (key[57])) + ((!g830) & (g2515) & (!g4740) & (g4742) & (key[57])) + ((!g830) & (g2515) & (g4740) & (!g4742) & (key[57])) + ((!g830) & (g2515) & (g4740) & (g4742) & (key[57])) + ((g830) & (!g2515) & (!g4740) & (g4742) & (!key[57])) + ((g830) & (!g2515) & (!g4740) & (g4742) & (key[57])) + ((g830) & (!g2515) & (g4740) & (!g4742) & (!key[57])) + ((g830) & (!g2515) & (g4740) & (!g4742) & (key[57])) + ((g830) & (!g2515) & (g4740) & (g4742) & (!key[57])) + ((g830) & (!g2515) & (g4740) & (g4742) & (key[57])) + ((g830) & (g2515) & (!g4740) & (!g4742) & (!key[57])) + ((g830) & (g2515) & (!g4740) & (!g4742) & (key[57])));
	assign g4744 = (((!g1967) & (!g1969) & (!g2434) & (g2533) & (!g4692)) + ((!g1967) & (!g1969) & (!g2434) & (g2533) & (g4692)) + ((!g1967) & (!g1969) & (g2434) & (!g2533) & (!g4692)) + ((!g1967) & (!g1969) & (g2434) & (g2533) & (g4692)) + ((!g1967) & (g1969) & (!g2434) & (!g2533) & (!g4692)) + ((!g1967) & (g1969) & (!g2434) & (!g2533) & (g4692)) + ((!g1967) & (g1969) & (g2434) & (!g2533) & (g4692)) + ((!g1967) & (g1969) & (g2434) & (g2533) & (!g4692)) + ((g1967) & (!g1969) & (!g2434) & (!g2533) & (!g4692)) + ((g1967) & (!g1969) & (!g2434) & (g2533) & (g4692)) + ((g1967) & (!g1969) & (g2434) & (!g2533) & (!g4692)) + ((g1967) & (!g1969) & (g2434) & (!g2533) & (g4692)) + ((g1967) & (g1969) & (!g2434) & (!g2533) & (g4692)) + ((g1967) & (g1969) & (!g2434) & (g2533) & (!g4692)) + ((g1967) & (g1969) & (g2434) & (g2533) & (!g4692)) + ((g1967) & (g1969) & (g2434) & (g2533) & (g4692)));
	assign g4745 = (((!g2827) & (!g2833) & (!g3770)) + ((!g2827) & (g2833) & (g3770)) + ((g2827) & (!g2833) & (g3770)) + ((g2827) & (g2833) & (!g3770)));
	assign g4746 = (((!g830) & (!g1914) & (!g2516) & (!g4744) & (!g4745) & (key[89])) + ((!g830) & (!g1914) & (!g2516) & (!g4744) & (g4745) & (key[89])) + ((!g830) & (!g1914) & (!g2516) & (g4744) & (!g4745) & (key[89])) + ((!g830) & (!g1914) & (!g2516) & (g4744) & (g4745) & (key[89])) + ((!g830) & (!g1914) & (g2516) & (!g4744) & (!g4745) & (key[89])) + ((!g830) & (!g1914) & (g2516) & (!g4744) & (g4745) & (key[89])) + ((!g830) & (!g1914) & (g2516) & (g4744) & (!g4745) & (key[89])) + ((!g830) & (!g1914) & (g2516) & (g4744) & (g4745) & (key[89])) + ((!g830) & (g1914) & (!g2516) & (!g4744) & (!g4745) & (key[89])) + ((!g830) & (g1914) & (!g2516) & (!g4744) & (g4745) & (key[89])) + ((!g830) & (g1914) & (!g2516) & (g4744) & (!g4745) & (key[89])) + ((!g830) & (g1914) & (!g2516) & (g4744) & (g4745) & (key[89])) + ((!g830) & (g1914) & (g2516) & (!g4744) & (!g4745) & (key[89])) + ((!g830) & (g1914) & (g2516) & (!g4744) & (g4745) & (key[89])) + ((!g830) & (g1914) & (g2516) & (g4744) & (!g4745) & (key[89])) + ((!g830) & (g1914) & (g2516) & (g4744) & (g4745) & (key[89])) + ((g830) & (!g1914) & (!g2516) & (!g4744) & (g4745) & (!key[89])) + ((g830) & (!g1914) & (!g2516) & (!g4744) & (g4745) & (key[89])) + ((g830) & (!g1914) & (!g2516) & (g4744) & (g4745) & (!key[89])) + ((g830) & (!g1914) & (!g2516) & (g4744) & (g4745) & (key[89])) + ((g830) & (!g1914) & (g2516) & (!g4744) & (!g4745) & (!key[89])) + ((g830) & (!g1914) & (g2516) & (!g4744) & (!g4745) & (key[89])) + ((g830) & (!g1914) & (g2516) & (g4744) & (!g4745) & (!key[89])) + ((g830) & (!g1914) & (g2516) & (g4744) & (!g4745) & (key[89])) + ((g830) & (g1914) & (!g2516) & (g4744) & (!g4745) & (!key[89])) + ((g830) & (g1914) & (!g2516) & (g4744) & (!g4745) & (key[89])) + ((g830) & (g1914) & (!g2516) & (g4744) & (g4745) & (!key[89])) + ((g830) & (g1914) & (!g2516) & (g4744) & (g4745) & (key[89])) + ((g830) & (g1914) & (g2516) & (!g4744) & (!g4745) & (!key[89])) + ((g830) & (g1914) & (g2516) & (!g4744) & (!g4745) & (key[89])) + ((g830) & (g1914) & (g2516) & (!g4744) & (g4745) & (!key[89])) + ((g830) & (g1914) & (g2516) & (!g4744) & (g4745) & (key[89])));
	assign g4747 = (((!g3419) & (g3420)) + ((g3419) & (!g3420)) + ((g3419) & (g3420)));
	assign g4748 = (((!g3402) & (g3403)) + ((g3402) & (!g3403)) + ((g3402) & (g3403)));
	assign g8313 = (((!g5560) & (g5611) & (!g4749)) + ((!g5560) & (g5611) & (g4749)) + ((g5560) & (!g5611) & (g4749)) + ((g5560) & (g5611) & (g4749)));
	assign g4750 = (((!g830) & (!g2518) & (!g6531) & (g4749)) + ((!g830) & (!g2518) & (g6531) & (g4749)) + ((!g830) & (g2518) & (!g6531) & (g4749)) + ((!g830) & (g2518) & (g6531) & (g4749)) + ((g830) & (!g2518) & (g6531) & (!g4749)) + ((g830) & (!g2518) & (g6531) & (g4749)) + ((g830) & (g2518) & (!g6531) & (!g4749)) + ((g830) & (g2518) & (!g6531) & (g4749)));
	assign g4751 = (((!g3477) & (!g2810) & (!g2833)) + ((!g3477) & (g2810) & (g2833)) + ((g3477) & (!g2810) & (g2833)) + ((g3477) & (g2810) & (!g2833)));
	assign g4752 = (((!g2003) & (!g2005) & (!g2468) & (g2523) & (!g4698)) + ((!g2003) & (!g2005) & (!g2468) & (g2523) & (g4698)) + ((!g2003) & (!g2005) & (g2468) & (!g2523) & (!g4698)) + ((!g2003) & (!g2005) & (g2468) & (g2523) & (g4698)) + ((!g2003) & (g2005) & (!g2468) & (!g2523) & (!g4698)) + ((!g2003) & (g2005) & (!g2468) & (!g2523) & (g4698)) + ((!g2003) & (g2005) & (g2468) & (!g2523) & (g4698)) + ((!g2003) & (g2005) & (g2468) & (g2523) & (!g4698)) + ((g2003) & (!g2005) & (!g2468) & (!g2523) & (!g4698)) + ((g2003) & (!g2005) & (!g2468) & (g2523) & (g4698)) + ((g2003) & (!g2005) & (g2468) & (!g2523) & (!g4698)) + ((g2003) & (!g2005) & (g2468) & (!g2523) & (g4698)) + ((g2003) & (g2005) & (!g2468) & (!g2523) & (g4698)) + ((g2003) & (g2005) & (!g2468) & (g2523) & (!g4698)) + ((g2003) & (g2005) & (g2468) & (g2523) & (!g4698)) + ((g2003) & (g2005) & (g2468) & (g2523) & (g4698)));
	assign g4753 = (((!g830) & (!g1914) & (!g2519) & (!g4751) & (!g4752) & (key[185])) + ((!g830) & (!g1914) & (!g2519) & (!g4751) & (g4752) & (key[185])) + ((!g830) & (!g1914) & (!g2519) & (g4751) & (!g4752) & (key[185])) + ((!g830) & (!g1914) & (!g2519) & (g4751) & (g4752) & (key[185])) + ((!g830) & (!g1914) & (g2519) & (!g4751) & (!g4752) & (key[185])) + ((!g830) & (!g1914) & (g2519) & (!g4751) & (g4752) & (key[185])) + ((!g830) & (!g1914) & (g2519) & (g4751) & (!g4752) & (key[185])) + ((!g830) & (!g1914) & (g2519) & (g4751) & (g4752) & (key[185])) + ((!g830) & (g1914) & (!g2519) & (!g4751) & (!g4752) & (key[185])) + ((!g830) & (g1914) & (!g2519) & (!g4751) & (g4752) & (key[185])) + ((!g830) & (g1914) & (!g2519) & (g4751) & (!g4752) & (key[185])) + ((!g830) & (g1914) & (!g2519) & (g4751) & (g4752) & (key[185])) + ((!g830) & (g1914) & (g2519) & (!g4751) & (!g4752) & (key[185])) + ((!g830) & (g1914) & (g2519) & (!g4751) & (g4752) & (key[185])) + ((!g830) & (g1914) & (g2519) & (g4751) & (!g4752) & (key[185])) + ((!g830) & (g1914) & (g2519) & (g4751) & (g4752) & (key[185])) + ((g830) & (!g1914) & (!g2519) & (!g4751) & (g4752) & (!key[185])) + ((g830) & (!g1914) & (!g2519) & (!g4751) & (g4752) & (key[185])) + ((g830) & (!g1914) & (!g2519) & (g4751) & (g4752) & (!key[185])) + ((g830) & (!g1914) & (!g2519) & (g4751) & (g4752) & (key[185])) + ((g830) & (!g1914) & (g2519) & (!g4751) & (!g4752) & (!key[185])) + ((g830) & (!g1914) & (g2519) & (!g4751) & (!g4752) & (key[185])) + ((g830) & (!g1914) & (g2519) & (g4751) & (!g4752) & (!key[185])) + ((g830) & (!g1914) & (g2519) & (g4751) & (!g4752) & (key[185])) + ((g830) & (g1914) & (!g2519) & (g4751) & (!g4752) & (!key[185])) + ((g830) & (g1914) & (!g2519) & (g4751) & (!g4752) & (key[185])) + ((g830) & (g1914) & (!g2519) & (g4751) & (g4752) & (!key[185])) + ((g830) & (g1914) & (!g2519) & (g4751) & (g4752) & (key[185])) + ((g830) & (g1914) & (g2519) & (!g4751) & (!g4752) & (!key[185])) + ((g830) & (g1914) & (g2519) & (!g4751) & (!g4752) & (key[185])) + ((g830) & (g1914) & (g2519) & (!g4751) & (g4752) & (!key[185])) + ((g830) & (g1914) & (g2519) & (!g4751) & (g4752) & (key[185])));
	assign g4754 = (((!g2518) & (g3116)) + ((g2518) & (!g3116)));
	assign g4755 = (((!g2378) & (!g2426) & (g3041) & (g3086) & (g4605) & (g4754)) + ((!g2378) & (g2426) & (!g3041) & (g3086) & (!g4605) & (g4754)) + ((!g2378) & (g2426) & (!g3041) & (g3086) & (g4605) & (g4754)) + ((!g2378) & (g2426) & (g3041) & (!g3086) & (g4605) & (g4754)) + ((!g2378) & (g2426) & (g3041) & (g3086) & (!g4605) & (g4754)) + ((!g2378) & (g2426) & (g3041) & (g3086) & (g4605) & (g4754)) + ((g2378) & (!g2426) & (!g3041) & (g3086) & (g4605) & (g4754)) + ((g2378) & (!g2426) & (g3041) & (g3086) & (!g4605) & (g4754)) + ((g2378) & (!g2426) & (g3041) & (g3086) & (g4605) & (g4754)) + ((g2378) & (g2426) & (!g3041) & (!g3086) & (g4605) & (g4754)) + ((g2378) & (g2426) & (!g3041) & (g3086) & (!g4605) & (g4754)) + ((g2378) & (g2426) & (!g3041) & (g3086) & (g4605) & (g4754)) + ((g2378) & (g2426) & (g3041) & (!g3086) & (!g4605) & (g4754)) + ((g2378) & (g2426) & (g3041) & (!g3086) & (g4605) & (g4754)) + ((g2378) & (g2426) & (g3041) & (g3086) & (!g4605) & (g4754)) + ((g2378) & (g2426) & (g3041) & (g3086) & (g4605) & (g4754)));
	assign g4756 = (((g2518) & (g3116)));
	assign g4757 = (((!g2555) & (!g3161) & (!g4755) & (g4756)) + ((!g2555) & (!g3161) & (g4755) & (!g4756)) + ((!g2555) & (!g3161) & (g4755) & (g4756)) + ((!g2555) & (g3161) & (!g4755) & (!g4756)) + ((g2555) & (!g3161) & (!g4755) & (!g4756)) + ((g2555) & (g3161) & (!g4755) & (g4756)) + ((g2555) & (g3161) & (g4755) & (!g4756)) + ((g2555) & (g3161) & (g4755) & (g4756)));
	assign g4758 = (((!g2423) & (!g2515) & (g3080) & (g3125) & (g4659)) + ((!g2423) & (g2515) & (!g3080) & (g3125) & (!g4659)) + ((!g2423) & (g2515) & (!g3080) & (g3125) & (g4659)) + ((!g2423) & (g2515) & (g3080) & (!g3125) & (g4659)) + ((!g2423) & (g2515) & (g3080) & (g3125) & (!g4659)) + ((!g2423) & (g2515) & (g3080) & (g3125) & (g4659)) + ((g2423) & (!g2515) & (!g3080) & (g3125) & (g4659)) + ((g2423) & (!g2515) & (g3080) & (g3125) & (!g4659)) + ((g2423) & (!g2515) & (g3080) & (g3125) & (g4659)) + ((g2423) & (g2515) & (!g3080) & (!g3125) & (g4659)) + ((g2423) & (g2515) & (!g3080) & (g3125) & (!g4659)) + ((g2423) & (g2515) & (!g3080) & (g3125) & (g4659)) + ((g2423) & (g2515) & (g3080) & (!g3125) & (!g4659)) + ((g2423) & (g2515) & (g3080) & (!g3125) & (g4659)) + ((g2423) & (g2515) & (g3080) & (g3125) & (!g4659)) + ((g2423) & (g2515) & (g3080) & (g3125) & (g4659)));
	assign g8314 = (((!g5560) & (g5613) & (!g4759)) + ((!g5560) & (g5613) & (g4759)) + ((g5560) & (!g5613) & (g4759)) + ((g5560) & (g5613) & (g4759)));
	assign g4760 = (((!g3122) & (g3131)) + ((g3122) & (!g3131)));
	assign g4761 = (((!g3047) & (!g3074) & (g3056) & (g3095) & (g4624) & (g4760)) + ((!g3047) & (g3074) & (!g3056) & (g3095) & (!g4624) & (g4760)) + ((!g3047) & (g3074) & (!g3056) & (g3095) & (g4624) & (g4760)) + ((!g3047) & (g3074) & (g3056) & (!g3095) & (g4624) & (g4760)) + ((!g3047) & (g3074) & (g3056) & (g3095) & (!g4624) & (g4760)) + ((!g3047) & (g3074) & (g3056) & (g3095) & (g4624) & (g4760)) + ((g3047) & (!g3074) & (!g3056) & (g3095) & (g4624) & (g4760)) + ((g3047) & (!g3074) & (g3056) & (g3095) & (!g4624) & (g4760)) + ((g3047) & (!g3074) & (g3056) & (g3095) & (g4624) & (g4760)) + ((g3047) & (g3074) & (!g3056) & (!g3095) & (g4624) & (g4760)) + ((g3047) & (g3074) & (!g3056) & (g3095) & (!g4624) & (g4760)) + ((g3047) & (g3074) & (!g3056) & (g3095) & (g4624) & (g4760)) + ((g3047) & (g3074) & (g3056) & (!g3095) & (!g4624) & (g4760)) + ((g3047) & (g3074) & (g3056) & (!g3095) & (g4624) & (g4760)) + ((g3047) & (g3074) & (g3056) & (g3095) & (!g4624) & (g4760)) + ((g3047) & (g3074) & (g3056) & (g3095) & (g4624) & (g4760)));
	assign g4762 = (((g3122) & (g3131)));
	assign g4763 = (((!g3149) & (!g3170) & (!g4761) & (g4762)) + ((!g3149) & (!g3170) & (g4761) & (!g4762)) + ((!g3149) & (!g3170) & (g4761) & (g4762)) + ((!g3149) & (g3170) & (!g4761) & (!g4762)) + ((g3149) & (!g3170) & (!g4761) & (!g4762)) + ((g3149) & (g3170) & (!g4761) & (g4762)) + ((g3149) & (g3170) & (g4761) & (!g4762)) + ((g3149) & (g3170) & (g4761) & (g4762)));
	assign g4764 = (((!g3084) & (!g3106) & (g3090) & (g3139) & (g4675)) + ((!g3084) & (g3106) & (!g3090) & (g3139) & (!g4675)) + ((!g3084) & (g3106) & (!g3090) & (g3139) & (g4675)) + ((!g3084) & (g3106) & (g3090) & (!g3139) & (g4675)) + ((!g3084) & (g3106) & (g3090) & (g3139) & (!g4675)) + ((!g3084) & (g3106) & (g3090) & (g3139) & (g4675)) + ((g3084) & (!g3106) & (!g3090) & (g3139) & (g4675)) + ((g3084) & (!g3106) & (g3090) & (g3139) & (!g4675)) + ((g3084) & (!g3106) & (g3090) & (g3139) & (g4675)) + ((g3084) & (g3106) & (!g3090) & (!g3139) & (g4675)) + ((g3084) & (g3106) & (!g3090) & (g3139) & (!g4675)) + ((g3084) & (g3106) & (!g3090) & (g3139) & (g4675)) + ((g3084) & (g3106) & (g3090) & (!g3139) & (!g4675)) + ((g3084) & (g3106) & (g3090) & (!g3139) & (g4675)) + ((g3084) & (g3106) & (g3090) & (g3139) & (!g4675)) + ((g3084) & (g3106) & (g3090) & (g3139) & (g4675)));
	assign g4765 = (((!g1983) & (!g2127) & (g3710)) + ((!g1983) & (g2127) & (!g3710)) + ((g1983) & (!g2127) & (!g3710)) + ((g1983) & (g2127) & (g3710)));
	assign g4766 = (((!g2110) & (!g2118) & (g3727)) + ((!g2110) & (g2118) & (!g3727)) + ((g2110) & (!g2118) & (!g3727)) + ((g2110) & (g2118) & (g3727)));
	assign g4767 = (((!g830) & (!g1914) & (!g2539) & (!g4765) & (!g4766) & (key[204])) + ((!g830) & (!g1914) & (!g2539) & (!g4765) & (g4766) & (key[204])) + ((!g830) & (!g1914) & (!g2539) & (g4765) & (!g4766) & (key[204])) + ((!g830) & (!g1914) & (!g2539) & (g4765) & (g4766) & (key[204])) + ((!g830) & (!g1914) & (g2539) & (!g4765) & (!g4766) & (key[204])) + ((!g830) & (!g1914) & (g2539) & (!g4765) & (g4766) & (key[204])) + ((!g830) & (!g1914) & (g2539) & (g4765) & (!g4766) & (key[204])) + ((!g830) & (!g1914) & (g2539) & (g4765) & (g4766) & (key[204])) + ((!g830) & (g1914) & (!g2539) & (!g4765) & (!g4766) & (key[204])) + ((!g830) & (g1914) & (!g2539) & (!g4765) & (g4766) & (key[204])) + ((!g830) & (g1914) & (!g2539) & (g4765) & (!g4766) & (key[204])) + ((!g830) & (g1914) & (!g2539) & (g4765) & (g4766) & (key[204])) + ((!g830) & (g1914) & (g2539) & (!g4765) & (!g4766) & (key[204])) + ((!g830) & (g1914) & (g2539) & (!g4765) & (g4766) & (key[204])) + ((!g830) & (g1914) & (g2539) & (g4765) & (!g4766) & (key[204])) + ((!g830) & (g1914) & (g2539) & (g4765) & (g4766) & (key[204])) + ((g830) & (!g1914) & (!g2539) & (!g4765) & (g4766) & (!key[204])) + ((g830) & (!g1914) & (!g2539) & (!g4765) & (g4766) & (key[204])) + ((g830) & (!g1914) & (!g2539) & (g4765) & (g4766) & (!key[204])) + ((g830) & (!g1914) & (!g2539) & (g4765) & (g4766) & (key[204])) + ((g830) & (!g1914) & (g2539) & (!g4765) & (!g4766) & (!key[204])) + ((g830) & (!g1914) & (g2539) & (!g4765) & (!g4766) & (key[204])) + ((g830) & (!g1914) & (g2539) & (g4765) & (!g4766) & (!key[204])) + ((g830) & (!g1914) & (g2539) & (g4765) & (!g4766) & (key[204])) + ((g830) & (g1914) & (!g2539) & (g4765) & (!g4766) & (!key[204])) + ((g830) & (g1914) & (!g2539) & (g4765) & (!g4766) & (key[204])) + ((g830) & (g1914) & (!g2539) & (g4765) & (g4766) & (!key[204])) + ((g830) & (g1914) & (!g2539) & (g4765) & (g4766) & (key[204])) + ((g830) & (g1914) & (g2539) & (!g4765) & (!g4766) & (!key[204])) + ((g830) & (g1914) & (g2539) & (!g4765) & (!g4766) & (key[204])) + ((g830) & (g1914) & (g2539) & (!g4765) & (g4766) & (!key[204])) + ((g830) & (g1914) & (g2539) & (!g4765) & (g4766) & (key[204])));
	assign g4768 = (((!g2116) & (!g2118) & (g3811)) + ((!g2116) & (g2118) & (!g3811)) + ((g2116) & (!g2118) & (!g3811)) + ((g2116) & (g2118) & (g3811)));
	assign g4769 = (((!g1945) & (!g2127) & (g3828)) + ((!g1945) & (g2127) & (!g3828)) + ((g1945) & (!g2127) & (!g3828)) + ((g1945) & (g2127) & (g3828)));
	assign g4770 = (((!g830) & (!g1914) & (!g2544) & (!g4768) & (!g4769) & (nonce[44])) + ((!g830) & (!g1914) & (!g2544) & (!g4768) & (g4769) & (nonce[44])) + ((!g830) & (!g1914) & (!g2544) & (g4768) & (!g4769) & (nonce[44])) + ((!g830) & (!g1914) & (!g2544) & (g4768) & (g4769) & (nonce[44])) + ((!g830) & (!g1914) & (g2544) & (!g4768) & (!g4769) & (nonce[44])) + ((!g830) & (!g1914) & (g2544) & (!g4768) & (g4769) & (nonce[44])) + ((!g830) & (!g1914) & (g2544) & (g4768) & (!g4769) & (nonce[44])) + ((!g830) & (!g1914) & (g2544) & (g4768) & (g4769) & (nonce[44])) + ((!g830) & (g1914) & (!g2544) & (!g4768) & (!g4769) & (nonce[44])) + ((!g830) & (g1914) & (!g2544) & (!g4768) & (g4769) & (nonce[44])) + ((!g830) & (g1914) & (!g2544) & (g4768) & (!g4769) & (nonce[44])) + ((!g830) & (g1914) & (!g2544) & (g4768) & (g4769) & (nonce[44])) + ((!g830) & (g1914) & (g2544) & (!g4768) & (!g4769) & (nonce[44])) + ((!g830) & (g1914) & (g2544) & (!g4768) & (g4769) & (nonce[44])) + ((!g830) & (g1914) & (g2544) & (g4768) & (!g4769) & (nonce[44])) + ((!g830) & (g1914) & (g2544) & (g4768) & (g4769) & (nonce[44])) + ((g830) & (!g1914) & (!g2544) & (!g4768) & (g4769) & (!nonce[44])) + ((g830) & (!g1914) & (!g2544) & (!g4768) & (g4769) & (nonce[44])) + ((g830) & (!g1914) & (!g2544) & (g4768) & (g4769) & (!nonce[44])) + ((g830) & (!g1914) & (!g2544) & (g4768) & (g4769) & (nonce[44])) + ((g830) & (!g1914) & (g2544) & (!g4768) & (!g4769) & (!nonce[44])) + ((g830) & (!g1914) & (g2544) & (!g4768) & (!g4769) & (nonce[44])) + ((g830) & (!g1914) & (g2544) & (g4768) & (!g4769) & (!nonce[44])) + ((g830) & (!g1914) & (g2544) & (g4768) & (!g4769) & (nonce[44])) + ((g830) & (g1914) & (!g2544) & (g4768) & (!g4769) & (!nonce[44])) + ((g830) & (g1914) & (!g2544) & (g4768) & (!g4769) & (nonce[44])) + ((g830) & (g1914) & (!g2544) & (g4768) & (g4769) & (!nonce[44])) + ((g830) & (g1914) & (!g2544) & (g4768) & (g4769) & (nonce[44])) + ((g830) & (g1914) & (g2544) & (!g4768) & (!g4769) & (!nonce[44])) + ((g830) & (g1914) & (g2544) & (!g4768) & (!g4769) & (nonce[44])) + ((g830) & (g1914) & (g2544) & (!g4768) & (g4769) & (!nonce[44])) + ((g830) & (g1914) & (g2544) & (!g4768) & (g4769) & (nonce[44])));
	assign g4771 = (((!g3136) & (g3139)) + ((g3136) & (!g3139)));
	assign g4772 = (((!g3061) & (!g3082) & (g3064) & (g3090) & (g4634) & (g4771)) + ((!g3061) & (g3082) & (!g3064) & (g3090) & (!g4634) & (g4771)) + ((!g3061) & (g3082) & (!g3064) & (g3090) & (g4634) & (g4771)) + ((!g3061) & (g3082) & (g3064) & (!g3090) & (g4634) & (g4771)) + ((!g3061) & (g3082) & (g3064) & (g3090) & (!g4634) & (g4771)) + ((!g3061) & (g3082) & (g3064) & (g3090) & (g4634) & (g4771)) + ((g3061) & (!g3082) & (!g3064) & (g3090) & (g4634) & (g4771)) + ((g3061) & (!g3082) & (g3064) & (g3090) & (!g4634) & (g4771)) + ((g3061) & (!g3082) & (g3064) & (g3090) & (g4634) & (g4771)) + ((g3061) & (g3082) & (!g3064) & (!g3090) & (g4634) & (g4771)) + ((g3061) & (g3082) & (!g3064) & (g3090) & (!g4634) & (g4771)) + ((g3061) & (g3082) & (!g3064) & (g3090) & (g4634) & (g4771)) + ((g3061) & (g3082) & (g3064) & (!g3090) & (!g4634) & (g4771)) + ((g3061) & (g3082) & (g3064) & (!g3090) & (g4634) & (g4771)) + ((g3061) & (g3082) & (g3064) & (g3090) & (!g4634) & (g4771)) + ((g3061) & (g3082) & (g3064) & (g3090) & (g4634) & (g4771)));
	assign g4773 = (((g3136) & (g3139)));
	assign g4774 = (((!g3157) & (!g3165) & (!g4772) & (g4773)) + ((!g3157) & (!g3165) & (g4772) & (!g4773)) + ((!g3157) & (!g3165) & (g4772) & (g4773)) + ((!g3157) & (g3165) & (!g4772) & (!g4773)) + ((g3157) & (!g3165) & (!g4772) & (!g4773)) + ((g3157) & (g3165) & (!g4772) & (g4773)) + ((g3157) & (g3165) & (g4772) & (!g4773)) + ((g3157) & (g3165) & (g4772) & (g4773)));
	assign g4775 = (((!g3093) & (!g3119) & (g3095) & (g3131) & (g4687)) + ((!g3093) & (g3119) & (!g3095) & (g3131) & (!g4687)) + ((!g3093) & (g3119) & (!g3095) & (g3131) & (g4687)) + ((!g3093) & (g3119) & (g3095) & (!g3131) & (g4687)) + ((!g3093) & (g3119) & (g3095) & (g3131) & (!g4687)) + ((!g3093) & (g3119) & (g3095) & (g3131) & (g4687)) + ((g3093) & (!g3119) & (!g3095) & (g3131) & (g4687)) + ((g3093) & (!g3119) & (g3095) & (g3131) & (!g4687)) + ((g3093) & (!g3119) & (g3095) & (g3131) & (g4687)) + ((g3093) & (g3119) & (!g3095) & (!g3131) & (g4687)) + ((g3093) & (g3119) & (!g3095) & (g3131) & (!g4687)) + ((g3093) & (g3119) & (!g3095) & (g3131) & (g4687)) + ((g3093) & (g3119) & (g3095) & (!g3131) & (!g4687)) + ((g3093) & (g3119) & (g3095) & (!g3131) & (g4687)) + ((g3093) & (g3119) & (g3095) & (g3131) & (!g4687)) + ((g3093) & (g3119) & (g3095) & (g3131) & (g4687)));
	assign g4776 = (((!g1370) & (!g1406) & (!g4739) & (!g2718) & (g2764)) + ((!g1370) & (!g1406) & (!g4739) & (g2718) & (!g2764)) + ((!g1370) & (!g1406) & (g4739) & (!g2718) & (g2764)) + ((!g1370) & (!g1406) & (g4739) & (g2718) & (g2764)) + ((!g1370) & (g1406) & (!g4739) & (!g2718) & (!g2764)) + ((!g1370) & (g1406) & (!g4739) & (g2718) & (g2764)) + ((!g1370) & (g1406) & (g4739) & (!g2718) & (!g2764)) + ((!g1370) & (g1406) & (g4739) & (g2718) & (!g2764)) + ((g1370) & (!g1406) & (!g4739) & (!g2718) & (!g2764)) + ((g1370) & (!g1406) & (!g4739) & (g2718) & (!g2764)) + ((g1370) & (!g1406) & (g4739) & (!g2718) & (g2764)) + ((g1370) & (!g1406) & (g4739) & (g2718) & (!g2764)) + ((g1370) & (g1406) & (!g4739) & (!g2718) & (g2764)) + ((g1370) & (g1406) & (!g4739) & (g2718) & (g2764)) + ((g1370) & (g1406) & (g4739) & (!g2718) & (!g2764)) + ((g1370) & (g1406) & (g4739) & (g2718) & (g2764)));
	assign g4777 = (((!g2703) & (!g2768) & (!g2713) & (g2783) & (!g4741)) + ((!g2703) & (!g2768) & (!g2713) & (g2783) & (g4741)) + ((!g2703) & (!g2768) & (g2713) & (!g2783) & (!g4741)) + ((!g2703) & (!g2768) & (g2713) & (g2783) & (g4741)) + ((!g2703) & (g2768) & (!g2713) & (!g2783) & (!g4741)) + ((!g2703) & (g2768) & (!g2713) & (!g2783) & (g4741)) + ((!g2703) & (g2768) & (g2713) & (!g2783) & (g4741)) + ((!g2703) & (g2768) & (g2713) & (g2783) & (!g4741)) + ((g2703) & (!g2768) & (!g2713) & (!g2783) & (!g4741)) + ((g2703) & (!g2768) & (!g2713) & (g2783) & (g4741)) + ((g2703) & (!g2768) & (g2713) & (!g2783) & (!g4741)) + ((g2703) & (!g2768) & (g2713) & (!g2783) & (g4741)) + ((g2703) & (g2768) & (!g2713) & (!g2783) & (g4741)) + ((g2703) & (g2768) & (!g2713) & (g2783) & (!g4741)) + ((g2703) & (g2768) & (g2713) & (g2783) & (!g4741)) + ((g2703) & (g2768) & (g2713) & (g2783) & (g4741)));
	assign g4778 = (((!g830) & (!g1914) & (!g2551) & (!g4776) & (!g4777) & (key[58])) + ((!g830) & (!g1914) & (!g2551) & (!g4776) & (g4777) & (key[58])) + ((!g830) & (!g1914) & (!g2551) & (g4776) & (!g4777) & (key[58])) + ((!g830) & (!g1914) & (!g2551) & (g4776) & (g4777) & (key[58])) + ((!g830) & (!g1914) & (g2551) & (!g4776) & (!g4777) & (key[58])) + ((!g830) & (!g1914) & (g2551) & (!g4776) & (g4777) & (key[58])) + ((!g830) & (!g1914) & (g2551) & (g4776) & (!g4777) & (key[58])) + ((!g830) & (!g1914) & (g2551) & (g4776) & (g4777) & (key[58])) + ((!g830) & (g1914) & (!g2551) & (!g4776) & (!g4777) & (key[58])) + ((!g830) & (g1914) & (!g2551) & (!g4776) & (g4777) & (key[58])) + ((!g830) & (g1914) & (!g2551) & (g4776) & (!g4777) & (key[58])) + ((!g830) & (g1914) & (!g2551) & (g4776) & (g4777) & (key[58])) + ((!g830) & (g1914) & (g2551) & (!g4776) & (!g4777) & (key[58])) + ((!g830) & (g1914) & (g2551) & (!g4776) & (g4777) & (key[58])) + ((!g830) & (g1914) & (g2551) & (g4776) & (!g4777) & (key[58])) + ((!g830) & (g1914) & (g2551) & (g4776) & (g4777) & (key[58])) + ((g830) & (!g1914) & (!g2551) & (!g4776) & (g4777) & (!key[58])) + ((g830) & (!g1914) & (!g2551) & (!g4776) & (g4777) & (key[58])) + ((g830) & (!g1914) & (!g2551) & (g4776) & (g4777) & (!key[58])) + ((g830) & (!g1914) & (!g2551) & (g4776) & (g4777) & (key[58])) + ((g830) & (!g1914) & (g2551) & (!g4776) & (!g4777) & (!key[58])) + ((g830) & (!g1914) & (g2551) & (!g4776) & (!g4777) & (key[58])) + ((g830) & (!g1914) & (g2551) & (g4776) & (!g4777) & (!key[58])) + ((g830) & (!g1914) & (g2551) & (g4776) & (!g4777) & (key[58])) + ((g830) & (g1914) & (!g2551) & (g4776) & (!g4777) & (!key[58])) + ((g830) & (g1914) & (!g2551) & (g4776) & (!g4777) & (key[58])) + ((g830) & (g1914) & (!g2551) & (g4776) & (g4777) & (!key[58])) + ((g830) & (g1914) & (!g2551) & (g4776) & (g4777) & (key[58])) + ((g830) & (g1914) & (g2551) & (!g4776) & (!g4777) & (!key[58])) + ((g830) & (g1914) & (g2551) & (!g4776) & (!g4777) & (key[58])) + ((g830) & (g1914) & (g2551) & (!g4776) & (g4777) & (!key[58])) + ((g830) & (g1914) & (g2551) & (!g4776) & (g4777) & (key[58])));
	assign g4779 = (((!g2827) & (g2833) & (!g3770)) + ((g2827) & (!g2833) & (!g3770)) + ((g2827) & (g2833) & (!g3770)) + ((g2827) & (g2833) & (g3770)));
	assign g4780 = (((!g1972) & (!g2559) & (!g3753)) + ((!g1972) & (g2559) & (g3753)) + ((g1972) & (!g2559) & (g3753)) + ((g1972) & (g2559) & (!g3753)));
	assign g4781 = (((!g1914) & (!g2851) & (!g2874) & (g4779) & (!g4780)) + ((!g1914) & (!g2851) & (!g2874) & (g4779) & (g4780)) + ((!g1914) & (!g2851) & (g2874) & (!g4779) & (!g4780)) + ((!g1914) & (!g2851) & (g2874) & (!g4779) & (g4780)) + ((!g1914) & (g2851) & (!g2874) & (!g4779) & (!g4780)) + ((!g1914) & (g2851) & (!g2874) & (!g4779) & (g4780)) + ((!g1914) & (g2851) & (g2874) & (g4779) & (!g4780)) + ((!g1914) & (g2851) & (g2874) & (g4779) & (g4780)) + ((g1914) & (!g2851) & (!g2874) & (!g4779) & (g4780)) + ((g1914) & (!g2851) & (!g2874) & (g4779) & (g4780)) + ((g1914) & (!g2851) & (g2874) & (!g4779) & (g4780)) + ((g1914) & (!g2851) & (g2874) & (g4779) & (g4780)) + ((g1914) & (g2851) & (!g2874) & (!g4779) & (g4780)) + ((g1914) & (g2851) & (!g2874) & (g4779) & (g4780)) + ((g1914) & (g2851) & (g2874) & (!g4779) & (g4780)) + ((g1914) & (g2851) & (g2874) & (g4779) & (g4780)));
	assign g4782 = (((!g830) & (!g2552) & (!g4781) & (key[90])) + ((!g830) & (!g2552) & (g4781) & (key[90])) + ((!g830) & (g2552) & (!g4781) & (key[90])) + ((!g830) & (g2552) & (g4781) & (key[90])) + ((g830) & (!g2552) & (g4781) & (!key[90])) + ((g830) & (!g2552) & (g4781) & (key[90])) + ((g830) & (g2552) & (!g4781) & (!key[90])) + ((g830) & (g2552) & (!g4781) & (key[90])));
	assign g4783 = (((!g4748) & (!g2703) & (!g2742) & (!g2768) & (g2772)) + ((!g4748) & (!g2703) & (!g2742) & (g2768) & (!g2772)) + ((!g4748) & (!g2703) & (g2742) & (!g2768) & (g2772)) + ((!g4748) & (!g2703) & (g2742) & (g2768) & (!g2772)) + ((!g4748) & (g2703) & (!g2742) & (!g2768) & (g2772)) + ((!g4748) & (g2703) & (!g2742) & (g2768) & (!g2772)) + ((!g4748) & (g2703) & (g2742) & (!g2768) & (!g2772)) + ((!g4748) & (g2703) & (g2742) & (g2768) & (g2772)) + ((g4748) & (!g2703) & (!g2742) & (!g2768) & (g2772)) + ((g4748) & (!g2703) & (!g2742) & (g2768) & (!g2772)) + ((g4748) & (!g2703) & (g2742) & (!g2768) & (!g2772)) + ((g4748) & (!g2703) & (g2742) & (g2768) & (g2772)) + ((g4748) & (g2703) & (!g2742) & (!g2768) & (!g2772)) + ((g4748) & (g2703) & (!g2742) & (g2768) & (g2772)) + ((g4748) & (g2703) & (g2742) & (!g2768) & (!g2772)) + ((g4748) & (g2703) & (g2742) & (g2768) & (g2772)));
	assign g8315 = (((!g5560) & (g5614) & (!g4784)) + ((!g5560) & (g5614) & (g4784)) + ((g5560) & (!g5614) & (g4784)) + ((g5560) & (g5614) & (g4784)));
	assign g4785 = (((!g830) & (!g2555) & (!g6442) & (g4784)) + ((!g830) & (!g2555) & (g6442) & (g4784)) + ((!g830) & (g2555) & (!g6442) & (g4784)) + ((!g830) & (g2555) & (g6442) & (g4784)) + ((g830) & (!g2555) & (g6442) & (!g4784)) + ((g830) & (!g2555) & (g6442) & (g4784)) + ((g830) & (g2555) & (!g6442) & (!g4784)) + ((g830) & (g2555) & (!g6442) & (g4784)));
	assign g4786 = (((!g3477) & (!g2810) & (g2833)) + ((!g3477) & (g2810) & (!g2833)) + ((!g3477) & (g2810) & (g2833)) + ((g3477) & (g2810) & (g2833)));
	assign g4787 = (((!g2011) & (!g2575) & (!g3491)) + ((!g2011) & (g2575) & (g3491)) + ((g2011) & (!g2575) & (g3491)) + ((g2011) & (g2575) & (!g3491)));
	assign g4788 = (((!g1914) & (!g4786) & (!g2868) & (!g2874) & (g4787)) + ((!g1914) & (!g4786) & (!g2868) & (g2874) & (g4787)) + ((!g1914) & (!g4786) & (g2868) & (!g2874) & (g4787)) + ((!g1914) & (!g4786) & (g2868) & (g2874) & (g4787)) + ((!g1914) & (g4786) & (!g2868) & (!g2874) & (g4787)) + ((!g1914) & (g4786) & (!g2868) & (g2874) & (g4787)) + ((!g1914) & (g4786) & (g2868) & (!g2874) & (g4787)) + ((!g1914) & (g4786) & (g2868) & (g2874) & (g4787)) + ((g1914) & (!g4786) & (!g2868) & (g2874) & (!g4787)) + ((g1914) & (!g4786) & (!g2868) & (g2874) & (g4787)) + ((g1914) & (!g4786) & (g2868) & (!g2874) & (!g4787)) + ((g1914) & (!g4786) & (g2868) & (!g2874) & (g4787)) + ((g1914) & (g4786) & (!g2868) & (!g2874) & (!g4787)) + ((g1914) & (g4786) & (!g2868) & (!g2874) & (g4787)) + ((g1914) & (g4786) & (g2868) & (g2874) & (!g4787)) + ((g1914) & (g4786) & (g2868) & (g2874) & (g4787)));
	assign g4789 = (((!g830) & (!g2556) & (!g4788) & (key[186])) + ((!g830) & (!g2556) & (g4788) & (key[186])) + ((!g830) & (g2556) & (!g4788) & (key[186])) + ((!g830) & (g2556) & (g4788) & (key[186])) + ((g830) & (!g2556) & (g4788) & (!key[186])) + ((g830) & (!g2556) & (g4788) & (key[186])) + ((g830) & (g2556) & (!g4788) & (!key[186])) + ((g830) & (g2556) & (!g4788) & (key[186])));
	assign g4790 = (((!g3623) & (g3624)) + ((g3623) & (!g3624)) + ((g3623) & (g3624)));
	assign g4791 = (((!g1914) & (!g1954) & (!g1031) & (!g1900) & (g1904) & (!g4790)) + ((!g1914) & (!g1954) & (!g1031) & (!g1900) & (g1904) & (g4790)) + ((!g1914) & (!g1954) & (!g1031) & (g1900) & (!g1904) & (!g4790)) + ((!g1914) & (!g1954) & (!g1031) & (g1900) & (!g1904) & (g4790)) + ((!g1914) & (!g1954) & (g1031) & (!g1900) & (g1904) & (!g4790)) + ((!g1914) & (!g1954) & (g1031) & (!g1900) & (g1904) & (g4790)) + ((!g1914) & (!g1954) & (g1031) & (g1900) & (!g1904) & (!g4790)) + ((!g1914) & (!g1954) & (g1031) & (g1900) & (!g1904) & (g4790)) + ((!g1914) & (g1954) & (!g1031) & (!g1900) & (g1904) & (!g4790)) + ((!g1914) & (g1954) & (!g1031) & (!g1900) & (g1904) & (g4790)) + ((!g1914) & (g1954) & (!g1031) & (g1900) & (!g1904) & (!g4790)) + ((!g1914) & (g1954) & (!g1031) & (g1900) & (!g1904) & (g4790)) + ((!g1914) & (g1954) & (g1031) & (!g1900) & (g1904) & (!g4790)) + ((!g1914) & (g1954) & (g1031) & (!g1900) & (g1904) & (g4790)) + ((!g1914) & (g1954) & (g1031) & (g1900) & (!g1904) & (!g4790)) + ((!g1914) & (g1954) & (g1031) & (g1900) & (!g1904) & (g4790)) + ((g1914) & (!g1954) & (!g1031) & (!g1900) & (!g1904) & (g4790)) + ((g1914) & (!g1954) & (!g1031) & (!g1900) & (g1904) & (g4790)) + ((g1914) & (!g1954) & (!g1031) & (g1900) & (!g1904) & (g4790)) + ((g1914) & (!g1954) & (!g1031) & (g1900) & (g1904) & (g4790)) + ((g1914) & (!g1954) & (g1031) & (!g1900) & (!g1904) & (!g4790)) + ((g1914) & (!g1954) & (g1031) & (!g1900) & (g1904) & (!g4790)) + ((g1914) & (!g1954) & (g1031) & (g1900) & (!g1904) & (!g4790)) + ((g1914) & (!g1954) & (g1031) & (g1900) & (g1904) & (!g4790)) + ((g1914) & (g1954) & (!g1031) & (!g1900) & (!g1904) & (!g4790)) + ((g1914) & (g1954) & (!g1031) & (!g1900) & (g1904) & (!g4790)) + ((g1914) & (g1954) & (!g1031) & (g1900) & (!g1904) & (!g4790)) + ((g1914) & (g1954) & (!g1031) & (g1900) & (g1904) & (!g4790)) + ((g1914) & (g1954) & (g1031) & (!g1900) & (!g1904) & (g4790)) + ((g1914) & (g1954) & (g1031) & (!g1900) & (g1904) & (g4790)) + ((g1914) & (g1954) & (g1031) & (g1900) & (!g1904) & (g4790)) + ((g1914) & (g1954) & (g1031) & (g1900) & (g1904) & (g4790)));
	assign g4792 = (((!g830) & (!g2559) & (!g4791) & (key[13])) + ((!g830) & (!g2559) & (g4791) & (key[13])) + ((!g830) & (g2559) & (!g4791) & (key[13])) + ((!g830) & (g2559) & (g4791) & (key[13])) + ((g830) & (!g2559) & (g4791) & (!key[13])) + ((g830) & (!g2559) & (g4791) & (key[13])) + ((g830) & (g2559) & (!g4791) & (!key[13])) + ((g830) & (g2559) & (!g4791) & (key[13])));
	assign g4793 = (((!g2555) & (!g2601) & (!g3161) & (g3187) & (!g4755) & (!g4756)) + ((!g2555) & (!g2601) & (!g3161) & (g3187) & (!g4755) & (g4756)) + ((!g2555) & (!g2601) & (!g3161) & (g3187) & (g4755) & (!g4756)) + ((!g2555) & (!g2601) & (!g3161) & (g3187) & (g4755) & (g4756)) + ((!g2555) & (!g2601) & (g3161) & (!g3187) & (!g4755) & (g4756)) + ((!g2555) & (!g2601) & (g3161) & (!g3187) & (g4755) & (!g4756)) + ((!g2555) & (!g2601) & (g3161) & (!g3187) & (g4755) & (g4756)) + ((!g2555) & (!g2601) & (g3161) & (g3187) & (!g4755) & (!g4756)) + ((!g2555) & (g2601) & (!g3161) & (!g3187) & (!g4755) & (!g4756)) + ((!g2555) & (g2601) & (!g3161) & (!g3187) & (!g4755) & (g4756)) + ((!g2555) & (g2601) & (!g3161) & (!g3187) & (g4755) & (!g4756)) + ((!g2555) & (g2601) & (!g3161) & (!g3187) & (g4755) & (g4756)) + ((!g2555) & (g2601) & (g3161) & (!g3187) & (!g4755) & (!g4756)) + ((!g2555) & (g2601) & (g3161) & (g3187) & (!g4755) & (g4756)) + ((!g2555) & (g2601) & (g3161) & (g3187) & (g4755) & (!g4756)) + ((!g2555) & (g2601) & (g3161) & (g3187) & (g4755) & (g4756)) + ((g2555) & (!g2601) & (!g3161) & (!g3187) & (!g4755) & (g4756)) + ((g2555) & (!g2601) & (!g3161) & (!g3187) & (g4755) & (!g4756)) + ((g2555) & (!g2601) & (!g3161) & (!g3187) & (g4755) & (g4756)) + ((g2555) & (!g2601) & (!g3161) & (g3187) & (!g4755) & (!g4756)) + ((g2555) & (!g2601) & (g3161) & (!g3187) & (!g4755) & (!g4756)) + ((g2555) & (!g2601) & (g3161) & (!g3187) & (!g4755) & (g4756)) + ((g2555) & (!g2601) & (g3161) & (!g3187) & (g4755) & (!g4756)) + ((g2555) & (!g2601) & (g3161) & (!g3187) & (g4755) & (g4756)) + ((g2555) & (g2601) & (!g3161) & (!g3187) & (!g4755) & (!g4756)) + ((g2555) & (g2601) & (!g3161) & (g3187) & (!g4755) & (g4756)) + ((g2555) & (g2601) & (!g3161) & (g3187) & (g4755) & (!g4756)) + ((g2555) & (g2601) & (!g3161) & (g3187) & (g4755) & (g4756)) + ((g2555) & (g2601) & (g3161) & (g3187) & (!g4755) & (!g4756)) + ((g2555) & (g2601) & (g3161) & (g3187) & (!g4755) & (g4756)) + ((g2555) & (g2601) & (g3161) & (g3187) & (g4755) & (!g4756)) + ((g2555) & (g2601) & (g3161) & (g3187) & (g4755) & (g4756)));
	assign g4794 = (((!g2551) & (!g2598) & (!g3155) & (g3196) & (!g4758)) + ((!g2551) & (!g2598) & (!g3155) & (g3196) & (g4758)) + ((!g2551) & (!g2598) & (g3155) & (!g3196) & (g4758)) + ((!g2551) & (!g2598) & (g3155) & (g3196) & (!g4758)) + ((!g2551) & (g2598) & (!g3155) & (!g3196) & (!g4758)) + ((!g2551) & (g2598) & (!g3155) & (!g3196) & (g4758)) + ((!g2551) & (g2598) & (g3155) & (!g3196) & (!g4758)) + ((!g2551) & (g2598) & (g3155) & (g3196) & (g4758)) + ((g2551) & (!g2598) & (!g3155) & (!g3196) & (g4758)) + ((g2551) & (!g2598) & (!g3155) & (g3196) & (!g4758)) + ((g2551) & (!g2598) & (g3155) & (!g3196) & (!g4758)) + ((g2551) & (!g2598) & (g3155) & (!g3196) & (g4758)) + ((g2551) & (g2598) & (!g3155) & (!g3196) & (!g4758)) + ((g2551) & (g2598) & (!g3155) & (g3196) & (g4758)) + ((g2551) & (g2598) & (g3155) & (g3196) & (!g4758)) + ((g2551) & (g2598) & (g3155) & (g3196) & (g4758)));
	assign g4795 = (((!g830) & (!g1914) & (!g2566) & (!g4793) & (!g4794)) + ((!g830) & (!g1914) & (!g2566) & (!g4793) & (g4794)) + ((!g830) & (!g1914) & (!g2566) & (g4793) & (!g4794)) + ((!g830) & (!g1914) & (!g2566) & (g4793) & (g4794)) + ((!g830) & (!g1914) & (g2566) & (!g4793) & (!g4794)) + ((!g830) & (!g1914) & (g2566) & (!g4793) & (g4794)) + ((!g830) & (!g1914) & (g2566) & (g4793) & (!g4794)) + ((!g830) & (!g1914) & (g2566) & (g4793) & (g4794)) + ((!g830) & (g1914) & (!g2566) & (!g4793) & (!g4794)) + ((!g830) & (g1914) & (!g2566) & (!g4793) & (g4794)) + ((!g830) & (g1914) & (!g2566) & (g4793) & (!g4794)) + ((!g830) & (g1914) & (!g2566) & (g4793) & (g4794)) + ((!g830) & (g1914) & (g2566) & (!g4793) & (!g4794)) + ((!g830) & (g1914) & (g2566) & (!g4793) & (g4794)) + ((!g830) & (g1914) & (g2566) & (g4793) & (!g4794)) + ((!g830) & (g1914) & (g2566) & (g4793) & (g4794)) + ((g830) & (!g1914) & (!g2566) & (!g4793) & (g4794)) + ((g830) & (!g1914) & (!g2566) & (g4793) & (g4794)) + ((g830) & (!g1914) & (g2566) & (!g4793) & (!g4794)) + ((g830) & (!g1914) & (g2566) & (g4793) & (!g4794)) + ((g830) & (g1914) & (!g2566) & (g4793) & (!g4794)) + ((g830) & (g1914) & (!g2566) & (g4793) & (g4794)) + ((g830) & (g1914) & (g2566) & (!g4793) & (!g4794)) + ((g830) & (g1914) & (g2566) & (!g4793) & (g4794)));
	assign g4796 = (((!g3671) & (g3672)) + ((g3671) & (!g3672)) + ((g3671) & (g3672)));
	assign g4797 = (((!g1914) & (!g1884) & (!g1908) & (!g2233) & (!g2239) & (g4796)) + ((!g1914) & (!g1884) & (!g1908) & (!g2233) & (g2239) & (!g4796)) + ((!g1914) & (!g1884) & (!g1908) & (g2233) & (!g2239) & (!g4796)) + ((!g1914) & (!g1884) & (!g1908) & (g2233) & (g2239) & (g4796)) + ((!g1914) & (!g1884) & (g1908) & (!g2233) & (!g2239) & (g4796)) + ((!g1914) & (!g1884) & (g1908) & (!g2233) & (g2239) & (!g4796)) + ((!g1914) & (!g1884) & (g1908) & (g2233) & (!g2239) & (!g4796)) + ((!g1914) & (!g1884) & (g1908) & (g2233) & (g2239) & (g4796)) + ((!g1914) & (g1884) & (!g1908) & (!g2233) & (!g2239) & (g4796)) + ((!g1914) & (g1884) & (!g1908) & (!g2233) & (g2239) & (!g4796)) + ((!g1914) & (g1884) & (!g1908) & (g2233) & (!g2239) & (!g4796)) + ((!g1914) & (g1884) & (!g1908) & (g2233) & (g2239) & (g4796)) + ((!g1914) & (g1884) & (g1908) & (!g2233) & (!g2239) & (g4796)) + ((!g1914) & (g1884) & (g1908) & (!g2233) & (g2239) & (!g4796)) + ((!g1914) & (g1884) & (g1908) & (g2233) & (!g2239) & (!g4796)) + ((!g1914) & (g1884) & (g1908) & (g2233) & (g2239) & (g4796)) + ((g1914) & (!g1884) & (g1908) & (!g2233) & (!g2239) & (!g4796)) + ((g1914) & (!g1884) & (g1908) & (!g2233) & (!g2239) & (g4796)) + ((g1914) & (!g1884) & (g1908) & (!g2233) & (g2239) & (!g4796)) + ((g1914) & (!g1884) & (g1908) & (!g2233) & (g2239) & (g4796)) + ((g1914) & (!g1884) & (g1908) & (g2233) & (!g2239) & (!g4796)) + ((g1914) & (!g1884) & (g1908) & (g2233) & (!g2239) & (g4796)) + ((g1914) & (!g1884) & (g1908) & (g2233) & (g2239) & (!g4796)) + ((g1914) & (!g1884) & (g1908) & (g2233) & (g2239) & (g4796)) + ((g1914) & (g1884) & (!g1908) & (!g2233) & (!g2239) & (!g4796)) + ((g1914) & (g1884) & (!g1908) & (!g2233) & (!g2239) & (g4796)) + ((g1914) & (g1884) & (!g1908) & (!g2233) & (g2239) & (!g4796)) + ((g1914) & (g1884) & (!g1908) & (!g2233) & (g2239) & (g4796)) + ((g1914) & (g1884) & (!g1908) & (g2233) & (!g2239) & (!g4796)) + ((g1914) & (g1884) & (!g1908) & (g2233) & (!g2239) & (g4796)) + ((g1914) & (g1884) & (!g1908) & (g2233) & (g2239) & (!g4796)) + ((g1914) & (g1884) & (!g1908) & (g2233) & (g2239) & (g4796)));
	assign g8316 = (((!g5560) & (g5615) & (!g4798)) + ((!g5560) & (g5615) & (g4798)) + ((g5560) & (!g5615) & (g4798)) + ((g5560) & (g5615) & (g4798)));
	assign g4799 = (((!g830) & (!g2569) & (!g4797) & (g4798)) + ((!g830) & (!g2569) & (g4797) & (g4798)) + ((!g830) & (g2569) & (!g4797) & (g4798)) + ((!g830) & (g2569) & (g4797) & (g4798)) + ((g830) & (!g2569) & (g4797) & (!g4798)) + ((g830) & (!g2569) & (g4797) & (g4798)) + ((g830) & (g2569) & (!g4797) & (!g4798)) + ((g830) & (g2569) & (!g4797) & (g4798)));
	assign g4800 = (((!g3780) & (g3781)) + ((g3780) & (!g3781)) + ((g3780) & (g3781)));
	assign g4801 = (((!g1914) & (!g1906) & (!g2224) & (g1910) & (!g2236) & (!g4800)) + ((!g1914) & (!g1906) & (!g2224) & (g1910) & (!g2236) & (g4800)) + ((!g1914) & (!g1906) & (!g2224) & (g1910) & (g2236) & (!g4800)) + ((!g1914) & (!g1906) & (!g2224) & (g1910) & (g2236) & (g4800)) + ((!g1914) & (!g1906) & (g2224) & (g1910) & (!g2236) & (!g4800)) + ((!g1914) & (!g1906) & (g2224) & (g1910) & (!g2236) & (g4800)) + ((!g1914) & (!g1906) & (g2224) & (g1910) & (g2236) & (!g4800)) + ((!g1914) & (!g1906) & (g2224) & (g1910) & (g2236) & (g4800)) + ((!g1914) & (g1906) & (!g2224) & (!g1910) & (!g2236) & (!g4800)) + ((!g1914) & (g1906) & (!g2224) & (!g1910) & (!g2236) & (g4800)) + ((!g1914) & (g1906) & (!g2224) & (!g1910) & (g2236) & (!g4800)) + ((!g1914) & (g1906) & (!g2224) & (!g1910) & (g2236) & (g4800)) + ((!g1914) & (g1906) & (g2224) & (!g1910) & (!g2236) & (!g4800)) + ((!g1914) & (g1906) & (g2224) & (!g1910) & (!g2236) & (g4800)) + ((!g1914) & (g1906) & (g2224) & (!g1910) & (g2236) & (!g4800)) + ((!g1914) & (g1906) & (g2224) & (!g1910) & (g2236) & (g4800)) + ((g1914) & (!g1906) & (!g2224) & (!g1910) & (!g2236) & (g4800)) + ((g1914) & (!g1906) & (!g2224) & (!g1910) & (g2236) & (!g4800)) + ((g1914) & (!g1906) & (!g2224) & (g1910) & (!g2236) & (g4800)) + ((g1914) & (!g1906) & (!g2224) & (g1910) & (g2236) & (!g4800)) + ((g1914) & (!g1906) & (g2224) & (!g1910) & (!g2236) & (!g4800)) + ((g1914) & (!g1906) & (g2224) & (!g1910) & (g2236) & (g4800)) + ((g1914) & (!g1906) & (g2224) & (g1910) & (!g2236) & (!g4800)) + ((g1914) & (!g1906) & (g2224) & (g1910) & (g2236) & (g4800)) + ((g1914) & (g1906) & (!g2224) & (!g1910) & (!g2236) & (g4800)) + ((g1914) & (g1906) & (!g2224) & (!g1910) & (g2236) & (!g4800)) + ((g1914) & (g1906) & (!g2224) & (g1910) & (!g2236) & (g4800)) + ((g1914) & (g1906) & (!g2224) & (g1910) & (g2236) & (!g4800)) + ((g1914) & (g1906) & (g2224) & (!g1910) & (!g2236) & (!g4800)) + ((g1914) & (g1906) & (g2224) & (!g1910) & (g2236) & (g4800)) + ((g1914) & (g1906) & (g2224) & (g1910) & (!g2236) & (!g4800)) + ((g1914) & (g1906) & (g2224) & (g1910) & (g2236) & (g4800)));
	assign g4802 = (((!g830) & (!g2572) & (!g4801) & (key[141])) + ((!g830) & (!g2572) & (g4801) & (key[141])) + ((!g830) & (g2572) & (!g4801) & (key[141])) + ((!g830) & (g2572) & (g4801) & (key[141])) + ((g830) & (!g2572) & (g4801) & (!key[141])) + ((g830) & (!g2572) & (g4801) & (key[141])) + ((g830) & (g2572) & (!g4801) & (!key[141])) + ((g830) & (g2572) & (!g4801) & (key[141])));
	assign g4803 = (((!g3446) & (g3447)) + ((g3446) & (!g3447)) + ((g3446) & (g3447)));
	assign g4804 = (((!g1914) & (!g1992) & (!g1031) & (!g1894) & (!g1910) & (g4803)) + ((!g1914) & (!g1992) & (!g1031) & (!g1894) & (g1910) & (g4803)) + ((!g1914) & (!g1992) & (!g1031) & (g1894) & (!g1910) & (g4803)) + ((!g1914) & (!g1992) & (!g1031) & (g1894) & (g1910) & (g4803)) + ((!g1914) & (!g1992) & (g1031) & (!g1894) & (!g1910) & (!g4803)) + ((!g1914) & (!g1992) & (g1031) & (!g1894) & (g1910) & (!g4803)) + ((!g1914) & (!g1992) & (g1031) & (g1894) & (!g1910) & (!g4803)) + ((!g1914) & (!g1992) & (g1031) & (g1894) & (g1910) & (!g4803)) + ((!g1914) & (g1992) & (!g1031) & (!g1894) & (!g1910) & (!g4803)) + ((!g1914) & (g1992) & (!g1031) & (!g1894) & (g1910) & (!g4803)) + ((!g1914) & (g1992) & (!g1031) & (g1894) & (!g1910) & (!g4803)) + ((!g1914) & (g1992) & (!g1031) & (g1894) & (g1910) & (!g4803)) + ((!g1914) & (g1992) & (g1031) & (!g1894) & (!g1910) & (g4803)) + ((!g1914) & (g1992) & (g1031) & (!g1894) & (g1910) & (g4803)) + ((!g1914) & (g1992) & (g1031) & (g1894) & (!g1910) & (g4803)) + ((!g1914) & (g1992) & (g1031) & (g1894) & (g1910) & (g4803)) + ((g1914) & (!g1992) & (!g1031) & (!g1894) & (g1910) & (!g4803)) + ((g1914) & (!g1992) & (!g1031) & (!g1894) & (g1910) & (g4803)) + ((g1914) & (!g1992) & (!g1031) & (g1894) & (!g1910) & (!g4803)) + ((g1914) & (!g1992) & (!g1031) & (g1894) & (!g1910) & (g4803)) + ((g1914) & (!g1992) & (g1031) & (!g1894) & (g1910) & (!g4803)) + ((g1914) & (!g1992) & (g1031) & (!g1894) & (g1910) & (g4803)) + ((g1914) & (!g1992) & (g1031) & (g1894) & (!g1910) & (!g4803)) + ((g1914) & (!g1992) & (g1031) & (g1894) & (!g1910) & (g4803)) + ((g1914) & (g1992) & (!g1031) & (!g1894) & (g1910) & (!g4803)) + ((g1914) & (g1992) & (!g1031) & (!g1894) & (g1910) & (g4803)) + ((g1914) & (g1992) & (!g1031) & (g1894) & (!g1910) & (!g4803)) + ((g1914) & (g1992) & (!g1031) & (g1894) & (!g1910) & (g4803)) + ((g1914) & (g1992) & (g1031) & (!g1894) & (g1910) & (!g4803)) + ((g1914) & (g1992) & (g1031) & (!g1894) & (g1910) & (g4803)) + ((g1914) & (g1992) & (g1031) & (g1894) & (!g1910) & (!g4803)) + ((g1914) & (g1992) & (g1031) & (g1894) & (!g1910) & (g4803)));
	assign g4805 = (((!g830) & (!g2575) & (!g4804) & (key[109])) + ((!g830) & (!g2575) & (g4804) & (key[109])) + ((!g830) & (g2575) & (!g4804) & (key[109])) + ((!g830) & (g2575) & (g4804) & (key[109])) + ((g830) & (!g2575) & (g4804) & (!key[109])) + ((g830) & (!g2575) & (g4804) & (key[109])) + ((g830) & (g2575) & (!g4804) & (!key[109])) + ((g830) & (g2575) & (!g4804) & (key[109])));
	assign g4806 = (((!g3557) & (g3558)) + ((g3557) & (!g3558)) + ((g3557) & (g3558)));
	assign g4807 = (((!g1914) & (!g1890) & (!g2217) & (g1896) & (!g4806) & (!g2239)) + ((!g1914) & (!g1890) & (!g2217) & (g1896) & (!g4806) & (g2239)) + ((!g1914) & (!g1890) & (!g2217) & (g1896) & (g4806) & (!g2239)) + ((!g1914) & (!g1890) & (!g2217) & (g1896) & (g4806) & (g2239)) + ((!g1914) & (!g1890) & (g2217) & (g1896) & (!g4806) & (!g2239)) + ((!g1914) & (!g1890) & (g2217) & (g1896) & (!g4806) & (g2239)) + ((!g1914) & (!g1890) & (g2217) & (g1896) & (g4806) & (!g2239)) + ((!g1914) & (!g1890) & (g2217) & (g1896) & (g4806) & (g2239)) + ((!g1914) & (g1890) & (!g2217) & (!g1896) & (!g4806) & (!g2239)) + ((!g1914) & (g1890) & (!g2217) & (!g1896) & (!g4806) & (g2239)) + ((!g1914) & (g1890) & (!g2217) & (!g1896) & (g4806) & (!g2239)) + ((!g1914) & (g1890) & (!g2217) & (!g1896) & (g4806) & (g2239)) + ((!g1914) & (g1890) & (g2217) & (!g1896) & (!g4806) & (!g2239)) + ((!g1914) & (g1890) & (g2217) & (!g1896) & (!g4806) & (g2239)) + ((!g1914) & (g1890) & (g2217) & (!g1896) & (g4806) & (!g2239)) + ((!g1914) & (g1890) & (g2217) & (!g1896) & (g4806) & (g2239)) + ((g1914) & (!g1890) & (!g2217) & (!g1896) & (!g4806) & (g2239)) + ((g1914) & (!g1890) & (!g2217) & (!g1896) & (g4806) & (!g2239)) + ((g1914) & (!g1890) & (!g2217) & (g1896) & (!g4806) & (g2239)) + ((g1914) & (!g1890) & (!g2217) & (g1896) & (g4806) & (!g2239)) + ((g1914) & (!g1890) & (g2217) & (!g1896) & (!g4806) & (!g2239)) + ((g1914) & (!g1890) & (g2217) & (!g1896) & (g4806) & (g2239)) + ((g1914) & (!g1890) & (g2217) & (g1896) & (!g4806) & (!g2239)) + ((g1914) & (!g1890) & (g2217) & (g1896) & (g4806) & (g2239)) + ((g1914) & (g1890) & (!g2217) & (!g1896) & (!g4806) & (g2239)) + ((g1914) & (g1890) & (!g2217) & (!g1896) & (g4806) & (!g2239)) + ((g1914) & (g1890) & (!g2217) & (g1896) & (!g4806) & (g2239)) + ((g1914) & (g1890) & (!g2217) & (g1896) & (g4806) & (!g2239)) + ((g1914) & (g1890) & (g2217) & (!g1896) & (!g4806) & (!g2239)) + ((g1914) & (g1890) & (g2217) & (!g1896) & (g4806) & (g2239)) + ((g1914) & (g1890) & (g2217) & (g1896) & (!g4806) & (!g2239)) + ((g1914) & (g1890) & (g2217) & (g1896) & (g4806) & (g2239)));
	assign g4808 = (((!g830) & (!g2578) & (!g4807) & (nonce[13])) + ((!g830) & (!g2578) & (g4807) & (nonce[13])) + ((!g830) & (g2578) & (!g4807) & (nonce[13])) + ((!g830) & (g2578) & (g4807) & (nonce[13])) + ((g830) & (!g2578) & (g4807) & (!nonce[13])) + ((g830) & (!g2578) & (g4807) & (nonce[13])) + ((g830) & (g2578) & (!g4807) & (!nonce[13])) + ((g830) & (g2578) & (!g4807) & (nonce[13])));
	assign g4809 = (((!g3149) & (!g3193) & (!g3170) & (g3202) & (!g4761) & (!g4762)) + ((!g3149) & (!g3193) & (!g3170) & (g3202) & (!g4761) & (g4762)) + ((!g3149) & (!g3193) & (!g3170) & (g3202) & (g4761) & (!g4762)) + ((!g3149) & (!g3193) & (!g3170) & (g3202) & (g4761) & (g4762)) + ((!g3149) & (!g3193) & (g3170) & (!g3202) & (!g4761) & (g4762)) + ((!g3149) & (!g3193) & (g3170) & (!g3202) & (g4761) & (!g4762)) + ((!g3149) & (!g3193) & (g3170) & (!g3202) & (g4761) & (g4762)) + ((!g3149) & (!g3193) & (g3170) & (g3202) & (!g4761) & (!g4762)) + ((!g3149) & (g3193) & (!g3170) & (!g3202) & (!g4761) & (!g4762)) + ((!g3149) & (g3193) & (!g3170) & (!g3202) & (!g4761) & (g4762)) + ((!g3149) & (g3193) & (!g3170) & (!g3202) & (g4761) & (!g4762)) + ((!g3149) & (g3193) & (!g3170) & (!g3202) & (g4761) & (g4762)) + ((!g3149) & (g3193) & (g3170) & (!g3202) & (!g4761) & (!g4762)) + ((!g3149) & (g3193) & (g3170) & (g3202) & (!g4761) & (g4762)) + ((!g3149) & (g3193) & (g3170) & (g3202) & (g4761) & (!g4762)) + ((!g3149) & (g3193) & (g3170) & (g3202) & (g4761) & (g4762)) + ((g3149) & (!g3193) & (!g3170) & (!g3202) & (!g4761) & (g4762)) + ((g3149) & (!g3193) & (!g3170) & (!g3202) & (g4761) & (!g4762)) + ((g3149) & (!g3193) & (!g3170) & (!g3202) & (g4761) & (g4762)) + ((g3149) & (!g3193) & (!g3170) & (g3202) & (!g4761) & (!g4762)) + ((g3149) & (!g3193) & (g3170) & (!g3202) & (!g4761) & (!g4762)) + ((g3149) & (!g3193) & (g3170) & (!g3202) & (!g4761) & (g4762)) + ((g3149) & (!g3193) & (g3170) & (!g3202) & (g4761) & (!g4762)) + ((g3149) & (!g3193) & (g3170) & (!g3202) & (g4761) & (g4762)) + ((g3149) & (g3193) & (!g3170) & (!g3202) & (!g4761) & (!g4762)) + ((g3149) & (g3193) & (!g3170) & (g3202) & (!g4761) & (g4762)) + ((g3149) & (g3193) & (!g3170) & (g3202) & (g4761) & (!g4762)) + ((g3149) & (g3193) & (!g3170) & (g3202) & (g4761) & (g4762)) + ((g3149) & (g3193) & (g3170) & (g3202) & (!g4761) & (!g4762)) + ((g3149) & (g3193) & (g3170) & (g3202) & (!g4761) & (g4762)) + ((g3149) & (g3193) & (g3170) & (g3202) & (g4761) & (!g4762)) + ((g3149) & (g3193) & (g3170) & (g3202) & (g4761) & (g4762)));
	assign g4810 = (((!g3159) & (!g3177) & (!g3165) & (g3210) & (!g4764)) + ((!g3159) & (!g3177) & (!g3165) & (g3210) & (g4764)) + ((!g3159) & (!g3177) & (g3165) & (!g3210) & (g4764)) + ((!g3159) & (!g3177) & (g3165) & (g3210) & (!g4764)) + ((!g3159) & (g3177) & (!g3165) & (!g3210) & (!g4764)) + ((!g3159) & (g3177) & (!g3165) & (!g3210) & (g4764)) + ((!g3159) & (g3177) & (g3165) & (!g3210) & (!g4764)) + ((!g3159) & (g3177) & (g3165) & (g3210) & (g4764)) + ((g3159) & (!g3177) & (!g3165) & (!g3210) & (g4764)) + ((g3159) & (!g3177) & (!g3165) & (g3210) & (!g4764)) + ((g3159) & (!g3177) & (g3165) & (!g3210) & (!g4764)) + ((g3159) & (!g3177) & (g3165) & (!g3210) & (g4764)) + ((g3159) & (g3177) & (!g3165) & (!g3210) & (!g4764)) + ((g3159) & (g3177) & (!g3165) & (g3210) & (g4764)) + ((g3159) & (g3177) & (g3165) & (g3210) & (!g4764)) + ((g3159) & (g3177) & (g3165) & (g3210) & (g4764)));
	assign g4811 = (((!g830) & (!g1914) & (!g2581) & (!g4809) & (!g4810)) + ((!g830) & (!g1914) & (!g2581) & (!g4809) & (g4810)) + ((!g830) & (!g1914) & (!g2581) & (g4809) & (!g4810)) + ((!g830) & (!g1914) & (!g2581) & (g4809) & (g4810)) + ((!g830) & (!g1914) & (g2581) & (!g4809) & (!g4810)) + ((!g830) & (!g1914) & (g2581) & (!g4809) & (g4810)) + ((!g830) & (!g1914) & (g2581) & (g4809) & (!g4810)) + ((!g830) & (!g1914) & (g2581) & (g4809) & (g4810)) + ((!g830) & (g1914) & (!g2581) & (!g4809) & (!g4810)) + ((!g830) & (g1914) & (!g2581) & (!g4809) & (g4810)) + ((!g830) & (g1914) & (!g2581) & (g4809) & (!g4810)) + ((!g830) & (g1914) & (!g2581) & (g4809) & (g4810)) + ((!g830) & (g1914) & (g2581) & (!g4809) & (!g4810)) + ((!g830) & (g1914) & (g2581) & (!g4809) & (g4810)) + ((!g830) & (g1914) & (g2581) & (g4809) & (!g4810)) + ((!g830) & (g1914) & (g2581) & (g4809) & (g4810)) + ((g830) & (!g1914) & (!g2581) & (!g4809) & (g4810)) + ((g830) & (!g1914) & (!g2581) & (g4809) & (g4810)) + ((g830) & (!g1914) & (g2581) & (!g4809) & (!g4810)) + ((g830) & (!g1914) & (g2581) & (g4809) & (!g4810)) + ((g830) & (g1914) & (!g2581) & (g4809) & (!g4810)) + ((g830) & (g1914) & (!g2581) & (g4809) & (g4810)) + ((g830) & (g1914) & (g2581) & (!g4809) & (!g4810)) + ((g830) & (g1914) & (g2581) & (!g4809) & (g4810)));
	assign g4812 = (((!g2116) & (g2118) & (g3811)) + ((g2116) & (!g2118) & (g3811)) + ((g2116) & (g2118) & (!g3811)) + ((g2116) & (g2118) & (g3811)));
	assign g4813 = (((g1914) & (!g2147) & (!g2159) & (g4812)) + ((g1914) & (!g2147) & (g2159) & (!g4812)) + ((g1914) & (g2147) & (!g2159) & (!g4812)) + ((g1914) & (g2147) & (g2159) & (g4812)));
	assign g4814 = (((!g1945) & (g2127) & (g3828)) + ((g1945) & (!g2127) & (g3828)) + ((g1945) & (g2127) & (!g3828)) + ((g1945) & (g2127) & (g3828)));
	assign g4815 = (((!g1914) & (!g1947) & (!g2173) & (g4814)) + ((!g1914) & (!g1947) & (g2173) & (!g4814)) + ((!g1914) & (g1947) & (!g2173) & (!g4814)) + ((!g1914) & (g1947) & (g2173) & (g4814)));
	assign g4816 = (((!g830) & (!g2584) & (!g4813) & (!g4815) & (nonce[45])) + ((!g830) & (!g2584) & (!g4813) & (g4815) & (nonce[45])) + ((!g830) & (!g2584) & (g4813) & (!g4815) & (nonce[45])) + ((!g830) & (!g2584) & (g4813) & (g4815) & (nonce[45])) + ((!g830) & (g2584) & (!g4813) & (!g4815) & (nonce[45])) + ((!g830) & (g2584) & (!g4813) & (g4815) & (nonce[45])) + ((!g830) & (g2584) & (g4813) & (!g4815) & (nonce[45])) + ((!g830) & (g2584) & (g4813) & (g4815) & (nonce[45])) + ((g830) & (!g2584) & (!g4813) & (g4815) & (!nonce[45])) + ((g830) & (!g2584) & (!g4813) & (g4815) & (nonce[45])) + ((g830) & (!g2584) & (g4813) & (!g4815) & (!nonce[45])) + ((g830) & (!g2584) & (g4813) & (!g4815) & (nonce[45])) + ((g830) & (!g2584) & (g4813) & (g4815) & (!nonce[45])) + ((g830) & (!g2584) & (g4813) & (g4815) & (nonce[45])) + ((g830) & (g2584) & (!g4813) & (!g4815) & (!nonce[45])) + ((g830) & (g2584) & (!g4813) & (!g4815) & (nonce[45])));
	assign g4817 = (((!g3604) & (g3605)) + ((g3604) & (!g3605)) + ((g3604) & (g3605)));
	assign g4818 = (((!g1914) & (!g1888) & (!g2224) & (!g2227) & (!g1904) & (g4817)) + ((!g1914) & (!g1888) & (!g2224) & (!g2227) & (g1904) & (g4817)) + ((!g1914) & (!g1888) & (!g2224) & (g2227) & (!g1904) & (!g4817)) + ((!g1914) & (!g1888) & (!g2224) & (g2227) & (g1904) & (!g4817)) + ((!g1914) & (!g1888) & (g2224) & (!g2227) & (!g1904) & (!g4817)) + ((!g1914) & (!g1888) & (g2224) & (!g2227) & (g1904) & (!g4817)) + ((!g1914) & (!g1888) & (g2224) & (g2227) & (!g1904) & (g4817)) + ((!g1914) & (!g1888) & (g2224) & (g2227) & (g1904) & (g4817)) + ((!g1914) & (g1888) & (!g2224) & (!g2227) & (!g1904) & (g4817)) + ((!g1914) & (g1888) & (!g2224) & (!g2227) & (g1904) & (g4817)) + ((!g1914) & (g1888) & (!g2224) & (g2227) & (!g1904) & (!g4817)) + ((!g1914) & (g1888) & (!g2224) & (g2227) & (g1904) & (!g4817)) + ((!g1914) & (g1888) & (g2224) & (!g2227) & (!g1904) & (!g4817)) + ((!g1914) & (g1888) & (g2224) & (!g2227) & (g1904) & (!g4817)) + ((!g1914) & (g1888) & (g2224) & (g2227) & (!g1904) & (g4817)) + ((!g1914) & (g1888) & (g2224) & (g2227) & (g1904) & (g4817)) + ((g1914) & (!g1888) & (!g2224) & (!g2227) & (g1904) & (!g4817)) + ((g1914) & (!g1888) & (!g2224) & (!g2227) & (g1904) & (g4817)) + ((g1914) & (!g1888) & (!g2224) & (g2227) & (g1904) & (!g4817)) + ((g1914) & (!g1888) & (!g2224) & (g2227) & (g1904) & (g4817)) + ((g1914) & (!g1888) & (g2224) & (!g2227) & (g1904) & (!g4817)) + ((g1914) & (!g1888) & (g2224) & (!g2227) & (g1904) & (g4817)) + ((g1914) & (!g1888) & (g2224) & (g2227) & (g1904) & (!g4817)) + ((g1914) & (!g1888) & (g2224) & (g2227) & (g1904) & (g4817)) + ((g1914) & (g1888) & (!g2224) & (!g2227) & (!g1904) & (!g4817)) + ((g1914) & (g1888) & (!g2224) & (!g2227) & (!g1904) & (g4817)) + ((g1914) & (g1888) & (!g2224) & (g2227) & (!g1904) & (!g4817)) + ((g1914) & (g1888) & (!g2224) & (g2227) & (!g1904) & (g4817)) + ((g1914) & (g1888) & (g2224) & (!g2227) & (!g1904) & (!g4817)) + ((g1914) & (g1888) & (g2224) & (!g2227) & (!g1904) & (g4817)) + ((g1914) & (g1888) & (g2224) & (g2227) & (!g1904) & (!g4817)) + ((g1914) & (g1888) & (g2224) & (g2227) & (!g1904) & (g4817)));
	assign g4819 = (((!g830) & (!g2589) & (!g4818) & (key[237])) + ((!g830) & (!g2589) & (g4818) & (key[237])) + ((!g830) & (g2589) & (!g4818) & (key[237])) + ((!g830) & (g2589) & (g4818) & (key[237])) + ((g830) & (!g2589) & (g4818) & (!key[237])) + ((g830) & (!g2589) & (g4818) & (key[237])) + ((g830) & (g2589) & (!g4818) & (!key[237])) + ((g830) & (g2589) & (!g4818) & (key[237])));
	assign g4820 = (((!g1983) & (g2127) & (g3710)) + ((g1983) & (!g2127) & (g3710)) + ((g1983) & (g2127) & (!g3710)) + ((g1983) & (g2127) & (g3710)));
	assign g4821 = (((g1914) & (!g1985) & (!g2173) & (g4820)) + ((g1914) & (!g1985) & (g2173) & (!g4820)) + ((g1914) & (g1985) & (!g2173) & (!g4820)) + ((g1914) & (g1985) & (g2173) & (g4820)));
	assign g4822 = (((!g2110) & (g2118) & (g3727)) + ((g2110) & (!g2118) & (g3727)) + ((g2110) & (g2118) & (!g3727)) + ((g2110) & (g2118) & (g3727)));
	assign g4823 = (((!g1914) & (!g2156) & (!g2159) & (g4822)) + ((!g1914) & (!g2156) & (g2159) & (!g4822)) + ((!g1914) & (g2156) & (!g2159) & (!g4822)) + ((!g1914) & (g2156) & (g2159) & (g4822)));
	assign g4824 = (((!g830) & (!g2592) & (!g4821) & (!g4823) & (key[205])) + ((!g830) & (!g2592) & (!g4821) & (g4823) & (key[205])) + ((!g830) & (!g2592) & (g4821) & (!g4823) & (key[205])) + ((!g830) & (!g2592) & (g4821) & (g4823) & (key[205])) + ((!g830) & (g2592) & (!g4821) & (!g4823) & (key[205])) + ((!g830) & (g2592) & (!g4821) & (g4823) & (key[205])) + ((!g830) & (g2592) & (g4821) & (!g4823) & (key[205])) + ((!g830) & (g2592) & (g4821) & (g4823) & (key[205])) + ((g830) & (!g2592) & (!g4821) & (g4823) & (!key[205])) + ((g830) & (!g2592) & (!g4821) & (g4823) & (key[205])) + ((g830) & (!g2592) & (g4821) & (!g4823) & (!key[205])) + ((g830) & (!g2592) & (g4821) & (!g4823) & (key[205])) + ((g830) & (!g2592) & (g4821) & (g4823) & (!key[205])) + ((g830) & (!g2592) & (g4821) & (g4823) & (key[205])) + ((g830) & (g2592) & (!g4821) & (!g4823) & (!key[205])) + ((g830) & (g2592) & (!g4821) & (!g4823) & (key[205])));
	assign g4825 = (((!g3157) & (!g3207) & (!g3165) & (g3210) & (!g4772) & (!g4773)) + ((!g3157) & (!g3207) & (!g3165) & (g3210) & (!g4772) & (g4773)) + ((!g3157) & (!g3207) & (!g3165) & (g3210) & (g4772) & (!g4773)) + ((!g3157) & (!g3207) & (!g3165) & (g3210) & (g4772) & (g4773)) + ((!g3157) & (!g3207) & (g3165) & (!g3210) & (!g4772) & (g4773)) + ((!g3157) & (!g3207) & (g3165) & (!g3210) & (g4772) & (!g4773)) + ((!g3157) & (!g3207) & (g3165) & (!g3210) & (g4772) & (g4773)) + ((!g3157) & (!g3207) & (g3165) & (g3210) & (!g4772) & (!g4773)) + ((!g3157) & (g3207) & (!g3165) & (!g3210) & (!g4772) & (!g4773)) + ((!g3157) & (g3207) & (!g3165) & (!g3210) & (!g4772) & (g4773)) + ((!g3157) & (g3207) & (!g3165) & (!g3210) & (g4772) & (!g4773)) + ((!g3157) & (g3207) & (!g3165) & (!g3210) & (g4772) & (g4773)) + ((!g3157) & (g3207) & (g3165) & (!g3210) & (!g4772) & (!g4773)) + ((!g3157) & (g3207) & (g3165) & (g3210) & (!g4772) & (g4773)) + ((!g3157) & (g3207) & (g3165) & (g3210) & (g4772) & (!g4773)) + ((!g3157) & (g3207) & (g3165) & (g3210) & (g4772) & (g4773)) + ((g3157) & (!g3207) & (!g3165) & (!g3210) & (!g4772) & (g4773)) + ((g3157) & (!g3207) & (!g3165) & (!g3210) & (g4772) & (!g4773)) + ((g3157) & (!g3207) & (!g3165) & (!g3210) & (g4772) & (g4773)) + ((g3157) & (!g3207) & (!g3165) & (g3210) & (!g4772) & (!g4773)) + ((g3157) & (!g3207) & (g3165) & (!g3210) & (!g4772) & (!g4773)) + ((g3157) & (!g3207) & (g3165) & (!g3210) & (!g4772) & (g4773)) + ((g3157) & (!g3207) & (g3165) & (!g3210) & (g4772) & (!g4773)) + ((g3157) & (!g3207) & (g3165) & (!g3210) & (g4772) & (g4773)) + ((g3157) & (g3207) & (!g3165) & (!g3210) & (!g4772) & (!g4773)) + ((g3157) & (g3207) & (!g3165) & (g3210) & (!g4772) & (g4773)) + ((g3157) & (g3207) & (!g3165) & (g3210) & (g4772) & (!g4773)) + ((g3157) & (g3207) & (!g3165) & (g3210) & (g4772) & (g4773)) + ((g3157) & (g3207) & (g3165) & (g3210) & (!g4772) & (!g4773)) + ((g3157) & (g3207) & (g3165) & (g3210) & (!g4772) & (g4773)) + ((g3157) & (g3207) & (g3165) & (g3210) & (g4772) & (!g4773)) + ((g3157) & (g3207) & (g3165) & (g3210) & (g4772) & (g4773)));
	assign g4826 = (((!g3168) & (!g3190) & (!g3170) & (g3202) & (!g4775)) + ((!g3168) & (!g3190) & (!g3170) & (g3202) & (g4775)) + ((!g3168) & (!g3190) & (g3170) & (!g3202) & (g4775)) + ((!g3168) & (!g3190) & (g3170) & (g3202) & (!g4775)) + ((!g3168) & (g3190) & (!g3170) & (!g3202) & (!g4775)) + ((!g3168) & (g3190) & (!g3170) & (!g3202) & (g4775)) + ((!g3168) & (g3190) & (g3170) & (!g3202) & (!g4775)) + ((!g3168) & (g3190) & (g3170) & (g3202) & (g4775)) + ((g3168) & (!g3190) & (!g3170) & (!g3202) & (g4775)) + ((g3168) & (!g3190) & (!g3170) & (g3202) & (!g4775)) + ((g3168) & (!g3190) & (g3170) & (!g3202) & (!g4775)) + ((g3168) & (!g3190) & (g3170) & (!g3202) & (g4775)) + ((g3168) & (g3190) & (!g3170) & (!g3202) & (!g4775)) + ((g3168) & (g3190) & (!g3170) & (g3202) & (g4775)) + ((g3168) & (g3190) & (g3170) & (g3202) & (!g4775)) + ((g3168) & (g3190) & (g3170) & (g3202) & (g4775)));
	assign g4827 = (((!g830) & (!g1914) & (!g2595) & (!g4825) & (!g4826)) + ((!g830) & (!g1914) & (!g2595) & (!g4825) & (g4826)) + ((!g830) & (!g1914) & (!g2595) & (g4825) & (!g4826)) + ((!g830) & (!g1914) & (!g2595) & (g4825) & (g4826)) + ((!g830) & (!g1914) & (g2595) & (!g4825) & (!g4826)) + ((!g830) & (!g1914) & (g2595) & (!g4825) & (g4826)) + ((!g830) & (!g1914) & (g2595) & (g4825) & (!g4826)) + ((!g830) & (!g1914) & (g2595) & (g4825) & (g4826)) + ((!g830) & (g1914) & (!g2595) & (!g4825) & (!g4826)) + ((!g830) & (g1914) & (!g2595) & (!g4825) & (g4826)) + ((!g830) & (g1914) & (!g2595) & (g4825) & (!g4826)) + ((!g830) & (g1914) & (!g2595) & (g4825) & (g4826)) + ((!g830) & (g1914) & (g2595) & (!g4825) & (!g4826)) + ((!g830) & (g1914) & (g2595) & (!g4825) & (g4826)) + ((!g830) & (g1914) & (g2595) & (g4825) & (!g4826)) + ((!g830) & (g1914) & (g2595) & (g4825) & (g4826)) + ((g830) & (!g1914) & (!g2595) & (!g4825) & (g4826)) + ((g830) & (!g1914) & (!g2595) & (g4825) & (g4826)) + ((g830) & (!g1914) & (g2595) & (!g4825) & (!g4826)) + ((g830) & (!g1914) & (g2595) & (g4825) & (!g4826)) + ((g830) & (g1914) & (!g2595) & (g4825) & (!g4826)) + ((g830) & (g1914) & (!g2595) & (g4825) & (g4826)) + ((g830) & (g1914) & (g2595) & (!g4825) & (!g4826)) + ((g830) & (g1914) & (g2595) & (!g4825) & (g4826)));
	assign g4828 = (((!g1439) & (!g3511) & (!g2813)) + ((!g1439) & (g3511) & (g2813)) + ((g1439) & (!g3511) & (g2813)) + ((g1439) & (g3511) & (!g2813)));
	assign g4829 = (((!g2804) & (!g2810) & (!g3528)) + ((!g2804) & (g2810) & (g3528)) + ((g2804) & (!g2810) & (g3528)) + ((g2804) & (g2810) & (!g3528)));
	assign g4830 = (((!g830) & (!g1914) & (!g2598) & (!g4828) & (!g4829) & (key[59])) + ((!g830) & (!g1914) & (!g2598) & (!g4828) & (g4829) & (key[59])) + ((!g830) & (!g1914) & (!g2598) & (g4828) & (!g4829) & (key[59])) + ((!g830) & (!g1914) & (!g2598) & (g4828) & (g4829) & (key[59])) + ((!g830) & (!g1914) & (g2598) & (!g4828) & (!g4829) & (key[59])) + ((!g830) & (!g1914) & (g2598) & (!g4828) & (g4829) & (key[59])) + ((!g830) & (!g1914) & (g2598) & (g4828) & (!g4829) & (key[59])) + ((!g830) & (!g1914) & (g2598) & (g4828) & (g4829) & (key[59])) + ((!g830) & (g1914) & (!g2598) & (!g4828) & (!g4829) & (key[59])) + ((!g830) & (g1914) & (!g2598) & (!g4828) & (g4829) & (key[59])) + ((!g830) & (g1914) & (!g2598) & (g4828) & (!g4829) & (key[59])) + ((!g830) & (g1914) & (!g2598) & (g4828) & (g4829) & (key[59])) + ((!g830) & (g1914) & (g2598) & (!g4828) & (!g4829) & (key[59])) + ((!g830) & (g1914) & (g2598) & (!g4828) & (g4829) & (key[59])) + ((!g830) & (g1914) & (g2598) & (g4828) & (!g4829) & (key[59])) + ((!g830) & (g1914) & (g2598) & (g4828) & (g4829) & (key[59])) + ((g830) & (!g1914) & (!g2598) & (!g4828) & (g4829) & (!key[59])) + ((g830) & (!g1914) & (!g2598) & (!g4828) & (g4829) & (key[59])) + ((g830) & (!g1914) & (!g2598) & (g4828) & (g4829) & (!key[59])) + ((g830) & (!g1914) & (!g2598) & (g4828) & (g4829) & (key[59])) + ((g830) & (!g1914) & (g2598) & (!g4828) & (!g4829) & (!key[59])) + ((g830) & (!g1914) & (g2598) & (!g4828) & (!g4829) & (key[59])) + ((g830) & (!g1914) & (g2598) & (g4828) & (!g4829) & (!key[59])) + ((g830) & (!g1914) & (g2598) & (g4828) & (!g4829) & (key[59])) + ((g830) & (g1914) & (!g2598) & (g4828) & (!g4829) & (!key[59])) + ((g830) & (g1914) & (!g2598) & (g4828) & (!g4829) & (key[59])) + ((g830) & (g1914) & (!g2598) & (g4828) & (g4829) & (!key[59])) + ((g830) & (g1914) & (!g2598) & (g4828) & (g4829) & (key[59])) + ((g830) & (g1914) & (g2598) & (!g4828) & (!g4829) & (!key[59])) + ((g830) & (g1914) & (g2598) & (!g4828) & (!g4829) & (key[59])) + ((g830) & (g1914) & (g2598) & (!g4828) & (g4829) & (!key[59])) + ((g830) & (g1914) & (g2598) & (!g4828) & (g4829) & (key[59])));
	assign g4831 = (((!g1972) & (!g1975) & (!g2559) & (g2623) & (!g3753)) + ((!g1972) & (!g1975) & (!g2559) & (g2623) & (g3753)) + ((!g1972) & (!g1975) & (g2559) & (!g2623) & (!g3753)) + ((!g1972) & (!g1975) & (g2559) & (g2623) & (g3753)) + ((!g1972) & (g1975) & (!g2559) & (!g2623) & (!g3753)) + ((!g1972) & (g1975) & (!g2559) & (!g2623) & (g3753)) + ((!g1972) & (g1975) & (g2559) & (!g2623) & (g3753)) + ((!g1972) & (g1975) & (g2559) & (g2623) & (!g3753)) + ((g1972) & (!g1975) & (!g2559) & (!g2623) & (!g3753)) + ((g1972) & (!g1975) & (!g2559) & (g2623) & (g3753)) + ((g1972) & (!g1975) & (g2559) & (!g2623) & (!g3753)) + ((g1972) & (!g1975) & (g2559) & (!g2623) & (g3753)) + ((g1972) & (g1975) & (!g2559) & (!g2623) & (g3753)) + ((g1972) & (g1975) & (!g2559) & (g2623) & (!g3753)) + ((g1972) & (g1975) & (g2559) & (g2623) & (!g3753)) + ((g1972) & (g1975) & (g2559) & (g2623) & (g3753)));
	assign g4832 = (((!g830) & (!g2599) & (!g6431) & (key[91])) + ((!g830) & (!g2599) & (g6431) & (key[91])) + ((!g830) & (g2599) & (!g6431) & (key[91])) + ((!g830) & (g2599) & (g6431) & (key[91])) + ((g830) & (!g2599) & (g6431) & (!key[91])) + ((g830) & (!g2599) & (g6431) & (key[91])) + ((g830) & (g2599) & (!g6431) & (!key[91])) + ((g830) & (g2599) & (!g6431) & (key[91])));
	assign g4833 = (((!g3404) & (!g2804) & (!g2827)) + ((!g3404) & (g2804) & (g2827)) + ((g3404) & (!g2804) & (g2827)) + ((g3404) & (g2804) & (!g2827)));
	assign g4834 = (((!g1439) & (!g3421) & (!g2797)) + ((!g1439) & (g3421) & (g2797)) + ((g1439) & (!g3421) & (g2797)) + ((g1439) & (g3421) & (!g2797)));
	assign g8317 = (((!g5560) & (g5617) & (!g4835)) + ((!g5560) & (g5617) & (g4835)) + ((g5560) & (!g5617) & (g4835)) + ((g5560) & (g5617) & (g4835)));
	assign g4836 = (((!g830) & (!g1914) & (!g2601) & (!g4833) & (!g4834) & (g4835)) + ((!g830) & (!g1914) & (!g2601) & (!g4833) & (g4834) & (g4835)) + ((!g830) & (!g1914) & (!g2601) & (g4833) & (!g4834) & (g4835)) + ((!g830) & (!g1914) & (!g2601) & (g4833) & (g4834) & (g4835)) + ((!g830) & (!g1914) & (g2601) & (!g4833) & (!g4834) & (g4835)) + ((!g830) & (!g1914) & (g2601) & (!g4833) & (g4834) & (g4835)) + ((!g830) & (!g1914) & (g2601) & (g4833) & (!g4834) & (g4835)) + ((!g830) & (!g1914) & (g2601) & (g4833) & (g4834) & (g4835)) + ((!g830) & (g1914) & (!g2601) & (!g4833) & (!g4834) & (g4835)) + ((!g830) & (g1914) & (!g2601) & (!g4833) & (g4834) & (g4835)) + ((!g830) & (g1914) & (!g2601) & (g4833) & (!g4834) & (g4835)) + ((!g830) & (g1914) & (!g2601) & (g4833) & (g4834) & (g4835)) + ((!g830) & (g1914) & (g2601) & (!g4833) & (!g4834) & (g4835)) + ((!g830) & (g1914) & (g2601) & (!g4833) & (g4834) & (g4835)) + ((!g830) & (g1914) & (g2601) & (g4833) & (!g4834) & (g4835)) + ((!g830) & (g1914) & (g2601) & (g4833) & (g4834) & (g4835)) + ((g830) & (!g1914) & (!g2601) & (!g4833) & (g4834) & (!g4835)) + ((g830) & (!g1914) & (!g2601) & (!g4833) & (g4834) & (g4835)) + ((g830) & (!g1914) & (!g2601) & (g4833) & (g4834) & (!g4835)) + ((g830) & (!g1914) & (!g2601) & (g4833) & (g4834) & (g4835)) + ((g830) & (!g1914) & (g2601) & (!g4833) & (!g4834) & (!g4835)) + ((g830) & (!g1914) & (g2601) & (!g4833) & (!g4834) & (g4835)) + ((g830) & (!g1914) & (g2601) & (g4833) & (!g4834) & (!g4835)) + ((g830) & (!g1914) & (g2601) & (g4833) & (!g4834) & (g4835)) + ((g830) & (g1914) & (!g2601) & (g4833) & (!g4834) & (!g4835)) + ((g830) & (g1914) & (!g2601) & (g4833) & (!g4834) & (g4835)) + ((g830) & (g1914) & (!g2601) & (g4833) & (g4834) & (!g4835)) + ((g830) & (g1914) & (!g2601) & (g4833) & (g4834) & (g4835)) + ((g830) & (g1914) & (g2601) & (!g4833) & (!g4834) & (!g4835)) + ((g830) & (g1914) & (g2601) & (!g4833) & (!g4834) & (g4835)) + ((g830) & (g1914) & (g2601) & (!g4833) & (g4834) & (!g4835)) + ((g830) & (g1914) & (g2601) & (!g4833) & (g4834) & (g4835)));
	assign g4837 = (((!g2011) & (!g2013) & (!g2575) & (g2607) & (!g3491)) + ((!g2011) & (!g2013) & (!g2575) & (g2607) & (g3491)) + ((!g2011) & (!g2013) & (g2575) & (!g2607) & (!g3491)) + ((!g2011) & (!g2013) & (g2575) & (g2607) & (g3491)) + ((!g2011) & (g2013) & (!g2575) & (!g2607) & (!g3491)) + ((!g2011) & (g2013) & (!g2575) & (!g2607) & (g3491)) + ((!g2011) & (g2013) & (g2575) & (!g2607) & (g3491)) + ((!g2011) & (g2013) & (g2575) & (g2607) & (!g3491)) + ((g2011) & (!g2013) & (!g2575) & (!g2607) & (!g3491)) + ((g2011) & (!g2013) & (!g2575) & (g2607) & (g3491)) + ((g2011) & (!g2013) & (g2575) & (!g2607) & (!g3491)) + ((g2011) & (!g2013) & (g2575) & (!g2607) & (g3491)) + ((g2011) & (g2013) & (!g2575) & (!g2607) & (g3491)) + ((g2011) & (g2013) & (!g2575) & (g2607) & (!g3491)) + ((g2011) & (g2013) & (g2575) & (g2607) & (!g3491)) + ((g2011) & (g2013) & (g2575) & (g2607) & (g3491)));
	assign g4838 = (((!g830) & (!g2602) & (!g6420) & (key[187])) + ((!g830) & (!g2602) & (g6420) & (key[187])) + ((!g830) & (g2602) & (!g6420) & (key[187])) + ((!g830) & (g2602) & (g6420) & (key[187])) + ((g830) & (!g2602) & (g6420) & (!key[187])) + ((g830) & (!g2602) & (g6420) & (key[187])) + ((g830) & (g2602) & (!g6420) & (!key[187])) + ((g830) & (g2602) & (!g6420) & (key[187])));
	assign g4839 = (((!g1894) & (!g1910) & (!g2034) & (g2038)) + ((!g1894) & (!g1910) & (g2034) & (!g2038)) + ((!g1894) & (g1910) & (!g2034) & (g2038)) + ((!g1894) & (g1910) & (g2034) & (!g2038)) + ((g1894) & (!g1910) & (!g2034) & (g2038)) + ((g1894) & (!g1910) & (g2034) & (!g2038)) + ((g1894) & (g1910) & (!g2034) & (!g2038)) + ((g1894) & (g1910) & (g2034) & (g2038)));
	assign g4840 = (((!g830) & (!g2607) & (!g6409) & (key[110])) + ((!g830) & (!g2607) & (g6409) & (key[110])) + ((!g830) & (g2607) & (!g6409) & (key[110])) + ((!g830) & (g2607) & (g6409) & (key[110])) + ((g830) & (!g2607) & (g6409) & (!key[110])) + ((g830) & (!g2607) & (g6409) & (key[110])) + ((g830) & (g2607) & (!g6409) & (!key[110])) + ((g830) & (g2607) & (!g6409) & (key[110])));
	assign g4841 = (((!g2555) & (!g2601) & (g3161) & (g3187) & (!g4755) & (g4756)) + ((!g2555) & (!g2601) & (g3161) & (g3187) & (g4755) & (!g4756)) + ((!g2555) & (!g2601) & (g3161) & (g3187) & (g4755) & (g4756)) + ((!g2555) & (g2601) & (!g3161) & (g3187) & (!g4755) & (!g4756)) + ((!g2555) & (g2601) & (!g3161) & (g3187) & (!g4755) & (g4756)) + ((!g2555) & (g2601) & (!g3161) & (g3187) & (g4755) & (!g4756)) + ((!g2555) & (g2601) & (!g3161) & (g3187) & (g4755) & (g4756)) + ((!g2555) & (g2601) & (g3161) & (!g3187) & (!g4755) & (g4756)) + ((!g2555) & (g2601) & (g3161) & (!g3187) & (g4755) & (!g4756)) + ((!g2555) & (g2601) & (g3161) & (!g3187) & (g4755) & (g4756)) + ((!g2555) & (g2601) & (g3161) & (g3187) & (!g4755) & (!g4756)) + ((!g2555) & (g2601) & (g3161) & (g3187) & (!g4755) & (g4756)) + ((!g2555) & (g2601) & (g3161) & (g3187) & (g4755) & (!g4756)) + ((!g2555) & (g2601) & (g3161) & (g3187) & (g4755) & (g4756)) + ((g2555) & (!g2601) & (!g3161) & (g3187) & (!g4755) & (g4756)) + ((g2555) & (!g2601) & (!g3161) & (g3187) & (g4755) & (!g4756)) + ((g2555) & (!g2601) & (!g3161) & (g3187) & (g4755) & (g4756)) + ((g2555) & (!g2601) & (g3161) & (g3187) & (!g4755) & (!g4756)) + ((g2555) & (!g2601) & (g3161) & (g3187) & (!g4755) & (g4756)) + ((g2555) & (!g2601) & (g3161) & (g3187) & (g4755) & (!g4756)) + ((g2555) & (!g2601) & (g3161) & (g3187) & (g4755) & (g4756)) + ((g2555) & (g2601) & (!g3161) & (!g3187) & (!g4755) & (g4756)) + ((g2555) & (g2601) & (!g3161) & (!g3187) & (g4755) & (!g4756)) + ((g2555) & (g2601) & (!g3161) & (!g3187) & (g4755) & (g4756)) + ((g2555) & (g2601) & (!g3161) & (g3187) & (!g4755) & (!g4756)) + ((g2555) & (g2601) & (!g3161) & (g3187) & (!g4755) & (g4756)) + ((g2555) & (g2601) & (!g3161) & (g3187) & (g4755) & (!g4756)) + ((g2555) & (g2601) & (!g3161) & (g3187) & (g4755) & (g4756)) + ((g2555) & (g2601) & (g3161) & (!g3187) & (!g4755) & (!g4756)) + ((g2555) & (g2601) & (g3161) & (!g3187) & (!g4755) & (g4756)) + ((g2555) & (g2601) & (g3161) & (!g3187) & (g4755) & (!g4756)) + ((g2555) & (g2601) & (g3161) & (!g3187) & (g4755) & (g4756)) + ((g2555) & (g2601) & (g3161) & (g3187) & (!g4755) & (!g4756)) + ((g2555) & (g2601) & (g3161) & (g3187) & (!g4755) & (g4756)) + ((g2555) & (g2601) & (g3161) & (g3187) & (g4755) & (!g4756)) + ((g2555) & (g2601) & (g3161) & (g3187) & (g4755) & (g4756)));
	assign g4842 = (((!g2551) & (!g2598) & (!g3155) & (!g3196) & (!g4758) & (!g5685)) + ((!g2551) & (!g2598) & (!g3155) & (!g3196) & (g4758) & (!g5685)) + ((!g2551) & (!g2598) & (!g3155) & (g3196) & (!g4758) & (!g5685)) + ((!g2551) & (!g2598) & (!g3155) & (g3196) & (g4758) & (!g5685)) + ((!g2551) & (!g2598) & (g3155) & (!g3196) & (!g4758) & (!g5685)) + ((!g2551) & (!g2598) & (g3155) & (!g3196) & (g4758) & (!g5685)) + ((!g2551) & (!g2598) & (g3155) & (g3196) & (!g4758) & (!g5685)) + ((!g2551) & (!g2598) & (g3155) & (g3196) & (g4758) & (g5685)) + ((!g2551) & (g2598) & (!g3155) & (!g3196) & (!g4758) & (!g5685)) + ((!g2551) & (g2598) & (!g3155) & (!g3196) & (g4758) & (!g5685)) + ((!g2551) & (g2598) & (!g3155) & (g3196) & (!g4758) & (g5685)) + ((!g2551) & (g2598) & (!g3155) & (g3196) & (g4758) & (g5685)) + ((!g2551) & (g2598) & (g3155) & (!g3196) & (!g4758) & (!g5685)) + ((!g2551) & (g2598) & (g3155) & (!g3196) & (g4758) & (g5685)) + ((!g2551) & (g2598) & (g3155) & (g3196) & (!g4758) & (g5685)) + ((!g2551) & (g2598) & (g3155) & (g3196) & (g4758) & (g5685)) + ((g2551) & (!g2598) & (!g3155) & (!g3196) & (!g4758) & (!g5685)) + ((g2551) & (!g2598) & (!g3155) & (!g3196) & (g4758) & (!g5685)) + ((g2551) & (!g2598) & (!g3155) & (g3196) & (!g4758) & (!g5685)) + ((g2551) & (!g2598) & (!g3155) & (g3196) & (g4758) & (g5685)) + ((g2551) & (!g2598) & (g3155) & (!g3196) & (!g4758) & (!g5685)) + ((g2551) & (!g2598) & (g3155) & (!g3196) & (g4758) & (!g5685)) + ((g2551) & (!g2598) & (g3155) & (g3196) & (!g4758) & (g5685)) + ((g2551) & (!g2598) & (g3155) & (g3196) & (g4758) & (g5685)) + ((g2551) & (g2598) & (!g3155) & (!g3196) & (!g4758) & (!g5685)) + ((g2551) & (g2598) & (!g3155) & (!g3196) & (g4758) & (g5685)) + ((g2551) & (g2598) & (!g3155) & (g3196) & (!g4758) & (g5685)) + ((g2551) & (g2598) & (!g3155) & (g3196) & (g4758) & (g5685)) + ((g2551) & (g2598) & (g3155) & (!g3196) & (!g4758) & (g5685)) + ((g2551) & (g2598) & (g3155) & (!g3196) & (g4758) & (g5685)) + ((g2551) & (g2598) & (g3155) & (g3196) & (!g4758) & (g5685)) + ((g2551) & (g2598) & (g3155) & (g3196) & (g4758) & (g5685)));
	assign g4843 = (((!g1890) & (!g1939) & (!g1896) & (g2041)) + ((!g1890) & (!g1939) & (g1896) & (g2041)) + ((!g1890) & (g1939) & (!g1896) & (!g2041)) + ((!g1890) & (g1939) & (g1896) & (!g2041)) + ((g1890) & (!g1939) & (!g1896) & (g2041)) + ((g1890) & (!g1939) & (g1896) & (!g2041)) + ((g1890) & (g1939) & (!g1896) & (!g2041)) + ((g1890) & (g1939) & (g1896) & (g2041)));
	assign g4844 = (((!g830) & (!g2617) & (!g6392) & (nonce[14])) + ((!g830) & (!g2617) & (g6392) & (nonce[14])) + ((!g830) & (g2617) & (!g6392) & (nonce[14])) + ((!g830) & (g2617) & (g6392) & (nonce[14])) + ((g830) & (!g2617) & (g6392) & (!nonce[14])) + ((g830) & (!g2617) & (g6392) & (nonce[14])) + ((g830) & (g2617) & (!g6392) & (!nonce[14])) + ((g830) & (g2617) & (!g6392) & (nonce[14])));
	assign g4845 = (((!g1888) & (!g1978) & (!g1904) & (g2043)) + ((!g1888) & (!g1978) & (g1904) & (g2043)) + ((!g1888) & (g1978) & (!g1904) & (!g2043)) + ((!g1888) & (g1978) & (g1904) & (!g2043)) + ((g1888) & (!g1978) & (!g1904) & (g2043)) + ((g1888) & (!g1978) & (g1904) & (!g2043)) + ((g1888) & (g1978) & (!g1904) & (!g2043)) + ((g1888) & (g1978) & (g1904) & (g2043)));
	assign g4846 = (((!g830) & (!g2620) & (!g6381) & (key[238])) + ((!g830) & (!g2620) & (g6381) & (key[238])) + ((!g830) & (g2620) & (!g6381) & (key[238])) + ((!g830) & (g2620) & (g6381) & (key[238])) + ((g830) & (!g2620) & (g6381) & (!key[238])) + ((g830) & (!g2620) & (g6381) & (key[238])) + ((g830) & (g2620) & (!g6381) & (!key[238])) + ((g830) & (g2620) & (!g6381) & (key[238])));
	assign g4847 = (((!g1900) & (!g2028) & (!g1904) & (g2043)) + ((!g1900) & (!g2028) & (g1904) & (g2043)) + ((!g1900) & (g2028) & (!g1904) & (!g2043)) + ((!g1900) & (g2028) & (g1904) & (!g2043)) + ((g1900) & (!g2028) & (!g1904) & (g2043)) + ((g1900) & (!g2028) & (g1904) & (!g2043)) + ((g1900) & (g2028) & (!g1904) & (!g2043)) + ((g1900) & (g2028) & (g1904) & (g2043)));
	assign g4848 = (((!g830) & (!g2623) & (!g6370) & (key[14])) + ((!g830) & (!g2623) & (g6370) & (key[14])) + ((!g830) & (g2623) & (!g6370) & (key[14])) + ((!g830) & (g2623) & (g6370) & (key[14])) + ((g830) & (!g2623) & (g6370) & (!key[14])) + ((g830) & (!g2623) & (g6370) & (key[14])) + ((g830) & (g2623) & (!g6370) & (!key[14])) + ((g830) & (g2623) & (!g6370) & (key[14])));
	assign g4849 = (((!g1884) & (!g1977) & (!g1908) & (g2030)) + ((!g1884) & (!g1977) & (g1908) & (g2030)) + ((!g1884) & (g1977) & (!g1908) & (!g2030)) + ((!g1884) & (g1977) & (g1908) & (!g2030)) + ((g1884) & (!g1977) & (!g1908) & (g2030)) + ((g1884) & (!g1977) & (g1908) & (!g2030)) + ((g1884) & (g1977) & (!g1908) & (!g2030)) + ((g1884) & (g1977) & (g1908) & (g2030)));
	assign g8318 = (((!g5560) & (g5619) & (!g4850)) + ((!g5560) & (g5619) & (g4850)) + ((g5560) & (!g5619) & (g4850)) + ((g5560) & (g5619) & (g4850)));
	assign g4851 = (((!g830) & (!g2626) & (!g6359) & (g4850)) + ((!g830) & (!g2626) & (g6359) & (g4850)) + ((!g830) & (g2626) & (!g6359) & (g4850)) + ((!g830) & (g2626) & (g6359) & (g4850)) + ((g830) & (!g2626) & (g6359) & (!g4850)) + ((g830) & (!g2626) & (g6359) & (g4850)) + ((g830) & (g2626) & (!g6359) & (!g4850)) + ((g830) & (g2626) & (!g6359) & (g4850)));
	assign g4852 = (((!g3149) & (!g3193) & (g3170) & (g3202) & (!g4761) & (g4762)) + ((!g3149) & (!g3193) & (g3170) & (g3202) & (g4761) & (!g4762)) + ((!g3149) & (!g3193) & (g3170) & (g3202) & (g4761) & (g4762)) + ((!g3149) & (g3193) & (!g3170) & (g3202) & (!g4761) & (!g4762)) + ((!g3149) & (g3193) & (!g3170) & (g3202) & (!g4761) & (g4762)) + ((!g3149) & (g3193) & (!g3170) & (g3202) & (g4761) & (!g4762)) + ((!g3149) & (g3193) & (!g3170) & (g3202) & (g4761) & (g4762)) + ((!g3149) & (g3193) & (g3170) & (!g3202) & (!g4761) & (g4762)) + ((!g3149) & (g3193) & (g3170) & (!g3202) & (g4761) & (!g4762)) + ((!g3149) & (g3193) & (g3170) & (!g3202) & (g4761) & (g4762)) + ((!g3149) & (g3193) & (g3170) & (g3202) & (!g4761) & (!g4762)) + ((!g3149) & (g3193) & (g3170) & (g3202) & (!g4761) & (g4762)) + ((!g3149) & (g3193) & (g3170) & (g3202) & (g4761) & (!g4762)) + ((!g3149) & (g3193) & (g3170) & (g3202) & (g4761) & (g4762)) + ((g3149) & (!g3193) & (!g3170) & (g3202) & (!g4761) & (g4762)) + ((g3149) & (!g3193) & (!g3170) & (g3202) & (g4761) & (!g4762)) + ((g3149) & (!g3193) & (!g3170) & (g3202) & (g4761) & (g4762)) + ((g3149) & (!g3193) & (g3170) & (g3202) & (!g4761) & (!g4762)) + ((g3149) & (!g3193) & (g3170) & (g3202) & (!g4761) & (g4762)) + ((g3149) & (!g3193) & (g3170) & (g3202) & (g4761) & (!g4762)) + ((g3149) & (!g3193) & (g3170) & (g3202) & (g4761) & (g4762)) + ((g3149) & (g3193) & (!g3170) & (!g3202) & (!g4761) & (g4762)) + ((g3149) & (g3193) & (!g3170) & (!g3202) & (g4761) & (!g4762)) + ((g3149) & (g3193) & (!g3170) & (!g3202) & (g4761) & (g4762)) + ((g3149) & (g3193) & (!g3170) & (g3202) & (!g4761) & (!g4762)) + ((g3149) & (g3193) & (!g3170) & (g3202) & (!g4761) & (g4762)) + ((g3149) & (g3193) & (!g3170) & (g3202) & (g4761) & (!g4762)) + ((g3149) & (g3193) & (!g3170) & (g3202) & (g4761) & (g4762)) + ((g3149) & (g3193) & (g3170) & (!g3202) & (!g4761) & (!g4762)) + ((g3149) & (g3193) & (g3170) & (!g3202) & (!g4761) & (g4762)) + ((g3149) & (g3193) & (g3170) & (!g3202) & (g4761) & (!g4762)) + ((g3149) & (g3193) & (g3170) & (!g3202) & (g4761) & (g4762)) + ((g3149) & (g3193) & (g3170) & (g3202) & (!g4761) & (!g4762)) + ((g3149) & (g3193) & (g3170) & (g3202) & (!g4761) & (g4762)) + ((g3149) & (g3193) & (g3170) & (g3202) & (g4761) & (!g4762)) + ((g3149) & (g3193) & (g3170) & (g3202) & (g4761) & (g4762)));
	assign g4853 = (((!g3159) & (!g3177) & (!g3165) & (!g3210) & (!g4764) & (!g5686)) + ((!g3159) & (!g3177) & (!g3165) & (!g3210) & (g4764) & (!g5686)) + ((!g3159) & (!g3177) & (!g3165) & (g3210) & (!g4764) & (!g5686)) + ((!g3159) & (!g3177) & (!g3165) & (g3210) & (g4764) & (!g5686)) + ((!g3159) & (!g3177) & (g3165) & (!g3210) & (!g4764) & (!g5686)) + ((!g3159) & (!g3177) & (g3165) & (!g3210) & (g4764) & (!g5686)) + ((!g3159) & (!g3177) & (g3165) & (g3210) & (!g4764) & (!g5686)) + ((!g3159) & (!g3177) & (g3165) & (g3210) & (g4764) & (g5686)) + ((!g3159) & (g3177) & (!g3165) & (!g3210) & (!g4764) & (!g5686)) + ((!g3159) & (g3177) & (!g3165) & (!g3210) & (g4764) & (!g5686)) + ((!g3159) & (g3177) & (!g3165) & (g3210) & (!g4764) & (g5686)) + ((!g3159) & (g3177) & (!g3165) & (g3210) & (g4764) & (g5686)) + ((!g3159) & (g3177) & (g3165) & (!g3210) & (!g4764) & (!g5686)) + ((!g3159) & (g3177) & (g3165) & (!g3210) & (g4764) & (g5686)) + ((!g3159) & (g3177) & (g3165) & (g3210) & (!g4764) & (g5686)) + ((!g3159) & (g3177) & (g3165) & (g3210) & (g4764) & (g5686)) + ((g3159) & (!g3177) & (!g3165) & (!g3210) & (!g4764) & (!g5686)) + ((g3159) & (!g3177) & (!g3165) & (!g3210) & (g4764) & (!g5686)) + ((g3159) & (!g3177) & (!g3165) & (g3210) & (!g4764) & (!g5686)) + ((g3159) & (!g3177) & (!g3165) & (g3210) & (g4764) & (g5686)) + ((g3159) & (!g3177) & (g3165) & (!g3210) & (!g4764) & (!g5686)) + ((g3159) & (!g3177) & (g3165) & (!g3210) & (g4764) & (!g5686)) + ((g3159) & (!g3177) & (g3165) & (g3210) & (!g4764) & (g5686)) + ((g3159) & (!g3177) & (g3165) & (g3210) & (g4764) & (g5686)) + ((g3159) & (g3177) & (!g3165) & (!g3210) & (!g4764) & (!g5686)) + ((g3159) & (g3177) & (!g3165) & (!g3210) & (g4764) & (g5686)) + ((g3159) & (g3177) & (!g3165) & (g3210) & (!g4764) & (g5686)) + ((g3159) & (g3177) & (!g3165) & (g3210) & (g4764) & (g5686)) + ((g3159) & (g3177) & (g3165) & (!g3210) & (!g4764) & (g5686)) + ((g3159) & (g3177) & (g3165) & (!g3210) & (g4764) & (g5686)) + ((g3159) & (g3177) & (g3165) & (g3210) & (!g4764) & (g5686)) + ((g3159) & (g3177) & (g3165) & (g3210) & (g4764) & (g5686)));
	assign g4854 = (((!g1985) & (!g1987) & (!g2173) & (g2207) & (!g4820)) + ((!g1985) & (!g1987) & (!g2173) & (g2207) & (g4820)) + ((!g1985) & (!g1987) & (g2173) & (!g2207) & (g4820)) + ((!g1985) & (!g1987) & (g2173) & (g2207) & (!g4820)) + ((!g1985) & (g1987) & (!g2173) & (!g2207) & (!g4820)) + ((!g1985) & (g1987) & (!g2173) & (!g2207) & (g4820)) + ((!g1985) & (g1987) & (g2173) & (!g2207) & (!g4820)) + ((!g1985) & (g1987) & (g2173) & (g2207) & (g4820)) + ((g1985) & (!g1987) & (!g2173) & (!g2207) & (g4820)) + ((g1985) & (!g1987) & (!g2173) & (g2207) & (!g4820)) + ((g1985) & (!g1987) & (g2173) & (!g2207) & (!g4820)) + ((g1985) & (!g1987) & (g2173) & (!g2207) & (g4820)) + ((g1985) & (g1987) & (!g2173) & (!g2207) & (!g4820)) + ((g1985) & (g1987) & (!g2173) & (g2207) & (g4820)) + ((g1985) & (g1987) & (g2173) & (g2207) & (!g4820)) + ((g1985) & (g1987) & (g2173) & (g2207) & (g4820)));
	assign g4855 = (((!g2156) & (!g2190) & (!g2159) & (g2198) & (!g4822)) + ((!g2156) & (!g2190) & (!g2159) & (g2198) & (g4822)) + ((!g2156) & (!g2190) & (g2159) & (!g2198) & (g4822)) + ((!g2156) & (!g2190) & (g2159) & (g2198) & (!g4822)) + ((!g2156) & (g2190) & (!g2159) & (!g2198) & (!g4822)) + ((!g2156) & (g2190) & (!g2159) & (!g2198) & (g4822)) + ((!g2156) & (g2190) & (g2159) & (!g2198) & (!g4822)) + ((!g2156) & (g2190) & (g2159) & (g2198) & (g4822)) + ((g2156) & (!g2190) & (!g2159) & (!g2198) & (g4822)) + ((g2156) & (!g2190) & (!g2159) & (g2198) & (!g4822)) + ((g2156) & (!g2190) & (g2159) & (!g2198) & (!g4822)) + ((g2156) & (!g2190) & (g2159) & (!g2198) & (g4822)) + ((g2156) & (g2190) & (!g2159) & (!g2198) & (!g4822)) + ((g2156) & (g2190) & (!g2159) & (g2198) & (g4822)) + ((g2156) & (g2190) & (g2159) & (g2198) & (!g4822)) + ((g2156) & (g2190) & (g2159) & (g2198) & (g4822)));
	assign g4856 = (((!g830) & (!g1914) & (!g2632) & (!g4854) & (!g4855) & (key[206])) + ((!g830) & (!g1914) & (!g2632) & (!g4854) & (g4855) & (key[206])) + ((!g830) & (!g1914) & (!g2632) & (g4854) & (!g4855) & (key[206])) + ((!g830) & (!g1914) & (!g2632) & (g4854) & (g4855) & (key[206])) + ((!g830) & (!g1914) & (g2632) & (!g4854) & (!g4855) & (key[206])) + ((!g830) & (!g1914) & (g2632) & (!g4854) & (g4855) & (key[206])) + ((!g830) & (!g1914) & (g2632) & (g4854) & (!g4855) & (key[206])) + ((!g830) & (!g1914) & (g2632) & (g4854) & (g4855) & (key[206])) + ((!g830) & (g1914) & (!g2632) & (!g4854) & (!g4855) & (key[206])) + ((!g830) & (g1914) & (!g2632) & (!g4854) & (g4855) & (key[206])) + ((!g830) & (g1914) & (!g2632) & (g4854) & (!g4855) & (key[206])) + ((!g830) & (g1914) & (!g2632) & (g4854) & (g4855) & (key[206])) + ((!g830) & (g1914) & (g2632) & (!g4854) & (!g4855) & (key[206])) + ((!g830) & (g1914) & (g2632) & (!g4854) & (g4855) & (key[206])) + ((!g830) & (g1914) & (g2632) & (g4854) & (!g4855) & (key[206])) + ((!g830) & (g1914) & (g2632) & (g4854) & (g4855) & (key[206])) + ((g830) & (!g1914) & (!g2632) & (!g4854) & (g4855) & (!key[206])) + ((g830) & (!g1914) & (!g2632) & (!g4854) & (g4855) & (key[206])) + ((g830) & (!g1914) & (!g2632) & (g4854) & (g4855) & (!key[206])) + ((g830) & (!g1914) & (!g2632) & (g4854) & (g4855) & (key[206])) + ((g830) & (!g1914) & (g2632) & (!g4854) & (!g4855) & (!key[206])) + ((g830) & (!g1914) & (g2632) & (!g4854) & (!g4855) & (key[206])) + ((g830) & (!g1914) & (g2632) & (g4854) & (!g4855) & (!key[206])) + ((g830) & (!g1914) & (g2632) & (g4854) & (!g4855) & (key[206])) + ((g830) & (g1914) & (!g2632) & (g4854) & (!g4855) & (!key[206])) + ((g830) & (g1914) & (!g2632) & (g4854) & (!g4855) & (key[206])) + ((g830) & (g1914) & (!g2632) & (g4854) & (g4855) & (!key[206])) + ((g830) & (g1914) & (!g2632) & (g4854) & (g4855) & (key[206])) + ((g830) & (g1914) & (g2632) & (!g4854) & (!g4855) & (!key[206])) + ((g830) & (g1914) & (g2632) & (!g4854) & (!g4855) & (key[206])) + ((g830) & (g1914) & (g2632) & (!g4854) & (g4855) & (!key[206])) + ((g830) & (g1914) & (g2632) & (!g4854) & (g4855) & (key[206])));
	assign g4857 = (((!g1906) & (!g1940) & (!g1910) & (g2038)) + ((!g1906) & (!g1940) & (g1910) & (g2038)) + ((!g1906) & (g1940) & (!g1910) & (!g2038)) + ((!g1906) & (g1940) & (g1910) & (!g2038)) + ((g1906) & (!g1940) & (!g1910) & (g2038)) + ((g1906) & (!g1940) & (g1910) & (!g2038)) + ((g1906) & (g1940) & (!g1910) & (!g2038)) + ((g1906) & (g1940) & (g1910) & (g2038)));
	assign g4858 = (((!g830) & (!g2637) & (!g6341) & (key[142])) + ((!g830) & (!g2637) & (g6341) & (key[142])) + ((!g830) & (g2637) & (!g6341) & (key[142])) + ((!g830) & (g2637) & (g6341) & (key[142])) + ((g830) & (!g2637) & (g6341) & (!key[142])) + ((g830) & (!g2637) & (g6341) & (key[142])) + ((g830) & (g2637) & (!g6341) & (!key[142])) + ((g830) & (g2637) & (!g6341) & (key[142])));
	assign g4859 = (((!g2147) & (!g2196) & (!g2159) & (g2198) & (!g4812)) + ((!g2147) & (!g2196) & (!g2159) & (g2198) & (g4812)) + ((!g2147) & (!g2196) & (g2159) & (!g2198) & (g4812)) + ((!g2147) & (!g2196) & (g2159) & (g2198) & (!g4812)) + ((!g2147) & (g2196) & (!g2159) & (!g2198) & (!g4812)) + ((!g2147) & (g2196) & (!g2159) & (!g2198) & (g4812)) + ((!g2147) & (g2196) & (g2159) & (!g2198) & (!g4812)) + ((!g2147) & (g2196) & (g2159) & (g2198) & (g4812)) + ((g2147) & (!g2196) & (!g2159) & (!g2198) & (g4812)) + ((g2147) & (!g2196) & (!g2159) & (g2198) & (!g4812)) + ((g2147) & (!g2196) & (g2159) & (!g2198) & (!g4812)) + ((g2147) & (!g2196) & (g2159) & (!g2198) & (g4812)) + ((g2147) & (g2196) & (!g2159) & (!g2198) & (!g4812)) + ((g2147) & (g2196) & (!g2159) & (g2198) & (g4812)) + ((g2147) & (g2196) & (g2159) & (g2198) & (!g4812)) + ((g2147) & (g2196) & (g2159) & (g2198) & (g4812)));
	assign g4860 = (((!g1947) & (!g1949) & (!g2173) & (g2207) & (!g4814)) + ((!g1947) & (!g1949) & (!g2173) & (g2207) & (g4814)) + ((!g1947) & (!g1949) & (g2173) & (!g2207) & (g4814)) + ((!g1947) & (!g1949) & (g2173) & (g2207) & (!g4814)) + ((!g1947) & (g1949) & (!g2173) & (!g2207) & (!g4814)) + ((!g1947) & (g1949) & (!g2173) & (!g2207) & (g4814)) + ((!g1947) & (g1949) & (g2173) & (!g2207) & (!g4814)) + ((!g1947) & (g1949) & (g2173) & (g2207) & (g4814)) + ((g1947) & (!g1949) & (!g2173) & (!g2207) & (g4814)) + ((g1947) & (!g1949) & (!g2173) & (g2207) & (!g4814)) + ((g1947) & (!g1949) & (g2173) & (!g2207) & (!g4814)) + ((g1947) & (!g1949) & (g2173) & (!g2207) & (g4814)) + ((g1947) & (g1949) & (!g2173) & (!g2207) & (!g4814)) + ((g1947) & (g1949) & (!g2173) & (g2207) & (g4814)) + ((g1947) & (g1949) & (g2173) & (g2207) & (!g4814)) + ((g1947) & (g1949) & (g2173) & (g2207) & (g4814)));
	assign g4861 = (((!g830) & (!g1914) & (!g2640) & (!g4859) & (!g4860) & (nonce[46])) + ((!g830) & (!g1914) & (!g2640) & (!g4859) & (g4860) & (nonce[46])) + ((!g830) & (!g1914) & (!g2640) & (g4859) & (!g4860) & (nonce[46])) + ((!g830) & (!g1914) & (!g2640) & (g4859) & (g4860) & (nonce[46])) + ((!g830) & (!g1914) & (g2640) & (!g4859) & (!g4860) & (nonce[46])) + ((!g830) & (!g1914) & (g2640) & (!g4859) & (g4860) & (nonce[46])) + ((!g830) & (!g1914) & (g2640) & (g4859) & (!g4860) & (nonce[46])) + ((!g830) & (!g1914) & (g2640) & (g4859) & (g4860) & (nonce[46])) + ((!g830) & (g1914) & (!g2640) & (!g4859) & (!g4860) & (nonce[46])) + ((!g830) & (g1914) & (!g2640) & (!g4859) & (g4860) & (nonce[46])) + ((!g830) & (g1914) & (!g2640) & (g4859) & (!g4860) & (nonce[46])) + ((!g830) & (g1914) & (!g2640) & (g4859) & (g4860) & (nonce[46])) + ((!g830) & (g1914) & (g2640) & (!g4859) & (!g4860) & (nonce[46])) + ((!g830) & (g1914) & (g2640) & (!g4859) & (g4860) & (nonce[46])) + ((!g830) & (g1914) & (g2640) & (g4859) & (!g4860) & (nonce[46])) + ((!g830) & (g1914) & (g2640) & (g4859) & (g4860) & (nonce[46])) + ((g830) & (!g1914) & (!g2640) & (!g4859) & (g4860) & (!nonce[46])) + ((g830) & (!g1914) & (!g2640) & (!g4859) & (g4860) & (nonce[46])) + ((g830) & (!g1914) & (!g2640) & (g4859) & (g4860) & (!nonce[46])) + ((g830) & (!g1914) & (!g2640) & (g4859) & (g4860) & (nonce[46])) + ((g830) & (!g1914) & (g2640) & (!g4859) & (!g4860) & (!nonce[46])) + ((g830) & (!g1914) & (g2640) & (!g4859) & (!g4860) & (nonce[46])) + ((g830) & (!g1914) & (g2640) & (g4859) & (!g4860) & (!nonce[46])) + ((g830) & (!g1914) & (g2640) & (g4859) & (!g4860) & (nonce[46])) + ((g830) & (g1914) & (!g2640) & (g4859) & (!g4860) & (!nonce[46])) + ((g830) & (g1914) & (!g2640) & (g4859) & (!g4860) & (nonce[46])) + ((g830) & (g1914) & (!g2640) & (g4859) & (g4860) & (!nonce[46])) + ((g830) & (g1914) & (!g2640) & (g4859) & (g4860) & (nonce[46])) + ((g830) & (g1914) & (g2640) & (!g4859) & (!g4860) & (!nonce[46])) + ((g830) & (g1914) & (g2640) & (!g4859) & (!g4860) & (nonce[46])) + ((g830) & (g1914) & (g2640) & (!g4859) & (g4860) & (!nonce[46])) + ((g830) & (g1914) & (g2640) & (!g4859) & (g4860) & (nonce[46])));
	assign g4862 = (((!g3157) & (!g3207) & (g3165) & (g3210) & (!g4772) & (g4773)) + ((!g3157) & (!g3207) & (g3165) & (g3210) & (g4772) & (!g4773)) + ((!g3157) & (!g3207) & (g3165) & (g3210) & (g4772) & (g4773)) + ((!g3157) & (g3207) & (!g3165) & (g3210) & (!g4772) & (!g4773)) + ((!g3157) & (g3207) & (!g3165) & (g3210) & (!g4772) & (g4773)) + ((!g3157) & (g3207) & (!g3165) & (g3210) & (g4772) & (!g4773)) + ((!g3157) & (g3207) & (!g3165) & (g3210) & (g4772) & (g4773)) + ((!g3157) & (g3207) & (g3165) & (!g3210) & (!g4772) & (g4773)) + ((!g3157) & (g3207) & (g3165) & (!g3210) & (g4772) & (!g4773)) + ((!g3157) & (g3207) & (g3165) & (!g3210) & (g4772) & (g4773)) + ((!g3157) & (g3207) & (g3165) & (g3210) & (!g4772) & (!g4773)) + ((!g3157) & (g3207) & (g3165) & (g3210) & (!g4772) & (g4773)) + ((!g3157) & (g3207) & (g3165) & (g3210) & (g4772) & (!g4773)) + ((!g3157) & (g3207) & (g3165) & (g3210) & (g4772) & (g4773)) + ((g3157) & (!g3207) & (!g3165) & (g3210) & (!g4772) & (g4773)) + ((g3157) & (!g3207) & (!g3165) & (g3210) & (g4772) & (!g4773)) + ((g3157) & (!g3207) & (!g3165) & (g3210) & (g4772) & (g4773)) + ((g3157) & (!g3207) & (g3165) & (g3210) & (!g4772) & (!g4773)) + ((g3157) & (!g3207) & (g3165) & (g3210) & (!g4772) & (g4773)) + ((g3157) & (!g3207) & (g3165) & (g3210) & (g4772) & (!g4773)) + ((g3157) & (!g3207) & (g3165) & (g3210) & (g4772) & (g4773)) + ((g3157) & (g3207) & (!g3165) & (!g3210) & (!g4772) & (g4773)) + ((g3157) & (g3207) & (!g3165) & (!g3210) & (g4772) & (!g4773)) + ((g3157) & (g3207) & (!g3165) & (!g3210) & (g4772) & (g4773)) + ((g3157) & (g3207) & (!g3165) & (g3210) & (!g4772) & (!g4773)) + ((g3157) & (g3207) & (!g3165) & (g3210) & (!g4772) & (g4773)) + ((g3157) & (g3207) & (!g3165) & (g3210) & (g4772) & (!g4773)) + ((g3157) & (g3207) & (!g3165) & (g3210) & (g4772) & (g4773)) + ((g3157) & (g3207) & (g3165) & (!g3210) & (!g4772) & (!g4773)) + ((g3157) & (g3207) & (g3165) & (!g3210) & (!g4772) & (g4773)) + ((g3157) & (g3207) & (g3165) & (!g3210) & (g4772) & (!g4773)) + ((g3157) & (g3207) & (g3165) & (!g3210) & (g4772) & (g4773)) + ((g3157) & (g3207) & (g3165) & (g3210) & (!g4772) & (!g4773)) + ((g3157) & (g3207) & (g3165) & (g3210) & (!g4772) & (g4773)) + ((g3157) & (g3207) & (g3165) & (g3210) & (g4772) & (!g4773)) + ((g3157) & (g3207) & (g3165) & (g3210) & (g4772) & (g4773)));
	assign g4863 = (((!g3168) & (!g3190) & (!g3170) & (!g3202) & (!g4775) & (!g5687)) + ((!g3168) & (!g3190) & (!g3170) & (!g3202) & (g4775) & (!g5687)) + ((!g3168) & (!g3190) & (!g3170) & (g3202) & (!g4775) & (!g5687)) + ((!g3168) & (!g3190) & (!g3170) & (g3202) & (g4775) & (!g5687)) + ((!g3168) & (!g3190) & (g3170) & (!g3202) & (!g4775) & (!g5687)) + ((!g3168) & (!g3190) & (g3170) & (!g3202) & (g4775) & (!g5687)) + ((!g3168) & (!g3190) & (g3170) & (g3202) & (!g4775) & (!g5687)) + ((!g3168) & (!g3190) & (g3170) & (g3202) & (g4775) & (g5687)) + ((!g3168) & (g3190) & (!g3170) & (!g3202) & (!g4775) & (!g5687)) + ((!g3168) & (g3190) & (!g3170) & (!g3202) & (g4775) & (!g5687)) + ((!g3168) & (g3190) & (!g3170) & (g3202) & (!g4775) & (g5687)) + ((!g3168) & (g3190) & (!g3170) & (g3202) & (g4775) & (g5687)) + ((!g3168) & (g3190) & (g3170) & (!g3202) & (!g4775) & (!g5687)) + ((!g3168) & (g3190) & (g3170) & (!g3202) & (g4775) & (g5687)) + ((!g3168) & (g3190) & (g3170) & (g3202) & (!g4775) & (g5687)) + ((!g3168) & (g3190) & (g3170) & (g3202) & (g4775) & (g5687)) + ((g3168) & (!g3190) & (!g3170) & (!g3202) & (!g4775) & (!g5687)) + ((g3168) & (!g3190) & (!g3170) & (!g3202) & (g4775) & (!g5687)) + ((g3168) & (!g3190) & (!g3170) & (g3202) & (!g4775) & (!g5687)) + ((g3168) & (!g3190) & (!g3170) & (g3202) & (g4775) & (g5687)) + ((g3168) & (!g3190) & (g3170) & (!g3202) & (!g4775) & (!g5687)) + ((g3168) & (!g3190) & (g3170) & (!g3202) & (g4775) & (!g5687)) + ((g3168) & (!g3190) & (g3170) & (g3202) & (!g4775) & (g5687)) + ((g3168) & (!g3190) & (g3170) & (g3202) & (g4775) & (g5687)) + ((g3168) & (g3190) & (!g3170) & (!g3202) & (!g4775) & (!g5687)) + ((g3168) & (g3190) & (!g3170) & (!g3202) & (g4775) & (g5687)) + ((g3168) & (g3190) & (!g3170) & (g3202) & (!g4775) & (g5687)) + ((g3168) & (g3190) & (!g3170) & (g3202) & (g4775) & (g5687)) + ((g3168) & (g3190) & (g3170) & (!g3202) & (!g4775) & (g5687)) + ((g3168) & (g3190) & (g3170) & (!g3202) & (g4775) & (g5687)) + ((g3168) & (g3190) & (g3170) & (g3202) & (!g4775) & (g5687)) + ((g3168) & (g3190) & (g3170) & (g3202) & (g4775) & (g5687)));
	assign g4864 = (((!g1439) & (!g3511) & (g2813)) + ((g1439) & (!g3511) & (!g2813)) + ((g1439) & (!g3511) & (g2813)) + ((g1439) & (g3511) & (g2813)));
	assign g4865 = (((g1914) & (!g1473) & (!g4864) & (g2838)) + ((g1914) & (!g1473) & (g4864) & (!g2838)) + ((g1914) & (g1473) & (!g4864) & (!g2838)) + ((g1914) & (g1473) & (g4864) & (g2838)));
	assign g4866 = (((!g2804) & (g2810) & (!g3528)) + ((g2804) & (!g2810) & (!g3528)) + ((g2804) & (g2810) & (!g3528)) + ((g2804) & (g2810) & (g3528)));
	assign g4867 = (((!g1914) & (!g2845) & (!g2868) & (g4866)) + ((!g1914) & (!g2845) & (g2868) & (!g4866)) + ((!g1914) & (g2845) & (!g2868) & (!g4866)) + ((!g1914) & (g2845) & (g2868) & (g4866)));
	assign g4868 = (((!g830) & (!g2647) & (!g4865) & (!g4867) & (key[60])) + ((!g830) & (!g2647) & (!g4865) & (g4867) & (key[60])) + ((!g830) & (!g2647) & (g4865) & (!g4867) & (key[60])) + ((!g830) & (!g2647) & (g4865) & (g4867) & (key[60])) + ((!g830) & (g2647) & (!g4865) & (!g4867) & (key[60])) + ((!g830) & (g2647) & (!g4865) & (g4867) & (key[60])) + ((!g830) & (g2647) & (g4865) & (!g4867) & (key[60])) + ((!g830) & (g2647) & (g4865) & (g4867) & (key[60])) + ((g830) & (!g2647) & (!g4865) & (g4867) & (!key[60])) + ((g830) & (!g2647) & (!g4865) & (g4867) & (key[60])) + ((g830) & (!g2647) & (g4865) & (!g4867) & (!key[60])) + ((g830) & (!g2647) & (g4865) & (!g4867) & (key[60])) + ((g830) & (!g2647) & (g4865) & (g4867) & (!key[60])) + ((g830) & (!g2647) & (g4865) & (g4867) & (key[60])) + ((g830) & (g2647) & (!g4865) & (!g4867) & (!key[60])) + ((g830) & (g2647) & (!g4865) & (!g4867) & (key[60])));
	assign g4869 = (((!g1972) & (!g1975) & (g2559) & (g2623) & (!g3753)) + ((!g1972) & (g1975) & (!g2559) & (g2623) & (!g3753)) + ((!g1972) & (g1975) & (!g2559) & (g2623) & (g3753)) + ((!g1972) & (g1975) & (g2559) & (!g2623) & (!g3753)) + ((!g1972) & (g1975) & (g2559) & (g2623) & (!g3753)) + ((!g1972) & (g1975) & (g2559) & (g2623) & (g3753)) + ((g1972) & (!g1975) & (!g2559) & (g2623) & (!g3753)) + ((g1972) & (!g1975) & (g2559) & (g2623) & (!g3753)) + ((g1972) & (!g1975) & (g2559) & (g2623) & (g3753)) + ((g1972) & (g1975) & (!g2559) & (!g2623) & (!g3753)) + ((g1972) & (g1975) & (!g2559) & (g2623) & (!g3753)) + ((g1972) & (g1975) & (!g2559) & (g2623) & (g3753)) + ((g1972) & (g1975) & (g2559) & (!g2623) & (!g3753)) + ((g1972) & (g1975) & (g2559) & (!g2623) & (g3753)) + ((g1972) & (g1975) & (g2559) & (g2623) & (!g3753)) + ((g1972) & (g1975) & (g2559) & (g2623) & (g3753)));
	assign g4870 = (((!g2047) & (!g2653) & (g4869)) + ((!g2047) & (g2653) & (!g4869)) + ((g2047) & (!g2653) & (!g4869)) + ((g2047) & (g2653) & (g4869)));
	assign g4871 = (((!g2944) & (!g2991) & (!g3772) & (g3773)) + ((!g2944) & (!g2991) & (g3772) & (!g3773)) + ((!g2944) & (!g2991) & (g3772) & (g3773)) + ((!g2944) & (g2991) & (!g3772) & (!g3773)) + ((g2944) & (!g2991) & (!g3772) & (!g3773)) + ((g2944) & (g2991) & (!g3772) & (g3773)) + ((g2944) & (g2991) & (g3772) & (!g3773)) + ((g2944) & (g2991) & (g3772) & (g3773)));
	assign g4872 = (((!g830) & (!g1914) & (!g2648) & (!g4870) & (!g4871) & (key[92])) + ((!g830) & (!g1914) & (!g2648) & (!g4870) & (g4871) & (key[92])) + ((!g830) & (!g1914) & (!g2648) & (g4870) & (!g4871) & (key[92])) + ((!g830) & (!g1914) & (!g2648) & (g4870) & (g4871) & (key[92])) + ((!g830) & (!g1914) & (g2648) & (!g4870) & (!g4871) & (key[92])) + ((!g830) & (!g1914) & (g2648) & (!g4870) & (g4871) & (key[92])) + ((!g830) & (!g1914) & (g2648) & (g4870) & (!g4871) & (key[92])) + ((!g830) & (!g1914) & (g2648) & (g4870) & (g4871) & (key[92])) + ((!g830) & (g1914) & (!g2648) & (!g4870) & (!g4871) & (key[92])) + ((!g830) & (g1914) & (!g2648) & (!g4870) & (g4871) & (key[92])) + ((!g830) & (g1914) & (!g2648) & (g4870) & (!g4871) & (key[92])) + ((!g830) & (g1914) & (!g2648) & (g4870) & (g4871) & (key[92])) + ((!g830) & (g1914) & (g2648) & (!g4870) & (!g4871) & (key[92])) + ((!g830) & (g1914) & (g2648) & (!g4870) & (g4871) & (key[92])) + ((!g830) & (g1914) & (g2648) & (g4870) & (!g4871) & (key[92])) + ((!g830) & (g1914) & (g2648) & (g4870) & (g4871) & (key[92])) + ((g830) & (!g1914) & (!g2648) & (!g4870) & (g4871) & (!key[92])) + ((g830) & (!g1914) & (!g2648) & (!g4870) & (g4871) & (key[92])) + ((g830) & (!g1914) & (!g2648) & (g4870) & (g4871) & (!key[92])) + ((g830) & (!g1914) & (!g2648) & (g4870) & (g4871) & (key[92])) + ((g830) & (!g1914) & (g2648) & (!g4870) & (!g4871) & (!key[92])) + ((g830) & (!g1914) & (g2648) & (!g4870) & (!g4871) & (key[92])) + ((g830) & (!g1914) & (g2648) & (g4870) & (!g4871) & (!key[92])) + ((g830) & (!g1914) & (g2648) & (g4870) & (!g4871) & (key[92])) + ((g830) & (g1914) & (!g2648) & (g4870) & (!g4871) & (!key[92])) + ((g830) & (g1914) & (!g2648) & (g4870) & (!g4871) & (key[92])) + ((g830) & (g1914) & (!g2648) & (g4870) & (g4871) & (!key[92])) + ((g830) & (g1914) & (!g2648) & (g4870) & (g4871) & (key[92])) + ((g830) & (g1914) & (g2648) & (!g4870) & (!g4871) & (!key[92])) + ((g830) & (g1914) & (g2648) & (!g4870) & (!g4871) & (key[92])) + ((g830) & (g1914) & (g2648) & (!g4870) & (g4871) & (!key[92])) + ((g830) & (g1914) & (g2648) & (!g4870) & (g4871) & (key[92])));
	assign g4873 = (((!g1439) & (!g3421) & (g2797)) + ((g1439) & (!g3421) & (!g2797)) + ((g1439) & (!g3421) & (g2797)) + ((g1439) & (g3421) & (g2797)));
	assign g4874 = (((!g3404) & (!g2804) & (g2827)) + ((!g3404) & (g2804) & (!g2827)) + ((!g3404) & (g2804) & (g2827)) + ((g3404) & (g2804) & (g2827)));
	assign g4875 = (((!g4874) & (!g2845) & (g2851)) + ((!g4874) & (g2845) & (!g2851)) + ((g4874) & (!g2845) & (!g2851)) + ((g4874) & (g2845) & (g2851)));
	assign g4876 = (((!g1914) & (!g1473) & (!g4873) & (g2854) & (!g4875)) + ((!g1914) & (!g1473) & (!g4873) & (g2854) & (g4875)) + ((!g1914) & (!g1473) & (g4873) & (!g2854) & (!g4875)) + ((!g1914) & (!g1473) & (g4873) & (!g2854) & (g4875)) + ((!g1914) & (g1473) & (!g4873) & (!g2854) & (!g4875)) + ((!g1914) & (g1473) & (!g4873) & (!g2854) & (g4875)) + ((!g1914) & (g1473) & (g4873) & (g2854) & (!g4875)) + ((!g1914) & (g1473) & (g4873) & (g2854) & (g4875)) + ((g1914) & (!g1473) & (!g4873) & (!g2854) & (g4875)) + ((g1914) & (!g1473) & (!g4873) & (g2854) & (g4875)) + ((g1914) & (!g1473) & (g4873) & (!g2854) & (g4875)) + ((g1914) & (!g1473) & (g4873) & (g2854) & (g4875)) + ((g1914) & (g1473) & (!g4873) & (!g2854) & (g4875)) + ((g1914) & (g1473) & (!g4873) & (g2854) & (g4875)) + ((g1914) & (g1473) & (g4873) & (!g2854) & (g4875)) + ((g1914) & (g1473) & (g4873) & (g2854) & (g4875)));
	assign g8319 = (((!g5560) & (g5620) & (!g4877)) + ((!g5560) & (g5620) & (g4877)) + ((g5560) & (!g5620) & (g4877)) + ((g5560) & (g5620) & (g4877)));
	assign g4878 = (((!g830) & (!g2649) & (!g4876) & (g4877)) + ((!g830) & (!g2649) & (g4876) & (g4877)) + ((!g830) & (g2649) & (!g4876) & (g4877)) + ((!g830) & (g2649) & (g4876) & (g4877)) + ((g830) & (!g2649) & (g4876) & (!g4877)) + ((g830) & (!g2649) & (g4876) & (g4877)) + ((g830) & (g2649) & (!g4876) & (!g4877)) + ((g830) & (g2649) & (!g4876) & (g4877)));
	assign g4879 = (((!g3479) & (!g3480) & (!g2979) & (g2991)) + ((!g3479) & (!g3480) & (g2979) & (!g2991)) + ((!g3479) & (g3480) & (!g2979) & (!g2991)) + ((!g3479) & (g3480) & (g2979) & (g2991)) + ((g3479) & (!g3480) & (!g2979) & (!g2991)) + ((g3479) & (!g3480) & (g2979) & (g2991)) + ((g3479) & (g3480) & (!g2979) & (!g2991)) + ((g3479) & (g3480) & (g2979) & (g2991)));
	assign g4880 = (((!g2011) & (!g2013) & (g2575) & (g2607) & (!g3491)) + ((!g2011) & (g2013) & (!g2575) & (g2607) & (!g3491)) + ((!g2011) & (g2013) & (!g2575) & (g2607) & (g3491)) + ((!g2011) & (g2013) & (g2575) & (!g2607) & (!g3491)) + ((!g2011) & (g2013) & (g2575) & (g2607) & (!g3491)) + ((!g2011) & (g2013) & (g2575) & (g2607) & (g3491)) + ((g2011) & (!g2013) & (!g2575) & (g2607) & (!g3491)) + ((g2011) & (!g2013) & (g2575) & (g2607) & (!g3491)) + ((g2011) & (!g2013) & (g2575) & (g2607) & (g3491)) + ((g2011) & (g2013) & (!g2575) & (!g2607) & (!g3491)) + ((g2011) & (g2013) & (!g2575) & (g2607) & (!g3491)) + ((g2011) & (g2013) & (!g2575) & (g2607) & (g3491)) + ((g2011) & (g2013) & (g2575) & (!g2607) & (!g3491)) + ((g2011) & (g2013) & (g2575) & (!g2607) & (g3491)) + ((g2011) & (g2013) & (g2575) & (g2607) & (!g3491)) + ((g2011) & (g2013) & (g2575) & (g2607) & (g3491)));
	assign g4881 = (((!g2051) & (!g2663) & (g4880)) + ((!g2051) & (g2663) & (!g4880)) + ((g2051) & (!g2663) & (!g4880)) + ((g2051) & (g2663) & (g4880)));
	assign g4882 = (((!g830) & (!g1914) & (!g2650) & (!g4879) & (!g4881) & (key[188])) + ((!g830) & (!g1914) & (!g2650) & (!g4879) & (g4881) & (key[188])) + ((!g830) & (!g1914) & (!g2650) & (g4879) & (!g4881) & (key[188])) + ((!g830) & (!g1914) & (!g2650) & (g4879) & (g4881) & (key[188])) + ((!g830) & (!g1914) & (g2650) & (!g4879) & (!g4881) & (key[188])) + ((!g830) & (!g1914) & (g2650) & (!g4879) & (g4881) & (key[188])) + ((!g830) & (!g1914) & (g2650) & (g4879) & (!g4881) & (key[188])) + ((!g830) & (!g1914) & (g2650) & (g4879) & (g4881) & (key[188])) + ((!g830) & (g1914) & (!g2650) & (!g4879) & (!g4881) & (key[188])) + ((!g830) & (g1914) & (!g2650) & (!g4879) & (g4881) & (key[188])) + ((!g830) & (g1914) & (!g2650) & (g4879) & (!g4881) & (key[188])) + ((!g830) & (g1914) & (!g2650) & (g4879) & (g4881) & (key[188])) + ((!g830) & (g1914) & (g2650) & (!g4879) & (!g4881) & (key[188])) + ((!g830) & (g1914) & (g2650) & (!g4879) & (g4881) & (key[188])) + ((!g830) & (g1914) & (g2650) & (g4879) & (!g4881) & (key[188])) + ((!g830) & (g1914) & (g2650) & (g4879) & (g4881) & (key[188])) + ((g830) & (!g1914) & (!g2650) & (!g4879) & (g4881) & (!key[188])) + ((g830) & (!g1914) & (!g2650) & (!g4879) & (g4881) & (key[188])) + ((g830) & (!g1914) & (!g2650) & (g4879) & (g4881) & (!key[188])) + ((g830) & (!g1914) & (!g2650) & (g4879) & (g4881) & (key[188])) + ((g830) & (!g1914) & (g2650) & (!g4879) & (!g4881) & (!key[188])) + ((g830) & (!g1914) & (g2650) & (!g4879) & (!g4881) & (key[188])) + ((g830) & (!g1914) & (g2650) & (g4879) & (!g4881) & (!key[188])) + ((g830) & (!g1914) & (g2650) & (g4879) & (!g4881) & (key[188])) + ((g830) & (g1914) & (!g2650) & (g4879) & (!g4881) & (!key[188])) + ((g830) & (g1914) & (!g2650) & (g4879) & (!g4881) & (key[188])) + ((g830) & (g1914) & (!g2650) & (g4879) & (g4881) & (!key[188])) + ((g830) & (g1914) & (!g2650) & (g4879) & (g4881) & (key[188])) + ((g830) & (g1914) & (g2650) & (!g4879) & (!g4881) & (!key[188])) + ((g830) & (g1914) & (g2650) & (!g4879) & (!g4881) & (key[188])) + ((g830) & (g1914) & (g2650) & (!g4879) & (g4881) & (!key[188])) + ((g830) & (g1914) & (g2650) & (!g4879) & (g4881) & (key[188])));
	assign g4883 = (((!g1959) & (!g1098) & (!g3625)) + ((!g1959) & (g1098) & (g3625)) + ((g1959) & (!g1098) & (g3625)) + ((g1959) & (g1098) & (!g3625)));
	assign g4884 = (((!g1900) & (!g2028) & (!g2074) & (!g1904) & (!g2043) & (g2080)) + ((!g1900) & (!g2028) & (!g2074) & (!g1904) & (g2043) & (g2080)) + ((!g1900) & (!g2028) & (!g2074) & (g1904) & (!g2043) & (g2080)) + ((!g1900) & (!g2028) & (!g2074) & (g1904) & (g2043) & (g2080)) + ((!g1900) & (!g2028) & (g2074) & (!g1904) & (!g2043) & (!g2080)) + ((!g1900) & (!g2028) & (g2074) & (!g1904) & (g2043) & (!g2080)) + ((!g1900) & (!g2028) & (g2074) & (g1904) & (!g2043) & (!g2080)) + ((!g1900) & (!g2028) & (g2074) & (g1904) & (g2043) & (!g2080)) + ((!g1900) & (g2028) & (!g2074) & (!g1904) & (!g2043) & (g2080)) + ((!g1900) & (g2028) & (!g2074) & (!g1904) & (g2043) & (!g2080)) + ((!g1900) & (g2028) & (!g2074) & (g1904) & (!g2043) & (g2080)) + ((!g1900) & (g2028) & (!g2074) & (g1904) & (g2043) & (!g2080)) + ((!g1900) & (g2028) & (g2074) & (!g1904) & (!g2043) & (!g2080)) + ((!g1900) & (g2028) & (g2074) & (!g1904) & (g2043) & (g2080)) + ((!g1900) & (g2028) & (g2074) & (g1904) & (!g2043) & (!g2080)) + ((!g1900) & (g2028) & (g2074) & (g1904) & (g2043) & (g2080)) + ((g1900) & (!g2028) & (!g2074) & (!g1904) & (!g2043) & (g2080)) + ((g1900) & (!g2028) & (!g2074) & (!g1904) & (g2043) & (g2080)) + ((g1900) & (!g2028) & (!g2074) & (g1904) & (!g2043) & (g2080)) + ((g1900) & (!g2028) & (!g2074) & (g1904) & (g2043) & (!g2080)) + ((g1900) & (!g2028) & (g2074) & (!g1904) & (!g2043) & (!g2080)) + ((g1900) & (!g2028) & (g2074) & (!g1904) & (g2043) & (!g2080)) + ((g1900) & (!g2028) & (g2074) & (g1904) & (!g2043) & (!g2080)) + ((g1900) & (!g2028) & (g2074) & (g1904) & (g2043) & (g2080)) + ((g1900) & (g2028) & (!g2074) & (!g1904) & (!g2043) & (g2080)) + ((g1900) & (g2028) & (!g2074) & (!g1904) & (g2043) & (!g2080)) + ((g1900) & (g2028) & (!g2074) & (g1904) & (!g2043) & (!g2080)) + ((g1900) & (g2028) & (!g2074) & (g1904) & (g2043) & (!g2080)) + ((g1900) & (g2028) & (g2074) & (!g1904) & (!g2043) & (!g2080)) + ((g1900) & (g2028) & (g2074) & (!g1904) & (g2043) & (g2080)) + ((g1900) & (g2028) & (g2074) & (g1904) & (!g2043) & (g2080)) + ((g1900) & (g2028) & (g2074) & (g1904) & (g2043) & (g2080)));
	assign g4885 = (((!g830) & (!g1914) & (!g2653) & (!g4883) & (!g4884) & (key[15])) + ((!g830) & (!g1914) & (!g2653) & (!g4883) & (g4884) & (key[15])) + ((!g830) & (!g1914) & (!g2653) & (g4883) & (!g4884) & (key[15])) + ((!g830) & (!g1914) & (!g2653) & (g4883) & (g4884) & (key[15])) + ((!g830) & (!g1914) & (g2653) & (!g4883) & (!g4884) & (key[15])) + ((!g830) & (!g1914) & (g2653) & (!g4883) & (g4884) & (key[15])) + ((!g830) & (!g1914) & (g2653) & (g4883) & (!g4884) & (key[15])) + ((!g830) & (!g1914) & (g2653) & (g4883) & (g4884) & (key[15])) + ((!g830) & (g1914) & (!g2653) & (!g4883) & (!g4884) & (key[15])) + ((!g830) & (g1914) & (!g2653) & (!g4883) & (g4884) & (key[15])) + ((!g830) & (g1914) & (!g2653) & (g4883) & (!g4884) & (key[15])) + ((!g830) & (g1914) & (!g2653) & (g4883) & (g4884) & (key[15])) + ((!g830) & (g1914) & (g2653) & (!g4883) & (!g4884) & (key[15])) + ((!g830) & (g1914) & (g2653) & (!g4883) & (g4884) & (key[15])) + ((!g830) & (g1914) & (g2653) & (g4883) & (!g4884) & (key[15])) + ((!g830) & (g1914) & (g2653) & (g4883) & (g4884) & (key[15])) + ((g830) & (!g1914) & (!g2653) & (!g4883) & (g4884) & (!key[15])) + ((g830) & (!g1914) & (!g2653) & (!g4883) & (g4884) & (key[15])) + ((g830) & (!g1914) & (!g2653) & (g4883) & (g4884) & (!key[15])) + ((g830) & (!g1914) & (!g2653) & (g4883) & (g4884) & (key[15])) + ((g830) & (!g1914) & (g2653) & (!g4883) & (!g4884) & (!key[15])) + ((g830) & (!g1914) & (g2653) & (!g4883) & (!g4884) & (key[15])) + ((g830) & (!g1914) & (g2653) & (g4883) & (!g4884) & (!key[15])) + ((g830) & (!g1914) & (g2653) & (g4883) & (!g4884) & (key[15])) + ((g830) & (g1914) & (!g2653) & (g4883) & (!g4884) & (!key[15])) + ((g830) & (g1914) & (!g2653) & (g4883) & (!g4884) & (key[15])) + ((g830) & (g1914) & (!g2653) & (g4883) & (g4884) & (!key[15])) + ((g830) & (g1914) & (!g2653) & (g4883) & (g4884) & (key[15])) + ((g830) & (g1914) & (g2653) & (!g4883) & (!g4884) & (!key[15])) + ((g830) & (g1914) & (g2653) & (!g4883) & (!g4884) & (key[15])) + ((g830) & (g1914) & (g2653) & (!g4883) & (g4884) & (!key[15])) + ((g830) & (g1914) & (g2653) & (!g4883) & (g4884) & (key[15])));
	assign g4886 = (((!g2647) & (g3240)) + ((g2647) & (!g3240)));
	assign g4887 = (((!g2551) & (!g2598) & (g3155) & (g3196) & (g4758) & (g4886)) + ((!g2551) & (g2598) & (!g3155) & (g3196) & (!g4758) & (g4886)) + ((!g2551) & (g2598) & (!g3155) & (g3196) & (g4758) & (g4886)) + ((!g2551) & (g2598) & (g3155) & (!g3196) & (g4758) & (g4886)) + ((!g2551) & (g2598) & (g3155) & (g3196) & (!g4758) & (g4886)) + ((!g2551) & (g2598) & (g3155) & (g3196) & (g4758) & (g4886)) + ((g2551) & (!g2598) & (!g3155) & (g3196) & (g4758) & (g4886)) + ((g2551) & (!g2598) & (g3155) & (g3196) & (!g4758) & (g4886)) + ((g2551) & (!g2598) & (g3155) & (g3196) & (g4758) & (g4886)) + ((g2551) & (g2598) & (!g3155) & (!g3196) & (g4758) & (g4886)) + ((g2551) & (g2598) & (!g3155) & (g3196) & (!g4758) & (g4886)) + ((g2551) & (g2598) & (!g3155) & (g3196) & (g4758) & (g4886)) + ((g2551) & (g2598) & (g3155) & (!g3196) & (!g4758) & (g4886)) + ((g2551) & (g2598) & (g3155) & (!g3196) & (g4758) & (g4886)) + ((g2551) & (g2598) & (g3155) & (g3196) & (!g4758) & (g4886)) + ((g2551) & (g2598) & (g3155) & (g3196) & (g4758) & (g4886)));
	assign g4888 = (((g2647) & (g3240)));
	assign g4889 = (((g830) & (!g1914) & (!g4887) & (!g4888) & (!g5710) & (!g5711)) + ((g830) & (!g1914) & (!g4887) & (!g4888) & (!g5710) & (g5711)) + ((g830) & (!g1914) & (!g4887) & (g4888) & (g5710) & (!g5711)) + ((g830) & (!g1914) & (!g4887) & (g4888) & (g5710) & (g5711)) + ((g830) & (!g1914) & (g4887) & (!g4888) & (g5710) & (!g5711)) + ((g830) & (!g1914) & (g4887) & (!g4888) & (g5710) & (g5711)) + ((g830) & (!g1914) & (g4887) & (g4888) & (g5710) & (!g5711)) + ((g830) & (!g1914) & (g4887) & (g4888) & (g5710) & (g5711)) + ((g830) & (g1914) & (!g4887) & (!g4888) & (!g5710) & (g5711)) + ((g830) & (g1914) & (!g4887) & (!g4888) & (g5710) & (g5711)) + ((g830) & (g1914) & (!g4887) & (g4888) & (!g5710) & (g5711)) + ((g830) & (g1914) & (!g4887) & (g4888) & (g5710) & (g5711)) + ((g830) & (g1914) & (g4887) & (!g4888) & (!g5710) & (g5711)) + ((g830) & (g1914) & (g4887) & (!g4888) & (g5710) & (g5711)) + ((g830) & (g1914) & (g4887) & (g4888) & (!g5710) & (g5711)) + ((g830) & (g1914) & (g4887) & (g4888) & (g5710) & (g5711)));
	assign g4890 = (((!g1884) & (!g1977) & (!g1979) & (!g1908) & (!g2030) & (g2085)) + ((!g1884) & (!g1977) & (!g1979) & (!g1908) & (g2030) & (g2085)) + ((!g1884) & (!g1977) & (!g1979) & (g1908) & (!g2030) & (g2085)) + ((!g1884) & (!g1977) & (!g1979) & (g1908) & (g2030) & (g2085)) + ((!g1884) & (!g1977) & (g1979) & (!g1908) & (!g2030) & (!g2085)) + ((!g1884) & (!g1977) & (g1979) & (!g1908) & (g2030) & (!g2085)) + ((!g1884) & (!g1977) & (g1979) & (g1908) & (!g2030) & (!g2085)) + ((!g1884) & (!g1977) & (g1979) & (g1908) & (g2030) & (!g2085)) + ((!g1884) & (g1977) & (!g1979) & (!g1908) & (!g2030) & (g2085)) + ((!g1884) & (g1977) & (!g1979) & (!g1908) & (g2030) & (!g2085)) + ((!g1884) & (g1977) & (!g1979) & (g1908) & (!g2030) & (g2085)) + ((!g1884) & (g1977) & (!g1979) & (g1908) & (g2030) & (!g2085)) + ((!g1884) & (g1977) & (g1979) & (!g1908) & (!g2030) & (!g2085)) + ((!g1884) & (g1977) & (g1979) & (!g1908) & (g2030) & (g2085)) + ((!g1884) & (g1977) & (g1979) & (g1908) & (!g2030) & (!g2085)) + ((!g1884) & (g1977) & (g1979) & (g1908) & (g2030) & (g2085)) + ((g1884) & (!g1977) & (!g1979) & (!g1908) & (!g2030) & (g2085)) + ((g1884) & (!g1977) & (!g1979) & (!g1908) & (g2030) & (g2085)) + ((g1884) & (!g1977) & (!g1979) & (g1908) & (!g2030) & (g2085)) + ((g1884) & (!g1977) & (!g1979) & (g1908) & (g2030) & (!g2085)) + ((g1884) & (!g1977) & (g1979) & (!g1908) & (!g2030) & (!g2085)) + ((g1884) & (!g1977) & (g1979) & (!g1908) & (g2030) & (!g2085)) + ((g1884) & (!g1977) & (g1979) & (g1908) & (!g2030) & (!g2085)) + ((g1884) & (!g1977) & (g1979) & (g1908) & (g2030) & (g2085)) + ((g1884) & (g1977) & (!g1979) & (!g1908) & (!g2030) & (g2085)) + ((g1884) & (g1977) & (!g1979) & (!g1908) & (g2030) & (!g2085)) + ((g1884) & (g1977) & (!g1979) & (g1908) & (!g2030) & (!g2085)) + ((g1884) & (g1977) & (!g1979) & (g1908) & (g2030) & (!g2085)) + ((g1884) & (g1977) & (g1979) & (!g1908) & (!g2030) & (!g2085)) + ((g1884) & (g1977) & (g1979) & (!g1908) & (g2030) & (g2085)) + ((g1884) & (g1977) & (g1979) & (g1908) & (!g2030) & (g2085)) + ((g1884) & (g1977) & (g1979) & (g1908) & (g2030) & (g2085)));
	assign g4891 = (((!g1914) & (!g2320) & (!g2326) & (!g3673) & (!g4890)) + ((!g1914) & (!g2320) & (!g2326) & (!g3673) & (g4890)) + ((!g1914) & (!g2320) & (g2326) & (g3673) & (!g4890)) + ((!g1914) & (!g2320) & (g2326) & (g3673) & (g4890)) + ((!g1914) & (g2320) & (!g2326) & (g3673) & (!g4890)) + ((!g1914) & (g2320) & (!g2326) & (g3673) & (g4890)) + ((!g1914) & (g2320) & (g2326) & (!g3673) & (!g4890)) + ((!g1914) & (g2320) & (g2326) & (!g3673) & (g4890)) + ((g1914) & (!g2320) & (!g2326) & (!g3673) & (g4890)) + ((g1914) & (!g2320) & (!g2326) & (g3673) & (g4890)) + ((g1914) & (!g2320) & (g2326) & (!g3673) & (g4890)) + ((g1914) & (!g2320) & (g2326) & (g3673) & (g4890)) + ((g1914) & (g2320) & (!g2326) & (!g3673) & (g4890)) + ((g1914) & (g2320) & (!g2326) & (g3673) & (g4890)) + ((g1914) & (g2320) & (g2326) & (!g3673) & (g4890)) + ((g1914) & (g2320) & (g2326) & (g3673) & (g4890)));
	assign g8320 = (((!g5560) & (g5622) & (!g4892)) + ((!g5560) & (g5622) & (g4892)) + ((g5560) & (!g5622) & (g4892)) + ((g5560) & (g5622) & (g4892)));
	assign g4893 = (((!g830) & (!g2659) & (!g4891) & (g4892)) + ((!g830) & (!g2659) & (g4891) & (g4892)) + ((!g830) & (g2659) & (!g4891) & (g4892)) + ((!g830) & (g2659) & (g4891) & (g4892)) + ((g830) & (!g2659) & (g4891) & (!g4892)) + ((g830) & (!g2659) & (g4891) & (g4892)) + ((g830) & (g2659) & (!g4891) & (!g4892)) + ((g830) & (g2659) & (!g4891) & (g4892)));
	assign g4894 = (((!g2311) & (!g2323) & (!g3782)) + ((!g2311) & (g2323) & (g3782)) + ((g2311) & (!g2323) & (g3782)) + ((g2311) & (g2323) & (!g3782)));
	assign g4895 = (((!g1906) & (!g1940) & (!g1942) & (!g1910) & (!g2038) & (g2088)) + ((!g1906) & (!g1940) & (!g1942) & (!g1910) & (g2038) & (g2088)) + ((!g1906) & (!g1940) & (!g1942) & (g1910) & (!g2038) & (g2088)) + ((!g1906) & (!g1940) & (!g1942) & (g1910) & (g2038) & (g2088)) + ((!g1906) & (!g1940) & (g1942) & (!g1910) & (!g2038) & (!g2088)) + ((!g1906) & (!g1940) & (g1942) & (!g1910) & (g2038) & (!g2088)) + ((!g1906) & (!g1940) & (g1942) & (g1910) & (!g2038) & (!g2088)) + ((!g1906) & (!g1940) & (g1942) & (g1910) & (g2038) & (!g2088)) + ((!g1906) & (g1940) & (!g1942) & (!g1910) & (!g2038) & (g2088)) + ((!g1906) & (g1940) & (!g1942) & (!g1910) & (g2038) & (!g2088)) + ((!g1906) & (g1940) & (!g1942) & (g1910) & (!g2038) & (g2088)) + ((!g1906) & (g1940) & (!g1942) & (g1910) & (g2038) & (!g2088)) + ((!g1906) & (g1940) & (g1942) & (!g1910) & (!g2038) & (!g2088)) + ((!g1906) & (g1940) & (g1942) & (!g1910) & (g2038) & (g2088)) + ((!g1906) & (g1940) & (g1942) & (g1910) & (!g2038) & (!g2088)) + ((!g1906) & (g1940) & (g1942) & (g1910) & (g2038) & (g2088)) + ((g1906) & (!g1940) & (!g1942) & (!g1910) & (!g2038) & (g2088)) + ((g1906) & (!g1940) & (!g1942) & (!g1910) & (g2038) & (g2088)) + ((g1906) & (!g1940) & (!g1942) & (g1910) & (!g2038) & (g2088)) + ((g1906) & (!g1940) & (!g1942) & (g1910) & (g2038) & (!g2088)) + ((g1906) & (!g1940) & (g1942) & (!g1910) & (!g2038) & (!g2088)) + ((g1906) & (!g1940) & (g1942) & (!g1910) & (g2038) & (!g2088)) + ((g1906) & (!g1940) & (g1942) & (g1910) & (!g2038) & (!g2088)) + ((g1906) & (!g1940) & (g1942) & (g1910) & (g2038) & (g2088)) + ((g1906) & (g1940) & (!g1942) & (!g1910) & (!g2038) & (g2088)) + ((g1906) & (g1940) & (!g1942) & (!g1910) & (g2038) & (!g2088)) + ((g1906) & (g1940) & (!g1942) & (g1910) & (!g2038) & (!g2088)) + ((g1906) & (g1940) & (!g1942) & (g1910) & (g2038) & (!g2088)) + ((g1906) & (g1940) & (g1942) & (!g1910) & (!g2038) & (!g2088)) + ((g1906) & (g1940) & (g1942) & (!g1910) & (g2038) & (g2088)) + ((g1906) & (g1940) & (g1942) & (g1910) & (!g2038) & (g2088)) + ((g1906) & (g1940) & (g1942) & (g1910) & (g2038) & (g2088)));
	assign g4896 = (((!g830) & (!g1914) & (!g2661) & (!g4894) & (!g4895) & (key[143])) + ((!g830) & (!g1914) & (!g2661) & (!g4894) & (g4895) & (key[143])) + ((!g830) & (!g1914) & (!g2661) & (g4894) & (!g4895) & (key[143])) + ((!g830) & (!g1914) & (!g2661) & (g4894) & (g4895) & (key[143])) + ((!g830) & (!g1914) & (g2661) & (!g4894) & (!g4895) & (key[143])) + ((!g830) & (!g1914) & (g2661) & (!g4894) & (g4895) & (key[143])) + ((!g830) & (!g1914) & (g2661) & (g4894) & (!g4895) & (key[143])) + ((!g830) & (!g1914) & (g2661) & (g4894) & (g4895) & (key[143])) + ((!g830) & (g1914) & (!g2661) & (!g4894) & (!g4895) & (key[143])) + ((!g830) & (g1914) & (!g2661) & (!g4894) & (g4895) & (key[143])) + ((!g830) & (g1914) & (!g2661) & (g4894) & (!g4895) & (key[143])) + ((!g830) & (g1914) & (!g2661) & (g4894) & (g4895) & (key[143])) + ((!g830) & (g1914) & (g2661) & (!g4894) & (!g4895) & (key[143])) + ((!g830) & (g1914) & (g2661) & (!g4894) & (g4895) & (key[143])) + ((!g830) & (g1914) & (g2661) & (g4894) & (!g4895) & (key[143])) + ((!g830) & (g1914) & (g2661) & (g4894) & (g4895) & (key[143])) + ((g830) & (!g1914) & (!g2661) & (!g4894) & (g4895) & (!key[143])) + ((g830) & (!g1914) & (!g2661) & (!g4894) & (g4895) & (key[143])) + ((g830) & (!g1914) & (!g2661) & (g4894) & (g4895) & (!key[143])) + ((g830) & (!g1914) & (!g2661) & (g4894) & (g4895) & (key[143])) + ((g830) & (!g1914) & (g2661) & (!g4894) & (!g4895) & (!key[143])) + ((g830) & (!g1914) & (g2661) & (!g4894) & (!g4895) & (key[143])) + ((g830) & (!g1914) & (g2661) & (g4894) & (!g4895) & (!key[143])) + ((g830) & (!g1914) & (g2661) & (g4894) & (!g4895) & (key[143])) + ((g830) & (g1914) & (!g2661) & (g4894) & (!g4895) & (!key[143])) + ((g830) & (g1914) & (!g2661) & (g4894) & (!g4895) & (key[143])) + ((g830) & (g1914) & (!g2661) & (g4894) & (g4895) & (!key[143])) + ((g830) & (g1914) & (!g2661) & (g4894) & (g4895) & (key[143])) + ((g830) & (g1914) & (g2661) & (!g4894) & (!g4895) & (!key[143])) + ((g830) & (g1914) & (g2661) & (!g4894) & (!g4895) & (key[143])) + ((g830) & (g1914) & (g2661) & (!g4894) & (g4895) & (!key[143])) + ((g830) & (g1914) & (g2661) & (!g4894) & (g4895) & (key[143])));
	assign g4897 = (((!g1894) & (!g1910) & (!g2034) & (!g2038) & (!g2065) & (g2088)) + ((!g1894) & (!g1910) & (!g2034) & (!g2038) & (g2065) & (!g2088)) + ((!g1894) & (!g1910) & (!g2034) & (g2038) & (!g2065) & (g2088)) + ((!g1894) & (!g1910) & (!g2034) & (g2038) & (g2065) & (!g2088)) + ((!g1894) & (!g1910) & (g2034) & (!g2038) & (!g2065) & (g2088)) + ((!g1894) & (!g1910) & (g2034) & (!g2038) & (g2065) & (!g2088)) + ((!g1894) & (!g1910) & (g2034) & (g2038) & (!g2065) & (!g2088)) + ((!g1894) & (!g1910) & (g2034) & (g2038) & (g2065) & (g2088)) + ((!g1894) & (g1910) & (!g2034) & (!g2038) & (!g2065) & (g2088)) + ((!g1894) & (g1910) & (!g2034) & (!g2038) & (g2065) & (!g2088)) + ((!g1894) & (g1910) & (!g2034) & (g2038) & (!g2065) & (g2088)) + ((!g1894) & (g1910) & (!g2034) & (g2038) & (g2065) & (!g2088)) + ((!g1894) & (g1910) & (g2034) & (!g2038) & (!g2065) & (g2088)) + ((!g1894) & (g1910) & (g2034) & (!g2038) & (g2065) & (!g2088)) + ((!g1894) & (g1910) & (g2034) & (g2038) & (!g2065) & (!g2088)) + ((!g1894) & (g1910) & (g2034) & (g2038) & (g2065) & (g2088)) + ((g1894) & (!g1910) & (!g2034) & (!g2038) & (!g2065) & (g2088)) + ((g1894) & (!g1910) & (!g2034) & (!g2038) & (g2065) & (!g2088)) + ((g1894) & (!g1910) & (!g2034) & (g2038) & (!g2065) & (g2088)) + ((g1894) & (!g1910) & (!g2034) & (g2038) & (g2065) & (!g2088)) + ((g1894) & (!g1910) & (g2034) & (!g2038) & (!g2065) & (g2088)) + ((g1894) & (!g1910) & (g2034) & (!g2038) & (g2065) & (!g2088)) + ((g1894) & (!g1910) & (g2034) & (g2038) & (!g2065) & (!g2088)) + ((g1894) & (!g1910) & (g2034) & (g2038) & (g2065) & (g2088)) + ((g1894) & (g1910) & (!g2034) & (!g2038) & (!g2065) & (g2088)) + ((g1894) & (g1910) & (!g2034) & (!g2038) & (g2065) & (!g2088)) + ((g1894) & (g1910) & (!g2034) & (g2038) & (!g2065) & (!g2088)) + ((g1894) & (g1910) & (!g2034) & (g2038) & (g2065) & (g2088)) + ((g1894) & (g1910) & (g2034) & (!g2038) & (!g2065) & (!g2088)) + ((g1894) & (g1910) & (g2034) & (!g2038) & (g2065) & (g2088)) + ((g1894) & (g1910) & (g2034) & (g2038) & (!g2065) & (!g2088)) + ((g1894) & (g1910) & (g2034) & (g2038) & (g2065) & (g2088)));
	assign g4898 = (((!g1997) & (!g1098) & (!g3448)) + ((!g1997) & (g1098) & (g3448)) + ((g1997) & (!g1098) & (g3448)) + ((g1997) & (g1098) & (!g3448)));
	assign g4899 = (((!g830) & (!g1914) & (!g2663) & (!g4897) & (!g4898) & (key[111])) + ((!g830) & (!g1914) & (!g2663) & (!g4897) & (g4898) & (key[111])) + ((!g830) & (!g1914) & (!g2663) & (g4897) & (!g4898) & (key[111])) + ((!g830) & (!g1914) & (!g2663) & (g4897) & (g4898) & (key[111])) + ((!g830) & (!g1914) & (g2663) & (!g4897) & (!g4898) & (key[111])) + ((!g830) & (!g1914) & (g2663) & (!g4897) & (g4898) & (key[111])) + ((!g830) & (!g1914) & (g2663) & (g4897) & (!g4898) & (key[111])) + ((!g830) & (!g1914) & (g2663) & (g4897) & (g4898) & (key[111])) + ((!g830) & (g1914) & (!g2663) & (!g4897) & (!g4898) & (key[111])) + ((!g830) & (g1914) & (!g2663) & (!g4897) & (g4898) & (key[111])) + ((!g830) & (g1914) & (!g2663) & (g4897) & (!g4898) & (key[111])) + ((!g830) & (g1914) & (!g2663) & (g4897) & (g4898) & (key[111])) + ((!g830) & (g1914) & (g2663) & (!g4897) & (!g4898) & (key[111])) + ((!g830) & (g1914) & (g2663) & (!g4897) & (g4898) & (key[111])) + ((!g830) & (g1914) & (g2663) & (g4897) & (!g4898) & (key[111])) + ((!g830) & (g1914) & (g2663) & (g4897) & (g4898) & (key[111])) + ((g830) & (!g1914) & (!g2663) & (!g4897) & (g4898) & (!key[111])) + ((g830) & (!g1914) & (!g2663) & (!g4897) & (g4898) & (key[111])) + ((g830) & (!g1914) & (!g2663) & (g4897) & (g4898) & (!key[111])) + ((g830) & (!g1914) & (!g2663) & (g4897) & (g4898) & (key[111])) + ((g830) & (!g1914) & (g2663) & (!g4897) & (!g4898) & (!key[111])) + ((g830) & (!g1914) & (g2663) & (!g4897) & (!g4898) & (key[111])) + ((g830) & (!g1914) & (g2663) & (g4897) & (!g4898) & (!key[111])) + ((g830) & (!g1914) & (g2663) & (g4897) & (!g4898) & (key[111])) + ((g830) & (g1914) & (!g2663) & (g4897) & (!g4898) & (!key[111])) + ((g830) & (g1914) & (!g2663) & (g4897) & (!g4898) & (key[111])) + ((g830) & (g1914) & (!g2663) & (g4897) & (g4898) & (!key[111])) + ((g830) & (g1914) & (!g2663) & (g4897) & (g4898) & (key[111])) + ((g830) & (g1914) & (g2663) & (!g4897) & (!g4898) & (!key[111])) + ((g830) & (g1914) & (g2663) & (!g4897) & (!g4898) & (key[111])) + ((g830) & (g1914) & (g2663) & (!g4897) & (g4898) & (!key[111])) + ((g830) & (g1914) & (g2663) & (!g4897) & (g4898) & (key[111])));
	assign g4900 = (((!g2304) & (!g3559) & (!g2326)) + ((!g2304) & (g3559) & (g2326)) + ((g2304) & (!g3559) & (g2326)) + ((g2304) & (g3559) & (!g2326)));
	assign g4901 = (((!g1890) & (!g1939) & (!g1941) & (!g1896) & (!g2041) & (g2068)) + ((!g1890) & (!g1939) & (!g1941) & (!g1896) & (g2041) & (g2068)) + ((!g1890) & (!g1939) & (!g1941) & (g1896) & (!g2041) & (g2068)) + ((!g1890) & (!g1939) & (!g1941) & (g1896) & (g2041) & (g2068)) + ((!g1890) & (!g1939) & (g1941) & (!g1896) & (!g2041) & (!g2068)) + ((!g1890) & (!g1939) & (g1941) & (!g1896) & (g2041) & (!g2068)) + ((!g1890) & (!g1939) & (g1941) & (g1896) & (!g2041) & (!g2068)) + ((!g1890) & (!g1939) & (g1941) & (g1896) & (g2041) & (!g2068)) + ((!g1890) & (g1939) & (!g1941) & (!g1896) & (!g2041) & (g2068)) + ((!g1890) & (g1939) & (!g1941) & (!g1896) & (g2041) & (!g2068)) + ((!g1890) & (g1939) & (!g1941) & (g1896) & (!g2041) & (g2068)) + ((!g1890) & (g1939) & (!g1941) & (g1896) & (g2041) & (!g2068)) + ((!g1890) & (g1939) & (g1941) & (!g1896) & (!g2041) & (!g2068)) + ((!g1890) & (g1939) & (g1941) & (!g1896) & (g2041) & (g2068)) + ((!g1890) & (g1939) & (g1941) & (g1896) & (!g2041) & (!g2068)) + ((!g1890) & (g1939) & (g1941) & (g1896) & (g2041) & (g2068)) + ((g1890) & (!g1939) & (!g1941) & (!g1896) & (!g2041) & (g2068)) + ((g1890) & (!g1939) & (!g1941) & (!g1896) & (g2041) & (g2068)) + ((g1890) & (!g1939) & (!g1941) & (g1896) & (!g2041) & (g2068)) + ((g1890) & (!g1939) & (!g1941) & (g1896) & (g2041) & (!g2068)) + ((g1890) & (!g1939) & (g1941) & (!g1896) & (!g2041) & (!g2068)) + ((g1890) & (!g1939) & (g1941) & (!g1896) & (g2041) & (!g2068)) + ((g1890) & (!g1939) & (g1941) & (g1896) & (!g2041) & (!g2068)) + ((g1890) & (!g1939) & (g1941) & (g1896) & (g2041) & (g2068)) + ((g1890) & (g1939) & (!g1941) & (!g1896) & (!g2041) & (g2068)) + ((g1890) & (g1939) & (!g1941) & (!g1896) & (g2041) & (!g2068)) + ((g1890) & (g1939) & (!g1941) & (g1896) & (!g2041) & (!g2068)) + ((g1890) & (g1939) & (!g1941) & (g1896) & (g2041) & (!g2068)) + ((g1890) & (g1939) & (g1941) & (!g1896) & (!g2041) & (!g2068)) + ((g1890) & (g1939) & (g1941) & (!g1896) & (g2041) & (g2068)) + ((g1890) & (g1939) & (g1941) & (g1896) & (!g2041) & (g2068)) + ((g1890) & (g1939) & (g1941) & (g1896) & (g2041) & (g2068)));
	assign g4902 = (((!g830) & (!g1914) & (!g2665) & (!g4900) & (!g4901) & (nonce[15])) + ((!g830) & (!g1914) & (!g2665) & (!g4900) & (g4901) & (nonce[15])) + ((!g830) & (!g1914) & (!g2665) & (g4900) & (!g4901) & (nonce[15])) + ((!g830) & (!g1914) & (!g2665) & (g4900) & (g4901) & (nonce[15])) + ((!g830) & (!g1914) & (g2665) & (!g4900) & (!g4901) & (nonce[15])) + ((!g830) & (!g1914) & (g2665) & (!g4900) & (g4901) & (nonce[15])) + ((!g830) & (!g1914) & (g2665) & (g4900) & (!g4901) & (nonce[15])) + ((!g830) & (!g1914) & (g2665) & (g4900) & (g4901) & (nonce[15])) + ((!g830) & (g1914) & (!g2665) & (!g4900) & (!g4901) & (nonce[15])) + ((!g830) & (g1914) & (!g2665) & (!g4900) & (g4901) & (nonce[15])) + ((!g830) & (g1914) & (!g2665) & (g4900) & (!g4901) & (nonce[15])) + ((!g830) & (g1914) & (!g2665) & (g4900) & (g4901) & (nonce[15])) + ((!g830) & (g1914) & (g2665) & (!g4900) & (!g4901) & (nonce[15])) + ((!g830) & (g1914) & (g2665) & (!g4900) & (g4901) & (nonce[15])) + ((!g830) & (g1914) & (g2665) & (g4900) & (!g4901) & (nonce[15])) + ((!g830) & (g1914) & (g2665) & (g4900) & (g4901) & (nonce[15])) + ((g830) & (!g1914) & (!g2665) & (!g4900) & (g4901) & (!nonce[15])) + ((g830) & (!g1914) & (!g2665) & (!g4900) & (g4901) & (nonce[15])) + ((g830) & (!g1914) & (!g2665) & (g4900) & (g4901) & (!nonce[15])) + ((g830) & (!g1914) & (!g2665) & (g4900) & (g4901) & (nonce[15])) + ((g830) & (!g1914) & (g2665) & (!g4900) & (!g4901) & (!nonce[15])) + ((g830) & (!g1914) & (g2665) & (!g4900) & (!g4901) & (nonce[15])) + ((g830) & (!g1914) & (g2665) & (g4900) & (!g4901) & (!nonce[15])) + ((g830) & (!g1914) & (g2665) & (g4900) & (!g4901) & (nonce[15])) + ((g830) & (g1914) & (!g2665) & (g4900) & (!g4901) & (!nonce[15])) + ((g830) & (g1914) & (!g2665) & (g4900) & (!g4901) & (nonce[15])) + ((g830) & (g1914) & (!g2665) & (g4900) & (g4901) & (!nonce[15])) + ((g830) & (g1914) & (!g2665) & (g4900) & (g4901) & (nonce[15])) + ((g830) & (g1914) & (g2665) & (!g4900) & (!g4901) & (!nonce[15])) + ((g830) & (g1914) & (g2665) & (!g4900) & (!g4901) & (nonce[15])) + ((g830) & (g1914) & (g2665) & (!g4900) & (g4901) & (!nonce[15])) + ((g830) & (g1914) & (g2665) & (!g4900) & (g4901) & (nonce[15])));
	assign g4903 = (((!g3250) & (g3265)) + ((g3250) & (!g3265)));
	assign g4904 = (((!g3159) & (!g3177) & (g3165) & (g3210) & (g4764) & (g4903)) + ((!g3159) & (g3177) & (!g3165) & (g3210) & (!g4764) & (g4903)) + ((!g3159) & (g3177) & (!g3165) & (g3210) & (g4764) & (g4903)) + ((!g3159) & (g3177) & (g3165) & (!g3210) & (g4764) & (g4903)) + ((!g3159) & (g3177) & (g3165) & (g3210) & (!g4764) & (g4903)) + ((!g3159) & (g3177) & (g3165) & (g3210) & (g4764) & (g4903)) + ((g3159) & (!g3177) & (!g3165) & (g3210) & (g4764) & (g4903)) + ((g3159) & (!g3177) & (g3165) & (g3210) & (!g4764) & (g4903)) + ((g3159) & (!g3177) & (g3165) & (g3210) & (g4764) & (g4903)) + ((g3159) & (g3177) & (!g3165) & (!g3210) & (g4764) & (g4903)) + ((g3159) & (g3177) & (!g3165) & (g3210) & (!g4764) & (g4903)) + ((g3159) & (g3177) & (!g3165) & (g3210) & (g4764) & (g4903)) + ((g3159) & (g3177) & (g3165) & (!g3210) & (!g4764) & (g4903)) + ((g3159) & (g3177) & (g3165) & (!g3210) & (g4764) & (g4903)) + ((g3159) & (g3177) & (g3165) & (g3210) & (!g4764) & (g4903)) + ((g3159) & (g3177) & (g3165) & (g3210) & (g4764) & (g4903)));
	assign g4905 = (((g3250) & (g3265)));
	assign g4906 = (((g830) & (!g1914) & (!g4904) & (!g4905) & (!g5712) & (!g5713)) + ((g830) & (!g1914) & (!g4904) & (!g4905) & (!g5712) & (g5713)) + ((g830) & (!g1914) & (!g4904) & (g4905) & (g5712) & (!g5713)) + ((g830) & (!g1914) & (!g4904) & (g4905) & (g5712) & (g5713)) + ((g830) & (!g1914) & (g4904) & (!g4905) & (g5712) & (!g5713)) + ((g830) & (!g1914) & (g4904) & (!g4905) & (g5712) & (g5713)) + ((g830) & (!g1914) & (g4904) & (g4905) & (g5712) & (!g5713)) + ((g830) & (!g1914) & (g4904) & (g4905) & (g5712) & (g5713)) + ((g830) & (g1914) & (!g4904) & (!g4905) & (!g5712) & (g5713)) + ((g830) & (g1914) & (!g4904) & (!g4905) & (g5712) & (g5713)) + ((g830) & (g1914) & (!g4904) & (g4905) & (!g5712) & (g5713)) + ((g830) & (g1914) & (!g4904) & (g4905) & (g5712) & (g5713)) + ((g830) & (g1914) & (g4904) & (!g4905) & (!g5712) & (g5713)) + ((g830) & (g1914) & (g4904) & (!g4905) & (g5712) & (g5713)) + ((g830) & (g1914) & (g4904) & (g4905) & (!g5712) & (g5713)) + ((g830) & (g1914) & (g4904) & (g4905) & (g5712) & (g5713)));
	assign g4907 = (((!g3813) & (!g3814)));
	assign g4908 = (((g1914) & (!g2227) & (!g2239) & (!g4907)) + ((g1914) & (!g2227) & (g2239) & (g4907)) + ((g1914) & (g2227) & (!g2239) & (g4907)) + ((g1914) & (g2227) & (g2239) & (!g4907)));
	assign g4909 = (((!g3830) & (!g3831)));
	assign g4910 = (((!g1914) & (!g1954) & (!g2253) & (!g4909)) + ((!g1914) & (!g1954) & (g2253) & (g4909)) + ((!g1914) & (g1954) & (!g2253) & (g4909)) + ((!g1914) & (g1954) & (g2253) & (!g4909)));
	assign g4911 = (((!g830) & (!g2669) & (!g4908) & (!g4910) & (nonce[47])) + ((!g830) & (!g2669) & (!g4908) & (g4910) & (nonce[47])) + ((!g830) & (!g2669) & (g4908) & (!g4910) & (nonce[47])) + ((!g830) & (!g2669) & (g4908) & (g4910) & (nonce[47])) + ((!g830) & (g2669) & (!g4908) & (!g4910) & (nonce[47])) + ((!g830) & (g2669) & (!g4908) & (g4910) & (nonce[47])) + ((!g830) & (g2669) & (g4908) & (!g4910) & (nonce[47])) + ((!g830) & (g2669) & (g4908) & (g4910) & (nonce[47])) + ((g830) & (!g2669) & (!g4908) & (g4910) & (!nonce[47])) + ((g830) & (!g2669) & (!g4908) & (g4910) & (nonce[47])) + ((g830) & (!g2669) & (g4908) & (!g4910) & (!nonce[47])) + ((g830) & (!g2669) & (g4908) & (!g4910) & (nonce[47])) + ((g830) & (!g2669) & (g4908) & (g4910) & (!nonce[47])) + ((g830) & (!g2669) & (g4908) & (g4910) & (nonce[47])) + ((g830) & (g2669) & (!g4908) & (!g4910) & (!nonce[47])) + ((g830) & (g2669) & (!g4908) & (!g4910) & (nonce[47])));
	assign g4912 = (((!g1888) & (!g1978) & (!g1980) & (!g1904) & (!g2043) & (g2080)) + ((!g1888) & (!g1978) & (!g1980) & (!g1904) & (g2043) & (g2080)) + ((!g1888) & (!g1978) & (!g1980) & (g1904) & (!g2043) & (g2080)) + ((!g1888) & (!g1978) & (!g1980) & (g1904) & (g2043) & (g2080)) + ((!g1888) & (!g1978) & (g1980) & (!g1904) & (!g2043) & (!g2080)) + ((!g1888) & (!g1978) & (g1980) & (!g1904) & (g2043) & (!g2080)) + ((!g1888) & (!g1978) & (g1980) & (g1904) & (!g2043) & (!g2080)) + ((!g1888) & (!g1978) & (g1980) & (g1904) & (g2043) & (!g2080)) + ((!g1888) & (g1978) & (!g1980) & (!g1904) & (!g2043) & (g2080)) + ((!g1888) & (g1978) & (!g1980) & (!g1904) & (g2043) & (!g2080)) + ((!g1888) & (g1978) & (!g1980) & (g1904) & (!g2043) & (g2080)) + ((!g1888) & (g1978) & (!g1980) & (g1904) & (g2043) & (!g2080)) + ((!g1888) & (g1978) & (g1980) & (!g1904) & (!g2043) & (!g2080)) + ((!g1888) & (g1978) & (g1980) & (!g1904) & (g2043) & (g2080)) + ((!g1888) & (g1978) & (g1980) & (g1904) & (!g2043) & (!g2080)) + ((!g1888) & (g1978) & (g1980) & (g1904) & (g2043) & (g2080)) + ((g1888) & (!g1978) & (!g1980) & (!g1904) & (!g2043) & (g2080)) + ((g1888) & (!g1978) & (!g1980) & (!g1904) & (g2043) & (g2080)) + ((g1888) & (!g1978) & (!g1980) & (g1904) & (!g2043) & (g2080)) + ((g1888) & (!g1978) & (!g1980) & (g1904) & (g2043) & (!g2080)) + ((g1888) & (!g1978) & (g1980) & (!g1904) & (!g2043) & (!g2080)) + ((g1888) & (!g1978) & (g1980) & (!g1904) & (g2043) & (!g2080)) + ((g1888) & (!g1978) & (g1980) & (g1904) & (!g2043) & (!g2080)) + ((g1888) & (!g1978) & (g1980) & (g1904) & (g2043) & (g2080)) + ((g1888) & (g1978) & (!g1980) & (!g1904) & (!g2043) & (g2080)) + ((g1888) & (g1978) & (!g1980) & (!g1904) & (g2043) & (!g2080)) + ((g1888) & (g1978) & (!g1980) & (g1904) & (!g2043) & (!g2080)) + ((g1888) & (g1978) & (!g1980) & (g1904) & (g2043) & (!g2080)) + ((g1888) & (g1978) & (g1980) & (!g1904) & (!g2043) & (!g2080)) + ((g1888) & (g1978) & (g1980) & (!g1904) & (g2043) & (g2080)) + ((g1888) & (g1978) & (g1980) & (g1904) & (!g2043) & (g2080)) + ((g1888) & (g1978) & (g1980) & (g1904) & (g2043) & (g2080)));
	assign g4913 = (((!g2311) & (!g2314) & (!g3606)) + ((!g2311) & (g2314) & (g3606)) + ((g2311) & (!g2314) & (g3606)) + ((g2311) & (g2314) & (!g3606)));
	assign g4914 = (((!g830) & (!g1914) & (!g2672) & (!g4912) & (!g4913) & (key[239])) + ((!g830) & (!g1914) & (!g2672) & (!g4912) & (g4913) & (key[239])) + ((!g830) & (!g1914) & (!g2672) & (g4912) & (!g4913) & (key[239])) + ((!g830) & (!g1914) & (!g2672) & (g4912) & (g4913) & (key[239])) + ((!g830) & (!g1914) & (g2672) & (!g4912) & (!g4913) & (key[239])) + ((!g830) & (!g1914) & (g2672) & (!g4912) & (g4913) & (key[239])) + ((!g830) & (!g1914) & (g2672) & (g4912) & (!g4913) & (key[239])) + ((!g830) & (!g1914) & (g2672) & (g4912) & (g4913) & (key[239])) + ((!g830) & (g1914) & (!g2672) & (!g4912) & (!g4913) & (key[239])) + ((!g830) & (g1914) & (!g2672) & (!g4912) & (g4913) & (key[239])) + ((!g830) & (g1914) & (!g2672) & (g4912) & (!g4913) & (key[239])) + ((!g830) & (g1914) & (!g2672) & (g4912) & (g4913) & (key[239])) + ((!g830) & (g1914) & (g2672) & (!g4912) & (!g4913) & (key[239])) + ((!g830) & (g1914) & (g2672) & (!g4912) & (g4913) & (key[239])) + ((!g830) & (g1914) & (g2672) & (g4912) & (!g4913) & (key[239])) + ((!g830) & (g1914) & (g2672) & (g4912) & (g4913) & (key[239])) + ((g830) & (!g1914) & (!g2672) & (!g4912) & (g4913) & (!key[239])) + ((g830) & (!g1914) & (!g2672) & (!g4912) & (g4913) & (key[239])) + ((g830) & (!g1914) & (!g2672) & (g4912) & (g4913) & (!key[239])) + ((g830) & (!g1914) & (!g2672) & (g4912) & (g4913) & (key[239])) + ((g830) & (!g1914) & (g2672) & (!g4912) & (!g4913) & (!key[239])) + ((g830) & (!g1914) & (g2672) & (!g4912) & (!g4913) & (key[239])) + ((g830) & (!g1914) & (g2672) & (g4912) & (!g4913) & (!key[239])) + ((g830) & (!g1914) & (g2672) & (g4912) & (!g4913) & (key[239])) + ((g830) & (g1914) & (!g2672) & (g4912) & (!g4913) & (!key[239])) + ((g830) & (g1914) & (!g2672) & (g4912) & (!g4913) & (key[239])) + ((g830) & (g1914) & (!g2672) & (g4912) & (g4913) & (!key[239])) + ((g830) & (g1914) & (!g2672) & (g4912) & (g4913) & (key[239])) + ((g830) & (g1914) & (g2672) & (!g4912) & (!g4913) & (!key[239])) + ((g830) & (g1914) & (g2672) & (!g4912) & (!g4913) & (key[239])) + ((g830) & (g1914) & (g2672) & (!g4912) & (g4913) & (!key[239])) + ((g830) & (g1914) & (g2672) & (!g4912) & (g4913) & (key[239])));
	assign g4915 = (((!g3712) & (!g3713)));
	assign g4916 = (((g1914) & (!g1992) & (!g2253) & (!g4915)) + ((g1914) & (!g1992) & (g2253) & (g4915)) + ((g1914) & (g1992) & (!g2253) & (g4915)) + ((g1914) & (g1992) & (g2253) & (!g4915)));
	assign g4917 = (((!g3729) & (!g3730)));
	assign g4918 = (((!g1914) & (!g2236) & (!g2239) & (!g4917)) + ((!g1914) & (!g2236) & (g2239) & (g4917)) + ((!g1914) & (g2236) & (!g2239) & (g4917)) + ((!g1914) & (g2236) & (g2239) & (!g4917)));
	assign g4919 = (((!g830) & (!g2674) & (!g4916) & (!g4918) & (key[207])) + ((!g830) & (!g2674) & (!g4916) & (g4918) & (key[207])) + ((!g830) & (!g2674) & (g4916) & (!g4918) & (key[207])) + ((!g830) & (!g2674) & (g4916) & (g4918) & (key[207])) + ((!g830) & (g2674) & (!g4916) & (!g4918) & (key[207])) + ((!g830) & (g2674) & (!g4916) & (g4918) & (key[207])) + ((!g830) & (g2674) & (g4916) & (!g4918) & (key[207])) + ((!g830) & (g2674) & (g4916) & (g4918) & (key[207])) + ((g830) & (!g2674) & (!g4916) & (g4918) & (!key[207])) + ((g830) & (!g2674) & (!g4916) & (g4918) & (key[207])) + ((g830) & (!g2674) & (g4916) & (!g4918) & (!key[207])) + ((g830) & (!g2674) & (g4916) & (!g4918) & (key[207])) + ((g830) & (!g2674) & (g4916) & (g4918) & (!key[207])) + ((g830) & (!g2674) & (g4916) & (g4918) & (key[207])) + ((g830) & (g2674) & (!g4916) & (!g4918) & (!key[207])) + ((g830) & (g2674) & (!g4916) & (!g4918) & (key[207])));
	assign g4920 = (((!g3274) & (g3279)) + ((g3274) & (!g3279)));
	assign g4921 = (((!g3168) & (!g3190) & (g3170) & (g3202) & (g4775) & (g4920)) + ((!g3168) & (g3190) & (!g3170) & (g3202) & (!g4775) & (g4920)) + ((!g3168) & (g3190) & (!g3170) & (g3202) & (g4775) & (g4920)) + ((!g3168) & (g3190) & (g3170) & (!g3202) & (g4775) & (g4920)) + ((!g3168) & (g3190) & (g3170) & (g3202) & (!g4775) & (g4920)) + ((!g3168) & (g3190) & (g3170) & (g3202) & (g4775) & (g4920)) + ((g3168) & (!g3190) & (!g3170) & (g3202) & (g4775) & (g4920)) + ((g3168) & (!g3190) & (g3170) & (g3202) & (!g4775) & (g4920)) + ((g3168) & (!g3190) & (g3170) & (g3202) & (g4775) & (g4920)) + ((g3168) & (g3190) & (!g3170) & (!g3202) & (g4775) & (g4920)) + ((g3168) & (g3190) & (!g3170) & (g3202) & (!g4775) & (g4920)) + ((g3168) & (g3190) & (!g3170) & (g3202) & (g4775) & (g4920)) + ((g3168) & (g3190) & (g3170) & (!g3202) & (!g4775) & (g4920)) + ((g3168) & (g3190) & (g3170) & (!g3202) & (g4775) & (g4920)) + ((g3168) & (g3190) & (g3170) & (g3202) & (!g4775) & (g4920)) + ((g3168) & (g3190) & (g3170) & (g3202) & (g4775) & (g4920)));
	assign g4922 = (((g3274) & (g3279)));
	assign g4923 = (((g830) & (!g1914) & (!g4921) & (!g4922) & (!g5714) & (!g5715)) + ((g830) & (!g1914) & (!g4921) & (!g4922) & (!g5714) & (g5715)) + ((g830) & (!g1914) & (!g4921) & (g4922) & (g5714) & (!g5715)) + ((g830) & (!g1914) & (!g4921) & (g4922) & (g5714) & (g5715)) + ((g830) & (!g1914) & (g4921) & (!g4922) & (g5714) & (!g5715)) + ((g830) & (!g1914) & (g4921) & (!g4922) & (g5714) & (g5715)) + ((g830) & (!g1914) & (g4921) & (g4922) & (g5714) & (!g5715)) + ((g830) & (!g1914) & (g4921) & (g4922) & (g5714) & (g5715)) + ((g830) & (g1914) & (!g4921) & (!g4922) & (!g5714) & (g5715)) + ((g830) & (g1914) & (!g4921) & (!g4922) & (g5714) & (g5715)) + ((g830) & (g1914) & (!g4921) & (g4922) & (!g5714) & (g5715)) + ((g830) & (g1914) & (!g4921) & (g4922) & (g5714) & (g5715)) + ((g830) & (g1914) & (g4921) & (!g4922) & (!g5714) & (g5715)) + ((g830) & (g1914) & (g4921) & (!g4922) & (g5714) & (g5715)) + ((g830) & (g1914) & (g4921) & (g4922) & (!g5714) & (g5715)) + ((g830) & (g1914) & (g4921) & (g4922) & (g5714) & (g5715)));
	assign g4924 = (((!g1473) & (!g1507) & (!g4864) & (!g2838) & (g2891)) + ((!g1473) & (!g1507) & (!g4864) & (g2838) & (g2891)) + ((!g1473) & (!g1507) & (g4864) & (!g2838) & (g2891)) + ((!g1473) & (!g1507) & (g4864) & (g2838) & (!g2891)) + ((!g1473) & (g1507) & (!g4864) & (!g2838) & (!g2891)) + ((!g1473) & (g1507) & (!g4864) & (g2838) & (!g2891)) + ((!g1473) & (g1507) & (g4864) & (!g2838) & (!g2891)) + ((!g1473) & (g1507) & (g4864) & (g2838) & (g2891)) + ((g1473) & (!g1507) & (!g4864) & (!g2838) & (g2891)) + ((g1473) & (!g1507) & (!g4864) & (g2838) & (!g2891)) + ((g1473) & (!g1507) & (g4864) & (!g2838) & (!g2891)) + ((g1473) & (!g1507) & (g4864) & (g2838) & (!g2891)) + ((g1473) & (g1507) & (!g4864) & (!g2838) & (!g2891)) + ((g1473) & (g1507) & (!g4864) & (g2838) & (g2891)) + ((g1473) & (g1507) & (g4864) & (!g2838) & (g2891)) + ((g1473) & (g1507) & (g4864) & (g2838) & (g2891)));
	assign g4925 = (((!g2845) & (!g2885) & (!g2868) & (g2889) & (!g4866)) + ((!g2845) & (!g2885) & (!g2868) & (g2889) & (g4866)) + ((!g2845) & (!g2885) & (g2868) & (!g2889) & (g4866)) + ((!g2845) & (!g2885) & (g2868) & (g2889) & (!g4866)) + ((!g2845) & (g2885) & (!g2868) & (!g2889) & (!g4866)) + ((!g2845) & (g2885) & (!g2868) & (!g2889) & (g4866)) + ((!g2845) & (g2885) & (g2868) & (!g2889) & (!g4866)) + ((!g2845) & (g2885) & (g2868) & (g2889) & (g4866)) + ((g2845) & (!g2885) & (!g2868) & (!g2889) & (g4866)) + ((g2845) & (!g2885) & (!g2868) & (g2889) & (!g4866)) + ((g2845) & (!g2885) & (g2868) & (!g2889) & (!g4866)) + ((g2845) & (!g2885) & (g2868) & (!g2889) & (g4866)) + ((g2845) & (g2885) & (!g2868) & (!g2889) & (!g4866)) + ((g2845) & (g2885) & (!g2868) & (g2889) & (g4866)) + ((g2845) & (g2885) & (g2868) & (g2889) & (!g4866)) + ((g2845) & (g2885) & (g2868) & (g2889) & (g4866)));
	assign g4926 = (((!g830) & (!g1914) & (!g2678) & (!g4924) & (!g4925) & (key[61])) + ((!g830) & (!g1914) & (!g2678) & (!g4924) & (g4925) & (key[61])) + ((!g830) & (!g1914) & (!g2678) & (g4924) & (!g4925) & (key[61])) + ((!g830) & (!g1914) & (!g2678) & (g4924) & (g4925) & (key[61])) + ((!g830) & (!g1914) & (g2678) & (!g4924) & (!g4925) & (key[61])) + ((!g830) & (!g1914) & (g2678) & (!g4924) & (g4925) & (key[61])) + ((!g830) & (!g1914) & (g2678) & (g4924) & (!g4925) & (key[61])) + ((!g830) & (!g1914) & (g2678) & (g4924) & (g4925) & (key[61])) + ((!g830) & (g1914) & (!g2678) & (!g4924) & (!g4925) & (key[61])) + ((!g830) & (g1914) & (!g2678) & (!g4924) & (g4925) & (key[61])) + ((!g830) & (g1914) & (!g2678) & (g4924) & (!g4925) & (key[61])) + ((!g830) & (g1914) & (!g2678) & (g4924) & (g4925) & (key[61])) + ((!g830) & (g1914) & (g2678) & (!g4924) & (!g4925) & (key[61])) + ((!g830) & (g1914) & (g2678) & (!g4924) & (g4925) & (key[61])) + ((!g830) & (g1914) & (g2678) & (g4924) & (!g4925) & (key[61])) + ((!g830) & (g1914) & (g2678) & (g4924) & (g4925) & (key[61])) + ((g830) & (!g1914) & (!g2678) & (!g4924) & (g4925) & (!key[61])) + ((g830) & (!g1914) & (!g2678) & (!g4924) & (g4925) & (key[61])) + ((g830) & (!g1914) & (!g2678) & (g4924) & (g4925) & (!key[61])) + ((g830) & (!g1914) & (!g2678) & (g4924) & (g4925) & (key[61])) + ((g830) & (!g1914) & (g2678) & (!g4924) & (!g4925) & (!key[61])) + ((g830) & (!g1914) & (g2678) & (!g4924) & (!g4925) & (key[61])) + ((g830) & (!g1914) & (g2678) & (g4924) & (!g4925) & (!key[61])) + ((g830) & (!g1914) & (g2678) & (g4924) & (!g4925) & (key[61])) + ((g830) & (g1914) & (!g2678) & (g4924) & (!g4925) & (!key[61])) + ((g830) & (g1914) & (!g2678) & (g4924) & (!g4925) & (key[61])) + ((g830) & (g1914) & (!g2678) & (g4924) & (g4925) & (!key[61])) + ((g830) & (g1914) & (!g2678) & (g4924) & (g4925) & (key[61])) + ((g830) & (g1914) & (g2678) & (!g4924) & (!g4925) & (!key[61])) + ((g830) & (g1914) & (g2678) & (!g4924) & (!g4925) & (key[61])) + ((g830) & (g1914) & (g2678) & (!g4924) & (g4925) & (!key[61])) + ((g830) & (g1914) & (g2678) & (!g4924) & (g4925) & (key[61])));
	assign g4927 = (((!g2944) & (g2991) & (!g3772) & (g3773)) + ((!g2944) & (g2991) & (g3772) & (!g3773)) + ((!g2944) & (g2991) & (g3772) & (g3773)) + ((g2944) & (!g2991) & (!g3772) & (g3773)) + ((g2944) & (!g2991) & (g3772) & (!g3773)) + ((g2944) & (!g2991) & (g3772) & (g3773)) + ((g2944) & (g2991) & (!g3772) & (!g3773)) + ((g2944) & (g2991) & (!g3772) & (g3773)) + ((g2944) & (g2991) & (g3772) & (!g3773)) + ((g2944) & (g2991) & (g3772) & (g3773)));
	assign g4928 = (((!g3755) & (g3756)) + ((g3755) & (!g3756)) + ((g3755) & (g3756)));
	assign g4929 = (((!g830) & (!g2679) & (!g6297) & (key[93])) + ((!g830) & (!g2679) & (g6297) & (key[93])) + ((!g830) & (g2679) & (!g6297) & (key[93])) + ((!g830) & (g2679) & (g6297) & (key[93])) + ((g830) & (!g2679) & (g6297) & (!key[93])) + ((g830) & (!g2679) & (g6297) & (key[93])) + ((g830) & (g2679) & (!g6297) & (!key[93])) + ((g830) & (g2679) & (!g6297) & (key[93])));
	assign g4930 = (((!g4874) & (!g2845) & (!g2851) & (!g2885) & (g2900)) + ((!g4874) & (!g2845) & (!g2851) & (g2885) & (!g2900)) + ((!g4874) & (!g2845) & (g2851) & (!g2885) & (g2900)) + ((!g4874) & (!g2845) & (g2851) & (g2885) & (!g2900)) + ((!g4874) & (g2845) & (!g2851) & (!g2885) & (g2900)) + ((!g4874) & (g2845) & (!g2851) & (g2885) & (!g2900)) + ((!g4874) & (g2845) & (g2851) & (!g2885) & (!g2900)) + ((!g4874) & (g2845) & (g2851) & (g2885) & (g2900)) + ((g4874) & (!g2845) & (!g2851) & (!g2885) & (g2900)) + ((g4874) & (!g2845) & (!g2851) & (g2885) & (!g2900)) + ((g4874) & (!g2845) & (g2851) & (!g2885) & (!g2900)) + ((g4874) & (!g2845) & (g2851) & (g2885) & (g2900)) + ((g4874) & (g2845) & (!g2851) & (!g2885) & (!g2900)) + ((g4874) & (g2845) & (!g2851) & (g2885) & (g2900)) + ((g4874) & (g2845) & (g2851) & (!g2885) & (!g2900)) + ((g4874) & (g2845) & (g2851) & (g2885) & (g2900)));
	assign g8321 = (((!g5560) & (g5624) & (!g4931)) + ((!g5560) & (g5624) & (g4931)) + ((g5560) & (!g5624) & (g4931)) + ((g5560) & (g5624) & (g4931)));
	assign g4932 = (((!g830) & (!g2683) & (!g6323) & (g4931)) + ((!g830) & (!g2683) & (g6323) & (g4931)) + ((!g830) & (g2683) & (!g6323) & (g4931)) + ((!g830) & (g2683) & (g6323) & (g4931)) + ((g830) & (!g2683) & (g6323) & (!g4931)) + ((g830) & (!g2683) & (g6323) & (g4931)) + ((g830) & (g2683) & (!g6323) & (!g4931)) + ((g830) & (g2683) & (!g6323) & (g4931)));
	assign g4933 = (((!g3479) & (!g3480) & (g2979) & (g2991)) + ((!g3479) & (g3480) & (!g2979) & (g2991)) + ((!g3479) & (g3480) & (g2979) & (!g2991)) + ((!g3479) & (g3480) & (g2979) & (g2991)) + ((g3479) & (!g3480) & (!g2979) & (g2991)) + ((g3479) & (!g3480) & (g2979) & (!g2991)) + ((g3479) & (!g3480) & (g2979) & (g2991)) + ((g3479) & (g3480) & (!g2979) & (g2991)) + ((g3479) & (g3480) & (g2979) & (!g2991)) + ((g3479) & (g3480) & (g2979) & (g2991)));
	assign g4934 = (((!g3493) & (g3494)) + ((g3493) & (!g3494)) + ((g3493) & (g3494)));
	assign g4935 = (((!g830) & (!g2684) & (!g6310) & (key[189])) + ((!g830) & (!g2684) & (g6310) & (key[189])) + ((!g830) & (g2684) & (!g6310) & (key[189])) + ((!g830) & (g2684) & (g6310) & (key[189])) + ((g830) & (!g2684) & (g6310) & (!key[189])) + ((g830) & (!g2684) & (g6310) & (key[189])) + ((g830) & (g2684) & (!g6310) & (!key[189])) + ((g830) & (g2684) & (!g6310) & (key[189])));
	assign g4936 = (((!g1997) & (g1098) & (!g3448)) + ((g1997) & (!g1098) & (!g3448)) + ((g1997) & (g1098) & (!g3448)) + ((g1997) & (g1098) & (g3448)));
	assign g4937 = (((!g3430) & (!g2116) & (g2120)) + ((!g3430) & (g2116) & (!g2120)) + ((g3430) & (!g2116) & (!g2120)) + ((g3430) & (g2116) & (g2120)));
	assign g4938 = (((!g1914) & (!g1999) & (!g1132) & (g4936) & (!g4937)) + ((!g1914) & (!g1999) & (!g1132) & (g4936) & (g4937)) + ((!g1914) & (!g1999) & (g1132) & (!g4936) & (!g4937)) + ((!g1914) & (!g1999) & (g1132) & (!g4936) & (g4937)) + ((!g1914) & (g1999) & (!g1132) & (!g4936) & (!g4937)) + ((!g1914) & (g1999) & (!g1132) & (!g4936) & (g4937)) + ((!g1914) & (g1999) & (g1132) & (g4936) & (!g4937)) + ((!g1914) & (g1999) & (g1132) & (g4936) & (g4937)) + ((g1914) & (!g1999) & (!g1132) & (!g4936) & (g4937)) + ((g1914) & (!g1999) & (!g1132) & (g4936) & (g4937)) + ((g1914) & (!g1999) & (g1132) & (!g4936) & (g4937)) + ((g1914) & (!g1999) & (g1132) & (g4936) & (g4937)) + ((g1914) & (g1999) & (!g1132) & (!g4936) & (g4937)) + ((g1914) & (g1999) & (!g1132) & (g4936) & (g4937)) + ((g1914) & (g1999) & (g1132) & (!g4936) & (g4937)) + ((g1914) & (g1999) & (g1132) & (g4936) & (g4937)));
	assign g4939 = (((!g830) & (!g2690) & (!g4938) & (key[112])) + ((!g830) & (!g2690) & (g4938) & (key[112])) + ((!g830) & (g2690) & (!g4938) & (key[112])) + ((!g830) & (g2690) & (g4938) & (key[112])) + ((g830) & (!g2690) & (g4938) & (!key[112])) + ((g830) & (!g2690) & (g4938) & (key[112])) + ((g830) & (g2690) & (!g4938) & (!key[112])) + ((g830) & (g2690) & (!g4938) & (key[112])));
	assign g4940 = (((!g2649) & (!g2683) & (g3255) & (g3297) & (g4841)) + ((!g2649) & (g2683) & (!g3255) & (g3297) & (!g4841)) + ((!g2649) & (g2683) & (!g3255) & (g3297) & (g4841)) + ((!g2649) & (g2683) & (g3255) & (!g3297) & (g4841)) + ((!g2649) & (g2683) & (g3255) & (g3297) & (!g4841)) + ((!g2649) & (g2683) & (g3255) & (g3297) & (g4841)) + ((g2649) & (!g2683) & (!g3255) & (g3297) & (g4841)) + ((g2649) & (!g2683) & (g3255) & (g3297) & (!g4841)) + ((g2649) & (!g2683) & (g3255) & (g3297) & (g4841)) + ((g2649) & (g2683) & (!g3255) & (!g3297) & (g4841)) + ((g2649) & (g2683) & (!g3255) & (g3297) & (!g4841)) + ((g2649) & (g2683) & (!g3255) & (g3297) & (g4841)) + ((g2649) & (g2683) & (g3255) & (!g3297) & (!g4841)) + ((g2649) & (g2683) & (g3255) & (!g3297) & (g4841)) + ((g2649) & (g2683) & (g3255) & (g3297) & (!g4841)) + ((g2649) & (g2683) & (g3255) & (g3297) & (g4841)));
	assign g4941 = (((!g2649) & (!g2683) & (!g3255) & (!g3297) & (!g4841) & (!g5717)) + ((!g2649) & (!g2683) & (!g3255) & (!g3297) & (g4841) & (!g5717)) + ((!g2649) & (!g2683) & (!g3255) & (g3297) & (!g4841) & (!g5717)) + ((!g2649) & (!g2683) & (!g3255) & (g3297) & (g4841) & (!g5717)) + ((!g2649) & (!g2683) & (g3255) & (!g3297) & (!g4841) & (!g5717)) + ((!g2649) & (!g2683) & (g3255) & (!g3297) & (g4841) & (!g5717)) + ((!g2649) & (!g2683) & (g3255) & (g3297) & (!g4841) & (!g5717)) + ((!g2649) & (!g2683) & (g3255) & (g3297) & (g4841) & (g5717)) + ((!g2649) & (g2683) & (!g3255) & (!g3297) & (!g4841) & (!g5717)) + ((!g2649) & (g2683) & (!g3255) & (!g3297) & (g4841) & (!g5717)) + ((!g2649) & (g2683) & (!g3255) & (g3297) & (!g4841) & (g5717)) + ((!g2649) & (g2683) & (!g3255) & (g3297) & (g4841) & (g5717)) + ((!g2649) & (g2683) & (g3255) & (!g3297) & (!g4841) & (!g5717)) + ((!g2649) & (g2683) & (g3255) & (!g3297) & (g4841) & (g5717)) + ((!g2649) & (g2683) & (g3255) & (g3297) & (!g4841) & (g5717)) + ((!g2649) & (g2683) & (g3255) & (g3297) & (g4841) & (g5717)) + ((g2649) & (!g2683) & (!g3255) & (!g3297) & (!g4841) & (!g5717)) + ((g2649) & (!g2683) & (!g3255) & (!g3297) & (g4841) & (!g5717)) + ((g2649) & (!g2683) & (!g3255) & (g3297) & (!g4841) & (!g5717)) + ((g2649) & (!g2683) & (!g3255) & (g3297) & (g4841) & (g5717)) + ((g2649) & (!g2683) & (g3255) & (!g3297) & (!g4841) & (!g5717)) + ((g2649) & (!g2683) & (g3255) & (!g3297) & (g4841) & (!g5717)) + ((g2649) & (!g2683) & (g3255) & (g3297) & (!g4841) & (g5717)) + ((g2649) & (!g2683) & (g3255) & (g3297) & (g4841) & (g5717)) + ((g2649) & (g2683) & (!g3255) & (!g3297) & (!g4841) & (!g5717)) + ((g2649) & (g2683) & (!g3255) & (!g3297) & (g4841) & (g5717)) + ((g2649) & (g2683) & (!g3255) & (g3297) & (!g4841) & (g5717)) + ((g2649) & (g2683) & (!g3255) & (g3297) & (g4841) & (g5717)) + ((g2649) & (g2683) & (g3255) & (!g3297) & (!g4841) & (g5717)) + ((g2649) & (g2683) & (g3255) & (!g3297) & (g4841) & (g5717)) + ((g2649) & (g2683) & (g3255) & (g3297) & (!g4841) & (g5717)) + ((g2649) & (g2683) & (g3255) & (g3297) & (g4841) & (g5717)));
	assign g4942 = (((!g2678) & (!g2758) & (!g3303) & (g3333) & (!g4887) & (!g4888)) + ((!g2678) & (!g2758) & (!g3303) & (g3333) & (!g4887) & (g4888)) + ((!g2678) & (!g2758) & (!g3303) & (g3333) & (g4887) & (!g4888)) + ((!g2678) & (!g2758) & (!g3303) & (g3333) & (g4887) & (g4888)) + ((!g2678) & (!g2758) & (g3303) & (!g3333) & (!g4887) & (g4888)) + ((!g2678) & (!g2758) & (g3303) & (!g3333) & (g4887) & (!g4888)) + ((!g2678) & (!g2758) & (g3303) & (!g3333) & (g4887) & (g4888)) + ((!g2678) & (!g2758) & (g3303) & (g3333) & (!g4887) & (!g4888)) + ((!g2678) & (g2758) & (!g3303) & (!g3333) & (!g4887) & (!g4888)) + ((!g2678) & (g2758) & (!g3303) & (!g3333) & (!g4887) & (g4888)) + ((!g2678) & (g2758) & (!g3303) & (!g3333) & (g4887) & (!g4888)) + ((!g2678) & (g2758) & (!g3303) & (!g3333) & (g4887) & (g4888)) + ((!g2678) & (g2758) & (g3303) & (!g3333) & (!g4887) & (!g4888)) + ((!g2678) & (g2758) & (g3303) & (g3333) & (!g4887) & (g4888)) + ((!g2678) & (g2758) & (g3303) & (g3333) & (g4887) & (!g4888)) + ((!g2678) & (g2758) & (g3303) & (g3333) & (g4887) & (g4888)) + ((g2678) & (!g2758) & (!g3303) & (!g3333) & (!g4887) & (g4888)) + ((g2678) & (!g2758) & (!g3303) & (!g3333) & (g4887) & (!g4888)) + ((g2678) & (!g2758) & (!g3303) & (!g3333) & (g4887) & (g4888)) + ((g2678) & (!g2758) & (!g3303) & (g3333) & (!g4887) & (!g4888)) + ((g2678) & (!g2758) & (g3303) & (!g3333) & (!g4887) & (!g4888)) + ((g2678) & (!g2758) & (g3303) & (!g3333) & (!g4887) & (g4888)) + ((g2678) & (!g2758) & (g3303) & (!g3333) & (g4887) & (!g4888)) + ((g2678) & (!g2758) & (g3303) & (!g3333) & (g4887) & (g4888)) + ((g2678) & (g2758) & (!g3303) & (!g3333) & (!g4887) & (!g4888)) + ((g2678) & (g2758) & (!g3303) & (g3333) & (!g4887) & (g4888)) + ((g2678) & (g2758) & (!g3303) & (g3333) & (g4887) & (!g4888)) + ((g2678) & (g2758) & (!g3303) & (g3333) & (g4887) & (g4888)) + ((g2678) & (g2758) & (g3303) & (g3333) & (!g4887) & (!g4888)) + ((g2678) & (g2758) & (g3303) & (g3333) & (!g4887) & (g4888)) + ((g2678) & (g2758) & (g3303) & (g3333) & (g4887) & (!g4888)) + ((g2678) & (g2758) & (g3303) & (g3333) & (g4887) & (g4888)));
	assign g4943 = (((g830) & (!g1914) & (!g2703) & (!g4941) & (g4942)) + ((g830) & (!g1914) & (!g2703) & (g4941) & (g4942)) + ((g830) & (!g1914) & (g2703) & (!g4941) & (!g4942)) + ((g830) & (!g1914) & (g2703) & (g4941) & (!g4942)) + ((g830) & (g1914) & (!g2703) & (g4941) & (!g4942)) + ((g830) & (g1914) & (!g2703) & (g4941) & (g4942)) + ((g830) & (g1914) & (g2703) & (!g4941) & (!g4942)) + ((g830) & (g1914) & (g2703) & (!g4941) & (g4942)));
	assign g4944 = (((!g2304) & (!g3559) & (g2326)) + ((g2304) & (!g3559) & (!g2326)) + ((g2304) & (!g3559) & (g2326)) + ((g2304) & (g3559) & (g2326)));
	assign g4945 = (((!g1944) & (!g2123) & (g3572)) + ((!g1944) & (g2123) & (!g3572)) + ((g1944) & (!g2123) & (!g3572)) + ((g1944) & (g2123) & (g3572)));
	assign g4946 = (((!g1914) & (!g2360) & (!g4944) & (!g2364) & (g4945)) + ((!g1914) & (!g2360) & (!g4944) & (g2364) & (g4945)) + ((!g1914) & (!g2360) & (g4944) & (!g2364) & (g4945)) + ((!g1914) & (!g2360) & (g4944) & (g2364) & (g4945)) + ((!g1914) & (g2360) & (!g4944) & (!g2364) & (g4945)) + ((!g1914) & (g2360) & (!g4944) & (g2364) & (g4945)) + ((!g1914) & (g2360) & (g4944) & (!g2364) & (g4945)) + ((!g1914) & (g2360) & (g4944) & (g2364) & (g4945)) + ((g1914) & (!g2360) & (!g4944) & (g2364) & (!g4945)) + ((g1914) & (!g2360) & (!g4944) & (g2364) & (g4945)) + ((g1914) & (!g2360) & (g4944) & (!g2364) & (!g4945)) + ((g1914) & (!g2360) & (g4944) & (!g2364) & (g4945)) + ((g1914) & (g2360) & (!g4944) & (!g2364) & (!g4945)) + ((g1914) & (g2360) & (!g4944) & (!g2364) & (g4945)) + ((g1914) & (g2360) & (g4944) & (g2364) & (!g4945)) + ((g1914) & (g2360) & (g4944) & (g2364) & (g4945)));
	assign g4947 = (((!g830) & (!g2708) & (!g4946) & (nonce[16])) + ((!g830) & (!g2708) & (g4946) & (nonce[16])) + ((!g830) & (g2708) & (!g4946) & (nonce[16])) + ((!g830) & (g2708) & (g4946) & (nonce[16])) + ((g830) & (!g2708) & (g4946) & (!nonce[16])) + ((g830) & (!g2708) & (g4946) & (nonce[16])) + ((g830) & (g2708) & (!g4946) & (!nonce[16])) + ((g830) & (g2708) & (!g4946) & (nonce[16])));
	assign g4948 = (((!g2311) & (g2314) & (!g3606)) + ((g2311) & (!g2314) & (!g3606)) + ((g2311) & (g2314) & (!g3606)) + ((g2311) & (g2314) & (g3606)));
	assign g4949 = (((!g1983) & (!g3588) & (g2125)) + ((!g1983) & (g3588) & (!g2125)) + ((g1983) & (!g3588) & (!g2125)) + ((g1983) & (g3588) & (g2125)));
	assign g4950 = (((!g1914) & (!g2354) & (!g2362) & (g4948) & (!g4949)) + ((!g1914) & (!g2354) & (!g2362) & (g4948) & (g4949)) + ((!g1914) & (!g2354) & (g2362) & (!g4948) & (!g4949)) + ((!g1914) & (!g2354) & (g2362) & (!g4948) & (g4949)) + ((!g1914) & (g2354) & (!g2362) & (!g4948) & (!g4949)) + ((!g1914) & (g2354) & (!g2362) & (!g4948) & (g4949)) + ((!g1914) & (g2354) & (g2362) & (g4948) & (!g4949)) + ((!g1914) & (g2354) & (g2362) & (g4948) & (g4949)) + ((g1914) & (!g2354) & (!g2362) & (!g4948) & (g4949)) + ((g1914) & (!g2354) & (!g2362) & (g4948) & (g4949)) + ((g1914) & (!g2354) & (g2362) & (!g4948) & (g4949)) + ((g1914) & (!g2354) & (g2362) & (g4948) & (g4949)) + ((g1914) & (g2354) & (!g2362) & (!g4948) & (g4949)) + ((g1914) & (g2354) & (!g2362) & (g4948) & (g4949)) + ((g1914) & (g2354) & (g2362) & (!g4948) & (g4949)) + ((g1914) & (g2354) & (g2362) & (g4948) & (g4949)));
	assign g4951 = (((!g830) & (!g2713) & (!g4950) & (key[240])) + ((!g830) & (!g2713) & (g4950) & (key[240])) + ((!g830) & (g2713) & (!g4950) & (key[240])) + ((!g830) & (g2713) & (g4950) & (key[240])) + ((g830) & (!g2713) & (g4950) & (!key[240])) + ((g830) & (!g2713) & (g4950) & (key[240])) + ((g830) & (g2713) & (!g4950) & (!key[240])) + ((g830) & (g2713) & (!g4950) & (key[240])));
	assign g4952 = (((!g1959) & (g1098) & (!g3625)) + ((g1959) & (!g1098) & (!g3625)) + ((g1959) & (g1098) & (!g3625)) + ((g1959) & (g1098) & (g3625)));
	assign g4953 = (((!g2110) & (!g2125) & (g3638)) + ((!g2110) & (g2125) & (!g3638)) + ((g2110) & (!g2125) & (!g3638)) + ((g2110) & (g2125) & (g3638)));
	assign g4954 = (((!g1914) & (!g1961) & (!g1132) & (!g4952) & (g4953)) + ((!g1914) & (!g1961) & (!g1132) & (g4952) & (g4953)) + ((!g1914) & (!g1961) & (g1132) & (!g4952) & (g4953)) + ((!g1914) & (!g1961) & (g1132) & (g4952) & (g4953)) + ((!g1914) & (g1961) & (!g1132) & (!g4952) & (g4953)) + ((!g1914) & (g1961) & (!g1132) & (g4952) & (g4953)) + ((!g1914) & (g1961) & (g1132) & (!g4952) & (g4953)) + ((!g1914) & (g1961) & (g1132) & (g4952) & (g4953)) + ((g1914) & (!g1961) & (!g1132) & (g4952) & (!g4953)) + ((g1914) & (!g1961) & (!g1132) & (g4952) & (g4953)) + ((g1914) & (!g1961) & (g1132) & (!g4952) & (!g4953)) + ((g1914) & (!g1961) & (g1132) & (!g4952) & (g4953)) + ((g1914) & (g1961) & (!g1132) & (!g4952) & (!g4953)) + ((g1914) & (g1961) & (!g1132) & (!g4952) & (g4953)) + ((g1914) & (g1961) & (g1132) & (g4952) & (!g4953)) + ((g1914) & (g1961) & (g1132) & (g4952) & (g4953)));
	assign g4955 = (((!g830) & (!g2718) & (!g4954) & (key[16])) + ((!g830) & (!g2718) & (g4954) & (key[16])) + ((!g830) & (g2718) & (!g4954) & (key[16])) + ((!g830) & (g2718) & (g4954) & (key[16])) + ((g830) & (!g2718) & (g4954) & (!key[16])) + ((g830) & (!g2718) & (g4954) & (key[16])) + ((g830) & (g2718) & (!g4954) & (!key[16])) + ((g830) & (g2718) & (!g4954) & (key[16])));
	assign g4956 = (((!g2320) & (g2326) & (!g3673)) + ((g2320) & (!g2326) & (!g3673)) + ((g2320) & (g2326) & (!g3673)) + ((g2320) & (g2326) & (g3673)));
	assign g4957 = (((!g1982) & (!g2112) & (g3654)) + ((!g1982) & (g2112) & (!g3654)) + ((g1982) & (!g2112) & (!g3654)) + ((g1982) & (g2112) & (g3654)));
	assign g4958 = (((!g1914) & (!g2350) & (!g2364) & (g4956) & (!g4957)) + ((!g1914) & (!g2350) & (!g2364) & (g4956) & (g4957)) + ((!g1914) & (!g2350) & (g2364) & (!g4956) & (!g4957)) + ((!g1914) & (!g2350) & (g2364) & (!g4956) & (g4957)) + ((!g1914) & (g2350) & (!g2364) & (!g4956) & (!g4957)) + ((!g1914) & (g2350) & (!g2364) & (!g4956) & (g4957)) + ((!g1914) & (g2350) & (g2364) & (g4956) & (!g4957)) + ((!g1914) & (g2350) & (g2364) & (g4956) & (g4957)) + ((g1914) & (!g2350) & (!g2364) & (!g4956) & (g4957)) + ((g1914) & (!g2350) & (!g2364) & (g4956) & (g4957)) + ((g1914) & (!g2350) & (g2364) & (!g4956) & (g4957)) + ((g1914) & (!g2350) & (g2364) & (g4956) & (g4957)) + ((g1914) & (g2350) & (!g2364) & (!g4956) & (g4957)) + ((g1914) & (g2350) & (!g2364) & (g4956) & (g4957)) + ((g1914) & (g2350) & (g2364) & (!g4956) & (g4957)) + ((g1914) & (g2350) & (g2364) & (g4956) & (g4957)));
	assign g8322 = (((!g5560) & (g5625) & (!g4959)) + ((!g5560) & (g5625) & (g4959)) + ((g5560) & (!g5625) & (g4959)) + ((g5560) & (g5625) & (g4959)));
	assign g4960 = (((!g830) & (!g2723) & (!g4958) & (g4959)) + ((!g830) & (!g2723) & (g4958) & (g4959)) + ((!g830) & (g2723) & (!g4958) & (g4959)) + ((!g830) & (g2723) & (g4958) & (g4959)) + ((g830) & (!g2723) & (g4958) & (!g4959)) + ((g830) & (!g2723) & (g4958) & (g4959)) + ((g830) & (g2723) & (!g4958) & (!g4959)) + ((g830) & (g2723) & (!g4958) & (g4959)));
	assign g4961 = (((!g3222) & (!g3301) & (g3279) & (g3307) & (g4852)) + ((!g3222) & (g3301) & (!g3279) & (g3307) & (!g4852)) + ((!g3222) & (g3301) & (!g3279) & (g3307) & (g4852)) + ((!g3222) & (g3301) & (g3279) & (!g3307) & (g4852)) + ((!g3222) & (g3301) & (g3279) & (g3307) & (!g4852)) + ((!g3222) & (g3301) & (g3279) & (g3307) & (g4852)) + ((g3222) & (!g3301) & (!g3279) & (g3307) & (g4852)) + ((g3222) & (!g3301) & (g3279) & (g3307) & (!g4852)) + ((g3222) & (!g3301) & (g3279) & (g3307) & (g4852)) + ((g3222) & (g3301) & (!g3279) & (!g3307) & (g4852)) + ((g3222) & (g3301) & (!g3279) & (g3307) & (!g4852)) + ((g3222) & (g3301) & (!g3279) & (g3307) & (g4852)) + ((g3222) & (g3301) & (g3279) & (!g3307) & (!g4852)) + ((g3222) & (g3301) & (g3279) & (!g3307) & (g4852)) + ((g3222) & (g3301) & (g3279) & (g3307) & (!g4852)) + ((g3222) & (g3301) & (g3279) & (g3307) & (g4852)));
	assign g4962 = (((!g3222) & (!g3301) & (!g3279) & (!g3307) & (!g4852) & (!g5718)) + ((!g3222) & (!g3301) & (!g3279) & (!g3307) & (g4852) & (!g5718)) + ((!g3222) & (!g3301) & (!g3279) & (g3307) & (!g4852) & (!g5718)) + ((!g3222) & (!g3301) & (!g3279) & (g3307) & (g4852) & (!g5718)) + ((!g3222) & (!g3301) & (g3279) & (!g3307) & (!g4852) & (!g5718)) + ((!g3222) & (!g3301) & (g3279) & (!g3307) & (g4852) & (!g5718)) + ((!g3222) & (!g3301) & (g3279) & (g3307) & (!g4852) & (!g5718)) + ((!g3222) & (!g3301) & (g3279) & (g3307) & (g4852) & (g5718)) + ((!g3222) & (g3301) & (!g3279) & (!g3307) & (!g4852) & (!g5718)) + ((!g3222) & (g3301) & (!g3279) & (!g3307) & (g4852) & (!g5718)) + ((!g3222) & (g3301) & (!g3279) & (g3307) & (!g4852) & (g5718)) + ((!g3222) & (g3301) & (!g3279) & (g3307) & (g4852) & (g5718)) + ((!g3222) & (g3301) & (g3279) & (!g3307) & (!g4852) & (!g5718)) + ((!g3222) & (g3301) & (g3279) & (!g3307) & (g4852) & (g5718)) + ((!g3222) & (g3301) & (g3279) & (g3307) & (!g4852) & (g5718)) + ((!g3222) & (g3301) & (g3279) & (g3307) & (g4852) & (g5718)) + ((g3222) & (!g3301) & (!g3279) & (!g3307) & (!g4852) & (!g5718)) + ((g3222) & (!g3301) & (!g3279) & (!g3307) & (g4852) & (!g5718)) + ((g3222) & (!g3301) & (!g3279) & (g3307) & (!g4852) & (!g5718)) + ((g3222) & (!g3301) & (!g3279) & (g3307) & (g4852) & (g5718)) + ((g3222) & (!g3301) & (g3279) & (!g3307) & (!g4852) & (!g5718)) + ((g3222) & (!g3301) & (g3279) & (!g3307) & (g4852) & (!g5718)) + ((g3222) & (!g3301) & (g3279) & (g3307) & (!g4852) & (g5718)) + ((g3222) & (!g3301) & (g3279) & (g3307) & (g4852) & (g5718)) + ((g3222) & (g3301) & (!g3279) & (!g3307) & (!g4852) & (!g5718)) + ((g3222) & (g3301) & (!g3279) & (!g3307) & (g4852) & (g5718)) + ((g3222) & (g3301) & (!g3279) & (g3307) & (!g4852) & (g5718)) + ((g3222) & (g3301) & (!g3279) & (g3307) & (g4852) & (g5718)) + ((g3222) & (g3301) & (g3279) & (!g3307) & (!g4852) & (g5718)) + ((g3222) & (g3301) & (g3279) & (!g3307) & (g4852) & (g5718)) + ((g3222) & (g3301) & (g3279) & (g3307) & (!g4852) & (g5718)) + ((g3222) & (g3301) & (g3279) & (g3307) & (g4852) & (g5718)));
	assign g4963 = (((!g3291) & (!g3339) & (!g3312) & (g3348) & (!g4904) & (!g4905)) + ((!g3291) & (!g3339) & (!g3312) & (g3348) & (!g4904) & (g4905)) + ((!g3291) & (!g3339) & (!g3312) & (g3348) & (g4904) & (!g4905)) + ((!g3291) & (!g3339) & (!g3312) & (g3348) & (g4904) & (g4905)) + ((!g3291) & (!g3339) & (g3312) & (!g3348) & (!g4904) & (g4905)) + ((!g3291) & (!g3339) & (g3312) & (!g3348) & (g4904) & (!g4905)) + ((!g3291) & (!g3339) & (g3312) & (!g3348) & (g4904) & (g4905)) + ((!g3291) & (!g3339) & (g3312) & (g3348) & (!g4904) & (!g4905)) + ((!g3291) & (g3339) & (!g3312) & (!g3348) & (!g4904) & (!g4905)) + ((!g3291) & (g3339) & (!g3312) & (!g3348) & (!g4904) & (g4905)) + ((!g3291) & (g3339) & (!g3312) & (!g3348) & (g4904) & (!g4905)) + ((!g3291) & (g3339) & (!g3312) & (!g3348) & (g4904) & (g4905)) + ((!g3291) & (g3339) & (g3312) & (!g3348) & (!g4904) & (!g4905)) + ((!g3291) & (g3339) & (g3312) & (g3348) & (!g4904) & (g4905)) + ((!g3291) & (g3339) & (g3312) & (g3348) & (g4904) & (!g4905)) + ((!g3291) & (g3339) & (g3312) & (g3348) & (g4904) & (g4905)) + ((g3291) & (!g3339) & (!g3312) & (!g3348) & (!g4904) & (g4905)) + ((g3291) & (!g3339) & (!g3312) & (!g3348) & (g4904) & (!g4905)) + ((g3291) & (!g3339) & (!g3312) & (!g3348) & (g4904) & (g4905)) + ((g3291) & (!g3339) & (!g3312) & (g3348) & (!g4904) & (!g4905)) + ((g3291) & (!g3339) & (g3312) & (!g3348) & (!g4904) & (!g4905)) + ((g3291) & (!g3339) & (g3312) & (!g3348) & (!g4904) & (g4905)) + ((g3291) & (!g3339) & (g3312) & (!g3348) & (g4904) & (!g4905)) + ((g3291) & (!g3339) & (g3312) & (!g3348) & (g4904) & (g4905)) + ((g3291) & (g3339) & (!g3312) & (!g3348) & (!g4904) & (!g4905)) + ((g3291) & (g3339) & (!g3312) & (g3348) & (!g4904) & (g4905)) + ((g3291) & (g3339) & (!g3312) & (g3348) & (g4904) & (!g4905)) + ((g3291) & (g3339) & (!g3312) & (g3348) & (g4904) & (g4905)) + ((g3291) & (g3339) & (g3312) & (g3348) & (!g4904) & (!g4905)) + ((g3291) & (g3339) & (g3312) & (g3348) & (!g4904) & (g4905)) + ((g3291) & (g3339) & (g3312) & (g3348) & (g4904) & (!g4905)) + ((g3291) & (g3339) & (g3312) & (g3348) & (g4904) & (g4905)));
	assign g4964 = (((g830) & (!g1914) & (!g2728) & (!g4962) & (g4963)) + ((g830) & (!g1914) & (!g2728) & (g4962) & (g4963)) + ((g830) & (!g1914) & (g2728) & (!g4962) & (!g4963)) + ((g830) & (!g1914) & (g2728) & (g4962) & (!g4963)) + ((g830) & (g1914) & (!g2728) & (g4962) & (!g4963)) + ((g830) & (g1914) & (!g2728) & (g4962) & (g4963)) + ((g830) & (g1914) & (g2728) & (!g4962) & (!g4963)) + ((g830) & (g1914) & (g2728) & (!g4962) & (g4963)));
	assign g4965 = (((!g1992) & (!g1994) & (!g2253) & (g2290) & (!g4915)) + ((!g1992) & (!g1994) & (!g2253) & (g2290) & (g4915)) + ((!g1992) & (!g1994) & (g2253) & (!g2290) & (!g4915)) + ((!g1992) & (!g1994) & (g2253) & (g2290) & (g4915)) + ((!g1992) & (g1994) & (!g2253) & (!g2290) & (!g4915)) + ((!g1992) & (g1994) & (!g2253) & (!g2290) & (g4915)) + ((!g1992) & (g1994) & (g2253) & (!g2290) & (g4915)) + ((!g1992) & (g1994) & (g2253) & (g2290) & (!g4915)) + ((g1992) & (!g1994) & (!g2253) & (!g2290) & (!g4915)) + ((g1992) & (!g1994) & (!g2253) & (g2290) & (g4915)) + ((g1992) & (!g1994) & (g2253) & (!g2290) & (!g4915)) + ((g1992) & (!g1994) & (g2253) & (!g2290) & (g4915)) + ((g1992) & (g1994) & (!g2253) & (!g2290) & (g4915)) + ((g1992) & (g1994) & (!g2253) & (g2290) & (!g4915)) + ((g1992) & (g1994) & (g2253) & (g2290) & (!g4915)) + ((g1992) & (g1994) & (g2253) & (g2290) & (g4915)));
	assign g4966 = (((!g2236) & (!g2273) & (!g2239) & (g2281) & (!g4917)) + ((!g2236) & (!g2273) & (!g2239) & (g2281) & (g4917)) + ((!g2236) & (!g2273) & (g2239) & (!g2281) & (!g4917)) + ((!g2236) & (!g2273) & (g2239) & (g2281) & (g4917)) + ((!g2236) & (g2273) & (!g2239) & (!g2281) & (!g4917)) + ((!g2236) & (g2273) & (!g2239) & (!g2281) & (g4917)) + ((!g2236) & (g2273) & (g2239) & (!g2281) & (g4917)) + ((!g2236) & (g2273) & (g2239) & (g2281) & (!g4917)) + ((g2236) & (!g2273) & (!g2239) & (!g2281) & (!g4917)) + ((g2236) & (!g2273) & (!g2239) & (g2281) & (g4917)) + ((g2236) & (!g2273) & (g2239) & (!g2281) & (!g4917)) + ((g2236) & (!g2273) & (g2239) & (!g2281) & (g4917)) + ((g2236) & (g2273) & (!g2239) & (!g2281) & (g4917)) + ((g2236) & (g2273) & (!g2239) & (g2281) & (!g4917)) + ((g2236) & (g2273) & (g2239) & (g2281) & (!g4917)) + ((g2236) & (g2273) & (g2239) & (g2281) & (g4917)));
	assign g4967 = (((!g830) & (!g1914) & (!g2733) & (!g4965) & (!g4966) & (key[208])) + ((!g830) & (!g1914) & (!g2733) & (!g4965) & (g4966) & (key[208])) + ((!g830) & (!g1914) & (!g2733) & (g4965) & (!g4966) & (key[208])) + ((!g830) & (!g1914) & (!g2733) & (g4965) & (g4966) & (key[208])) + ((!g830) & (!g1914) & (g2733) & (!g4965) & (!g4966) & (key[208])) + ((!g830) & (!g1914) & (g2733) & (!g4965) & (g4966) & (key[208])) + ((!g830) & (!g1914) & (g2733) & (g4965) & (!g4966) & (key[208])) + ((!g830) & (!g1914) & (g2733) & (g4965) & (g4966) & (key[208])) + ((!g830) & (g1914) & (!g2733) & (!g4965) & (!g4966) & (key[208])) + ((!g830) & (g1914) & (!g2733) & (!g4965) & (g4966) & (key[208])) + ((!g830) & (g1914) & (!g2733) & (g4965) & (!g4966) & (key[208])) + ((!g830) & (g1914) & (!g2733) & (g4965) & (g4966) & (key[208])) + ((!g830) & (g1914) & (g2733) & (!g4965) & (!g4966) & (key[208])) + ((!g830) & (g1914) & (g2733) & (!g4965) & (g4966) & (key[208])) + ((!g830) & (g1914) & (g2733) & (g4965) & (!g4966) & (key[208])) + ((!g830) & (g1914) & (g2733) & (g4965) & (g4966) & (key[208])) + ((g830) & (!g1914) & (!g2733) & (!g4965) & (g4966) & (!key[208])) + ((g830) & (!g1914) & (!g2733) & (!g4965) & (g4966) & (key[208])) + ((g830) & (!g1914) & (!g2733) & (g4965) & (g4966) & (!key[208])) + ((g830) & (!g1914) & (!g2733) & (g4965) & (g4966) & (key[208])) + ((g830) & (!g1914) & (g2733) & (!g4965) & (!g4966) & (!key[208])) + ((g830) & (!g1914) & (g2733) & (!g4965) & (!g4966) & (key[208])) + ((g830) & (!g1914) & (g2733) & (g4965) & (!g4966) & (!key[208])) + ((g830) & (!g1914) & (g2733) & (g4965) & (!g4966) & (key[208])) + ((g830) & (g1914) & (!g2733) & (g4965) & (!g4966) & (!key[208])) + ((g830) & (g1914) & (!g2733) & (g4965) & (!g4966) & (key[208])) + ((g830) & (g1914) & (!g2733) & (g4965) & (g4966) & (!key[208])) + ((g830) & (g1914) & (!g2733) & (g4965) & (g4966) & (key[208])) + ((g830) & (g1914) & (g2733) & (!g4965) & (!g4966) & (!key[208])) + ((g830) & (g1914) & (g2733) & (!g4965) & (!g4966) & (key[208])) + ((g830) & (g1914) & (g2733) & (!g4965) & (g4966) & (!key[208])) + ((g830) & (g1914) & (g2733) & (!g4965) & (g4966) & (key[208])));
	assign g4968 = (((!g2311) & (g2323) & (!g3782)) + ((g2311) & (!g2323) & (!g3782)) + ((g2311) & (g2323) & (!g3782)) + ((g2311) & (g2323) & (g3782)));
	assign g4969 = (((!g1945) & (!g2120) & (g3795)) + ((!g1945) & (g2120) & (!g3795)) + ((g1945) & (!g2120) & (!g3795)) + ((g1945) & (g2120) & (g3795)));
	assign g4970 = (((!g1914) & (!g2354) & (!g2356) & (!g4968) & (g4969)) + ((!g1914) & (!g2354) & (!g2356) & (g4968) & (g4969)) + ((!g1914) & (!g2354) & (g2356) & (!g4968) & (g4969)) + ((!g1914) & (!g2354) & (g2356) & (g4968) & (g4969)) + ((!g1914) & (g2354) & (!g2356) & (!g4968) & (g4969)) + ((!g1914) & (g2354) & (!g2356) & (g4968) & (g4969)) + ((!g1914) & (g2354) & (g2356) & (!g4968) & (g4969)) + ((!g1914) & (g2354) & (g2356) & (g4968) & (g4969)) + ((g1914) & (!g2354) & (!g2356) & (g4968) & (!g4969)) + ((g1914) & (!g2354) & (!g2356) & (g4968) & (g4969)) + ((g1914) & (!g2354) & (g2356) & (!g4968) & (!g4969)) + ((g1914) & (!g2354) & (g2356) & (!g4968) & (g4969)) + ((g1914) & (g2354) & (!g2356) & (!g4968) & (!g4969)) + ((g1914) & (g2354) & (!g2356) & (!g4968) & (g4969)) + ((g1914) & (g2354) & (g2356) & (g4968) & (!g4969)) + ((g1914) & (g2354) & (g2356) & (g4968) & (g4969)));
	assign g4971 = (((!g830) & (!g2742) & (!g4970) & (key[144])) + ((!g830) & (!g2742) & (g4970) & (key[144])) + ((!g830) & (g2742) & (!g4970) & (key[144])) + ((!g830) & (g2742) & (g4970) & (key[144])) + ((g830) & (!g2742) & (g4970) & (!key[144])) + ((g830) & (!g2742) & (g4970) & (key[144])) + ((g830) & (g2742) & (!g4970) & (!key[144])) + ((g830) & (g2742) & (!g4970) & (key[144])));
	assign g4972 = (((!g2227) & (!g2279) & (!g2239) & (g2281) & (!g4907)) + ((!g2227) & (!g2279) & (!g2239) & (g2281) & (g4907)) + ((!g2227) & (!g2279) & (g2239) & (!g2281) & (!g4907)) + ((!g2227) & (!g2279) & (g2239) & (g2281) & (g4907)) + ((!g2227) & (g2279) & (!g2239) & (!g2281) & (!g4907)) + ((!g2227) & (g2279) & (!g2239) & (!g2281) & (g4907)) + ((!g2227) & (g2279) & (g2239) & (!g2281) & (g4907)) + ((!g2227) & (g2279) & (g2239) & (g2281) & (!g4907)) + ((g2227) & (!g2279) & (!g2239) & (!g2281) & (!g4907)) + ((g2227) & (!g2279) & (!g2239) & (g2281) & (g4907)) + ((g2227) & (!g2279) & (g2239) & (!g2281) & (!g4907)) + ((g2227) & (!g2279) & (g2239) & (!g2281) & (g4907)) + ((g2227) & (g2279) & (!g2239) & (!g2281) & (g4907)) + ((g2227) & (g2279) & (!g2239) & (g2281) & (!g4907)) + ((g2227) & (g2279) & (g2239) & (g2281) & (!g4907)) + ((g2227) & (g2279) & (g2239) & (g2281) & (g4907)));
	assign g4973 = (((!g1954) & (!g1956) & (!g2253) & (g2290) & (!g4909)) + ((!g1954) & (!g1956) & (!g2253) & (g2290) & (g4909)) + ((!g1954) & (!g1956) & (g2253) & (!g2290) & (!g4909)) + ((!g1954) & (!g1956) & (g2253) & (g2290) & (g4909)) + ((!g1954) & (g1956) & (!g2253) & (!g2290) & (!g4909)) + ((!g1954) & (g1956) & (!g2253) & (!g2290) & (g4909)) + ((!g1954) & (g1956) & (g2253) & (!g2290) & (g4909)) + ((!g1954) & (g1956) & (g2253) & (g2290) & (!g4909)) + ((g1954) & (!g1956) & (!g2253) & (!g2290) & (!g4909)) + ((g1954) & (!g1956) & (!g2253) & (g2290) & (g4909)) + ((g1954) & (!g1956) & (g2253) & (!g2290) & (!g4909)) + ((g1954) & (!g1956) & (g2253) & (!g2290) & (g4909)) + ((g1954) & (g1956) & (!g2253) & (!g2290) & (g4909)) + ((g1954) & (g1956) & (!g2253) & (g2290) & (!g4909)) + ((g1954) & (g1956) & (g2253) & (g2290) & (!g4909)) + ((g1954) & (g1956) & (g2253) & (g2290) & (g4909)));
	assign g4974 = (((!g830) & (!g1914) & (!g2747) & (!g4972) & (!g4973) & (nonce[48])) + ((!g830) & (!g1914) & (!g2747) & (!g4972) & (g4973) & (nonce[48])) + ((!g830) & (!g1914) & (!g2747) & (g4972) & (!g4973) & (nonce[48])) + ((!g830) & (!g1914) & (!g2747) & (g4972) & (g4973) & (nonce[48])) + ((!g830) & (!g1914) & (g2747) & (!g4972) & (!g4973) & (nonce[48])) + ((!g830) & (!g1914) & (g2747) & (!g4972) & (g4973) & (nonce[48])) + ((!g830) & (!g1914) & (g2747) & (g4972) & (!g4973) & (nonce[48])) + ((!g830) & (!g1914) & (g2747) & (g4972) & (g4973) & (nonce[48])) + ((!g830) & (g1914) & (!g2747) & (!g4972) & (!g4973) & (nonce[48])) + ((!g830) & (g1914) & (!g2747) & (!g4972) & (g4973) & (nonce[48])) + ((!g830) & (g1914) & (!g2747) & (g4972) & (!g4973) & (nonce[48])) + ((!g830) & (g1914) & (!g2747) & (g4972) & (g4973) & (nonce[48])) + ((!g830) & (g1914) & (g2747) & (!g4972) & (!g4973) & (nonce[48])) + ((!g830) & (g1914) & (g2747) & (!g4972) & (g4973) & (nonce[48])) + ((!g830) & (g1914) & (g2747) & (g4972) & (!g4973) & (nonce[48])) + ((!g830) & (g1914) & (g2747) & (g4972) & (g4973) & (nonce[48])) + ((g830) & (!g1914) & (!g2747) & (!g4972) & (g4973) & (!nonce[48])) + ((g830) & (!g1914) & (!g2747) & (!g4972) & (g4973) & (nonce[48])) + ((g830) & (!g1914) & (!g2747) & (g4972) & (g4973) & (!nonce[48])) + ((g830) & (!g1914) & (!g2747) & (g4972) & (g4973) & (nonce[48])) + ((g830) & (!g1914) & (g2747) & (!g4972) & (!g4973) & (!nonce[48])) + ((g830) & (!g1914) & (g2747) & (!g4972) & (!g4973) & (nonce[48])) + ((g830) & (!g1914) & (g2747) & (g4972) & (!g4973) & (!nonce[48])) + ((g830) & (!g1914) & (g2747) & (g4972) & (!g4973) & (nonce[48])) + ((g830) & (g1914) & (!g2747) & (g4972) & (!g4973) & (!nonce[48])) + ((g830) & (g1914) & (!g2747) & (g4972) & (!g4973) & (nonce[48])) + ((g830) & (g1914) & (!g2747) & (g4972) & (g4973) & (!nonce[48])) + ((g830) & (g1914) & (!g2747) & (g4972) & (g4973) & (nonce[48])) + ((g830) & (g1914) & (g2747) & (!g4972) & (!g4973) & (!nonce[48])) + ((g830) & (g1914) & (g2747) & (!g4972) & (!g4973) & (nonce[48])) + ((g830) & (g1914) & (g2747) & (!g4972) & (g4973) & (!nonce[48])) + ((g830) & (g1914) & (g2747) & (!g4972) & (g4973) & (nonce[48])));
	assign g4975 = (((!g3245) & (!g3310) & (g3265) & (g3312) & (g4862)) + ((!g3245) & (g3310) & (!g3265) & (g3312) & (!g4862)) + ((!g3245) & (g3310) & (!g3265) & (g3312) & (g4862)) + ((!g3245) & (g3310) & (g3265) & (!g3312) & (g4862)) + ((!g3245) & (g3310) & (g3265) & (g3312) & (!g4862)) + ((!g3245) & (g3310) & (g3265) & (g3312) & (g4862)) + ((g3245) & (!g3310) & (!g3265) & (g3312) & (g4862)) + ((g3245) & (!g3310) & (g3265) & (g3312) & (!g4862)) + ((g3245) & (!g3310) & (g3265) & (g3312) & (g4862)) + ((g3245) & (g3310) & (!g3265) & (!g3312) & (g4862)) + ((g3245) & (g3310) & (!g3265) & (g3312) & (!g4862)) + ((g3245) & (g3310) & (!g3265) & (g3312) & (g4862)) + ((g3245) & (g3310) & (g3265) & (!g3312) & (!g4862)) + ((g3245) & (g3310) & (g3265) & (!g3312) & (g4862)) + ((g3245) & (g3310) & (g3265) & (g3312) & (!g4862)) + ((g3245) & (g3310) & (g3265) & (g3312) & (g4862)));
	assign g4976 = (((!g3245) & (!g3310) & (!g3265) & (!g3312) & (!g4862) & (!g5719)) + ((!g3245) & (!g3310) & (!g3265) & (!g3312) & (g4862) & (!g5719)) + ((!g3245) & (!g3310) & (!g3265) & (g3312) & (!g4862) & (!g5719)) + ((!g3245) & (!g3310) & (!g3265) & (g3312) & (g4862) & (!g5719)) + ((!g3245) & (!g3310) & (g3265) & (!g3312) & (!g4862) & (!g5719)) + ((!g3245) & (!g3310) & (g3265) & (!g3312) & (g4862) & (!g5719)) + ((!g3245) & (!g3310) & (g3265) & (g3312) & (!g4862) & (!g5719)) + ((!g3245) & (!g3310) & (g3265) & (g3312) & (g4862) & (g5719)) + ((!g3245) & (g3310) & (!g3265) & (!g3312) & (!g4862) & (!g5719)) + ((!g3245) & (g3310) & (!g3265) & (!g3312) & (g4862) & (!g5719)) + ((!g3245) & (g3310) & (!g3265) & (g3312) & (!g4862) & (g5719)) + ((!g3245) & (g3310) & (!g3265) & (g3312) & (g4862) & (g5719)) + ((!g3245) & (g3310) & (g3265) & (!g3312) & (!g4862) & (!g5719)) + ((!g3245) & (g3310) & (g3265) & (!g3312) & (g4862) & (g5719)) + ((!g3245) & (g3310) & (g3265) & (g3312) & (!g4862) & (g5719)) + ((!g3245) & (g3310) & (g3265) & (g3312) & (g4862) & (g5719)) + ((g3245) & (!g3310) & (!g3265) & (!g3312) & (!g4862) & (!g5719)) + ((g3245) & (!g3310) & (!g3265) & (!g3312) & (g4862) & (!g5719)) + ((g3245) & (!g3310) & (!g3265) & (g3312) & (!g4862) & (!g5719)) + ((g3245) & (!g3310) & (!g3265) & (g3312) & (g4862) & (g5719)) + ((g3245) & (!g3310) & (g3265) & (!g3312) & (!g4862) & (!g5719)) + ((g3245) & (!g3310) & (g3265) & (!g3312) & (g4862) & (!g5719)) + ((g3245) & (!g3310) & (g3265) & (g3312) & (!g4862) & (g5719)) + ((g3245) & (!g3310) & (g3265) & (g3312) & (g4862) & (g5719)) + ((g3245) & (g3310) & (!g3265) & (!g3312) & (!g4862) & (!g5719)) + ((g3245) & (g3310) & (!g3265) & (!g3312) & (g4862) & (g5719)) + ((g3245) & (g3310) & (!g3265) & (g3312) & (!g4862) & (g5719)) + ((g3245) & (g3310) & (!g3265) & (g3312) & (g4862) & (g5719)) + ((g3245) & (g3310) & (g3265) & (!g3312) & (!g4862) & (g5719)) + ((g3245) & (g3310) & (g3265) & (!g3312) & (g4862) & (g5719)) + ((g3245) & (g3310) & (g3265) & (g3312) & (!g4862) & (g5719)) + ((g3245) & (g3310) & (g3265) & (g3312) & (g4862) & (g5719)));
	assign g4977 = (((!g3299) & (!g3353) & (!g3307) & (g3356) & (!g4921) & (!g4922)) + ((!g3299) & (!g3353) & (!g3307) & (g3356) & (!g4921) & (g4922)) + ((!g3299) & (!g3353) & (!g3307) & (g3356) & (g4921) & (!g4922)) + ((!g3299) & (!g3353) & (!g3307) & (g3356) & (g4921) & (g4922)) + ((!g3299) & (!g3353) & (g3307) & (!g3356) & (!g4921) & (g4922)) + ((!g3299) & (!g3353) & (g3307) & (!g3356) & (g4921) & (!g4922)) + ((!g3299) & (!g3353) & (g3307) & (!g3356) & (g4921) & (g4922)) + ((!g3299) & (!g3353) & (g3307) & (g3356) & (!g4921) & (!g4922)) + ((!g3299) & (g3353) & (!g3307) & (!g3356) & (!g4921) & (!g4922)) + ((!g3299) & (g3353) & (!g3307) & (!g3356) & (!g4921) & (g4922)) + ((!g3299) & (g3353) & (!g3307) & (!g3356) & (g4921) & (!g4922)) + ((!g3299) & (g3353) & (!g3307) & (!g3356) & (g4921) & (g4922)) + ((!g3299) & (g3353) & (g3307) & (!g3356) & (!g4921) & (!g4922)) + ((!g3299) & (g3353) & (g3307) & (g3356) & (!g4921) & (g4922)) + ((!g3299) & (g3353) & (g3307) & (g3356) & (g4921) & (!g4922)) + ((!g3299) & (g3353) & (g3307) & (g3356) & (g4921) & (g4922)) + ((g3299) & (!g3353) & (!g3307) & (!g3356) & (!g4921) & (g4922)) + ((g3299) & (!g3353) & (!g3307) & (!g3356) & (g4921) & (!g4922)) + ((g3299) & (!g3353) & (!g3307) & (!g3356) & (g4921) & (g4922)) + ((g3299) & (!g3353) & (!g3307) & (g3356) & (!g4921) & (!g4922)) + ((g3299) & (!g3353) & (g3307) & (!g3356) & (!g4921) & (!g4922)) + ((g3299) & (!g3353) & (g3307) & (!g3356) & (!g4921) & (g4922)) + ((g3299) & (!g3353) & (g3307) & (!g3356) & (g4921) & (!g4922)) + ((g3299) & (!g3353) & (g3307) & (!g3356) & (g4921) & (g4922)) + ((g3299) & (g3353) & (!g3307) & (!g3356) & (!g4921) & (!g4922)) + ((g3299) & (g3353) & (!g3307) & (g3356) & (!g4921) & (g4922)) + ((g3299) & (g3353) & (!g3307) & (g3356) & (g4921) & (!g4922)) + ((g3299) & (g3353) & (!g3307) & (g3356) & (g4921) & (g4922)) + ((g3299) & (g3353) & (g3307) & (g3356) & (!g4921) & (!g4922)) + ((g3299) & (g3353) & (g3307) & (g3356) & (!g4921) & (g4922)) + ((g3299) & (g3353) & (g3307) & (g3356) & (g4921) & (!g4922)) + ((g3299) & (g3353) & (g3307) & (g3356) & (g4921) & (g4922)));
	assign g4978 = (((g830) & (!g1914) & (!g2752) & (!g4976) & (g4977)) + ((g830) & (!g1914) & (!g2752) & (g4976) & (g4977)) + ((g830) & (!g1914) & (g2752) & (!g4976) & (!g4977)) + ((g830) & (!g1914) & (g2752) & (g4976) & (!g4977)) + ((g830) & (g1914) & (!g2752) & (g4976) & (!g4977)) + ((g830) & (g1914) & (!g2752) & (g4976) & (g4977)) + ((g830) & (g1914) & (g2752) & (!g4976) & (!g4977)) + ((g830) & (g1914) & (g2752) & (!g4976) & (g4977)));
	assign g4979 = (((!g1540) & (!g3513) & (!g3514) & (g2916)) + ((!g1540) & (!g3513) & (g3514) & (!g2916)) + ((!g1540) & (g3513) & (!g3514) & (!g2916)) + ((!g1540) & (g3513) & (g3514) & (!g2916)) + ((g1540) & (!g3513) & (!g3514) & (!g2916)) + ((g1540) & (!g3513) & (g3514) & (g2916)) + ((g1540) & (g3513) & (!g3514) & (g2916)) + ((g1540) & (g3513) & (g3514) & (g2916)));
	assign g4980 = (((!g2932) & (!g2979) & (!g3530) & (g3531)) + ((!g2932) & (!g2979) & (g3530) & (!g3531)) + ((!g2932) & (!g2979) & (g3530) & (g3531)) + ((!g2932) & (g2979) & (!g3530) & (!g3531)) + ((g2932) & (!g2979) & (!g3530) & (!g3531)) + ((g2932) & (g2979) & (!g3530) & (g3531)) + ((g2932) & (g2979) & (g3530) & (!g3531)) + ((g2932) & (g2979) & (g3530) & (g3531)));
	assign g4981 = (((!g830) & (!g1914) & (!g2758) & (!g4979) & (!g4980) & (key[62])) + ((!g830) & (!g1914) & (!g2758) & (!g4979) & (g4980) & (key[62])) + ((!g830) & (!g1914) & (!g2758) & (g4979) & (!g4980) & (key[62])) + ((!g830) & (!g1914) & (!g2758) & (g4979) & (g4980) & (key[62])) + ((!g830) & (!g1914) & (g2758) & (!g4979) & (!g4980) & (key[62])) + ((!g830) & (!g1914) & (g2758) & (!g4979) & (g4980) & (key[62])) + ((!g830) & (!g1914) & (g2758) & (g4979) & (!g4980) & (key[62])) + ((!g830) & (!g1914) & (g2758) & (g4979) & (g4980) & (key[62])) + ((!g830) & (g1914) & (!g2758) & (!g4979) & (!g4980) & (key[62])) + ((!g830) & (g1914) & (!g2758) & (!g4979) & (g4980) & (key[62])) + ((!g830) & (g1914) & (!g2758) & (g4979) & (!g4980) & (key[62])) + ((!g830) & (g1914) & (!g2758) & (g4979) & (g4980) & (key[62])) + ((!g830) & (g1914) & (g2758) & (!g4979) & (!g4980) & (key[62])) + ((!g830) & (g1914) & (g2758) & (!g4979) & (g4980) & (key[62])) + ((!g830) & (g1914) & (g2758) & (g4979) & (!g4980) & (key[62])) + ((!g830) & (g1914) & (g2758) & (g4979) & (g4980) & (key[62])) + ((g830) & (!g1914) & (!g2758) & (!g4979) & (g4980) & (!key[62])) + ((g830) & (!g1914) & (!g2758) & (!g4979) & (g4980) & (key[62])) + ((g830) & (!g1914) & (!g2758) & (g4979) & (g4980) & (!key[62])) + ((g830) & (!g1914) & (!g2758) & (g4979) & (g4980) & (key[62])) + ((g830) & (!g1914) & (g2758) & (!g4979) & (!g4980) & (!key[62])) + ((g830) & (!g1914) & (g2758) & (!g4979) & (!g4980) & (key[62])) + ((g830) & (!g1914) & (g2758) & (g4979) & (!g4980) & (!key[62])) + ((g830) & (!g1914) & (g2758) & (g4979) & (!g4980) & (key[62])) + ((g830) & (g1914) & (!g2758) & (g4979) & (!g4980) & (!key[62])) + ((g830) & (g1914) & (!g2758) & (g4979) & (!g4980) & (key[62])) + ((g830) & (g1914) & (!g2758) & (g4979) & (g4980) & (!key[62])) + ((g830) & (g1914) & (!g2758) & (g4979) & (g4980) & (key[62])) + ((g830) & (g1914) & (g2758) & (!g4979) & (!g4980) & (!key[62])) + ((g830) & (g1914) & (g2758) & (!g4979) & (!g4980) & (key[62])) + ((g830) & (g1914) & (g2758) & (!g4979) & (g4980) & (!key[62])) + ((g830) & (g1914) & (g2758) & (!g4979) & (g4980) & (key[62])));
	assign g4982 = (((!g2098) & (!g2129) & (!g2718) & (g2764) & (!g4928)) + ((!g2098) & (!g2129) & (!g2718) & (g2764) & (g4928)) + ((!g2098) & (!g2129) & (g2718) & (!g2764) & (g4928)) + ((!g2098) & (!g2129) & (g2718) & (g2764) & (!g4928)) + ((!g2098) & (g2129) & (!g2718) & (!g2764) & (!g4928)) + ((!g2098) & (g2129) & (!g2718) & (!g2764) & (g4928)) + ((!g2098) & (g2129) & (g2718) & (!g2764) & (!g4928)) + ((!g2098) & (g2129) & (g2718) & (g2764) & (g4928)) + ((g2098) & (!g2129) & (!g2718) & (!g2764) & (g4928)) + ((g2098) & (!g2129) & (!g2718) & (g2764) & (!g4928)) + ((g2098) & (!g2129) & (g2718) & (!g2764) & (!g4928)) + ((g2098) & (!g2129) & (g2718) & (!g2764) & (g4928)) + ((g2098) & (g2129) & (!g2718) & (!g2764) & (!g4928)) + ((g2098) & (g2129) & (!g2718) & (g2764) & (g4928)) + ((g2098) & (g2129) & (g2718) & (g2764) & (!g4928)) + ((g2098) & (g2129) & (g2718) & (g2764) & (g4928)));
	assign g4983 = (((!g1914) & (!g3044) & (!g3067) & (!g3774) & (!g4982)) + ((!g1914) & (!g3044) & (!g3067) & (!g3774) & (g4982)) + ((!g1914) & (!g3044) & (g3067) & (g3774) & (!g4982)) + ((!g1914) & (!g3044) & (g3067) & (g3774) & (g4982)) + ((!g1914) & (g3044) & (!g3067) & (g3774) & (!g4982)) + ((!g1914) & (g3044) & (!g3067) & (g3774) & (g4982)) + ((!g1914) & (g3044) & (g3067) & (!g3774) & (!g4982)) + ((!g1914) & (g3044) & (g3067) & (!g3774) & (g4982)) + ((g1914) & (!g3044) & (!g3067) & (!g3774) & (g4982)) + ((g1914) & (!g3044) & (!g3067) & (g3774) & (g4982)) + ((g1914) & (!g3044) & (g3067) & (!g3774) & (g4982)) + ((g1914) & (!g3044) & (g3067) & (g3774) & (g4982)) + ((g1914) & (g3044) & (!g3067) & (!g3774) & (g4982)) + ((g1914) & (g3044) & (!g3067) & (g3774) & (g4982)) + ((g1914) & (g3044) & (g3067) & (!g3774) & (g4982)) + ((g1914) & (g3044) & (g3067) & (g3774) & (g4982)));
	assign g4984 = (((!g830) & (!g2759) & (!g4983) & (key[94])) + ((!g830) & (!g2759) & (g4983) & (key[94])) + ((!g830) & (g2759) & (!g4983) & (key[94])) + ((!g830) & (g2759) & (g4983) & (key[94])) + ((g830) & (!g2759) & (g4983) & (!key[94])) + ((g830) & (!g2759) & (g4983) & (key[94])) + ((g830) & (g2759) & (!g4983) & (!key[94])) + ((g830) & (g2759) & (!g4983) & (key[94])));
	assign g4985 = (((!g3423) & (g3424)) + ((g3423) & (!g3424)) + ((g3423) & (g3424)));
	assign g4986 = (((!g3406) & (g3407)) + ((g3406) & (!g3407)) + ((g3406) & (g3407)));
	assign g8323 = (((!g5560) & (g5626) & (!g4987)) + ((!g5560) & (g5626) & (g4987)) + ((g5560) & (!g5626) & (g4987)) + ((g5560) & (g5626) & (g4987)));
	assign g4988 = (((!g830) & (!g2760) & (!g6284) & (g4987)) + ((!g830) & (!g2760) & (g6284) & (g4987)) + ((!g830) & (g2760) & (!g6284) & (g4987)) + ((!g830) & (g2760) & (g6284) & (g4987)) + ((g830) & (!g2760) & (g6284) & (!g4987)) + ((g830) & (!g2760) & (g6284) & (g4987)) + ((g830) & (g2760) & (!g6284) & (!g4987)) + ((g830) & (g2760) & (!g6284) & (g4987)));
	assign g4989 = (((!g2100) & (!g2133) & (!g2690) & (g2774) & (!g4934)) + ((!g2100) & (!g2133) & (!g2690) & (g2774) & (g4934)) + ((!g2100) & (!g2133) & (g2690) & (!g2774) & (g4934)) + ((!g2100) & (!g2133) & (g2690) & (g2774) & (!g4934)) + ((!g2100) & (g2133) & (!g2690) & (!g2774) & (!g4934)) + ((!g2100) & (g2133) & (!g2690) & (!g2774) & (g4934)) + ((!g2100) & (g2133) & (g2690) & (!g2774) & (!g4934)) + ((!g2100) & (g2133) & (g2690) & (g2774) & (g4934)) + ((g2100) & (!g2133) & (!g2690) & (!g2774) & (g4934)) + ((g2100) & (!g2133) & (!g2690) & (g2774) & (!g4934)) + ((g2100) & (!g2133) & (g2690) & (!g2774) & (!g4934)) + ((g2100) & (!g2133) & (g2690) & (!g2774) & (g4934)) + ((g2100) & (g2133) & (!g2690) & (!g2774) & (!g4934)) + ((g2100) & (g2133) & (!g2690) & (g2774) & (g4934)) + ((g2100) & (g2133) & (g2690) & (g2774) & (!g4934)) + ((g2100) & (g2133) & (g2690) & (g2774) & (g4934)));
	assign g4990 = (((!g1914) & (!g3481) & (!g3061) & (!g3067) & (g4989)) + ((!g1914) & (!g3481) & (!g3061) & (g3067) & (g4989)) + ((!g1914) & (!g3481) & (g3061) & (!g3067) & (g4989)) + ((!g1914) & (!g3481) & (g3061) & (g3067) & (g4989)) + ((!g1914) & (g3481) & (!g3061) & (!g3067) & (g4989)) + ((!g1914) & (g3481) & (!g3061) & (g3067) & (g4989)) + ((!g1914) & (g3481) & (g3061) & (!g3067) & (g4989)) + ((!g1914) & (g3481) & (g3061) & (g3067) & (g4989)) + ((g1914) & (!g3481) & (!g3061) & (!g3067) & (!g4989)) + ((g1914) & (!g3481) & (!g3061) & (!g3067) & (g4989)) + ((g1914) & (!g3481) & (g3061) & (g3067) & (!g4989)) + ((g1914) & (!g3481) & (g3061) & (g3067) & (g4989)) + ((g1914) & (g3481) & (!g3061) & (g3067) & (!g4989)) + ((g1914) & (g3481) & (!g3061) & (g3067) & (g4989)) + ((g1914) & (g3481) & (g3061) & (!g3067) & (!g4989)) + ((g1914) & (g3481) & (g3061) & (!g3067) & (g4989)));
	assign g4991 = (((!g830) & (!g2761) & (!g4990) & (key[190])) + ((!g830) & (!g2761) & (g4990) & (key[190])) + ((!g830) & (g2761) & (!g4990) & (key[190])) + ((!g830) & (g2761) & (g4990) & (key[190])) + ((g830) & (!g2761) & (g4990) & (!key[190])) + ((g830) & (!g2761) & (g4990) & (key[190])) + ((g830) & (g2761) & (!g4990) & (!key[190])) + ((g830) & (g2761) & (!g4990) & (key[190])));
	assign g4992 = (((!g2110) & (g2125) & (g3638)) + ((g2110) & (!g2125) & (g3638)) + ((g2110) & (g2125) & (!g3638)) + ((g2110) & (g2125) & (g3638)));
	assign g4993 = (((!g2156) & (!g2162) & (g4992)) + ((!g2156) & (g2162) & (!g4992)) + ((g2156) & (!g2162) & (!g4992)) + ((g2156) & (g2162) & (g4992)));
	assign g4994 = (((!g830) & (!g2764) & (!g6273) & (key[17])) + ((!g830) & (!g2764) & (g6273) & (key[17])) + ((!g830) & (g2764) & (!g6273) & (key[17])) + ((!g830) & (g2764) & (g6273) & (key[17])) + ((g830) & (!g2764) & (g6273) & (!key[17])) + ((g830) & (!g2764) & (g6273) & (key[17])) + ((g830) & (g2764) & (!g6273) & (!key[17])) + ((g830) & (g2764) & (!g6273) & (key[17])));
	assign g4995 = (((!g2760) & (!g2793) & (!g3342) & (g3372) & (!g4940)) + ((!g2760) & (!g2793) & (!g3342) & (g3372) & (g4940)) + ((!g2760) & (!g2793) & (g3342) & (!g3372) & (g4940)) + ((!g2760) & (!g2793) & (g3342) & (g3372) & (!g4940)) + ((!g2760) & (g2793) & (!g3342) & (!g3372) & (!g4940)) + ((!g2760) & (g2793) & (!g3342) & (!g3372) & (g4940)) + ((!g2760) & (g2793) & (g3342) & (!g3372) & (!g4940)) + ((!g2760) & (g2793) & (g3342) & (g3372) & (g4940)) + ((g2760) & (!g2793) & (!g3342) & (!g3372) & (g4940)) + ((g2760) & (!g2793) & (!g3342) & (g3372) & (!g4940)) + ((g2760) & (!g2793) & (g3342) & (!g3372) & (!g4940)) + ((g2760) & (!g2793) & (g3342) & (!g3372) & (g4940)) + ((g2760) & (g2793) & (!g3342) & (!g3372) & (!g4940)) + ((g2760) & (g2793) & (!g3342) & (g3372) & (g4940)) + ((g2760) & (g2793) & (g3342) & (g3372) & (!g4940)) + ((g2760) & (g2793) & (g3342) & (g3372) & (g4940)));
	assign g4996 = (((!g2678) & (!g2758) & (g3303) & (g3333) & (!g4887) & (g4888)) + ((!g2678) & (!g2758) & (g3303) & (g3333) & (g4887) & (!g4888)) + ((!g2678) & (!g2758) & (g3303) & (g3333) & (g4887) & (g4888)) + ((!g2678) & (g2758) & (!g3303) & (g3333) & (!g4887) & (!g4888)) + ((!g2678) & (g2758) & (!g3303) & (g3333) & (!g4887) & (g4888)) + ((!g2678) & (g2758) & (!g3303) & (g3333) & (g4887) & (!g4888)) + ((!g2678) & (g2758) & (!g3303) & (g3333) & (g4887) & (g4888)) + ((!g2678) & (g2758) & (g3303) & (!g3333) & (!g4887) & (g4888)) + ((!g2678) & (g2758) & (g3303) & (!g3333) & (g4887) & (!g4888)) + ((!g2678) & (g2758) & (g3303) & (!g3333) & (g4887) & (g4888)) + ((!g2678) & (g2758) & (g3303) & (g3333) & (!g4887) & (!g4888)) + ((!g2678) & (g2758) & (g3303) & (g3333) & (!g4887) & (g4888)) + ((!g2678) & (g2758) & (g3303) & (g3333) & (g4887) & (!g4888)) + ((!g2678) & (g2758) & (g3303) & (g3333) & (g4887) & (g4888)) + ((g2678) & (!g2758) & (!g3303) & (g3333) & (!g4887) & (g4888)) + ((g2678) & (!g2758) & (!g3303) & (g3333) & (g4887) & (!g4888)) + ((g2678) & (!g2758) & (!g3303) & (g3333) & (g4887) & (g4888)) + ((g2678) & (!g2758) & (g3303) & (g3333) & (!g4887) & (!g4888)) + ((g2678) & (!g2758) & (g3303) & (g3333) & (!g4887) & (g4888)) + ((g2678) & (!g2758) & (g3303) & (g3333) & (g4887) & (!g4888)) + ((g2678) & (!g2758) & (g3303) & (g3333) & (g4887) & (g4888)) + ((g2678) & (g2758) & (!g3303) & (!g3333) & (!g4887) & (g4888)) + ((g2678) & (g2758) & (!g3303) & (!g3333) & (g4887) & (!g4888)) + ((g2678) & (g2758) & (!g3303) & (!g3333) & (g4887) & (g4888)) + ((g2678) & (g2758) & (!g3303) & (g3333) & (!g4887) & (!g4888)) + ((g2678) & (g2758) & (!g3303) & (g3333) & (!g4887) & (g4888)) + ((g2678) & (g2758) & (!g3303) & (g3333) & (g4887) & (!g4888)) + ((g2678) & (g2758) & (!g3303) & (g3333) & (g4887) & (g4888)) + ((g2678) & (g2758) & (g3303) & (!g3333) & (!g4887) & (!g4888)) + ((g2678) & (g2758) & (g3303) & (!g3333) & (!g4887) & (g4888)) + ((g2678) & (g2758) & (g3303) & (!g3333) & (g4887) & (!g4888)) + ((g2678) & (g2758) & (g3303) & (!g3333) & (g4887) & (g4888)) + ((g2678) & (g2758) & (g3303) & (g3333) & (!g4887) & (!g4888)) + ((g2678) & (g2758) & (g3303) & (g3333) & (!g4887) & (g4888)) + ((g2678) & (g2758) & (g3303) & (g3333) & (g4887) & (!g4888)) + ((g2678) & (g2758) & (g3303) & (g3333) & (g4887) & (g4888)));
	assign g4997 = (((!g1982) & (g2112) & (g3654)) + ((g1982) & (!g2112) & (g3654)) + ((g1982) & (g2112) & (!g3654)) + ((g1982) & (g2112) & (g3654)));
	assign g4998 = (((!g1984) & (!g2167) & (g4997)) + ((!g1984) & (g2167) & (!g4997)) + ((g1984) & (!g2167) & (!g4997)) + ((g1984) & (g2167) & (g4997)));
	assign g8324 = (((!g5560) & (g5627) & (!g4999)) + ((!g5560) & (g5627) & (g4999)) + ((g5560) & (!g5627) & (g4999)) + ((g5560) & (g5627) & (g4999)));
	assign g5000 = (((!g830) & (!g2770) & (!g6255) & (g4999)) + ((!g830) & (!g2770) & (g6255) & (g4999)) + ((!g830) & (g2770) & (!g6255) & (g4999)) + ((!g830) & (g2770) & (g6255) & (g4999)) + ((g830) & (!g2770) & (g6255) & (!g4999)) + ((g830) & (!g2770) & (g6255) & (g4999)) + ((g830) & (g2770) & (!g6255) & (!g4999)) + ((g830) & (g2770) & (!g6255) & (g4999)));
	assign g5001 = (((!g1945) & (g2120) & (g3795)) + ((g1945) & (!g2120) & (g3795)) + ((g1945) & (g2120) & (!g3795)) + ((g1945) & (g2120) & (g3795)));
	assign g5002 = (((!g1947) & (!g2170) & (g5001)) + ((!g1947) & (g2170) & (!g5001)) + ((g1947) & (!g2170) & (!g5001)) + ((g1947) & (g2170) & (g5001)));
	assign g5003 = (((!g830) & (!g2772) & (!g6244) & (key[145])) + ((!g830) & (!g2772) & (g6244) & (key[145])) + ((!g830) & (g2772) & (!g6244) & (key[145])) + ((!g830) & (g2772) & (g6244) & (key[145])) + ((g830) & (!g2772) & (g6244) & (!key[145])) + ((g830) & (!g2772) & (g6244) & (key[145])) + ((g830) & (g2772) & (!g6244) & (!key[145])) + ((g830) & (g2772) & (!g6244) & (key[145])));
	assign g5004 = (((!g3430) & (g2116) & (g2120)) + ((g3430) & (!g2116) & (g2120)) + ((g3430) & (g2116) & (!g2120)) + ((g3430) & (g2116) & (g2120)));
	assign g5005 = (((!g5004) & (!g2147) & (g2170)) + ((!g5004) & (g2147) & (!g2170)) + ((g5004) & (!g2147) & (!g2170)) + ((g5004) & (g2147) & (g2170)));
	assign g5006 = (((!g830) & (!g2774) & (!g6233) & (key[113])) + ((!g830) & (!g2774) & (g6233) & (key[113])) + ((!g830) & (g2774) & (!g6233) & (key[113])) + ((!g830) & (g2774) & (g6233) & (key[113])) + ((g830) & (!g2774) & (g6233) & (!key[113])) + ((g830) & (!g2774) & (g6233) & (key[113])) + ((g830) & (g2774) & (!g6233) & (!key[113])) + ((g830) & (g2774) & (!g6233) & (key[113])));
	assign g5007 = (((!g1944) & (g2123) & (g3572)) + ((g1944) & (!g2123) & (g3572)) + ((g1944) & (g2123) & (!g3572)) + ((g1944) & (g2123) & (g3572)));
	assign g5008 = (((!g1946) & (!g2150) & (g5007)) + ((!g1946) & (g2150) & (!g5007)) + ((g1946) & (!g2150) & (!g5007)) + ((g1946) & (g2150) & (g5007)));
	assign g5009 = (((!g830) & (!g2776) & (!g6222) & (nonce[17])) + ((!g830) & (!g2776) & (g6222) & (nonce[17])) + ((!g830) & (g2776) & (!g6222) & (nonce[17])) + ((!g830) & (g2776) & (g6222) & (nonce[17])) + ((g830) & (!g2776) & (g6222) & (!nonce[17])) + ((g830) & (!g2776) & (g6222) & (nonce[17])) + ((g830) & (g2776) & (!g6222) & (!nonce[17])) + ((g830) & (g2776) & (!g6222) & (nonce[17])));
	assign g5010 = (((!g3323) & (!g3376) & (!g3356) & (g3382) & (!g4961)) + ((!g3323) & (!g3376) & (!g3356) & (g3382) & (g4961)) + ((!g3323) & (!g3376) & (g3356) & (!g3382) & (g4961)) + ((!g3323) & (!g3376) & (g3356) & (g3382) & (!g4961)) + ((!g3323) & (g3376) & (!g3356) & (!g3382) & (!g4961)) + ((!g3323) & (g3376) & (!g3356) & (!g3382) & (g4961)) + ((!g3323) & (g3376) & (g3356) & (!g3382) & (!g4961)) + ((!g3323) & (g3376) & (g3356) & (g3382) & (g4961)) + ((g3323) & (!g3376) & (!g3356) & (!g3382) & (g4961)) + ((g3323) & (!g3376) & (!g3356) & (g3382) & (!g4961)) + ((g3323) & (!g3376) & (g3356) & (!g3382) & (!g4961)) + ((g3323) & (!g3376) & (g3356) & (!g3382) & (g4961)) + ((g3323) & (g3376) & (!g3356) & (!g3382) & (!g4961)) + ((g3323) & (g3376) & (!g3356) & (g3382) & (g4961)) + ((g3323) & (g3376) & (g3356) & (g3382) & (!g4961)) + ((g3323) & (g3376) & (g3356) & (g3382) & (g4961)));
	assign g5011 = (((!g3291) & (!g3339) & (g3312) & (g3348) & (!g4904) & (g4905)) + ((!g3291) & (!g3339) & (g3312) & (g3348) & (g4904) & (!g4905)) + ((!g3291) & (!g3339) & (g3312) & (g3348) & (g4904) & (g4905)) + ((!g3291) & (g3339) & (!g3312) & (g3348) & (!g4904) & (!g4905)) + ((!g3291) & (g3339) & (!g3312) & (g3348) & (!g4904) & (g4905)) + ((!g3291) & (g3339) & (!g3312) & (g3348) & (g4904) & (!g4905)) + ((!g3291) & (g3339) & (!g3312) & (g3348) & (g4904) & (g4905)) + ((!g3291) & (g3339) & (g3312) & (!g3348) & (!g4904) & (g4905)) + ((!g3291) & (g3339) & (g3312) & (!g3348) & (g4904) & (!g4905)) + ((!g3291) & (g3339) & (g3312) & (!g3348) & (g4904) & (g4905)) + ((!g3291) & (g3339) & (g3312) & (g3348) & (!g4904) & (!g4905)) + ((!g3291) & (g3339) & (g3312) & (g3348) & (!g4904) & (g4905)) + ((!g3291) & (g3339) & (g3312) & (g3348) & (g4904) & (!g4905)) + ((!g3291) & (g3339) & (g3312) & (g3348) & (g4904) & (g4905)) + ((g3291) & (!g3339) & (!g3312) & (g3348) & (!g4904) & (g4905)) + ((g3291) & (!g3339) & (!g3312) & (g3348) & (g4904) & (!g4905)) + ((g3291) & (!g3339) & (!g3312) & (g3348) & (g4904) & (g4905)) + ((g3291) & (!g3339) & (g3312) & (g3348) & (!g4904) & (!g4905)) + ((g3291) & (!g3339) & (g3312) & (g3348) & (!g4904) & (g4905)) + ((g3291) & (!g3339) & (g3312) & (g3348) & (g4904) & (!g4905)) + ((g3291) & (!g3339) & (g3312) & (g3348) & (g4904) & (g4905)) + ((g3291) & (g3339) & (!g3312) & (!g3348) & (!g4904) & (g4905)) + ((g3291) & (g3339) & (!g3312) & (!g3348) & (g4904) & (!g4905)) + ((g3291) & (g3339) & (!g3312) & (!g3348) & (g4904) & (g4905)) + ((g3291) & (g3339) & (!g3312) & (g3348) & (!g4904) & (!g4905)) + ((g3291) & (g3339) & (!g3312) & (g3348) & (!g4904) & (g4905)) + ((g3291) & (g3339) & (!g3312) & (g3348) & (g4904) & (!g4905)) + ((g3291) & (g3339) & (!g3312) & (g3348) & (g4904) & (g4905)) + ((g3291) & (g3339) & (g3312) & (!g3348) & (!g4904) & (!g4905)) + ((g3291) & (g3339) & (g3312) & (!g3348) & (!g4904) & (g4905)) + ((g3291) & (g3339) & (g3312) & (!g3348) & (g4904) & (!g4905)) + ((g3291) & (g3339) & (g3312) & (!g3348) & (g4904) & (g4905)) + ((g3291) & (g3339) & (g3312) & (g3348) & (!g4904) & (!g4905)) + ((g3291) & (g3339) & (g3312) & (g3348) & (!g4904) & (g4905)) + ((g3291) & (g3339) & (g3312) & (g3348) & (g4904) & (!g4905)) + ((g3291) & (g3339) & (g3312) & (g3348) & (g4904) & (g4905)));
	assign g5012 = (((!g2314) & (!g2326) & (!g3815)) + ((!g2314) & (g2326) & (g3815)) + ((g2314) & (!g2326) & (g3815)) + ((g2314) & (g2326) & (!g3815)));
	assign g5013 = (((!g1959) & (!g2340) & (!g3832)) + ((!g1959) & (g2340) & (g3832)) + ((g1959) & (!g2340) & (g3832)) + ((g1959) & (g2340) & (!g3832)));
	assign g5014 = (((!g830) & (!g1914) & (!g2780) & (!g5012) & (!g5013) & (nonce[49])) + ((!g830) & (!g1914) & (!g2780) & (!g5012) & (g5013) & (nonce[49])) + ((!g830) & (!g1914) & (!g2780) & (g5012) & (!g5013) & (nonce[49])) + ((!g830) & (!g1914) & (!g2780) & (g5012) & (g5013) & (nonce[49])) + ((!g830) & (!g1914) & (g2780) & (!g5012) & (!g5013) & (nonce[49])) + ((!g830) & (!g1914) & (g2780) & (!g5012) & (g5013) & (nonce[49])) + ((!g830) & (!g1914) & (g2780) & (g5012) & (!g5013) & (nonce[49])) + ((!g830) & (!g1914) & (g2780) & (g5012) & (g5013) & (nonce[49])) + ((!g830) & (g1914) & (!g2780) & (!g5012) & (!g5013) & (nonce[49])) + ((!g830) & (g1914) & (!g2780) & (!g5012) & (g5013) & (nonce[49])) + ((!g830) & (g1914) & (!g2780) & (g5012) & (!g5013) & (nonce[49])) + ((!g830) & (g1914) & (!g2780) & (g5012) & (g5013) & (nonce[49])) + ((!g830) & (g1914) & (g2780) & (!g5012) & (!g5013) & (nonce[49])) + ((!g830) & (g1914) & (g2780) & (!g5012) & (g5013) & (nonce[49])) + ((!g830) & (g1914) & (g2780) & (g5012) & (!g5013) & (nonce[49])) + ((!g830) & (g1914) & (g2780) & (g5012) & (g5013) & (nonce[49])) + ((g830) & (!g1914) & (!g2780) & (!g5012) & (g5013) & (!nonce[49])) + ((g830) & (!g1914) & (!g2780) & (!g5012) & (g5013) & (nonce[49])) + ((g830) & (!g1914) & (!g2780) & (g5012) & (g5013) & (!nonce[49])) + ((g830) & (!g1914) & (!g2780) & (g5012) & (g5013) & (nonce[49])) + ((g830) & (!g1914) & (g2780) & (!g5012) & (!g5013) & (!nonce[49])) + ((g830) & (!g1914) & (g2780) & (!g5012) & (!g5013) & (nonce[49])) + ((g830) & (!g1914) & (g2780) & (g5012) & (!g5013) & (!nonce[49])) + ((g830) & (!g1914) & (g2780) & (g5012) & (!g5013) & (nonce[49])) + ((g830) & (g1914) & (!g2780) & (g5012) & (!g5013) & (!nonce[49])) + ((g830) & (g1914) & (!g2780) & (g5012) & (!g5013) & (nonce[49])) + ((g830) & (g1914) & (!g2780) & (g5012) & (g5013) & (!nonce[49])) + ((g830) & (g1914) & (!g2780) & (g5012) & (g5013) & (nonce[49])) + ((g830) & (g1914) & (g2780) & (!g5012) & (!g5013) & (!nonce[49])) + ((g830) & (g1914) & (g2780) & (!g5012) & (!g5013) & (nonce[49])) + ((g830) & (g1914) & (g2780) & (!g5012) & (g5013) & (!nonce[49])) + ((g830) & (g1914) & (g2780) & (!g5012) & (g5013) & (nonce[49])));
	assign g5015 = (((!g1983) & (g3588) & (g2125)) + ((g1983) & (!g3588) & (g2125)) + ((g1983) & (g3588) & (!g2125)) + ((g1983) & (g3588) & (g2125)));
	assign g5016 = (((!g1985) & (!g5015) & (g2162)) + ((!g1985) & (g5015) & (!g2162)) + ((g1985) & (!g5015) & (!g2162)) + ((g1985) & (g5015) & (g2162)));
	assign g5017 = (((!g830) & (!g2783) & (!g6205) & (key[241])) + ((!g830) & (!g2783) & (g6205) & (key[241])) + ((!g830) & (g2783) & (!g6205) & (key[241])) + ((!g830) & (g2783) & (g6205) & (key[241])) + ((g830) & (!g2783) & (g6205) & (!key[241])) + ((g830) & (!g2783) & (g6205) & (key[241])) + ((g830) & (g2783) & (!g6205) & (!key[241])) + ((g830) & (g2783) & (!g6205) & (key[241])));
	assign g5018 = (((!g1997) & (!g2340) & (!g3714)) + ((!g1997) & (g2340) & (g3714)) + ((g1997) & (!g2340) & (g3714)) + ((g1997) & (g2340) & (!g3714)));
	assign g5019 = (((!g2323) & (!g2326) & (!g3731)) + ((!g2323) & (g2326) & (g3731)) + ((g2323) & (!g2326) & (g3731)) + ((g2323) & (g2326) & (!g3731)));
	assign g5020 = (((!g830) & (!g1914) & (!g2785) & (!g5018) & (!g5019) & (key[209])) + ((!g830) & (!g1914) & (!g2785) & (!g5018) & (g5019) & (key[209])) + ((!g830) & (!g1914) & (!g2785) & (g5018) & (!g5019) & (key[209])) + ((!g830) & (!g1914) & (!g2785) & (g5018) & (g5019) & (key[209])) + ((!g830) & (!g1914) & (g2785) & (!g5018) & (!g5019) & (key[209])) + ((!g830) & (!g1914) & (g2785) & (!g5018) & (g5019) & (key[209])) + ((!g830) & (!g1914) & (g2785) & (g5018) & (!g5019) & (key[209])) + ((!g830) & (!g1914) & (g2785) & (g5018) & (g5019) & (key[209])) + ((!g830) & (g1914) & (!g2785) & (!g5018) & (!g5019) & (key[209])) + ((!g830) & (g1914) & (!g2785) & (!g5018) & (g5019) & (key[209])) + ((!g830) & (g1914) & (!g2785) & (g5018) & (!g5019) & (key[209])) + ((!g830) & (g1914) & (!g2785) & (g5018) & (g5019) & (key[209])) + ((!g830) & (g1914) & (g2785) & (!g5018) & (!g5019) & (key[209])) + ((!g830) & (g1914) & (g2785) & (!g5018) & (g5019) & (key[209])) + ((!g830) & (g1914) & (g2785) & (g5018) & (!g5019) & (key[209])) + ((!g830) & (g1914) & (g2785) & (g5018) & (g5019) & (key[209])) + ((g830) & (!g1914) & (!g2785) & (!g5018) & (g5019) & (!key[209])) + ((g830) & (!g1914) & (!g2785) & (!g5018) & (g5019) & (key[209])) + ((g830) & (!g1914) & (!g2785) & (g5018) & (g5019) & (!key[209])) + ((g830) & (!g1914) & (!g2785) & (g5018) & (g5019) & (key[209])) + ((g830) & (!g1914) & (g2785) & (!g5018) & (!g5019) & (!key[209])) + ((g830) & (!g1914) & (g2785) & (!g5018) & (!g5019) & (key[209])) + ((g830) & (!g1914) & (g2785) & (g5018) & (!g5019) & (!key[209])) + ((g830) & (!g1914) & (g2785) & (g5018) & (!g5019) & (key[209])) + ((g830) & (g1914) & (!g2785) & (g5018) & (!g5019) & (!key[209])) + ((g830) & (g1914) & (!g2785) & (g5018) & (!g5019) & (key[209])) + ((g830) & (g1914) & (!g2785) & (g5018) & (g5019) & (!key[209])) + ((g830) & (g1914) & (!g2785) & (g5018) & (g5019) & (key[209])) + ((g830) & (g1914) & (g2785) & (!g5018) & (!g5019) & (!key[209])) + ((g830) & (g1914) & (g2785) & (!g5018) & (!g5019) & (key[209])) + ((g830) & (g1914) & (g2785) & (!g5018) & (g5019) & (!key[209])) + ((g830) & (g1914) & (g2785) & (!g5018) & (g5019) & (key[209])));
	assign g5021 = (((!g3336) & (!g3385) & (!g3348) & (g3387) & (!g4975)) + ((!g3336) & (!g3385) & (!g3348) & (g3387) & (g4975)) + ((!g3336) & (!g3385) & (g3348) & (!g3387) & (g4975)) + ((!g3336) & (!g3385) & (g3348) & (g3387) & (!g4975)) + ((!g3336) & (g3385) & (!g3348) & (!g3387) & (!g4975)) + ((!g3336) & (g3385) & (!g3348) & (!g3387) & (g4975)) + ((!g3336) & (g3385) & (g3348) & (!g3387) & (!g4975)) + ((!g3336) & (g3385) & (g3348) & (g3387) & (g4975)) + ((g3336) & (!g3385) & (!g3348) & (!g3387) & (g4975)) + ((g3336) & (!g3385) & (!g3348) & (g3387) & (!g4975)) + ((g3336) & (!g3385) & (g3348) & (!g3387) & (!g4975)) + ((g3336) & (!g3385) & (g3348) & (!g3387) & (g4975)) + ((g3336) & (g3385) & (!g3348) & (!g3387) & (!g4975)) + ((g3336) & (g3385) & (!g3348) & (g3387) & (g4975)) + ((g3336) & (g3385) & (g3348) & (g3387) & (!g4975)) + ((g3336) & (g3385) & (g3348) & (g3387) & (g4975)));
	assign g5022 = (((!g3299) & (!g3353) & (g3307) & (g3356) & (!g4921) & (g4922)) + ((!g3299) & (!g3353) & (g3307) & (g3356) & (g4921) & (!g4922)) + ((!g3299) & (!g3353) & (g3307) & (g3356) & (g4921) & (g4922)) + ((!g3299) & (g3353) & (!g3307) & (g3356) & (!g4921) & (!g4922)) + ((!g3299) & (g3353) & (!g3307) & (g3356) & (!g4921) & (g4922)) + ((!g3299) & (g3353) & (!g3307) & (g3356) & (g4921) & (!g4922)) + ((!g3299) & (g3353) & (!g3307) & (g3356) & (g4921) & (g4922)) + ((!g3299) & (g3353) & (g3307) & (!g3356) & (!g4921) & (g4922)) + ((!g3299) & (g3353) & (g3307) & (!g3356) & (g4921) & (!g4922)) + ((!g3299) & (g3353) & (g3307) & (!g3356) & (g4921) & (g4922)) + ((!g3299) & (g3353) & (g3307) & (g3356) & (!g4921) & (!g4922)) + ((!g3299) & (g3353) & (g3307) & (g3356) & (!g4921) & (g4922)) + ((!g3299) & (g3353) & (g3307) & (g3356) & (g4921) & (!g4922)) + ((!g3299) & (g3353) & (g3307) & (g3356) & (g4921) & (g4922)) + ((g3299) & (!g3353) & (!g3307) & (g3356) & (!g4921) & (g4922)) + ((g3299) & (!g3353) & (!g3307) & (g3356) & (g4921) & (!g4922)) + ((g3299) & (!g3353) & (!g3307) & (g3356) & (g4921) & (g4922)) + ((g3299) & (!g3353) & (g3307) & (g3356) & (!g4921) & (!g4922)) + ((g3299) & (!g3353) & (g3307) & (g3356) & (!g4921) & (g4922)) + ((g3299) & (!g3353) & (g3307) & (g3356) & (g4921) & (!g4922)) + ((g3299) & (!g3353) & (g3307) & (g3356) & (g4921) & (g4922)) + ((g3299) & (g3353) & (!g3307) & (!g3356) & (!g4921) & (g4922)) + ((g3299) & (g3353) & (!g3307) & (!g3356) & (g4921) & (!g4922)) + ((g3299) & (g3353) & (!g3307) & (!g3356) & (g4921) & (g4922)) + ((g3299) & (g3353) & (!g3307) & (g3356) & (!g4921) & (!g4922)) + ((g3299) & (g3353) & (!g3307) & (g3356) & (!g4921) & (g4922)) + ((g3299) & (g3353) & (!g3307) & (g3356) & (g4921) & (!g4922)) + ((g3299) & (g3353) & (!g3307) & (g3356) & (g4921) & (g4922)) + ((g3299) & (g3353) & (g3307) & (!g3356) & (!g4921) & (!g4922)) + ((g3299) & (g3353) & (g3307) & (!g3356) & (!g4921) & (g4922)) + ((g3299) & (g3353) & (g3307) & (!g3356) & (g4921) & (!g4922)) + ((g3299) & (g3353) & (g3307) & (!g3356) & (g4921) & (g4922)) + ((g3299) & (g3353) & (g3307) & (g3356) & (!g4921) & (!g4922)) + ((g3299) & (g3353) & (g3307) & (g3356) & (!g4921) & (g4922)) + ((g3299) & (g3353) & (g3307) & (g3356) & (g4921) & (!g4922)) + ((g3299) & (g3353) & (g3307) & (g3356) & (g4921) & (g4922)));
	assign g5023 = (((!g1540) & (!g3513) & (!g3514) & (!g2916)) + ((!g1540) & (!g3513) & (!g3514) & (g2916)) + ((!g1540) & (!g3513) & (g3514) & (!g2916)) + ((!g1540) & (g3513) & (!g3514) & (!g2916)) + ((!g1540) & (g3513) & (g3514) & (!g2916)) + ((g1540) & (!g3513) & (!g3514) & (!g2916)));
	assign g5024 = (((g1914) & (!g1577) & (!g5023) & (!g3009)) + ((g1914) & (!g1577) & (g5023) & (g3009)) + ((g1914) & (g1577) & (!g5023) & (g3009)) + ((g1914) & (g1577) & (g5023) & (!g3009)));
	assign g5025 = (((!g2932) & (!g2979) & (!g3530) & (!g3531)) + ((!g2932) & (!g2979) & (!g3530) & (g3531)) + ((!g2932) & (!g2979) & (g3530) & (!g3531)) + ((!g2932) & (!g2979) & (g3530) & (g3531)) + ((!g2932) & (g2979) & (!g3530) & (!g3531)) + ((g2932) & (!g2979) & (!g3530) & (!g3531)));
	assign g5026 = (((!g1914) & (!g3003) & (!g3007) & (!g5025)) + ((!g1914) & (!g3003) & (g3007) & (g5025)) + ((!g1914) & (g3003) & (!g3007) & (g5025)) + ((!g1914) & (g3003) & (g3007) & (!g5025)));
	assign g5027 = (((!g830) & (!g2789) & (!g5024) & (!g5026) & (key[63])) + ((!g830) & (!g2789) & (!g5024) & (g5026) & (key[63])) + ((!g830) & (!g2789) & (g5024) & (!g5026) & (key[63])) + ((!g830) & (!g2789) & (g5024) & (g5026) & (key[63])) + ((!g830) & (g2789) & (!g5024) & (!g5026) & (key[63])) + ((!g830) & (g2789) & (!g5024) & (g5026) & (key[63])) + ((!g830) & (g2789) & (g5024) & (!g5026) & (key[63])) + ((!g830) & (g2789) & (g5024) & (g5026) & (key[63])) + ((g830) & (!g2789) & (!g5024) & (g5026) & (!key[63])) + ((g830) & (!g2789) & (!g5024) & (g5026) & (key[63])) + ((g830) & (!g2789) & (g5024) & (!g5026) & (!key[63])) + ((g830) & (!g2789) & (g5024) & (!g5026) & (key[63])) + ((g830) & (!g2789) & (g5024) & (g5026) & (!key[63])) + ((g830) & (!g2789) & (g5024) & (g5026) & (key[63])) + ((g830) & (g2789) & (!g5024) & (!g5026) & (!key[63])) + ((g830) & (g2789) & (!g5024) & (!g5026) & (key[63])));
	assign g5028 = (((!g2177) & (!g2813) & (!g3757)) + ((!g2177) & (g2813) & (g3757)) + ((g2177) & (!g2813) & (g3757)) + ((g2177) & (g2813) & (!g3757)));
	assign g5029 = (((!g1914) & (!g3097) & (!g3775) & (g3093) & (!g5028)) + ((!g1914) & (!g3097) & (!g3775) & (g3093) & (g5028)) + ((!g1914) & (!g3097) & (g3775) & (!g3093) & (!g5028)) + ((!g1914) & (!g3097) & (g3775) & (!g3093) & (g5028)) + ((!g1914) & (g3097) & (!g3775) & (!g3093) & (!g5028)) + ((!g1914) & (g3097) & (!g3775) & (!g3093) & (g5028)) + ((!g1914) & (g3097) & (g3775) & (g3093) & (!g5028)) + ((!g1914) & (g3097) & (g3775) & (g3093) & (g5028)) + ((g1914) & (!g3097) & (!g3775) & (!g3093) & (g5028)) + ((g1914) & (!g3097) & (!g3775) & (g3093) & (g5028)) + ((g1914) & (!g3097) & (g3775) & (!g3093) & (g5028)) + ((g1914) & (!g3097) & (g3775) & (g3093) & (g5028)) + ((g1914) & (g3097) & (!g3775) & (!g3093) & (g5028)) + ((g1914) & (g3097) & (!g3775) & (g3093) & (g5028)) + ((g1914) & (g3097) & (g3775) & (!g3093) & (g5028)) + ((g1914) & (g3097) & (g3775) & (g3093) & (g5028)));
	assign g5030 = (((!g830) & (!g2790) & (!g5029) & (key[95])) + ((!g830) & (!g2790) & (g5029) & (key[95])) + ((!g830) & (g2790) & (!g5029) & (key[95])) + ((!g830) & (g2790) & (g5029) & (key[95])) + ((g830) & (!g2790) & (g5029) & (!key[95])) + ((g830) & (!g2790) & (g5029) & (key[95])) + ((g830) & (g2790) & (!g5029) & (!key[95])) + ((g830) & (g2790) & (!g5029) & (key[95])));
	assign g5031 = (((!g4986) & (!g2932) & (!g2944) & (!g3003) & (g3018)) + ((!g4986) & (!g2932) & (!g2944) & (g3003) & (!g3018)) + ((!g4986) & (!g2932) & (g2944) & (!g3003) & (g3018)) + ((!g4986) & (!g2932) & (g2944) & (g3003) & (!g3018)) + ((!g4986) & (g2932) & (!g2944) & (!g3003) & (g3018)) + ((!g4986) & (g2932) & (!g2944) & (g3003) & (!g3018)) + ((!g4986) & (g2932) & (g2944) & (!g3003) & (!g3018)) + ((!g4986) & (g2932) & (g2944) & (g3003) & (g3018)) + ((g4986) & (!g2932) & (!g2944) & (!g3003) & (g3018)) + ((g4986) & (!g2932) & (!g2944) & (g3003) & (!g3018)) + ((g4986) & (!g2932) & (g2944) & (!g3003) & (!g3018)) + ((g4986) & (!g2932) & (g2944) & (g3003) & (g3018)) + ((g4986) & (g2932) & (!g2944) & (!g3003) & (!g3018)) + ((g4986) & (g2932) & (!g2944) & (g3003) & (g3018)) + ((g4986) & (g2932) & (g2944) & (!g3003) & (!g3018)) + ((g4986) & (g2932) & (g2944) & (g3003) & (g3018)));
	assign g5032 = (((!g1540) & (!g1577) & (!g4985) & (!g2950) & (g2999)) + ((!g1540) & (!g1577) & (!g4985) & (g2950) & (g2999)) + ((!g1540) & (!g1577) & (g4985) & (!g2950) & (g2999)) + ((!g1540) & (!g1577) & (g4985) & (g2950) & (!g2999)) + ((!g1540) & (g1577) & (!g4985) & (!g2950) & (!g2999)) + ((!g1540) & (g1577) & (!g4985) & (g2950) & (!g2999)) + ((!g1540) & (g1577) & (g4985) & (!g2950) & (!g2999)) + ((!g1540) & (g1577) & (g4985) & (g2950) & (g2999)) + ((g1540) & (!g1577) & (!g4985) & (!g2950) & (g2999)) + ((g1540) & (!g1577) & (!g4985) & (g2950) & (!g2999)) + ((g1540) & (!g1577) & (g4985) & (!g2950) & (!g2999)) + ((g1540) & (!g1577) & (g4985) & (g2950) & (!g2999)) + ((g1540) & (g1577) & (!g4985) & (!g2950) & (!g2999)) + ((g1540) & (g1577) & (!g4985) & (g2950) & (g2999)) + ((g1540) & (g1577) & (g4985) & (!g2950) & (g2999)) + ((g1540) & (g1577) & (g4985) & (g2950) & (g2999)));
	assign g8325 = (((!g5560) & (g5628) & (!g5033)) + ((!g5560) & (g5628) & (g5033)) + ((g5560) & (!g5628) & (g5033)) + ((g5560) & (g5628) & (g5033)));
	assign g5034 = (((!g830) & (!g1914) & (!g2793) & (!g5031) & (!g5032) & (g5033)) + ((!g830) & (!g1914) & (!g2793) & (!g5031) & (g5032) & (g5033)) + ((!g830) & (!g1914) & (!g2793) & (g5031) & (!g5032) & (g5033)) + ((!g830) & (!g1914) & (!g2793) & (g5031) & (g5032) & (g5033)) + ((!g830) & (!g1914) & (g2793) & (!g5031) & (!g5032) & (g5033)) + ((!g830) & (!g1914) & (g2793) & (!g5031) & (g5032) & (g5033)) + ((!g830) & (!g1914) & (g2793) & (g5031) & (!g5032) & (g5033)) + ((!g830) & (!g1914) & (g2793) & (g5031) & (g5032) & (g5033)) + ((!g830) & (g1914) & (!g2793) & (!g5031) & (!g5032) & (g5033)) + ((!g830) & (g1914) & (!g2793) & (!g5031) & (g5032) & (g5033)) + ((!g830) & (g1914) & (!g2793) & (g5031) & (!g5032) & (g5033)) + ((!g830) & (g1914) & (!g2793) & (g5031) & (g5032) & (g5033)) + ((!g830) & (g1914) & (g2793) & (!g5031) & (!g5032) & (g5033)) + ((!g830) & (g1914) & (g2793) & (!g5031) & (g5032) & (g5033)) + ((!g830) & (g1914) & (g2793) & (g5031) & (!g5032) & (g5033)) + ((!g830) & (g1914) & (g2793) & (g5031) & (g5032) & (g5033)) + ((g830) & (!g1914) & (!g2793) & (!g5031) & (g5032) & (!g5033)) + ((g830) & (!g1914) & (!g2793) & (!g5031) & (g5032) & (g5033)) + ((g830) & (!g1914) & (!g2793) & (g5031) & (g5032) & (!g5033)) + ((g830) & (!g1914) & (!g2793) & (g5031) & (g5032) & (g5033)) + ((g830) & (!g1914) & (g2793) & (!g5031) & (!g5032) & (!g5033)) + ((g830) & (!g1914) & (g2793) & (!g5031) & (!g5032) & (g5033)) + ((g830) & (!g1914) & (g2793) & (g5031) & (!g5032) & (!g5033)) + ((g830) & (!g1914) & (g2793) & (g5031) & (!g5032) & (g5033)) + ((g830) & (g1914) & (!g2793) & (g5031) & (!g5032) & (!g5033)) + ((g830) & (g1914) & (!g2793) & (g5031) & (!g5032) & (g5033)) + ((g830) & (g1914) & (!g2793) & (g5031) & (g5032) & (!g5033)) + ((g830) & (g1914) & (!g2793) & (g5031) & (g5032) & (g5033)) + ((g830) & (g1914) & (g2793) & (!g5031) & (!g5032) & (!g5033)) + ((g830) & (g1914) & (g2793) & (!g5031) & (!g5032) & (g5033)) + ((g830) & (g1914) & (g2793) & (!g5031) & (g5032) & (!g5033)) + ((g830) & (g1914) & (g2793) & (!g5031) & (g5032) & (g5033)));
	assign g5035 = (((!g2180) & (!g2797) & (!g3495)) + ((!g2180) & (g2797) & (g3495)) + ((g2180) & (!g2797) & (g3495)) + ((g2180) & (g2797) & (!g3495)));
	assign g5036 = (((!g1914) & (!g3482) & (!g3082) & (!g3097) & (g5035)) + ((!g1914) & (!g3482) & (!g3082) & (g3097) & (g5035)) + ((!g1914) & (!g3482) & (g3082) & (!g3097) & (g5035)) + ((!g1914) & (!g3482) & (g3082) & (g3097) & (g5035)) + ((!g1914) & (g3482) & (!g3082) & (!g3097) & (g5035)) + ((!g1914) & (g3482) & (!g3082) & (g3097) & (g5035)) + ((!g1914) & (g3482) & (g3082) & (!g3097) & (g5035)) + ((!g1914) & (g3482) & (g3082) & (g3097) & (g5035)) + ((g1914) & (!g3482) & (!g3082) & (g3097) & (!g5035)) + ((g1914) & (!g3482) & (!g3082) & (g3097) & (g5035)) + ((g1914) & (!g3482) & (g3082) & (!g3097) & (!g5035)) + ((g1914) & (!g3482) & (g3082) & (!g3097) & (g5035)) + ((g1914) & (g3482) & (!g3082) & (!g3097) & (!g5035)) + ((g1914) & (g3482) & (!g3082) & (!g3097) & (g5035)) + ((g1914) & (g3482) & (g3082) & (g3097) & (!g5035)) + ((g1914) & (g3482) & (g3082) & (g3097) & (g5035)));
	assign g5037 = (((!g830) & (!g2794) & (!g5036) & (key[191])) + ((!g830) & (!g2794) & (g5036) & (key[191])) + ((!g830) & (g2794) & (!g5036) & (key[191])) + ((!g830) & (g2794) & (g5036) & (key[191])) + ((g830) & (!g2794) & (g5036) & (!key[191])) + ((g830) & (!g2794) & (g5036) & (key[191])) + ((g830) & (g2794) & (!g5036) & (!key[191])) + ((g830) & (g2794) & (!g5036) & (key[191])));
	assign g5038 = (((!g3450) & (!g3451)));
	assign g5039 = (((!g5004) & (!g2147) & (!g2170) & (!g2196) & (g2200)) + ((!g5004) & (!g2147) & (!g2170) & (g2196) & (!g2200)) + ((!g5004) & (!g2147) & (g2170) & (!g2196) & (g2200)) + ((!g5004) & (!g2147) & (g2170) & (g2196) & (!g2200)) + ((!g5004) & (g2147) & (!g2170) & (!g2196) & (g2200)) + ((!g5004) & (g2147) & (!g2170) & (g2196) & (!g2200)) + ((!g5004) & (g2147) & (g2170) & (!g2196) & (!g2200)) + ((!g5004) & (g2147) & (g2170) & (g2196) & (g2200)) + ((g5004) & (!g2147) & (!g2170) & (!g2196) & (g2200)) + ((g5004) & (!g2147) & (!g2170) & (g2196) & (!g2200)) + ((g5004) & (!g2147) & (g2170) & (!g2196) & (!g2200)) + ((g5004) & (!g2147) & (g2170) & (g2196) & (g2200)) + ((g5004) & (g2147) & (!g2170) & (!g2196) & (!g2200)) + ((g5004) & (g2147) & (!g2170) & (g2196) & (g2200)) + ((g5004) & (g2147) & (g2170) & (!g2196) & (!g2200)) + ((g5004) & (g2147) & (g2170) & (g2196) & (g2200)));
	assign g5040 = (((!g1914) & (!g2004) & (!g1199) & (!g5038) & (!g5039)) + ((!g1914) & (!g2004) & (!g1199) & (!g5038) & (g5039)) + ((!g1914) & (!g2004) & (g1199) & (g5038) & (!g5039)) + ((!g1914) & (!g2004) & (g1199) & (g5038) & (g5039)) + ((!g1914) & (g2004) & (!g1199) & (g5038) & (!g5039)) + ((!g1914) & (g2004) & (!g1199) & (g5038) & (g5039)) + ((!g1914) & (g2004) & (g1199) & (!g5038) & (!g5039)) + ((!g1914) & (g2004) & (g1199) & (!g5038) & (g5039)) + ((g1914) & (!g2004) & (!g1199) & (!g5038) & (g5039)) + ((g1914) & (!g2004) & (!g1199) & (g5038) & (g5039)) + ((g1914) & (!g2004) & (g1199) & (!g5038) & (g5039)) + ((g1914) & (!g2004) & (g1199) & (g5038) & (g5039)) + ((g1914) & (g2004) & (!g1199) & (!g5038) & (g5039)) + ((g1914) & (g2004) & (!g1199) & (g5038) & (g5039)) + ((g1914) & (g2004) & (g1199) & (!g5038) & (g5039)) + ((g1914) & (g2004) & (g1199) & (g5038) & (g5039)));
	assign g5041 = (((!g830) & (!g2797) & (!g5040) & (key[114])) + ((!g830) & (!g2797) & (g5040) & (key[114])) + ((!g830) & (g2797) & (!g5040) & (key[114])) + ((!g830) & (g2797) & (g5040) & (key[114])) + ((g830) & (!g2797) & (g5040) & (!key[114])) + ((g830) & (!g2797) & (g5040) & (key[114])) + ((g830) & (g2797) & (!g5040) & (!key[114])) + ((g830) & (g2797) & (!g5040) & (key[114])));
	assign g5042 = (((!g3560) & (!g3561)));
	assign g5043 = (((!g1946) & (!g1948) & (!g2150) & (g2203) & (!g5007)) + ((!g1946) & (!g1948) & (!g2150) & (g2203) & (g5007)) + ((!g1946) & (!g1948) & (g2150) & (!g2203) & (g5007)) + ((!g1946) & (!g1948) & (g2150) & (g2203) & (!g5007)) + ((!g1946) & (g1948) & (!g2150) & (!g2203) & (!g5007)) + ((!g1946) & (g1948) & (!g2150) & (!g2203) & (g5007)) + ((!g1946) & (g1948) & (g2150) & (!g2203) & (!g5007)) + ((!g1946) & (g1948) & (g2150) & (g2203) & (g5007)) + ((g1946) & (!g1948) & (!g2150) & (!g2203) & (g5007)) + ((g1946) & (!g1948) & (!g2150) & (g2203) & (!g5007)) + ((g1946) & (!g1948) & (g2150) & (!g2203) & (!g5007)) + ((g1946) & (!g1948) & (g2150) & (!g2203) & (g5007)) + ((g1946) & (g1948) & (!g2150) & (!g2203) & (!g5007)) + ((g1946) & (g1948) & (!g2150) & (g2203) & (g5007)) + ((g1946) & (g1948) & (g2150) & (g2203) & (!g5007)) + ((g1946) & (g1948) & (g2150) & (g2203) & (g5007)));
	assign g5044 = (((!g1914) & (!g2468) & (!g5042) & (!g2480) & (g5043)) + ((!g1914) & (!g2468) & (!g5042) & (g2480) & (g5043)) + ((!g1914) & (!g2468) & (g5042) & (!g2480) & (g5043)) + ((!g1914) & (!g2468) & (g5042) & (g2480) & (g5043)) + ((!g1914) & (g2468) & (!g5042) & (!g2480) & (g5043)) + ((!g1914) & (g2468) & (!g5042) & (g2480) & (g5043)) + ((!g1914) & (g2468) & (g5042) & (!g2480) & (g5043)) + ((!g1914) & (g2468) & (g5042) & (g2480) & (g5043)) + ((g1914) & (!g2468) & (!g5042) & (!g2480) & (!g5043)) + ((g1914) & (!g2468) & (!g5042) & (!g2480) & (g5043)) + ((g1914) & (!g2468) & (g5042) & (g2480) & (!g5043)) + ((g1914) & (!g2468) & (g5042) & (g2480) & (g5043)) + ((g1914) & (g2468) & (!g5042) & (g2480) & (!g5043)) + ((g1914) & (g2468) & (!g5042) & (g2480) & (g5043)) + ((g1914) & (g2468) & (g5042) & (!g2480) & (!g5043)) + ((g1914) & (g2468) & (g5042) & (!g2480) & (g5043)));
	assign g5045 = (((!g830) & (!g2807) & (!g5044) & (nonce[18])) + ((!g830) & (!g2807) & (g5044) & (nonce[18])) + ((!g830) & (g2807) & (!g5044) & (nonce[18])) + ((!g830) & (g2807) & (g5044) & (nonce[18])) + ((g830) & (!g2807) & (g5044) & (!nonce[18])) + ((g830) & (!g2807) & (g5044) & (nonce[18])) + ((g830) & (g2807) & (!g5044) & (!nonce[18])) + ((g830) & (g2807) & (!g5044) & (nonce[18])));
	assign g5046 = (((!g3608) & (!g3609)));
	assign g5047 = (((!g1985) & (!g1987) & (!g5015) & (!g2162) & (g2205)) + ((!g1985) & (!g1987) & (!g5015) & (g2162) & (g2205)) + ((!g1985) & (!g1987) & (g5015) & (!g2162) & (g2205)) + ((!g1985) & (!g1987) & (g5015) & (g2162) & (!g2205)) + ((!g1985) & (g1987) & (!g5015) & (!g2162) & (!g2205)) + ((!g1985) & (g1987) & (!g5015) & (g2162) & (!g2205)) + ((!g1985) & (g1987) & (g5015) & (!g2162) & (!g2205)) + ((!g1985) & (g1987) & (g5015) & (g2162) & (g2205)) + ((g1985) & (!g1987) & (!g5015) & (!g2162) & (g2205)) + ((g1985) & (!g1987) & (!g5015) & (g2162) & (!g2205)) + ((g1985) & (!g1987) & (g5015) & (!g2162) & (!g2205)) + ((g1985) & (!g1987) & (g5015) & (g2162) & (!g2205)) + ((g1985) & (g1987) & (!g5015) & (!g2162) & (!g2205)) + ((g1985) & (g1987) & (!g5015) & (g2162) & (g2205)) + ((g1985) & (g1987) & (g5015) & (!g2162) & (g2205)) + ((g1985) & (g1987) & (g5015) & (g2162) & (g2205)));
	assign g5048 = (((!g1914) & (!g2450) & (!g2474) & (!g5046) & (!g5047)) + ((!g1914) & (!g2450) & (!g2474) & (!g5046) & (g5047)) + ((!g1914) & (!g2450) & (g2474) & (g5046) & (!g5047)) + ((!g1914) & (!g2450) & (g2474) & (g5046) & (g5047)) + ((!g1914) & (g2450) & (!g2474) & (g5046) & (!g5047)) + ((!g1914) & (g2450) & (!g2474) & (g5046) & (g5047)) + ((!g1914) & (g2450) & (g2474) & (!g5046) & (!g5047)) + ((!g1914) & (g2450) & (g2474) & (!g5046) & (g5047)) + ((g1914) & (!g2450) & (!g2474) & (!g5046) & (g5047)) + ((g1914) & (!g2450) & (!g2474) & (g5046) & (g5047)) + ((g1914) & (!g2450) & (g2474) & (!g5046) & (g5047)) + ((g1914) & (!g2450) & (g2474) & (g5046) & (g5047)) + ((g1914) & (g2450) & (!g2474) & (!g5046) & (g5047)) + ((g1914) & (g2450) & (!g2474) & (g5046) & (g5047)) + ((g1914) & (g2450) & (g2474) & (!g5046) & (g5047)) + ((g1914) & (g2450) & (g2474) & (g5046) & (g5047)));
	assign g5049 = (((!g830) & (!g2810) & (!g5048) & (key[242])) + ((!g830) & (!g2810) & (g5048) & (key[242])) + ((!g830) & (g2810) & (!g5048) & (key[242])) + ((!g830) & (g2810) & (g5048) & (key[242])) + ((g830) & (!g2810) & (g5048) & (!key[242])) + ((g830) & (!g2810) & (g5048) & (key[242])) + ((g830) & (g2810) & (!g5048) & (!key[242])) + ((g830) & (g2810) & (!g5048) & (key[242])));
	assign g5050 = (((!g3627) & (!g3628)));
	assign g5051 = (((!g2156) & (!g2190) & (!g2162) & (g2205) & (!g4992)) + ((!g2156) & (!g2190) & (!g2162) & (g2205) & (g4992)) + ((!g2156) & (!g2190) & (g2162) & (!g2205) & (g4992)) + ((!g2156) & (!g2190) & (g2162) & (g2205) & (!g4992)) + ((!g2156) & (g2190) & (!g2162) & (!g2205) & (!g4992)) + ((!g2156) & (g2190) & (!g2162) & (!g2205) & (g4992)) + ((!g2156) & (g2190) & (g2162) & (!g2205) & (!g4992)) + ((!g2156) & (g2190) & (g2162) & (g2205) & (g4992)) + ((g2156) & (!g2190) & (!g2162) & (!g2205) & (g4992)) + ((g2156) & (!g2190) & (!g2162) & (g2205) & (!g4992)) + ((g2156) & (!g2190) & (g2162) & (!g2205) & (!g4992)) + ((g2156) & (!g2190) & (g2162) & (!g2205) & (g4992)) + ((g2156) & (g2190) & (!g2162) & (!g2205) & (!g4992)) + ((g2156) & (g2190) & (!g2162) & (g2205) & (g4992)) + ((g2156) & (g2190) & (g2162) & (g2205) & (!g4992)) + ((g2156) & (g2190) & (g2162) & (g2205) & (g4992)));
	assign g5052 = (((!g1914) & (!g1968) & (!g1199) & (!g5050) & (g5051)) + ((!g1914) & (!g1968) & (!g1199) & (g5050) & (g5051)) + ((!g1914) & (!g1968) & (g1199) & (!g5050) & (g5051)) + ((!g1914) & (!g1968) & (g1199) & (g5050) & (g5051)) + ((!g1914) & (g1968) & (!g1199) & (!g5050) & (g5051)) + ((!g1914) & (g1968) & (!g1199) & (g5050) & (g5051)) + ((!g1914) & (g1968) & (g1199) & (!g5050) & (g5051)) + ((!g1914) & (g1968) & (g1199) & (g5050) & (g5051)) + ((g1914) & (!g1968) & (!g1199) & (!g5050) & (!g5051)) + ((g1914) & (!g1968) & (!g1199) & (!g5050) & (g5051)) + ((g1914) & (!g1968) & (g1199) & (g5050) & (!g5051)) + ((g1914) & (!g1968) & (g1199) & (g5050) & (g5051)) + ((g1914) & (g1968) & (!g1199) & (g5050) & (!g5051)) + ((g1914) & (g1968) & (!g1199) & (g5050) & (g5051)) + ((g1914) & (g1968) & (g1199) & (!g5050) & (!g5051)) + ((g1914) & (g1968) & (g1199) & (!g5050) & (g5051)));
	assign g5053 = (((!g830) & (!g2813) & (!g5052) & (key[18])) + ((!g830) & (!g2813) & (g5052) & (key[18])) + ((!g830) & (g2813) & (!g5052) & (key[18])) + ((!g830) & (g2813) & (g5052) & (key[18])) + ((g830) & (!g2813) & (g5052) & (!key[18])) + ((g830) & (!g2813) & (g5052) & (key[18])) + ((g830) & (g2813) & (!g5052) & (!key[18])) + ((g830) & (g2813) & (!g5052) & (key[18])));
	assign g5054 = (((!g3675) & (!g3676)));
	assign g5055 = (((!g1984) & (!g1986) & (!g2167) & (g2192) & (!g4997)) + ((!g1984) & (!g1986) & (!g2167) & (g2192) & (g4997)) + ((!g1984) & (!g1986) & (g2167) & (!g2192) & (g4997)) + ((!g1984) & (!g1986) & (g2167) & (g2192) & (!g4997)) + ((!g1984) & (g1986) & (!g2167) & (!g2192) & (!g4997)) + ((!g1984) & (g1986) & (!g2167) & (!g2192) & (g4997)) + ((!g1984) & (g1986) & (g2167) & (!g2192) & (!g4997)) + ((!g1984) & (g1986) & (g2167) & (g2192) & (g4997)) + ((g1984) & (!g1986) & (!g2167) & (!g2192) & (g4997)) + ((g1984) & (!g1986) & (!g2167) & (g2192) & (!g4997)) + ((g1984) & (!g1986) & (g2167) & (!g2192) & (!g4997)) + ((g1984) & (!g1986) & (g2167) & (!g2192) & (g4997)) + ((g1984) & (g1986) & (!g2167) & (!g2192) & (!g4997)) + ((g1984) & (g1986) & (!g2167) & (g2192) & (g4997)) + ((g1984) & (g1986) & (g2167) & (g2192) & (!g4997)) + ((g1984) & (g1986) & (g2167) & (g2192) & (g4997)));
	assign g5056 = (((!g1914) & (!g2434) & (!g2480) & (!g5054) & (!g5055)) + ((!g1914) & (!g2434) & (!g2480) & (!g5054) & (g5055)) + ((!g1914) & (!g2434) & (g2480) & (g5054) & (!g5055)) + ((!g1914) & (!g2434) & (g2480) & (g5054) & (g5055)) + ((!g1914) & (g2434) & (!g2480) & (g5054) & (!g5055)) + ((!g1914) & (g2434) & (!g2480) & (g5054) & (g5055)) + ((!g1914) & (g2434) & (g2480) & (!g5054) & (!g5055)) + ((!g1914) & (g2434) & (g2480) & (!g5054) & (g5055)) + ((g1914) & (!g2434) & (!g2480) & (!g5054) & (g5055)) + ((g1914) & (!g2434) & (!g2480) & (g5054) & (g5055)) + ((g1914) & (!g2434) & (g2480) & (!g5054) & (g5055)) + ((g1914) & (!g2434) & (g2480) & (g5054) & (g5055)) + ((g1914) & (g2434) & (!g2480) & (!g5054) & (g5055)) + ((g1914) & (g2434) & (!g2480) & (g5054) & (g5055)) + ((g1914) & (g2434) & (g2480) & (!g5054) & (g5055)) + ((g1914) & (g2434) & (g2480) & (g5054) & (g5055)));
	assign g8326 = (((!g5560) & (g5629) & (!g5057)) + ((!g5560) & (g5629) & (g5057)) + ((g5560) & (!g5629) & (g5057)) + ((g5560) & (g5629) & (g5057)));
	assign g5058 = (((!g830) & (!g2816) & (!g5056) & (g5057)) + ((!g830) & (!g2816) & (g5056) & (g5057)) + ((!g830) & (g2816) & (!g5056) & (g5057)) + ((!g830) & (g2816) & (g5056) & (g5057)) + ((g830) & (!g2816) & (g5056) & (!g5057)) + ((g830) & (!g2816) & (g5056) & (g5057)) + ((g830) & (g2816) & (!g5056) & (!g5057)) + ((g830) & (g2816) & (!g5056) & (g5057)));
	assign g5059 = (((!g1997) & (g2340) & (!g3714)) + ((g1997) & (!g2340) & (!g3714)) + ((g1997) & (g2340) & (!g3714)) + ((g1997) & (g2340) & (g3714)));
	assign g5060 = (((g1914) & (!g1999) & (!g2373) & (g5059)) + ((g1914) & (!g1999) & (g2373) & (!g5059)) + ((g1914) & (g1999) & (!g2373) & (!g5059)) + ((g1914) & (g1999) & (g2373) & (g5059)));
	assign g5061 = (((!g2323) & (g2326) & (!g3731)) + ((g2323) & (!g2326) & (!g3731)) + ((g2323) & (g2326) & (!g3731)) + ((g2323) & (g2326) & (g3731)));
	assign g5062 = (((!g1914) & (!g2356) & (!g2364) & (g5061)) + ((!g1914) & (!g2356) & (g2364) & (!g5061)) + ((!g1914) & (g2356) & (!g2364) & (!g5061)) + ((!g1914) & (g2356) & (g2364) & (g5061)));
	assign g5063 = (((!g830) & (!g2822) & (!g5060) & (!g5062) & (key[210])) + ((!g830) & (!g2822) & (!g5060) & (g5062) & (key[210])) + ((!g830) & (!g2822) & (g5060) & (!g5062) & (key[210])) + ((!g830) & (!g2822) & (g5060) & (g5062) & (key[210])) + ((!g830) & (g2822) & (!g5060) & (!g5062) & (key[210])) + ((!g830) & (g2822) & (!g5060) & (g5062) & (key[210])) + ((!g830) & (g2822) & (g5060) & (!g5062) & (key[210])) + ((!g830) & (g2822) & (g5060) & (g5062) & (key[210])) + ((g830) & (!g2822) & (!g5060) & (g5062) & (!key[210])) + ((g830) & (!g2822) & (!g5060) & (g5062) & (key[210])) + ((g830) & (!g2822) & (g5060) & (!g5062) & (!key[210])) + ((g830) & (!g2822) & (g5060) & (!g5062) & (key[210])) + ((g830) & (!g2822) & (g5060) & (g5062) & (!key[210])) + ((g830) & (!g2822) & (g5060) & (g5062) & (key[210])) + ((g830) & (g2822) & (!g5060) & (!g5062) & (!key[210])) + ((g830) & (g2822) & (!g5060) & (!g5062) & (key[210])));
	assign g5064 = (((!g3784) & (!g3785)));
	assign g5065 = (((!g1947) & (!g1949) & (!g2170) & (g2200) & (!g5001)) + ((!g1947) & (!g1949) & (!g2170) & (g2200) & (g5001)) + ((!g1947) & (!g1949) & (g2170) & (!g2200) & (g5001)) + ((!g1947) & (!g1949) & (g2170) & (g2200) & (!g5001)) + ((!g1947) & (g1949) & (!g2170) & (!g2200) & (!g5001)) + ((!g1947) & (g1949) & (!g2170) & (!g2200) & (g5001)) + ((!g1947) & (g1949) & (g2170) & (!g2200) & (!g5001)) + ((!g1947) & (g1949) & (g2170) & (g2200) & (g5001)) + ((g1947) & (!g1949) & (!g2170) & (!g2200) & (g5001)) + ((g1947) & (!g1949) & (!g2170) & (g2200) & (!g5001)) + ((g1947) & (!g1949) & (g2170) & (!g2200) & (!g5001)) + ((g1947) & (!g1949) & (g2170) & (!g2200) & (g5001)) + ((g1947) & (g1949) & (!g2170) & (!g2200) & (!g5001)) + ((g1947) & (g1949) & (!g2170) & (g2200) & (g5001)) + ((g1947) & (g1949) & (g2170) & (g2200) & (!g5001)) + ((g1947) & (g1949) & (g2170) & (g2200) & (g5001)));
	assign g5066 = (((!g1914) & (!g2450) & (!g2456) & (!g5064) & (g5065)) + ((!g1914) & (!g2450) & (!g2456) & (g5064) & (g5065)) + ((!g1914) & (!g2450) & (g2456) & (!g5064) & (g5065)) + ((!g1914) & (!g2450) & (g2456) & (g5064) & (g5065)) + ((!g1914) & (g2450) & (!g2456) & (!g5064) & (g5065)) + ((!g1914) & (g2450) & (!g2456) & (g5064) & (g5065)) + ((!g1914) & (g2450) & (g2456) & (!g5064) & (g5065)) + ((!g1914) & (g2450) & (g2456) & (g5064) & (g5065)) + ((g1914) & (!g2450) & (!g2456) & (!g5064) & (!g5065)) + ((g1914) & (!g2450) & (!g2456) & (!g5064) & (g5065)) + ((g1914) & (!g2450) & (g2456) & (g5064) & (!g5065)) + ((g1914) & (!g2450) & (g2456) & (g5064) & (g5065)) + ((g1914) & (g2450) & (!g2456) & (g5064) & (!g5065)) + ((g1914) & (g2450) & (!g2456) & (g5064) & (g5065)) + ((g1914) & (g2450) & (g2456) & (!g5064) & (!g5065)) + ((g1914) & (g2450) & (g2456) & (!g5064) & (g5065)));
	assign g5067 = (((!g830) & (!g2827) & (!g5066) & (key[146])) + ((!g830) & (!g2827) & (g5066) & (key[146])) + ((!g830) & (g2827) & (!g5066) & (key[146])) + ((!g830) & (g2827) & (g5066) & (key[146])) + ((g830) & (!g2827) & (g5066) & (!key[146])) + ((g830) & (!g2827) & (g5066) & (key[146])) + ((g830) & (g2827) & (!g5066) & (!key[146])) + ((g830) & (g2827) & (!g5066) & (key[146])));
	assign g5068 = (((!g2314) & (g2326) & (!g3815)) + ((g2314) & (!g2326) & (!g3815)) + ((g2314) & (g2326) & (!g3815)) + ((g2314) & (g2326) & (g3815)));
	assign g5069 = (((g1914) & (!g2362) & (!g2364) & (g5068)) + ((g1914) & (!g2362) & (g2364) & (!g5068)) + ((g1914) & (g2362) & (!g2364) & (!g5068)) + ((g1914) & (g2362) & (g2364) & (g5068)));
	assign g5070 = (((!g1959) & (g2340) & (!g3832)) + ((g1959) & (!g2340) & (!g3832)) + ((g1959) & (g2340) & (!g3832)) + ((g1959) & (g2340) & (g3832)));
	assign g5071 = (((!g1914) & (!g1961) & (!g2373) & (g5070)) + ((!g1914) & (!g1961) & (g2373) & (!g5070)) + ((!g1914) & (g1961) & (!g2373) & (!g5070)) + ((!g1914) & (g1961) & (g2373) & (g5070)));
	assign g5072 = (((!g830) & (!g2830) & (!g5069) & (!g5071) & (nonce[50])) + ((!g830) & (!g2830) & (!g5069) & (g5071) & (nonce[50])) + ((!g830) & (!g2830) & (g5069) & (!g5071) & (nonce[50])) + ((!g830) & (!g2830) & (g5069) & (g5071) & (nonce[50])) + ((!g830) & (g2830) & (!g5069) & (!g5071) & (nonce[50])) + ((!g830) & (g2830) & (!g5069) & (g5071) & (nonce[50])) + ((!g830) & (g2830) & (g5069) & (!g5071) & (nonce[50])) + ((!g830) & (g2830) & (g5069) & (g5071) & (nonce[50])) + ((g830) & (!g2830) & (!g5069) & (g5071) & (!nonce[50])) + ((g830) & (!g2830) & (!g5069) & (g5071) & (nonce[50])) + ((g830) & (!g2830) & (g5069) & (!g5071) & (!nonce[50])) + ((g830) & (!g2830) & (g5069) & (!g5071) & (nonce[50])) + ((g830) & (!g2830) & (g5069) & (g5071) & (!nonce[50])) + ((g830) & (!g2830) & (g5069) & (g5071) & (nonce[50])) + ((g830) & (g2830) & (!g5069) & (!g5071) & (!nonce[50])) + ((g830) & (g2830) & (!g5069) & (!g5071) & (nonce[50])));
	assign g5073 = (((!g1968) & (!g1970) & (!g1199) & (g1236) & (!g5050)) + ((!g1968) & (!g1970) & (!g1199) & (g1236) & (g5050)) + ((!g1968) & (!g1970) & (g1199) & (!g1236) & (!g5050)) + ((!g1968) & (!g1970) & (g1199) & (g1236) & (g5050)) + ((!g1968) & (g1970) & (!g1199) & (!g1236) & (!g5050)) + ((!g1968) & (g1970) & (!g1199) & (!g1236) & (g5050)) + ((!g1968) & (g1970) & (g1199) & (!g1236) & (g5050)) + ((!g1968) & (g1970) & (g1199) & (g1236) & (!g5050)) + ((g1968) & (!g1970) & (!g1199) & (!g1236) & (!g5050)) + ((g1968) & (!g1970) & (!g1199) & (g1236) & (g5050)) + ((g1968) & (!g1970) & (g1199) & (!g1236) & (!g5050)) + ((g1968) & (!g1970) & (g1199) & (!g1236) & (g5050)) + ((g1968) & (g1970) & (!g1199) & (!g1236) & (g5050)) + ((g1968) & (g1970) & (!g1199) & (g1236) & (!g5050)) + ((g1968) & (g1970) & (g1199) & (g1236) & (!g5050)) + ((g1968) & (g1970) & (g1199) & (g1236) & (g5050)));
	assign g5074 = (((!g3640) & (!g3641)));
	assign g5075 = (((!g2236) & (!g2242) & (!g5074)) + ((!g2236) & (g2242) & (g5074)) + ((g2236) & (!g2242) & (g5074)) + ((g2236) & (g2242) & (!g5074)));
	assign g5076 = (((!g830) & (!g1914) & (!g2838) & (!g5073) & (!g5075) & (key[19])) + ((!g830) & (!g1914) & (!g2838) & (!g5073) & (g5075) & (key[19])) + ((!g830) & (!g1914) & (!g2838) & (g5073) & (!g5075) & (key[19])) + ((!g830) & (!g1914) & (!g2838) & (g5073) & (g5075) & (key[19])) + ((!g830) & (!g1914) & (g2838) & (!g5073) & (!g5075) & (key[19])) + ((!g830) & (!g1914) & (g2838) & (!g5073) & (g5075) & (key[19])) + ((!g830) & (!g1914) & (g2838) & (g5073) & (!g5075) & (key[19])) + ((!g830) & (!g1914) & (g2838) & (g5073) & (g5075) & (key[19])) + ((!g830) & (g1914) & (!g2838) & (!g5073) & (!g5075) & (key[19])) + ((!g830) & (g1914) & (!g2838) & (!g5073) & (g5075) & (key[19])) + ((!g830) & (g1914) & (!g2838) & (g5073) & (!g5075) & (key[19])) + ((!g830) & (g1914) & (!g2838) & (g5073) & (g5075) & (key[19])) + ((!g830) & (g1914) & (g2838) & (!g5073) & (!g5075) & (key[19])) + ((!g830) & (g1914) & (g2838) & (!g5073) & (g5075) & (key[19])) + ((!g830) & (g1914) & (g2838) & (g5073) & (!g5075) & (key[19])) + ((!g830) & (g1914) & (g2838) & (g5073) & (g5075) & (key[19])) + ((g830) & (!g1914) & (!g2838) & (!g5073) & (g5075) & (!key[19])) + ((g830) & (!g1914) & (!g2838) & (!g5073) & (g5075) & (key[19])) + ((g830) & (!g1914) & (!g2838) & (g5073) & (g5075) & (!key[19])) + ((g830) & (!g1914) & (!g2838) & (g5073) & (g5075) & (key[19])) + ((g830) & (!g1914) & (g2838) & (!g5073) & (!g5075) & (!key[19])) + ((g830) & (!g1914) & (g2838) & (!g5073) & (!g5075) & (key[19])) + ((g830) & (!g1914) & (g2838) & (g5073) & (!g5075) & (!key[19])) + ((g830) & (!g1914) & (g2838) & (g5073) & (!g5075) & (key[19])) + ((g830) & (g1914) & (!g2838) & (g5073) & (!g5075) & (!key[19])) + ((g830) & (g1914) & (!g2838) & (g5073) & (!g5075) & (key[19])) + ((g830) & (g1914) & (!g2838) & (g5073) & (g5075) & (!key[19])) + ((g830) & (g1914) & (!g2838) & (g5073) & (g5075) & (key[19])) + ((g830) & (g1914) & (g2838) & (!g5073) & (!g5075) & (!key[19])) + ((g830) & (g1914) & (g2838) & (!g5073) & (!g5075) & (key[19])) + ((g830) & (g1914) & (g2838) & (!g5073) & (g5075) & (!key[19])) + ((g830) & (g1914) & (g2838) & (!g5073) & (g5075) & (key[19])));
	assign g5077 = (((!g1884) & (!g1977) & (!g1900) & (g2028)) + ((!g1884) & (!g1977) & (g1900) & (g2028)) + ((!g1884) & (g1977) & (!g1900) & (!g2028)) + ((!g1884) & (g1977) & (g1900) & (!g2028)) + ((g1884) & (!g1977) & (!g1900) & (g2028)) + ((g1884) & (!g1977) & (g1900) & (!g2028)) + ((g1884) & (g1977) & (!g1900) & (!g2028)) + ((g1884) & (g1977) & (g1900) & (g2028)));
	assign g5078 = (((!g1890) & (!g1939) & (!g1894) & (g2034)) + ((!g1890) & (!g1939) & (g1894) & (g2034)) + ((!g1890) & (g1939) & (!g1894) & (!g2034)) + ((!g1890) & (g1939) & (g1894) & (!g2034)) + ((g1890) & (!g1939) & (!g1894) & (g2034)) + ((g1890) & (!g1939) & (g1894) & (!g2034)) + ((g1890) & (g1939) & (!g1894) & (!g2034)) + ((g1890) & (g1939) & (g1894) & (g2034)));
	assign g5079 = (((g830) & (!g1914) & (!g2845) & (!g5077) & (g5078)) + ((g830) & (!g1914) & (!g2845) & (g5077) & (g5078)) + ((g830) & (!g1914) & (g2845) & (!g5077) & (!g5078)) + ((g830) & (!g1914) & (g2845) & (g5077) & (!g5078)) + ((g830) & (g1914) & (!g2845) & (g5077) & (!g5078)) + ((g830) & (g1914) & (!g2845) & (g5077) & (g5078)) + ((g830) & (g1914) & (g2845) & (!g5077) & (!g5078)) + ((g830) & (g1914) & (g2845) & (!g5077) & (g5078)));
	assign g5080 = (((!g3656) & (!g3657)));
	assign g5081 = (((!g2434) & (!g2533) & (!g2480) & (g2537) & (!g5054)) + ((!g2434) & (!g2533) & (!g2480) & (g2537) & (g5054)) + ((!g2434) & (!g2533) & (g2480) & (!g2537) & (!g5054)) + ((!g2434) & (!g2533) & (g2480) & (g2537) & (g5054)) + ((!g2434) & (g2533) & (!g2480) & (!g2537) & (!g5054)) + ((!g2434) & (g2533) & (!g2480) & (!g2537) & (g5054)) + ((!g2434) & (g2533) & (g2480) & (!g2537) & (g5054)) + ((!g2434) & (g2533) & (g2480) & (g2537) & (!g5054)) + ((g2434) & (!g2533) & (!g2480) & (!g2537) & (!g5054)) + ((g2434) & (!g2533) & (!g2480) & (g2537) & (g5054)) + ((g2434) & (!g2533) & (g2480) & (!g2537) & (!g5054)) + ((g2434) & (!g2533) & (g2480) & (!g2537) & (g5054)) + ((g2434) & (g2533) & (!g2480) & (!g2537) & (g5054)) + ((g2434) & (g2533) & (!g2480) & (g2537) & (!g5054)) + ((g2434) & (g2533) & (g2480) & (g2537) & (!g5054)) + ((g2434) & (g2533) & (g2480) & (g2537) & (g5054)));
	assign g5082 = (((!g1914) & (!g1991) & (!g2247) & (!g5080) & (g5081)) + ((!g1914) & (!g1991) & (!g2247) & (g5080) & (g5081)) + ((!g1914) & (!g1991) & (g2247) & (!g5080) & (g5081)) + ((!g1914) & (!g1991) & (g2247) & (g5080) & (g5081)) + ((!g1914) & (g1991) & (!g2247) & (!g5080) & (g5081)) + ((!g1914) & (g1991) & (!g2247) & (g5080) & (g5081)) + ((!g1914) & (g1991) & (g2247) & (!g5080) & (g5081)) + ((!g1914) & (g1991) & (g2247) & (g5080) & (g5081)) + ((g1914) & (!g1991) & (!g2247) & (!g5080) & (!g5081)) + ((g1914) & (!g1991) & (!g2247) & (!g5080) & (g5081)) + ((g1914) & (!g1991) & (g2247) & (g5080) & (!g5081)) + ((g1914) & (!g1991) & (g2247) & (g5080) & (g5081)) + ((g1914) & (g1991) & (!g2247) & (g5080) & (!g5081)) + ((g1914) & (g1991) & (!g2247) & (g5080) & (g5081)) + ((g1914) & (g1991) & (g2247) & (!g5080) & (!g5081)) + ((g1914) & (g1991) & (g2247) & (!g5080) & (g5081)));
	assign g8327 = (((!g5560) & (g5631) & (!g5083)) + ((!g5560) & (g5631) & (g5083)) + ((g5560) & (!g5631) & (g5083)) + ((g5560) & (g5631) & (g5083)));
	assign g5084 = (((!g830) & (!g2848) & (!g5082) & (g5083)) + ((!g830) & (!g2848) & (g5082) & (g5083)) + ((!g830) & (g2848) & (!g5082) & (g5083)) + ((!g830) & (g2848) & (g5082) & (g5083)) + ((g830) & (!g2848) & (g5082) & (!g5083)) + ((g830) & (!g2848) & (g5082) & (g5083)) + ((g830) & (g2848) & (!g5082) & (!g5083)) + ((g830) & (g2848) & (!g5082) & (g5083)));
	assign g5085 = (((!g2450) & (!g2527) & (!g2456) & (g2535) & (!g5064)) + ((!g2450) & (!g2527) & (!g2456) & (g2535) & (g5064)) + ((!g2450) & (!g2527) & (g2456) & (!g2535) & (!g5064)) + ((!g2450) & (!g2527) & (g2456) & (g2535) & (g5064)) + ((!g2450) & (g2527) & (!g2456) & (!g2535) & (!g5064)) + ((!g2450) & (g2527) & (!g2456) & (!g2535) & (g5064)) + ((!g2450) & (g2527) & (g2456) & (!g2535) & (g5064)) + ((!g2450) & (g2527) & (g2456) & (g2535) & (!g5064)) + ((g2450) & (!g2527) & (!g2456) & (!g2535) & (!g5064)) + ((g2450) & (!g2527) & (!g2456) & (g2535) & (g5064)) + ((g2450) & (!g2527) & (g2456) & (!g2535) & (!g5064)) + ((g2450) & (!g2527) & (g2456) & (!g2535) & (g5064)) + ((g2450) & (g2527) & (!g2456) & (!g2535) & (g5064)) + ((g2450) & (g2527) & (!g2456) & (g2535) & (!g5064)) + ((g2450) & (g2527) & (g2456) & (g2535) & (!g5064)) + ((g2450) & (g2527) & (g2456) & (g2535) & (g5064)));
	assign g5086 = (((!g3797) & (!g3798)));
	assign g5087 = (((!g1954) & (!g2250) & (!g5086)) + ((!g1954) & (g2250) & (g5086)) + ((g1954) & (!g2250) & (g5086)) + ((g1954) & (g2250) & (!g5086)));
	assign g5088 = (((!g830) & (!g1914) & (!g2851) & (!g5085) & (!g5087) & (key[147])) + ((!g830) & (!g1914) & (!g2851) & (!g5085) & (g5087) & (key[147])) + ((!g830) & (!g1914) & (!g2851) & (g5085) & (!g5087) & (key[147])) + ((!g830) & (!g1914) & (!g2851) & (g5085) & (g5087) & (key[147])) + ((!g830) & (!g1914) & (g2851) & (!g5085) & (!g5087) & (key[147])) + ((!g830) & (!g1914) & (g2851) & (!g5085) & (g5087) & (key[147])) + ((!g830) & (!g1914) & (g2851) & (g5085) & (!g5087) & (key[147])) + ((!g830) & (!g1914) & (g2851) & (g5085) & (g5087) & (key[147])) + ((!g830) & (g1914) & (!g2851) & (!g5085) & (!g5087) & (key[147])) + ((!g830) & (g1914) & (!g2851) & (!g5085) & (g5087) & (key[147])) + ((!g830) & (g1914) & (!g2851) & (g5085) & (!g5087) & (key[147])) + ((!g830) & (g1914) & (!g2851) & (g5085) & (g5087) & (key[147])) + ((!g830) & (g1914) & (g2851) & (!g5085) & (!g5087) & (key[147])) + ((!g830) & (g1914) & (g2851) & (!g5085) & (g5087) & (key[147])) + ((!g830) & (g1914) & (g2851) & (g5085) & (!g5087) & (key[147])) + ((!g830) & (g1914) & (g2851) & (g5085) & (g5087) & (key[147])) + ((g830) & (!g1914) & (!g2851) & (!g5085) & (g5087) & (!key[147])) + ((g830) & (!g1914) & (!g2851) & (!g5085) & (g5087) & (key[147])) + ((g830) & (!g1914) & (!g2851) & (g5085) & (g5087) & (!key[147])) + ((g830) & (!g1914) & (!g2851) & (g5085) & (g5087) & (key[147])) + ((g830) & (!g1914) & (g2851) & (!g5085) & (!g5087) & (!key[147])) + ((g830) & (!g1914) & (g2851) & (!g5085) & (!g5087) & (key[147])) + ((g830) & (!g1914) & (g2851) & (g5085) & (!g5087) & (!key[147])) + ((g830) & (!g1914) & (g2851) & (g5085) & (!g5087) & (key[147])) + ((g830) & (g1914) & (!g2851) & (g5085) & (!g5087) & (!key[147])) + ((g830) & (g1914) & (!g2851) & (g5085) & (!g5087) & (key[147])) + ((g830) & (g1914) & (!g2851) & (g5085) & (g5087) & (!key[147])) + ((g830) & (g1914) & (!g2851) & (g5085) & (g5087) & (key[147])) + ((g830) & (g1914) & (g2851) & (!g5085) & (!g5087) & (!key[147])) + ((g830) & (g1914) & (g2851) & (!g5085) & (!g5087) & (key[147])) + ((g830) & (g1914) & (g2851) & (!g5085) & (g5087) & (!key[147])) + ((g830) & (g1914) & (g2851) & (!g5085) & (g5087) & (key[147])));
	assign g5089 = (((!g3432) & (!g3433)));
	assign g5090 = (((!g5089) & (!g2227) & (!g2250)) + ((!g5089) & (g2227) & (g2250)) + ((g5089) & (!g2227) & (g2250)) + ((g5089) & (g2227) & (!g2250)));
	assign g5091 = (((!g2004) & (!g2006) & (!g1199) & (g1236) & (!g5038)) + ((!g2004) & (!g2006) & (!g1199) & (g1236) & (g5038)) + ((!g2004) & (!g2006) & (g1199) & (!g1236) & (!g5038)) + ((!g2004) & (!g2006) & (g1199) & (g1236) & (g5038)) + ((!g2004) & (g2006) & (!g1199) & (!g1236) & (!g5038)) + ((!g2004) & (g2006) & (!g1199) & (!g1236) & (g5038)) + ((!g2004) & (g2006) & (g1199) & (!g1236) & (g5038)) + ((!g2004) & (g2006) & (g1199) & (g1236) & (!g5038)) + ((g2004) & (!g2006) & (!g1199) & (!g1236) & (!g5038)) + ((g2004) & (!g2006) & (!g1199) & (g1236) & (g5038)) + ((g2004) & (!g2006) & (g1199) & (!g1236) & (!g5038)) + ((g2004) & (!g2006) & (g1199) & (!g1236) & (g5038)) + ((g2004) & (g2006) & (!g1199) & (!g1236) & (g5038)) + ((g2004) & (g2006) & (!g1199) & (g1236) & (!g5038)) + ((g2004) & (g2006) & (g1199) & (g1236) & (!g5038)) + ((g2004) & (g2006) & (g1199) & (g1236) & (g5038)));
	assign g5092 = (((!g830) & (!g1914) & (!g2854) & (!g5090) & (!g5091) & (key[115])) + ((!g830) & (!g1914) & (!g2854) & (!g5090) & (g5091) & (key[115])) + ((!g830) & (!g1914) & (!g2854) & (g5090) & (!g5091) & (key[115])) + ((!g830) & (!g1914) & (!g2854) & (g5090) & (g5091) & (key[115])) + ((!g830) & (!g1914) & (g2854) & (!g5090) & (!g5091) & (key[115])) + ((!g830) & (!g1914) & (g2854) & (!g5090) & (g5091) & (key[115])) + ((!g830) & (!g1914) & (g2854) & (g5090) & (!g5091) & (key[115])) + ((!g830) & (!g1914) & (g2854) & (g5090) & (g5091) & (key[115])) + ((!g830) & (g1914) & (!g2854) & (!g5090) & (!g5091) & (key[115])) + ((!g830) & (g1914) & (!g2854) & (!g5090) & (g5091) & (key[115])) + ((!g830) & (g1914) & (!g2854) & (g5090) & (!g5091) & (key[115])) + ((!g830) & (g1914) & (!g2854) & (g5090) & (g5091) & (key[115])) + ((!g830) & (g1914) & (g2854) & (!g5090) & (!g5091) & (key[115])) + ((!g830) & (g1914) & (g2854) & (!g5090) & (g5091) & (key[115])) + ((!g830) & (g1914) & (g2854) & (g5090) & (!g5091) & (key[115])) + ((!g830) & (g1914) & (g2854) & (g5090) & (g5091) & (key[115])) + ((g830) & (!g1914) & (!g2854) & (!g5090) & (g5091) & (!key[115])) + ((g830) & (!g1914) & (!g2854) & (!g5090) & (g5091) & (key[115])) + ((g830) & (!g1914) & (!g2854) & (g5090) & (g5091) & (!key[115])) + ((g830) & (!g1914) & (!g2854) & (g5090) & (g5091) & (key[115])) + ((g830) & (!g1914) & (g2854) & (!g5090) & (!g5091) & (!key[115])) + ((g830) & (!g1914) & (g2854) & (!g5090) & (!g5091) & (key[115])) + ((g830) & (!g1914) & (g2854) & (g5090) & (!g5091) & (!key[115])) + ((g830) & (!g1914) & (g2854) & (g5090) & (!g5091) & (key[115])) + ((g830) & (g1914) & (!g2854) & (g5090) & (!g5091) & (!key[115])) + ((g830) & (g1914) & (!g2854) & (g5090) & (!g5091) & (key[115])) + ((g830) & (g1914) & (!g2854) & (g5090) & (g5091) & (!key[115])) + ((g830) & (g1914) & (!g2854) & (g5090) & (g5091) & (key[115])) + ((g830) & (g1914) & (g2854) & (!g5090) & (!g5091) & (!key[115])) + ((g830) & (g1914) & (g2854) & (!g5090) & (!g5091) & (key[115])) + ((g830) & (g1914) & (g2854) & (!g5090) & (g5091) & (!key[115])) + ((g830) & (g1914) & (g2854) & (!g5090) & (g5091) & (key[115])));
	assign g5093 = (((!g2468) & (!g2523) & (!g5042) & (!g2480) & (g2537)) + ((!g2468) & (!g2523) & (!g5042) & (g2480) & (!g2537)) + ((!g2468) & (!g2523) & (g5042) & (!g2480) & (g2537)) + ((!g2468) & (!g2523) & (g5042) & (g2480) & (g2537)) + ((!g2468) & (g2523) & (!g5042) & (!g2480) & (!g2537)) + ((!g2468) & (g2523) & (!g5042) & (g2480) & (g2537)) + ((!g2468) & (g2523) & (g5042) & (!g2480) & (!g2537)) + ((!g2468) & (g2523) & (g5042) & (g2480) & (!g2537)) + ((g2468) & (!g2523) & (!g5042) & (!g2480) & (!g2537)) + ((g2468) & (!g2523) & (!g5042) & (g2480) & (!g2537)) + ((g2468) & (!g2523) & (g5042) & (!g2480) & (g2537)) + ((g2468) & (!g2523) & (g5042) & (g2480) & (!g2537)) + ((g2468) & (g2523) & (!g5042) & (!g2480) & (g2537)) + ((g2468) & (g2523) & (!g5042) & (g2480) & (g2537)) + ((g2468) & (g2523) & (g5042) & (!g2480) & (!g2537)) + ((g2468) & (g2523) & (g5042) & (g2480) & (g2537)));
	assign g5094 = (((!g3574) & (!g3575)));
	assign g5095 = (((!g1953) & (!g2230) & (!g5094)) + ((!g1953) & (g2230) & (g5094)) + ((g1953) & (!g2230) & (g5094)) + ((g1953) & (g2230) & (!g5094)));
	assign g5096 = (((!g830) & (!g1914) & (!g2857) & (!g5093) & (!g5095) & (nonce[19])) + ((!g830) & (!g1914) & (!g2857) & (!g5093) & (g5095) & (nonce[19])) + ((!g830) & (!g1914) & (!g2857) & (g5093) & (!g5095) & (nonce[19])) + ((!g830) & (!g1914) & (!g2857) & (g5093) & (g5095) & (nonce[19])) + ((!g830) & (!g1914) & (g2857) & (!g5093) & (!g5095) & (nonce[19])) + ((!g830) & (!g1914) & (g2857) & (!g5093) & (g5095) & (nonce[19])) + ((!g830) & (!g1914) & (g2857) & (g5093) & (!g5095) & (nonce[19])) + ((!g830) & (!g1914) & (g2857) & (g5093) & (g5095) & (nonce[19])) + ((!g830) & (g1914) & (!g2857) & (!g5093) & (!g5095) & (nonce[19])) + ((!g830) & (g1914) & (!g2857) & (!g5093) & (g5095) & (nonce[19])) + ((!g830) & (g1914) & (!g2857) & (g5093) & (!g5095) & (nonce[19])) + ((!g830) & (g1914) & (!g2857) & (g5093) & (g5095) & (nonce[19])) + ((!g830) & (g1914) & (g2857) & (!g5093) & (!g5095) & (nonce[19])) + ((!g830) & (g1914) & (g2857) & (!g5093) & (g5095) & (nonce[19])) + ((!g830) & (g1914) & (g2857) & (g5093) & (!g5095) & (nonce[19])) + ((!g830) & (g1914) & (g2857) & (g5093) & (g5095) & (nonce[19])) + ((g830) & (!g1914) & (!g2857) & (!g5093) & (g5095) & (!nonce[19])) + ((g830) & (!g1914) & (!g2857) & (!g5093) & (g5095) & (nonce[19])) + ((g830) & (!g1914) & (!g2857) & (g5093) & (g5095) & (!nonce[19])) + ((g830) & (!g1914) & (!g2857) & (g5093) & (g5095) & (nonce[19])) + ((g830) & (!g1914) & (g2857) & (!g5093) & (!g5095) & (!nonce[19])) + ((g830) & (!g1914) & (g2857) & (!g5093) & (!g5095) & (nonce[19])) + ((g830) & (!g1914) & (g2857) & (g5093) & (!g5095) & (!nonce[19])) + ((g830) & (!g1914) & (g2857) & (g5093) & (!g5095) & (nonce[19])) + ((g830) & (g1914) & (!g2857) & (g5093) & (!g5095) & (!nonce[19])) + ((g830) & (g1914) & (!g2857) & (g5093) & (!g5095) & (nonce[19])) + ((g830) & (g1914) & (!g2857) & (g5093) & (g5095) & (!nonce[19])) + ((g830) & (g1914) & (!g2857) & (g5093) & (g5095) & (nonce[19])) + ((g830) & (g1914) & (g2857) & (!g5093) & (!g5095) & (!nonce[19])) + ((g830) & (g1914) & (g2857) & (!g5093) & (!g5095) & (nonce[19])) + ((g830) & (g1914) & (g2857) & (!g5093) & (g5095) & (!nonce[19])) + ((g830) & (g1914) & (g2857) & (!g5093) & (g5095) & (nonce[19])));
	assign g5097 = (((!g1886) & (!g2032) & (!g1910) & (g2038)) + ((!g1886) & (!g2032) & (g1910) & (g2038)) + ((!g1886) & (g2032) & (!g1910) & (!g2038)) + ((!g1886) & (g2032) & (g1910) & (!g2038)) + ((g1886) & (!g2032) & (!g1910) & (g2038)) + ((g1886) & (!g2032) & (g1910) & (!g2038)) + ((g1886) & (g2032) & (!g1910) & (!g2038)) + ((g1886) & (g2032) & (g1910) & (g2038)));
	assign g5098 = (((!g1898) & (!g2022) & (!g1904) & (g2043)) + ((!g1898) & (!g2022) & (g1904) & (g2043)) + ((!g1898) & (g2022) & (!g1904) & (!g2043)) + ((!g1898) & (g2022) & (g1904) & (!g2043)) + ((g1898) & (!g2022) & (!g1904) & (g2043)) + ((g1898) & (!g2022) & (g1904) & (!g2043)) + ((g1898) & (g2022) & (!g1904) & (!g2043)) + ((g1898) & (g2022) & (g1904) & (g2043)));
	assign g5099 = (((g830) & (!g1914) & (!g2860) & (!g5097) & (g5098)) + ((g830) & (!g1914) & (!g2860) & (g5097) & (g5098)) + ((g830) & (!g1914) & (g2860) & (!g5097) & (!g5098)) + ((g830) & (!g1914) & (g2860) & (g5097) & (!g5098)) + ((g830) & (g1914) & (!g2860) & (g5097) & (!g5098)) + ((g830) & (g1914) & (!g2860) & (g5097) & (g5098)) + ((g830) & (g1914) & (g2860) & (!g5097) & (!g5098)) + ((g830) & (g1914) & (g2860) & (!g5097) & (g5098)));
	assign g5100 = (((!g2362) & (!g2393) & (!g2364) & (g2405) & (!g5068)) + ((!g2362) & (!g2393) & (!g2364) & (g2405) & (g5068)) + ((!g2362) & (!g2393) & (g2364) & (!g2405) & (g5068)) + ((!g2362) & (!g2393) & (g2364) & (g2405) & (!g5068)) + ((!g2362) & (g2393) & (!g2364) & (!g2405) & (!g5068)) + ((!g2362) & (g2393) & (!g2364) & (!g2405) & (g5068)) + ((!g2362) & (g2393) & (g2364) & (!g2405) & (!g5068)) + ((!g2362) & (g2393) & (g2364) & (g2405) & (g5068)) + ((g2362) & (!g2393) & (!g2364) & (!g2405) & (g5068)) + ((g2362) & (!g2393) & (!g2364) & (g2405) & (!g5068)) + ((g2362) & (!g2393) & (g2364) & (!g2405) & (!g5068)) + ((g2362) & (!g2393) & (g2364) & (!g2405) & (g5068)) + ((g2362) & (g2393) & (!g2364) & (!g2405) & (!g5068)) + ((g2362) & (g2393) & (!g2364) & (g2405) & (g5068)) + ((g2362) & (g2393) & (g2364) & (g2405) & (!g5068)) + ((g2362) & (g2393) & (g2364) & (g2405) & (g5068)));
	assign g5101 = (((!g1961) & (!g1963) & (!g2373) & (g2419) & (!g5070)) + ((!g1961) & (!g1963) & (!g2373) & (g2419) & (g5070)) + ((!g1961) & (!g1963) & (g2373) & (!g2419) & (g5070)) + ((!g1961) & (!g1963) & (g2373) & (g2419) & (!g5070)) + ((!g1961) & (g1963) & (!g2373) & (!g2419) & (!g5070)) + ((!g1961) & (g1963) & (!g2373) & (!g2419) & (g5070)) + ((!g1961) & (g1963) & (g2373) & (!g2419) & (!g5070)) + ((!g1961) & (g1963) & (g2373) & (g2419) & (g5070)) + ((g1961) & (!g1963) & (!g2373) & (!g2419) & (g5070)) + ((g1961) & (!g1963) & (!g2373) & (g2419) & (!g5070)) + ((g1961) & (!g1963) & (g2373) & (!g2419) & (!g5070)) + ((g1961) & (!g1963) & (g2373) & (!g2419) & (g5070)) + ((g1961) & (g1963) & (!g2373) & (!g2419) & (!g5070)) + ((g1961) & (g1963) & (!g2373) & (g2419) & (g5070)) + ((g1961) & (g1963) & (g2373) & (g2419) & (!g5070)) + ((g1961) & (g1963) & (g2373) & (g2419) & (g5070)));
	assign g5102 = (((!g830) & (!g1914) & (!g2863) & (!g5100) & (!g5101) & (nonce[51])) + ((!g830) & (!g1914) & (!g2863) & (!g5100) & (g5101) & (nonce[51])) + ((!g830) & (!g1914) & (!g2863) & (g5100) & (!g5101) & (nonce[51])) + ((!g830) & (!g1914) & (!g2863) & (g5100) & (g5101) & (nonce[51])) + ((!g830) & (!g1914) & (g2863) & (!g5100) & (!g5101) & (nonce[51])) + ((!g830) & (!g1914) & (g2863) & (!g5100) & (g5101) & (nonce[51])) + ((!g830) & (!g1914) & (g2863) & (g5100) & (!g5101) & (nonce[51])) + ((!g830) & (!g1914) & (g2863) & (g5100) & (g5101) & (nonce[51])) + ((!g830) & (g1914) & (!g2863) & (!g5100) & (!g5101) & (nonce[51])) + ((!g830) & (g1914) & (!g2863) & (!g5100) & (g5101) & (nonce[51])) + ((!g830) & (g1914) & (!g2863) & (g5100) & (!g5101) & (nonce[51])) + ((!g830) & (g1914) & (!g2863) & (g5100) & (g5101) & (nonce[51])) + ((!g830) & (g1914) & (g2863) & (!g5100) & (!g5101) & (nonce[51])) + ((!g830) & (g1914) & (g2863) & (!g5100) & (g5101) & (nonce[51])) + ((!g830) & (g1914) & (g2863) & (g5100) & (!g5101) & (nonce[51])) + ((!g830) & (g1914) & (g2863) & (g5100) & (g5101) & (nonce[51])) + ((g830) & (!g1914) & (!g2863) & (!g5100) & (g5101) & (!nonce[51])) + ((g830) & (!g1914) & (!g2863) & (!g5100) & (g5101) & (nonce[51])) + ((g830) & (!g1914) & (!g2863) & (g5100) & (g5101) & (!nonce[51])) + ((g830) & (!g1914) & (!g2863) & (g5100) & (g5101) & (nonce[51])) + ((g830) & (!g1914) & (g2863) & (!g5100) & (!g5101) & (!nonce[51])) + ((g830) & (!g1914) & (g2863) & (!g5100) & (!g5101) & (nonce[51])) + ((g830) & (!g1914) & (g2863) & (g5100) & (!g5101) & (!nonce[51])) + ((g830) & (!g1914) & (g2863) & (g5100) & (!g5101) & (nonce[51])) + ((g830) & (g1914) & (!g2863) & (g5100) & (!g5101) & (!nonce[51])) + ((g830) & (g1914) & (!g2863) & (g5100) & (!g5101) & (nonce[51])) + ((g830) & (g1914) & (!g2863) & (g5100) & (g5101) & (!nonce[51])) + ((g830) & (g1914) & (!g2863) & (g5100) & (g5101) & (nonce[51])) + ((g830) & (g1914) & (g2863) & (!g5100) & (!g5101) & (!nonce[51])) + ((g830) & (g1914) & (g2863) & (!g5100) & (!g5101) & (nonce[51])) + ((g830) & (g1914) & (g2863) & (!g5100) & (g5101) & (!nonce[51])) + ((g830) & (g1914) & (g2863) & (!g5100) & (g5101) & (nonce[51])));
	assign g5103 = (((!g3590) & (!g3591)));
	assign g5104 = (((!g1992) & (!g5103) & (!g2242)) + ((!g1992) & (g5103) & (g2242)) + ((g1992) & (!g5103) & (g2242)) + ((g1992) & (g5103) & (!g2242)));
	assign g5105 = (((!g2450) & (!g2527) & (!g2474) & (g2529) & (!g5046)) + ((!g2450) & (!g2527) & (!g2474) & (g2529) & (g5046)) + ((!g2450) & (!g2527) & (g2474) & (!g2529) & (!g5046)) + ((!g2450) & (!g2527) & (g2474) & (g2529) & (g5046)) + ((!g2450) & (g2527) & (!g2474) & (!g2529) & (!g5046)) + ((!g2450) & (g2527) & (!g2474) & (!g2529) & (g5046)) + ((!g2450) & (g2527) & (g2474) & (!g2529) & (g5046)) + ((!g2450) & (g2527) & (g2474) & (g2529) & (!g5046)) + ((g2450) & (!g2527) & (!g2474) & (!g2529) & (!g5046)) + ((g2450) & (!g2527) & (!g2474) & (g2529) & (g5046)) + ((g2450) & (!g2527) & (g2474) & (!g2529) & (!g5046)) + ((g2450) & (!g2527) & (g2474) & (!g2529) & (g5046)) + ((g2450) & (g2527) & (!g2474) & (!g2529) & (g5046)) + ((g2450) & (g2527) & (!g2474) & (g2529) & (!g5046)) + ((g2450) & (g2527) & (g2474) & (g2529) & (!g5046)) + ((g2450) & (g2527) & (g2474) & (g2529) & (g5046)));
	assign g5106 = (((!g830) & (!g1914) & (!g2868) & (!g5104) & (!g5105) & (key[243])) + ((!g830) & (!g1914) & (!g2868) & (!g5104) & (g5105) & (key[243])) + ((!g830) & (!g1914) & (!g2868) & (g5104) & (!g5105) & (key[243])) + ((!g830) & (!g1914) & (!g2868) & (g5104) & (g5105) & (key[243])) + ((!g830) & (!g1914) & (g2868) & (!g5104) & (!g5105) & (key[243])) + ((!g830) & (!g1914) & (g2868) & (!g5104) & (g5105) & (key[243])) + ((!g830) & (!g1914) & (g2868) & (g5104) & (!g5105) & (key[243])) + ((!g830) & (!g1914) & (g2868) & (g5104) & (g5105) & (key[243])) + ((!g830) & (g1914) & (!g2868) & (!g5104) & (!g5105) & (key[243])) + ((!g830) & (g1914) & (!g2868) & (!g5104) & (g5105) & (key[243])) + ((!g830) & (g1914) & (!g2868) & (g5104) & (!g5105) & (key[243])) + ((!g830) & (g1914) & (!g2868) & (g5104) & (g5105) & (key[243])) + ((!g830) & (g1914) & (g2868) & (!g5104) & (!g5105) & (key[243])) + ((!g830) & (g1914) & (g2868) & (!g5104) & (g5105) & (key[243])) + ((!g830) & (g1914) & (g2868) & (g5104) & (!g5105) & (key[243])) + ((!g830) & (g1914) & (g2868) & (g5104) & (g5105) & (key[243])) + ((g830) & (!g1914) & (!g2868) & (!g5104) & (g5105) & (!key[243])) + ((g830) & (!g1914) & (!g2868) & (!g5104) & (g5105) & (key[243])) + ((g830) & (!g1914) & (!g2868) & (g5104) & (g5105) & (!key[243])) + ((g830) & (!g1914) & (!g2868) & (g5104) & (g5105) & (key[243])) + ((g830) & (!g1914) & (g2868) & (!g5104) & (!g5105) & (!key[243])) + ((g830) & (!g1914) & (g2868) & (!g5104) & (!g5105) & (key[243])) + ((g830) & (!g1914) & (g2868) & (g5104) & (!g5105) & (!key[243])) + ((g830) & (!g1914) & (g2868) & (g5104) & (!g5105) & (key[243])) + ((g830) & (g1914) & (!g2868) & (g5104) & (!g5105) & (!key[243])) + ((g830) & (g1914) & (!g2868) & (g5104) & (!g5105) & (key[243])) + ((g830) & (g1914) & (!g2868) & (g5104) & (g5105) & (!key[243])) + ((g830) & (g1914) & (!g2868) & (g5104) & (g5105) & (key[243])) + ((g830) & (g1914) & (g2868) & (!g5104) & (!g5105) & (!key[243])) + ((g830) & (g1914) & (g2868) & (!g5104) & (!g5105) & (key[243])) + ((g830) & (g1914) & (g2868) & (!g5104) & (g5105) & (!key[243])) + ((g830) & (g1914) & (g2868) & (!g5104) & (g5105) & (key[243])));
	assign g5107 = (((!g1999) & (!g2002) & (!g2373) & (g2419) & (!g5059)) + ((!g1999) & (!g2002) & (!g2373) & (g2419) & (g5059)) + ((!g1999) & (!g2002) & (g2373) & (!g2419) & (g5059)) + ((!g1999) & (!g2002) & (g2373) & (g2419) & (!g5059)) + ((!g1999) & (g2002) & (!g2373) & (!g2419) & (!g5059)) + ((!g1999) & (g2002) & (!g2373) & (!g2419) & (g5059)) + ((!g1999) & (g2002) & (g2373) & (!g2419) & (!g5059)) + ((!g1999) & (g2002) & (g2373) & (g2419) & (g5059)) + ((g1999) & (!g2002) & (!g2373) & (!g2419) & (g5059)) + ((g1999) & (!g2002) & (!g2373) & (g2419) & (!g5059)) + ((g1999) & (!g2002) & (g2373) & (!g2419) & (!g5059)) + ((g1999) & (!g2002) & (g2373) & (!g2419) & (g5059)) + ((g1999) & (g2002) & (!g2373) & (!g2419) & (!g5059)) + ((g1999) & (g2002) & (!g2373) & (g2419) & (g5059)) + ((g1999) & (g2002) & (g2373) & (g2419) & (!g5059)) + ((g1999) & (g2002) & (g2373) & (g2419) & (g5059)));
	assign g5108 = (((!g2356) & (!g2402) & (!g2364) & (g2405) & (!g5061)) + ((!g2356) & (!g2402) & (!g2364) & (g2405) & (g5061)) + ((!g2356) & (!g2402) & (g2364) & (!g2405) & (g5061)) + ((!g2356) & (!g2402) & (g2364) & (g2405) & (!g5061)) + ((!g2356) & (g2402) & (!g2364) & (!g2405) & (!g5061)) + ((!g2356) & (g2402) & (!g2364) & (!g2405) & (g5061)) + ((!g2356) & (g2402) & (g2364) & (!g2405) & (!g5061)) + ((!g2356) & (g2402) & (g2364) & (g2405) & (g5061)) + ((g2356) & (!g2402) & (!g2364) & (!g2405) & (g5061)) + ((g2356) & (!g2402) & (!g2364) & (g2405) & (!g5061)) + ((g2356) & (!g2402) & (g2364) & (!g2405) & (!g5061)) + ((g2356) & (!g2402) & (g2364) & (!g2405) & (g5061)) + ((g2356) & (g2402) & (!g2364) & (!g2405) & (!g5061)) + ((g2356) & (g2402) & (!g2364) & (g2405) & (g5061)) + ((g2356) & (g2402) & (g2364) & (g2405) & (!g5061)) + ((g2356) & (g2402) & (g2364) & (g2405) & (g5061)));
	assign g5109 = (((!g830) & (!g1914) & (!g2871) & (!g5107) & (!g5108) & (key[211])) + ((!g830) & (!g1914) & (!g2871) & (!g5107) & (g5108) & (key[211])) + ((!g830) & (!g1914) & (!g2871) & (g5107) & (!g5108) & (key[211])) + ((!g830) & (!g1914) & (!g2871) & (g5107) & (g5108) & (key[211])) + ((!g830) & (!g1914) & (g2871) & (!g5107) & (!g5108) & (key[211])) + ((!g830) & (!g1914) & (g2871) & (!g5107) & (g5108) & (key[211])) + ((!g830) & (!g1914) & (g2871) & (g5107) & (!g5108) & (key[211])) + ((!g830) & (!g1914) & (g2871) & (g5107) & (g5108) & (key[211])) + ((!g830) & (g1914) & (!g2871) & (!g5107) & (!g5108) & (key[211])) + ((!g830) & (g1914) & (!g2871) & (!g5107) & (g5108) & (key[211])) + ((!g830) & (g1914) & (!g2871) & (g5107) & (!g5108) & (key[211])) + ((!g830) & (g1914) & (!g2871) & (g5107) & (g5108) & (key[211])) + ((!g830) & (g1914) & (g2871) & (!g5107) & (!g5108) & (key[211])) + ((!g830) & (g1914) & (g2871) & (!g5107) & (g5108) & (key[211])) + ((!g830) & (g1914) & (g2871) & (g5107) & (!g5108) & (key[211])) + ((!g830) & (g1914) & (g2871) & (g5107) & (g5108) & (key[211])) + ((g830) & (!g1914) & (!g2871) & (!g5107) & (g5108) & (!key[211])) + ((g830) & (!g1914) & (!g2871) & (!g5107) & (g5108) & (key[211])) + ((g830) & (!g1914) & (!g2871) & (g5107) & (g5108) & (!key[211])) + ((g830) & (!g1914) & (!g2871) & (g5107) & (g5108) & (key[211])) + ((g830) & (!g1914) & (g2871) & (!g5107) & (!g5108) & (!key[211])) + ((g830) & (!g1914) & (g2871) & (!g5107) & (!g5108) & (key[211])) + ((g830) & (!g1914) & (g2871) & (g5107) & (!g5108) & (!key[211])) + ((g830) & (!g1914) & (g2871) & (g5107) & (!g5108) & (key[211])) + ((g830) & (g1914) & (!g2871) & (g5107) & (!g5108) & (!key[211])) + ((g830) & (g1914) & (!g2871) & (g5107) & (!g5108) & (key[211])) + ((g830) & (g1914) & (!g2871) & (g5107) & (g5108) & (!key[211])) + ((g830) & (g1914) & (!g2871) & (g5107) & (g5108) & (key[211])) + ((g830) & (g1914) & (g2871) & (!g5107) & (!g5108) & (!key[211])) + ((g830) & (g1914) & (g2871) & (!g5107) & (!g5108) & (key[211])) + ((g830) & (g1914) & (g2871) & (!g5107) & (g5108) & (!key[211])) + ((g830) & (g1914) & (g2871) & (!g5107) & (g5108) & (key[211])));
	assign g5110 = (((!g1896) & (!g2041) & (!g1904) & (g2043)) + ((!g1896) & (!g2041) & (g1904) & (g2043)) + ((!g1896) & (g2041) & (!g1904) & (!g2043)) + ((!g1896) & (g2041) & (g1904) & (!g2043)) + ((g1896) & (!g2041) & (!g1904) & (g2043)) + ((g1896) & (!g2041) & (g1904) & (!g2043)) + ((g1896) & (g2041) & (!g1904) & (!g2043)) + ((g1896) & (g2041) & (g1904) & (g2043)));
	assign g5111 = (((!g1908) & (!g2030) & (!g1910) & (g2038)) + ((!g1908) & (!g2030) & (g1910) & (g2038)) + ((!g1908) & (g2030) & (!g1910) & (!g2038)) + ((!g1908) & (g2030) & (g1910) & (!g2038)) + ((g1908) & (!g2030) & (!g1910) & (g2038)) + ((g1908) & (!g2030) & (g1910) & (!g2038)) + ((g1908) & (g2030) & (!g1910) & (!g2038)) + ((g1908) & (g2030) & (g1910) & (g2038)));
	assign g5112 = (((g830) & (!g1914) & (!g2874) & (!g5110) & (g5111)) + ((g830) & (!g1914) & (!g2874) & (g5110) & (g5111)) + ((g830) & (!g1914) & (g2874) & (!g5110) & (!g5111)) + ((g830) & (!g1914) & (g2874) & (g5110) & (!g5111)) + ((g830) & (g1914) & (!g2874) & (g5110) & (!g5111)) + ((g830) & (g1914) & (!g2874) & (g5110) & (g5111)) + ((g830) & (g1914) & (g2874) & (!g5110) & (!g5111)) + ((g830) & (g1914) & (g2874) & (!g5110) & (g5111)));
	assign g5113 = (((!g5089) & (!g2227) & (!g2250) & (!g2279) & (g2283)) + ((!g5089) & (!g2227) & (!g2250) & (g2279) & (!g2283)) + ((!g5089) & (!g2227) & (g2250) & (!g2279) & (!g2283)) + ((!g5089) & (!g2227) & (g2250) & (g2279) & (g2283)) + ((!g5089) & (g2227) & (!g2250) & (!g2279) & (!g2283)) + ((!g5089) & (g2227) & (!g2250) & (g2279) & (g2283)) + ((!g5089) & (g2227) & (g2250) & (!g2279) & (!g2283)) + ((!g5089) & (g2227) & (g2250) & (g2279) & (g2283)) + ((g5089) & (!g2227) & (!g2250) & (!g2279) & (g2283)) + ((g5089) & (!g2227) & (!g2250) & (g2279) & (!g2283)) + ((g5089) & (!g2227) & (g2250) & (!g2279) & (g2283)) + ((g5089) & (!g2227) & (g2250) & (g2279) & (!g2283)) + ((g5089) & (g2227) & (!g2250) & (!g2279) & (g2283)) + ((g5089) & (g2227) & (!g2250) & (g2279) & (!g2283)) + ((g5089) & (g2227) & (g2250) & (!g2279) & (!g2283)) + ((g5089) & (g2227) & (g2250) & (g2279) & (g2283)));
	assign g5114 = (((!g2012) & (!g1269) & (!g3452)) + ((!g2012) & (g1269) & (g3452)) + ((g2012) & (!g1269) & (g3452)) + ((g2012) & (g1269) & (!g3452)));
	assign g5115 = (((!g830) & (!g1914) & (!g2881) & (!g5113) & (!g5114) & (key[116])) + ((!g830) & (!g1914) & (!g2881) & (!g5113) & (g5114) & (key[116])) + ((!g830) & (!g1914) & (!g2881) & (g5113) & (!g5114) & (key[116])) + ((!g830) & (!g1914) & (!g2881) & (g5113) & (g5114) & (key[116])) + ((!g830) & (!g1914) & (g2881) & (!g5113) & (!g5114) & (key[116])) + ((!g830) & (!g1914) & (g2881) & (!g5113) & (g5114) & (key[116])) + ((!g830) & (!g1914) & (g2881) & (g5113) & (!g5114) & (key[116])) + ((!g830) & (!g1914) & (g2881) & (g5113) & (g5114) & (key[116])) + ((!g830) & (g1914) & (!g2881) & (!g5113) & (!g5114) & (key[116])) + ((!g830) & (g1914) & (!g2881) & (!g5113) & (g5114) & (key[116])) + ((!g830) & (g1914) & (!g2881) & (g5113) & (!g5114) & (key[116])) + ((!g830) & (g1914) & (!g2881) & (g5113) & (g5114) & (key[116])) + ((!g830) & (g1914) & (g2881) & (!g5113) & (!g5114) & (key[116])) + ((!g830) & (g1914) & (g2881) & (!g5113) & (g5114) & (key[116])) + ((!g830) & (g1914) & (g2881) & (g5113) & (!g5114) & (key[116])) + ((!g830) & (g1914) & (g2881) & (g5113) & (g5114) & (key[116])) + ((g830) & (!g1914) & (!g2881) & (!g5113) & (g5114) & (!key[116])) + ((g830) & (!g1914) & (!g2881) & (!g5113) & (g5114) & (key[116])) + ((g830) & (!g1914) & (!g2881) & (g5113) & (g5114) & (!key[116])) + ((g830) & (!g1914) & (!g2881) & (g5113) & (g5114) & (key[116])) + ((g830) & (!g1914) & (g2881) & (!g5113) & (!g5114) & (!key[116])) + ((g830) & (!g1914) & (g2881) & (!g5113) & (!g5114) & (key[116])) + ((g830) & (!g1914) & (g2881) & (g5113) & (!g5114) & (!key[116])) + ((g830) & (!g1914) & (g2881) & (g5113) & (!g5114) & (key[116])) + ((g830) & (g1914) & (!g2881) & (g5113) & (!g5114) & (!key[116])) + ((g830) & (g1914) & (!g2881) & (g5113) & (!g5114) & (key[116])) + ((g830) & (g1914) & (!g2881) & (g5113) & (g5114) & (!key[116])) + ((g830) & (g1914) & (!g2881) & (g5113) & (g5114) & (key[116])) + ((g830) & (g1914) & (g2881) & (!g5113) & (!g5114) & (!key[116])) + ((g830) & (g1914) & (g2881) & (!g5113) & (!g5114) & (key[116])) + ((g830) & (g1914) & (g2881) & (!g5113) & (g5114) & (!key[116])) + ((g830) & (g1914) & (g2881) & (!g5113) & (g5114) & (key[116])));
	assign g5116 = (((!g1884) & (g1977) & (!g1900) & (g2028)) + ((!g1884) & (g1977) & (g1900) & (g2028)) + ((g1884) & (!g1977) & (g1900) & (g2028)) + ((g1884) & (g1977) & (!g1900) & (g2028)) + ((g1884) & (g1977) & (g1900) & (!g2028)) + ((g1884) & (g1977) & (g1900) & (g2028)));
	assign g5117 = (((g1914) & (!g1979) & (!g5116) & (g2074)) + ((g1914) & (!g1979) & (g5116) & (!g2074)) + ((g1914) & (g1979) & (!g5116) & (!g2074)) + ((g1914) & (g1979) & (g5116) & (g2074)));
	assign g5118 = (((!g1890) & (g1939) & (!g1894) & (g2034)) + ((!g1890) & (g1939) & (g1894) & (g2034)) + ((g1890) & (!g1939) & (g1894) & (g2034)) + ((g1890) & (g1939) & (!g1894) & (g2034)) + ((g1890) & (g1939) & (g1894) & (!g2034)) + ((g1890) & (g1939) & (g1894) & (g2034)));
	assign g5119 = (((!g1914) & (!g1941) & (!g2065) & (g5118)) + ((!g1914) & (!g1941) & (g2065) & (!g5118)) + ((!g1914) & (g1941) & (!g2065) & (!g5118)) + ((!g1914) & (g1941) & (g2065) & (g5118)));
	assign g5120 = (((g830) & (!g2885) & (!g5117) & (g5119)) + ((g830) & (!g2885) & (g5117) & (!g5119)) + ((g830) & (!g2885) & (g5117) & (g5119)) + ((g830) & (g2885) & (!g5117) & (!g5119)));
	assign g5121 = (((!g2575) & (!g3562) & (!g2581)) + ((!g2575) & (g3562) & (g2581)) + ((g2575) & (!g3562) & (g2581)) + ((g2575) & (g3562) & (!g2581)));
	assign g5122 = (((!g1953) & (!g1955) & (!g2230) & (g2286) & (!g5094)) + ((!g1953) & (!g1955) & (!g2230) & (g2286) & (g5094)) + ((!g1953) & (!g1955) & (g2230) & (!g2286) & (!g5094)) + ((!g1953) & (!g1955) & (g2230) & (g2286) & (g5094)) + ((!g1953) & (g1955) & (!g2230) & (!g2286) & (!g5094)) + ((!g1953) & (g1955) & (!g2230) & (!g2286) & (g5094)) + ((!g1953) & (g1955) & (g2230) & (!g2286) & (g5094)) + ((!g1953) & (g1955) & (g2230) & (g2286) & (!g5094)) + ((g1953) & (!g1955) & (!g2230) & (!g2286) & (!g5094)) + ((g1953) & (!g1955) & (!g2230) & (g2286) & (g5094)) + ((g1953) & (!g1955) & (g2230) & (!g2286) & (!g5094)) + ((g1953) & (!g1955) & (g2230) & (!g2286) & (g5094)) + ((g1953) & (g1955) & (!g2230) & (!g2286) & (g5094)) + ((g1953) & (g1955) & (!g2230) & (g2286) & (!g5094)) + ((g1953) & (g1955) & (g2230) & (g2286) & (!g5094)) + ((g1953) & (g1955) & (g2230) & (g2286) & (g5094)));
	assign g5123 = (((!g830) & (!g1914) & (!g2887) & (!g5121) & (!g5122) & (nonce[20])) + ((!g830) & (!g1914) & (!g2887) & (!g5121) & (g5122) & (nonce[20])) + ((!g830) & (!g1914) & (!g2887) & (g5121) & (!g5122) & (nonce[20])) + ((!g830) & (!g1914) & (!g2887) & (g5121) & (g5122) & (nonce[20])) + ((!g830) & (!g1914) & (g2887) & (!g5121) & (!g5122) & (nonce[20])) + ((!g830) & (!g1914) & (g2887) & (!g5121) & (g5122) & (nonce[20])) + ((!g830) & (!g1914) & (g2887) & (g5121) & (!g5122) & (nonce[20])) + ((!g830) & (!g1914) & (g2887) & (g5121) & (g5122) & (nonce[20])) + ((!g830) & (g1914) & (!g2887) & (!g5121) & (!g5122) & (nonce[20])) + ((!g830) & (g1914) & (!g2887) & (!g5121) & (g5122) & (nonce[20])) + ((!g830) & (g1914) & (!g2887) & (g5121) & (!g5122) & (nonce[20])) + ((!g830) & (g1914) & (!g2887) & (g5121) & (g5122) & (nonce[20])) + ((!g830) & (g1914) & (g2887) & (!g5121) & (!g5122) & (nonce[20])) + ((!g830) & (g1914) & (g2887) & (!g5121) & (g5122) & (nonce[20])) + ((!g830) & (g1914) & (g2887) & (g5121) & (!g5122) & (nonce[20])) + ((!g830) & (g1914) & (g2887) & (g5121) & (g5122) & (nonce[20])) + ((g830) & (!g1914) & (!g2887) & (!g5121) & (g5122) & (!nonce[20])) + ((g830) & (!g1914) & (!g2887) & (!g5121) & (g5122) & (nonce[20])) + ((g830) & (!g1914) & (!g2887) & (g5121) & (g5122) & (!nonce[20])) + ((g830) & (!g1914) & (!g2887) & (g5121) & (g5122) & (nonce[20])) + ((g830) & (!g1914) & (g2887) & (!g5121) & (!g5122) & (!nonce[20])) + ((g830) & (!g1914) & (g2887) & (!g5121) & (!g5122) & (nonce[20])) + ((g830) & (!g1914) & (g2887) & (g5121) & (!g5122) & (!nonce[20])) + ((g830) & (!g1914) & (g2887) & (g5121) & (!g5122) & (nonce[20])) + ((g830) & (g1914) & (!g2887) & (g5121) & (!g5122) & (!nonce[20])) + ((g830) & (g1914) & (!g2887) & (g5121) & (!g5122) & (nonce[20])) + ((g830) & (g1914) & (!g2887) & (g5121) & (g5122) & (!nonce[20])) + ((g830) & (g1914) & (!g2887) & (g5121) & (g5122) & (nonce[20])) + ((g830) & (g1914) & (g2887) & (!g5121) & (!g5122) & (!nonce[20])) + ((g830) & (g1914) & (g2887) & (!g5121) & (!g5122) & (nonce[20])) + ((g830) & (g1914) & (g2887) & (!g5121) & (g5122) & (!nonce[20])) + ((g830) & (g1914) & (g2887) & (!g5121) & (g5122) & (nonce[20])));
	assign g5124 = (((!g1992) & (!g1994) & (!g5103) & (!g2242) & (g2288)) + ((!g1992) & (!g1994) & (!g5103) & (g2242) & (!g2288)) + ((!g1992) & (!g1994) & (g5103) & (!g2242) & (g2288)) + ((!g1992) & (!g1994) & (g5103) & (g2242) & (g2288)) + ((!g1992) & (g1994) & (!g5103) & (!g2242) & (!g2288)) + ((!g1992) & (g1994) & (!g5103) & (g2242) & (g2288)) + ((!g1992) & (g1994) & (g5103) & (!g2242) & (!g2288)) + ((!g1992) & (g1994) & (g5103) & (g2242) & (!g2288)) + ((g1992) & (!g1994) & (!g5103) & (!g2242) & (!g2288)) + ((g1992) & (!g1994) & (!g5103) & (g2242) & (!g2288)) + ((g1992) & (!g1994) & (g5103) & (!g2242) & (g2288)) + ((g1992) & (!g1994) & (g5103) & (g2242) & (!g2288)) + ((g1992) & (g1994) & (!g5103) & (!g2242) & (g2288)) + ((g1992) & (g1994) & (!g5103) & (g2242) & (g2288)) + ((g1992) & (g1994) & (g5103) & (!g2242) & (!g2288)) + ((g1992) & (g1994) & (g5103) & (g2242) & (g2288)));
	assign g5125 = (((!g2566) & (!g2578) & (!g3610)) + ((!g2566) & (g2578) & (g3610)) + ((g2566) & (!g2578) & (g3610)) + ((g2566) & (g2578) & (!g3610)));
	assign g5126 = (((!g830) & (!g1914) & (!g2889) & (!g5124) & (!g5125) & (key[244])) + ((!g830) & (!g1914) & (!g2889) & (!g5124) & (g5125) & (key[244])) + ((!g830) & (!g1914) & (!g2889) & (g5124) & (!g5125) & (key[244])) + ((!g830) & (!g1914) & (!g2889) & (g5124) & (g5125) & (key[244])) + ((!g830) & (!g1914) & (g2889) & (!g5124) & (!g5125) & (key[244])) + ((!g830) & (!g1914) & (g2889) & (!g5124) & (g5125) & (key[244])) + ((!g830) & (!g1914) & (g2889) & (g5124) & (!g5125) & (key[244])) + ((!g830) & (!g1914) & (g2889) & (g5124) & (g5125) & (key[244])) + ((!g830) & (g1914) & (!g2889) & (!g5124) & (!g5125) & (key[244])) + ((!g830) & (g1914) & (!g2889) & (!g5124) & (g5125) & (key[244])) + ((!g830) & (g1914) & (!g2889) & (g5124) & (!g5125) & (key[244])) + ((!g830) & (g1914) & (!g2889) & (g5124) & (g5125) & (key[244])) + ((!g830) & (g1914) & (g2889) & (!g5124) & (!g5125) & (key[244])) + ((!g830) & (g1914) & (g2889) & (!g5124) & (g5125) & (key[244])) + ((!g830) & (g1914) & (g2889) & (g5124) & (!g5125) & (key[244])) + ((!g830) & (g1914) & (g2889) & (g5124) & (g5125) & (key[244])) + ((g830) & (!g1914) & (!g2889) & (!g5124) & (g5125) & (!key[244])) + ((g830) & (!g1914) & (!g2889) & (!g5124) & (g5125) & (key[244])) + ((g830) & (!g1914) & (!g2889) & (g5124) & (g5125) & (!key[244])) + ((g830) & (!g1914) & (!g2889) & (g5124) & (g5125) & (key[244])) + ((g830) & (!g1914) & (g2889) & (!g5124) & (!g5125) & (!key[244])) + ((g830) & (!g1914) & (g2889) & (!g5124) & (!g5125) & (key[244])) + ((g830) & (!g1914) & (g2889) & (g5124) & (!g5125) & (!key[244])) + ((g830) & (!g1914) & (g2889) & (g5124) & (!g5125) & (key[244])) + ((g830) & (g1914) & (!g2889) & (g5124) & (!g5125) & (!key[244])) + ((g830) & (g1914) & (!g2889) & (g5124) & (!g5125) & (key[244])) + ((g830) & (g1914) & (!g2889) & (g5124) & (g5125) & (!key[244])) + ((g830) & (g1914) & (!g2889) & (g5124) & (g5125) & (key[244])) + ((g830) & (g1914) & (g2889) & (!g5124) & (!g5125) & (!key[244])) + ((g830) & (g1914) & (g2889) & (!g5124) & (!g5125) & (key[244])) + ((g830) & (g1914) & (g2889) & (!g5124) & (g5125) & (!key[244])) + ((g830) & (g1914) & (g2889) & (!g5124) & (g5125) & (key[244])));
	assign g5127 = (((!g1973) & (!g1269) & (!g3629)) + ((!g1973) & (g1269) & (g3629)) + ((g1973) & (!g1269) & (g3629)) + ((g1973) & (g1269) & (!g3629)));
	assign g5128 = (((!g2236) & (!g2273) & (!g2242) & (g2288) & (!g5074)) + ((!g2236) & (!g2273) & (!g2242) & (g2288) & (g5074)) + ((!g2236) & (!g2273) & (g2242) & (!g2288) & (!g5074)) + ((!g2236) & (!g2273) & (g2242) & (g2288) & (g5074)) + ((!g2236) & (g2273) & (!g2242) & (!g2288) & (!g5074)) + ((!g2236) & (g2273) & (!g2242) & (!g2288) & (g5074)) + ((!g2236) & (g2273) & (g2242) & (!g2288) & (g5074)) + ((!g2236) & (g2273) & (g2242) & (g2288) & (!g5074)) + ((g2236) & (!g2273) & (!g2242) & (!g2288) & (!g5074)) + ((g2236) & (!g2273) & (!g2242) & (g2288) & (g5074)) + ((g2236) & (!g2273) & (g2242) & (!g2288) & (!g5074)) + ((g2236) & (!g2273) & (g2242) & (!g2288) & (g5074)) + ((g2236) & (g2273) & (!g2242) & (!g2288) & (g5074)) + ((g2236) & (g2273) & (!g2242) & (g2288) & (!g5074)) + ((g2236) & (g2273) & (g2242) & (g2288) & (!g5074)) + ((g2236) & (g2273) & (g2242) & (g2288) & (g5074)));
	assign g5129 = (((!g830) & (!g1914) & (!g2891) & (!g5127) & (!g5128) & (key[20])) + ((!g830) & (!g1914) & (!g2891) & (!g5127) & (g5128) & (key[20])) + ((!g830) & (!g1914) & (!g2891) & (g5127) & (!g5128) & (key[20])) + ((!g830) & (!g1914) & (!g2891) & (g5127) & (g5128) & (key[20])) + ((!g830) & (!g1914) & (g2891) & (!g5127) & (!g5128) & (key[20])) + ((!g830) & (!g1914) & (g2891) & (!g5127) & (g5128) & (key[20])) + ((!g830) & (!g1914) & (g2891) & (g5127) & (!g5128) & (key[20])) + ((!g830) & (!g1914) & (g2891) & (g5127) & (g5128) & (key[20])) + ((!g830) & (g1914) & (!g2891) & (!g5127) & (!g5128) & (key[20])) + ((!g830) & (g1914) & (!g2891) & (!g5127) & (g5128) & (key[20])) + ((!g830) & (g1914) & (!g2891) & (g5127) & (!g5128) & (key[20])) + ((!g830) & (g1914) & (!g2891) & (g5127) & (g5128) & (key[20])) + ((!g830) & (g1914) & (g2891) & (!g5127) & (!g5128) & (key[20])) + ((!g830) & (g1914) & (g2891) & (!g5127) & (g5128) & (key[20])) + ((!g830) & (g1914) & (g2891) & (g5127) & (!g5128) & (key[20])) + ((!g830) & (g1914) & (g2891) & (g5127) & (g5128) & (key[20])) + ((g830) & (!g1914) & (!g2891) & (!g5127) & (g5128) & (!key[20])) + ((g830) & (!g1914) & (!g2891) & (!g5127) & (g5128) & (key[20])) + ((g830) & (!g1914) & (!g2891) & (g5127) & (g5128) & (!key[20])) + ((g830) & (!g1914) & (!g2891) & (g5127) & (g5128) & (key[20])) + ((g830) & (!g1914) & (g2891) & (!g5127) & (!g5128) & (!key[20])) + ((g830) & (!g1914) & (g2891) & (!g5127) & (!g5128) & (key[20])) + ((g830) & (!g1914) & (g2891) & (g5127) & (!g5128) & (!key[20])) + ((g830) & (!g1914) & (g2891) & (g5127) & (!g5128) & (key[20])) + ((g830) & (g1914) & (!g2891) & (g5127) & (!g5128) & (!key[20])) + ((g830) & (g1914) & (!g2891) & (g5127) & (!g5128) & (key[20])) + ((g830) & (g1914) & (!g2891) & (g5127) & (g5128) & (!key[20])) + ((g830) & (g1914) & (!g2891) & (g5127) & (g5128) & (key[20])) + ((g830) & (g1914) & (g2891) & (!g5127) & (!g5128) & (!key[20])) + ((g830) & (g1914) & (g2891) & (!g5127) & (!g5128) & (key[20])) + ((g830) & (g1914) & (g2891) & (!g5127) & (g5128) & (!key[20])) + ((g830) & (g1914) & (g2891) & (!g5127) & (g5128) & (key[20])));
	assign g5130 = (((!g1991) & (!g1993) & (!g2247) & (g2275) & (!g5080)) + ((!g1991) & (!g1993) & (!g2247) & (g2275) & (g5080)) + ((!g1991) & (!g1993) & (g2247) & (!g2275) & (!g5080)) + ((!g1991) & (!g1993) & (g2247) & (g2275) & (g5080)) + ((!g1991) & (g1993) & (!g2247) & (!g2275) & (!g5080)) + ((!g1991) & (g1993) & (!g2247) & (!g2275) & (g5080)) + ((!g1991) & (g1993) & (g2247) & (!g2275) & (g5080)) + ((!g1991) & (g1993) & (g2247) & (g2275) & (!g5080)) + ((g1991) & (!g1993) & (!g2247) & (!g2275) & (!g5080)) + ((g1991) & (!g1993) & (!g2247) & (g2275) & (g5080)) + ((g1991) & (!g1993) & (g2247) & (!g2275) & (!g5080)) + ((g1991) & (!g1993) & (g2247) & (!g2275) & (g5080)) + ((g1991) & (g1993) & (!g2247) & (!g2275) & (g5080)) + ((g1991) & (g1993) & (!g2247) & (g2275) & (!g5080)) + ((g1991) & (g1993) & (g2247) & (g2275) & (!g5080)) + ((g1991) & (g1993) & (g2247) & (g2275) & (g5080)));
	assign g5131 = (((!g1914) & (!g2559) & (!g2581) & (!g3677) & (!g5130)) + ((!g1914) & (!g2559) & (!g2581) & (!g3677) & (g5130)) + ((!g1914) & (!g2559) & (g2581) & (g3677) & (!g5130)) + ((!g1914) & (!g2559) & (g2581) & (g3677) & (g5130)) + ((!g1914) & (g2559) & (!g2581) & (g3677) & (!g5130)) + ((!g1914) & (g2559) & (!g2581) & (g3677) & (g5130)) + ((!g1914) & (g2559) & (g2581) & (!g3677) & (!g5130)) + ((!g1914) & (g2559) & (g2581) & (!g3677) & (g5130)) + ((g1914) & (!g2559) & (!g2581) & (!g3677) & (g5130)) + ((g1914) & (!g2559) & (!g2581) & (g3677) & (g5130)) + ((g1914) & (!g2559) & (g2581) & (!g3677) & (g5130)) + ((g1914) & (!g2559) & (g2581) & (g3677) & (g5130)) + ((g1914) & (g2559) & (!g2581) & (!g3677) & (g5130)) + ((g1914) & (g2559) & (!g2581) & (g3677) & (g5130)) + ((g1914) & (g2559) & (g2581) & (!g3677) & (g5130)) + ((g1914) & (g2559) & (g2581) & (g3677) & (g5130)));
	assign g8328 = (((!g5560) & (g5632) & (!g5132)) + ((!g5560) & (g5632) & (g5132)) + ((g5560) & (!g5632) & (g5132)) + ((g5560) & (g5632) & (g5132)));
	assign g5133 = (((!g830) & (!g2893) & (!g5131) & (g5132)) + ((!g830) & (!g2893) & (g5131) & (g5132)) + ((!g830) & (g2893) & (!g5131) & (g5132)) + ((!g830) & (g2893) & (g5131) & (g5132)) + ((g830) & (!g2893) & (g5131) & (!g5132)) + ((g830) & (!g2893) & (g5131) & (g5132)) + ((g830) & (g2893) & (!g5131) & (!g5132)) + ((g830) & (g2893) & (!g5131) & (g5132)));
	assign g5134 = (((!g1886) & (g2032) & (!g1910) & (g2038)) + ((!g1886) & (g2032) & (g1910) & (g2038)) + ((g1886) & (!g2032) & (g1910) & (g2038)) + ((g1886) & (g2032) & (!g1910) & (g2038)) + ((g1886) & (g2032) & (g1910) & (!g2038)) + ((g1886) & (g2032) & (g1910) & (g2038)));
	assign g5135 = (((g1914) & (!g2055) & (!g2088) & (g5134)) + ((g1914) & (!g2055) & (g2088) & (!g5134)) + ((g1914) & (g2055) & (!g2088) & (!g5134)) + ((g1914) & (g2055) & (g2088) & (g5134)));
	assign g5136 = (((!g1898) & (g2022) & (!g1904) & (g2043)) + ((!g1898) & (g2022) & (g1904) & (g2043)) + ((g1898) & (!g2022) & (g1904) & (g2043)) + ((g1898) & (g2022) & (!g1904) & (g2043)) + ((g1898) & (g2022) & (g1904) & (!g2043)) + ((g1898) & (g2022) & (g1904) & (g2043)));
	assign g5137 = (((!g1914) & (!g2071) & (!g2080) & (g5136)) + ((!g1914) & (!g2071) & (g2080) & (!g5136)) + ((!g1914) & (g2071) & (!g2080) & (!g5136)) + ((!g1914) & (g2071) & (g2080) & (g5136)));
	assign g5138 = (((g830) & (!g2895) & (!g5135) & (g5137)) + ((g830) & (!g2895) & (g5135) & (!g5137)) + ((g830) & (!g2895) & (g5135) & (g5137)) + ((g830) & (g2895) & (!g5135) & (!g5137)));
	assign g5139 = (((!g3716) & (!g3717)));
	assign g5140 = (((g1914) & (!g2004) & (!g2509) & (!g5139)) + ((g1914) & (!g2004) & (g2509) & (g5139)) + ((g1914) & (g2004) & (!g2509) & (g5139)) + ((g1914) & (g2004) & (g2509) & (!g5139)));
	assign g5141 = (((!g3733) & (!g3734)));
	assign g5142 = (((!g1914) & (!g2456) & (!g2480) & (!g5141)) + ((!g1914) & (!g2456) & (g2480) & (g5141)) + ((!g1914) & (g2456) & (!g2480) & (g5141)) + ((!g1914) & (g2456) & (g2480) & (!g5141)));
	assign g5143 = (((!g830) & (!g2897) & (!g5140) & (!g5142) & (key[212])) + ((!g830) & (!g2897) & (!g5140) & (g5142) & (key[212])) + ((!g830) & (!g2897) & (g5140) & (!g5142) & (key[212])) + ((!g830) & (!g2897) & (g5140) & (g5142) & (key[212])) + ((!g830) & (g2897) & (!g5140) & (!g5142) & (key[212])) + ((!g830) & (g2897) & (!g5140) & (g5142) & (key[212])) + ((!g830) & (g2897) & (g5140) & (!g5142) & (key[212])) + ((!g830) & (g2897) & (g5140) & (g5142) & (key[212])) + ((g830) & (!g2897) & (!g5140) & (g5142) & (!key[212])) + ((g830) & (!g2897) & (!g5140) & (g5142) & (key[212])) + ((g830) & (!g2897) & (g5140) & (!g5142) & (!key[212])) + ((g830) & (!g2897) & (g5140) & (!g5142) & (key[212])) + ((g830) & (!g2897) & (g5140) & (g5142) & (!key[212])) + ((g830) & (!g2897) & (g5140) & (g5142) & (key[212])) + ((g830) & (g2897) & (!g5140) & (!g5142) & (!key[212])) + ((g830) & (g2897) & (!g5140) & (!g5142) & (key[212])));
	assign g5144 = (((!g2566) & (!g2569) & (!g3786)) + ((!g2566) & (g2569) & (g3786)) + ((g2566) & (!g2569) & (g3786)) + ((g2566) & (g2569) & (!g3786)));
	assign g5145 = (((!g1954) & (!g1956) & (!g2250) & (g2283) & (!g5086)) + ((!g1954) & (!g1956) & (!g2250) & (g2283) & (g5086)) + ((!g1954) & (!g1956) & (g2250) & (!g2283) & (!g5086)) + ((!g1954) & (!g1956) & (g2250) & (g2283) & (g5086)) + ((!g1954) & (g1956) & (!g2250) & (!g2283) & (!g5086)) + ((!g1954) & (g1956) & (!g2250) & (!g2283) & (g5086)) + ((!g1954) & (g1956) & (g2250) & (!g2283) & (g5086)) + ((!g1954) & (g1956) & (g2250) & (g2283) & (!g5086)) + ((g1954) & (!g1956) & (!g2250) & (!g2283) & (!g5086)) + ((g1954) & (!g1956) & (!g2250) & (g2283) & (g5086)) + ((g1954) & (!g1956) & (g2250) & (!g2283) & (!g5086)) + ((g1954) & (!g1956) & (g2250) & (!g2283) & (g5086)) + ((g1954) & (g1956) & (!g2250) & (!g2283) & (g5086)) + ((g1954) & (g1956) & (!g2250) & (g2283) & (!g5086)) + ((g1954) & (g1956) & (g2250) & (g2283) & (!g5086)) + ((g1954) & (g1956) & (g2250) & (g2283) & (g5086)));
	assign g5146 = (((!g830) & (!g1914) & (!g2900) & (!g5144) & (!g5145) & (key[148])) + ((!g830) & (!g1914) & (!g2900) & (!g5144) & (g5145) & (key[148])) + ((!g830) & (!g1914) & (!g2900) & (g5144) & (!g5145) & (key[148])) + ((!g830) & (!g1914) & (!g2900) & (g5144) & (g5145) & (key[148])) + ((!g830) & (!g1914) & (g2900) & (!g5144) & (!g5145) & (key[148])) + ((!g830) & (!g1914) & (g2900) & (!g5144) & (g5145) & (key[148])) + ((!g830) & (!g1914) & (g2900) & (g5144) & (!g5145) & (key[148])) + ((!g830) & (!g1914) & (g2900) & (g5144) & (g5145) & (key[148])) + ((!g830) & (g1914) & (!g2900) & (!g5144) & (!g5145) & (key[148])) + ((!g830) & (g1914) & (!g2900) & (!g5144) & (g5145) & (key[148])) + ((!g830) & (g1914) & (!g2900) & (g5144) & (!g5145) & (key[148])) + ((!g830) & (g1914) & (!g2900) & (g5144) & (g5145) & (key[148])) + ((!g830) & (g1914) & (g2900) & (!g5144) & (!g5145) & (key[148])) + ((!g830) & (g1914) & (g2900) & (!g5144) & (g5145) & (key[148])) + ((!g830) & (g1914) & (g2900) & (g5144) & (!g5145) & (key[148])) + ((!g830) & (g1914) & (g2900) & (g5144) & (g5145) & (key[148])) + ((g830) & (!g1914) & (!g2900) & (!g5144) & (g5145) & (!key[148])) + ((g830) & (!g1914) & (!g2900) & (!g5144) & (g5145) & (key[148])) + ((g830) & (!g1914) & (!g2900) & (g5144) & (g5145) & (!key[148])) + ((g830) & (!g1914) & (!g2900) & (g5144) & (g5145) & (key[148])) + ((g830) & (!g1914) & (g2900) & (!g5144) & (!g5145) & (!key[148])) + ((g830) & (!g1914) & (g2900) & (!g5144) & (!g5145) & (key[148])) + ((g830) & (!g1914) & (g2900) & (g5144) & (!g5145) & (!key[148])) + ((g830) & (!g1914) & (g2900) & (g5144) & (!g5145) & (key[148])) + ((g830) & (g1914) & (!g2900) & (g5144) & (!g5145) & (!key[148])) + ((g830) & (g1914) & (!g2900) & (g5144) & (!g5145) & (key[148])) + ((g830) & (g1914) & (!g2900) & (g5144) & (g5145) & (!key[148])) + ((g830) & (g1914) & (!g2900) & (g5144) & (g5145) & (key[148])) + ((g830) & (g1914) & (g2900) & (!g5144) & (!g5145) & (!key[148])) + ((g830) & (g1914) & (g2900) & (!g5144) & (!g5145) & (key[148])) + ((g830) & (g1914) & (g2900) & (!g5144) & (g5145) & (!key[148])) + ((g830) & (g1914) & (g2900) & (!g5144) & (g5145) & (key[148])));
	assign g5147 = (((!g3817) & (!g3818)));
	assign g5148 = (((g1914) & (!g2474) & (!g2480) & (!g5147)) + ((g1914) & (!g2474) & (g2480) & (g5147)) + ((g1914) & (g2474) & (!g2480) & (g5147)) + ((g1914) & (g2474) & (g2480) & (!g5147)));
	assign g5149 = (((!g3834) & (!g3835)));
	assign g5150 = (((!g1914) & (!g1968) & (!g2509) & (!g5149)) + ((!g1914) & (!g1968) & (g2509) & (g5149)) + ((!g1914) & (g1968) & (!g2509) & (g5149)) + ((!g1914) & (g1968) & (g2509) & (!g5149)));
	assign g5151 = (((!g830) & (!g2902) & (!g5148) & (!g5150) & (nonce[52])) + ((!g830) & (!g2902) & (!g5148) & (g5150) & (nonce[52])) + ((!g830) & (!g2902) & (g5148) & (!g5150) & (nonce[52])) + ((!g830) & (!g2902) & (g5148) & (g5150) & (nonce[52])) + ((!g830) & (g2902) & (!g5148) & (!g5150) & (nonce[52])) + ((!g830) & (g2902) & (!g5148) & (g5150) & (nonce[52])) + ((!g830) & (g2902) & (g5148) & (!g5150) & (nonce[52])) + ((!g830) & (g2902) & (g5148) & (g5150) & (nonce[52])) + ((g830) & (!g2902) & (!g5148) & (g5150) & (!nonce[52])) + ((g830) & (!g2902) & (!g5148) & (g5150) & (nonce[52])) + ((g830) & (!g2902) & (g5148) & (!g5150) & (!nonce[52])) + ((g830) & (!g2902) & (g5148) & (!g5150) & (nonce[52])) + ((g830) & (!g2902) & (g5148) & (g5150) & (!nonce[52])) + ((g830) & (!g2902) & (g5148) & (g5150) & (nonce[52])) + ((g830) & (g2902) & (!g5148) & (!g5150) & (!nonce[52])) + ((g830) & (g2902) & (!g5148) & (!g5150) & (nonce[52])));
	assign g5152 = (((!g1896) & (g2041) & (!g1904) & (g2043)) + ((!g1896) & (g2041) & (g1904) & (g2043)) + ((g1896) & (!g2041) & (g1904) & (g2043)) + ((g1896) & (g2041) & (!g1904) & (g2043)) + ((g1896) & (g2041) & (g1904) & (!g2043)) + ((g1896) & (g2041) & (g1904) & (g2043)));
	assign g5153 = (((g1914) & (!g2068) & (!g2080) & (g5152)) + ((g1914) & (!g2068) & (g2080) & (!g5152)) + ((g1914) & (g2068) & (!g2080) & (!g5152)) + ((g1914) & (g2068) & (g2080) & (g5152)));
	assign g5154 = (((!g1908) & (g2030) & (!g1910) & (g2038)) + ((!g1908) & (g2030) & (g1910) & (g2038)) + ((g1908) & (!g2030) & (g1910) & (g2038)) + ((g1908) & (g2030) & (!g1910) & (g2038)) + ((g1908) & (g2030) & (g1910) & (!g2038)) + ((g1908) & (g2030) & (g1910) & (g2038)));
	assign g5155 = (((!g1914) & (!g2085) & (!g2088) & (g5154)) + ((!g1914) & (!g2085) & (g2088) & (!g5154)) + ((!g1914) & (g2085) & (!g2088) & (!g5154)) + ((!g1914) & (g2085) & (g2088) & (g5154)));
	assign g5156 = (((g830) & (!g2904) & (!g5153) & (g5155)) + ((g830) & (!g2904) & (g5153) & (!g5155)) + ((g830) & (!g2904) & (g5153) & (g5155)) + ((g830) & (g2904) & (!g5153) & (!g5155)));
	assign g5157 = (((!g1973) & (g1269) & (!g3629)) + ((g1973) & (!g1269) & (!g3629)) + ((g1973) & (g1269) & (!g3629)) + ((g1973) & (g1269) & (g3629)));
	assign g5158 = (((!g2323) & (!g2329) & (!g3642)) + ((!g2323) & (g2329) & (g3642)) + ((g2323) & (!g2329) & (g3642)) + ((g2323) & (g2329) & (!g3642)));
	assign g5159 = (((!g1914) & (!g1976) & (!g1303) & (!g5157) & (g5158)) + ((!g1914) & (!g1976) & (!g1303) & (g5157) & (g5158)) + ((!g1914) & (!g1976) & (g1303) & (!g5157) & (g5158)) + ((!g1914) & (!g1976) & (g1303) & (g5157) & (g5158)) + ((!g1914) & (g1976) & (!g1303) & (!g5157) & (g5158)) + ((!g1914) & (g1976) & (!g1303) & (g5157) & (g5158)) + ((!g1914) & (g1976) & (g1303) & (!g5157) & (g5158)) + ((!g1914) & (g1976) & (g1303) & (g5157) & (g5158)) + ((g1914) & (!g1976) & (!g1303) & (g5157) & (!g5158)) + ((g1914) & (!g1976) & (!g1303) & (g5157) & (g5158)) + ((g1914) & (!g1976) & (g1303) & (!g5157) & (!g5158)) + ((g1914) & (!g1976) & (g1303) & (!g5157) & (g5158)) + ((g1914) & (g1976) & (!g1303) & (!g5157) & (!g5158)) + ((g1914) & (g1976) & (!g1303) & (!g5157) & (g5158)) + ((g1914) & (g1976) & (g1303) & (g5157) & (!g5158)) + ((g1914) & (g1976) & (g1303) & (g5157) & (g5158)));
	assign g5160 = (((!g830) & (!g2916) & (!g5159) & (key[21])) + ((!g830) & (!g2916) & (g5159) & (key[21])) + ((!g830) & (g2916) & (!g5159) & (key[21])) + ((!g830) & (g2916) & (g5159) & (key[21])) + ((g830) & (!g2916) & (g5159) & (!key[21])) + ((g830) & (!g2916) & (g5159) & (key[21])) + ((g830) & (g2916) & (!g5159) & (!key[21])) + ((g830) & (g2916) & (!g5159) & (key[21])));
	assign g5161 = (((!g1944) & (!g2116) & (g3544)) + ((!g1944) & (g2116) & (!g3544)) + ((g1944) & (!g2116) & (!g3544)) + ((g1944) & (g2116) & (g3544)));
	assign g5162 = (((!g2559) & (g2581) & (!g3677)) + ((g2559) & (!g2581) & (!g3677)) + ((g2559) & (g2581) & (!g3677)) + ((g2559) & (g2581) & (g3677)));
	assign g5163 = (((!g1996) & (!g2334) & (!g3658)) + ((!g1996) & (g2334) & (g3658)) + ((g1996) & (!g2334) & (g3658)) + ((g1996) & (g2334) & (!g3658)));
	assign g5164 = (((!g1914) & (!g2623) & (!g2629) & (g5162) & (!g5163)) + ((!g1914) & (!g2623) & (!g2629) & (g5162) & (g5163)) + ((!g1914) & (!g2623) & (g2629) & (!g5162) & (!g5163)) + ((!g1914) & (!g2623) & (g2629) & (!g5162) & (g5163)) + ((!g1914) & (g2623) & (!g2629) & (!g5162) & (!g5163)) + ((!g1914) & (g2623) & (!g2629) & (!g5162) & (g5163)) + ((!g1914) & (g2623) & (g2629) & (g5162) & (!g5163)) + ((!g1914) & (g2623) & (g2629) & (g5162) & (g5163)) + ((g1914) & (!g2623) & (!g2629) & (!g5162) & (g5163)) + ((g1914) & (!g2623) & (!g2629) & (g5162) & (g5163)) + ((g1914) & (!g2623) & (g2629) & (!g5162) & (g5163)) + ((g1914) & (!g2623) & (g2629) & (g5162) & (g5163)) + ((g1914) & (g2623) & (!g2629) & (!g5162) & (g5163)) + ((g1914) & (g2623) & (!g2629) & (g5162) & (g5163)) + ((g1914) & (g2623) & (g2629) & (!g5162) & (g5163)) + ((g1914) & (g2623) & (g2629) & (g5162) & (g5163)));
	assign g8329 = (((!g5560) & (g5634) & (!g5165)) + ((!g5560) & (g5634) & (g5165)) + ((g5560) & (!g5634) & (g5165)) + ((g5560) & (g5634) & (g5165)));
	assign g5166 = (((!g830) & (!g2938) & (!g5164) & (g5165)) + ((!g830) & (!g2938) & (g5164) & (g5165)) + ((!g830) & (g2938) & (!g5164) & (g5165)) + ((!g830) & (g2938) & (g5164) & (g5165)) + ((g830) & (!g2938) & (g5164) & (!g5165)) + ((g830) & (!g2938) & (g5164) & (g5165)) + ((g830) & (g2938) & (!g5164) & (!g5165)) + ((g830) & (g2938) & (!g5164) & (g5165)));
	assign g5167 = (((!g2566) & (g2569) & (!g3786)) + ((g2566) & (!g2569) & (!g3786)) + ((g2566) & (g2569) & (!g3786)) + ((g2566) & (g2569) & (g3786)));
	assign g5168 = (((!g1959) & (!g2337) & (!g3799)) + ((!g1959) & (g2337) & (g3799)) + ((g1959) & (!g2337) & (g3799)) + ((g1959) & (g2337) & (!g3799)));
	assign g5169 = (((!g1914) & (!g2614) & (!g2626) & (!g5167) & (g5168)) + ((!g1914) & (!g2614) & (!g2626) & (g5167) & (g5168)) + ((!g1914) & (!g2614) & (g2626) & (!g5167) & (g5168)) + ((!g1914) & (!g2614) & (g2626) & (g5167) & (g5168)) + ((!g1914) & (g2614) & (!g2626) & (!g5167) & (g5168)) + ((!g1914) & (g2614) & (!g2626) & (g5167) & (g5168)) + ((!g1914) & (g2614) & (g2626) & (!g5167) & (g5168)) + ((!g1914) & (g2614) & (g2626) & (g5167) & (g5168)) + ((g1914) & (!g2614) & (!g2626) & (g5167) & (!g5168)) + ((g1914) & (!g2614) & (!g2626) & (g5167) & (g5168)) + ((g1914) & (!g2614) & (g2626) & (!g5167) & (!g5168)) + ((g1914) & (!g2614) & (g2626) & (!g5167) & (g5168)) + ((g1914) & (g2614) & (!g2626) & (!g5167) & (!g5168)) + ((g1914) & (g2614) & (!g2626) & (!g5167) & (g5168)) + ((g1914) & (g2614) & (g2626) & (g5167) & (!g5168)) + ((g1914) & (g2614) & (g2626) & (g5167) & (g5168)));
	assign g5170 = (((!g830) & (!g2944) & (!g5169) & (key[149])) + ((!g830) & (!g2944) & (g5169) & (key[149])) + ((!g830) & (g2944) & (!g5169) & (key[149])) + ((!g830) & (g2944) & (g5169) & (key[149])) + ((g830) & (!g2944) & (g5169) & (!key[149])) + ((g830) & (!g2944) & (g5169) & (key[149])) + ((g830) & (g2944) & (!g5169) & (!key[149])) + ((g830) & (g2944) & (!g5169) & (key[149])));
	assign g5171 = (((!g2012) & (g1269) & (!g3452)) + ((g2012) & (!g1269) & (!g3452)) + ((g2012) & (g1269) & (!g3452)) + ((g2012) & (g1269) & (g3452)));
	assign g5172 = (((!g3434) & (!g2314) & (!g2337)) + ((!g3434) & (g2314) & (g2337)) + ((g3434) & (!g2314) & (g2337)) + ((g3434) & (g2314) & (!g2337)));
	assign g5173 = (((!g1914) & (!g2014) & (!g1303) & (g5171) & (!g5172)) + ((!g1914) & (!g2014) & (!g1303) & (g5171) & (g5172)) + ((!g1914) & (!g2014) & (g1303) & (!g5171) & (!g5172)) + ((!g1914) & (!g2014) & (g1303) & (!g5171) & (g5172)) + ((!g1914) & (g2014) & (!g1303) & (!g5171) & (!g5172)) + ((!g1914) & (g2014) & (!g1303) & (!g5171) & (g5172)) + ((!g1914) & (g2014) & (g1303) & (g5171) & (!g5172)) + ((!g1914) & (g2014) & (g1303) & (g5171) & (g5172)) + ((g1914) & (!g2014) & (!g1303) & (!g5171) & (g5172)) + ((g1914) & (!g2014) & (!g1303) & (g5171) & (g5172)) + ((g1914) & (!g2014) & (g1303) & (!g5171) & (g5172)) + ((g1914) & (!g2014) & (g1303) & (g5171) & (g5172)) + ((g1914) & (g2014) & (!g1303) & (!g5171) & (g5172)) + ((g1914) & (g2014) & (!g1303) & (g5171) & (g5172)) + ((g1914) & (g2014) & (g1303) & (!g5171) & (g5172)) + ((g1914) & (g2014) & (g1303) & (g5171) & (g5172)));
	assign g5174 = (((!g830) & (!g2950) & (!g5173) & (key[117])) + ((!g830) & (!g2950) & (g5173) & (key[117])) + ((!g830) & (g2950) & (!g5173) & (key[117])) + ((!g830) & (g2950) & (g5173) & (key[117])) + ((g830) & (!g2950) & (g5173) & (!key[117])) + ((g830) & (!g2950) & (g5173) & (key[117])) + ((g830) & (g2950) & (!g5173) & (!key[117])) + ((g830) & (g2950) & (!g5173) & (key[117])));
	assign g5175 = (((!g2575) & (!g3562) & (g2581)) + ((g2575) & (!g3562) & (!g2581)) + ((g2575) & (!g3562) & (g2581)) + ((g2575) & (g3562) & (g2581)));
	assign g5176 = (((!g1958) & (!g2317) & (!g3576)) + ((!g1958) & (g2317) & (g3576)) + ((g1958) & (!g2317) & (g3576)) + ((g1958) & (g2317) & (!g3576)));
	assign g5177 = (((!g1914) & (!g2607) & (!g5175) & (!g2629) & (g5176)) + ((!g1914) & (!g2607) & (!g5175) & (g2629) & (g5176)) + ((!g1914) & (!g2607) & (g5175) & (!g2629) & (g5176)) + ((!g1914) & (!g2607) & (g5175) & (g2629) & (g5176)) + ((!g1914) & (g2607) & (!g5175) & (!g2629) & (g5176)) + ((!g1914) & (g2607) & (!g5175) & (g2629) & (g5176)) + ((!g1914) & (g2607) & (g5175) & (!g2629) & (g5176)) + ((!g1914) & (g2607) & (g5175) & (g2629) & (g5176)) + ((g1914) & (!g2607) & (!g5175) & (g2629) & (!g5176)) + ((g1914) & (!g2607) & (!g5175) & (g2629) & (g5176)) + ((g1914) & (!g2607) & (g5175) & (!g2629) & (!g5176)) + ((g1914) & (!g2607) & (g5175) & (!g2629) & (g5176)) + ((g1914) & (g2607) & (!g5175) & (!g2629) & (!g5176)) + ((g1914) & (g2607) & (!g5175) & (!g2629) & (g5176)) + ((g1914) & (g2607) & (g5175) & (g2629) & (!g5176)) + ((g1914) & (g2607) & (g5175) & (g2629) & (g5176)));
	assign g5178 = (((!g830) & (!g2956) & (!g5177) & (nonce[21])) + ((!g830) & (!g2956) & (g5177) & (nonce[21])) + ((!g830) & (g2956) & (!g5177) & (nonce[21])) + ((!g830) & (g2956) & (g5177) & (nonce[21])) + ((g830) & (!g2956) & (g5177) & (!nonce[21])) + ((g830) & (!g2956) & (g5177) & (nonce[21])) + ((g830) & (g2956) & (!g5177) & (!nonce[21])) + ((g830) & (g2956) & (!g5177) & (nonce[21])));
	assign g5179 = (((!g2104) & (!g2125) & (g3699)) + ((!g2104) & (g2125) & (!g3699)) + ((g2104) & (!g2125) & (!g3699)) + ((g2104) & (g2125) & (g3699)));
	assign g5180 = (((!g2474) & (!g2529) & (!g2480) & (g2537) & (!g5147)) + ((!g2474) & (!g2529) & (!g2480) & (g2537) & (g5147)) + ((!g2474) & (!g2529) & (g2480) & (!g2537) & (!g5147)) + ((!g2474) & (!g2529) & (g2480) & (g2537) & (g5147)) + ((!g2474) & (g2529) & (!g2480) & (!g2537) & (!g5147)) + ((!g2474) & (g2529) & (!g2480) & (!g2537) & (g5147)) + ((!g2474) & (g2529) & (g2480) & (!g2537) & (g5147)) + ((!g2474) & (g2529) & (g2480) & (g2537) & (!g5147)) + ((g2474) & (!g2529) & (!g2480) & (!g2537) & (!g5147)) + ((g2474) & (!g2529) & (!g2480) & (g2537) & (g5147)) + ((g2474) & (!g2529) & (g2480) & (!g2537) & (!g5147)) + ((g2474) & (!g2529) & (g2480) & (!g2537) & (g5147)) + ((g2474) & (g2529) & (!g2480) & (!g2537) & (g5147)) + ((g2474) & (g2529) & (!g2480) & (g2537) & (!g5147)) + ((g2474) & (g2529) & (g2480) & (g2537) & (!g5147)) + ((g2474) & (g2529) & (g2480) & (g2537) & (g5147)));
	assign g5181 = (((!g1968) & (!g1970) & (!g2509) & (g2546) & (!g5149)) + ((!g1968) & (!g1970) & (!g2509) & (g2546) & (g5149)) + ((!g1968) & (!g1970) & (g2509) & (!g2546) & (!g5149)) + ((!g1968) & (!g1970) & (g2509) & (g2546) & (g5149)) + ((!g1968) & (g1970) & (!g2509) & (!g2546) & (!g5149)) + ((!g1968) & (g1970) & (!g2509) & (!g2546) & (g5149)) + ((!g1968) & (g1970) & (g2509) & (!g2546) & (g5149)) + ((!g1968) & (g1970) & (g2509) & (g2546) & (!g5149)) + ((g1968) & (!g1970) & (!g2509) & (!g2546) & (!g5149)) + ((g1968) & (!g1970) & (!g2509) & (g2546) & (g5149)) + ((g1968) & (!g1970) & (g2509) & (!g2546) & (!g5149)) + ((g1968) & (!g1970) & (g2509) & (!g2546) & (g5149)) + ((g1968) & (g1970) & (!g2509) & (!g2546) & (g5149)) + ((g1968) & (g1970) & (!g2509) & (g2546) & (!g5149)) + ((g1968) & (g1970) & (g2509) & (g2546) & (!g5149)) + ((g1968) & (g1970) & (g2509) & (g2546) & (g5149)));
	assign g5182 = (((!g830) & (!g1914) & (!g2968) & (!g5180) & (!g5181) & (nonce[53])) + ((!g830) & (!g1914) & (!g2968) & (!g5180) & (g5181) & (nonce[53])) + ((!g830) & (!g1914) & (!g2968) & (g5180) & (!g5181) & (nonce[53])) + ((!g830) & (!g1914) & (!g2968) & (g5180) & (g5181) & (nonce[53])) + ((!g830) & (!g1914) & (g2968) & (!g5180) & (!g5181) & (nonce[53])) + ((!g830) & (!g1914) & (g2968) & (!g5180) & (g5181) & (nonce[53])) + ((!g830) & (!g1914) & (g2968) & (g5180) & (!g5181) & (nonce[53])) + ((!g830) & (!g1914) & (g2968) & (g5180) & (g5181) & (nonce[53])) + ((!g830) & (g1914) & (!g2968) & (!g5180) & (!g5181) & (nonce[53])) + ((!g830) & (g1914) & (!g2968) & (!g5180) & (g5181) & (nonce[53])) + ((!g830) & (g1914) & (!g2968) & (g5180) & (!g5181) & (nonce[53])) + ((!g830) & (g1914) & (!g2968) & (g5180) & (g5181) & (nonce[53])) + ((!g830) & (g1914) & (g2968) & (!g5180) & (!g5181) & (nonce[53])) + ((!g830) & (g1914) & (g2968) & (!g5180) & (g5181) & (nonce[53])) + ((!g830) & (g1914) & (g2968) & (g5180) & (!g5181) & (nonce[53])) + ((!g830) & (g1914) & (g2968) & (g5180) & (g5181) & (nonce[53])) + ((g830) & (!g1914) & (!g2968) & (!g5180) & (g5181) & (!nonce[53])) + ((g830) & (!g1914) & (!g2968) & (!g5180) & (g5181) & (nonce[53])) + ((g830) & (!g1914) & (!g2968) & (g5180) & (g5181) & (!nonce[53])) + ((g830) & (!g1914) & (!g2968) & (g5180) & (g5181) & (nonce[53])) + ((g830) & (!g1914) & (g2968) & (!g5180) & (!g5181) & (!nonce[53])) + ((g830) & (!g1914) & (g2968) & (!g5180) & (!g5181) & (nonce[53])) + ((g830) & (!g1914) & (g2968) & (g5180) & (!g5181) & (!nonce[53])) + ((g830) & (!g1914) & (g2968) & (g5180) & (!g5181) & (nonce[53])) + ((g830) & (g1914) & (!g2968) & (g5180) & (!g5181) & (!nonce[53])) + ((g830) & (g1914) & (!g2968) & (g5180) & (!g5181) & (nonce[53])) + ((g830) & (g1914) & (!g2968) & (g5180) & (g5181) & (!nonce[53])) + ((g830) & (g1914) & (!g2968) & (g5180) & (g5181) & (nonce[53])) + ((g830) & (g1914) & (g2968) & (!g5180) & (!g5181) & (!nonce[53])) + ((g830) & (g1914) & (g2968) & (!g5180) & (!g5181) & (nonce[53])) + ((g830) & (g1914) & (g2968) & (!g5180) & (g5181) & (!nonce[53])) + ((g830) & (g1914) & (g2968) & (!g5180) & (g5181) & (nonce[53])));
	assign g5183 = (((!g2566) & (g2578) & (!g3610)) + ((g2566) & (!g2578) & (!g3610)) + ((g2566) & (g2578) & (!g3610)) + ((g2566) & (g2578) & (g3610)));
	assign g5184 = (((!g1997) & (!g3592) & (!g2329)) + ((!g1997) & (g3592) & (g2329)) + ((g1997) & (!g3592) & (g2329)) + ((g1997) & (g3592) & (!g2329)));
	assign g5185 = (((!g1914) & (!g2614) & (!g2617) & (g5183) & (!g5184)) + ((!g1914) & (!g2614) & (!g2617) & (g5183) & (g5184)) + ((!g1914) & (!g2614) & (g2617) & (!g5183) & (!g5184)) + ((!g1914) & (!g2614) & (g2617) & (!g5183) & (g5184)) + ((!g1914) & (g2614) & (!g2617) & (!g5183) & (!g5184)) + ((!g1914) & (g2614) & (!g2617) & (!g5183) & (g5184)) + ((!g1914) & (g2614) & (g2617) & (g5183) & (!g5184)) + ((!g1914) & (g2614) & (g2617) & (g5183) & (g5184)) + ((g1914) & (!g2614) & (!g2617) & (!g5183) & (g5184)) + ((g1914) & (!g2614) & (!g2617) & (g5183) & (g5184)) + ((g1914) & (!g2614) & (g2617) & (!g5183) & (g5184)) + ((g1914) & (!g2614) & (g2617) & (g5183) & (g5184)) + ((g1914) & (g2614) & (!g2617) & (!g5183) & (g5184)) + ((g1914) & (g2614) & (!g2617) & (g5183) & (g5184)) + ((g1914) & (g2614) & (g2617) & (!g5183) & (g5184)) + ((g1914) & (g2614) & (g2617) & (g5183) & (g5184)));
	assign g5186 = (((!g830) & (!g2979) & (!g5185) & (key[245])) + ((!g830) & (!g2979) & (g5185) & (key[245])) + ((!g830) & (g2979) & (!g5185) & (key[245])) + ((!g830) & (g2979) & (g5185) & (key[245])) + ((g830) & (!g2979) & (g5185) & (!key[245])) + ((g830) & (!g2979) & (g5185) & (key[245])) + ((g830) & (g2979) & (!g5185) & (!key[245])) + ((g830) & (g2979) & (!g5185) & (key[245])));
	assign g5187 = (((!g2004) & (!g2006) & (!g2509) & (g2546) & (!g5139)) + ((!g2004) & (!g2006) & (!g2509) & (g2546) & (g5139)) + ((!g2004) & (!g2006) & (g2509) & (!g2546) & (!g5139)) + ((!g2004) & (!g2006) & (g2509) & (g2546) & (g5139)) + ((!g2004) & (g2006) & (!g2509) & (!g2546) & (!g5139)) + ((!g2004) & (g2006) & (!g2509) & (!g2546) & (g5139)) + ((!g2004) & (g2006) & (g2509) & (!g2546) & (g5139)) + ((!g2004) & (g2006) & (g2509) & (g2546) & (!g5139)) + ((g2004) & (!g2006) & (!g2509) & (!g2546) & (!g5139)) + ((g2004) & (!g2006) & (!g2509) & (g2546) & (g5139)) + ((g2004) & (!g2006) & (g2509) & (!g2546) & (!g5139)) + ((g2004) & (!g2006) & (g2509) & (!g2546) & (g5139)) + ((g2004) & (g2006) & (!g2509) & (!g2546) & (g5139)) + ((g2004) & (g2006) & (!g2509) & (g2546) & (!g5139)) + ((g2004) & (g2006) & (g2509) & (g2546) & (!g5139)) + ((g2004) & (g2006) & (g2509) & (g2546) & (g5139)));
	assign g5188 = (((!g2456) & (!g2535) & (!g2480) & (g2537) & (!g5141)) + ((!g2456) & (!g2535) & (!g2480) & (g2537) & (g5141)) + ((!g2456) & (!g2535) & (g2480) & (!g2537) & (!g5141)) + ((!g2456) & (!g2535) & (g2480) & (g2537) & (g5141)) + ((!g2456) & (g2535) & (!g2480) & (!g2537) & (!g5141)) + ((!g2456) & (g2535) & (!g2480) & (!g2537) & (g5141)) + ((!g2456) & (g2535) & (g2480) & (!g2537) & (g5141)) + ((!g2456) & (g2535) & (g2480) & (g2537) & (!g5141)) + ((g2456) & (!g2535) & (!g2480) & (!g2537) & (!g5141)) + ((g2456) & (!g2535) & (!g2480) & (g2537) & (g5141)) + ((g2456) & (!g2535) & (g2480) & (!g2537) & (!g5141)) + ((g2456) & (!g2535) & (g2480) & (!g2537) & (g5141)) + ((g2456) & (g2535) & (!g2480) & (!g2537) & (g5141)) + ((g2456) & (g2535) & (!g2480) & (g2537) & (!g5141)) + ((g2456) & (g2535) & (g2480) & (g2537) & (!g5141)) + ((g2456) & (g2535) & (g2480) & (g2537) & (g5141)));
	assign g5189 = (((!g830) & (!g1914) & (!g2985) & (!g5187) & (!g5188) & (key[213])) + ((!g830) & (!g1914) & (!g2985) & (!g5187) & (g5188) & (key[213])) + ((!g830) & (!g1914) & (!g2985) & (g5187) & (!g5188) & (key[213])) + ((!g830) & (!g1914) & (!g2985) & (g5187) & (g5188) & (key[213])) + ((!g830) & (!g1914) & (g2985) & (!g5187) & (!g5188) & (key[213])) + ((!g830) & (!g1914) & (g2985) & (!g5187) & (g5188) & (key[213])) + ((!g830) & (!g1914) & (g2985) & (g5187) & (!g5188) & (key[213])) + ((!g830) & (!g1914) & (g2985) & (g5187) & (g5188) & (key[213])) + ((!g830) & (g1914) & (!g2985) & (!g5187) & (!g5188) & (key[213])) + ((!g830) & (g1914) & (!g2985) & (!g5187) & (g5188) & (key[213])) + ((!g830) & (g1914) & (!g2985) & (g5187) & (!g5188) & (key[213])) + ((!g830) & (g1914) & (!g2985) & (g5187) & (g5188) & (key[213])) + ((!g830) & (g1914) & (g2985) & (!g5187) & (!g5188) & (key[213])) + ((!g830) & (g1914) & (g2985) & (!g5187) & (g5188) & (key[213])) + ((!g830) & (g1914) & (g2985) & (g5187) & (!g5188) & (key[213])) + ((!g830) & (g1914) & (g2985) & (g5187) & (g5188) & (key[213])) + ((g830) & (!g1914) & (!g2985) & (!g5187) & (g5188) & (!key[213])) + ((g830) & (!g1914) & (!g2985) & (!g5187) & (g5188) & (key[213])) + ((g830) & (!g1914) & (!g2985) & (g5187) & (g5188) & (!key[213])) + ((g830) & (!g1914) & (!g2985) & (g5187) & (g5188) & (key[213])) + ((g830) & (!g1914) & (g2985) & (!g5187) & (!g5188) & (!key[213])) + ((g830) & (!g1914) & (g2985) & (!g5187) & (!g5188) & (key[213])) + ((g830) & (!g1914) & (g2985) & (g5187) & (!g5188) & (!key[213])) + ((g830) & (!g1914) & (g2985) & (g5187) & (!g5188) & (key[213])) + ((g830) & (g1914) & (!g2985) & (g5187) & (!g5188) & (!key[213])) + ((g830) & (g1914) & (!g2985) & (g5187) & (!g5188) & (key[213])) + ((g830) & (g1914) & (!g2985) & (g5187) & (g5188) & (!key[213])) + ((g830) & (g1914) & (!g2985) & (g5187) & (g5188) & (key[213])) + ((g830) & (g1914) & (g2985) & (!g5187) & (!g5188) & (!key[213])) + ((g830) & (g1914) & (g2985) & (!g5187) & (!g5188) & (key[213])) + ((g830) & (g1914) & (g2985) & (!g5187) & (g5188) & (!key[213])) + ((g830) & (g1914) & (g2985) & (!g5187) & (g5188) & (key[213])));
	assign g5190 = (((!g2112) & (!g2120) & (g3856)) + ((!g2112) & (g2120) & (!g3856)) + ((g2112) & (!g2120) & (!g3856)) + ((g2112) & (g2120) & (g3856)));
	assign g5191 = (((!g3434) & (!g2314) & (g2337)) + ((!g3434) & (g2314) & (!g2337)) + ((!g3434) & (g2314) & (g2337)) + ((g3434) & (g2314) & (g2337)));
	assign g5192 = (((!g5191) & (!g2362) & (g2366)) + ((!g5191) & (g2362) & (!g2366)) + ((g5191) & (!g2362) & (!g2366)) + ((g5191) & (g2362) & (g2366)));
	assign g5193 = (((!g830) & (!g2999) & (!g6149) & (key[118])) + ((!g830) & (!g2999) & (g6149) & (key[118])) + ((!g830) & (g2999) & (!g6149) & (key[118])) + ((!g830) & (g2999) & (g6149) & (key[118])) + ((g830) & (!g2999) & (g6149) & (!key[118])) + ((g830) & (!g2999) & (g6149) & (key[118])) + ((g830) & (g2999) & (!g6149) & (!key[118])) + ((g830) & (g2999) & (!g6149) & (key[118])));
	assign g5194 = (((!g1982) & (g3535) & (g2110)) + ((g1982) & (!g3535) & (g2110)) + ((g1982) & (g3535) & (!g2110)) + ((g1982) & (g3535) & (g2110)));
	assign g5195 = (((g1914) & (!g1984) & (!g5194) & (g2156)) + ((g1914) & (!g1984) & (g5194) & (!g2156)) + ((g1914) & (g1984) & (!g5194) & (!g2156)) + ((g1914) & (g1984) & (g5194) & (g2156)));
	assign g5196 = (((!g1944) & (g2116) & (g3544)) + ((g1944) & (!g2116) & (g3544)) + ((g1944) & (g2116) & (!g3544)) + ((g1944) & (g2116) & (g3544)));
	assign g5197 = (((!g1914) & (!g1946) & (!g2147) & (g5196)) + ((!g1914) & (!g1946) & (g2147) & (!g5196)) + ((!g1914) & (g1946) & (!g2147) & (!g5196)) + ((!g1914) & (g1946) & (g2147) & (g5196)));
	assign g5198 = (((!g830) & (!g3003) & (!g5195) & (!g5197)) + ((!g830) & (!g3003) & (!g5195) & (g5197)) + ((!g830) & (!g3003) & (g5195) & (!g5197)) + ((!g830) & (!g3003) & (g5195) & (g5197)) + ((!g830) & (g3003) & (!g5195) & (!g5197)) + ((!g830) & (g3003) & (!g5195) & (g5197)) + ((!g830) & (g3003) & (g5195) & (!g5197)) + ((!g830) & (g3003) & (g5195) & (g5197)) + ((g830) & (!g3003) & (!g5195) & (g5197)) + ((g830) & (!g3003) & (g5195) & (!g5197)) + ((g830) & (!g3003) & (g5195) & (g5197)) + ((g830) & (g3003) & (!g5195) & (!g5197)));
	assign g5199 = (((!g1958) & (g2317) & (!g3576)) + ((g1958) & (!g2317) & (!g3576)) + ((g1958) & (g2317) & (!g3576)) + ((g1958) & (g2317) & (g3576)));
	assign g5200 = (((!g1960) & (!g2369) & (g5199)) + ((!g1960) & (g2369) & (!g5199)) + ((g1960) & (!g2369) & (!g5199)) + ((g1960) & (g2369) & (g5199)));
	assign g5201 = (((!g830) & (!g3005) & (!g6138) & (nonce[22])) + ((!g830) & (!g3005) & (g6138) & (nonce[22])) + ((!g830) & (g3005) & (!g6138) & (nonce[22])) + ((!g830) & (g3005) & (g6138) & (nonce[22])) + ((g830) & (!g3005) & (g6138) & (!nonce[22])) + ((g830) & (!g3005) & (g6138) & (nonce[22])) + ((g830) & (g3005) & (!g6138) & (!nonce[22])) + ((g830) & (g3005) & (!g6138) & (nonce[22])));
	assign g5202 = (((!g1997) & (!g3592) & (g2329)) + ((g1997) & (!g3592) & (!g2329)) + ((g1997) & (!g3592) & (g2329)) + ((g1997) & (g3592) & (g2329)));
	assign g5203 = (((!g1999) & (!g5202) & (g2371)) + ((!g1999) & (g5202) & (!g2371)) + ((g1999) & (!g5202) & (!g2371)) + ((g1999) & (g5202) & (g2371)));
	assign g5204 = (((!g830) & (!g3007) & (!g6127) & (key[246])) + ((!g830) & (!g3007) & (g6127) & (key[246])) + ((!g830) & (g3007) & (!g6127) & (key[246])) + ((!g830) & (g3007) & (g6127) & (key[246])) + ((g830) & (!g3007) & (g6127) & (!key[246])) + ((g830) & (!g3007) & (g6127) & (key[246])) + ((g830) & (g3007) & (!g6127) & (!key[246])) + ((g830) & (g3007) & (!g6127) & (key[246])));
	assign g5205 = (((!g2323) & (g2329) & (!g3642)) + ((g2323) & (!g2329) & (!g3642)) + ((g2323) & (g2329) & (!g3642)) + ((g2323) & (g2329) & (g3642)));
	assign g5206 = (((!g2356) & (!g2371) & (g5205)) + ((!g2356) & (g2371) & (!g5205)) + ((g2356) & (!g2371) & (!g5205)) + ((g2356) & (g2371) & (g5205)));
	assign g5207 = (((!g830) & (!g3009) & (!g6116) & (key[22])) + ((!g830) & (!g3009) & (g6116) & (key[22])) + ((!g830) & (g3009) & (!g6116) & (key[22])) + ((!g830) & (g3009) & (g6116) & (key[22])) + ((g830) & (!g3009) & (g6116) & (!key[22])) + ((g830) & (!g3009) & (g6116) & (key[22])) + ((g830) & (g3009) & (!g6116) & (!key[22])) + ((g830) & (g3009) & (!g6116) & (key[22])));
	assign g5208 = (((!g1996) & (g2334) & (!g3658)) + ((g1996) & (!g2334) & (!g3658)) + ((g1996) & (g2334) & (!g3658)) + ((g1996) & (g2334) & (g3658)));
	assign g5209 = (((!g1998) & (!g2358) & (g5208)) + ((!g1998) & (g2358) & (!g5208)) + ((g1998) & (!g2358) & (!g5208)) + ((g1998) & (g2358) & (g5208)));
	assign g8330 = (((!g5560) & (g5635) & (!g5210)) + ((!g5560) & (g5635) & (g5210)) + ((g5560) & (!g5635) & (g5210)) + ((g5560) & (g5635) & (g5210)));
	assign g5211 = (((!g830) & (!g3011) & (!g6105) & (g5210)) + ((!g830) & (!g3011) & (g6105) & (g5210)) + ((!g830) & (g3011) & (!g6105) & (g5210)) + ((!g830) & (g3011) & (g6105) & (g5210)) + ((g830) & (!g3011) & (g6105) & (!g5210)) + ((g830) & (!g3011) & (g6105) & (g5210)) + ((g830) & (g3011) & (!g6105) & (!g5210)) + ((g830) & (g3011) & (!g6105) & (g5210)));
	assign g5212 = (((!g2114) & (g2120) & (g3689)) + ((g2114) & (!g2120) & (g3689)) + ((g2114) & (g2120) & (!g3689)) + ((g2114) & (g2120) & (g3689)));
	assign g5213 = (((g1914) & (!g2137) & (!g2170) & (g5212)) + ((g1914) & (!g2137) & (g2170) & (!g5212)) + ((g1914) & (g2137) & (!g2170) & (!g5212)) + ((g1914) & (g2137) & (g2170) & (g5212)));
	assign g5214 = (((!g2104) & (g2125) & (g3699)) + ((g2104) & (!g2125) & (g3699)) + ((g2104) & (g2125) & (!g3699)) + ((g2104) & (g2125) & (g3699)));
	assign g5215 = (((!g1914) & (!g2153) & (!g2162) & (g5214)) + ((!g1914) & (!g2153) & (g2162) & (!g5214)) + ((!g1914) & (g2153) & (!g2162) & (!g5214)) + ((!g1914) & (g2153) & (g2162) & (g5214)));
	assign g5216 = (((g830) & (!g3013) & (!g5213) & (g5215)) + ((g830) & (!g3013) & (g5213) & (!g5215)) + ((g830) & (!g3013) & (g5213) & (g5215)) + ((g830) & (g3013) & (!g5213) & (!g5215)));
	assign g5217 = (((!g2012) & (!g2595) & (!g3718)) + ((!g2012) & (g2595) & (g3718)) + ((g2012) & (!g2595) & (g3718)) + ((g2012) & (g2595) & (!g3718)));
	assign g5218 = (((!g2569) & (!g2581) & (!g3735)) + ((!g2569) & (g2581) & (g3735)) + ((g2569) & (!g2581) & (g3735)) + ((g2569) & (g2581) & (!g3735)));
	assign g5219 = (((!g830) & (!g1914) & (!g3015) & (!g5217) & (!g5218) & (key[214])) + ((!g830) & (!g1914) & (!g3015) & (!g5217) & (g5218) & (key[214])) + ((!g830) & (!g1914) & (!g3015) & (g5217) & (!g5218) & (key[214])) + ((!g830) & (!g1914) & (!g3015) & (g5217) & (g5218) & (key[214])) + ((!g830) & (!g1914) & (g3015) & (!g5217) & (!g5218) & (key[214])) + ((!g830) & (!g1914) & (g3015) & (!g5217) & (g5218) & (key[214])) + ((!g830) & (!g1914) & (g3015) & (g5217) & (!g5218) & (key[214])) + ((!g830) & (!g1914) & (g3015) & (g5217) & (g5218) & (key[214])) + ((!g830) & (g1914) & (!g3015) & (!g5217) & (!g5218) & (key[214])) + ((!g830) & (g1914) & (!g3015) & (!g5217) & (g5218) & (key[214])) + ((!g830) & (g1914) & (!g3015) & (g5217) & (!g5218) & (key[214])) + ((!g830) & (g1914) & (!g3015) & (g5217) & (g5218) & (key[214])) + ((!g830) & (g1914) & (g3015) & (!g5217) & (!g5218) & (key[214])) + ((!g830) & (g1914) & (g3015) & (!g5217) & (g5218) & (key[214])) + ((!g830) & (g1914) & (g3015) & (g5217) & (!g5218) & (key[214])) + ((!g830) & (g1914) & (g3015) & (g5217) & (g5218) & (key[214])) + ((g830) & (!g1914) & (!g3015) & (!g5217) & (g5218) & (!key[214])) + ((g830) & (!g1914) & (!g3015) & (!g5217) & (g5218) & (key[214])) + ((g830) & (!g1914) & (!g3015) & (g5217) & (g5218) & (!key[214])) + ((g830) & (!g1914) & (!g3015) & (g5217) & (g5218) & (key[214])) + ((g830) & (!g1914) & (g3015) & (!g5217) & (!g5218) & (!key[214])) + ((g830) & (!g1914) & (g3015) & (!g5217) & (!g5218) & (key[214])) + ((g830) & (!g1914) & (g3015) & (g5217) & (!g5218) & (!key[214])) + ((g830) & (!g1914) & (g3015) & (g5217) & (!g5218) & (key[214])) + ((g830) & (g1914) & (!g3015) & (g5217) & (!g5218) & (!key[214])) + ((g830) & (g1914) & (!g3015) & (g5217) & (!g5218) & (key[214])) + ((g830) & (g1914) & (!g3015) & (g5217) & (g5218) & (!key[214])) + ((g830) & (g1914) & (!g3015) & (g5217) & (g5218) & (key[214])) + ((g830) & (g1914) & (g3015) & (!g5217) & (!g5218) & (!key[214])) + ((g830) & (g1914) & (g3015) & (!g5217) & (!g5218) & (key[214])) + ((g830) & (g1914) & (g3015) & (!g5217) & (g5218) & (!key[214])) + ((g830) & (g1914) & (g3015) & (!g5217) & (g5218) & (key[214])));
	assign g5220 = (((!g1959) & (g2337) & (!g3799)) + ((g1959) & (!g2337) & (!g3799)) + ((g1959) & (g2337) & (!g3799)) + ((g1959) & (g2337) & (g3799)));
	assign g5221 = (((!g1961) & (!g2366) & (g5220)) + ((!g1961) & (g2366) & (!g5220)) + ((g1961) & (!g2366) & (!g5220)) + ((g1961) & (g2366) & (g5220)));
	assign g5222 = (((!g830) & (!g3018) & (!g6094) & (key[150])) + ((!g830) & (!g3018) & (g6094) & (key[150])) + ((!g830) & (g3018) & (!g6094) & (key[150])) + ((!g830) & (g3018) & (g6094) & (key[150])) + ((g830) & (!g3018) & (g6094) & (!key[150])) + ((g830) & (!g3018) & (g6094) & (key[150])) + ((g830) & (g3018) & (!g6094) & (!key[150])) + ((g830) & (g3018) & (!g6094) & (key[150])));
	assign g5223 = (((!g2578) & (!g2581) & (!g3819)) + ((!g2578) & (g2581) & (g3819)) + ((g2578) & (!g2581) & (g3819)) + ((g2578) & (g2581) & (!g3819)));
	assign g5224 = (((!g1973) & (!g2595) & (!g3836)) + ((!g1973) & (g2595) & (g3836)) + ((g1973) & (!g2595) & (g3836)) + ((g1973) & (g2595) & (!g3836)));
	assign g5225 = (((!g830) & (!g1914) & (!g3020) & (!g5223) & (!g5224) & (nonce[54])) + ((!g830) & (!g1914) & (!g3020) & (!g5223) & (g5224) & (nonce[54])) + ((!g830) & (!g1914) & (!g3020) & (g5223) & (!g5224) & (nonce[54])) + ((!g830) & (!g1914) & (!g3020) & (g5223) & (g5224) & (nonce[54])) + ((!g830) & (!g1914) & (g3020) & (!g5223) & (!g5224) & (nonce[54])) + ((!g830) & (!g1914) & (g3020) & (!g5223) & (g5224) & (nonce[54])) + ((!g830) & (!g1914) & (g3020) & (g5223) & (!g5224) & (nonce[54])) + ((!g830) & (!g1914) & (g3020) & (g5223) & (g5224) & (nonce[54])) + ((!g830) & (g1914) & (!g3020) & (!g5223) & (!g5224) & (nonce[54])) + ((!g830) & (g1914) & (!g3020) & (!g5223) & (g5224) & (nonce[54])) + ((!g830) & (g1914) & (!g3020) & (g5223) & (!g5224) & (nonce[54])) + ((!g830) & (g1914) & (!g3020) & (g5223) & (g5224) & (nonce[54])) + ((!g830) & (g1914) & (g3020) & (!g5223) & (!g5224) & (nonce[54])) + ((!g830) & (g1914) & (g3020) & (!g5223) & (g5224) & (nonce[54])) + ((!g830) & (g1914) & (g3020) & (g5223) & (!g5224) & (nonce[54])) + ((!g830) & (g1914) & (g3020) & (g5223) & (g5224) & (nonce[54])) + ((g830) & (!g1914) & (!g3020) & (!g5223) & (g5224) & (!nonce[54])) + ((g830) & (!g1914) & (!g3020) & (!g5223) & (g5224) & (nonce[54])) + ((g830) & (!g1914) & (!g3020) & (g5223) & (g5224) & (!nonce[54])) + ((g830) & (!g1914) & (!g3020) & (g5223) & (g5224) & (nonce[54])) + ((g830) & (!g1914) & (g3020) & (!g5223) & (!g5224) & (!nonce[54])) + ((g830) & (!g1914) & (g3020) & (!g5223) & (!g5224) & (nonce[54])) + ((g830) & (!g1914) & (g3020) & (g5223) & (!g5224) & (!nonce[54])) + ((g830) & (!g1914) & (g3020) & (g5223) & (!g5224) & (nonce[54])) + ((g830) & (g1914) & (!g3020) & (g5223) & (!g5224) & (!nonce[54])) + ((g830) & (g1914) & (!g3020) & (g5223) & (!g5224) & (nonce[54])) + ((g830) & (g1914) & (!g3020) & (g5223) & (g5224) & (!nonce[54])) + ((g830) & (g1914) & (!g3020) & (g5223) & (g5224) & (nonce[54])) + ((g830) & (g1914) & (g3020) & (!g5223) & (!g5224) & (!nonce[54])) + ((g830) & (g1914) & (g3020) & (!g5223) & (!g5224) & (nonce[54])) + ((g830) & (g1914) & (g3020) & (!g5223) & (g5224) & (!nonce[54])) + ((g830) & (g1914) & (g3020) & (!g5223) & (g5224) & (nonce[54])));
	assign g5226 = (((!g2123) & (g2125) & (g3846)) + ((g2123) & (!g2125) & (g3846)) + ((g2123) & (g2125) & (!g3846)) + ((g2123) & (g2125) & (g3846)));
	assign g5227 = (((g1914) & (!g2150) & (!g2162) & (g5226)) + ((g1914) & (!g2150) & (g2162) & (!g5226)) + ((g1914) & (g2150) & (!g2162) & (!g5226)) + ((g1914) & (g2150) & (g2162) & (g5226)));
	assign g5228 = (((!g2112) & (g2120) & (g3856)) + ((g2112) & (!g2120) & (g3856)) + ((g2112) & (g2120) & (!g3856)) + ((g2112) & (g2120) & (g3856)));
	assign g5229 = (((!g1914) & (!g2167) & (!g2170) & (g5228)) + ((!g1914) & (!g2167) & (g2170) & (!g5228)) + ((!g1914) & (g2167) & (!g2170) & (!g5228)) + ((!g1914) & (g2167) & (g2170) & (g5228)));
	assign g5230 = (((g830) & (!g3022) & (!g5227) & (g5229)) + ((g830) & (!g3022) & (g5227) & (!g5229)) + ((g830) & (!g3022) & (g5227) & (g5229)) + ((g830) & (g3022) & (!g5227) & (!g5229)));
	assign g5231 = (((!g3630) & (g3631)) + ((g3630) & (!g3631)) + ((g3630) & (g3631)));
	assign g5232 = (((!g2356) & (!g2402) & (!g2371) & (g2408) & (!g5205)) + ((!g2356) & (!g2402) & (!g2371) & (g2408) & (g5205)) + ((!g2356) & (!g2402) & (g2371) & (!g2408) & (g5205)) + ((!g2356) & (!g2402) & (g2371) & (g2408) & (!g5205)) + ((!g2356) & (g2402) & (!g2371) & (!g2408) & (!g5205)) + ((!g2356) & (g2402) & (!g2371) & (!g2408) & (g5205)) + ((!g2356) & (g2402) & (g2371) & (!g2408) & (!g5205)) + ((!g2356) & (g2402) & (g2371) & (g2408) & (g5205)) + ((g2356) & (!g2402) & (!g2371) & (!g2408) & (g5205)) + ((g2356) & (!g2402) & (!g2371) & (g2408) & (!g5205)) + ((g2356) & (!g2402) & (g2371) & (!g2408) & (!g5205)) + ((g2356) & (!g2402) & (g2371) & (!g2408) & (g5205)) + ((g2356) & (g2402) & (!g2371) & (!g2408) & (!g5205)) + ((g2356) & (g2402) & (!g2371) & (g2408) & (g5205)) + ((g2356) & (g2402) & (g2371) & (g2408) & (!g5205)) + ((g2356) & (g2402) & (g2371) & (g2408) & (g5205)));
	assign g5233 = (((!g1914) & (!g2099) & (!g1370) & (!g5231) & (g5232)) + ((!g1914) & (!g2099) & (!g1370) & (g5231) & (g5232)) + ((!g1914) & (!g2099) & (g1370) & (!g5231) & (g5232)) + ((!g1914) & (!g2099) & (g1370) & (g5231) & (g5232)) + ((!g1914) & (g2099) & (!g1370) & (!g5231) & (g5232)) + ((!g1914) & (g2099) & (!g1370) & (g5231) & (g5232)) + ((!g1914) & (g2099) & (g1370) & (!g5231) & (g5232)) + ((!g1914) & (g2099) & (g1370) & (g5231) & (g5232)) + ((g1914) & (!g2099) & (!g1370) & (g5231) & (!g5232)) + ((g1914) & (!g2099) & (!g1370) & (g5231) & (g5232)) + ((g1914) & (!g2099) & (g1370) & (!g5231) & (!g5232)) + ((g1914) & (!g2099) & (g1370) & (!g5231) & (g5232)) + ((g1914) & (g2099) & (!g1370) & (!g5231) & (!g5232)) + ((g1914) & (g2099) & (!g1370) & (!g5231) & (g5232)) + ((g1914) & (g2099) & (g1370) & (g5231) & (!g5232)) + ((g1914) & (g2099) & (g1370) & (g5231) & (g5232)));
	assign g5234 = (((!g830) & (!g3031) & (!g5233) & (key[23])) + ((!g830) & (!g3031) & (g5233) & (key[23])) + ((!g830) & (g3031) & (!g5233) & (key[23])) + ((!g830) & (g3031) & (g5233) & (key[23])) + ((g830) & (!g3031) & (g5233) & (!key[23])) + ((g830) & (!g3031) & (g5233) & (key[23])) + ((g830) & (g3031) & (!g5233) & (!key[23])) + ((g830) & (g3031) & (!g5233) & (key[23])));
	assign g5235 = (((!g1984) & (!g1986) & (!g5194) & (!g2156) & (g2190)) + ((!g1984) & (!g1986) & (!g5194) & (g2156) & (g2190)) + ((!g1984) & (!g1986) & (g5194) & (!g2156) & (g2190)) + ((!g1984) & (!g1986) & (g5194) & (g2156) & (!g2190)) + ((!g1984) & (g1986) & (!g5194) & (!g2156) & (!g2190)) + ((!g1984) & (g1986) & (!g5194) & (g2156) & (!g2190)) + ((!g1984) & (g1986) & (g5194) & (!g2156) & (!g2190)) + ((!g1984) & (g1986) & (g5194) & (g2156) & (g2190)) + ((g1984) & (!g1986) & (!g5194) & (!g2156) & (g2190)) + ((g1984) & (!g1986) & (!g5194) & (g2156) & (!g2190)) + ((g1984) & (!g1986) & (g5194) & (!g2156) & (!g2190)) + ((g1984) & (!g1986) & (g5194) & (g2156) & (!g2190)) + ((g1984) & (g1986) & (!g5194) & (!g2156) & (!g2190)) + ((g1984) & (g1986) & (!g5194) & (g2156) & (g2190)) + ((g1984) & (g1986) & (g5194) & (!g2156) & (g2190)) + ((g1984) & (g1986) & (g5194) & (g2156) & (g2190)));
	assign g5236 = (((!g1946) & (!g1948) & (!g2147) & (g2196) & (!g5196)) + ((!g1946) & (!g1948) & (!g2147) & (g2196) & (g5196)) + ((!g1946) & (!g1948) & (g2147) & (!g2196) & (g5196)) + ((!g1946) & (!g1948) & (g2147) & (g2196) & (!g5196)) + ((!g1946) & (g1948) & (!g2147) & (!g2196) & (!g5196)) + ((!g1946) & (g1948) & (!g2147) & (!g2196) & (g5196)) + ((!g1946) & (g1948) & (g2147) & (!g2196) & (!g5196)) + ((!g1946) & (g1948) & (g2147) & (g2196) & (g5196)) + ((g1946) & (!g1948) & (!g2147) & (!g2196) & (g5196)) + ((g1946) & (!g1948) & (!g2147) & (g2196) & (!g5196)) + ((g1946) & (!g1948) & (g2147) & (!g2196) & (!g5196)) + ((g1946) & (!g1948) & (g2147) & (!g2196) & (g5196)) + ((g1946) & (g1948) & (!g2147) & (!g2196) & (!g5196)) + ((g1946) & (g1948) & (!g2147) & (g2196) & (g5196)) + ((g1946) & (g1948) & (g2147) & (g2196) & (!g5196)) + ((g1946) & (g1948) & (g2147) & (g2196) & (g5196)));
	assign g5237 = (((g830) & (!g1914) & (!g3038) & (!g5235) & (g5236)) + ((g830) & (!g1914) & (!g3038) & (g5235) & (g5236)) + ((g830) & (!g1914) & (g3038) & (!g5235) & (!g5236)) + ((g830) & (!g1914) & (g3038) & (g5235) & (!g5236)) + ((g830) & (g1914) & (!g3038) & (g5235) & (!g5236)) + ((g830) & (g1914) & (!g3038) & (g5235) & (g5236)) + ((g830) & (g1914) & (g3038) & (!g5235) & (!g5236)) + ((g830) & (g1914) & (g3038) & (!g5235) & (g5236)));
	assign g5238 = (((!g3678) & (g3679)) + ((g3678) & (!g3679)) + ((g3678) & (g3679)));
	assign g5239 = (((!g1998) & (!g2001) & (!g2358) & (g2413) & (!g5208)) + ((!g1998) & (!g2001) & (!g2358) & (g2413) & (g5208)) + ((!g1998) & (!g2001) & (g2358) & (!g2413) & (g5208)) + ((!g1998) & (!g2001) & (g2358) & (g2413) & (!g5208)) + ((!g1998) & (g2001) & (!g2358) & (!g2413) & (!g5208)) + ((!g1998) & (g2001) & (!g2358) & (!g2413) & (g5208)) + ((!g1998) & (g2001) & (g2358) & (!g2413) & (!g5208)) + ((!g1998) & (g2001) & (g2358) & (g2413) & (g5208)) + ((g1998) & (!g2001) & (!g2358) & (!g2413) & (g5208)) + ((g1998) & (!g2001) & (!g2358) & (g2413) & (!g5208)) + ((g1998) & (!g2001) & (g2358) & (!g2413) & (!g5208)) + ((g1998) & (!g2001) & (g2358) & (!g2413) & (g5208)) + ((g1998) & (g2001) & (!g2358) & (!g2413) & (!g5208)) + ((g1998) & (g2001) & (!g2358) & (g2413) & (g5208)) + ((g1998) & (g2001) & (g2358) & (g2413) & (!g5208)) + ((g1998) & (g2001) & (g2358) & (g2413) & (g5208)));
	assign g5240 = (((!g1914) & (!g2718) & (!g2728) & (g5238) & (!g5239)) + ((!g1914) & (!g2718) & (!g2728) & (g5238) & (g5239)) + ((!g1914) & (!g2718) & (g2728) & (!g5238) & (!g5239)) + ((!g1914) & (!g2718) & (g2728) & (!g5238) & (g5239)) + ((!g1914) & (g2718) & (!g2728) & (!g5238) & (!g5239)) + ((!g1914) & (g2718) & (!g2728) & (!g5238) & (g5239)) + ((!g1914) & (g2718) & (g2728) & (g5238) & (!g5239)) + ((!g1914) & (g2718) & (g2728) & (g5238) & (g5239)) + ((g1914) & (!g2718) & (!g2728) & (!g5238) & (g5239)) + ((g1914) & (!g2718) & (!g2728) & (g5238) & (g5239)) + ((g1914) & (!g2718) & (g2728) & (!g5238) & (g5239)) + ((g1914) & (!g2718) & (g2728) & (g5238) & (g5239)) + ((g1914) & (g2718) & (!g2728) & (!g5238) & (g5239)) + ((g1914) & (g2718) & (!g2728) & (g5238) & (g5239)) + ((g1914) & (g2718) & (g2728) & (!g5238) & (g5239)) + ((g1914) & (g2718) & (g2728) & (g5238) & (g5239)));
	assign g8331 = (((!g5560) & (g5636) & (!g5241)) + ((!g5560) & (g5636) & (g5241)) + ((g5560) & (!g5636) & (g5241)) + ((g5560) & (g5636) & (g5241)));
	assign g5242 = (((!g830) & (!g3041) & (!g5240) & (g5241)) + ((!g830) & (!g3041) & (g5240) & (g5241)) + ((!g830) & (g3041) & (!g5240) & (g5241)) + ((!g830) & (g3041) & (g5240) & (g5241)) + ((g830) & (!g3041) & (g5240) & (!g5241)) + ((g830) & (!g3041) & (g5240) & (g5241)) + ((g830) & (g3041) & (!g5240) & (!g5241)) + ((g830) & (g3041) & (!g5240) & (g5241)));
	assign g5243 = (((!g3787) & (g3788)) + ((g3787) & (!g3788)) + ((g3787) & (g3788)));
	assign g5244 = (((!g1961) & (!g1963) & (!g2366) & (g2416) & (!g5220)) + ((!g1961) & (!g1963) & (!g2366) & (g2416) & (g5220)) + ((!g1961) & (!g1963) & (g2366) & (!g2416) & (g5220)) + ((!g1961) & (!g1963) & (g2366) & (g2416) & (!g5220)) + ((!g1961) & (g1963) & (!g2366) & (!g2416) & (!g5220)) + ((!g1961) & (g1963) & (!g2366) & (!g2416) & (g5220)) + ((!g1961) & (g1963) & (g2366) & (!g2416) & (!g5220)) + ((!g1961) & (g1963) & (g2366) & (g2416) & (g5220)) + ((g1961) & (!g1963) & (!g2366) & (!g2416) & (g5220)) + ((g1961) & (!g1963) & (!g2366) & (g2416) & (!g5220)) + ((g1961) & (!g1963) & (g2366) & (!g2416) & (!g5220)) + ((g1961) & (!g1963) & (g2366) & (!g2416) & (g5220)) + ((g1961) & (g1963) & (!g2366) & (!g2416) & (!g5220)) + ((g1961) & (g1963) & (!g2366) & (g2416) & (g5220)) + ((g1961) & (g1963) & (g2366) & (g2416) & (!g5220)) + ((g1961) & (g1963) & (g2366) & (g2416) & (g5220)));
	assign g5245 = (((!g1914) & (!g2703) & (!g2723) & (!g5243) & (g5244)) + ((!g1914) & (!g2703) & (!g2723) & (g5243) & (g5244)) + ((!g1914) & (!g2703) & (g2723) & (!g5243) & (g5244)) + ((!g1914) & (!g2703) & (g2723) & (g5243) & (g5244)) + ((!g1914) & (g2703) & (!g2723) & (!g5243) & (g5244)) + ((!g1914) & (g2703) & (!g2723) & (g5243) & (g5244)) + ((!g1914) & (g2703) & (g2723) & (!g5243) & (g5244)) + ((!g1914) & (g2703) & (g2723) & (g5243) & (g5244)) + ((g1914) & (!g2703) & (!g2723) & (g5243) & (!g5244)) + ((g1914) & (!g2703) & (!g2723) & (g5243) & (g5244)) + ((g1914) & (!g2703) & (g2723) & (!g5243) & (!g5244)) + ((g1914) & (!g2703) & (g2723) & (!g5243) & (g5244)) + ((g1914) & (g2703) & (!g2723) & (!g5243) & (!g5244)) + ((g1914) & (g2703) & (!g2723) & (!g5243) & (g5244)) + ((g1914) & (g2703) & (g2723) & (g5243) & (!g5244)) + ((g1914) & (g2703) & (g2723) & (g5243) & (g5244)));
	assign g5246 = (((!g830) & (!g3044) & (!g5245) & (key[151])) + ((!g830) & (!g3044) & (g5245) & (key[151])) + ((!g830) & (g3044) & (!g5245) & (key[151])) + ((!g830) & (g3044) & (g5245) & (key[151])) + ((g830) & (!g3044) & (g5245) & (!key[151])) + ((g830) & (!g3044) & (g5245) & (key[151])) + ((g830) & (g3044) & (!g5245) & (!key[151])) + ((g830) & (g3044) & (!g5245) & (key[151])));
	assign g5247 = (((!g3453) & (g3454)) + ((g3453) & (!g3454)) + ((g3453) & (g3454)));
	assign g5248 = (((!g5191) & (!g2362) & (!g2366) & (!g2393) & (g2416)) + ((!g5191) & (!g2362) & (!g2366) & (g2393) & (!g2416)) + ((!g5191) & (!g2362) & (g2366) & (!g2393) & (g2416)) + ((!g5191) & (!g2362) & (g2366) & (g2393) & (!g2416)) + ((!g5191) & (g2362) & (!g2366) & (!g2393) & (g2416)) + ((!g5191) & (g2362) & (!g2366) & (g2393) & (!g2416)) + ((!g5191) & (g2362) & (g2366) & (!g2393) & (!g2416)) + ((!g5191) & (g2362) & (g2366) & (g2393) & (g2416)) + ((g5191) & (!g2362) & (!g2366) & (!g2393) & (g2416)) + ((g5191) & (!g2362) & (!g2366) & (g2393) & (!g2416)) + ((g5191) & (!g2362) & (g2366) & (!g2393) & (!g2416)) + ((g5191) & (!g2362) & (g2366) & (g2393) & (g2416)) + ((g5191) & (g2362) & (!g2366) & (!g2393) & (!g2416)) + ((g5191) & (g2362) & (!g2366) & (g2393) & (g2416)) + ((g5191) & (g2362) & (g2366) & (!g2393) & (!g2416)) + ((g5191) & (g2362) & (g2366) & (g2393) & (g2416)));
	assign g5249 = (((!g1914) & (!g2101) & (!g1370) & (g5247) & (!g5248)) + ((!g1914) & (!g2101) & (!g1370) & (g5247) & (g5248)) + ((!g1914) & (!g2101) & (g1370) & (!g5247) & (!g5248)) + ((!g1914) & (!g2101) & (g1370) & (!g5247) & (g5248)) + ((!g1914) & (g2101) & (!g1370) & (!g5247) & (!g5248)) + ((!g1914) & (g2101) & (!g1370) & (!g5247) & (g5248)) + ((!g1914) & (g2101) & (g1370) & (g5247) & (!g5248)) + ((!g1914) & (g2101) & (g1370) & (g5247) & (g5248)) + ((g1914) & (!g2101) & (!g1370) & (!g5247) & (g5248)) + ((g1914) & (!g2101) & (!g1370) & (g5247) & (g5248)) + ((g1914) & (!g2101) & (g1370) & (!g5247) & (g5248)) + ((g1914) & (!g2101) & (g1370) & (g5247) & (g5248)) + ((g1914) & (g2101) & (!g1370) & (!g5247) & (g5248)) + ((g1914) & (g2101) & (!g1370) & (g5247) & (g5248)) + ((g1914) & (g2101) & (g1370) & (!g5247) & (g5248)) + ((g1914) & (g2101) & (g1370) & (g5247) & (g5248)));
	assign g5250 = (((!g830) & (!g3047) & (!g5249) & (key[119])) + ((!g830) & (!g3047) & (g5249) & (key[119])) + ((!g830) & (g3047) & (!g5249) & (key[119])) + ((!g830) & (g3047) & (g5249) & (key[119])) + ((g830) & (!g3047) & (g5249) & (!key[119])) + ((g830) & (!g3047) & (g5249) & (key[119])) + ((g830) & (g3047) & (!g5249) & (!key[119])) + ((g830) & (g3047) & (!g5249) & (key[119])));
	assign g5251 = (((!g3564) & (g3565)) + ((g3564) & (!g3565)) + ((g3564) & (g3565)));
	assign g5252 = (((!g1960) & (!g1962) & (!g2369) & (g2396) & (!g5199)) + ((!g1960) & (!g1962) & (!g2369) & (g2396) & (g5199)) + ((!g1960) & (!g1962) & (g2369) & (!g2396) & (g5199)) + ((!g1960) & (!g1962) & (g2369) & (g2396) & (!g5199)) + ((!g1960) & (g1962) & (!g2369) & (!g2396) & (!g5199)) + ((!g1960) & (g1962) & (!g2369) & (!g2396) & (g5199)) + ((!g1960) & (g1962) & (g2369) & (!g2396) & (!g5199)) + ((!g1960) & (g1962) & (g2369) & (g2396) & (g5199)) + ((g1960) & (!g1962) & (!g2369) & (!g2396) & (g5199)) + ((g1960) & (!g1962) & (!g2369) & (g2396) & (!g5199)) + ((g1960) & (!g1962) & (g2369) & (!g2396) & (!g5199)) + ((g1960) & (!g1962) & (g2369) & (!g2396) & (g5199)) + ((g1960) & (g1962) & (!g2369) & (!g2396) & (!g5199)) + ((g1960) & (g1962) & (!g2369) & (g2396) & (g5199)) + ((g1960) & (g1962) & (g2369) & (g2396) & (!g5199)) + ((g1960) & (g1962) & (g2369) & (g2396) & (g5199)));
	assign g5253 = (((!g1914) & (!g2690) & (!g5251) & (!g2728) & (g5252)) + ((!g1914) & (!g2690) & (!g5251) & (g2728) & (g5252)) + ((!g1914) & (!g2690) & (g5251) & (!g2728) & (g5252)) + ((!g1914) & (!g2690) & (g5251) & (g2728) & (g5252)) + ((!g1914) & (g2690) & (!g5251) & (!g2728) & (g5252)) + ((!g1914) & (g2690) & (!g5251) & (g2728) & (g5252)) + ((!g1914) & (g2690) & (g5251) & (!g2728) & (g5252)) + ((!g1914) & (g2690) & (g5251) & (g2728) & (g5252)) + ((g1914) & (!g2690) & (!g5251) & (g2728) & (!g5252)) + ((g1914) & (!g2690) & (!g5251) & (g2728) & (g5252)) + ((g1914) & (!g2690) & (g5251) & (!g2728) & (!g5252)) + ((g1914) & (!g2690) & (g5251) & (!g2728) & (g5252)) + ((g1914) & (g2690) & (!g5251) & (!g2728) & (!g5252)) + ((g1914) & (g2690) & (!g5251) & (!g2728) & (g5252)) + ((g1914) & (g2690) & (g5251) & (g2728) & (!g5252)) + ((g1914) & (g2690) & (g5251) & (g2728) & (g5252)));
	assign g5254 = (((!g830) & (!g3050) & (!g5253) & (nonce[23])) + ((!g830) & (!g3050) & (g5253) & (nonce[23])) + ((!g830) & (g3050) & (!g5253) & (nonce[23])) + ((!g830) & (g3050) & (g5253) & (nonce[23])) + ((g830) & (!g3050) & (g5253) & (!nonce[23])) + ((g830) & (!g3050) & (g5253) & (nonce[23])) + ((g830) & (g3050) & (!g5253) & (!nonce[23])) + ((g830) & (g3050) & (!g5253) & (nonce[23])));
	assign g5255 = (((!g2137) & (!g2194) & (!g2170) & (g2200) & (!g5212)) + ((!g2137) & (!g2194) & (!g2170) & (g2200) & (g5212)) + ((!g2137) & (!g2194) & (g2170) & (!g2200) & (g5212)) + ((!g2137) & (!g2194) & (g2170) & (g2200) & (!g5212)) + ((!g2137) & (g2194) & (!g2170) & (!g2200) & (!g5212)) + ((!g2137) & (g2194) & (!g2170) & (!g2200) & (g5212)) + ((!g2137) & (g2194) & (g2170) & (!g2200) & (!g5212)) + ((!g2137) & (g2194) & (g2170) & (g2200) & (g5212)) + ((g2137) & (!g2194) & (!g2170) & (!g2200) & (g5212)) + ((g2137) & (!g2194) & (!g2170) & (g2200) & (!g5212)) + ((g2137) & (!g2194) & (g2170) & (!g2200) & (!g5212)) + ((g2137) & (!g2194) & (g2170) & (!g2200) & (g5212)) + ((g2137) & (g2194) & (!g2170) & (!g2200) & (!g5212)) + ((g2137) & (g2194) & (!g2170) & (g2200) & (g5212)) + ((g2137) & (g2194) & (g2170) & (g2200) & (!g5212)) + ((g2137) & (g2194) & (g2170) & (g2200) & (g5212)));
	assign g5256 = (((!g2153) & (!g2184) & (!g2162) & (g2205) & (!g5214)) + ((!g2153) & (!g2184) & (!g2162) & (g2205) & (g5214)) + ((!g2153) & (!g2184) & (g2162) & (!g2205) & (g5214)) + ((!g2153) & (!g2184) & (g2162) & (g2205) & (!g5214)) + ((!g2153) & (g2184) & (!g2162) & (!g2205) & (!g5214)) + ((!g2153) & (g2184) & (!g2162) & (!g2205) & (g5214)) + ((!g2153) & (g2184) & (g2162) & (!g2205) & (!g5214)) + ((!g2153) & (g2184) & (g2162) & (g2205) & (g5214)) + ((g2153) & (!g2184) & (!g2162) & (!g2205) & (g5214)) + ((g2153) & (!g2184) & (!g2162) & (g2205) & (!g5214)) + ((g2153) & (!g2184) & (g2162) & (!g2205) & (!g5214)) + ((g2153) & (!g2184) & (g2162) & (!g2205) & (g5214)) + ((g2153) & (g2184) & (!g2162) & (!g2205) & (!g5214)) + ((g2153) & (g2184) & (!g2162) & (g2205) & (g5214)) + ((g2153) & (g2184) & (g2162) & (g2205) & (!g5214)) + ((g2153) & (g2184) & (g2162) & (g2205) & (g5214)));
	assign g5257 = (((g830) & (!g1914) & (!g3053) & (!g5255) & (g5256)) + ((g830) & (!g1914) & (!g3053) & (g5255) & (g5256)) + ((g830) & (!g1914) & (g3053) & (!g5255) & (!g5256)) + ((g830) & (!g1914) & (g3053) & (g5255) & (!g5256)) + ((g830) & (g1914) & (!g3053) & (g5255) & (!g5256)) + ((g830) & (g1914) & (!g3053) & (g5255) & (g5256)) + ((g830) & (g1914) & (g3053) & (!g5255) & (!g5256)) + ((g830) & (g1914) & (g3053) & (!g5255) & (g5256)));
	assign g5258 = (((!g2578) & (g2581) & (!g3819)) + ((g2578) & (!g2581) & (!g3819)) + ((g2578) & (g2581) & (!g3819)) + ((g2578) & (g2581) & (g3819)));
	assign g5259 = (((g1914) & (!g2617) & (!g2629) & (g5258)) + ((g1914) & (!g2617) & (g2629) & (!g5258)) + ((g1914) & (g2617) & (!g2629) & (!g5258)) + ((g1914) & (g2617) & (g2629) & (g5258)));
	assign g5260 = (((!g1973) & (g2595) & (!g3836)) + ((g1973) & (!g2595) & (!g3836)) + ((g1973) & (g2595) & (!g3836)) + ((g1973) & (g2595) & (g3836)));
	assign g5261 = (((!g1914) & (!g1976) & (!g2643) & (g5260)) + ((!g1914) & (!g1976) & (g2643) & (!g5260)) + ((!g1914) & (g1976) & (!g2643) & (!g5260)) + ((!g1914) & (g1976) & (g2643) & (g5260)));
	assign g5262 = (((!g830) & (!g3056) & (!g5259) & (!g5261) & (nonce[55])) + ((!g830) & (!g3056) & (!g5259) & (g5261) & (nonce[55])) + ((!g830) & (!g3056) & (g5259) & (!g5261) & (nonce[55])) + ((!g830) & (!g3056) & (g5259) & (g5261) & (nonce[55])) + ((!g830) & (g3056) & (!g5259) & (!g5261) & (nonce[55])) + ((!g830) & (g3056) & (!g5259) & (g5261) & (nonce[55])) + ((!g830) & (g3056) & (g5259) & (!g5261) & (nonce[55])) + ((!g830) & (g3056) & (g5259) & (g5261) & (nonce[55])) + ((g830) & (!g3056) & (!g5259) & (g5261) & (!nonce[55])) + ((g830) & (!g3056) & (!g5259) & (g5261) & (nonce[55])) + ((g830) & (!g3056) & (g5259) & (!g5261) & (!nonce[55])) + ((g830) & (!g3056) & (g5259) & (!g5261) & (nonce[55])) + ((g830) & (!g3056) & (g5259) & (g5261) & (!nonce[55])) + ((g830) & (!g3056) & (g5259) & (g5261) & (nonce[55])) + ((g830) & (g3056) & (!g5259) & (!g5261) & (!nonce[55])) + ((g830) & (g3056) & (!g5259) & (!g5261) & (nonce[55])));
	assign g5263 = (((!g3611) & (g3612)) + ((g3611) & (!g3612)) + ((g3611) & (g3612)));
	assign g5264 = (((!g1999) & (!g2002) & (!g5202) & (!g2371) & (g2408)) + ((!g1999) & (!g2002) & (!g5202) & (g2371) & (g2408)) + ((!g1999) & (!g2002) & (g5202) & (!g2371) & (g2408)) + ((!g1999) & (!g2002) & (g5202) & (g2371) & (!g2408)) + ((!g1999) & (g2002) & (!g5202) & (!g2371) & (!g2408)) + ((!g1999) & (g2002) & (!g5202) & (g2371) & (!g2408)) + ((!g1999) & (g2002) & (g5202) & (!g2371) & (!g2408)) + ((!g1999) & (g2002) & (g5202) & (g2371) & (g2408)) + ((g1999) & (!g2002) & (!g5202) & (!g2371) & (g2408)) + ((g1999) & (!g2002) & (!g5202) & (g2371) & (!g2408)) + ((g1999) & (!g2002) & (g5202) & (!g2371) & (!g2408)) + ((g1999) & (!g2002) & (g5202) & (g2371) & (!g2408)) + ((g1999) & (g2002) & (!g5202) & (!g2371) & (!g2408)) + ((g1999) & (g2002) & (!g5202) & (g2371) & (g2408)) + ((g1999) & (g2002) & (g5202) & (!g2371) & (g2408)) + ((g1999) & (g2002) & (g5202) & (g2371) & (g2408)));
	assign g5265 = (((!g1914) & (!g2703) & (!g2708) & (g5263) & (!g5264)) + ((!g1914) & (!g2703) & (!g2708) & (g5263) & (g5264)) + ((!g1914) & (!g2703) & (g2708) & (!g5263) & (!g5264)) + ((!g1914) & (!g2703) & (g2708) & (!g5263) & (g5264)) + ((!g1914) & (g2703) & (!g2708) & (!g5263) & (!g5264)) + ((!g1914) & (g2703) & (!g2708) & (!g5263) & (g5264)) + ((!g1914) & (g2703) & (g2708) & (g5263) & (!g5264)) + ((!g1914) & (g2703) & (g2708) & (g5263) & (g5264)) + ((g1914) & (!g2703) & (!g2708) & (!g5263) & (g5264)) + ((g1914) & (!g2703) & (!g2708) & (g5263) & (g5264)) + ((g1914) & (!g2703) & (g2708) & (!g5263) & (g5264)) + ((g1914) & (!g2703) & (g2708) & (g5263) & (g5264)) + ((g1914) & (g2703) & (!g2708) & (!g5263) & (g5264)) + ((g1914) & (g2703) & (!g2708) & (g5263) & (g5264)) + ((g1914) & (g2703) & (g2708) & (!g5263) & (g5264)) + ((g1914) & (g2703) & (g2708) & (g5263) & (g5264)));
	assign g5266 = (((!g830) & (!g3061) & (!g5265) & (key[247])) + ((!g830) & (!g3061) & (g5265) & (key[247])) + ((!g830) & (g3061) & (!g5265) & (key[247])) + ((!g830) & (g3061) & (g5265) & (key[247])) + ((g830) & (!g3061) & (g5265) & (!key[247])) + ((g830) & (!g3061) & (g5265) & (key[247])) + ((g830) & (g3061) & (!g5265) & (!key[247])) + ((g830) & (g3061) & (!g5265) & (key[247])));
	assign g5267 = (((!g2012) & (g2595) & (!g3718)) + ((g2012) & (!g2595) & (!g3718)) + ((g2012) & (g2595) & (!g3718)) + ((g2012) & (g2595) & (g3718)));
	assign g5268 = (((g1914) & (!g2014) & (!g2643) & (g5267)) + ((g1914) & (!g2014) & (g2643) & (!g5267)) + ((g1914) & (g2014) & (!g2643) & (!g5267)) + ((g1914) & (g2014) & (g2643) & (g5267)));
	assign g5269 = (((!g2569) & (g2581) & (!g3735)) + ((g2569) & (!g2581) & (!g3735)) + ((g2569) & (g2581) & (!g3735)) + ((g2569) & (g2581) & (g3735)));
	assign g5270 = (((!g1914) & (!g2626) & (!g2629) & (g5269)) + ((!g1914) & (!g2626) & (g2629) & (!g5269)) + ((!g1914) & (g2626) & (!g2629) & (!g5269)) + ((!g1914) & (g2626) & (g2629) & (g5269)));
	assign g5271 = (((!g830) & (!g3064) & (!g5268) & (!g5270) & (key[215])) + ((!g830) & (!g3064) & (!g5268) & (g5270) & (key[215])) + ((!g830) & (!g3064) & (g5268) & (!g5270) & (key[215])) + ((!g830) & (!g3064) & (g5268) & (g5270) & (key[215])) + ((!g830) & (g3064) & (!g5268) & (!g5270) & (key[215])) + ((!g830) & (g3064) & (!g5268) & (g5270) & (key[215])) + ((!g830) & (g3064) & (g5268) & (!g5270) & (key[215])) + ((!g830) & (g3064) & (g5268) & (g5270) & (key[215])) + ((g830) & (!g3064) & (!g5268) & (g5270) & (!key[215])) + ((g830) & (!g3064) & (!g5268) & (g5270) & (key[215])) + ((g830) & (!g3064) & (g5268) & (!g5270) & (!key[215])) + ((g830) & (!g3064) & (g5268) & (!g5270) & (key[215])) + ((g830) & (!g3064) & (g5268) & (g5270) & (!key[215])) + ((g830) & (!g3064) & (g5268) & (g5270) & (key[215])) + ((g830) & (g3064) & (!g5268) & (!g5270) & (!key[215])) + ((g830) & (g3064) & (!g5268) & (!g5270) & (key[215])));
	assign g5272 = (((!g2150) & (!g2203) & (!g2162) & (g2205) & (!g5226)) + ((!g2150) & (!g2203) & (!g2162) & (g2205) & (g5226)) + ((!g2150) & (!g2203) & (g2162) & (!g2205) & (g5226)) + ((!g2150) & (!g2203) & (g2162) & (g2205) & (!g5226)) + ((!g2150) & (g2203) & (!g2162) & (!g2205) & (!g5226)) + ((!g2150) & (g2203) & (!g2162) & (!g2205) & (g5226)) + ((!g2150) & (g2203) & (g2162) & (!g2205) & (!g5226)) + ((!g2150) & (g2203) & (g2162) & (g2205) & (g5226)) + ((g2150) & (!g2203) & (!g2162) & (!g2205) & (g5226)) + ((g2150) & (!g2203) & (!g2162) & (g2205) & (!g5226)) + ((g2150) & (!g2203) & (g2162) & (!g2205) & (!g5226)) + ((g2150) & (!g2203) & (g2162) & (!g2205) & (g5226)) + ((g2150) & (g2203) & (!g2162) & (!g2205) & (!g5226)) + ((g2150) & (g2203) & (!g2162) & (g2205) & (g5226)) + ((g2150) & (g2203) & (g2162) & (g2205) & (!g5226)) + ((g2150) & (g2203) & (g2162) & (g2205) & (g5226)));
	assign g5273 = (((!g2167) & (!g2192) & (!g2170) & (g2200) & (!g5228)) + ((!g2167) & (!g2192) & (!g2170) & (g2200) & (g5228)) + ((!g2167) & (!g2192) & (g2170) & (!g2200) & (g5228)) + ((!g2167) & (!g2192) & (g2170) & (g2200) & (!g5228)) + ((!g2167) & (g2192) & (!g2170) & (!g2200) & (!g5228)) + ((!g2167) & (g2192) & (!g2170) & (!g2200) & (g5228)) + ((!g2167) & (g2192) & (g2170) & (!g2200) & (!g5228)) + ((!g2167) & (g2192) & (g2170) & (g2200) & (g5228)) + ((g2167) & (!g2192) & (!g2170) & (!g2200) & (g5228)) + ((g2167) & (!g2192) & (!g2170) & (g2200) & (!g5228)) + ((g2167) & (!g2192) & (g2170) & (!g2200) & (!g5228)) + ((g2167) & (!g2192) & (g2170) & (!g2200) & (g5228)) + ((g2167) & (g2192) & (!g2170) & (!g2200) & (!g5228)) + ((g2167) & (g2192) & (!g2170) & (g2200) & (g5228)) + ((g2167) & (g2192) & (g2170) & (g2200) & (!g5228)) + ((g2167) & (g2192) & (g2170) & (g2200) & (g5228)));
	assign g5274 = (((g830) & (!g1914) & (!g3067) & (!g5272) & (g5273)) + ((g830) & (!g1914) & (!g3067) & (g5272) & (g5273)) + ((g830) & (!g1914) & (g3067) & (!g5272) & (!g5273)) + ((g830) & (!g1914) & (g3067) & (g5272) & (!g5273)) + ((g830) & (g1914) & (!g3067) & (g5272) & (!g5273)) + ((g830) & (g1914) & (!g3067) & (g5272) & (g5273)) + ((g830) & (g1914) & (g3067) & (!g5272) & (!g5273)) + ((g830) & (g1914) & (g3067) & (!g5272) & (g5273)));
	assign g5275 = (((!g3436) & (!g3437)));
	assign g5276 = (((!g5275) & (!g2474) & (!g2486)) + ((!g5275) & (g2474) & (g2486)) + ((g5275) & (!g2474) & (g2486)) + ((g5275) & (g2474) & (!g2486)));
	assign g5277 = (((!g830) & (!g3074) & (!g6083) & (key[120])) + ((!g830) & (!g3074) & (g6083) & (key[120])) + ((!g830) & (g3074) & (!g6083) & (key[120])) + ((!g830) & (g3074) & (g6083) & (key[120])) + ((g830) & (!g3074) & (g6083) & (!key[120])) + ((g830) & (!g3074) & (g6083) & (key[120])) + ((g830) & (g3074) & (!g6083) & (!key[120])) + ((g830) & (g3074) & (!g6083) & (key[120])));
	assign g5278 = (((!g3537) & (!g3538)));
	assign g5279 = (((g1914) & (!g1991) & (!g5278) & (!g2236)) + ((g1914) & (!g1991) & (g5278) & (g2236)) + ((g1914) & (g1991) & (!g5278) & (g2236)) + ((g1914) & (g1991) & (g5278) & (!g2236)));
	assign g5280 = (((!g3546) & (!g3547)));
	assign g5281 = (((!g1914) & (!g1953) & (!g2227) & (!g5280)) + ((!g1914) & (!g1953) & (g2227) & (g5280)) + ((!g1914) & (g1953) & (!g2227) & (g5280)) + ((!g1914) & (g1953) & (g2227) & (!g5280)));
	assign g5282 = (((!g830) & (!g3078) & (!g5279) & (!g5281)) + ((!g830) & (!g3078) & (!g5279) & (g5281)) + ((!g830) & (!g3078) & (g5279) & (!g5281)) + ((!g830) & (!g3078) & (g5279) & (g5281)) + ((!g830) & (g3078) & (!g5279) & (!g5281)) + ((!g830) & (g3078) & (!g5279) & (g5281)) + ((!g830) & (g3078) & (g5279) & (!g5281)) + ((!g830) & (g3078) & (g5279) & (g5281)) + ((g830) & (!g3078) & (!g5279) & (g5281)) + ((g830) & (!g3078) & (g5279) & (!g5281)) + ((g830) & (!g3078) & (g5279) & (g5281)) + ((g830) & (g3078) & (!g5279) & (!g5281)));
	assign g5283 = (((!g3578) & (!g3579)));
	assign g5284 = (((!g1967) & (!g2497) & (!g5283)) + ((!g1967) & (g2497) & (g5283)) + ((g1967) & (!g2497) & (g5283)) + ((g1967) & (g2497) & (!g5283)));
	assign g5285 = (((!g830) & (!g3080) & (!g6072) & (nonce[24])) + ((!g830) & (!g3080) & (g6072) & (nonce[24])) + ((!g830) & (g3080) & (!g6072) & (nonce[24])) + ((!g830) & (g3080) & (g6072) & (nonce[24])) + ((g830) & (!g3080) & (g6072) & (!nonce[24])) + ((g830) & (!g3080) & (g6072) & (nonce[24])) + ((g830) & (g3080) & (!g6072) & (!nonce[24])) + ((g830) & (g3080) & (!g6072) & (nonce[24])));
	assign g5286 = (((!g3594) & (!g3595)));
	assign g5287 = (((!g2004) & (!g5286) & (!g2503)) + ((!g2004) & (g5286) & (g2503)) + ((g2004) & (!g5286) & (g2503)) + ((g2004) & (g5286) & (!g2503)));
	assign g5288 = (((!g830) & (!g3082) & (!g6061) & (key[248])) + ((!g830) & (!g3082) & (g6061) & (key[248])) + ((!g830) & (g3082) & (!g6061) & (key[248])) + ((!g830) & (g3082) & (g6061) & (key[248])) + ((g830) & (!g3082) & (g6061) & (!key[248])) + ((g830) & (!g3082) & (g6061) & (key[248])) + ((g830) & (g3082) & (!g6061) & (!key[248])) + ((g830) & (g3082) & (!g6061) & (key[248])));
	assign g5289 = (((!g3644) & (!g3645)));
	assign g5290 = (((!g2456) & (!g2503) & (!g5289)) + ((!g2456) & (g2503) & (g5289)) + ((g2456) & (!g2503) & (g5289)) + ((g2456) & (g2503) & (!g5289)));
	assign g5291 = (((!g830) & (!g3084) & (!g6050) & (key[24])) + ((!g830) & (!g3084) & (g6050) & (key[24])) + ((!g830) & (g3084) & (!g6050) & (key[24])) + ((!g830) & (g3084) & (g6050) & (key[24])) + ((g830) & (!g3084) & (g6050) & (!key[24])) + ((g830) & (!g3084) & (g6050) & (key[24])) + ((g830) & (g3084) & (!g6050) & (!key[24])) + ((g830) & (g3084) & (!g6050) & (key[24])));
	assign g5292 = (((!g3660) & (!g3661)));
	assign g5293 = (((!g2003) & (!g2462) & (!g5292)) + ((!g2003) & (g2462) & (g5292)) + ((g2003) & (!g2462) & (g5292)) + ((g2003) & (g2462) & (!g5292)));
	assign g8332 = (((!g5560) & (g5638) & (!g5294)) + ((!g5560) & (g5638) & (g5294)) + ((g5560) & (!g5638) & (g5294)) + ((g5560) & (g5638) & (g5294)));
	assign g5295 = (((!g830) & (!g3086) & (!g6039) & (g5294)) + ((!g830) & (!g3086) & (g6039) & (g5294)) + ((!g830) & (g3086) & (!g6039) & (g5294)) + ((!g830) & (g3086) & (g6039) & (g5294)) + ((g830) & (!g3086) & (g6039) & (!g5294)) + ((g830) & (!g3086) & (g6039) & (g5294)) + ((g830) & (g3086) & (!g6039) & (!g5294)) + ((g830) & (g3086) & (!g6039) & (g5294)));
	assign g5296 = (((!g3691) & (!g3692)));
	assign g5297 = (((g1914) & (!g2217) & (!g2250) & (!g5296)) + ((g1914) & (!g2217) & (g2250) & (g5296)) + ((g1914) & (g2217) & (!g2250) & (g5296)) + ((g1914) & (g2217) & (g2250) & (!g5296)));
	assign g5298 = (((!g3701) & (!g3702)));
	assign g5299 = (((!g1914) & (!g2233) & (!g2242) & (!g5298)) + ((!g1914) & (!g2233) & (g2242) & (g5298)) + ((!g1914) & (g2233) & (!g2242) & (g5298)) + ((!g1914) & (g2233) & (g2242) & (!g5298)));
	assign g5300 = (((!g830) & (!g3088) & (!g5297) & (!g5299)) + ((!g830) & (!g3088) & (!g5297) & (g5299)) + ((!g830) & (!g3088) & (g5297) & (!g5299)) + ((!g830) & (!g3088) & (g5297) & (g5299)) + ((!g830) & (g3088) & (!g5297) & (!g5299)) + ((!g830) & (g3088) & (!g5297) & (g5299)) + ((!g830) & (g3088) & (g5297) & (!g5299)) + ((!g830) & (g3088) & (g5297) & (g5299)) + ((g830) & (!g3088) & (!g5297) & (g5299)) + ((g830) & (!g3088) & (g5297) & (!g5299)) + ((g830) & (!g3088) & (g5297) & (g5299)) + ((g830) & (g3088) & (!g5297) & (!g5299)));
	assign g5301 = (((!g2014) & (!g2052) & (!g2643) & (g2676) & (!g5267)) + ((!g2014) & (!g2052) & (!g2643) & (g2676) & (g5267)) + ((!g2014) & (!g2052) & (g2643) & (!g2676) & (g5267)) + ((!g2014) & (!g2052) & (g2643) & (g2676) & (!g5267)) + ((!g2014) & (g2052) & (!g2643) & (!g2676) & (!g5267)) + ((!g2014) & (g2052) & (!g2643) & (!g2676) & (g5267)) + ((!g2014) & (g2052) & (g2643) & (!g2676) & (!g5267)) + ((!g2014) & (g2052) & (g2643) & (g2676) & (g5267)) + ((g2014) & (!g2052) & (!g2643) & (!g2676) & (g5267)) + ((g2014) & (!g2052) & (!g2643) & (g2676) & (!g5267)) + ((g2014) & (!g2052) & (g2643) & (!g2676) & (!g5267)) + ((g2014) & (!g2052) & (g2643) & (!g2676) & (g5267)) + ((g2014) & (g2052) & (!g2643) & (!g2676) & (!g5267)) + ((g2014) & (g2052) & (!g2643) & (g2676) & (g5267)) + ((g2014) & (g2052) & (g2643) & (g2676) & (!g5267)) + ((g2014) & (g2052) & (g2643) & (g2676) & (g5267)));
	assign g5302 = (((!g2626) & (!g2629) & (!g2667) & (g2659) & (!g5269)) + ((!g2626) & (!g2629) & (!g2667) & (g2659) & (g5269)) + ((!g2626) & (!g2629) & (g2667) & (!g2659) & (!g5269)) + ((!g2626) & (!g2629) & (g2667) & (!g2659) & (g5269)) + ((!g2626) & (g2629) & (!g2667) & (!g2659) & (g5269)) + ((!g2626) & (g2629) & (!g2667) & (g2659) & (!g5269)) + ((!g2626) & (g2629) & (g2667) & (!g2659) & (!g5269)) + ((!g2626) & (g2629) & (g2667) & (g2659) & (g5269)) + ((g2626) & (!g2629) & (!g2667) & (!g2659) & (g5269)) + ((g2626) & (!g2629) & (!g2667) & (g2659) & (!g5269)) + ((g2626) & (!g2629) & (g2667) & (!g2659) & (!g5269)) + ((g2626) & (!g2629) & (g2667) & (g2659) & (g5269)) + ((g2626) & (g2629) & (!g2667) & (!g2659) & (!g5269)) + ((g2626) & (g2629) & (!g2667) & (!g2659) & (g5269)) + ((g2626) & (g2629) & (g2667) & (g2659) & (!g5269)) + ((g2626) & (g2629) & (g2667) & (g2659) & (g5269)));
	assign g5303 = (((!g830) & (!g1914) & (!g3090) & (!g5301) & (!g5302) & (key[216])) + ((!g830) & (!g1914) & (!g3090) & (!g5301) & (g5302) & (key[216])) + ((!g830) & (!g1914) & (!g3090) & (g5301) & (!g5302) & (key[216])) + ((!g830) & (!g1914) & (!g3090) & (g5301) & (g5302) & (key[216])) + ((!g830) & (!g1914) & (g3090) & (!g5301) & (!g5302) & (key[216])) + ((!g830) & (!g1914) & (g3090) & (!g5301) & (g5302) & (key[216])) + ((!g830) & (!g1914) & (g3090) & (g5301) & (!g5302) & (key[216])) + ((!g830) & (!g1914) & (g3090) & (g5301) & (g5302) & (key[216])) + ((!g830) & (g1914) & (!g3090) & (!g5301) & (!g5302) & (key[216])) + ((!g830) & (g1914) & (!g3090) & (!g5301) & (g5302) & (key[216])) + ((!g830) & (g1914) & (!g3090) & (g5301) & (!g5302) & (key[216])) + ((!g830) & (g1914) & (!g3090) & (g5301) & (g5302) & (key[216])) + ((!g830) & (g1914) & (g3090) & (!g5301) & (!g5302) & (key[216])) + ((!g830) & (g1914) & (g3090) & (!g5301) & (g5302) & (key[216])) + ((!g830) & (g1914) & (g3090) & (g5301) & (!g5302) & (key[216])) + ((!g830) & (g1914) & (g3090) & (g5301) & (g5302) & (key[216])) + ((g830) & (!g1914) & (!g3090) & (!g5301) & (g5302) & (!key[216])) + ((g830) & (!g1914) & (!g3090) & (!g5301) & (g5302) & (key[216])) + ((g830) & (!g1914) & (!g3090) & (g5301) & (g5302) & (!key[216])) + ((g830) & (!g1914) & (!g3090) & (g5301) & (g5302) & (key[216])) + ((g830) & (!g1914) & (g3090) & (!g5301) & (!g5302) & (!key[216])) + ((g830) & (!g1914) & (g3090) & (!g5301) & (!g5302) & (key[216])) + ((g830) & (!g1914) & (g3090) & (g5301) & (!g5302) & (!key[216])) + ((g830) & (!g1914) & (g3090) & (g5301) & (!g5302) & (key[216])) + ((g830) & (g1914) & (!g3090) & (g5301) & (!g5302) & (!key[216])) + ((g830) & (g1914) & (!g3090) & (g5301) & (!g5302) & (key[216])) + ((g830) & (g1914) & (!g3090) & (g5301) & (g5302) & (!key[216])) + ((g830) & (g1914) & (!g3090) & (g5301) & (g5302) & (key[216])) + ((g830) & (g1914) & (g3090) & (!g5301) & (!g5302) & (!key[216])) + ((g830) & (g1914) & (g3090) & (!g5301) & (!g5302) & (key[216])) + ((g830) & (g1914) & (g3090) & (!g5301) & (g5302) & (!key[216])) + ((g830) & (g1914) & (g3090) & (!g5301) & (g5302) & (key[216])));
	assign g5304 = (((!g3801) & (!g3802)));
	assign g5305 = (((!g1968) & (!g2486) & (!g5304)) + ((!g1968) & (g2486) & (g5304)) + ((g1968) & (!g2486) & (g5304)) + ((g1968) & (g2486) & (!g5304)));
	assign g5306 = (((!g830) & (!g3093) & (!g6028) & (key[152])) + ((!g830) & (!g3093) & (g6028) & (key[152])) + ((!g830) & (g3093) & (!g6028) & (key[152])) + ((!g830) & (g3093) & (g6028) & (key[152])) + ((g830) & (!g3093) & (g6028) & (!key[152])) + ((g830) & (!g3093) & (g6028) & (key[152])) + ((g830) & (g3093) & (!g6028) & (!key[152])) + ((g830) & (g3093) & (!g6028) & (key[152])));
	assign g5307 = (((!g2617) & (!g2665) & (!g2629) & (g2667) & (!g5258)) + ((!g2617) & (!g2665) & (!g2629) & (g2667) & (g5258)) + ((!g2617) & (!g2665) & (g2629) & (!g2667) & (g5258)) + ((!g2617) & (!g2665) & (g2629) & (g2667) & (!g5258)) + ((!g2617) & (g2665) & (!g2629) & (!g2667) & (!g5258)) + ((!g2617) & (g2665) & (!g2629) & (!g2667) & (g5258)) + ((!g2617) & (g2665) & (g2629) & (!g2667) & (!g5258)) + ((!g2617) & (g2665) & (g2629) & (g2667) & (g5258)) + ((g2617) & (!g2665) & (!g2629) & (!g2667) & (g5258)) + ((g2617) & (!g2665) & (!g2629) & (g2667) & (!g5258)) + ((g2617) & (!g2665) & (g2629) & (!g2667) & (!g5258)) + ((g2617) & (!g2665) & (g2629) & (!g2667) & (g5258)) + ((g2617) & (g2665) & (!g2629) & (!g2667) & (!g5258)) + ((g2617) & (g2665) & (!g2629) & (g2667) & (g5258)) + ((g2617) & (g2665) & (g2629) & (g2667) & (!g5258)) + ((g2617) & (g2665) & (g2629) & (g2667) & (g5258)));
	assign g5308 = (((!g1976) & (!g2048) & (!g2643) & (g2676) & (!g5260)) + ((!g1976) & (!g2048) & (!g2643) & (g2676) & (g5260)) + ((!g1976) & (!g2048) & (g2643) & (!g2676) & (g5260)) + ((!g1976) & (!g2048) & (g2643) & (g2676) & (!g5260)) + ((!g1976) & (g2048) & (!g2643) & (!g2676) & (!g5260)) + ((!g1976) & (g2048) & (!g2643) & (!g2676) & (g5260)) + ((!g1976) & (g2048) & (g2643) & (!g2676) & (!g5260)) + ((!g1976) & (g2048) & (g2643) & (g2676) & (g5260)) + ((g1976) & (!g2048) & (!g2643) & (!g2676) & (g5260)) + ((g1976) & (!g2048) & (!g2643) & (g2676) & (!g5260)) + ((g1976) & (!g2048) & (g2643) & (!g2676) & (!g5260)) + ((g1976) & (!g2048) & (g2643) & (!g2676) & (g5260)) + ((g1976) & (g2048) & (!g2643) & (!g2676) & (!g5260)) + ((g1976) & (g2048) & (!g2643) & (g2676) & (g5260)) + ((g1976) & (g2048) & (g2643) & (g2676) & (!g5260)) + ((g1976) & (g2048) & (g2643) & (g2676) & (g5260)));
	assign g5309 = (((!g830) & (!g1914) & (!g3095) & (!g5307) & (!g5308) & (nonce[56])) + ((!g830) & (!g1914) & (!g3095) & (!g5307) & (g5308) & (nonce[56])) + ((!g830) & (!g1914) & (!g3095) & (g5307) & (!g5308) & (nonce[56])) + ((!g830) & (!g1914) & (!g3095) & (g5307) & (g5308) & (nonce[56])) + ((!g830) & (!g1914) & (g3095) & (!g5307) & (!g5308) & (nonce[56])) + ((!g830) & (!g1914) & (g3095) & (!g5307) & (g5308) & (nonce[56])) + ((!g830) & (!g1914) & (g3095) & (g5307) & (!g5308) & (nonce[56])) + ((!g830) & (!g1914) & (g3095) & (g5307) & (g5308) & (nonce[56])) + ((!g830) & (g1914) & (!g3095) & (!g5307) & (!g5308) & (nonce[56])) + ((!g830) & (g1914) & (!g3095) & (!g5307) & (g5308) & (nonce[56])) + ((!g830) & (g1914) & (!g3095) & (g5307) & (!g5308) & (nonce[56])) + ((!g830) & (g1914) & (!g3095) & (g5307) & (g5308) & (nonce[56])) + ((!g830) & (g1914) & (g3095) & (!g5307) & (!g5308) & (nonce[56])) + ((!g830) & (g1914) & (g3095) & (!g5307) & (g5308) & (nonce[56])) + ((!g830) & (g1914) & (g3095) & (g5307) & (!g5308) & (nonce[56])) + ((!g830) & (g1914) & (g3095) & (g5307) & (g5308) & (nonce[56])) + ((g830) & (!g1914) & (!g3095) & (!g5307) & (g5308) & (!nonce[56])) + ((g830) & (!g1914) & (!g3095) & (!g5307) & (g5308) & (nonce[56])) + ((g830) & (!g1914) & (!g3095) & (g5307) & (g5308) & (!nonce[56])) + ((g830) & (!g1914) & (!g3095) & (g5307) & (g5308) & (nonce[56])) + ((g830) & (!g1914) & (g3095) & (!g5307) & (!g5308) & (!nonce[56])) + ((g830) & (!g1914) & (g3095) & (!g5307) & (!g5308) & (nonce[56])) + ((g830) & (!g1914) & (g3095) & (g5307) & (!g5308) & (!nonce[56])) + ((g830) & (!g1914) & (g3095) & (g5307) & (!g5308) & (nonce[56])) + ((g830) & (g1914) & (!g3095) & (g5307) & (!g5308) & (!nonce[56])) + ((g830) & (g1914) & (!g3095) & (g5307) & (!g5308) & (nonce[56])) + ((g830) & (g1914) & (!g3095) & (g5307) & (g5308) & (!nonce[56])) + ((g830) & (g1914) & (!g3095) & (g5307) & (g5308) & (nonce[56])) + ((g830) & (g1914) & (g3095) & (!g5307) & (!g5308) & (!nonce[56])) + ((g830) & (g1914) & (g3095) & (!g5307) & (!g5308) & (nonce[56])) + ((g830) & (g1914) & (g3095) & (!g5307) & (g5308) & (!nonce[56])) + ((g830) & (g1914) & (g3095) & (!g5307) & (g5308) & (nonce[56])));
	assign g5310 = (((!g3848) & (!g3849)));
	assign g5311 = (((g1914) & (!g2230) & (!g2242) & (!g5310)) + ((g1914) & (!g2230) & (g2242) & (g5310)) + ((g1914) & (g2230) & (!g2242) & (g5310)) + ((g1914) & (g2230) & (g2242) & (!g5310)));
	assign g5312 = (((!g3858) & (!g3859)));
	assign g5313 = (((!g1914) & (!g2247) & (!g2250) & (!g5312)) + ((!g1914) & (!g2247) & (g2250) & (g5312)) + ((!g1914) & (g2247) & (!g2250) & (g5312)) + ((!g1914) & (g2247) & (g2250) & (!g5312)));
	assign g5314 = (((!g830) & (!g3097) & (!g5311) & (!g5313)) + ((!g830) & (!g3097) & (!g5311) & (g5313)) + ((!g830) & (!g3097) & (g5311) & (!g5313)) + ((!g830) & (!g3097) & (g5311) & (g5313)) + ((!g830) & (g3097) & (!g5311) & (!g5313)) + ((!g830) & (g3097) & (!g5311) & (g5313)) + ((!g830) & (g3097) & (g5311) & (!g5313)) + ((!g830) & (g3097) & (g5311) & (g5313)) + ((g830) & (!g3097) & (!g5311) & (g5313)) + ((g830) & (!g3097) & (g5311) & (!g5313)) + ((g830) & (!g3097) & (g5311) & (g5313)) + ((g830) & (g3097) & (!g5311) & (!g5313)));
	assign g5315 = (((!g2178) & (!g1439) & (!g3632)) + ((!g2178) & (g1439) & (g3632)) + ((g2178) & (!g1439) & (g3632)) + ((g2178) & (g1439) & (!g3632)));
	assign g5316 = (((!g2456) & (!g2535) & (!g2503) & (g2539) & (!g5289)) + ((!g2456) & (!g2535) & (!g2503) & (g2539) & (g5289)) + ((!g2456) & (!g2535) & (g2503) & (!g2539) & (!g5289)) + ((!g2456) & (!g2535) & (g2503) & (g2539) & (g5289)) + ((!g2456) & (g2535) & (!g2503) & (!g2539) & (!g5289)) + ((!g2456) & (g2535) & (!g2503) & (!g2539) & (g5289)) + ((!g2456) & (g2535) & (g2503) & (!g2539) & (g5289)) + ((!g2456) & (g2535) & (g2503) & (g2539) & (!g5289)) + ((g2456) & (!g2535) & (!g2503) & (!g2539) & (!g5289)) + ((g2456) & (!g2535) & (!g2503) & (g2539) & (g5289)) + ((g2456) & (!g2535) & (g2503) & (!g2539) & (!g5289)) + ((g2456) & (!g2535) & (g2503) & (!g2539) & (g5289)) + ((g2456) & (g2535) & (!g2503) & (!g2539) & (g5289)) + ((g2456) & (g2535) & (!g2503) & (g2539) & (!g5289)) + ((g2456) & (g2535) & (g2503) & (g2539) & (!g5289)) + ((g2456) & (g2535) & (g2503) & (g2539) & (g5289)));
	assign g5317 = (((!g830) & (!g1914) & (!g3106) & (!g5315) & (!g5316) & (key[25])) + ((!g830) & (!g1914) & (!g3106) & (!g5315) & (g5316) & (key[25])) + ((!g830) & (!g1914) & (!g3106) & (g5315) & (!g5316) & (key[25])) + ((!g830) & (!g1914) & (!g3106) & (g5315) & (g5316) & (key[25])) + ((!g830) & (!g1914) & (g3106) & (!g5315) & (!g5316) & (key[25])) + ((!g830) & (!g1914) & (g3106) & (!g5315) & (g5316) & (key[25])) + ((!g830) & (!g1914) & (g3106) & (g5315) & (!g5316) & (key[25])) + ((!g830) & (!g1914) & (g3106) & (g5315) & (g5316) & (key[25])) + ((!g830) & (g1914) & (!g3106) & (!g5315) & (!g5316) & (key[25])) + ((!g830) & (g1914) & (!g3106) & (!g5315) & (g5316) & (key[25])) + ((!g830) & (g1914) & (!g3106) & (g5315) & (!g5316) & (key[25])) + ((!g830) & (g1914) & (!g3106) & (g5315) & (g5316) & (key[25])) + ((!g830) & (g1914) & (g3106) & (!g5315) & (!g5316) & (key[25])) + ((!g830) & (g1914) & (g3106) & (!g5315) & (g5316) & (key[25])) + ((!g830) & (g1914) & (g3106) & (g5315) & (!g5316) & (key[25])) + ((!g830) & (g1914) & (g3106) & (g5315) & (g5316) & (key[25])) + ((g830) & (!g1914) & (!g3106) & (!g5315) & (g5316) & (!key[25])) + ((g830) & (!g1914) & (!g3106) & (!g5315) & (g5316) & (key[25])) + ((g830) & (!g1914) & (!g3106) & (g5315) & (g5316) & (!key[25])) + ((g830) & (!g1914) & (!g3106) & (g5315) & (g5316) & (key[25])) + ((g830) & (!g1914) & (g3106) & (!g5315) & (!g5316) & (!key[25])) + ((g830) & (!g1914) & (g3106) & (!g5315) & (!g5316) & (key[25])) + ((g830) & (!g1914) & (g3106) & (g5315) & (!g5316) & (!key[25])) + ((g830) & (!g1914) & (g3106) & (g5315) & (!g5316) & (key[25])) + ((g830) & (g1914) & (!g3106) & (g5315) & (!g5316) & (!key[25])) + ((g830) & (g1914) & (!g3106) & (g5315) & (!g5316) & (key[25])) + ((g830) & (g1914) & (!g3106) & (g5315) & (g5316) & (!key[25])) + ((g830) & (g1914) & (!g3106) & (g5315) & (g5316) & (key[25])) + ((g830) & (g1914) & (g3106) & (!g5315) & (!g5316) & (!key[25])) + ((g830) & (g1914) & (g3106) & (!g5315) & (!g5316) & (key[25])) + ((g830) & (g1914) & (g3106) & (!g5315) & (g5316) & (!key[25])) + ((g830) & (g1914) & (g3106) & (!g5315) & (g5316) & (key[25])));
	assign g5318 = (((!g1991) & (!g1993) & (!g5278) & (!g2236) & (g2273)) + ((!g1991) & (!g1993) & (!g5278) & (g2236) & (!g2273)) + ((!g1991) & (!g1993) & (g5278) & (!g2236) & (g2273)) + ((!g1991) & (!g1993) & (g5278) & (g2236) & (g2273)) + ((!g1991) & (g1993) & (!g5278) & (!g2236) & (!g2273)) + ((!g1991) & (g1993) & (!g5278) & (g2236) & (g2273)) + ((!g1991) & (g1993) & (g5278) & (!g2236) & (!g2273)) + ((!g1991) & (g1993) & (g5278) & (g2236) & (!g2273)) + ((g1991) & (!g1993) & (!g5278) & (!g2236) & (!g2273)) + ((g1991) & (!g1993) & (!g5278) & (g2236) & (!g2273)) + ((g1991) & (!g1993) & (g5278) & (!g2236) & (g2273)) + ((g1991) & (!g1993) & (g5278) & (g2236) & (!g2273)) + ((g1991) & (g1993) & (!g5278) & (!g2236) & (g2273)) + ((g1991) & (g1993) & (!g5278) & (g2236) & (g2273)) + ((g1991) & (g1993) & (g5278) & (!g2236) & (!g2273)) + ((g1991) & (g1993) & (g5278) & (g2236) & (g2273)));
	assign g5319 = (((!g1953) & (!g1955) & (!g2227) & (g2279) & (!g5280)) + ((!g1953) & (!g1955) & (!g2227) & (g2279) & (g5280)) + ((!g1953) & (!g1955) & (g2227) & (!g2279) & (!g5280)) + ((!g1953) & (!g1955) & (g2227) & (g2279) & (g5280)) + ((!g1953) & (g1955) & (!g2227) & (!g2279) & (!g5280)) + ((!g1953) & (g1955) & (!g2227) & (!g2279) & (g5280)) + ((!g1953) & (g1955) & (g2227) & (!g2279) & (g5280)) + ((!g1953) & (g1955) & (g2227) & (g2279) & (!g5280)) + ((g1953) & (!g1955) & (!g2227) & (!g2279) & (!g5280)) + ((g1953) & (!g1955) & (!g2227) & (g2279) & (g5280)) + ((g1953) & (!g1955) & (g2227) & (!g2279) & (!g5280)) + ((g1953) & (!g1955) & (g2227) & (!g2279) & (g5280)) + ((g1953) & (g1955) & (!g2227) & (!g2279) & (g5280)) + ((g1953) & (g1955) & (!g2227) & (g2279) & (!g5280)) + ((g1953) & (g1955) & (g2227) & (g2279) & (!g5280)) + ((g1953) & (g1955) & (g2227) & (g2279) & (g5280)));
	assign g5320 = (((g830) & (!g1914) & (!g3113) & (!g5318) & (g5319)) + ((g830) & (!g1914) & (!g3113) & (g5318) & (g5319)) + ((g830) & (!g1914) & (g3113) & (!g5318) & (!g5319)) + ((g830) & (!g1914) & (g3113) & (g5318) & (!g5319)) + ((g830) & (g1914) & (!g3113) & (g5318) & (!g5319)) + ((g830) & (g1914) & (!g3113) & (g5318) & (g5319)) + ((g830) & (g1914) & (g3113) & (!g5318) & (!g5319)) + ((g830) & (g1914) & (g3113) & (!g5318) & (g5319)));
	assign g5321 = (((!g2003) & (!g2005) & (!g2462) & (g2542) & (!g5292)) + ((!g2003) & (!g2005) & (!g2462) & (g2542) & (g5292)) + ((!g2003) & (!g2005) & (g2462) & (!g2542) & (!g5292)) + ((!g2003) & (!g2005) & (g2462) & (g2542) & (g5292)) + ((!g2003) & (g2005) & (!g2462) & (!g2542) & (!g5292)) + ((!g2003) & (g2005) & (!g2462) & (!g2542) & (g5292)) + ((!g2003) & (g2005) & (g2462) & (!g2542) & (g5292)) + ((!g2003) & (g2005) & (g2462) & (g2542) & (!g5292)) + ((g2003) & (!g2005) & (!g2462) & (!g2542) & (!g5292)) + ((g2003) & (!g2005) & (!g2462) & (g2542) & (g5292)) + ((g2003) & (!g2005) & (g2462) & (!g2542) & (!g5292)) + ((g2003) & (!g2005) & (g2462) & (!g2542) & (g5292)) + ((g2003) & (g2005) & (!g2462) & (!g2542) & (g5292)) + ((g2003) & (g2005) & (!g2462) & (g2542) & (!g5292)) + ((g2003) & (g2005) & (g2462) & (g2542) & (!g5292)) + ((g2003) & (g2005) & (g2462) & (g2542) & (g5292)));
	assign g5322 = (((!g1914) & (!g2813) & (!g2819) & (!g3680) & (!g5321)) + ((!g1914) & (!g2813) & (!g2819) & (!g3680) & (g5321)) + ((!g1914) & (!g2813) & (g2819) & (g3680) & (!g5321)) + ((!g1914) & (!g2813) & (g2819) & (g3680) & (g5321)) + ((!g1914) & (g2813) & (!g2819) & (g3680) & (!g5321)) + ((!g1914) & (g2813) & (!g2819) & (g3680) & (g5321)) + ((!g1914) & (g2813) & (g2819) & (!g3680) & (!g5321)) + ((!g1914) & (g2813) & (g2819) & (!g3680) & (g5321)) + ((g1914) & (!g2813) & (!g2819) & (!g3680) & (g5321)) + ((g1914) & (!g2813) & (!g2819) & (g3680) & (g5321)) + ((g1914) & (!g2813) & (g2819) & (!g3680) & (g5321)) + ((g1914) & (!g2813) & (g2819) & (g3680) & (g5321)) + ((g1914) & (g2813) & (!g2819) & (!g3680) & (g5321)) + ((g1914) & (g2813) & (!g2819) & (g3680) & (g5321)) + ((g1914) & (g2813) & (g2819) & (!g3680) & (g5321)) + ((g1914) & (g2813) & (g2819) & (g3680) & (g5321)));
	assign g8333 = (((!g5560) & (g5639) & (!g5323)) + ((!g5560) & (g5639) & (g5323)) + ((g5560) & (!g5639) & (g5323)) + ((g5560) & (g5639) & (g5323)));
	assign g5324 = (((!g830) & (!g3116) & (!g5322) & (g5323)) + ((!g830) & (!g3116) & (g5322) & (g5323)) + ((!g830) & (g3116) & (!g5322) & (g5323)) + ((!g830) & (g3116) & (g5322) & (g5323)) + ((g830) & (!g3116) & (g5322) & (!g5323)) + ((g830) & (!g3116) & (g5322) & (g5323)) + ((g830) & (g3116) & (!g5322) & (!g5323)) + ((g830) & (g3116) & (!g5322) & (g5323)));
	assign g5325 = (((!g2804) & (!g2816) & (!g3789)) + ((!g2804) & (g2816) & (g3789)) + ((g2804) & (!g2816) & (g3789)) + ((g2804) & (g2816) & (!g3789)));
	assign g5326 = (((!g1968) & (!g1970) & (!g2486) & (g2544) & (!g5304)) + ((!g1968) & (!g1970) & (!g2486) & (g2544) & (g5304)) + ((!g1968) & (!g1970) & (g2486) & (!g2544) & (!g5304)) + ((!g1968) & (!g1970) & (g2486) & (g2544) & (g5304)) + ((!g1968) & (g1970) & (!g2486) & (!g2544) & (!g5304)) + ((!g1968) & (g1970) & (!g2486) & (!g2544) & (g5304)) + ((!g1968) & (g1970) & (g2486) & (!g2544) & (g5304)) + ((!g1968) & (g1970) & (g2486) & (g2544) & (!g5304)) + ((g1968) & (!g1970) & (!g2486) & (!g2544) & (!g5304)) + ((g1968) & (!g1970) & (!g2486) & (g2544) & (g5304)) + ((g1968) & (!g1970) & (g2486) & (!g2544) & (!g5304)) + ((g1968) & (!g1970) & (g2486) & (!g2544) & (g5304)) + ((g1968) & (g1970) & (!g2486) & (!g2544) & (g5304)) + ((g1968) & (g1970) & (!g2486) & (g2544) & (!g5304)) + ((g1968) & (g1970) & (g2486) & (g2544) & (!g5304)) + ((g1968) & (g1970) & (g2486) & (g2544) & (g5304)));
	assign g5327 = (((!g830) & (!g1914) & (!g3119) & (!g5325) & (!g5326) & (key[153])) + ((!g830) & (!g1914) & (!g3119) & (!g5325) & (g5326) & (key[153])) + ((!g830) & (!g1914) & (!g3119) & (g5325) & (!g5326) & (key[153])) + ((!g830) & (!g1914) & (!g3119) & (g5325) & (g5326) & (key[153])) + ((!g830) & (!g1914) & (g3119) & (!g5325) & (!g5326) & (key[153])) + ((!g830) & (!g1914) & (g3119) & (!g5325) & (g5326) & (key[153])) + ((!g830) & (!g1914) & (g3119) & (g5325) & (!g5326) & (key[153])) + ((!g830) & (!g1914) & (g3119) & (g5325) & (g5326) & (key[153])) + ((!g830) & (g1914) & (!g3119) & (!g5325) & (!g5326) & (key[153])) + ((!g830) & (g1914) & (!g3119) & (!g5325) & (g5326) & (key[153])) + ((!g830) & (g1914) & (!g3119) & (g5325) & (!g5326) & (key[153])) + ((!g830) & (g1914) & (!g3119) & (g5325) & (g5326) & (key[153])) + ((!g830) & (g1914) & (g3119) & (!g5325) & (!g5326) & (key[153])) + ((!g830) & (g1914) & (g3119) & (!g5325) & (g5326) & (key[153])) + ((!g830) & (g1914) & (g3119) & (g5325) & (!g5326) & (key[153])) + ((!g830) & (g1914) & (g3119) & (g5325) & (g5326) & (key[153])) + ((g830) & (!g1914) & (!g3119) & (!g5325) & (g5326) & (!key[153])) + ((g830) & (!g1914) & (!g3119) & (!g5325) & (g5326) & (key[153])) + ((g830) & (!g1914) & (!g3119) & (g5325) & (g5326) & (!key[153])) + ((g830) & (!g1914) & (!g3119) & (g5325) & (g5326) & (key[153])) + ((g830) & (!g1914) & (g3119) & (!g5325) & (!g5326) & (!key[153])) + ((g830) & (!g1914) & (g3119) & (!g5325) & (!g5326) & (key[153])) + ((g830) & (!g1914) & (g3119) & (g5325) & (!g5326) & (!key[153])) + ((g830) & (!g1914) & (g3119) & (g5325) & (!g5326) & (key[153])) + ((g830) & (g1914) & (!g3119) & (g5325) & (!g5326) & (!key[153])) + ((g830) & (g1914) & (!g3119) & (g5325) & (!g5326) & (key[153])) + ((g830) & (g1914) & (!g3119) & (g5325) & (g5326) & (!key[153])) + ((g830) & (g1914) & (!g3119) & (g5325) & (g5326) & (key[153])) + ((g830) & (g1914) & (g3119) & (!g5325) & (!g5326) & (!key[153])) + ((g830) & (g1914) & (g3119) & (!g5325) & (!g5326) & (key[153])) + ((g830) & (g1914) & (g3119) & (!g5325) & (g5326) & (!key[153])) + ((g830) & (g1914) & (g3119) & (!g5325) & (g5326) & (key[153])));
	assign g5328 = (((!g5275) & (!g2474) & (!g2486) & (!g2529) & (g2544)) + ((!g5275) & (!g2474) & (!g2486) & (g2529) & (!g2544)) + ((!g5275) & (!g2474) & (g2486) & (!g2529) & (!g2544)) + ((!g5275) & (!g2474) & (g2486) & (g2529) & (g2544)) + ((!g5275) & (g2474) & (!g2486) & (!g2529) & (!g2544)) + ((!g5275) & (g2474) & (!g2486) & (g2529) & (g2544)) + ((!g5275) & (g2474) & (g2486) & (!g2529) & (!g2544)) + ((!g5275) & (g2474) & (g2486) & (g2529) & (g2544)) + ((g5275) & (!g2474) & (!g2486) & (!g2529) & (g2544)) + ((g5275) & (!g2474) & (!g2486) & (g2529) & (!g2544)) + ((g5275) & (!g2474) & (g2486) & (!g2529) & (g2544)) + ((g5275) & (!g2474) & (g2486) & (g2529) & (!g2544)) + ((g5275) & (g2474) & (!g2486) & (!g2529) & (g2544)) + ((g5275) & (g2474) & (!g2486) & (g2529) & (!g2544)) + ((g5275) & (g2474) & (g2486) & (!g2529) & (!g2544)) + ((g5275) & (g2474) & (g2486) & (g2529) & (g2544)));
	assign g5329 = (((!g2181) & (!g1439) & (!g3455)) + ((!g2181) & (g1439) & (g3455)) + ((g2181) & (!g1439) & (g3455)) + ((g2181) & (g1439) & (!g3455)));
	assign g5330 = (((!g830) & (!g1914) & (!g3122) & (!g5328) & (!g5329) & (key[121])) + ((!g830) & (!g1914) & (!g3122) & (!g5328) & (g5329) & (key[121])) + ((!g830) & (!g1914) & (!g3122) & (g5328) & (!g5329) & (key[121])) + ((!g830) & (!g1914) & (!g3122) & (g5328) & (g5329) & (key[121])) + ((!g830) & (!g1914) & (g3122) & (!g5328) & (!g5329) & (key[121])) + ((!g830) & (!g1914) & (g3122) & (!g5328) & (g5329) & (key[121])) + ((!g830) & (!g1914) & (g3122) & (g5328) & (!g5329) & (key[121])) + ((!g830) & (!g1914) & (g3122) & (g5328) & (g5329) & (key[121])) + ((!g830) & (g1914) & (!g3122) & (!g5328) & (!g5329) & (key[121])) + ((!g830) & (g1914) & (!g3122) & (!g5328) & (g5329) & (key[121])) + ((!g830) & (g1914) & (!g3122) & (g5328) & (!g5329) & (key[121])) + ((!g830) & (g1914) & (!g3122) & (g5328) & (g5329) & (key[121])) + ((!g830) & (g1914) & (g3122) & (!g5328) & (!g5329) & (key[121])) + ((!g830) & (g1914) & (g3122) & (!g5328) & (g5329) & (key[121])) + ((!g830) & (g1914) & (g3122) & (g5328) & (!g5329) & (key[121])) + ((!g830) & (g1914) & (g3122) & (g5328) & (g5329) & (key[121])) + ((g830) & (!g1914) & (!g3122) & (!g5328) & (g5329) & (!key[121])) + ((g830) & (!g1914) & (!g3122) & (!g5328) & (g5329) & (key[121])) + ((g830) & (!g1914) & (!g3122) & (g5328) & (g5329) & (!key[121])) + ((g830) & (!g1914) & (!g3122) & (g5328) & (g5329) & (key[121])) + ((g830) & (!g1914) & (g3122) & (!g5328) & (!g5329) & (!key[121])) + ((g830) & (!g1914) & (g3122) & (!g5328) & (!g5329) & (key[121])) + ((g830) & (!g1914) & (g3122) & (g5328) & (!g5329) & (!key[121])) + ((g830) & (!g1914) & (g3122) & (g5328) & (!g5329) & (key[121])) + ((g830) & (g1914) & (!g3122) & (g5328) & (!g5329) & (!key[121])) + ((g830) & (g1914) & (!g3122) & (g5328) & (!g5329) & (key[121])) + ((g830) & (g1914) & (!g3122) & (g5328) & (g5329) & (!key[121])) + ((g830) & (g1914) & (!g3122) & (g5328) & (g5329) & (key[121])) + ((g830) & (g1914) & (g3122) & (!g5328) & (!g5329) & (!key[121])) + ((g830) & (g1914) & (g3122) & (!g5328) & (!g5329) & (key[121])) + ((g830) & (g1914) & (g3122) & (!g5328) & (g5329) & (!key[121])) + ((g830) & (g1914) & (g3122) & (!g5328) & (g5329) & (key[121])));
	assign g5331 = (((!g2797) & (!g3566) & (!g2819)) + ((!g2797) & (g3566) & (g2819)) + ((g2797) & (!g3566) & (g2819)) + ((g2797) & (g3566) & (!g2819)));
	assign g5332 = (((!g1967) & (!g1969) & (!g2497) & (g2531) & (!g5283)) + ((!g1967) & (!g1969) & (!g2497) & (g2531) & (g5283)) + ((!g1967) & (!g1969) & (g2497) & (!g2531) & (!g5283)) + ((!g1967) & (!g1969) & (g2497) & (g2531) & (g5283)) + ((!g1967) & (g1969) & (!g2497) & (!g2531) & (!g5283)) + ((!g1967) & (g1969) & (!g2497) & (!g2531) & (g5283)) + ((!g1967) & (g1969) & (g2497) & (!g2531) & (g5283)) + ((!g1967) & (g1969) & (g2497) & (g2531) & (!g5283)) + ((g1967) & (!g1969) & (!g2497) & (!g2531) & (!g5283)) + ((g1967) & (!g1969) & (!g2497) & (g2531) & (g5283)) + ((g1967) & (!g1969) & (g2497) & (!g2531) & (!g5283)) + ((g1967) & (!g1969) & (g2497) & (!g2531) & (g5283)) + ((g1967) & (g1969) & (!g2497) & (!g2531) & (g5283)) + ((g1967) & (g1969) & (!g2497) & (g2531) & (!g5283)) + ((g1967) & (g1969) & (g2497) & (g2531) & (!g5283)) + ((g1967) & (g1969) & (g2497) & (g2531) & (g5283)));
	assign g5333 = (((!g830) & (!g1914) & (!g3125) & (!g5331) & (!g5332) & (nonce[25])) + ((!g830) & (!g1914) & (!g3125) & (!g5331) & (g5332) & (nonce[25])) + ((!g830) & (!g1914) & (!g3125) & (g5331) & (!g5332) & (nonce[25])) + ((!g830) & (!g1914) & (!g3125) & (g5331) & (g5332) & (nonce[25])) + ((!g830) & (!g1914) & (g3125) & (!g5331) & (!g5332) & (nonce[25])) + ((!g830) & (!g1914) & (g3125) & (!g5331) & (g5332) & (nonce[25])) + ((!g830) & (!g1914) & (g3125) & (g5331) & (!g5332) & (nonce[25])) + ((!g830) & (!g1914) & (g3125) & (g5331) & (g5332) & (nonce[25])) + ((!g830) & (g1914) & (!g3125) & (!g5331) & (!g5332) & (nonce[25])) + ((!g830) & (g1914) & (!g3125) & (!g5331) & (g5332) & (nonce[25])) + ((!g830) & (g1914) & (!g3125) & (g5331) & (!g5332) & (nonce[25])) + ((!g830) & (g1914) & (!g3125) & (g5331) & (g5332) & (nonce[25])) + ((!g830) & (g1914) & (g3125) & (!g5331) & (!g5332) & (nonce[25])) + ((!g830) & (g1914) & (g3125) & (!g5331) & (g5332) & (nonce[25])) + ((!g830) & (g1914) & (g3125) & (g5331) & (!g5332) & (nonce[25])) + ((!g830) & (g1914) & (g3125) & (g5331) & (g5332) & (nonce[25])) + ((g830) & (!g1914) & (!g3125) & (!g5331) & (g5332) & (!nonce[25])) + ((g830) & (!g1914) & (!g3125) & (!g5331) & (g5332) & (nonce[25])) + ((g830) & (!g1914) & (!g3125) & (g5331) & (g5332) & (!nonce[25])) + ((g830) & (!g1914) & (!g3125) & (g5331) & (g5332) & (nonce[25])) + ((g830) & (!g1914) & (g3125) & (!g5331) & (!g5332) & (!nonce[25])) + ((g830) & (!g1914) & (g3125) & (!g5331) & (!g5332) & (nonce[25])) + ((g830) & (!g1914) & (g3125) & (g5331) & (!g5332) & (!nonce[25])) + ((g830) & (!g1914) & (g3125) & (g5331) & (!g5332) & (nonce[25])) + ((g830) & (g1914) & (!g3125) & (g5331) & (!g5332) & (!nonce[25])) + ((g830) & (g1914) & (!g3125) & (g5331) & (!g5332) & (nonce[25])) + ((g830) & (g1914) & (!g3125) & (g5331) & (g5332) & (!nonce[25])) + ((g830) & (g1914) & (!g3125) & (g5331) & (g5332) & (nonce[25])) + ((g830) & (g1914) & (g3125) & (!g5331) & (!g5332) & (!nonce[25])) + ((g830) & (g1914) & (g3125) & (!g5331) & (!g5332) & (nonce[25])) + ((g830) & (g1914) & (g3125) & (!g5331) & (g5332) & (!nonce[25])) + ((g830) & (g1914) & (g3125) & (!g5331) & (g5332) & (nonce[25])));
	assign g5334 = (((!g2217) & (!g2277) & (!g2250) & (g2283) & (!g5296)) + ((!g2217) & (!g2277) & (!g2250) & (g2283) & (g5296)) + ((!g2217) & (!g2277) & (g2250) & (!g2283) & (!g5296)) + ((!g2217) & (!g2277) & (g2250) & (g2283) & (g5296)) + ((!g2217) & (g2277) & (!g2250) & (!g2283) & (!g5296)) + ((!g2217) & (g2277) & (!g2250) & (!g2283) & (g5296)) + ((!g2217) & (g2277) & (g2250) & (!g2283) & (g5296)) + ((!g2217) & (g2277) & (g2250) & (g2283) & (!g5296)) + ((g2217) & (!g2277) & (!g2250) & (!g2283) & (!g5296)) + ((g2217) & (!g2277) & (!g2250) & (g2283) & (g5296)) + ((g2217) & (!g2277) & (g2250) & (!g2283) & (!g5296)) + ((g2217) & (!g2277) & (g2250) & (!g2283) & (g5296)) + ((g2217) & (g2277) & (!g2250) & (!g2283) & (g5296)) + ((g2217) & (g2277) & (!g2250) & (g2283) & (!g5296)) + ((g2217) & (g2277) & (g2250) & (g2283) & (!g5296)) + ((g2217) & (g2277) & (g2250) & (g2283) & (g5296)));
	assign g5335 = (((!g2233) & (!g2267) & (!g2242) & (g2288) & (!g5298)) + ((!g2233) & (!g2267) & (!g2242) & (g2288) & (g5298)) + ((!g2233) & (!g2267) & (g2242) & (!g2288) & (!g5298)) + ((!g2233) & (!g2267) & (g2242) & (g2288) & (g5298)) + ((!g2233) & (g2267) & (!g2242) & (!g2288) & (!g5298)) + ((!g2233) & (g2267) & (!g2242) & (!g2288) & (g5298)) + ((!g2233) & (g2267) & (g2242) & (!g2288) & (g5298)) + ((!g2233) & (g2267) & (g2242) & (g2288) & (!g5298)) + ((g2233) & (!g2267) & (!g2242) & (!g2288) & (!g5298)) + ((g2233) & (!g2267) & (!g2242) & (g2288) & (g5298)) + ((g2233) & (!g2267) & (g2242) & (!g2288) & (!g5298)) + ((g2233) & (!g2267) & (g2242) & (!g2288) & (g5298)) + ((g2233) & (g2267) & (!g2242) & (!g2288) & (g5298)) + ((g2233) & (g2267) & (!g2242) & (g2288) & (!g5298)) + ((g2233) & (g2267) & (g2242) & (g2288) & (!g5298)) + ((g2233) & (g2267) & (g2242) & (g2288) & (g5298)));
	assign g5336 = (((!g830) & (!g1914) & (!g3128) & (!g5334) & (!g5335)) + ((!g830) & (!g1914) & (!g3128) & (!g5334) & (g5335)) + ((!g830) & (!g1914) & (!g3128) & (g5334) & (!g5335)) + ((!g830) & (!g1914) & (!g3128) & (g5334) & (g5335)) + ((!g830) & (!g1914) & (g3128) & (!g5334) & (!g5335)) + ((!g830) & (!g1914) & (g3128) & (!g5334) & (g5335)) + ((!g830) & (!g1914) & (g3128) & (g5334) & (!g5335)) + ((!g830) & (!g1914) & (g3128) & (g5334) & (g5335)) + ((!g830) & (g1914) & (!g3128) & (!g5334) & (!g5335)) + ((!g830) & (g1914) & (!g3128) & (!g5334) & (g5335)) + ((!g830) & (g1914) & (!g3128) & (g5334) & (!g5335)) + ((!g830) & (g1914) & (!g3128) & (g5334) & (g5335)) + ((!g830) & (g1914) & (g3128) & (!g5334) & (!g5335)) + ((!g830) & (g1914) & (g3128) & (!g5334) & (g5335)) + ((!g830) & (g1914) & (g3128) & (g5334) & (!g5335)) + ((!g830) & (g1914) & (g3128) & (g5334) & (g5335)) + ((g830) & (!g1914) & (!g3128) & (!g5334) & (g5335)) + ((g830) & (!g1914) & (!g3128) & (g5334) & (g5335)) + ((g830) & (!g1914) & (g3128) & (!g5334) & (!g5335)) + ((g830) & (!g1914) & (g3128) & (g5334) & (!g5335)) + ((g830) & (g1914) & (!g3128) & (g5334) & (!g5335)) + ((g830) & (g1914) & (!g3128) & (g5334) & (g5335)) + ((g830) & (g1914) & (g3128) & (!g5334) & (!g5335)) + ((g830) & (g1914) & (g3128) & (!g5334) & (g5335)));
	assign g5337 = (((!g3820) & (!g3821)));
	assign g5338 = (((g1914) & (!g2708) & (!g2728) & (!g5337)) + ((g1914) & (!g2708) & (g2728) & (g5337)) + ((g1914) & (g2708) & (!g2728) & (g5337)) + ((g1914) & (g2708) & (g2728) & (!g5337)));
	assign g5339 = (((!g3837) & (!g3838)));
	assign g5340 = (((!g1914) & (!g2099) & (!g2752) & (!g5339)) + ((!g1914) & (!g2099) & (g2752) & (g5339)) + ((!g1914) & (g2099) & (!g2752) & (g5339)) + ((!g1914) & (g2099) & (g2752) & (!g5339)));
	assign g5341 = (((!g830) & (!g3131) & (!g5338) & (!g5340) & (nonce[57])) + ((!g830) & (!g3131) & (!g5338) & (g5340) & (nonce[57])) + ((!g830) & (!g3131) & (g5338) & (!g5340) & (nonce[57])) + ((!g830) & (!g3131) & (g5338) & (g5340) & (nonce[57])) + ((!g830) & (g3131) & (!g5338) & (!g5340) & (nonce[57])) + ((!g830) & (g3131) & (!g5338) & (g5340) & (nonce[57])) + ((!g830) & (g3131) & (g5338) & (!g5340) & (nonce[57])) + ((!g830) & (g3131) & (g5338) & (g5340) & (nonce[57])) + ((g830) & (!g3131) & (!g5338) & (g5340) & (!nonce[57])) + ((g830) & (!g3131) & (!g5338) & (g5340) & (nonce[57])) + ((g830) & (!g3131) & (g5338) & (!g5340) & (!nonce[57])) + ((g830) & (!g3131) & (g5338) & (!g5340) & (nonce[57])) + ((g830) & (!g3131) & (g5338) & (g5340) & (!nonce[57])) + ((g830) & (!g3131) & (g5338) & (g5340) & (nonce[57])) + ((g830) & (g3131) & (!g5338) & (!g5340) & (!nonce[57])) + ((g830) & (g3131) & (!g5338) & (!g5340) & (nonce[57])));
	assign g5342 = (((!g2004) & (!g2006) & (!g5286) & (!g2503) & (g2539)) + ((!g2004) & (!g2006) & (!g5286) & (g2503) & (!g2539)) + ((!g2004) & (!g2006) & (g5286) & (!g2503) & (g2539)) + ((!g2004) & (!g2006) & (g5286) & (g2503) & (g2539)) + ((!g2004) & (g2006) & (!g5286) & (!g2503) & (!g2539)) + ((!g2004) & (g2006) & (!g5286) & (g2503) & (g2539)) + ((!g2004) & (g2006) & (g5286) & (!g2503) & (!g2539)) + ((!g2004) & (g2006) & (g5286) & (g2503) & (!g2539)) + ((g2004) & (!g2006) & (!g5286) & (!g2503) & (!g2539)) + ((g2004) & (!g2006) & (!g5286) & (g2503) & (!g2539)) + ((g2004) & (!g2006) & (g5286) & (!g2503) & (g2539)) + ((g2004) & (!g2006) & (g5286) & (g2503) & (!g2539)) + ((g2004) & (g2006) & (!g5286) & (!g2503) & (g2539)) + ((g2004) & (g2006) & (!g5286) & (g2503) & (g2539)) + ((g2004) & (g2006) & (g5286) & (!g2503) & (!g2539)) + ((g2004) & (g2006) & (g5286) & (g2503) & (g2539)));
	assign g5343 = (((!g2804) & (!g2807) & (!g3613)) + ((!g2804) & (g2807) & (g3613)) + ((g2804) & (!g2807) & (g3613)) + ((g2804) & (g2807) & (!g3613)));
	assign g5344 = (((!g830) & (!g1914) & (!g3136) & (!g5342) & (!g5343) & (key[249])) + ((!g830) & (!g1914) & (!g3136) & (!g5342) & (g5343) & (key[249])) + ((!g830) & (!g1914) & (!g3136) & (g5342) & (!g5343) & (key[249])) + ((!g830) & (!g1914) & (!g3136) & (g5342) & (g5343) & (key[249])) + ((!g830) & (!g1914) & (g3136) & (!g5342) & (!g5343) & (key[249])) + ((!g830) & (!g1914) & (g3136) & (!g5342) & (g5343) & (key[249])) + ((!g830) & (!g1914) & (g3136) & (g5342) & (!g5343) & (key[249])) + ((!g830) & (!g1914) & (g3136) & (g5342) & (g5343) & (key[249])) + ((!g830) & (g1914) & (!g3136) & (!g5342) & (!g5343) & (key[249])) + ((!g830) & (g1914) & (!g3136) & (!g5342) & (g5343) & (key[249])) + ((!g830) & (g1914) & (!g3136) & (g5342) & (!g5343) & (key[249])) + ((!g830) & (g1914) & (!g3136) & (g5342) & (g5343) & (key[249])) + ((!g830) & (g1914) & (g3136) & (!g5342) & (!g5343) & (key[249])) + ((!g830) & (g1914) & (g3136) & (!g5342) & (g5343) & (key[249])) + ((!g830) & (g1914) & (g3136) & (g5342) & (!g5343) & (key[249])) + ((!g830) & (g1914) & (g3136) & (g5342) & (g5343) & (key[249])) + ((g830) & (!g1914) & (!g3136) & (!g5342) & (g5343) & (!key[249])) + ((g830) & (!g1914) & (!g3136) & (!g5342) & (g5343) & (key[249])) + ((g830) & (!g1914) & (!g3136) & (g5342) & (g5343) & (!key[249])) + ((g830) & (!g1914) & (!g3136) & (g5342) & (g5343) & (key[249])) + ((g830) & (!g1914) & (g3136) & (!g5342) & (!g5343) & (!key[249])) + ((g830) & (!g1914) & (g3136) & (!g5342) & (!g5343) & (key[249])) + ((g830) & (!g1914) & (g3136) & (g5342) & (!g5343) & (!key[249])) + ((g830) & (!g1914) & (g3136) & (g5342) & (!g5343) & (key[249])) + ((g830) & (g1914) & (!g3136) & (g5342) & (!g5343) & (!key[249])) + ((g830) & (g1914) & (!g3136) & (g5342) & (!g5343) & (key[249])) + ((g830) & (g1914) & (!g3136) & (g5342) & (g5343) & (!key[249])) + ((g830) & (g1914) & (!g3136) & (g5342) & (g5343) & (key[249])) + ((g830) & (g1914) & (g3136) & (!g5342) & (!g5343) & (!key[249])) + ((g830) & (g1914) & (g3136) & (!g5342) & (!g5343) & (key[249])) + ((g830) & (g1914) & (g3136) & (!g5342) & (g5343) & (!key[249])) + ((g830) & (g1914) & (g3136) & (!g5342) & (g5343) & (key[249])));
	assign g5345 = (((!g3719) & (!g3720)));
	assign g5346 = (((g1914) & (!g2101) & (!g2752) & (!g5345)) + ((g1914) & (!g2101) & (g2752) & (g5345)) + ((g1914) & (g2101) & (!g2752) & (g5345)) + ((g1914) & (g2101) & (g2752) & (!g5345)));
	assign g5347 = (((!g3736) & (!g3737)));
	assign g5348 = (((!g1914) & (!g2728) & (!g2723) & (!g5347)) + ((!g1914) & (!g2728) & (g2723) & (g5347)) + ((!g1914) & (g2728) & (!g2723) & (g5347)) + ((!g1914) & (g2728) & (g2723) & (!g5347)));
	assign g5349 = (((!g830) & (!g3139) & (!g5346) & (!g5348) & (key[217])) + ((!g830) & (!g3139) & (!g5346) & (g5348) & (key[217])) + ((!g830) & (!g3139) & (g5346) & (!g5348) & (key[217])) + ((!g830) & (!g3139) & (g5346) & (g5348) & (key[217])) + ((!g830) & (g3139) & (!g5346) & (!g5348) & (key[217])) + ((!g830) & (g3139) & (!g5346) & (g5348) & (key[217])) + ((!g830) & (g3139) & (g5346) & (!g5348) & (key[217])) + ((!g830) & (g3139) & (g5346) & (g5348) & (key[217])) + ((g830) & (!g3139) & (!g5346) & (g5348) & (!key[217])) + ((g830) & (!g3139) & (!g5346) & (g5348) & (key[217])) + ((g830) & (!g3139) & (g5346) & (!g5348) & (!key[217])) + ((g830) & (!g3139) & (g5346) & (!g5348) & (key[217])) + ((g830) & (!g3139) & (g5346) & (g5348) & (!key[217])) + ((g830) & (!g3139) & (g5346) & (g5348) & (key[217])) + ((g830) & (g3139) & (!g5346) & (!g5348) & (!key[217])) + ((g830) & (g3139) & (!g5346) & (!g5348) & (key[217])));
	assign g5350 = (((!g2230) & (!g2286) & (!g2242) & (g2288) & (!g5310)) + ((!g2230) & (!g2286) & (!g2242) & (g2288) & (g5310)) + ((!g2230) & (!g2286) & (g2242) & (!g2288) & (!g5310)) + ((!g2230) & (!g2286) & (g2242) & (g2288) & (g5310)) + ((!g2230) & (g2286) & (!g2242) & (!g2288) & (!g5310)) + ((!g2230) & (g2286) & (!g2242) & (!g2288) & (g5310)) + ((!g2230) & (g2286) & (g2242) & (!g2288) & (g5310)) + ((!g2230) & (g2286) & (g2242) & (g2288) & (!g5310)) + ((g2230) & (!g2286) & (!g2242) & (!g2288) & (!g5310)) + ((g2230) & (!g2286) & (!g2242) & (g2288) & (g5310)) + ((g2230) & (!g2286) & (g2242) & (!g2288) & (!g5310)) + ((g2230) & (!g2286) & (g2242) & (!g2288) & (g5310)) + ((g2230) & (g2286) & (!g2242) & (!g2288) & (g5310)) + ((g2230) & (g2286) & (!g2242) & (g2288) & (!g5310)) + ((g2230) & (g2286) & (g2242) & (g2288) & (!g5310)) + ((g2230) & (g2286) & (g2242) & (g2288) & (g5310)));
	assign g5351 = (((!g2247) & (!g2275) & (!g2250) & (g2283) & (!g5312)) + ((!g2247) & (!g2275) & (!g2250) & (g2283) & (g5312)) + ((!g2247) & (!g2275) & (g2250) & (!g2283) & (!g5312)) + ((!g2247) & (!g2275) & (g2250) & (g2283) & (g5312)) + ((!g2247) & (g2275) & (!g2250) & (!g2283) & (!g5312)) + ((!g2247) & (g2275) & (!g2250) & (!g2283) & (g5312)) + ((!g2247) & (g2275) & (g2250) & (!g2283) & (g5312)) + ((!g2247) & (g2275) & (g2250) & (g2283) & (!g5312)) + ((g2247) & (!g2275) & (!g2250) & (!g2283) & (!g5312)) + ((g2247) & (!g2275) & (!g2250) & (g2283) & (g5312)) + ((g2247) & (!g2275) & (g2250) & (!g2283) & (!g5312)) + ((g2247) & (!g2275) & (g2250) & (!g2283) & (g5312)) + ((g2247) & (g2275) & (!g2250) & (!g2283) & (g5312)) + ((g2247) & (g2275) & (!g2250) & (g2283) & (!g5312)) + ((g2247) & (g2275) & (g2250) & (g2283) & (!g5312)) + ((g2247) & (g2275) & (g2250) & (g2283) & (g5312)));
	assign g5352 = (((!g830) & (!g1914) & (!g3142) & (!g5350) & (!g5351)) + ((!g830) & (!g1914) & (!g3142) & (!g5350) & (g5351)) + ((!g830) & (!g1914) & (!g3142) & (g5350) & (!g5351)) + ((!g830) & (!g1914) & (!g3142) & (g5350) & (g5351)) + ((!g830) & (!g1914) & (g3142) & (!g5350) & (!g5351)) + ((!g830) & (!g1914) & (g3142) & (!g5350) & (g5351)) + ((!g830) & (!g1914) & (g3142) & (g5350) & (!g5351)) + ((!g830) & (!g1914) & (g3142) & (g5350) & (g5351)) + ((!g830) & (g1914) & (!g3142) & (!g5350) & (!g5351)) + ((!g830) & (g1914) & (!g3142) & (!g5350) & (g5351)) + ((!g830) & (g1914) & (!g3142) & (g5350) & (!g5351)) + ((!g830) & (g1914) & (!g3142) & (g5350) & (g5351)) + ((!g830) & (g1914) & (g3142) & (!g5350) & (!g5351)) + ((!g830) & (g1914) & (g3142) & (!g5350) & (g5351)) + ((!g830) & (g1914) & (g3142) & (g5350) & (!g5351)) + ((!g830) & (g1914) & (g3142) & (g5350) & (g5351)) + ((g830) & (!g1914) & (!g3142) & (!g5350) & (g5351)) + ((g830) & (!g1914) & (!g3142) & (g5350) & (g5351)) + ((g830) & (!g1914) & (g3142) & (!g5350) & (!g5351)) + ((g830) & (!g1914) & (g3142) & (g5350) & (!g5351)) + ((g830) & (g1914) & (!g3142) & (g5350) & (!g5351)) + ((g830) & (g1914) & (!g3142) & (g5350) & (g5351)) + ((g830) & (g1914) & (g3142) & (!g5350) & (!g5351)) + ((g830) & (g1914) & (g3142) & (!g5350) & (g5351)));
	assign g5353 = (((!g2181) & (g1439) & (!g3455)) + ((g2181) & (!g1439) & (!g3455)) + ((g2181) & (g1439) & (!g3455)) + ((g2181) & (g1439) & (g3455)));
	assign g5354 = (((!g3438) & (!g2578) & (!g2584)) + ((!g3438) & (g2578) & (g2584)) + ((g3438) & (!g2578) & (g2584)) + ((g3438) & (g2578) & (!g2584)));
	assign g5355 = (((!g1914) & (!g2213) & (!g1473) & (g5353) & (!g5354)) + ((!g1914) & (!g2213) & (!g1473) & (g5353) & (g5354)) + ((!g1914) & (!g2213) & (g1473) & (!g5353) & (!g5354)) + ((!g1914) & (!g2213) & (g1473) & (!g5353) & (g5354)) + ((!g1914) & (g2213) & (!g1473) & (!g5353) & (!g5354)) + ((!g1914) & (g2213) & (!g1473) & (!g5353) & (g5354)) + ((!g1914) & (g2213) & (g1473) & (g5353) & (!g5354)) + ((!g1914) & (g2213) & (g1473) & (g5353) & (g5354)) + ((g1914) & (!g2213) & (!g1473) & (!g5353) & (g5354)) + ((g1914) & (!g2213) & (!g1473) & (g5353) & (g5354)) + ((g1914) & (!g2213) & (g1473) & (!g5353) & (g5354)) + ((g1914) & (!g2213) & (g1473) & (g5353) & (g5354)) + ((g1914) & (g2213) & (!g1473) & (!g5353) & (g5354)) + ((g1914) & (g2213) & (!g1473) & (g5353) & (g5354)) + ((g1914) & (g2213) & (g1473) & (!g5353) & (g5354)) + ((g1914) & (g2213) & (g1473) & (g5353) & (g5354)));
	assign g5356 = (((!g830) & (!g3149) & (!g5355) & (key[122])) + ((!g830) & (!g3149) & (g5355) & (key[122])) + ((!g830) & (g3149) & (!g5355) & (key[122])) + ((!g830) & (g3149) & (g5355) & (key[122])) + ((g830) & (!g3149) & (g5355) & (!key[122])) + ((g830) & (!g3149) & (g5355) & (key[122])) + ((g830) & (g3149) & (!g5355) & (!key[122])) + ((g830) & (g3149) & (!g5355) & (key[122])));
	assign g5357 = (((!g1958) & (!g2314) & (!g3548)) + ((!g1958) & (g2314) & (g3548)) + ((g1958) & (!g2314) & (g3548)) + ((g1958) & (g2314) & (!g3548)));
	assign g5358 = (((!g2797) & (!g3566) & (g2819)) + ((g2797) & (!g3566) & (!g2819)) + ((g2797) & (!g3566) & (g2819)) + ((g2797) & (g3566) & (g2819)));
	assign g5359 = (((!g1972) & (!g2589) & (!g3580)) + ((!g1972) & (g2589) & (g3580)) + ((g1972) & (!g2589) & (g3580)) + ((g1972) & (g2589) & (!g3580)));
	assign g5360 = (((!g1914) & (!g2854) & (!g5358) & (!g2860) & (g5359)) + ((!g1914) & (!g2854) & (!g5358) & (g2860) & (g5359)) + ((!g1914) & (!g2854) & (g5358) & (!g2860) & (g5359)) + ((!g1914) & (!g2854) & (g5358) & (g2860) & (g5359)) + ((!g1914) & (g2854) & (!g5358) & (!g2860) & (g5359)) + ((!g1914) & (g2854) & (!g5358) & (g2860) & (g5359)) + ((!g1914) & (g2854) & (g5358) & (!g2860) & (g5359)) + ((!g1914) & (g2854) & (g5358) & (g2860) & (g5359)) + ((g1914) & (!g2854) & (!g5358) & (g2860) & (!g5359)) + ((g1914) & (!g2854) & (!g5358) & (g2860) & (g5359)) + ((g1914) & (!g2854) & (g5358) & (!g2860) & (!g5359)) + ((g1914) & (!g2854) & (g5358) & (!g2860) & (g5359)) + ((g1914) & (g2854) & (!g5358) & (!g2860) & (!g5359)) + ((g1914) & (g2854) & (!g5358) & (!g2860) & (g5359)) + ((g1914) & (g2854) & (g5358) & (g2860) & (!g5359)) + ((g1914) & (g2854) & (g5358) & (g2860) & (g5359)));
	assign g5361 = (((!g830) & (!g3155) & (!g5360) & (nonce[26])) + ((!g830) & (!g3155) & (g5360) & (nonce[26])) + ((!g830) & (g3155) & (!g5360) & (nonce[26])) + ((!g830) & (g3155) & (g5360) & (nonce[26])) + ((g830) & (!g3155) & (g5360) & (!nonce[26])) + ((g830) & (!g3155) & (g5360) & (nonce[26])) + ((g830) & (g3155) & (!g5360) & (!nonce[26])) + ((g830) & (g3155) & (!g5360) & (nonce[26])));
	assign g5362 = (((!g2804) & (g2807) & (!g3613)) + ((g2804) & (!g2807) & (!g3613)) + ((g2804) & (g2807) & (!g3613)) + ((g2804) & (g2807) & (g3613)));
	assign g5363 = (((!g2012) & (!g3596) & (!g2592)) + ((!g2012) & (g3596) & (g2592)) + ((g2012) & (!g3596) & (g2592)) + ((g2012) & (g3596) & (!g2592)));
	assign g5364 = (((!g1914) & (!g2845) & (!g2857) & (g5362) & (!g5363)) + ((!g1914) & (!g2845) & (!g2857) & (g5362) & (g5363)) + ((!g1914) & (!g2845) & (g2857) & (!g5362) & (!g5363)) + ((!g1914) & (!g2845) & (g2857) & (!g5362) & (g5363)) + ((!g1914) & (g2845) & (!g2857) & (!g5362) & (!g5363)) + ((!g1914) & (g2845) & (!g2857) & (!g5362) & (g5363)) + ((!g1914) & (g2845) & (g2857) & (g5362) & (!g5363)) + ((!g1914) & (g2845) & (g2857) & (g5362) & (g5363)) + ((g1914) & (!g2845) & (!g2857) & (!g5362) & (g5363)) + ((g1914) & (!g2845) & (!g2857) & (g5362) & (g5363)) + ((g1914) & (!g2845) & (g2857) & (!g5362) & (g5363)) + ((g1914) & (!g2845) & (g2857) & (g5362) & (g5363)) + ((g1914) & (g2845) & (!g2857) & (!g5362) & (g5363)) + ((g1914) & (g2845) & (!g2857) & (g5362) & (g5363)) + ((g1914) & (g2845) & (g2857) & (!g5362) & (g5363)) + ((g1914) & (g2845) & (g2857) & (g5362) & (g5363)));
	assign g5365 = (((!g830) & (!g3157) & (!g5364) & (key[250])) + ((!g830) & (!g3157) & (g5364) & (key[250])) + ((!g830) & (g3157) & (!g5364) & (key[250])) + ((!g830) & (g3157) & (g5364) & (key[250])) + ((g830) & (!g3157) & (g5364) & (!key[250])) + ((g830) & (!g3157) & (g5364) & (key[250])) + ((g830) & (g3157) & (!g5364) & (!key[250])) + ((g830) & (g3157) & (!g5364) & (key[250])));
	assign g5366 = (((!g2178) & (g1439) & (!g3632)) + ((g2178) & (!g1439) & (!g3632)) + ((g2178) & (g1439) & (!g3632)) + ((g2178) & (g1439) & (g3632)));
	assign g5367 = (((!g2569) & (!g2592) & (!g3646)) + ((!g2569) & (g2592) & (g3646)) + ((g2569) & (!g2592) & (g3646)) + ((g2569) & (g2592) & (!g3646)));
	assign g5368 = (((!g1914) & (!g2211) & (!g1473) & (!g5366) & (g5367)) + ((!g1914) & (!g2211) & (!g1473) & (g5366) & (g5367)) + ((!g1914) & (!g2211) & (g1473) & (!g5366) & (g5367)) + ((!g1914) & (!g2211) & (g1473) & (g5366) & (g5367)) + ((!g1914) & (g2211) & (!g1473) & (!g5366) & (g5367)) + ((!g1914) & (g2211) & (!g1473) & (g5366) & (g5367)) + ((!g1914) & (g2211) & (g1473) & (!g5366) & (g5367)) + ((!g1914) & (g2211) & (g1473) & (g5366) & (g5367)) + ((g1914) & (!g2211) & (!g1473) & (g5366) & (!g5367)) + ((g1914) & (!g2211) & (!g1473) & (g5366) & (g5367)) + ((g1914) & (!g2211) & (g1473) & (!g5366) & (!g5367)) + ((g1914) & (!g2211) & (g1473) & (!g5366) & (g5367)) + ((g1914) & (g2211) & (!g1473) & (!g5366) & (!g5367)) + ((g1914) & (g2211) & (!g1473) & (!g5366) & (g5367)) + ((g1914) & (g2211) & (g1473) & (g5366) & (!g5367)) + ((g1914) & (g2211) & (g1473) & (g5366) & (g5367)));
	assign g5369 = (((!g830) & (!g3159) & (!g5368) & (key[26])) + ((!g830) & (!g3159) & (g5368) & (key[26])) + ((!g830) & (g3159) & (!g5368) & (key[26])) + ((!g830) & (g3159) & (g5368) & (key[26])) + ((g830) & (!g3159) & (g5368) & (!key[26])) + ((g830) & (!g3159) & (g5368) & (key[26])) + ((g830) & (g3159) & (!g5368) & (!key[26])) + ((g830) & (g3159) & (!g5368) & (key[26])));
	assign g5370 = (((!g2813) & (g2819) & (!g3680)) + ((g2813) & (!g2819) & (!g3680)) + ((g2813) & (g2819) & (!g3680)) + ((g2813) & (g2819) & (g3680)));
	assign g5371 = (((!g2011) & (!g2572) & (!g3662)) + ((!g2011) & (g2572) & (g3662)) + ((g2011) & (!g2572) & (g3662)) + ((g2011) & (g2572) & (!g3662)));
	assign g5372 = (((!g1914) & (!g2838) & (!g2860) & (g5370) & (!g5371)) + ((!g1914) & (!g2838) & (!g2860) & (g5370) & (g5371)) + ((!g1914) & (!g2838) & (g2860) & (!g5370) & (!g5371)) + ((!g1914) & (!g2838) & (g2860) & (!g5370) & (g5371)) + ((!g1914) & (g2838) & (!g2860) & (!g5370) & (!g5371)) + ((!g1914) & (g2838) & (!g2860) & (!g5370) & (g5371)) + ((!g1914) & (g2838) & (g2860) & (g5370) & (!g5371)) + ((!g1914) & (g2838) & (g2860) & (g5370) & (g5371)) + ((g1914) & (!g2838) & (!g2860) & (!g5370) & (g5371)) + ((g1914) & (!g2838) & (!g2860) & (g5370) & (g5371)) + ((g1914) & (!g2838) & (g2860) & (!g5370) & (g5371)) + ((g1914) & (!g2838) & (g2860) & (g5370) & (g5371)) + ((g1914) & (g2838) & (!g2860) & (!g5370) & (g5371)) + ((g1914) & (g2838) & (!g2860) & (g5370) & (g5371)) + ((g1914) & (g2838) & (g2860) & (!g5370) & (g5371)) + ((g1914) & (g2838) & (g2860) & (g5370) & (g5371)));
	assign g8334 = (((!g5560) & (g5640) & (!g5373)) + ((!g5560) & (g5640) & (g5373)) + ((g5560) & (!g5640) & (g5373)) + ((g5560) & (g5640) & (g5373)));
	assign g5374 = (((!g830) & (!g3161) & (!g5372) & (g5373)) + ((!g830) & (!g3161) & (g5372) & (g5373)) + ((!g830) & (g3161) & (!g5372) & (g5373)) + ((!g830) & (g3161) & (g5372) & (g5373)) + ((g830) & (!g3161) & (g5372) & (!g5373)) + ((g830) & (!g3161) & (g5372) & (g5373)) + ((g830) & (g3161) & (!g5372) & (!g5373)) + ((g830) & (g3161) & (!g5372) & (g5373)));
	assign g5375 = (((!g2320) & (!g2329) & (!g3703)) + ((!g2320) & (g2329) & (g3703)) + ((g2320) & (!g2329) & (g3703)) + ((g2320) & (g2329) & (!g3703)));
	assign g5376 = (((!g2101) & (!g2134) & (!g2752) & (g2787) & (!g5345)) + ((!g2101) & (!g2134) & (!g2752) & (g2787) & (g5345)) + ((!g2101) & (!g2134) & (g2752) & (!g2787) & (!g5345)) + ((!g2101) & (!g2134) & (g2752) & (g2787) & (g5345)) + ((!g2101) & (g2134) & (!g2752) & (!g2787) & (!g5345)) + ((!g2101) & (g2134) & (!g2752) & (!g2787) & (g5345)) + ((!g2101) & (g2134) & (g2752) & (!g2787) & (g5345)) + ((!g2101) & (g2134) & (g2752) & (g2787) & (!g5345)) + ((g2101) & (!g2134) & (!g2752) & (!g2787) & (!g5345)) + ((g2101) & (!g2134) & (!g2752) & (g2787) & (g5345)) + ((g2101) & (!g2134) & (g2752) & (!g2787) & (!g5345)) + ((g2101) & (!g2134) & (g2752) & (!g2787) & (g5345)) + ((g2101) & (g2134) & (!g2752) & (!g2787) & (g5345)) + ((g2101) & (g2134) & (!g2752) & (g2787) & (!g5345)) + ((g2101) & (g2134) & (g2752) & (g2787) & (!g5345)) + ((g2101) & (g2134) & (g2752) & (g2787) & (g5345)));
	assign g5377 = (((!g2728) & (!g2778) & (!g2723) & (g2770) & (!g5347)) + ((!g2728) & (!g2778) & (!g2723) & (g2770) & (g5347)) + ((!g2728) & (!g2778) & (g2723) & (!g2770) & (!g5347)) + ((!g2728) & (!g2778) & (g2723) & (g2770) & (g5347)) + ((!g2728) & (g2778) & (!g2723) & (!g2770) & (!g5347)) + ((!g2728) & (g2778) & (!g2723) & (!g2770) & (g5347)) + ((!g2728) & (g2778) & (g2723) & (!g2770) & (g5347)) + ((!g2728) & (g2778) & (g2723) & (g2770) & (!g5347)) + ((g2728) & (!g2778) & (!g2723) & (!g2770) & (!g5347)) + ((g2728) & (!g2778) & (!g2723) & (g2770) & (g5347)) + ((g2728) & (!g2778) & (g2723) & (!g2770) & (!g5347)) + ((g2728) & (!g2778) & (g2723) & (!g2770) & (g5347)) + ((g2728) & (g2778) & (!g2723) & (!g2770) & (g5347)) + ((g2728) & (g2778) & (!g2723) & (g2770) & (!g5347)) + ((g2728) & (g2778) & (g2723) & (g2770) & (!g5347)) + ((g2728) & (g2778) & (g2723) & (g2770) & (g5347)));
	assign g5378 = (((!g830) & (!g1914) & (!g3165) & (!g5376) & (!g5377) & (key[218])) + ((!g830) & (!g1914) & (!g3165) & (!g5376) & (g5377) & (key[218])) + ((!g830) & (!g1914) & (!g3165) & (g5376) & (!g5377) & (key[218])) + ((!g830) & (!g1914) & (!g3165) & (g5376) & (g5377) & (key[218])) + ((!g830) & (!g1914) & (g3165) & (!g5376) & (!g5377) & (key[218])) + ((!g830) & (!g1914) & (g3165) & (!g5376) & (g5377) & (key[218])) + ((!g830) & (!g1914) & (g3165) & (g5376) & (!g5377) & (key[218])) + ((!g830) & (!g1914) & (g3165) & (g5376) & (g5377) & (key[218])) + ((!g830) & (g1914) & (!g3165) & (!g5376) & (!g5377) & (key[218])) + ((!g830) & (g1914) & (!g3165) & (!g5376) & (g5377) & (key[218])) + ((!g830) & (g1914) & (!g3165) & (g5376) & (!g5377) & (key[218])) + ((!g830) & (g1914) & (!g3165) & (g5376) & (g5377) & (key[218])) + ((!g830) & (g1914) & (g3165) & (!g5376) & (!g5377) & (key[218])) + ((!g830) & (g1914) & (g3165) & (!g5376) & (g5377) & (key[218])) + ((!g830) & (g1914) & (g3165) & (g5376) & (!g5377) & (key[218])) + ((!g830) & (g1914) & (g3165) & (g5376) & (g5377) & (key[218])) + ((g830) & (!g1914) & (!g3165) & (!g5376) & (g5377) & (!key[218])) + ((g830) & (!g1914) & (!g3165) & (!g5376) & (g5377) & (key[218])) + ((g830) & (!g1914) & (!g3165) & (g5376) & (g5377) & (!key[218])) + ((g830) & (!g1914) & (!g3165) & (g5376) & (g5377) & (key[218])) + ((g830) & (!g1914) & (g3165) & (!g5376) & (!g5377) & (!key[218])) + ((g830) & (!g1914) & (g3165) & (!g5376) & (!g5377) & (key[218])) + ((g830) & (!g1914) & (g3165) & (g5376) & (!g5377) & (!key[218])) + ((g830) & (!g1914) & (g3165) & (g5376) & (!g5377) & (key[218])) + ((g830) & (g1914) & (!g3165) & (g5376) & (!g5377) & (!key[218])) + ((g830) & (g1914) & (!g3165) & (g5376) & (!g5377) & (key[218])) + ((g830) & (g1914) & (!g3165) & (g5376) & (g5377) & (!key[218])) + ((g830) & (g1914) & (!g3165) & (g5376) & (g5377) & (key[218])) + ((g830) & (g1914) & (g3165) & (!g5376) & (!g5377) & (!key[218])) + ((g830) & (g1914) & (g3165) & (!g5376) & (!g5377) & (key[218])) + ((g830) & (g1914) & (g3165) & (!g5376) & (g5377) & (!key[218])) + ((g830) & (g1914) & (g3165) & (!g5376) & (g5377) & (key[218])));
	assign g5379 = (((!g2804) & (g2816) & (!g3789)) + ((g2804) & (!g2816) & (!g3789)) + ((g2804) & (g2816) & (!g3789)) + ((g2804) & (g2816) & (g3789)));
	assign g5380 = (((!g1973) & (!g2584) & (!g3803)) + ((!g1973) & (g2584) & (g3803)) + ((g1973) & (!g2584) & (g3803)) + ((g1973) & (g2584) & (!g3803)));
	assign g5381 = (((!g1914) & (!g2845) & (!g2848) & (!g5379) & (g5380)) + ((!g1914) & (!g2845) & (!g2848) & (g5379) & (g5380)) + ((!g1914) & (!g2845) & (g2848) & (!g5379) & (g5380)) + ((!g1914) & (!g2845) & (g2848) & (g5379) & (g5380)) + ((!g1914) & (g2845) & (!g2848) & (!g5379) & (g5380)) + ((!g1914) & (g2845) & (!g2848) & (g5379) & (g5380)) + ((!g1914) & (g2845) & (g2848) & (!g5379) & (g5380)) + ((!g1914) & (g2845) & (g2848) & (g5379) & (g5380)) + ((g1914) & (!g2845) & (!g2848) & (g5379) & (!g5380)) + ((g1914) & (!g2845) & (!g2848) & (g5379) & (g5380)) + ((g1914) & (!g2845) & (g2848) & (!g5379) & (!g5380)) + ((g1914) & (!g2845) & (g2848) & (!g5379) & (g5380)) + ((g1914) & (g2845) & (!g2848) & (!g5379) & (!g5380)) + ((g1914) & (g2845) & (!g2848) & (!g5379) & (g5380)) + ((g1914) & (g2845) & (g2848) & (g5379) & (!g5380)) + ((g1914) & (g2845) & (g2848) & (g5379) & (g5380)));
	assign g5382 = (((!g830) & (!g3168) & (!g5381) & (key[154])) + ((!g830) & (!g3168) & (g5381) & (key[154])) + ((!g830) & (g3168) & (!g5381) & (key[154])) + ((!g830) & (g3168) & (g5381) & (key[154])) + ((g830) & (!g3168) & (g5381) & (!key[154])) + ((g830) & (!g3168) & (g5381) & (key[154])) + ((g830) & (g3168) & (!g5381) & (!key[154])) + ((g830) & (g3168) & (!g5381) & (key[154])));
	assign g5383 = (((!g2708) & (!g2776) & (!g2728) & (g2778) & (!g5337)) + ((!g2708) & (!g2776) & (!g2728) & (g2778) & (g5337)) + ((!g2708) & (!g2776) & (g2728) & (!g2778) & (!g5337)) + ((!g2708) & (!g2776) & (g2728) & (g2778) & (g5337)) + ((!g2708) & (g2776) & (!g2728) & (!g2778) & (!g5337)) + ((!g2708) & (g2776) & (!g2728) & (!g2778) & (g5337)) + ((!g2708) & (g2776) & (g2728) & (!g2778) & (g5337)) + ((!g2708) & (g2776) & (g2728) & (g2778) & (!g5337)) + ((g2708) & (!g2776) & (!g2728) & (!g2778) & (!g5337)) + ((g2708) & (!g2776) & (!g2728) & (g2778) & (g5337)) + ((g2708) & (!g2776) & (g2728) & (!g2778) & (!g5337)) + ((g2708) & (!g2776) & (g2728) & (!g2778) & (g5337)) + ((g2708) & (g2776) & (!g2728) & (!g2778) & (g5337)) + ((g2708) & (g2776) & (!g2728) & (g2778) & (!g5337)) + ((g2708) & (g2776) & (g2728) & (g2778) & (!g5337)) + ((g2708) & (g2776) & (g2728) & (g2778) & (g5337)));
	assign g5384 = (((!g2099) & (!g2130) & (!g2752) & (g2787) & (!g5339)) + ((!g2099) & (!g2130) & (!g2752) & (g2787) & (g5339)) + ((!g2099) & (!g2130) & (g2752) & (!g2787) & (!g5339)) + ((!g2099) & (!g2130) & (g2752) & (g2787) & (g5339)) + ((!g2099) & (g2130) & (!g2752) & (!g2787) & (!g5339)) + ((!g2099) & (g2130) & (!g2752) & (!g2787) & (g5339)) + ((!g2099) & (g2130) & (g2752) & (!g2787) & (g5339)) + ((!g2099) & (g2130) & (g2752) & (g2787) & (!g5339)) + ((g2099) & (!g2130) & (!g2752) & (!g2787) & (!g5339)) + ((g2099) & (!g2130) & (!g2752) & (g2787) & (g5339)) + ((g2099) & (!g2130) & (g2752) & (!g2787) & (!g5339)) + ((g2099) & (!g2130) & (g2752) & (!g2787) & (g5339)) + ((g2099) & (g2130) & (!g2752) & (!g2787) & (g5339)) + ((g2099) & (g2130) & (!g2752) & (g2787) & (!g5339)) + ((g2099) & (g2130) & (g2752) & (g2787) & (!g5339)) + ((g2099) & (g2130) & (g2752) & (g2787) & (g5339)));
	assign g5385 = (((!g830) & (!g1914) & (!g3170) & (!g5383) & (!g5384) & (nonce[58])) + ((!g830) & (!g1914) & (!g3170) & (!g5383) & (g5384) & (nonce[58])) + ((!g830) & (!g1914) & (!g3170) & (g5383) & (!g5384) & (nonce[58])) + ((!g830) & (!g1914) & (!g3170) & (g5383) & (g5384) & (nonce[58])) + ((!g830) & (!g1914) & (g3170) & (!g5383) & (!g5384) & (nonce[58])) + ((!g830) & (!g1914) & (g3170) & (!g5383) & (g5384) & (nonce[58])) + ((!g830) & (!g1914) & (g3170) & (g5383) & (!g5384) & (nonce[58])) + ((!g830) & (!g1914) & (g3170) & (g5383) & (g5384) & (nonce[58])) + ((!g830) & (g1914) & (!g3170) & (!g5383) & (!g5384) & (nonce[58])) + ((!g830) & (g1914) & (!g3170) & (!g5383) & (g5384) & (nonce[58])) + ((!g830) & (g1914) & (!g3170) & (g5383) & (!g5384) & (nonce[58])) + ((!g830) & (g1914) & (!g3170) & (g5383) & (g5384) & (nonce[58])) + ((!g830) & (g1914) & (g3170) & (!g5383) & (!g5384) & (nonce[58])) + ((!g830) & (g1914) & (g3170) & (!g5383) & (g5384) & (nonce[58])) + ((!g830) & (g1914) & (g3170) & (g5383) & (!g5384) & (nonce[58])) + ((!g830) & (g1914) & (g3170) & (g5383) & (g5384) & (nonce[58])) + ((g830) & (!g1914) & (!g3170) & (!g5383) & (g5384) & (!nonce[58])) + ((g830) & (!g1914) & (!g3170) & (!g5383) & (g5384) & (nonce[58])) + ((g830) & (!g1914) & (!g3170) & (g5383) & (g5384) & (!nonce[58])) + ((g830) & (!g1914) & (!g3170) & (g5383) & (g5384) & (nonce[58])) + ((g830) & (!g1914) & (g3170) & (!g5383) & (!g5384) & (!nonce[58])) + ((g830) & (!g1914) & (g3170) & (!g5383) & (!g5384) & (nonce[58])) + ((g830) & (!g1914) & (g3170) & (g5383) & (!g5384) & (!nonce[58])) + ((g830) & (!g1914) & (g3170) & (g5383) & (!g5384) & (nonce[58])) + ((g830) & (g1914) & (!g3170) & (g5383) & (!g5384) & (!nonce[58])) + ((g830) & (g1914) & (!g3170) & (g5383) & (!g5384) & (nonce[58])) + ((g830) & (g1914) & (!g3170) & (g5383) & (g5384) & (!nonce[58])) + ((g830) & (g1914) & (!g3170) & (g5383) & (g5384) & (nonce[58])) + ((g830) & (g1914) & (g3170) & (!g5383) & (!g5384) & (!nonce[58])) + ((g830) & (g1914) & (g3170) & (!g5383) & (!g5384) & (nonce[58])) + ((g830) & (g1914) & (g3170) & (!g5383) & (g5384) & (!nonce[58])) + ((g830) & (g1914) & (g3170) & (!g5383) & (g5384) & (nonce[58])));
	assign g5386 = (((!g2334) & (!g2337) & (!g3860)) + ((!g2334) & (g2337) & (g3860)) + ((g2334) & (!g2337) & (g3860)) + ((g2334) & (g2337) & (!g3860)));
	assign g5387 = (((!g2569) & (!g2626) & (!g2592) & (g2632) & (!g3646)) + ((!g2569) & (!g2626) & (!g2592) & (g2632) & (g3646)) + ((!g2569) & (!g2626) & (g2592) & (!g2632) & (!g3646)) + ((!g2569) & (!g2626) & (g2592) & (g2632) & (g3646)) + ((!g2569) & (g2626) & (!g2592) & (!g2632) & (!g3646)) + ((!g2569) & (g2626) & (!g2592) & (!g2632) & (g3646)) + ((!g2569) & (g2626) & (g2592) & (!g2632) & (g3646)) + ((!g2569) & (g2626) & (g2592) & (g2632) & (!g3646)) + ((g2569) & (!g2626) & (!g2592) & (!g2632) & (!g3646)) + ((g2569) & (!g2626) & (!g2592) & (g2632) & (g3646)) + ((g2569) & (!g2626) & (g2592) & (!g2632) & (!g3646)) + ((g2569) & (!g2626) & (g2592) & (!g2632) & (g3646)) + ((g2569) & (g2626) & (!g2592) & (!g2632) & (g3646)) + ((g2569) & (g2626) & (!g2592) & (g2632) & (!g3646)) + ((g2569) & (g2626) & (g2592) & (g2632) & (!g3646)) + ((g2569) & (g2626) & (g2592) & (g2632) & (g3646)));
	assign g5388 = (((!g830) & (!g3177) & (!g5999) & (key[27])) + ((!g830) & (!g3177) & (g5999) & (key[27])) + ((!g830) & (g3177) & (!g5999) & (key[27])) + ((!g830) & (g3177) & (g5999) & (key[27])) + ((g830) & (!g3177) & (g5999) & (!key[27])) + ((g830) & (!g3177) & (g5999) & (key[27])) + ((g830) & (g3177) & (!g5999) & (!key[27])) + ((g830) & (g3177) & (!g5999) & (key[27])));
	assign g5389 = (((!g1996) & (g3539) & (g2323)) + ((g1996) & (!g3539) & (g2323)) + ((g1996) & (g3539) & (!g2323)) + ((g1996) & (g3539) & (g2323)));
	assign g5390 = (((!g1958) & (!g1960) & (!g2314) & (g2362) & (!g3548)) + ((!g1958) & (!g1960) & (!g2314) & (g2362) & (g3548)) + ((!g1958) & (!g1960) & (g2314) & (!g2362) & (!g3548)) + ((!g1958) & (!g1960) & (g2314) & (g2362) & (g3548)) + ((!g1958) & (g1960) & (!g2314) & (!g2362) & (!g3548)) + ((!g1958) & (g1960) & (!g2314) & (!g2362) & (g3548)) + ((!g1958) & (g1960) & (g2314) & (!g2362) & (g3548)) + ((!g1958) & (g1960) & (g2314) & (g2362) & (!g3548)) + ((g1958) & (!g1960) & (!g2314) & (!g2362) & (!g3548)) + ((g1958) & (!g1960) & (!g2314) & (g2362) & (g3548)) + ((g1958) & (!g1960) & (g2314) & (!g2362) & (!g3548)) + ((g1958) & (!g1960) & (g2314) & (!g2362) & (g3548)) + ((g1958) & (g1960) & (!g2314) & (!g2362) & (g3548)) + ((g1958) & (g1960) & (!g2314) & (g2362) & (!g3548)) + ((g1958) & (g1960) & (g2314) & (g2362) & (!g3548)) + ((g1958) & (g1960) & (g2314) & (g2362) & (g3548)));
	assign g5391 = (((!g2011) & (!g2013) & (!g2572) & (g2637) & (!g3662)) + ((!g2011) & (!g2013) & (!g2572) & (g2637) & (g3662)) + ((!g2011) & (!g2013) & (g2572) & (!g2637) & (!g3662)) + ((!g2011) & (!g2013) & (g2572) & (g2637) & (g3662)) + ((!g2011) & (g2013) & (!g2572) & (!g2637) & (!g3662)) + ((!g2011) & (g2013) & (!g2572) & (!g2637) & (g3662)) + ((!g2011) & (g2013) & (g2572) & (!g2637) & (g3662)) + ((!g2011) & (g2013) & (g2572) & (g2637) & (!g3662)) + ((g2011) & (!g2013) & (!g2572) & (!g2637) & (!g3662)) + ((g2011) & (!g2013) & (!g2572) & (g2637) & (g3662)) + ((g2011) & (!g2013) & (g2572) & (!g2637) & (!g3662)) + ((g2011) & (!g2013) & (g2572) & (!g2637) & (g3662)) + ((g2011) & (g2013) & (!g2572) & (!g2637) & (g3662)) + ((g2011) & (g2013) & (!g2572) & (g2637) & (!g3662)) + ((g2011) & (g2013) & (g2572) & (g2637) & (!g3662)) + ((g2011) & (g2013) & (g2572) & (g2637) & (g3662)));
	assign g5392 = (((!g2838) & (!g2891) & (!g2860) & (g2895) & (!g5370)) + ((!g2838) & (!g2891) & (!g2860) & (g2895) & (g5370)) + ((!g2838) & (!g2891) & (g2860) & (!g2895) & (g5370)) + ((!g2838) & (!g2891) & (g2860) & (g2895) & (!g5370)) + ((!g2838) & (g2891) & (!g2860) & (!g2895) & (!g5370)) + ((!g2838) & (g2891) & (!g2860) & (!g2895) & (g5370)) + ((!g2838) & (g2891) & (g2860) & (!g2895) & (!g5370)) + ((!g2838) & (g2891) & (g2860) & (g2895) & (g5370)) + ((g2838) & (!g2891) & (!g2860) & (!g2895) & (g5370)) + ((g2838) & (!g2891) & (!g2860) & (g2895) & (!g5370)) + ((g2838) & (!g2891) & (g2860) & (!g2895) & (!g5370)) + ((g2838) & (!g2891) & (g2860) & (!g2895) & (g5370)) + ((g2838) & (g2891) & (!g2860) & (!g2895) & (!g5370)) + ((g2838) & (g2891) & (!g2860) & (g2895) & (g5370)) + ((g2838) & (g2891) & (g2860) & (g2895) & (!g5370)) + ((g2838) & (g2891) & (g2860) & (g2895) & (g5370)));
	assign g8335 = (((!g5560) & (g5642) & (!g5393)) + ((!g5560) & (g5642) & (g5393)) + ((g5560) & (!g5642) & (g5393)) + ((g5560) & (g5642) & (g5393)));
	assign g5394 = (((!g830) & (!g1914) & (!g3187) & (!g5391) & (!g5392) & (g5393)) + ((!g830) & (!g1914) & (!g3187) & (!g5391) & (g5392) & (g5393)) + ((!g830) & (!g1914) & (!g3187) & (g5391) & (!g5392) & (g5393)) + ((!g830) & (!g1914) & (!g3187) & (g5391) & (g5392) & (g5393)) + ((!g830) & (!g1914) & (g3187) & (!g5391) & (!g5392) & (g5393)) + ((!g830) & (!g1914) & (g3187) & (!g5391) & (g5392) & (g5393)) + ((!g830) & (!g1914) & (g3187) & (g5391) & (!g5392) & (g5393)) + ((!g830) & (!g1914) & (g3187) & (g5391) & (g5392) & (g5393)) + ((!g830) & (g1914) & (!g3187) & (!g5391) & (!g5392) & (g5393)) + ((!g830) & (g1914) & (!g3187) & (!g5391) & (g5392) & (g5393)) + ((!g830) & (g1914) & (!g3187) & (g5391) & (!g5392) & (g5393)) + ((!g830) & (g1914) & (!g3187) & (g5391) & (g5392) & (g5393)) + ((!g830) & (g1914) & (g3187) & (!g5391) & (!g5392) & (g5393)) + ((!g830) & (g1914) & (g3187) & (!g5391) & (g5392) & (g5393)) + ((!g830) & (g1914) & (g3187) & (g5391) & (!g5392) & (g5393)) + ((!g830) & (g1914) & (g3187) & (g5391) & (g5392) & (g5393)) + ((g830) & (!g1914) & (!g3187) & (!g5391) & (g5392) & (!g5393)) + ((g830) & (!g1914) & (!g3187) & (!g5391) & (g5392) & (g5393)) + ((g830) & (!g1914) & (!g3187) & (g5391) & (g5392) & (!g5393)) + ((g830) & (!g1914) & (!g3187) & (g5391) & (g5392) & (g5393)) + ((g830) & (!g1914) & (g3187) & (!g5391) & (!g5392) & (!g5393)) + ((g830) & (!g1914) & (g3187) & (!g5391) & (!g5392) & (g5393)) + ((g830) & (!g1914) & (g3187) & (g5391) & (!g5392) & (!g5393)) + ((g830) & (!g1914) & (g3187) & (g5391) & (!g5392) & (g5393)) + ((g830) & (g1914) & (!g3187) & (g5391) & (!g5392) & (!g5393)) + ((g830) & (g1914) & (!g3187) & (g5391) & (!g5392) & (g5393)) + ((g830) & (g1914) & (!g3187) & (g5391) & (g5392) & (!g5393)) + ((g830) & (g1914) & (!g3187) & (g5391) & (g5392) & (g5393)) + ((g830) & (g1914) & (g3187) & (!g5391) & (!g5392) & (!g5393)) + ((g830) & (g1914) & (g3187) & (!g5391) & (!g5392) & (g5393)) + ((g830) & (g1914) & (g3187) & (!g5391) & (g5392) & (!g5393)) + ((g830) & (g1914) & (g3187) & (!g5391) & (g5392) & (g5393)));
	assign g5395 = (((!g1973) & (!g1976) & (!g2584) & (g2640) & (!g3803)) + ((!g1973) & (!g1976) & (!g2584) & (g2640) & (g3803)) + ((!g1973) & (!g1976) & (g2584) & (!g2640) & (!g3803)) + ((!g1973) & (!g1976) & (g2584) & (g2640) & (g3803)) + ((!g1973) & (g1976) & (!g2584) & (!g2640) & (!g3803)) + ((!g1973) & (g1976) & (!g2584) & (!g2640) & (g3803)) + ((!g1973) & (g1976) & (g2584) & (!g2640) & (g3803)) + ((!g1973) & (g1976) & (g2584) & (g2640) & (!g3803)) + ((g1973) & (!g1976) & (!g2584) & (!g2640) & (!g3803)) + ((g1973) & (!g1976) & (!g2584) & (g2640) & (g3803)) + ((g1973) & (!g1976) & (g2584) & (!g2640) & (!g3803)) + ((g1973) & (!g1976) & (g2584) & (!g2640) & (g3803)) + ((g1973) & (g1976) & (!g2584) & (!g2640) & (g3803)) + ((g1973) & (g1976) & (!g2584) & (g2640) & (!g3803)) + ((g1973) & (g1976) & (g2584) & (g2640) & (!g3803)) + ((g1973) & (g1976) & (g2584) & (g2640) & (g3803)));
	assign g5396 = (((!g830) & (!g3190) & (!g5981) & (key[155])) + ((!g830) & (!g3190) & (g5981) & (key[155])) + ((!g830) & (g3190) & (!g5981) & (key[155])) + ((!g830) & (g3190) & (g5981) & (key[155])) + ((g830) & (!g3190) & (g5981) & (!key[155])) + ((g830) & (!g3190) & (g5981) & (key[155])) + ((g830) & (g3190) & (!g5981) & (!key[155])) + ((g830) & (g3190) & (!g5981) & (key[155])));
	assign g5397 = (((!g3438) & (!g2578) & (!g2584) & (!g2617) & (g2640)) + ((!g3438) & (!g2578) & (!g2584) & (g2617) & (!g2640)) + ((!g3438) & (!g2578) & (g2584) & (!g2617) & (!g2640)) + ((!g3438) & (!g2578) & (g2584) & (g2617) & (g2640)) + ((!g3438) & (g2578) & (!g2584) & (!g2617) & (!g2640)) + ((!g3438) & (g2578) & (!g2584) & (g2617) & (g2640)) + ((!g3438) & (g2578) & (g2584) & (!g2617) & (!g2640)) + ((!g3438) & (g2578) & (g2584) & (g2617) & (g2640)) + ((g3438) & (!g2578) & (!g2584) & (!g2617) & (g2640)) + ((g3438) & (!g2578) & (!g2584) & (g2617) & (!g2640)) + ((g3438) & (!g2578) & (g2584) & (!g2617) & (g2640)) + ((g3438) & (!g2578) & (g2584) & (g2617) & (!g2640)) + ((g3438) & (g2578) & (!g2584) & (!g2617) & (g2640)) + ((g3438) & (g2578) & (!g2584) & (g2617) & (!g2640)) + ((g3438) & (g2578) & (g2584) & (!g2617) & (!g2640)) + ((g3438) & (g2578) & (g2584) & (g2617) & (g2640)));
	assign g5398 = (((!g830) & (!g3193) & (!g5970) & (key[123])) + ((!g830) & (!g3193) & (g5970) & (key[123])) + ((!g830) & (g3193) & (!g5970) & (key[123])) + ((!g830) & (g3193) & (g5970) & (key[123])) + ((g830) & (!g3193) & (g5970) & (!key[123])) + ((g830) & (!g3193) & (g5970) & (key[123])) + ((g830) & (g3193) & (!g5970) & (!key[123])) + ((g830) & (g3193) & (!g5970) & (key[123])));
	assign g5399 = (((!g1972) & (!g1975) & (!g2589) & (g2620) & (!g3580)) + ((!g1972) & (!g1975) & (!g2589) & (g2620) & (g3580)) + ((!g1972) & (!g1975) & (g2589) & (!g2620) & (!g3580)) + ((!g1972) & (!g1975) & (g2589) & (g2620) & (g3580)) + ((!g1972) & (g1975) & (!g2589) & (!g2620) & (!g3580)) + ((!g1972) & (g1975) & (!g2589) & (!g2620) & (g3580)) + ((!g1972) & (g1975) & (g2589) & (!g2620) & (g3580)) + ((!g1972) & (g1975) & (g2589) & (g2620) & (!g3580)) + ((g1972) & (!g1975) & (!g2589) & (!g2620) & (!g3580)) + ((g1972) & (!g1975) & (!g2589) & (g2620) & (g3580)) + ((g1972) & (!g1975) & (g2589) & (!g2620) & (!g3580)) + ((g1972) & (!g1975) & (g2589) & (!g2620) & (g3580)) + ((g1972) & (g1975) & (!g2589) & (!g2620) & (g3580)) + ((g1972) & (g1975) & (!g2589) & (g2620) & (!g3580)) + ((g1972) & (g1975) & (g2589) & (g2620) & (!g3580)) + ((g1972) & (g1975) & (g2589) & (g2620) & (g3580)));
	assign g5400 = (((!g830) & (!g3196) & (!g5959) & (nonce[27])) + ((!g830) & (!g3196) & (g5959) & (nonce[27])) + ((!g830) & (g3196) & (!g5959) & (nonce[27])) + ((!g830) & (g3196) & (g5959) & (nonce[27])) + ((g830) & (!g3196) & (g5959) & (!nonce[27])) + ((g830) & (!g3196) & (g5959) & (nonce[27])) + ((g830) & (g3196) & (!g5959) & (!nonce[27])) + ((g830) & (g3196) & (!g5959) & (nonce[27])));
	assign g5401 = (((!g2304) & (g2337) & (g3693)) + ((g2304) & (!g2337) & (g3693)) + ((g2304) & (g2337) & (!g3693)) + ((g2304) & (g2337) & (g3693)));
	assign g5402 = (((!g2320) & (!g2350) & (!g2329) & (g2371) & (!g3703)) + ((!g2320) & (!g2350) & (!g2329) & (g2371) & (g3703)) + ((!g2320) & (!g2350) & (g2329) & (!g2371) & (!g3703)) + ((!g2320) & (!g2350) & (g2329) & (g2371) & (g3703)) + ((!g2320) & (g2350) & (!g2329) & (!g2371) & (!g3703)) + ((!g2320) & (g2350) & (!g2329) & (!g2371) & (g3703)) + ((!g2320) & (g2350) & (g2329) & (!g2371) & (g3703)) + ((!g2320) & (g2350) & (g2329) & (g2371) & (!g3703)) + ((g2320) & (!g2350) & (!g2329) & (!g2371) & (!g3703)) + ((g2320) & (!g2350) & (!g2329) & (g2371) & (g3703)) + ((g2320) & (!g2350) & (g2329) & (!g2371) & (!g3703)) + ((g2320) & (!g2350) & (g2329) & (!g2371) & (g3703)) + ((g2320) & (g2350) & (!g2329) & (!g2371) & (g3703)) + ((g2320) & (g2350) & (!g2329) & (g2371) & (!g3703)) + ((g2320) & (g2350) & (g2329) & (g2371) & (!g3703)) + ((g2320) & (g2350) & (g2329) & (g2371) & (g3703)));
	assign g5403 = (((!g2807) & (!g2819) & (!g3822)) + ((!g2807) & (g2819) & (g3822)) + ((g2807) & (!g2819) & (g3822)) + ((g2807) & (g2819) & (!g3822)));
	assign g5404 = (((!g2178) & (!g2833) & (!g3839)) + ((!g2178) & (g2833) & (g3839)) + ((g2178) & (!g2833) & (g3839)) + ((g2178) & (g2833) & (!g3839)));
	assign g5405 = (((!g830) & (!g1914) & (!g3202) & (!g5403) & (!g5404) & (nonce[59])) + ((!g830) & (!g1914) & (!g3202) & (!g5403) & (g5404) & (nonce[59])) + ((!g830) & (!g1914) & (!g3202) & (g5403) & (!g5404) & (nonce[59])) + ((!g830) & (!g1914) & (!g3202) & (g5403) & (g5404) & (nonce[59])) + ((!g830) & (!g1914) & (g3202) & (!g5403) & (!g5404) & (nonce[59])) + ((!g830) & (!g1914) & (g3202) & (!g5403) & (g5404) & (nonce[59])) + ((!g830) & (!g1914) & (g3202) & (g5403) & (!g5404) & (nonce[59])) + ((!g830) & (!g1914) & (g3202) & (g5403) & (g5404) & (nonce[59])) + ((!g830) & (g1914) & (!g3202) & (!g5403) & (!g5404) & (nonce[59])) + ((!g830) & (g1914) & (!g3202) & (!g5403) & (g5404) & (nonce[59])) + ((!g830) & (g1914) & (!g3202) & (g5403) & (!g5404) & (nonce[59])) + ((!g830) & (g1914) & (!g3202) & (g5403) & (g5404) & (nonce[59])) + ((!g830) & (g1914) & (g3202) & (!g5403) & (!g5404) & (nonce[59])) + ((!g830) & (g1914) & (g3202) & (!g5403) & (g5404) & (nonce[59])) + ((!g830) & (g1914) & (g3202) & (g5403) & (!g5404) & (nonce[59])) + ((!g830) & (g1914) & (g3202) & (g5403) & (g5404) & (nonce[59])) + ((g830) & (!g1914) & (!g3202) & (!g5403) & (g5404) & (!nonce[59])) + ((g830) & (!g1914) & (!g3202) & (!g5403) & (g5404) & (nonce[59])) + ((g830) & (!g1914) & (!g3202) & (g5403) & (g5404) & (!nonce[59])) + ((g830) & (!g1914) & (!g3202) & (g5403) & (g5404) & (nonce[59])) + ((g830) & (!g1914) & (g3202) & (!g5403) & (!g5404) & (!nonce[59])) + ((g830) & (!g1914) & (g3202) & (!g5403) & (!g5404) & (nonce[59])) + ((g830) & (!g1914) & (g3202) & (g5403) & (!g5404) & (!nonce[59])) + ((g830) & (!g1914) & (g3202) & (g5403) & (!g5404) & (nonce[59])) + ((g830) & (g1914) & (!g3202) & (g5403) & (!g5404) & (!nonce[59])) + ((g830) & (g1914) & (!g3202) & (g5403) & (!g5404) & (nonce[59])) + ((g830) & (g1914) & (!g3202) & (g5403) & (g5404) & (!nonce[59])) + ((g830) & (g1914) & (!g3202) & (g5403) & (g5404) & (nonce[59])) + ((g830) & (g1914) & (g3202) & (!g5403) & (!g5404) & (!nonce[59])) + ((g830) & (g1914) & (g3202) & (!g5403) & (!g5404) & (nonce[59])) + ((g830) & (g1914) & (g3202) & (!g5403) & (g5404) & (!nonce[59])) + ((g830) & (g1914) & (g3202) & (!g5403) & (g5404) & (nonce[59])));
	assign g5406 = (((!g2012) & (!g2014) & (!g3596) & (!g2592) & (g2632)) + ((!g2012) & (!g2014) & (!g3596) & (g2592) & (!g2632)) + ((!g2012) & (!g2014) & (g3596) & (!g2592) & (g2632)) + ((!g2012) & (!g2014) & (g3596) & (g2592) & (g2632)) + ((!g2012) & (g2014) & (!g3596) & (!g2592) & (!g2632)) + ((!g2012) & (g2014) & (!g3596) & (g2592) & (g2632)) + ((!g2012) & (g2014) & (g3596) & (!g2592) & (!g2632)) + ((!g2012) & (g2014) & (g3596) & (g2592) & (!g2632)) + ((g2012) & (!g2014) & (!g3596) & (!g2592) & (!g2632)) + ((g2012) & (!g2014) & (!g3596) & (g2592) & (!g2632)) + ((g2012) & (!g2014) & (g3596) & (!g2592) & (g2632)) + ((g2012) & (!g2014) & (g3596) & (g2592) & (!g2632)) + ((g2012) & (g2014) & (!g3596) & (!g2592) & (g2632)) + ((g2012) & (g2014) & (!g3596) & (g2592) & (g2632)) + ((g2012) & (g2014) & (g3596) & (!g2592) & (!g2632)) + ((g2012) & (g2014) & (g3596) & (g2592) & (g2632)));
	assign g5407 = (((!g830) & (!g3207) & (!g5942) & (key[251])) + ((!g830) & (!g3207) & (g5942) & (key[251])) + ((!g830) & (g3207) & (!g5942) & (key[251])) + ((!g830) & (g3207) & (g5942) & (key[251])) + ((g830) & (!g3207) & (g5942) & (!key[251])) + ((g830) & (!g3207) & (g5942) & (key[251])) + ((g830) & (g3207) & (!g5942) & (!key[251])) + ((g830) & (g3207) & (!g5942) & (key[251])));
	assign g5408 = (((!g2181) & (!g2833) & (!g3721)) + ((!g2181) & (g2833) & (g3721)) + ((g2181) & (!g2833) & (g3721)) + ((g2181) & (g2833) & (!g3721)));
	assign g5409 = (((!g2819) & (!g2816) & (!g3738)) + ((!g2819) & (g2816) & (g3738)) + ((g2819) & (!g2816) & (g3738)) + ((g2819) & (g2816) & (!g3738)));
	assign g5410 = (((!g830) & (!g1914) & (!g3210) & (!g5408) & (!g5409) & (key[219])) + ((!g830) & (!g1914) & (!g3210) & (!g5408) & (g5409) & (key[219])) + ((!g830) & (!g1914) & (!g3210) & (g5408) & (!g5409) & (key[219])) + ((!g830) & (!g1914) & (!g3210) & (g5408) & (g5409) & (key[219])) + ((!g830) & (!g1914) & (g3210) & (!g5408) & (!g5409) & (key[219])) + ((!g830) & (!g1914) & (g3210) & (!g5408) & (g5409) & (key[219])) + ((!g830) & (!g1914) & (g3210) & (g5408) & (!g5409) & (key[219])) + ((!g830) & (!g1914) & (g3210) & (g5408) & (g5409) & (key[219])) + ((!g830) & (g1914) & (!g3210) & (!g5408) & (!g5409) & (key[219])) + ((!g830) & (g1914) & (!g3210) & (!g5408) & (g5409) & (key[219])) + ((!g830) & (g1914) & (!g3210) & (g5408) & (!g5409) & (key[219])) + ((!g830) & (g1914) & (!g3210) & (g5408) & (g5409) & (key[219])) + ((!g830) & (g1914) & (g3210) & (!g5408) & (!g5409) & (key[219])) + ((!g830) & (g1914) & (g3210) & (!g5408) & (g5409) & (key[219])) + ((!g830) & (g1914) & (g3210) & (g5408) & (!g5409) & (key[219])) + ((!g830) & (g1914) & (g3210) & (g5408) & (g5409) & (key[219])) + ((g830) & (!g1914) & (!g3210) & (!g5408) & (g5409) & (!key[219])) + ((g830) & (!g1914) & (!g3210) & (!g5408) & (g5409) & (key[219])) + ((g830) & (!g1914) & (!g3210) & (g5408) & (g5409) & (!key[219])) + ((g830) & (!g1914) & (!g3210) & (g5408) & (g5409) & (key[219])) + ((g830) & (!g1914) & (g3210) & (!g5408) & (!g5409) & (!key[219])) + ((g830) & (!g1914) & (g3210) & (!g5408) & (!g5409) & (key[219])) + ((g830) & (!g1914) & (g3210) & (g5408) & (!g5409) & (!key[219])) + ((g830) & (!g1914) & (g3210) & (g5408) & (!g5409) & (key[219])) + ((g830) & (g1914) & (!g3210) & (g5408) & (!g5409) & (!key[219])) + ((g830) & (g1914) & (!g3210) & (g5408) & (!g5409) & (key[219])) + ((g830) & (g1914) & (!g3210) & (g5408) & (g5409) & (!key[219])) + ((g830) & (g1914) & (!g3210) & (g5408) & (g5409) & (key[219])) + ((g830) & (g1914) & (g3210) & (!g5408) & (!g5409) & (!key[219])) + ((g830) & (g1914) & (g3210) & (!g5408) & (!g5409) & (key[219])) + ((g830) & (g1914) & (g3210) & (!g5408) & (g5409) & (!key[219])) + ((g830) & (g1914) & (g3210) & (!g5408) & (g5409) & (key[219])));
	assign g5411 = (((!g2317) & (g2329) & (g3850)) + ((g2317) & (!g2329) & (g3850)) + ((g2317) & (g2329) & (!g3850)) + ((g2317) & (g2329) & (g3850)));
	assign g5412 = (((!g2334) & (!g2358) & (!g2337) & (g2366) & (!g3860)) + ((!g2334) & (!g2358) & (!g2337) & (g2366) & (g3860)) + ((!g2334) & (!g2358) & (g2337) & (!g2366) & (!g3860)) + ((!g2334) & (!g2358) & (g2337) & (g2366) & (g3860)) + ((!g2334) & (g2358) & (!g2337) & (!g2366) & (!g3860)) + ((!g2334) & (g2358) & (!g2337) & (!g2366) & (g3860)) + ((!g2334) & (g2358) & (g2337) & (!g2366) & (g3860)) + ((!g2334) & (g2358) & (g2337) & (g2366) & (!g3860)) + ((g2334) & (!g2358) & (!g2337) & (!g2366) & (!g3860)) + ((g2334) & (!g2358) & (!g2337) & (g2366) & (g3860)) + ((g2334) & (!g2358) & (g2337) & (!g2366) & (!g3860)) + ((g2334) & (!g2358) & (g2337) & (!g2366) & (g3860)) + ((g2334) & (g2358) & (!g2337) & (!g2366) & (g3860)) + ((g2334) & (g2358) & (!g2337) & (g2366) & (!g3860)) + ((g2334) & (g2358) & (g2337) & (g2366) & (!g3860)) + ((g2334) & (g2358) & (g2337) & (g2366) & (g3860)));
	assign g5413 = (((!g3438) & (!g2578) & (!g2584) & (g2617) & (g2640)) + ((!g3438) & (!g2578) & (g2584) & (!g2617) & (g2640)) + ((!g3438) & (!g2578) & (g2584) & (g2617) & (!g2640)) + ((!g3438) & (!g2578) & (g2584) & (g2617) & (g2640)) + ((!g3438) & (g2578) & (!g2584) & (!g2617) & (g2640)) + ((!g3438) & (g2578) & (!g2584) & (g2617) & (!g2640)) + ((!g3438) & (g2578) & (!g2584) & (g2617) & (g2640)) + ((!g3438) & (g2578) & (g2584) & (!g2617) & (g2640)) + ((!g3438) & (g2578) & (g2584) & (g2617) & (!g2640)) + ((!g3438) & (g2578) & (g2584) & (g2617) & (g2640)) + ((g3438) & (!g2578) & (!g2584) & (g2617) & (g2640)) + ((g3438) & (!g2578) & (g2584) & (g2617) & (g2640)) + ((g3438) & (g2578) & (!g2584) & (g2617) & (g2640)) + ((g3438) & (g2578) & (g2584) & (!g2617) & (g2640)) + ((g3438) & (g2578) & (g2584) & (g2617) & (!g2640)) + ((g3438) & (g2578) & (g2584) & (g2617) & (g2640)));
	assign g5414 = (((!g5413) & (!g2665) & (g2669)) + ((!g5413) & (g2665) & (!g2669)) + ((g5413) & (!g2665) & (!g2669)) + ((g5413) & (g2665) & (g2669)));
	assign g5415 = (((!g2299) & (!g1540) & (!g3457) & (g3458)) + ((!g2299) & (!g1540) & (g3457) & (!g3458)) + ((!g2299) & (!g1540) & (g3457) & (g3458)) + ((!g2299) & (g1540) & (!g3457) & (!g3458)) + ((g2299) & (!g1540) & (!g3457) & (!g3458)) + ((g2299) & (g1540) & (!g3457) & (g3458)) + ((g2299) & (g1540) & (g3457) & (!g3458)) + ((g2299) & (g1540) & (g3457) & (g3458)));
	assign g5416 = (((!g830) & (!g1914) & (!g3222) & (!g5414) & (!g5415) & (key[124])) + ((!g830) & (!g1914) & (!g3222) & (!g5414) & (g5415) & (key[124])) + ((!g830) & (!g1914) & (!g3222) & (g5414) & (!g5415) & (key[124])) + ((!g830) & (!g1914) & (!g3222) & (g5414) & (g5415) & (key[124])) + ((!g830) & (!g1914) & (g3222) & (!g5414) & (!g5415) & (key[124])) + ((!g830) & (!g1914) & (g3222) & (!g5414) & (g5415) & (key[124])) + ((!g830) & (!g1914) & (g3222) & (g5414) & (!g5415) & (key[124])) + ((!g830) & (!g1914) & (g3222) & (g5414) & (g5415) & (key[124])) + ((!g830) & (g1914) & (!g3222) & (!g5414) & (!g5415) & (key[124])) + ((!g830) & (g1914) & (!g3222) & (!g5414) & (g5415) & (key[124])) + ((!g830) & (g1914) & (!g3222) & (g5414) & (!g5415) & (key[124])) + ((!g830) & (g1914) & (!g3222) & (g5414) & (g5415) & (key[124])) + ((!g830) & (g1914) & (g3222) & (!g5414) & (!g5415) & (key[124])) + ((!g830) & (g1914) & (g3222) & (!g5414) & (g5415) & (key[124])) + ((!g830) & (g1914) & (g3222) & (g5414) & (!g5415) & (key[124])) + ((!g830) & (g1914) & (g3222) & (g5414) & (g5415) & (key[124])) + ((g830) & (!g1914) & (!g3222) & (!g5414) & (g5415) & (!key[124])) + ((g830) & (!g1914) & (!g3222) & (!g5414) & (g5415) & (key[124])) + ((g830) & (!g1914) & (!g3222) & (g5414) & (g5415) & (!key[124])) + ((g830) & (!g1914) & (!g3222) & (g5414) & (g5415) & (key[124])) + ((g830) & (!g1914) & (g3222) & (!g5414) & (!g5415) & (!key[124])) + ((g830) & (!g1914) & (g3222) & (!g5414) & (!g5415) & (key[124])) + ((g830) & (!g1914) & (g3222) & (g5414) & (!g5415) & (!key[124])) + ((g830) & (!g1914) & (g3222) & (g5414) & (!g5415) & (key[124])) + ((g830) & (g1914) & (!g3222) & (g5414) & (!g5415) & (!key[124])) + ((g830) & (g1914) & (!g3222) & (g5414) & (!g5415) & (key[124])) + ((g830) & (g1914) & (!g3222) & (g5414) & (g5415) & (!key[124])) + ((g830) & (g1914) & (!g3222) & (g5414) & (g5415) & (key[124])) + ((g830) & (g1914) & (g3222) & (!g5414) & (!g5415) & (!key[124])) + ((g830) & (g1914) & (g3222) & (!g5414) & (!g5415) & (key[124])) + ((g830) & (g1914) & (g3222) & (!g5414) & (g5415) & (!key[124])) + ((g830) & (g1914) & (g3222) & (!g5414) & (g5415) & (key[124])));
	assign g5417 = (((!g1998) & (!g2001) & (!g5389) & (!g2356) & (g2402)) + ((!g1998) & (!g2001) & (!g5389) & (g2356) & (g2402)) + ((!g1998) & (!g2001) & (g5389) & (!g2356) & (g2402)) + ((!g1998) & (!g2001) & (g5389) & (g2356) & (!g2402)) + ((!g1998) & (g2001) & (!g5389) & (!g2356) & (!g2402)) + ((!g1998) & (g2001) & (!g5389) & (g2356) & (!g2402)) + ((!g1998) & (g2001) & (g5389) & (!g2356) & (!g2402)) + ((!g1998) & (g2001) & (g5389) & (g2356) & (g2402)) + ((g1998) & (!g2001) & (!g5389) & (!g2356) & (g2402)) + ((g1998) & (!g2001) & (!g5389) & (g2356) & (!g2402)) + ((g1998) & (!g2001) & (g5389) & (!g2356) & (!g2402)) + ((g1998) & (!g2001) & (g5389) & (g2356) & (!g2402)) + ((g1998) & (g2001) & (!g5389) & (!g2356) & (!g2402)) + ((g1998) & (g2001) & (!g5389) & (g2356) & (g2402)) + ((g1998) & (g2001) & (g5389) & (!g2356) & (g2402)) + ((g1998) & (g2001) & (g5389) & (g2356) & (g2402)));
	assign g5418 = (((!g2950) & (!g3568) & (!g3569) & (g2962)) + ((!g2950) & (!g3568) & (g3569) & (!g2962)) + ((!g2950) & (g3568) & (!g3569) & (!g2962)) + ((!g2950) & (g3568) & (g3569) & (!g2962)) + ((g2950) & (!g3568) & (!g3569) & (!g2962)) + ((g2950) & (!g3568) & (g3569) & (g2962)) + ((g2950) & (g3568) & (!g3569) & (g2962)) + ((g2950) & (g3568) & (g3569) & (g2962)));
	assign g5419 = (((!g1972) & (!g1975) & (g2589) & (g2620) & (!g3580)) + ((!g1972) & (g1975) & (!g2589) & (g2620) & (!g3580)) + ((!g1972) & (g1975) & (!g2589) & (g2620) & (g3580)) + ((!g1972) & (g1975) & (g2589) & (!g2620) & (!g3580)) + ((!g1972) & (g1975) & (g2589) & (g2620) & (!g3580)) + ((!g1972) & (g1975) & (g2589) & (g2620) & (g3580)) + ((g1972) & (!g1975) & (!g2589) & (g2620) & (!g3580)) + ((g1972) & (!g1975) & (g2589) & (g2620) & (!g3580)) + ((g1972) & (!g1975) & (g2589) & (g2620) & (g3580)) + ((g1972) & (g1975) & (!g2589) & (!g2620) & (!g3580)) + ((g1972) & (g1975) & (!g2589) & (g2620) & (!g3580)) + ((g1972) & (g1975) & (!g2589) & (g2620) & (g3580)) + ((g1972) & (g1975) & (g2589) & (!g2620) & (!g3580)) + ((g1972) & (g1975) & (g2589) & (!g2620) & (g3580)) + ((g1972) & (g1975) & (g2589) & (g2620) & (!g3580)) + ((g1972) & (g1975) & (g2589) & (g2620) & (g3580)));
	assign g5420 = (((!g2047) & (!g2672) & (g5419)) + ((!g2047) & (g2672) & (!g5419)) + ((g2047) & (!g2672) & (!g5419)) + ((g2047) & (g2672) & (g5419)));
	assign g5421 = (((!g830) & (!g1914) & (!g3240) & (!g5418) & (!g5420) & (nonce[28])) + ((!g830) & (!g1914) & (!g3240) & (!g5418) & (g5420) & (nonce[28])) + ((!g830) & (!g1914) & (!g3240) & (g5418) & (!g5420) & (nonce[28])) + ((!g830) & (!g1914) & (!g3240) & (g5418) & (g5420) & (nonce[28])) + ((!g830) & (!g1914) & (g3240) & (!g5418) & (!g5420) & (nonce[28])) + ((!g830) & (!g1914) & (g3240) & (!g5418) & (g5420) & (nonce[28])) + ((!g830) & (!g1914) & (g3240) & (g5418) & (!g5420) & (nonce[28])) + ((!g830) & (!g1914) & (g3240) & (g5418) & (g5420) & (nonce[28])) + ((!g830) & (g1914) & (!g3240) & (!g5418) & (!g5420) & (nonce[28])) + ((!g830) & (g1914) & (!g3240) & (!g5418) & (g5420) & (nonce[28])) + ((!g830) & (g1914) & (!g3240) & (g5418) & (!g5420) & (nonce[28])) + ((!g830) & (g1914) & (!g3240) & (g5418) & (g5420) & (nonce[28])) + ((!g830) & (g1914) & (g3240) & (!g5418) & (!g5420) & (nonce[28])) + ((!g830) & (g1914) & (g3240) & (!g5418) & (g5420) & (nonce[28])) + ((!g830) & (g1914) & (g3240) & (g5418) & (!g5420) & (nonce[28])) + ((!g830) & (g1914) & (g3240) & (g5418) & (g5420) & (nonce[28])) + ((g830) & (!g1914) & (!g3240) & (!g5418) & (g5420) & (!nonce[28])) + ((g830) & (!g1914) & (!g3240) & (!g5418) & (g5420) & (nonce[28])) + ((g830) & (!g1914) & (!g3240) & (g5418) & (g5420) & (!nonce[28])) + ((g830) & (!g1914) & (!g3240) & (g5418) & (g5420) & (nonce[28])) + ((g830) & (!g1914) & (g3240) & (!g5418) & (!g5420) & (!nonce[28])) + ((g830) & (!g1914) & (g3240) & (!g5418) & (!g5420) & (nonce[28])) + ((g830) & (!g1914) & (g3240) & (g5418) & (!g5420) & (!nonce[28])) + ((g830) & (!g1914) & (g3240) & (g5418) & (!g5420) & (nonce[28])) + ((g830) & (g1914) & (!g3240) & (g5418) & (!g5420) & (!nonce[28])) + ((g830) & (g1914) & (!g3240) & (g5418) & (!g5420) & (nonce[28])) + ((g830) & (g1914) & (!g3240) & (g5418) & (g5420) & (!nonce[28])) + ((g830) & (g1914) & (!g3240) & (g5418) & (g5420) & (nonce[28])) + ((g830) & (g1914) & (g3240) & (!g5418) & (!g5420) & (!nonce[28])) + ((g830) & (g1914) & (g3240) & (!g5418) & (!g5420) & (nonce[28])) + ((g830) & (g1914) & (g3240) & (!g5418) & (g5420) & (!nonce[28])) + ((g830) & (g1914) & (g3240) & (!g5418) & (g5420) & (nonce[28])));
	assign g5422 = (((!g2012) & (!g2014) & (!g3596) & (g2592) & (g2632)) + ((!g2012) & (g2014) & (!g3596) & (!g2592) & (g2632)) + ((!g2012) & (g2014) & (!g3596) & (g2592) & (!g2632)) + ((!g2012) & (g2014) & (!g3596) & (g2592) & (g2632)) + ((!g2012) & (g2014) & (g3596) & (!g2592) & (g2632)) + ((!g2012) & (g2014) & (g3596) & (g2592) & (g2632)) + ((g2012) & (!g2014) & (!g3596) & (!g2592) & (g2632)) + ((g2012) & (!g2014) & (!g3596) & (g2592) & (g2632)) + ((g2012) & (!g2014) & (g3596) & (g2592) & (g2632)) + ((g2012) & (g2014) & (!g3596) & (!g2592) & (!g2632)) + ((g2012) & (g2014) & (!g3596) & (!g2592) & (g2632)) + ((g2012) & (g2014) & (!g3596) & (g2592) & (!g2632)) + ((g2012) & (g2014) & (!g3596) & (g2592) & (g2632)) + ((g2012) & (g2014) & (g3596) & (!g2592) & (g2632)) + ((g2012) & (g2014) & (g3596) & (g2592) & (!g2632)) + ((g2012) & (g2014) & (g3596) & (g2592) & (g2632)));
	assign g5423 = (((!g2052) & (!g5422) & (g2674)) + ((!g2052) & (g5422) & (!g2674)) + ((g2052) & (!g5422) & (!g2674)) + ((g2052) & (g5422) & (g2674)));
	assign g5424 = (((!g2932) & (!g3615) & (!g3616) & (g2956)) + ((!g2932) & (!g3615) & (g3616) & (!g2956)) + ((!g2932) & (g3615) & (!g3616) & (!g2956)) + ((!g2932) & (g3615) & (g3616) & (!g2956)) + ((g2932) & (!g3615) & (!g3616) & (!g2956)) + ((g2932) & (!g3615) & (g3616) & (g2956)) + ((g2932) & (g3615) & (!g3616) & (g2956)) + ((g2932) & (g3615) & (g3616) & (g2956)));
	assign g5425 = (((!g830) & (!g1914) & (!g3245) & (!g5423) & (!g5424) & (key[252])) + ((!g830) & (!g1914) & (!g3245) & (!g5423) & (g5424) & (key[252])) + ((!g830) & (!g1914) & (!g3245) & (g5423) & (!g5424) & (key[252])) + ((!g830) & (!g1914) & (!g3245) & (g5423) & (g5424) & (key[252])) + ((!g830) & (!g1914) & (g3245) & (!g5423) & (!g5424) & (key[252])) + ((!g830) & (!g1914) & (g3245) & (!g5423) & (g5424) & (key[252])) + ((!g830) & (!g1914) & (g3245) & (g5423) & (!g5424) & (key[252])) + ((!g830) & (!g1914) & (g3245) & (g5423) & (g5424) & (key[252])) + ((!g830) & (g1914) & (!g3245) & (!g5423) & (!g5424) & (key[252])) + ((!g830) & (g1914) & (!g3245) & (!g5423) & (g5424) & (key[252])) + ((!g830) & (g1914) & (!g3245) & (g5423) & (!g5424) & (key[252])) + ((!g830) & (g1914) & (!g3245) & (g5423) & (g5424) & (key[252])) + ((!g830) & (g1914) & (g3245) & (!g5423) & (!g5424) & (key[252])) + ((!g830) & (g1914) & (g3245) & (!g5423) & (g5424) & (key[252])) + ((!g830) & (g1914) & (g3245) & (g5423) & (!g5424) & (key[252])) + ((!g830) & (g1914) & (g3245) & (g5423) & (g5424) & (key[252])) + ((g830) & (!g1914) & (!g3245) & (!g5423) & (g5424) & (!key[252])) + ((g830) & (!g1914) & (!g3245) & (!g5423) & (g5424) & (key[252])) + ((g830) & (!g1914) & (!g3245) & (g5423) & (g5424) & (!key[252])) + ((g830) & (!g1914) & (!g3245) & (g5423) & (g5424) & (key[252])) + ((g830) & (!g1914) & (g3245) & (!g5423) & (!g5424) & (!key[252])) + ((g830) & (!g1914) & (g3245) & (!g5423) & (!g5424) & (key[252])) + ((g830) & (!g1914) & (g3245) & (g5423) & (!g5424) & (!key[252])) + ((g830) & (!g1914) & (g3245) & (g5423) & (!g5424) & (key[252])) + ((g830) & (g1914) & (!g3245) & (g5423) & (!g5424) & (!key[252])) + ((g830) & (g1914) & (!g3245) & (g5423) & (!g5424) & (key[252])) + ((g830) & (g1914) & (!g3245) & (g5423) & (g5424) & (!key[252])) + ((g830) & (g1914) & (!g3245) & (g5423) & (g5424) & (key[252])) + ((g830) & (g1914) & (g3245) & (!g5423) & (!g5424) & (!key[252])) + ((g830) & (g1914) & (g3245) & (!g5423) & (!g5424) & (key[252])) + ((g830) & (g1914) & (g3245) & (!g5423) & (g5424) & (!key[252])) + ((g830) & (g1914) & (g3245) & (!g5423) & (g5424) & (key[252])));
	assign g5426 = (((!g2296) & (!g1540) & (!g3634) & (g3635)) + ((!g2296) & (!g1540) & (g3634) & (!g3635)) + ((!g2296) & (!g1540) & (g3634) & (g3635)) + ((!g2296) & (g1540) & (!g3634) & (!g3635)) + ((g2296) & (!g1540) & (!g3634) & (!g3635)) + ((g2296) & (g1540) & (!g3634) & (g3635)) + ((g2296) & (g1540) & (g3634) & (!g3635)) + ((g2296) & (g1540) & (g3634) & (g3635)));
	assign g5427 = (((!g2569) & (!g2626) & (g2592) & (g2632) & (!g3646)) + ((!g2569) & (g2626) & (!g2592) & (g2632) & (!g3646)) + ((!g2569) & (g2626) & (!g2592) & (g2632) & (g3646)) + ((!g2569) & (g2626) & (g2592) & (!g2632) & (!g3646)) + ((!g2569) & (g2626) & (g2592) & (g2632) & (!g3646)) + ((!g2569) & (g2626) & (g2592) & (g2632) & (g3646)) + ((g2569) & (!g2626) & (!g2592) & (g2632) & (!g3646)) + ((g2569) & (!g2626) & (g2592) & (g2632) & (!g3646)) + ((g2569) & (!g2626) & (g2592) & (g2632) & (g3646)) + ((g2569) & (g2626) & (!g2592) & (!g2632) & (!g3646)) + ((g2569) & (g2626) & (!g2592) & (g2632) & (!g3646)) + ((g2569) & (g2626) & (!g2592) & (g2632) & (g3646)) + ((g2569) & (g2626) & (g2592) & (!g2632) & (!g3646)) + ((g2569) & (g2626) & (g2592) & (!g2632) & (g3646)) + ((g2569) & (g2626) & (g2592) & (g2632) & (!g3646)) + ((g2569) & (g2626) & (g2592) & (g2632) & (g3646)));
	assign g5428 = (((!g2674) & (!g5427) & (g2659)) + ((!g2674) & (g5427) & (!g2659)) + ((g2674) & (!g5427) & (!g2659)) + ((g2674) & (g5427) & (g2659)));
	assign g5429 = (((!g830) & (!g1914) & (!g3250) & (!g5426) & (!g5428) & (key[28])) + ((!g830) & (!g1914) & (!g3250) & (!g5426) & (g5428) & (key[28])) + ((!g830) & (!g1914) & (!g3250) & (g5426) & (!g5428) & (key[28])) + ((!g830) & (!g1914) & (!g3250) & (g5426) & (g5428) & (key[28])) + ((!g830) & (!g1914) & (g3250) & (!g5426) & (!g5428) & (key[28])) + ((!g830) & (!g1914) & (g3250) & (!g5426) & (g5428) & (key[28])) + ((!g830) & (!g1914) & (g3250) & (g5426) & (!g5428) & (key[28])) + ((!g830) & (!g1914) & (g3250) & (g5426) & (g5428) & (key[28])) + ((!g830) & (g1914) & (!g3250) & (!g5426) & (!g5428) & (key[28])) + ((!g830) & (g1914) & (!g3250) & (!g5426) & (g5428) & (key[28])) + ((!g830) & (g1914) & (!g3250) & (g5426) & (!g5428) & (key[28])) + ((!g830) & (g1914) & (!g3250) & (g5426) & (g5428) & (key[28])) + ((!g830) & (g1914) & (g3250) & (!g5426) & (!g5428) & (key[28])) + ((!g830) & (g1914) & (g3250) & (!g5426) & (g5428) & (key[28])) + ((!g830) & (g1914) & (g3250) & (g5426) & (!g5428) & (key[28])) + ((!g830) & (g1914) & (g3250) & (g5426) & (g5428) & (key[28])) + ((g830) & (!g1914) & (!g3250) & (!g5426) & (g5428) & (!key[28])) + ((g830) & (!g1914) & (!g3250) & (!g5426) & (g5428) & (key[28])) + ((g830) & (!g1914) & (!g3250) & (g5426) & (g5428) & (!key[28])) + ((g830) & (!g1914) & (!g3250) & (g5426) & (g5428) & (key[28])) + ((g830) & (!g1914) & (g3250) & (!g5426) & (!g5428) & (!key[28])) + ((g830) & (!g1914) & (g3250) & (!g5426) & (!g5428) & (key[28])) + ((g830) & (!g1914) & (g3250) & (g5426) & (!g5428) & (!key[28])) + ((g830) & (!g1914) & (g3250) & (g5426) & (!g5428) & (key[28])) + ((g830) & (g1914) & (!g3250) & (g5426) & (!g5428) & (!key[28])) + ((g830) & (g1914) & (!g3250) & (g5426) & (!g5428) & (key[28])) + ((g830) & (g1914) & (!g3250) & (g5426) & (g5428) & (!key[28])) + ((g830) & (g1914) & (!g3250) & (g5426) & (g5428) & (key[28])) + ((g830) & (g1914) & (g3250) & (!g5426) & (!g5428) & (!key[28])) + ((g830) & (g1914) & (g3250) & (!g5426) & (!g5428) & (key[28])) + ((g830) & (g1914) & (g3250) & (!g5426) & (g5428) & (!key[28])) + ((g830) & (g1914) & (g3250) & (!g5426) & (g5428) & (key[28])));
	assign g5430 = (((!g2011) & (!g2013) & (g2572) & (g2637) & (!g3662)) + ((!g2011) & (g2013) & (!g2572) & (g2637) & (!g3662)) + ((!g2011) & (g2013) & (!g2572) & (g2637) & (g3662)) + ((!g2011) & (g2013) & (g2572) & (!g2637) & (!g3662)) + ((!g2011) & (g2013) & (g2572) & (g2637) & (!g3662)) + ((!g2011) & (g2013) & (g2572) & (g2637) & (g3662)) + ((g2011) & (!g2013) & (!g2572) & (g2637) & (!g3662)) + ((g2011) & (!g2013) & (g2572) & (g2637) & (!g3662)) + ((g2011) & (!g2013) & (g2572) & (g2637) & (g3662)) + ((g2011) & (g2013) & (!g2572) & (!g2637) & (!g3662)) + ((g2011) & (g2013) & (!g2572) & (g2637) & (!g3662)) + ((g2011) & (g2013) & (!g2572) & (g2637) & (g3662)) + ((g2011) & (g2013) & (g2572) & (!g2637) & (!g3662)) + ((g2011) & (g2013) & (g2572) & (!g2637) & (g3662)) + ((g2011) & (g2013) & (g2572) & (g2637) & (!g3662)) + ((g2011) & (g2013) & (g2572) & (g2637) & (g3662)));
	assign g5431 = (((!g2051) & (!g2661) & (g5430)) + ((!g2051) & (g2661) & (!g5430)) + ((g2051) & (!g2661) & (!g5430)) + ((g2051) & (g2661) & (g5430)));
	assign g5432 = (((!g3682) & (!g3683)));
	assign g5433 = (((!g2916) & (!g2962) & (!g5432)) + ((!g2916) & (g2962) & (g5432)) + ((g2916) & (!g2962) & (g5432)) + ((g2916) & (g2962) & (!g5432)));
	assign g8336 = (((!g5560) & (g5643) & (!g5434)) + ((!g5560) & (g5643) & (g5434)) + ((g5560) & (!g5643) & (g5434)) + ((g5560) & (g5643) & (g5434)));
	assign g5435 = (((!g830) & (!g1914) & (!g3255) & (!g5431) & (!g5433) & (g5434)) + ((!g830) & (!g1914) & (!g3255) & (!g5431) & (g5433) & (g5434)) + ((!g830) & (!g1914) & (!g3255) & (g5431) & (!g5433) & (g5434)) + ((!g830) & (!g1914) & (!g3255) & (g5431) & (g5433) & (g5434)) + ((!g830) & (!g1914) & (g3255) & (!g5431) & (!g5433) & (g5434)) + ((!g830) & (!g1914) & (g3255) & (!g5431) & (g5433) & (g5434)) + ((!g830) & (!g1914) & (g3255) & (g5431) & (!g5433) & (g5434)) + ((!g830) & (!g1914) & (g3255) & (g5431) & (g5433) & (g5434)) + ((!g830) & (g1914) & (!g3255) & (!g5431) & (!g5433) & (g5434)) + ((!g830) & (g1914) & (!g3255) & (!g5431) & (g5433) & (g5434)) + ((!g830) & (g1914) & (!g3255) & (g5431) & (!g5433) & (g5434)) + ((!g830) & (g1914) & (!g3255) & (g5431) & (g5433) & (g5434)) + ((!g830) & (g1914) & (g3255) & (!g5431) & (!g5433) & (g5434)) + ((!g830) & (g1914) & (g3255) & (!g5431) & (g5433) & (g5434)) + ((!g830) & (g1914) & (g3255) & (g5431) & (!g5433) & (g5434)) + ((!g830) & (g1914) & (g3255) & (g5431) & (g5433) & (g5434)) + ((g830) & (!g1914) & (!g3255) & (!g5431) & (g5433) & (!g5434)) + ((g830) & (!g1914) & (!g3255) & (!g5431) & (g5433) & (g5434)) + ((g830) & (!g1914) & (!g3255) & (g5431) & (g5433) & (!g5434)) + ((g830) & (!g1914) & (!g3255) & (g5431) & (g5433) & (g5434)) + ((g830) & (!g1914) & (g3255) & (!g5431) & (!g5433) & (!g5434)) + ((g830) & (!g1914) & (g3255) & (!g5431) & (!g5433) & (g5434)) + ((g830) & (!g1914) & (g3255) & (g5431) & (!g5433) & (!g5434)) + ((g830) & (!g1914) & (g3255) & (g5431) & (!g5433) & (g5434)) + ((g830) & (g1914) & (!g3255) & (g5431) & (!g5433) & (!g5434)) + ((g830) & (g1914) & (!g3255) & (g5431) & (!g5433) & (g5434)) + ((g830) & (g1914) & (!g3255) & (g5431) & (g5433) & (!g5434)) + ((g830) & (g1914) & (!g3255) & (g5431) & (g5433) & (g5434)) + ((g830) & (g1914) & (g3255) & (!g5431) & (!g5433) & (!g5434)) + ((g830) & (g1914) & (g3255) & (!g5431) & (!g5433) & (g5434)) + ((g830) & (g1914) & (g3255) & (!g5431) & (g5433) & (!g5434)) + ((g830) & (g1914) & (g3255) & (!g5431) & (g5433) & (g5434)));
	assign g5436 = (((!g2360) & (!g2383) & (!g2366) & (g2416) & (!g5401)) + ((!g2360) & (!g2383) & (!g2366) & (g2416) & (g5401)) + ((!g2360) & (!g2383) & (g2366) & (!g2416) & (g5401)) + ((!g2360) & (!g2383) & (g2366) & (g2416) & (!g5401)) + ((!g2360) & (g2383) & (!g2366) & (!g2416) & (!g5401)) + ((!g2360) & (g2383) & (!g2366) & (!g2416) & (g5401)) + ((!g2360) & (g2383) & (g2366) & (!g2416) & (!g5401)) + ((!g2360) & (g2383) & (g2366) & (g2416) & (g5401)) + ((g2360) & (!g2383) & (!g2366) & (!g2416) & (g5401)) + ((g2360) & (!g2383) & (!g2366) & (g2416) & (!g5401)) + ((g2360) & (!g2383) & (g2366) & (!g2416) & (!g5401)) + ((g2360) & (!g2383) & (g2366) & (!g2416) & (g5401)) + ((g2360) & (g2383) & (!g2366) & (!g2416) & (!g5401)) + ((g2360) & (g2383) & (!g2366) & (g2416) & (g5401)) + ((g2360) & (g2383) & (g2366) & (g2416) & (!g5401)) + ((g2360) & (g2383) & (g2366) & (g2416) & (g5401)));
	assign g5437 = (((!g2181) & (g2833) & (!g3721)) + ((g2181) & (!g2833) & (!g3721)) + ((g2181) & (g2833) & (!g3721)) + ((g2181) & (g2833) & (g3721)));
	assign g5438 = (((g1914) & (!g2213) & (!g2874) & (g5437)) + ((g1914) & (!g2213) & (g2874) & (!g5437)) + ((g1914) & (g2213) & (!g2874) & (!g5437)) + ((g1914) & (g2213) & (g2874) & (g5437)));
	assign g5439 = (((!g2819) & (g2816) & (!g3738)) + ((g2819) & (!g2816) & (!g3738)) + ((g2819) & (g2816) & (!g3738)) + ((g2819) & (g2816) & (g3738)));
	assign g5440 = (((!g1914) & (!g2860) & (!g2848) & (g5439)) + ((!g1914) & (!g2860) & (g2848) & (!g5439)) + ((!g1914) & (g2860) & (!g2848) & (!g5439)) + ((!g1914) & (g2860) & (g2848) & (g5439)));
	assign g5441 = (((!g830) & (!g3265) & (!g5438) & (!g5440) & (key[220])) + ((!g830) & (!g3265) & (!g5438) & (g5440) & (key[220])) + ((!g830) & (!g3265) & (g5438) & (!g5440) & (key[220])) + ((!g830) & (!g3265) & (g5438) & (g5440) & (key[220])) + ((!g830) & (g3265) & (!g5438) & (!g5440) & (key[220])) + ((!g830) & (g3265) & (!g5438) & (g5440) & (key[220])) + ((!g830) & (g3265) & (g5438) & (!g5440) & (key[220])) + ((!g830) & (g3265) & (g5438) & (g5440) & (key[220])) + ((g830) & (!g3265) & (!g5438) & (g5440) & (!key[220])) + ((g830) & (!g3265) & (!g5438) & (g5440) & (key[220])) + ((g830) & (!g3265) & (g5438) & (!g5440) & (!key[220])) + ((g830) & (!g3265) & (g5438) & (!g5440) & (key[220])) + ((g830) & (!g3265) & (g5438) & (g5440) & (!key[220])) + ((g830) & (!g3265) & (g5438) & (g5440) & (key[220])) + ((g830) & (g3265) & (!g5438) & (!g5440) & (!key[220])) + ((g830) & (g3265) & (!g5438) & (!g5440) & (key[220])));
	assign g5442 = (((!g2932) & (!g2938) & (!g3791) & (g3792)) + ((!g2932) & (!g2938) & (g3791) & (!g3792)) + ((!g2932) & (!g2938) & (g3791) & (g3792)) + ((!g2932) & (g2938) & (!g3791) & (!g3792)) + ((g2932) & (!g2938) & (!g3791) & (!g3792)) + ((g2932) & (g2938) & (!g3791) & (g3792)) + ((g2932) & (g2938) & (g3791) & (!g3792)) + ((g2932) & (g2938) & (g3791) & (g3792)));
	assign g5443 = (((!g1973) & (!g1976) & (g2584) & (g2640) & (!g3803)) + ((!g1973) & (g1976) & (!g2584) & (g2640) & (!g3803)) + ((!g1973) & (g1976) & (!g2584) & (g2640) & (g3803)) + ((!g1973) & (g1976) & (g2584) & (!g2640) & (!g3803)) + ((!g1973) & (g1976) & (g2584) & (g2640) & (!g3803)) + ((!g1973) & (g1976) & (g2584) & (g2640) & (g3803)) + ((g1973) & (!g1976) & (!g2584) & (g2640) & (!g3803)) + ((g1973) & (!g1976) & (g2584) & (g2640) & (!g3803)) + ((g1973) & (!g1976) & (g2584) & (g2640) & (g3803)) + ((g1973) & (g1976) & (!g2584) & (!g2640) & (!g3803)) + ((g1973) & (g1976) & (!g2584) & (g2640) & (!g3803)) + ((g1973) & (g1976) & (!g2584) & (g2640) & (g3803)) + ((g1973) & (g1976) & (g2584) & (!g2640) & (!g3803)) + ((g1973) & (g1976) & (g2584) & (!g2640) & (g3803)) + ((g1973) & (g1976) & (g2584) & (g2640) & (!g3803)) + ((g1973) & (g1976) & (g2584) & (g2640) & (g3803)));
	assign g5444 = (((!g2048) & (!g2669) & (g5443)) + ((!g2048) & (g2669) & (!g5443)) + ((g2048) & (!g2669) & (!g5443)) + ((g2048) & (g2669) & (g5443)));
	assign g5445 = (((!g830) & (!g1914) & (!g3274) & (!g5442) & (!g5444) & (key[156])) + ((!g830) & (!g1914) & (!g3274) & (!g5442) & (g5444) & (key[156])) + ((!g830) & (!g1914) & (!g3274) & (g5442) & (!g5444) & (key[156])) + ((!g830) & (!g1914) & (!g3274) & (g5442) & (g5444) & (key[156])) + ((!g830) & (!g1914) & (g3274) & (!g5442) & (!g5444) & (key[156])) + ((!g830) & (!g1914) & (g3274) & (!g5442) & (g5444) & (key[156])) + ((!g830) & (!g1914) & (g3274) & (g5442) & (!g5444) & (key[156])) + ((!g830) & (!g1914) & (g3274) & (g5442) & (g5444) & (key[156])) + ((!g830) & (g1914) & (!g3274) & (!g5442) & (!g5444) & (key[156])) + ((!g830) & (g1914) & (!g3274) & (!g5442) & (g5444) & (key[156])) + ((!g830) & (g1914) & (!g3274) & (g5442) & (!g5444) & (key[156])) + ((!g830) & (g1914) & (!g3274) & (g5442) & (g5444) & (key[156])) + ((!g830) & (g1914) & (g3274) & (!g5442) & (!g5444) & (key[156])) + ((!g830) & (g1914) & (g3274) & (!g5442) & (g5444) & (key[156])) + ((!g830) & (g1914) & (g3274) & (g5442) & (!g5444) & (key[156])) + ((!g830) & (g1914) & (g3274) & (g5442) & (g5444) & (key[156])) + ((g830) & (!g1914) & (!g3274) & (!g5442) & (g5444) & (!key[156])) + ((g830) & (!g1914) & (!g3274) & (!g5442) & (g5444) & (key[156])) + ((g830) & (!g1914) & (!g3274) & (g5442) & (g5444) & (!key[156])) + ((g830) & (!g1914) & (!g3274) & (g5442) & (g5444) & (key[156])) + ((g830) & (!g1914) & (g3274) & (!g5442) & (!g5444) & (!key[156])) + ((g830) & (!g1914) & (g3274) & (!g5442) & (!g5444) & (key[156])) + ((g830) & (!g1914) & (g3274) & (g5442) & (!g5444) & (!key[156])) + ((g830) & (!g1914) & (g3274) & (g5442) & (!g5444) & (key[156])) + ((g830) & (g1914) & (!g3274) & (g5442) & (!g5444) & (!key[156])) + ((g830) & (g1914) & (!g3274) & (g5442) & (!g5444) & (key[156])) + ((g830) & (g1914) & (!g3274) & (g5442) & (g5444) & (!key[156])) + ((g830) & (g1914) & (!g3274) & (g5442) & (g5444) & (key[156])) + ((g830) & (g1914) & (g3274) & (!g5442) & (!g5444) & (!key[156])) + ((g830) & (g1914) & (g3274) & (!g5442) & (!g5444) & (key[156])) + ((g830) & (g1914) & (g3274) & (!g5442) & (g5444) & (!key[156])) + ((g830) & (g1914) & (g3274) & (!g5442) & (g5444) & (key[156])));
	assign g5446 = (((!g2807) & (g2819) & (!g3822)) + ((g2807) & (!g2819) & (!g3822)) + ((g2807) & (g2819) & (!g3822)) + ((g2807) & (g2819) & (g3822)));
	assign g5447 = (((g1914) & (!g2857) & (!g2860) & (g5446)) + ((g1914) & (!g2857) & (g2860) & (!g5446)) + ((g1914) & (g2857) & (!g2860) & (!g5446)) + ((g1914) & (g2857) & (g2860) & (g5446)));
	assign g5448 = (((!g2178) & (g2833) & (!g3839)) + ((g2178) & (!g2833) & (!g3839)) + ((g2178) & (g2833) & (!g3839)) + ((g2178) & (g2833) & (g3839)));
	assign g5449 = (((!g1914) & (!g2211) & (!g2874) & (g5448)) + ((!g1914) & (!g2211) & (g2874) & (!g5448)) + ((!g1914) & (g2211) & (!g2874) & (!g5448)) + ((!g1914) & (g2211) & (g2874) & (g5448)));
	assign g5450 = (((!g830) & (!g3279) & (!g5447) & (!g5449) & (nonce[60])) + ((!g830) & (!g3279) & (!g5447) & (g5449) & (nonce[60])) + ((!g830) & (!g3279) & (g5447) & (!g5449) & (nonce[60])) + ((!g830) & (!g3279) & (g5447) & (g5449) & (nonce[60])) + ((!g830) & (g3279) & (!g5447) & (!g5449) & (nonce[60])) + ((!g830) & (g3279) & (!g5447) & (g5449) & (nonce[60])) + ((!g830) & (g3279) & (g5447) & (!g5449) & (nonce[60])) + ((!g830) & (g3279) & (g5447) & (g5449) & (nonce[60])) + ((g830) & (!g3279) & (!g5447) & (g5449) & (!nonce[60])) + ((g830) & (!g3279) & (!g5447) & (g5449) & (nonce[60])) + ((g830) & (!g3279) & (g5447) & (!g5449) & (!nonce[60])) + ((g830) & (!g3279) & (g5447) & (!g5449) & (nonce[60])) + ((g830) & (!g3279) & (g5447) & (g5449) & (!nonce[60])) + ((g830) & (!g3279) & (g5447) & (g5449) & (nonce[60])) + ((g830) & (g3279) & (!g5447) & (!g5449) & (!nonce[60])) + ((g830) & (g3279) & (!g5447) & (!g5449) & (nonce[60])));
	assign g5451 = (((!g2369) & (!g2396) & (!g2371) & (g2408) & (!g5411)) + ((!g2369) & (!g2396) & (!g2371) & (g2408) & (g5411)) + ((!g2369) & (!g2396) & (g2371) & (!g2408) & (g5411)) + ((!g2369) & (!g2396) & (g2371) & (g2408) & (!g5411)) + ((!g2369) & (g2396) & (!g2371) & (!g2408) & (!g5411)) + ((!g2369) & (g2396) & (!g2371) & (!g2408) & (g5411)) + ((!g2369) & (g2396) & (g2371) & (!g2408) & (!g5411)) + ((!g2369) & (g2396) & (g2371) & (g2408) & (g5411)) + ((g2369) & (!g2396) & (!g2371) & (!g2408) & (g5411)) + ((g2369) & (!g2396) & (!g2371) & (g2408) & (!g5411)) + ((g2369) & (!g2396) & (g2371) & (!g2408) & (!g5411)) + ((g2369) & (!g2396) & (g2371) & (!g2408) & (g5411)) + ((g2369) & (g2396) & (!g2371) & (!g2408) & (!g5411)) + ((g2369) & (g2396) & (!g2371) & (g2408) & (g5411)) + ((g2369) & (g2396) & (g2371) & (g2408) & (!g5411)) + ((g2369) & (g2396) & (g2371) & (g2408) & (g5411)));
	assign g5452 = (((!g2296) & (g1540) & (!g3634) & (g3635)) + ((!g2296) & (g1540) & (g3634) & (!g3635)) + ((!g2296) & (g1540) & (g3634) & (g3635)) + ((g2296) & (!g1540) & (!g3634) & (g3635)) + ((g2296) & (!g1540) & (g3634) & (!g3635)) + ((g2296) & (!g1540) & (g3634) & (g3635)) + ((g2296) & (g1540) & (!g3634) & (!g3635)) + ((g2296) & (g1540) & (!g3634) & (g3635)) + ((g2296) & (g1540) & (g3634) & (!g3635)) + ((g2296) & (g1540) & (g3634) & (g3635)));
	assign g5453 = (((!g3648) & (g3649)) + ((g3648) & (!g3649)) + ((g3648) & (g3649)));
	assign g5454 = (((!g830) & (!g3291) & (!g5902) & (key[29])) + ((!g830) & (!g3291) & (g5902) & (key[29])) + ((!g830) & (g3291) & (!g5902) & (key[29])) + ((!g830) & (g3291) & (g5902) & (key[29])) + ((g830) & (!g3291) & (g5902) & (!key[29])) + ((g830) & (!g3291) & (g5902) & (key[29])) + ((g830) & (g3291) & (!g5902) & (!key[29])) + ((g830) & (g3291) & (!g5902) & (key[29])));
	assign g5455 = (((!g3540) & (!g3541)));
	assign g5456 = (((g1914) & (!g2003) & (!g5455) & (!g2456)) + ((g1914) & (!g2003) & (g5455) & (g2456)) + ((g1914) & (g2003) & (!g5455) & (g2456)) + ((g1914) & (g2003) & (g5455) & (!g2456)));
	assign g5457 = (((!g1962) & (g2393) & (g3549)) + ((g1962) & (!g2393) & (g3549)) + ((g1962) & (g2393) & (!g3549)) + ((g1962) & (g2393) & (g3549)));
	assign g5458 = (((!g1914) & (!g1967) & (!g2474) & (g5457)) + ((!g1914) & (!g1967) & (g2474) & (!g5457)) + ((!g1914) & (g1967) & (!g2474) & (!g5457)) + ((!g1914) & (g1967) & (g2474) & (g5457)));
	assign g5459 = (((!g830) & (!g3295) & (!g5456) & (!g5458)) + ((!g830) & (!g3295) & (!g5456) & (g5458)) + ((!g830) & (!g3295) & (g5456) & (!g5458)) + ((!g830) & (!g3295) & (g5456) & (g5458)) + ((!g830) & (g3295) & (!g5456) & (!g5458)) + ((!g830) & (g3295) & (!g5456) & (g5458)) + ((!g830) & (g3295) & (g5456) & (!g5458)) + ((!g830) & (g3295) & (g5456) & (g5458)) + ((g830) & (!g3295) & (!g5456) & (g5458)) + ((g830) & (!g3295) & (g5456) & (!g5458)) + ((g830) & (!g3295) & (g5456) & (g5458)) + ((g830) & (g3295) & (!g5456) & (!g5458)));
	assign g5460 = (((!g3664) & (!g3665)));
	assign g5461 = (((!g2100) & (!g2742) & (!g5460)) + ((!g2100) & (g2742) & (g5460)) + ((g2100) & (!g2742) & (g5460)) + ((g2100) & (g2742) & (!g5460)));
	assign g5462 = (((!g2916) & (!g3009) & (!g2962) & (g3013) & (!g5432)) + ((!g2916) & (!g3009) & (!g2962) & (g3013) & (g5432)) + ((!g2916) & (!g3009) & (g2962) & (!g3013) & (!g5432)) + ((!g2916) & (!g3009) & (g2962) & (g3013) & (g5432)) + ((!g2916) & (g3009) & (!g2962) & (!g3013) & (!g5432)) + ((!g2916) & (g3009) & (!g2962) & (!g3013) & (g5432)) + ((!g2916) & (g3009) & (g2962) & (!g3013) & (g5432)) + ((!g2916) & (g3009) & (g2962) & (g3013) & (!g5432)) + ((g2916) & (!g3009) & (!g2962) & (!g3013) & (!g5432)) + ((g2916) & (!g3009) & (!g2962) & (g3013) & (g5432)) + ((g2916) & (!g3009) & (g2962) & (!g3013) & (!g5432)) + ((g2916) & (!g3009) & (g2962) & (!g3013) & (g5432)) + ((g2916) & (g3009) & (!g2962) & (!g3013) & (g5432)) + ((g2916) & (g3009) & (!g2962) & (g3013) & (!g5432)) + ((g2916) & (g3009) & (g2962) & (g3013) & (!g5432)) + ((g2916) & (g3009) & (g2962) & (g3013) & (g5432)));
	assign g8337 = (((!g5560) & (g5645) & (!g5463)) + ((!g5560) & (g5645) & (g5463)) + ((g5560) & (!g5645) & (g5463)) + ((g5560) & (g5645) & (g5463)));
	assign g5464 = (((!g830) & (!g1914) & (!g3297) & (!g5461) & (!g5462) & (g5463)) + ((!g830) & (!g1914) & (!g3297) & (!g5461) & (g5462) & (g5463)) + ((!g830) & (!g1914) & (!g3297) & (g5461) & (!g5462) & (g5463)) + ((!g830) & (!g1914) & (!g3297) & (g5461) & (g5462) & (g5463)) + ((!g830) & (!g1914) & (g3297) & (!g5461) & (!g5462) & (g5463)) + ((!g830) & (!g1914) & (g3297) & (!g5461) & (g5462) & (g5463)) + ((!g830) & (!g1914) & (g3297) & (g5461) & (!g5462) & (g5463)) + ((!g830) & (!g1914) & (g3297) & (g5461) & (g5462) & (g5463)) + ((!g830) & (g1914) & (!g3297) & (!g5461) & (!g5462) & (g5463)) + ((!g830) & (g1914) & (!g3297) & (!g5461) & (g5462) & (g5463)) + ((!g830) & (g1914) & (!g3297) & (g5461) & (!g5462) & (g5463)) + ((!g830) & (g1914) & (!g3297) & (g5461) & (g5462) & (g5463)) + ((!g830) & (g1914) & (g3297) & (!g5461) & (!g5462) & (g5463)) + ((!g830) & (g1914) & (g3297) & (!g5461) & (g5462) & (g5463)) + ((!g830) & (g1914) & (g3297) & (g5461) & (!g5462) & (g5463)) + ((!g830) & (g1914) & (g3297) & (g5461) & (g5462) & (g5463)) + ((g830) & (!g1914) & (!g3297) & (!g5461) & (g5462) & (!g5463)) + ((g830) & (!g1914) & (!g3297) & (!g5461) & (g5462) & (g5463)) + ((g830) & (!g1914) & (!g3297) & (g5461) & (g5462) & (!g5463)) + ((g830) & (!g1914) & (!g3297) & (g5461) & (g5462) & (g5463)) + ((g830) & (!g1914) & (g3297) & (!g5461) & (!g5462) & (!g5463)) + ((g830) & (!g1914) & (g3297) & (!g5461) & (!g5462) & (g5463)) + ((g830) & (!g1914) & (g3297) & (g5461) & (!g5462) & (!g5463)) + ((g830) & (!g1914) & (g3297) & (g5461) & (!g5462) & (g5463)) + ((g830) & (g1914) & (!g3297) & (g5461) & (!g5462) & (!g5463)) + ((g830) & (g1914) & (!g3297) & (g5461) & (!g5462) & (g5463)) + ((g830) & (g1914) & (!g3297) & (g5461) & (g5462) & (!g5463)) + ((g830) & (g1914) & (!g3297) & (g5461) & (g5462) & (g5463)) + ((g830) & (g1914) & (g3297) & (!g5461) & (!g5462) & (!g5463)) + ((g830) & (g1914) & (g3297) & (!g5461) & (!g5462) & (g5463)) + ((g830) & (g1914) & (g3297) & (!g5461) & (g5462) & (!g5463)) + ((g830) & (g1914) & (g3297) & (!g5461) & (g5462) & (g5463)));
	assign g5465 = (((!g2932) & (g2938) & (!g3791) & (g3792)) + ((!g2932) & (g2938) & (g3791) & (!g3792)) + ((!g2932) & (g2938) & (g3791) & (g3792)) + ((g2932) & (!g2938) & (!g3791) & (g3792)) + ((g2932) & (!g2938) & (g3791) & (!g3792)) + ((g2932) & (!g2938) & (g3791) & (g3792)) + ((g2932) & (g2938) & (!g3791) & (!g3792)) + ((g2932) & (g2938) & (!g3791) & (g3792)) + ((g2932) & (g2938) & (g3791) & (!g3792)) + ((g2932) & (g2938) & (g3791) & (g3792)));
	assign g5466 = (((!g3805) & (g3806)) + ((g3805) & (!g3806)) + ((g3805) & (g3806)));
	assign g5467 = (((!g830) & (!g3299) & (!g5889) & (key[157])) + ((!g830) & (!g3299) & (g5889) & (key[157])) + ((!g830) & (g3299) & (!g5889) & (key[157])) + ((!g830) & (g3299) & (g5889) & (key[157])) + ((g830) & (!g3299) & (g5889) & (!key[157])) + ((g830) & (!g3299) & (g5889) & (key[157])) + ((g830) & (g3299) & (!g5889) & (!key[157])) + ((g830) & (g3299) & (!g5889) & (key[157])));
	assign g5468 = (((!g2299) & (g1540) & (!g3457) & (g3458)) + ((!g2299) & (g1540) & (g3457) & (!g3458)) + ((!g2299) & (g1540) & (g3457) & (g3458)) + ((g2299) & (!g1540) & (!g3457) & (g3458)) + ((g2299) & (!g1540) & (g3457) & (!g3458)) + ((g2299) & (!g1540) & (g3457) & (g3458)) + ((g2299) & (g1540) & (!g3457) & (!g3458)) + ((g2299) & (g1540) & (!g3457) & (g3458)) + ((g2299) & (g1540) & (g3457) & (!g3458)) + ((g2299) & (g1540) & (g3457) & (g3458)));
	assign g5469 = (((!g3440) & (g3441)) + ((g3440) & (!g3441)) + ((g3440) & (g3441)));
	assign g5470 = (((!g830) & (!g3301) & (!g5876) & (key[125])) + ((!g830) & (!g3301) & (g5876) & (key[125])) + ((!g830) & (g3301) & (!g5876) & (key[125])) + ((!g830) & (g3301) & (g5876) & (key[125])) + ((g830) & (!g3301) & (g5876) & (!key[125])) + ((g830) & (!g3301) & (g5876) & (key[125])) + ((g830) & (g3301) & (!g5876) & (!key[125])) + ((g830) & (g3301) & (!g5876) & (key[125])));
	assign g5471 = (((!g2950) & (!g3568) & (g3569) & (g2962)) + ((!g2950) & (g3568) & (!g3569) & (g2962)) + ((!g2950) & (g3568) & (g3569) & (g2962)) + ((g2950) & (!g3568) & (!g3569) & (g2962)) + ((g2950) & (!g3568) & (g3569) & (!g2962)) + ((g2950) & (!g3568) & (g3569) & (g2962)) + ((g2950) & (g3568) & (!g3569) & (!g2962)) + ((g2950) & (g3568) & (!g3569) & (g2962)) + ((g2950) & (g3568) & (g3569) & (!g2962)) + ((g2950) & (g3568) & (g3569) & (g2962)));
	assign g5472 = (((!g3582) & (g3583)) + ((g3582) & (!g3583)) + ((g3582) & (g3583)));
	assign g5473 = (((!g830) & (!g3303) & (!g5863) & (nonce[29])) + ((!g830) & (!g3303) & (g5863) & (nonce[29])) + ((!g830) & (g3303) & (!g5863) & (nonce[29])) + ((!g830) & (g3303) & (g5863) & (nonce[29])) + ((g830) & (!g3303) & (g5863) & (!nonce[29])) + ((g830) & (!g3303) & (g5863) & (nonce[29])) + ((g830) & (g3303) & (!g5863) & (!nonce[29])) + ((g830) & (g3303) & (!g5863) & (nonce[29])));
	assign g5474 = (((!g3695) & (!g3696)));
	assign g5475 = (((g1914) & (!g2468) & (!g2486) & (!g5474)) + ((g1914) & (!g2468) & (g2486) & (g5474)) + ((g1914) & (g2468) & (!g2486) & (g5474)) + ((g1914) & (g2468) & (g2486) & (!g5474)));
	assign g5476 = (((!g2399) & (g2408) & (g3704)) + ((g2399) & (!g2408) & (g3704)) + ((g2399) & (g2408) & (!g3704)) + ((g2399) & (g2408) & (g3704)));
	assign g5477 = (((!g1914) & (!g2434) & (!g2503) & (g5476)) + ((!g1914) & (!g2434) & (g2503) & (!g5476)) + ((!g1914) & (g2434) & (!g2503) & (!g5476)) + ((!g1914) & (g2434) & (g2503) & (g5476)));
	assign g5478 = (((!g830) & (!g3305) & (!g5475) & (!g5477)) + ((!g830) & (!g3305) & (!g5475) & (g5477)) + ((!g830) & (!g3305) & (g5475) & (!g5477)) + ((!g830) & (!g3305) & (g5475) & (g5477)) + ((!g830) & (g3305) & (!g5475) & (!g5477)) + ((!g830) & (g3305) & (!g5475) & (g5477)) + ((!g830) & (g3305) & (g5475) & (!g5477)) + ((!g830) & (g3305) & (g5475) & (g5477)) + ((g830) & (!g3305) & (!g5475) & (g5477)) + ((g830) & (!g3305) & (g5475) & (!g5477)) + ((g830) & (!g3305) & (g5475) & (g5477)) + ((g830) & (g3305) & (!g5475) & (!g5477)));
	assign g5479 = (((!g2857) & (!g2860) & (!g2895) & (g2887) & (!g5446)) + ((!g2857) & (!g2860) & (!g2895) & (g2887) & (g5446)) + ((!g2857) & (!g2860) & (g2895) & (!g2887) & (!g5446)) + ((!g2857) & (!g2860) & (g2895) & (!g2887) & (g5446)) + ((!g2857) & (g2860) & (!g2895) & (!g2887) & (g5446)) + ((!g2857) & (g2860) & (!g2895) & (g2887) & (!g5446)) + ((!g2857) & (g2860) & (g2895) & (!g2887) & (!g5446)) + ((!g2857) & (g2860) & (g2895) & (g2887) & (g5446)) + ((g2857) & (!g2860) & (!g2895) & (!g2887) & (g5446)) + ((g2857) & (!g2860) & (!g2895) & (g2887) & (!g5446)) + ((g2857) & (!g2860) & (g2895) & (!g2887) & (!g5446)) + ((g2857) & (!g2860) & (g2895) & (g2887) & (g5446)) + ((g2857) & (g2860) & (!g2895) & (!g2887) & (!g5446)) + ((g2857) & (g2860) & (!g2895) & (!g2887) & (g5446)) + ((g2857) & (g2860) & (g2895) & (g2887) & (!g5446)) + ((g2857) & (g2860) & (g2895) & (g2887) & (g5446)));
	assign g5480 = (((!g2211) & (!g2257) & (!g2874) & (g2904) & (!g5448)) + ((!g2211) & (!g2257) & (!g2874) & (g2904) & (g5448)) + ((!g2211) & (!g2257) & (g2874) & (!g2904) & (g5448)) + ((!g2211) & (!g2257) & (g2874) & (g2904) & (!g5448)) + ((!g2211) & (g2257) & (!g2874) & (!g2904) & (!g5448)) + ((!g2211) & (g2257) & (!g2874) & (!g2904) & (g5448)) + ((!g2211) & (g2257) & (g2874) & (!g2904) & (!g5448)) + ((!g2211) & (g2257) & (g2874) & (g2904) & (g5448)) + ((g2211) & (!g2257) & (!g2874) & (!g2904) & (g5448)) + ((g2211) & (!g2257) & (!g2874) & (g2904) & (!g5448)) + ((g2211) & (!g2257) & (g2874) & (!g2904) & (!g5448)) + ((g2211) & (!g2257) & (g2874) & (!g2904) & (g5448)) + ((g2211) & (g2257) & (!g2874) & (!g2904) & (!g5448)) + ((g2211) & (g2257) & (!g2874) & (g2904) & (g5448)) + ((g2211) & (g2257) & (g2874) & (g2904) & (!g5448)) + ((g2211) & (g2257) & (g2874) & (g2904) & (g5448)));
	assign g5481 = (((!g830) & (!g1914) & (!g3307) & (!g5479) & (!g5480) & (nonce[61])) + ((!g830) & (!g1914) & (!g3307) & (!g5479) & (g5480) & (nonce[61])) + ((!g830) & (!g1914) & (!g3307) & (g5479) & (!g5480) & (nonce[61])) + ((!g830) & (!g1914) & (!g3307) & (g5479) & (g5480) & (nonce[61])) + ((!g830) & (!g1914) & (g3307) & (!g5479) & (!g5480) & (nonce[61])) + ((!g830) & (!g1914) & (g3307) & (!g5479) & (g5480) & (nonce[61])) + ((!g830) & (!g1914) & (g3307) & (g5479) & (!g5480) & (nonce[61])) + ((!g830) & (!g1914) & (g3307) & (g5479) & (g5480) & (nonce[61])) + ((!g830) & (g1914) & (!g3307) & (!g5479) & (!g5480) & (nonce[61])) + ((!g830) & (g1914) & (!g3307) & (!g5479) & (g5480) & (nonce[61])) + ((!g830) & (g1914) & (!g3307) & (g5479) & (!g5480) & (nonce[61])) + ((!g830) & (g1914) & (!g3307) & (g5479) & (g5480) & (nonce[61])) + ((!g830) & (g1914) & (g3307) & (!g5479) & (!g5480) & (nonce[61])) + ((!g830) & (g1914) & (g3307) & (!g5479) & (g5480) & (nonce[61])) + ((!g830) & (g1914) & (g3307) & (g5479) & (!g5480) & (nonce[61])) + ((!g830) & (g1914) & (g3307) & (g5479) & (g5480) & (nonce[61])) + ((g830) & (!g1914) & (!g3307) & (!g5479) & (g5480) & (!nonce[61])) + ((g830) & (!g1914) & (!g3307) & (!g5479) & (g5480) & (nonce[61])) + ((g830) & (!g1914) & (!g3307) & (g5479) & (g5480) & (!nonce[61])) + ((g830) & (!g1914) & (!g3307) & (g5479) & (g5480) & (nonce[61])) + ((g830) & (!g1914) & (g3307) & (!g5479) & (!g5480) & (!nonce[61])) + ((g830) & (!g1914) & (g3307) & (!g5479) & (!g5480) & (nonce[61])) + ((g830) & (!g1914) & (g3307) & (g5479) & (!g5480) & (!nonce[61])) + ((g830) & (!g1914) & (g3307) & (g5479) & (!g5480) & (nonce[61])) + ((g830) & (g1914) & (!g3307) & (g5479) & (!g5480) & (!nonce[61])) + ((g830) & (g1914) & (!g3307) & (g5479) & (!g5480) & (nonce[61])) + ((g830) & (g1914) & (!g3307) & (g5479) & (g5480) & (!nonce[61])) + ((g830) & (g1914) & (!g3307) & (g5479) & (g5480) & (nonce[61])) + ((g830) & (g1914) & (g3307) & (!g5479) & (!g5480) & (!nonce[61])) + ((g830) & (g1914) & (g3307) & (!g5479) & (!g5480) & (nonce[61])) + ((g830) & (g1914) & (g3307) & (!g5479) & (g5480) & (!nonce[61])) + ((g830) & (g1914) & (g3307) & (!g5479) & (g5480) & (nonce[61])));
	assign g5482 = (((!g2932) & (!g3615) & (g3616) & (g2956)) + ((!g2932) & (g3615) & (!g3616) & (g2956)) + ((!g2932) & (g3615) & (g3616) & (g2956)) + ((g2932) & (!g3615) & (!g3616) & (g2956)) + ((g2932) & (!g3615) & (g3616) & (!g2956)) + ((g2932) & (!g3615) & (g3616) & (g2956)) + ((g2932) & (g3615) & (!g3616) & (!g2956)) + ((g2932) & (g3615) & (!g3616) & (g2956)) + ((g2932) & (g3615) & (g3616) & (!g2956)) + ((g2932) & (g3615) & (g3616) & (g2956)));
	assign g5483 = (((!g3598) & (g3599)) + ((g3598) & (!g3599)) + ((g3598) & (g3599)));
	assign g5484 = (((!g830) & (!g3310) & (!g5850) & (key[253])) + ((!g830) & (!g3310) & (g5850) & (key[253])) + ((!g830) & (g3310) & (!g5850) & (key[253])) + ((!g830) & (g3310) & (g5850) & (key[253])) + ((g830) & (!g3310) & (g5850) & (!key[253])) + ((g830) & (!g3310) & (g5850) & (key[253])) + ((g830) & (g3310) & (!g5850) & (!key[253])) + ((g830) & (g3310) & (!g5850) & (key[253])));
	assign g5485 = (((!g2213) & (!g2263) & (!g2874) & (g2904) & (!g5437)) + ((!g2213) & (!g2263) & (!g2874) & (g2904) & (g5437)) + ((!g2213) & (!g2263) & (g2874) & (!g2904) & (g5437)) + ((!g2213) & (!g2263) & (g2874) & (g2904) & (!g5437)) + ((!g2213) & (g2263) & (!g2874) & (!g2904) & (!g5437)) + ((!g2213) & (g2263) & (!g2874) & (!g2904) & (g5437)) + ((!g2213) & (g2263) & (g2874) & (!g2904) & (!g5437)) + ((!g2213) & (g2263) & (g2874) & (g2904) & (g5437)) + ((g2213) & (!g2263) & (!g2874) & (!g2904) & (g5437)) + ((g2213) & (!g2263) & (!g2874) & (g2904) & (!g5437)) + ((g2213) & (!g2263) & (g2874) & (!g2904) & (!g5437)) + ((g2213) & (!g2263) & (g2874) & (!g2904) & (g5437)) + ((g2213) & (g2263) & (!g2874) & (!g2904) & (!g5437)) + ((g2213) & (g2263) & (!g2874) & (g2904) & (g5437)) + ((g2213) & (g2263) & (g2874) & (g2904) & (!g5437)) + ((g2213) & (g2263) & (g2874) & (g2904) & (g5437)));
	assign g5486 = (((!g2860) & (!g2895) & (!g2848) & (!g5439) & (g2893)) + ((!g2860) & (!g2895) & (!g2848) & (g5439) & (g2893)) + ((!g2860) & (!g2895) & (g2848) & (!g5439) & (g2893)) + ((!g2860) & (!g2895) & (g2848) & (g5439) & (!g2893)) + ((!g2860) & (g2895) & (!g2848) & (!g5439) & (!g2893)) + ((!g2860) & (g2895) & (!g2848) & (g5439) & (!g2893)) + ((!g2860) & (g2895) & (g2848) & (!g5439) & (!g2893)) + ((!g2860) & (g2895) & (g2848) & (g5439) & (g2893)) + ((g2860) & (!g2895) & (!g2848) & (!g5439) & (g2893)) + ((g2860) & (!g2895) & (!g2848) & (g5439) & (!g2893)) + ((g2860) & (!g2895) & (g2848) & (!g5439) & (!g2893)) + ((g2860) & (!g2895) & (g2848) & (g5439) & (!g2893)) + ((g2860) & (g2895) & (!g2848) & (!g5439) & (!g2893)) + ((g2860) & (g2895) & (!g2848) & (g5439) & (g2893)) + ((g2860) & (g2895) & (g2848) & (!g5439) & (g2893)) + ((g2860) & (g2895) & (g2848) & (g5439) & (g2893)));
	assign g5487 = (((!g830) & (!g1914) & (!g3312) & (!g5485) & (!g5486) & (key[221])) + ((!g830) & (!g1914) & (!g3312) & (!g5485) & (g5486) & (key[221])) + ((!g830) & (!g1914) & (!g3312) & (g5485) & (!g5486) & (key[221])) + ((!g830) & (!g1914) & (!g3312) & (g5485) & (g5486) & (key[221])) + ((!g830) & (!g1914) & (g3312) & (!g5485) & (!g5486) & (key[221])) + ((!g830) & (!g1914) & (g3312) & (!g5485) & (g5486) & (key[221])) + ((!g830) & (!g1914) & (g3312) & (g5485) & (!g5486) & (key[221])) + ((!g830) & (!g1914) & (g3312) & (g5485) & (g5486) & (key[221])) + ((!g830) & (g1914) & (!g3312) & (!g5485) & (!g5486) & (key[221])) + ((!g830) & (g1914) & (!g3312) & (!g5485) & (g5486) & (key[221])) + ((!g830) & (g1914) & (!g3312) & (g5485) & (!g5486) & (key[221])) + ((!g830) & (g1914) & (!g3312) & (g5485) & (g5486) & (key[221])) + ((!g830) & (g1914) & (g3312) & (!g5485) & (!g5486) & (key[221])) + ((!g830) & (g1914) & (g3312) & (!g5485) & (g5486) & (key[221])) + ((!g830) & (g1914) & (g3312) & (g5485) & (!g5486) & (key[221])) + ((!g830) & (g1914) & (g3312) & (g5485) & (g5486) & (key[221])) + ((g830) & (!g1914) & (!g3312) & (!g5485) & (g5486) & (!key[221])) + ((g830) & (!g1914) & (!g3312) & (!g5485) & (g5486) & (key[221])) + ((g830) & (!g1914) & (!g3312) & (g5485) & (g5486) & (!key[221])) + ((g830) & (!g1914) & (!g3312) & (g5485) & (g5486) & (key[221])) + ((g830) & (!g1914) & (g3312) & (!g5485) & (!g5486) & (!key[221])) + ((g830) & (!g1914) & (g3312) & (!g5485) & (!g5486) & (key[221])) + ((g830) & (!g1914) & (g3312) & (g5485) & (!g5486) & (!key[221])) + ((g830) & (!g1914) & (g3312) & (g5485) & (!g5486) & (key[221])) + ((g830) & (g1914) & (!g3312) & (g5485) & (!g5486) & (!key[221])) + ((g830) & (g1914) & (!g3312) & (g5485) & (!g5486) & (key[221])) + ((g830) & (g1914) & (!g3312) & (g5485) & (g5486) & (!key[221])) + ((g830) & (g1914) & (!g3312) & (g5485) & (g5486) & (key[221])) + ((g830) & (g1914) & (g3312) & (!g5485) & (!g5486) & (!key[221])) + ((g830) & (g1914) & (g3312) & (!g5485) & (!g5486) & (key[221])) + ((g830) & (g1914) & (g3312) & (!g5485) & (g5486) & (!key[221])) + ((g830) & (g1914) & (g3312) & (!g5485) & (g5486) & (key[221])));
	assign g5488 = (((!g3852) & (!g3853)));
	assign g5489 = (((g1914) & (!g2497) & (!g2503) & (!g5488)) + ((g1914) & (!g2497) & (g2503) & (g5488)) + ((g1914) & (g2497) & (!g2503) & (g5488)) + ((g1914) & (g2497) & (g2503) & (!g5488)));
	assign g5490 = (((!g2413) & (g2416) & (g3861)) + ((g2413) & (!g2416) & (g3861)) + ((g2413) & (g2416) & (!g3861)) + ((g2413) & (g2416) & (g3861)));
	assign g5491 = (((!g1914) & (!g2462) & (!g2486) & (g5490)) + ((!g1914) & (!g2462) & (g2486) & (!g5490)) + ((!g1914) & (g2462) & (!g2486) & (!g5490)) + ((!g1914) & (g2462) & (g2486) & (g5490)));
	assign g5492 = (((!g830) & (!g3314) & (!g5489) & (!g5491)) + ((!g830) & (!g3314) & (!g5489) & (g5491)) + ((!g830) & (!g3314) & (g5489) & (!g5491)) + ((!g830) & (!g3314) & (g5489) & (g5491)) + ((!g830) & (g3314) & (!g5489) & (!g5491)) + ((!g830) & (g3314) & (!g5489) & (g5491)) + ((!g830) & (g3314) & (g5489) & (!g5491)) + ((!g830) & (g3314) & (g5489) & (g5491)) + ((g830) & (!g3314) & (!g5489) & (g5491)) + ((g830) & (!g3314) & (g5489) & (!g5491)) + ((g830) & (!g3314) & (g5489) & (g5491)) + ((g830) & (g3314) & (!g5489) & (!g5491)));
	assign g5493 = (((!g5469) & (!g2708) & (!g2747) & (!g2776) & (g2780)) + ((!g5469) & (!g2708) & (!g2747) & (g2776) & (!g2780)) + ((!g5469) & (!g2708) & (g2747) & (!g2776) & (g2780)) + ((!g5469) & (!g2708) & (g2747) & (g2776) & (!g2780)) + ((!g5469) & (g2708) & (!g2747) & (!g2776) & (g2780)) + ((!g5469) & (g2708) & (!g2747) & (g2776) & (!g2780)) + ((!g5469) & (g2708) & (g2747) & (!g2776) & (!g2780)) + ((!g5469) & (g2708) & (g2747) & (g2776) & (g2780)) + ((g5469) & (!g2708) & (!g2747) & (!g2776) & (g2780)) + ((g5469) & (!g2708) & (!g2747) & (g2776) & (!g2780)) + ((g5469) & (!g2708) & (g2747) & (!g2776) & (!g2780)) + ((g5469) & (!g2708) & (g2747) & (g2776) & (g2780)) + ((g5469) & (g2708) & (!g2747) & (!g2776) & (!g2780)) + ((g5469) & (g2708) & (!g2747) & (g2776) & (g2780)) + ((g5469) & (g2708) & (g2747) & (!g2776) & (!g2780)) + ((g5469) & (g2708) & (g2747) & (g2776) & (g2780)));
	assign g5494 = (((!g1914) & (!g2379) & (!g1610) & (!g3459) & (!g5493)) + ((!g1914) & (!g2379) & (!g1610) & (!g3459) & (g5493)) + ((!g1914) & (!g2379) & (g1610) & (g3459) & (!g5493)) + ((!g1914) & (!g2379) & (g1610) & (g3459) & (g5493)) + ((!g1914) & (g2379) & (!g1610) & (g3459) & (!g5493)) + ((!g1914) & (g2379) & (!g1610) & (g3459) & (g5493)) + ((!g1914) & (g2379) & (g1610) & (!g3459) & (!g5493)) + ((!g1914) & (g2379) & (g1610) & (!g3459) & (g5493)) + ((g1914) & (!g2379) & (!g1610) & (!g3459) & (g5493)) + ((g1914) & (!g2379) & (!g1610) & (g3459) & (g5493)) + ((g1914) & (!g2379) & (g1610) & (!g3459) & (g5493)) + ((g1914) & (!g2379) & (g1610) & (g3459) & (g5493)) + ((g1914) & (g2379) & (!g1610) & (!g3459) & (g5493)) + ((g1914) & (g2379) & (!g1610) & (g3459) & (g5493)) + ((g1914) & (g2379) & (g1610) & (!g3459) & (g5493)) + ((g1914) & (g2379) & (g1610) & (g3459) & (g5493)));
	assign g5495 = (((!g830) & (!g3323) & (!g5494) & (key[126])) + ((!g830) & (!g3323) & (g5494) & (key[126])) + ((!g830) & (g3323) & (!g5494) & (key[126])) + ((!g830) & (g3323) & (g5494) & (key[126])) + ((g830) & (!g3323) & (g5494) & (!key[126])) + ((g830) & (!g3323) & (g5494) & (key[126])) + ((g830) & (g3323) & (!g5494) & (!key[126])) + ((g830) & (g3323) & (!g5494) & (key[126])));
	assign g5496 = (((!g2003) & (!g2005) & (!g5455) & (!g2456) & (g2535)) + ((!g2003) & (!g2005) & (!g5455) & (g2456) & (!g2535)) + ((!g2003) & (!g2005) & (g5455) & (!g2456) & (g2535)) + ((!g2003) & (!g2005) & (g5455) & (g2456) & (g2535)) + ((!g2003) & (g2005) & (!g5455) & (!g2456) & (!g2535)) + ((!g2003) & (g2005) & (!g5455) & (g2456) & (g2535)) + ((!g2003) & (g2005) & (g5455) & (!g2456) & (!g2535)) + ((!g2003) & (g2005) & (g5455) & (g2456) & (!g2535)) + ((g2003) & (!g2005) & (!g5455) & (!g2456) & (!g2535)) + ((g2003) & (!g2005) & (!g5455) & (g2456) & (!g2535)) + ((g2003) & (!g2005) & (g5455) & (!g2456) & (g2535)) + ((g2003) & (!g2005) & (g5455) & (g2456) & (!g2535)) + ((g2003) & (g2005) & (!g5455) & (!g2456) & (g2535)) + ((g2003) & (g2005) & (!g5455) & (g2456) & (g2535)) + ((g2003) & (g2005) & (g5455) & (!g2456) & (!g2535)) + ((g2003) & (g2005) & (g5455) & (g2456) & (g2535)));
	assign g5497 = (((!g1967) & (!g1969) & (!g2474) & (g2529) & (!g5457)) + ((!g1967) & (!g1969) & (!g2474) & (g2529) & (g5457)) + ((!g1967) & (!g1969) & (g2474) & (!g2529) & (g5457)) + ((!g1967) & (!g1969) & (g2474) & (g2529) & (!g5457)) + ((!g1967) & (g1969) & (!g2474) & (!g2529) & (!g5457)) + ((!g1967) & (g1969) & (!g2474) & (!g2529) & (g5457)) + ((!g1967) & (g1969) & (g2474) & (!g2529) & (!g5457)) + ((!g1967) & (g1969) & (g2474) & (g2529) & (g5457)) + ((g1967) & (!g1969) & (!g2474) & (!g2529) & (g5457)) + ((g1967) & (!g1969) & (!g2474) & (g2529) & (!g5457)) + ((g1967) & (!g1969) & (g2474) & (!g2529) & (!g5457)) + ((g1967) & (!g1969) & (g2474) & (!g2529) & (g5457)) + ((g1967) & (g1969) & (!g2474) & (!g2529) & (!g5457)) + ((g1967) & (g1969) & (!g2474) & (g2529) & (g5457)) + ((g1967) & (g1969) & (g2474) & (g2529) & (!g5457)) + ((g1967) & (g1969) & (g2474) & (g2529) & (g5457)));
	assign g5498 = (((!g830) & (!g1914) & (!g3330) & (!g5496) & (!g5497)) + ((!g830) & (!g1914) & (!g3330) & (!g5496) & (g5497)) + ((!g830) & (!g1914) & (!g3330) & (g5496) & (!g5497)) + ((!g830) & (!g1914) & (!g3330) & (g5496) & (g5497)) + ((!g830) & (!g1914) & (g3330) & (!g5496) & (!g5497)) + ((!g830) & (!g1914) & (g3330) & (!g5496) & (g5497)) + ((!g830) & (!g1914) & (g3330) & (g5496) & (!g5497)) + ((!g830) & (!g1914) & (g3330) & (g5496) & (g5497)) + ((!g830) & (g1914) & (!g3330) & (!g5496) & (!g5497)) + ((!g830) & (g1914) & (!g3330) & (!g5496) & (g5497)) + ((!g830) & (g1914) & (!g3330) & (g5496) & (!g5497)) + ((!g830) & (g1914) & (!g3330) & (g5496) & (g5497)) + ((!g830) & (g1914) & (g3330) & (!g5496) & (!g5497)) + ((!g830) & (g1914) & (g3330) & (!g5496) & (g5497)) + ((!g830) & (g1914) & (g3330) & (g5496) & (!g5497)) + ((!g830) & (g1914) & (g3330) & (g5496) & (g5497)) + ((g830) & (!g1914) & (!g3330) & (!g5496) & (g5497)) + ((g830) & (!g1914) & (!g3330) & (g5496) & (g5497)) + ((g830) & (!g1914) & (g3330) & (!g5496) & (!g5497)) + ((g830) & (!g1914) & (g3330) & (g5496) & (!g5497)) + ((g830) & (g1914) & (!g3330) & (g5496) & (!g5497)) + ((g830) & (g1914) & (!g3330) & (g5496) & (g5497)) + ((g830) & (g1914) & (g3330) & (!g5496) & (!g5497)) + ((g830) & (g1914) & (g3330) & (!g5496) & (g5497)));
	assign g5499 = (((!g2098) & (!g2129) & (!g2713) & (g2783) & (!g5472)) + ((!g2098) & (!g2129) & (!g2713) & (g2783) & (g5472)) + ((!g2098) & (!g2129) & (g2713) & (!g2783) & (g5472)) + ((!g2098) & (!g2129) & (g2713) & (g2783) & (!g5472)) + ((!g2098) & (g2129) & (!g2713) & (!g2783) & (!g5472)) + ((!g2098) & (g2129) & (!g2713) & (!g2783) & (g5472)) + ((!g2098) & (g2129) & (g2713) & (!g2783) & (!g5472)) + ((!g2098) & (g2129) & (g2713) & (g2783) & (g5472)) + ((g2098) & (!g2129) & (!g2713) & (!g2783) & (g5472)) + ((g2098) & (!g2129) & (!g2713) & (g2783) & (!g5472)) + ((g2098) & (!g2129) & (g2713) & (!g2783) & (!g5472)) + ((g2098) & (!g2129) & (g2713) & (!g2783) & (g5472)) + ((g2098) & (g2129) & (!g2713) & (!g2783) & (!g5472)) + ((g2098) & (g2129) & (!g2713) & (g2783) & (g5472)) + ((g2098) & (g2129) & (g2713) & (g2783) & (!g5472)) + ((g2098) & (g2129) & (g2713) & (g2783) & (g5472)));
	assign g5500 = (((!g1914) & (!g3047) & (!g3570) & (!g3053) & (g5499)) + ((!g1914) & (!g3047) & (!g3570) & (g3053) & (g5499)) + ((!g1914) & (!g3047) & (g3570) & (!g3053) & (g5499)) + ((!g1914) & (!g3047) & (g3570) & (g3053) & (g5499)) + ((!g1914) & (g3047) & (!g3570) & (!g3053) & (g5499)) + ((!g1914) & (g3047) & (!g3570) & (g3053) & (g5499)) + ((!g1914) & (g3047) & (g3570) & (!g3053) & (g5499)) + ((!g1914) & (g3047) & (g3570) & (g3053) & (g5499)) + ((g1914) & (!g3047) & (!g3570) & (!g3053) & (!g5499)) + ((g1914) & (!g3047) & (!g3570) & (!g3053) & (g5499)) + ((g1914) & (!g3047) & (g3570) & (g3053) & (!g5499)) + ((g1914) & (!g3047) & (g3570) & (g3053) & (g5499)) + ((g1914) & (g3047) & (!g3570) & (g3053) & (!g5499)) + ((g1914) & (g3047) & (!g3570) & (g3053) & (g5499)) + ((g1914) & (g3047) & (g3570) & (!g3053) & (!g5499)) + ((g1914) & (g3047) & (g3570) & (!g3053) & (g5499)));
	assign g5501 = (((!g830) & (!g3333) & (!g5500) & (nonce[30])) + ((!g830) & (!g3333) & (g5500) & (nonce[30])) + ((!g830) & (g3333) & (!g5500) & (nonce[30])) + ((!g830) & (g3333) & (g5500) & (nonce[30])) + ((g830) & (!g3333) & (g5500) & (!nonce[30])) + ((g830) & (!g3333) & (g5500) & (nonce[30])) + ((g830) & (g3333) & (!g5500) & (!nonce[30])) + ((g830) & (g3333) & (!g5500) & (nonce[30])));
	assign g5502 = (((!g2101) & (!g2134) & (!g5483) & (!g2733) & (g2785)) + ((!g2101) & (!g2134) & (!g5483) & (g2733) & (g2785)) + ((!g2101) & (!g2134) & (g5483) & (!g2733) & (g2785)) + ((!g2101) & (!g2134) & (g5483) & (g2733) & (!g2785)) + ((!g2101) & (g2134) & (!g5483) & (!g2733) & (!g2785)) + ((!g2101) & (g2134) & (!g5483) & (g2733) & (!g2785)) + ((!g2101) & (g2134) & (g5483) & (!g2733) & (!g2785)) + ((!g2101) & (g2134) & (g5483) & (g2733) & (g2785)) + ((g2101) & (!g2134) & (!g5483) & (!g2733) & (g2785)) + ((g2101) & (!g2134) & (!g5483) & (g2733) & (!g2785)) + ((g2101) & (!g2134) & (g5483) & (!g2733) & (!g2785)) + ((g2101) & (!g2134) & (g5483) & (g2733) & (!g2785)) + ((g2101) & (g2134) & (!g5483) & (!g2733) & (!g2785)) + ((g2101) & (g2134) & (!g5483) & (g2733) & (g2785)) + ((g2101) & (g2134) & (g5483) & (!g2733) & (g2785)) + ((g2101) & (g2134) & (g5483) & (g2733) & (g2785)));
	assign g5503 = (((!g1914) & (!g3038) & (!g3617) & (!g3050) & (!g5502)) + ((!g1914) & (!g3038) & (!g3617) & (!g3050) & (g5502)) + ((!g1914) & (!g3038) & (g3617) & (g3050) & (!g5502)) + ((!g1914) & (!g3038) & (g3617) & (g3050) & (g5502)) + ((!g1914) & (g3038) & (!g3617) & (g3050) & (!g5502)) + ((!g1914) & (g3038) & (!g3617) & (g3050) & (g5502)) + ((!g1914) & (g3038) & (g3617) & (!g3050) & (!g5502)) + ((!g1914) & (g3038) & (g3617) & (!g3050) & (g5502)) + ((g1914) & (!g3038) & (!g3617) & (!g3050) & (g5502)) + ((g1914) & (!g3038) & (!g3617) & (g3050) & (g5502)) + ((g1914) & (!g3038) & (g3617) & (!g3050) & (g5502)) + ((g1914) & (!g3038) & (g3617) & (g3050) & (g5502)) + ((g1914) & (g3038) & (!g3617) & (!g3050) & (g5502)) + ((g1914) & (g3038) & (!g3617) & (g3050) & (g5502)) + ((g1914) & (g3038) & (g3617) & (!g3050) & (g5502)) + ((g1914) & (g3038) & (g3617) & (g3050) & (g5502)));
	assign g5504 = (((!g830) & (!g3336) & (!g5503) & (key[254])) + ((!g830) & (!g3336) & (g5503) & (key[254])) + ((!g830) & (g3336) & (!g5503) & (key[254])) + ((!g830) & (g3336) & (g5503) & (key[254])) + ((g830) & (!g3336) & (g5503) & (!key[254])) + ((g830) & (!g3336) & (g5503) & (key[254])) + ((g830) & (g3336) & (!g5503) & (!key[254])) + ((g830) & (g3336) & (!g5503) & (key[254])));
	assign g5505 = (((!g2733) & (!g2785) & (!g5453) & (!g2723) & (g2770)) + ((!g2733) & (!g2785) & (!g5453) & (g2723) & (g2770)) + ((!g2733) & (!g2785) & (g5453) & (!g2723) & (g2770)) + ((!g2733) & (!g2785) & (g5453) & (g2723) & (!g2770)) + ((!g2733) & (g2785) & (!g5453) & (!g2723) & (!g2770)) + ((!g2733) & (g2785) & (!g5453) & (g2723) & (!g2770)) + ((!g2733) & (g2785) & (g5453) & (!g2723) & (!g2770)) + ((!g2733) & (g2785) & (g5453) & (g2723) & (g2770)) + ((g2733) & (!g2785) & (!g5453) & (!g2723) & (g2770)) + ((g2733) & (!g2785) & (!g5453) & (g2723) & (!g2770)) + ((g2733) & (!g2785) & (g5453) & (!g2723) & (!g2770)) + ((g2733) & (!g2785) & (g5453) & (g2723) & (!g2770)) + ((g2733) & (g2785) & (!g5453) & (!g2723) & (!g2770)) + ((g2733) & (g2785) & (!g5453) & (g2723) & (g2770)) + ((g2733) & (g2785) & (g5453) & (!g2723) & (g2770)) + ((g2733) & (g2785) & (g5453) & (g2723) & (g2770)));
	assign g5506 = (((!g1914) & (!g2377) & (!g1610) & (!g3636) & (g5505)) + ((!g1914) & (!g2377) & (!g1610) & (g3636) & (g5505)) + ((!g1914) & (!g2377) & (g1610) & (!g3636) & (g5505)) + ((!g1914) & (!g2377) & (g1610) & (g3636) & (g5505)) + ((!g1914) & (g2377) & (!g1610) & (!g3636) & (g5505)) + ((!g1914) & (g2377) & (!g1610) & (g3636) & (g5505)) + ((!g1914) & (g2377) & (g1610) & (!g3636) & (g5505)) + ((!g1914) & (g2377) & (g1610) & (g3636) & (g5505)) + ((g1914) & (!g2377) & (!g1610) & (!g3636) & (!g5505)) + ((g1914) & (!g2377) & (!g1610) & (!g3636) & (g5505)) + ((g1914) & (!g2377) & (g1610) & (g3636) & (!g5505)) + ((g1914) & (!g2377) & (g1610) & (g3636) & (g5505)) + ((g1914) & (g2377) & (!g1610) & (g3636) & (!g5505)) + ((g1914) & (g2377) & (!g1610) & (g3636) & (g5505)) + ((g1914) & (g2377) & (g1610) & (!g3636) & (!g5505)) + ((g1914) & (g2377) & (g1610) & (!g3636) & (g5505)));
	assign g5507 = (((!g830) & (!g3339) & (!g5506) & (key[30])) + ((!g830) & (!g3339) & (g5506) & (key[30])) + ((!g830) & (g3339) & (!g5506) & (key[30])) + ((!g830) & (g3339) & (g5506) & (key[30])) + ((g830) & (!g3339) & (g5506) & (!key[30])) + ((g830) & (!g3339) & (g5506) & (key[30])) + ((g830) & (g3339) & (!g5506) & (!key[30])) + ((g830) & (g3339) & (!g5506) & (key[30])));
	assign g5508 = (((!g2100) & (!g2133) & (!g2742) & (g2772) & (!g5460)) + ((!g2100) & (!g2133) & (!g2742) & (g2772) & (g5460)) + ((!g2100) & (!g2133) & (g2742) & (!g2772) & (!g5460)) + ((!g2100) & (!g2133) & (g2742) & (g2772) & (g5460)) + ((!g2100) & (g2133) & (!g2742) & (!g2772) & (!g5460)) + ((!g2100) & (g2133) & (!g2742) & (!g2772) & (g5460)) + ((!g2100) & (g2133) & (g2742) & (!g2772) & (g5460)) + ((!g2100) & (g2133) & (g2742) & (g2772) & (!g5460)) + ((g2100) & (!g2133) & (!g2742) & (!g2772) & (!g5460)) + ((g2100) & (!g2133) & (!g2742) & (g2772) & (g5460)) + ((g2100) & (!g2133) & (g2742) & (!g2772) & (!g5460)) + ((g2100) & (!g2133) & (g2742) & (!g2772) & (g5460)) + ((g2100) & (g2133) & (!g2742) & (!g2772) & (g5460)) + ((g2100) & (g2133) & (!g2742) & (g2772) & (!g5460)) + ((g2100) & (g2133) & (g2742) & (g2772) & (!g5460)) + ((g2100) & (g2133) & (g2742) & (g2772) & (g5460)));
	assign g5509 = (((!g3031) & (!g3053) & (!g3684)) + ((!g3031) & (g3053) & (g3684)) + ((g3031) & (!g3053) & (g3684)) + ((g3031) & (g3053) & (!g3684)));
	assign g8338 = (((!g5560) & (g5646) & (!g5510)) + ((!g5560) & (g5646) & (g5510)) + ((g5560) & (!g5646) & (g5510)) + ((g5560) & (g5646) & (g5510)));
	assign g5511 = (((!g830) & (!g1914) & (!g3342) & (!g5508) & (!g5509) & (g5510)) + ((!g830) & (!g1914) & (!g3342) & (!g5508) & (g5509) & (g5510)) + ((!g830) & (!g1914) & (!g3342) & (g5508) & (!g5509) & (g5510)) + ((!g830) & (!g1914) & (!g3342) & (g5508) & (g5509) & (g5510)) + ((!g830) & (!g1914) & (g3342) & (!g5508) & (!g5509) & (g5510)) + ((!g830) & (!g1914) & (g3342) & (!g5508) & (g5509) & (g5510)) + ((!g830) & (!g1914) & (g3342) & (g5508) & (!g5509) & (g5510)) + ((!g830) & (!g1914) & (g3342) & (g5508) & (g5509) & (g5510)) + ((!g830) & (g1914) & (!g3342) & (!g5508) & (!g5509) & (g5510)) + ((!g830) & (g1914) & (!g3342) & (!g5508) & (g5509) & (g5510)) + ((!g830) & (g1914) & (!g3342) & (g5508) & (!g5509) & (g5510)) + ((!g830) & (g1914) & (!g3342) & (g5508) & (g5509) & (g5510)) + ((!g830) & (g1914) & (g3342) & (!g5508) & (!g5509) & (g5510)) + ((!g830) & (g1914) & (g3342) & (!g5508) & (g5509) & (g5510)) + ((!g830) & (g1914) & (g3342) & (g5508) & (!g5509) & (g5510)) + ((!g830) & (g1914) & (g3342) & (g5508) & (g5509) & (g5510)) + ((g830) & (!g1914) & (!g3342) & (!g5508) & (g5509) & (!g5510)) + ((g830) & (!g1914) & (!g3342) & (!g5508) & (g5509) & (g5510)) + ((g830) & (!g1914) & (!g3342) & (g5508) & (g5509) & (!g5510)) + ((g830) & (!g1914) & (!g3342) & (g5508) & (g5509) & (g5510)) + ((g830) & (!g1914) & (g3342) & (!g5508) & (!g5509) & (!g5510)) + ((g830) & (!g1914) & (g3342) & (!g5508) & (!g5509) & (g5510)) + ((g830) & (!g1914) & (g3342) & (g5508) & (!g5509) & (!g5510)) + ((g830) & (!g1914) & (g3342) & (g5508) & (!g5509) & (g5510)) + ((g830) & (g1914) & (!g3342) & (g5508) & (!g5509) & (!g5510)) + ((g830) & (g1914) & (!g3342) & (g5508) & (!g5509) & (g5510)) + ((g830) & (g1914) & (!g3342) & (g5508) & (g5509) & (!g5510)) + ((g830) & (g1914) & (!g3342) & (g5508) & (g5509) & (g5510)) + ((g830) & (g1914) & (g3342) & (!g5508) & (!g5509) & (!g5510)) + ((g830) & (g1914) & (g3342) & (!g5508) & (!g5509) & (g5510)) + ((g830) & (g1914) & (g3342) & (!g5508) & (g5509) & (!g5510)) + ((g830) & (g1914) & (g3342) & (!g5508) & (g5509) & (g5510)));
	assign g5512 = (((!g2468) & (!g2523) & (!g2486) & (g2544) & (!g5474)) + ((!g2468) & (!g2523) & (!g2486) & (g2544) & (g5474)) + ((!g2468) & (!g2523) & (g2486) & (!g2544) & (!g5474)) + ((!g2468) & (!g2523) & (g2486) & (g2544) & (g5474)) + ((!g2468) & (g2523) & (!g2486) & (!g2544) & (!g5474)) + ((!g2468) & (g2523) & (!g2486) & (!g2544) & (g5474)) + ((!g2468) & (g2523) & (g2486) & (!g2544) & (g5474)) + ((!g2468) & (g2523) & (g2486) & (g2544) & (!g5474)) + ((g2468) & (!g2523) & (!g2486) & (!g2544) & (!g5474)) + ((g2468) & (!g2523) & (!g2486) & (g2544) & (g5474)) + ((g2468) & (!g2523) & (g2486) & (!g2544) & (!g5474)) + ((g2468) & (!g2523) & (g2486) & (!g2544) & (g5474)) + ((g2468) & (g2523) & (!g2486) & (!g2544) & (g5474)) + ((g2468) & (g2523) & (!g2486) & (g2544) & (!g5474)) + ((g2468) & (g2523) & (g2486) & (g2544) & (!g5474)) + ((g2468) & (g2523) & (g2486) & (g2544) & (g5474)));
	assign g5513 = (((!g2434) & (!g2533) & (!g2503) & (g2539) & (!g5476)) + ((!g2434) & (!g2533) & (!g2503) & (g2539) & (g5476)) + ((!g2434) & (!g2533) & (g2503) & (!g2539) & (g5476)) + ((!g2434) & (!g2533) & (g2503) & (g2539) & (!g5476)) + ((!g2434) & (g2533) & (!g2503) & (!g2539) & (!g5476)) + ((!g2434) & (g2533) & (!g2503) & (!g2539) & (g5476)) + ((!g2434) & (g2533) & (g2503) & (!g2539) & (!g5476)) + ((!g2434) & (g2533) & (g2503) & (g2539) & (g5476)) + ((g2434) & (!g2533) & (!g2503) & (!g2539) & (g5476)) + ((g2434) & (!g2533) & (!g2503) & (g2539) & (!g5476)) + ((g2434) & (!g2533) & (g2503) & (!g2539) & (!g5476)) + ((g2434) & (!g2533) & (g2503) & (!g2539) & (g5476)) + ((g2434) & (g2533) & (!g2503) & (!g2539) & (!g5476)) + ((g2434) & (g2533) & (!g2503) & (g2539) & (g5476)) + ((g2434) & (g2533) & (g2503) & (g2539) & (!g5476)) + ((g2434) & (g2533) & (g2503) & (g2539) & (g5476)));
	assign g5514 = (((g830) & (!g1914) & (!g3345) & (!g5512) & (g5513)) + ((g830) & (!g1914) & (!g3345) & (g5512) & (g5513)) + ((g830) & (!g1914) & (g3345) & (!g5512) & (!g5513)) + ((g830) & (!g1914) & (g3345) & (g5512) & (!g5513)) + ((g830) & (g1914) & (!g3345) & (g5512) & (!g5513)) + ((g830) & (g1914) & (!g3345) & (g5512) & (g5513)) + ((g830) & (g1914) & (g3345) & (!g5512) & (!g5513)) + ((g830) & (g1914) & (g3345) & (!g5512) & (g5513)));
	assign g5515 = (((!g2299) & (!g2991) & (!g3723) & (g3724)) + ((!g2299) & (!g2991) & (g3723) & (!g3724)) + ((!g2299) & (!g2991) & (g3723) & (g3724)) + ((!g2299) & (g2991) & (!g3723) & (!g3724)) + ((g2299) & (!g2991) & (!g3723) & (!g3724)) + ((g2299) & (g2991) & (!g3723) & (g3724)) + ((g2299) & (g2991) & (g3723) & (!g3724)) + ((g2299) & (g2991) & (g3723) & (g3724)));
	assign g5516 = (((!g2962) & (!g3740) & (!g3741) & (g2938)) + ((!g2962) & (!g3740) & (g3741) & (!g2938)) + ((!g2962) & (g3740) & (!g3741) & (!g2938)) + ((!g2962) & (g3740) & (g3741) & (!g2938)) + ((g2962) & (!g3740) & (!g3741) & (!g2938)) + ((g2962) & (!g3740) & (g3741) & (g2938)) + ((g2962) & (g3740) & (!g3741) & (g2938)) + ((g2962) & (g3740) & (g3741) & (g2938)));
	assign g5517 = (((!g830) & (!g1914) & (!g3348) & (!g5515) & (!g5516) & (key[222])) + ((!g830) & (!g1914) & (!g3348) & (!g5515) & (g5516) & (key[222])) + ((!g830) & (!g1914) & (!g3348) & (g5515) & (!g5516) & (key[222])) + ((!g830) & (!g1914) & (!g3348) & (g5515) & (g5516) & (key[222])) + ((!g830) & (!g1914) & (g3348) & (!g5515) & (!g5516) & (key[222])) + ((!g830) & (!g1914) & (g3348) & (!g5515) & (g5516) & (key[222])) + ((!g830) & (!g1914) & (g3348) & (g5515) & (!g5516) & (key[222])) + ((!g830) & (!g1914) & (g3348) & (g5515) & (g5516) & (key[222])) + ((!g830) & (g1914) & (!g3348) & (!g5515) & (!g5516) & (key[222])) + ((!g830) & (g1914) & (!g3348) & (!g5515) & (g5516) & (key[222])) + ((!g830) & (g1914) & (!g3348) & (g5515) & (!g5516) & (key[222])) + ((!g830) & (g1914) & (!g3348) & (g5515) & (g5516) & (key[222])) + ((!g830) & (g1914) & (g3348) & (!g5515) & (!g5516) & (key[222])) + ((!g830) & (g1914) & (g3348) & (!g5515) & (g5516) & (key[222])) + ((!g830) & (g1914) & (g3348) & (g5515) & (!g5516) & (key[222])) + ((!g830) & (g1914) & (g3348) & (g5515) & (g5516) & (key[222])) + ((g830) & (!g1914) & (!g3348) & (!g5515) & (g5516) & (!key[222])) + ((g830) & (!g1914) & (!g3348) & (!g5515) & (g5516) & (key[222])) + ((g830) & (!g1914) & (!g3348) & (g5515) & (g5516) & (!key[222])) + ((g830) & (!g1914) & (!g3348) & (g5515) & (g5516) & (key[222])) + ((g830) & (!g1914) & (g3348) & (!g5515) & (!g5516) & (!key[222])) + ((g830) & (!g1914) & (g3348) & (!g5515) & (!g5516) & (key[222])) + ((g830) & (!g1914) & (g3348) & (g5515) & (!g5516) & (!key[222])) + ((g830) & (!g1914) & (g3348) & (g5515) & (!g5516) & (key[222])) + ((g830) & (g1914) & (!g3348) & (g5515) & (!g5516) & (!key[222])) + ((g830) & (g1914) & (!g3348) & (g5515) & (!g5516) & (key[222])) + ((g830) & (g1914) & (!g3348) & (g5515) & (g5516) & (!key[222])) + ((g830) & (g1914) & (!g3348) & (g5515) & (g5516) & (key[222])) + ((g830) & (g1914) & (g3348) & (!g5515) & (!g5516) & (!key[222])) + ((g830) & (g1914) & (g3348) & (!g5515) & (!g5516) & (key[222])) + ((g830) & (g1914) & (g3348) & (!g5515) & (g5516) & (!key[222])) + ((g830) & (g1914) & (g3348) & (!g5515) & (g5516) & (key[222])));
	assign g5518 = (((!g2099) & (!g2130) & (!g2747) & (g2780) & (!g5466)) + ((!g2099) & (!g2130) & (!g2747) & (g2780) & (g5466)) + ((!g2099) & (!g2130) & (g2747) & (!g2780) & (g5466)) + ((!g2099) & (!g2130) & (g2747) & (g2780) & (!g5466)) + ((!g2099) & (g2130) & (!g2747) & (!g2780) & (!g5466)) + ((!g2099) & (g2130) & (!g2747) & (!g2780) & (g5466)) + ((!g2099) & (g2130) & (g2747) & (!g2780) & (!g5466)) + ((!g2099) & (g2130) & (g2747) & (g2780) & (g5466)) + ((g2099) & (!g2130) & (!g2747) & (!g2780) & (g5466)) + ((g2099) & (!g2130) & (!g2747) & (g2780) & (!g5466)) + ((g2099) & (!g2130) & (g2747) & (!g2780) & (!g5466)) + ((g2099) & (!g2130) & (g2747) & (!g2780) & (g5466)) + ((g2099) & (g2130) & (!g2747) & (!g2780) & (!g5466)) + ((g2099) & (g2130) & (!g2747) & (g2780) & (g5466)) + ((g2099) & (g2130) & (g2747) & (g2780) & (!g5466)) + ((g2099) & (g2130) & (g2747) & (g2780) & (g5466)));
	assign g5519 = (((!g1914) & (!g3038) & (!g3041) & (!g3793) & (g5518)) + ((!g1914) & (!g3038) & (!g3041) & (g3793) & (g5518)) + ((!g1914) & (!g3038) & (g3041) & (!g3793) & (g5518)) + ((!g1914) & (!g3038) & (g3041) & (g3793) & (g5518)) + ((!g1914) & (g3038) & (!g3041) & (!g3793) & (g5518)) + ((!g1914) & (g3038) & (!g3041) & (g3793) & (g5518)) + ((!g1914) & (g3038) & (g3041) & (!g3793) & (g5518)) + ((!g1914) & (g3038) & (g3041) & (g3793) & (g5518)) + ((g1914) & (!g3038) & (!g3041) & (!g3793) & (!g5518)) + ((g1914) & (!g3038) & (!g3041) & (!g3793) & (g5518)) + ((g1914) & (!g3038) & (g3041) & (g3793) & (!g5518)) + ((g1914) & (!g3038) & (g3041) & (g3793) & (g5518)) + ((g1914) & (g3038) & (!g3041) & (g3793) & (!g5518)) + ((g1914) & (g3038) & (!g3041) & (g3793) & (g5518)) + ((g1914) & (g3038) & (g3041) & (!g3793) & (!g5518)) + ((g1914) & (g3038) & (g3041) & (!g3793) & (g5518)));
	assign g5520 = (((!g830) & (!g3353) & (!g5519) & (key[158])) + ((!g830) & (!g3353) & (g5519) & (key[158])) + ((!g830) & (g3353) & (!g5519) & (key[158])) + ((!g830) & (g3353) & (g5519) & (key[158])) + ((g830) & (!g3353) & (g5519) & (!key[158])) + ((g830) & (!g3353) & (g5519) & (key[158])) + ((g830) & (g3353) & (!g5519) & (!key[158])) + ((g830) & (g3353) & (!g5519) & (key[158])));
	assign g5521 = (((!g2962) & (!g2956) & (!g3824) & (g3825)) + ((!g2962) & (!g2956) & (g3824) & (!g3825)) + ((!g2962) & (!g2956) & (g3824) & (g3825)) + ((!g2962) & (g2956) & (!g3824) & (!g3825)) + ((g2962) & (!g2956) & (!g3824) & (!g3825)) + ((g2962) & (g2956) & (!g3824) & (g3825)) + ((g2962) & (g2956) & (g3824) & (!g3825)) + ((g2962) & (g2956) & (g3824) & (g3825)));
	assign g5522 = (((!g2296) & (!g2991) & (!g3841) & (g3842)) + ((!g2296) & (!g2991) & (g3841) & (!g3842)) + ((!g2296) & (!g2991) & (g3841) & (g3842)) + ((!g2296) & (g2991) & (!g3841) & (!g3842)) + ((g2296) & (!g2991) & (!g3841) & (!g3842)) + ((g2296) & (g2991) & (!g3841) & (g3842)) + ((g2296) & (g2991) & (g3841) & (!g3842)) + ((g2296) & (g2991) & (g3841) & (g3842)));
	assign g5523 = (((!g830) & (!g1914) & (!g3356) & (!g5521) & (!g5522) & (nonce[62])) + ((!g830) & (!g1914) & (!g3356) & (!g5521) & (g5522) & (nonce[62])) + ((!g830) & (!g1914) & (!g3356) & (g5521) & (!g5522) & (nonce[62])) + ((!g830) & (!g1914) & (!g3356) & (g5521) & (g5522) & (nonce[62])) + ((!g830) & (!g1914) & (g3356) & (!g5521) & (!g5522) & (nonce[62])) + ((!g830) & (!g1914) & (g3356) & (!g5521) & (g5522) & (nonce[62])) + ((!g830) & (!g1914) & (g3356) & (g5521) & (!g5522) & (nonce[62])) + ((!g830) & (!g1914) & (g3356) & (g5521) & (g5522) & (nonce[62])) + ((!g830) & (g1914) & (!g3356) & (!g5521) & (!g5522) & (nonce[62])) + ((!g830) & (g1914) & (!g3356) & (!g5521) & (g5522) & (nonce[62])) + ((!g830) & (g1914) & (!g3356) & (g5521) & (!g5522) & (nonce[62])) + ((!g830) & (g1914) & (!g3356) & (g5521) & (g5522) & (nonce[62])) + ((!g830) & (g1914) & (g3356) & (!g5521) & (!g5522) & (nonce[62])) + ((!g830) & (g1914) & (g3356) & (!g5521) & (g5522) & (nonce[62])) + ((!g830) & (g1914) & (g3356) & (g5521) & (!g5522) & (nonce[62])) + ((!g830) & (g1914) & (g3356) & (g5521) & (g5522) & (nonce[62])) + ((g830) & (!g1914) & (!g3356) & (!g5521) & (g5522) & (!nonce[62])) + ((g830) & (!g1914) & (!g3356) & (!g5521) & (g5522) & (nonce[62])) + ((g830) & (!g1914) & (!g3356) & (g5521) & (g5522) & (!nonce[62])) + ((g830) & (!g1914) & (!g3356) & (g5521) & (g5522) & (nonce[62])) + ((g830) & (!g1914) & (g3356) & (!g5521) & (!g5522) & (!nonce[62])) + ((g830) & (!g1914) & (g3356) & (!g5521) & (!g5522) & (nonce[62])) + ((g830) & (!g1914) & (g3356) & (g5521) & (!g5522) & (!nonce[62])) + ((g830) & (!g1914) & (g3356) & (g5521) & (!g5522) & (nonce[62])) + ((g830) & (g1914) & (!g3356) & (g5521) & (!g5522) & (!nonce[62])) + ((g830) & (g1914) & (!g3356) & (g5521) & (!g5522) & (nonce[62])) + ((g830) & (g1914) & (!g3356) & (g5521) & (g5522) & (!nonce[62])) + ((g830) & (g1914) & (!g3356) & (g5521) & (g5522) & (nonce[62])) + ((g830) & (g1914) & (g3356) & (!g5521) & (!g5522) & (!nonce[62])) + ((g830) & (g1914) & (g3356) & (!g5521) & (!g5522) & (nonce[62])) + ((g830) & (g1914) & (g3356) & (!g5521) & (g5522) & (!nonce[62])) + ((g830) & (g1914) & (g3356) & (!g5521) & (g5522) & (nonce[62])));
	assign g5524 = (((!g2497) & (!g2531) & (!g2503) & (g2539) & (!g5488)) + ((!g2497) & (!g2531) & (!g2503) & (g2539) & (g5488)) + ((!g2497) & (!g2531) & (g2503) & (!g2539) & (!g5488)) + ((!g2497) & (!g2531) & (g2503) & (g2539) & (g5488)) + ((!g2497) & (g2531) & (!g2503) & (!g2539) & (!g5488)) + ((!g2497) & (g2531) & (!g2503) & (!g2539) & (g5488)) + ((!g2497) & (g2531) & (g2503) & (!g2539) & (g5488)) + ((!g2497) & (g2531) & (g2503) & (g2539) & (!g5488)) + ((g2497) & (!g2531) & (!g2503) & (!g2539) & (!g5488)) + ((g2497) & (!g2531) & (!g2503) & (g2539) & (g5488)) + ((g2497) & (!g2531) & (g2503) & (!g2539) & (!g5488)) + ((g2497) & (!g2531) & (g2503) & (!g2539) & (g5488)) + ((g2497) & (g2531) & (!g2503) & (!g2539) & (g5488)) + ((g2497) & (g2531) & (!g2503) & (g2539) & (!g5488)) + ((g2497) & (g2531) & (g2503) & (g2539) & (!g5488)) + ((g2497) & (g2531) & (g2503) & (g2539) & (g5488)));
	assign g5525 = (((!g2462) & (!g2542) & (!g2486) & (g2544) & (!g5490)) + ((!g2462) & (!g2542) & (!g2486) & (g2544) & (g5490)) + ((!g2462) & (!g2542) & (g2486) & (!g2544) & (g5490)) + ((!g2462) & (!g2542) & (g2486) & (g2544) & (!g5490)) + ((!g2462) & (g2542) & (!g2486) & (!g2544) & (!g5490)) + ((!g2462) & (g2542) & (!g2486) & (!g2544) & (g5490)) + ((!g2462) & (g2542) & (g2486) & (!g2544) & (!g5490)) + ((!g2462) & (g2542) & (g2486) & (g2544) & (g5490)) + ((g2462) & (!g2542) & (!g2486) & (!g2544) & (g5490)) + ((g2462) & (!g2542) & (!g2486) & (g2544) & (!g5490)) + ((g2462) & (!g2542) & (g2486) & (!g2544) & (!g5490)) + ((g2462) & (!g2542) & (g2486) & (!g2544) & (g5490)) + ((g2462) & (g2542) & (!g2486) & (!g2544) & (!g5490)) + ((g2462) & (g2542) & (!g2486) & (g2544) & (g5490)) + ((g2462) & (g2542) & (g2486) & (g2544) & (!g5490)) + ((g2462) & (g2542) & (g2486) & (g2544) & (g5490)));
	assign g5526 = (((!g830) & (!g1914) & (!g3359) & (!g5524) & (!g5525)) + ((!g830) & (!g1914) & (!g3359) & (!g5524) & (g5525)) + ((!g830) & (!g1914) & (!g3359) & (g5524) & (!g5525)) + ((!g830) & (!g1914) & (!g3359) & (g5524) & (g5525)) + ((!g830) & (!g1914) & (g3359) & (!g5524) & (!g5525)) + ((!g830) & (!g1914) & (g3359) & (!g5524) & (g5525)) + ((!g830) & (!g1914) & (g3359) & (g5524) & (!g5525)) + ((!g830) & (!g1914) & (g3359) & (g5524) & (g5525)) + ((!g830) & (g1914) & (!g3359) & (!g5524) & (!g5525)) + ((!g830) & (g1914) & (!g3359) & (!g5524) & (g5525)) + ((!g830) & (g1914) & (!g3359) & (g5524) & (!g5525)) + ((!g830) & (g1914) & (!g3359) & (g5524) & (g5525)) + ((!g830) & (g1914) & (g3359) & (!g5524) & (!g5525)) + ((!g830) & (g1914) & (g3359) & (!g5524) & (g5525)) + ((!g830) & (g1914) & (g3359) & (g5524) & (!g5525)) + ((!g830) & (g1914) & (g3359) & (g5524) & (g5525)) + ((g830) & (!g1914) & (!g3359) & (!g5524) & (g5525)) + ((g830) & (!g1914) & (!g3359) & (g5524) & (g5525)) + ((g830) & (!g1914) & (g3359) & (!g5524) & (!g5525)) + ((g830) & (!g1914) & (g3359) & (g5524) & (!g5525)) + ((g830) & (g1914) & (!g3359) & (g5524) & (!g5525)) + ((g830) & (g1914) & (!g3359) & (g5524) & (g5525)) + ((g830) & (g1914) & (g3359) & (!g5524) & (!g5525)) + ((g830) & (g1914) & (g3359) & (!g5524) & (g5525)));
	assign g5527 = (((!g2822) & (!g3650) & (!g2816)) + ((!g2822) & (g3650) & (g2816)) + ((g2822) & (!g3650) & (g2816)) + ((g2822) & (g3650) & (!g2816)));
	assign g5528 = (((!g1914) & (!g2424) & (!g1644) & (!g3637) & (g5527)) + ((!g1914) & (!g2424) & (!g1644) & (g3637) & (g5527)) + ((!g1914) & (!g2424) & (g1644) & (!g3637) & (g5527)) + ((!g1914) & (!g2424) & (g1644) & (g3637) & (g5527)) + ((!g1914) & (g2424) & (!g1644) & (!g3637) & (g5527)) + ((!g1914) & (g2424) & (!g1644) & (g3637) & (g5527)) + ((!g1914) & (g2424) & (g1644) & (!g3637) & (g5527)) + ((!g1914) & (g2424) & (g1644) & (g3637) & (g5527)) + ((g1914) & (!g2424) & (!g1644) & (g3637) & (!g5527)) + ((g1914) & (!g2424) & (!g1644) & (g3637) & (g5527)) + ((g1914) & (!g2424) & (g1644) & (!g3637) & (!g5527)) + ((g1914) & (!g2424) & (g1644) & (!g3637) & (g5527)) + ((g1914) & (g2424) & (!g1644) & (!g3637) & (!g5527)) + ((g1914) & (g2424) & (!g1644) & (!g3637) & (g5527)) + ((g1914) & (g2424) & (g1644) & (g3637) & (!g5527)) + ((g1914) & (g2424) & (g1644) & (g3637) & (g5527)));
	assign g5529 = (((!g830) & (!g3366) & (!g5528) & (key[31])) + ((!g830) & (!g3366) & (g5528) & (key[31])) + ((!g830) & (g3366) & (!g5528) & (key[31])) + ((!g830) & (g3366) & (g5528) & (key[31])) + ((g830) & (!g3366) & (g5528) & (!key[31])) + ((g830) & (!g3366) & (g5528) & (key[31])) + ((g830) & (g3366) & (!g5528) & (!key[31])) + ((g830) & (g3366) & (!g5528) & (key[31])));
	assign g5530 = (((!g1972) & (!g2578) & (!g3553)) + ((!g1972) & (g2578) & (g3553)) + ((g1972) & (!g2578) & (g3553)) + ((g1972) & (g2578) & (!g3553)));
	assign g5531 = (((!g2180) & (!g2827) & (!g3666)) + ((!g2180) & (g2827) & (g3666)) + ((g2180) & (!g2827) & (g3666)) + ((g2180) & (g2827) & (!g3666)));
	assign g5532 = (((!g1914) & (!g3088) & (!g3685) & (g3084) & (!g5531)) + ((!g1914) & (!g3088) & (!g3685) & (g3084) & (g5531)) + ((!g1914) & (!g3088) & (g3685) & (!g3084) & (!g5531)) + ((!g1914) & (!g3088) & (g3685) & (!g3084) & (g5531)) + ((!g1914) & (g3088) & (!g3685) & (!g3084) & (!g5531)) + ((!g1914) & (g3088) & (!g3685) & (!g3084) & (g5531)) + ((!g1914) & (g3088) & (g3685) & (g3084) & (!g5531)) + ((!g1914) & (g3088) & (g3685) & (g3084) & (g5531)) + ((g1914) & (!g3088) & (!g3685) & (!g3084) & (g5531)) + ((g1914) & (!g3088) & (!g3685) & (g3084) & (g5531)) + ((g1914) & (!g3088) & (g3685) & (!g3084) & (g5531)) + ((g1914) & (!g3088) & (g3685) & (g3084) & (g5531)) + ((g1914) & (g3088) & (!g3685) & (!g3084) & (g5531)) + ((g1914) & (g3088) & (!g3685) & (g3084) & (g5531)) + ((g1914) & (g3088) & (g3685) & (!g3084) & (g5531)) + ((g1914) & (g3088) & (g3685) & (g3084) & (g5531)));
	assign g8339 = (((!g5560) & (g5647) & (!g5533)) + ((!g5560) & (g5647) & (g5533)) + ((g5560) & (!g5647) & (g5533)) + ((g5560) & (g5647) & (g5533)));
	assign g5534 = (((!g830) & (!g3372) & (!g5532) & (g5533)) + ((!g830) & (!g3372) & (g5532) & (g5533)) + ((!g830) & (g3372) & (!g5532) & (g5533)) + ((!g830) & (g3372) & (g5532) & (g5533)) + ((g830) & (!g3372) & (g5532) & (!g5533)) + ((g830) & (!g3372) & (g5532) & (g5533)) + ((g830) & (g3372) & (!g5532) & (!g5533)) + ((g830) & (g3372) & (!g5532) & (g5533)));
	assign g5535 = (((!g2178) & (!g2830) & (!g3807)) + ((!g2178) & (g2830) & (g3807)) + ((g2178) & (!g2830) & (g3807)) + ((g2178) & (g2830) & (!g3807)));
	assign g5536 = (((!g1914) & (!g3078) & (!g3794) & (!g3086) & (g5535)) + ((!g1914) & (!g3078) & (!g3794) & (g3086) & (g5535)) + ((!g1914) & (!g3078) & (g3794) & (!g3086) & (g5535)) + ((!g1914) & (!g3078) & (g3794) & (g3086) & (g5535)) + ((!g1914) & (g3078) & (!g3794) & (!g3086) & (g5535)) + ((!g1914) & (g3078) & (!g3794) & (g3086) & (g5535)) + ((!g1914) & (g3078) & (g3794) & (!g3086) & (g5535)) + ((!g1914) & (g3078) & (g3794) & (g3086) & (g5535)) + ((g1914) & (!g3078) & (!g3794) & (g3086) & (!g5535)) + ((g1914) & (!g3078) & (!g3794) & (g3086) & (g5535)) + ((g1914) & (!g3078) & (g3794) & (!g3086) & (!g5535)) + ((g1914) & (!g3078) & (g3794) & (!g3086) & (g5535)) + ((g1914) & (g3078) & (!g3794) & (!g3086) & (!g5535)) + ((g1914) & (g3078) & (!g3794) & (!g3086) & (g5535)) + ((g1914) & (g3078) & (g3794) & (g3086) & (!g5535)) + ((g1914) & (g3078) & (g3794) & (g3086) & (g5535)));
	assign g5537 = (((!g830) & (!g3374) & (!g5536) & (key[159])) + ((!g830) & (!g3374) & (g5536) & (key[159])) + ((!g830) & (g3374) & (!g5536) & (key[159])) + ((!g830) & (g3374) & (g5536) & (key[159])) + ((g830) & (!g3374) & (g5536) & (!key[159])) + ((g830) & (!g3374) & (g5536) & (key[159])) + ((g830) & (g3374) & (!g5536) & (!key[159])) + ((g830) & (g3374) & (!g5536) & (key[159])));
	assign g5538 = (((!g3442) & (!g2807) & (!g2830)) + ((!g3442) & (g2807) & (g2830)) + ((g3442) & (!g2807) & (g2830)) + ((g3442) & (g2807) & (!g2830)));
	assign g5539 = (((!g1914) & (!g2427) & (!g1644) & (g3460) & (!g5538)) + ((!g1914) & (!g2427) & (!g1644) & (g3460) & (g5538)) + ((!g1914) & (!g2427) & (g1644) & (!g3460) & (!g5538)) + ((!g1914) & (!g2427) & (g1644) & (!g3460) & (g5538)) + ((!g1914) & (g2427) & (!g1644) & (!g3460) & (!g5538)) + ((!g1914) & (g2427) & (!g1644) & (!g3460) & (g5538)) + ((!g1914) & (g2427) & (g1644) & (g3460) & (!g5538)) + ((!g1914) & (g2427) & (g1644) & (g3460) & (g5538)) + ((g1914) & (!g2427) & (!g1644) & (!g3460) & (g5538)) + ((g1914) & (!g2427) & (!g1644) & (g3460) & (g5538)) + ((g1914) & (!g2427) & (g1644) & (!g3460) & (g5538)) + ((g1914) & (!g2427) & (g1644) & (g3460) & (g5538)) + ((g1914) & (g2427) & (!g1644) & (!g3460) & (g5538)) + ((g1914) & (g2427) & (!g1644) & (g3460) & (g5538)) + ((g1914) & (g2427) & (g1644) & (!g3460) & (g5538)) + ((g1914) & (g2427) & (g1644) & (g3460) & (g5538)));
	assign g5540 = (((!g830) & (!g3376) & (!g5539) & (key[127])) + ((!g830) & (!g3376) & (g5539) & (key[127])) + ((!g830) & (g3376) & (!g5539) & (key[127])) + ((!g830) & (g3376) & (g5539) & (key[127])) + ((g830) & (!g3376) & (g5539) & (!key[127])) + ((g830) & (!g3376) & (g5539) & (key[127])) + ((g830) & (g3376) & (!g5539) & (!key[127])) + ((g830) & (g3376) & (!g5539) & (key[127])));
	assign g5541 = (((!g2177) & (!g2810) & (!g3584)) + ((!g2177) & (g2810) & (g3584)) + ((g2177) & (!g2810) & (g3584)) + ((g2177) & (g2810) & (!g3584)));
	assign g5542 = (((!g1914) & (!g3571) & (!g3074) & (!g3088) & (g5541)) + ((!g1914) & (!g3571) & (!g3074) & (g3088) & (g5541)) + ((!g1914) & (!g3571) & (g3074) & (!g3088) & (g5541)) + ((!g1914) & (!g3571) & (g3074) & (g3088) & (g5541)) + ((!g1914) & (g3571) & (!g3074) & (!g3088) & (g5541)) + ((!g1914) & (g3571) & (!g3074) & (g3088) & (g5541)) + ((!g1914) & (g3571) & (g3074) & (!g3088) & (g5541)) + ((!g1914) & (g3571) & (g3074) & (g3088) & (g5541)) + ((g1914) & (!g3571) & (!g3074) & (g3088) & (!g5541)) + ((g1914) & (!g3571) & (!g3074) & (g3088) & (g5541)) + ((g1914) & (!g3571) & (g3074) & (!g3088) & (!g5541)) + ((g1914) & (!g3571) & (g3074) & (!g3088) & (g5541)) + ((g1914) & (g3571) & (!g3074) & (!g3088) & (!g5541)) + ((g1914) & (g3571) & (!g3074) & (!g3088) & (g5541)) + ((g1914) & (g3571) & (g3074) & (g3088) & (!g5541)) + ((g1914) & (g3571) & (g3074) & (g3088) & (g5541)));
	assign g5543 = (((!g830) & (!g3378) & (!g5542) & (nonce[31])) + ((!g830) & (!g3378) & (g5542) & (nonce[31])) + ((!g830) & (g3378) & (!g5542) & (nonce[31])) + ((!g830) & (g3378) & (g5542) & (nonce[31])) + ((g830) & (!g3378) & (g5542) & (!nonce[31])) + ((g830) & (!g3378) & (g5542) & (nonce[31])) + ((g830) & (g3378) & (!g5542) & (!nonce[31])) + ((g830) & (g3378) & (!g5542) & (nonce[31])));
	assign g5544 = (((!g2559) & (!g2592) & (!g3708)) + ((!g2559) & (g2592) & (g3708)) + ((g2559) & (!g2592) & (g3708)) + ((g2559) & (g2592) & (!g3708)));
	assign g5545 = (((!g2962) & (!g2956) & (!g3824) & (!g3825)) + ((!g2962) & (!g2956) & (!g3824) & (g3825)) + ((!g2962) & (!g2956) & (g3824) & (!g3825)) + ((!g2962) & (!g2956) & (g3824) & (g3825)) + ((!g2962) & (g2956) & (!g3824) & (!g3825)) + ((g2962) & (!g2956) & (!g3824) & (!g3825)));
	assign g5546 = (((g1914) & (!g3013) & (!g3005) & (!g5545)) + ((g1914) & (!g3013) & (g3005) & (g5545)) + ((g1914) & (g3013) & (!g3005) & (g5545)) + ((g1914) & (g3013) & (g3005) & (!g5545)));
	assign g5547 = (((!g2296) & (!g2991) & (!g3841) & (!g3842)) + ((!g2296) & (!g2991) & (!g3841) & (g3842)) + ((!g2296) & (!g2991) & (g3841) & (!g3842)) + ((!g2296) & (!g2991) & (g3841) & (g3842)) + ((!g2296) & (g2991) & (!g3841) & (!g3842)) + ((g2296) & (!g2991) & (!g3841) & (!g3842)));
	assign g5548 = (((!g1914) & (!g2344) & (!g3022) & (!g5547)) + ((!g1914) & (!g2344) & (g3022) & (g5547)) + ((!g1914) & (g2344) & (!g3022) & (g5547)) + ((!g1914) & (g2344) & (g3022) & (!g5547)));
	assign g5549 = (((!g830) & (!g3382) & (!g5546) & (!g5548) & (nonce[63])) + ((!g830) & (!g3382) & (!g5546) & (g5548) & (nonce[63])) + ((!g830) & (!g3382) & (g5546) & (!g5548) & (nonce[63])) + ((!g830) & (!g3382) & (g5546) & (g5548) & (nonce[63])) + ((!g830) & (g3382) & (!g5546) & (!g5548) & (nonce[63])) + ((!g830) & (g3382) & (!g5546) & (g5548) & (nonce[63])) + ((!g830) & (g3382) & (g5546) & (!g5548) & (nonce[63])) + ((!g830) & (g3382) & (g5546) & (g5548) & (nonce[63])) + ((g830) & (!g3382) & (!g5546) & (g5548) & (!nonce[63])) + ((g830) & (!g3382) & (!g5546) & (g5548) & (nonce[63])) + ((g830) & (!g3382) & (g5546) & (!g5548) & (!nonce[63])) + ((g830) & (!g3382) & (g5546) & (!g5548) & (nonce[63])) + ((g830) & (!g3382) & (g5546) & (g5548) & (!nonce[63])) + ((g830) & (!g3382) & (g5546) & (g5548) & (nonce[63])) + ((g830) & (g3382) & (!g5546) & (!g5548) & (!nonce[63])) + ((g830) & (g3382) & (!g5546) & (!g5548) & (nonce[63])));
	assign g5550 = (((!g2181) & (!g3600) & (!g2822)) + ((!g2181) & (g3600) & (g2822)) + ((g2181) & (!g3600) & (g2822)) + ((g2181) & (g3600) & (!g2822)));
	assign g5551 = (((!g1914) & (!g3618) & (!g3078) & (g3080) & (!g5550)) + ((!g1914) & (!g3618) & (!g3078) & (g3080) & (g5550)) + ((!g1914) & (!g3618) & (g3078) & (!g3080) & (!g5550)) + ((!g1914) & (!g3618) & (g3078) & (!g3080) & (g5550)) + ((!g1914) & (g3618) & (!g3078) & (!g3080) & (!g5550)) + ((!g1914) & (g3618) & (!g3078) & (!g3080) & (g5550)) + ((!g1914) & (g3618) & (g3078) & (g3080) & (!g5550)) + ((!g1914) & (g3618) & (g3078) & (g3080) & (g5550)) + ((g1914) & (!g3618) & (!g3078) & (!g3080) & (g5550)) + ((g1914) & (!g3618) & (!g3078) & (g3080) & (g5550)) + ((g1914) & (!g3618) & (g3078) & (!g3080) & (g5550)) + ((g1914) & (!g3618) & (g3078) & (g3080) & (g5550)) + ((g1914) & (g3618) & (!g3078) & (!g3080) & (g5550)) + ((g1914) & (g3618) & (!g3078) & (g3080) & (g5550)) + ((g1914) & (g3618) & (g3078) & (!g3080) & (g5550)) + ((g1914) & (g3618) & (g3078) & (g3080) & (g5550)));
	assign g5552 = (((!g830) & (!g3385) & (!g5551) & (key[255])) + ((!g830) & (!g3385) & (g5551) & (key[255])) + ((!g830) & (g3385) & (!g5551) & (key[255])) + ((!g830) & (g3385) & (g5551) & (key[255])) + ((g830) & (!g3385) & (g5551) & (!key[255])) + ((g830) & (!g3385) & (g5551) & (key[255])) + ((g830) & (g3385) & (!g5551) & (!key[255])) + ((g830) & (g3385) & (!g5551) & (key[255])));
	assign g5553 = (((!g2299) & (!g2991) & (!g3723) & (!g3724)) + ((!g2299) & (!g2991) & (!g3723) & (g3724)) + ((!g2299) & (!g2991) & (g3723) & (!g3724)) + ((!g2299) & (!g2991) & (g3723) & (g3724)) + ((!g2299) & (g2991) & (!g3723) & (!g3724)) + ((g2299) & (!g2991) & (!g3723) & (!g3724)));
	assign g5554 = (((g1914) & (!g2348) & (!g3022) & (!g5553)) + ((g1914) & (!g2348) & (g3022) & (g5553)) + ((g1914) & (g2348) & (!g3022) & (g5553)) + ((g1914) & (g2348) & (g3022) & (!g5553)));
	assign g5555 = (((!g2962) & (!g3740) & (!g3741) & (!g2938)) + ((!g2962) & (!g3740) & (!g3741) & (g2938)) + ((!g2962) & (!g3740) & (g3741) & (!g2938)) + ((!g2962) & (g3740) & (!g3741) & (!g2938)) + ((!g2962) & (g3740) & (g3741) & (!g2938)) + ((g2962) & (!g3740) & (!g3741) & (!g2938)));
	assign g5556 = (((!g1914) & (!g3013) & (!g5555) & (!g3011)) + ((!g1914) & (!g3013) & (g5555) & (g3011)) + ((!g1914) & (g3013) & (!g5555) & (g3011)) + ((!g1914) & (g3013) & (g5555) & (!g3011)));
	assign g5557 = (((!g830) & (!g3387) & (!g5554) & (!g5556) & (key[223])) + ((!g830) & (!g3387) & (!g5554) & (g5556) & (key[223])) + ((!g830) & (!g3387) & (g5554) & (!g5556) & (key[223])) + ((!g830) & (!g3387) & (g5554) & (g5556) & (key[223])) + ((!g830) & (g3387) & (!g5554) & (!g5556) & (key[223])) + ((!g830) & (g3387) & (!g5554) & (g5556) & (key[223])) + ((!g830) & (g3387) & (g5554) & (!g5556) & (key[223])) + ((!g830) & (g3387) & (g5554) & (g5556) & (key[223])) + ((g830) & (!g3387) & (!g5554) & (g5556) & (!key[223])) + ((g830) & (!g3387) & (!g5554) & (g5556) & (key[223])) + ((g830) & (!g3387) & (g5554) & (!g5556) & (!key[223])) + ((g830) & (!g3387) & (g5554) & (!g5556) & (key[223])) + ((g830) & (!g3387) & (g5554) & (g5556) & (!key[223])) + ((g830) & (!g3387) & (g5554) & (g5556) & (key[223])) + ((g830) & (g3387) & (!g5554) & (!g5556) & (!key[223])) + ((g830) & (g3387) & (!g5554) & (!g5556) & (key[223])));
	assign g5558 = (((!g2572) & (!g2584) & (!g3865)) + ((!g2572) & (g2584) & (g3865)) + ((g2572) & (!g2584) & (g3865)) + ((g2572) & (g2584) & (!g3865)));
	assign g5559 = (((g827) & (!g3427)));
	assign g5560 = (((!reset) & (!g830) & (g831)) + ((!reset) & (g830) & (!g831)) + ((!reset) & (g830) & (g831)) + ((reset) & (!g830) & (!g831)) + ((reset) & (!g830) & (g831)) + ((reset) & (g830) & (!g831)) + ((reset) & (g830) & (g831)));
	assign g5561 = (((g3427) & (g4000) & (g4010) & (g4027) & (g4036)));
	assign g5562 = (((g4046) & (g4053) & (g4060) & (g5561)));
	assign g5563 = (((g4068) & (g4075) & (g4083) & (g4046) & (g5561) & (g5716)));
	assign g5564 = (((g4091) & (g4098) & (g4104) & (g4110) & (g4177) & (g5563)));
	assign g5565 = (((g4252) & (g4315) & (g4377) & (g4426) & (g4482) & (g5564)));
	assign g5566 = (((g4545) & (g4596) & (g4649) & (g4696) & (g4749) & (g5565)));
	assign g5567 = (((g4784) & (g4835) & (g4877) & (g4931) & (g4987) & (g5566)));
	assign g5568 = (((g5033) & (g5567)));
	assign g5569 = (((g827) & (!g3687) & (g5568)) + ((g827) & (g3687) & (!g5568)));
	assign g5570 = (((g827) & (!g3427) & (g4000)) + ((g827) & (g3427) & (!g4000)));
	assign g5571 = (((g827) & (!g3427) & (!g4000) & (g4010)) + ((g827) & (!g3427) & (g4000) & (g4010)) + ((g827) & (g3427) & (!g4000) & (g4010)) + ((g827) & (g3427) & (g4000) & (!g4010)));
	assign g5572 = (((g827) & (!g3427) & (!g4000) & (!g4010) & (g4027)) + ((g827) & (!g3427) & (!g4000) & (g4010) & (g4027)) + ((g827) & (!g3427) & (g4000) & (!g4010) & (g4027)) + ((g827) & (!g3427) & (g4000) & (g4010) & (g4027)) + ((g827) & (g3427) & (!g4000) & (!g4010) & (g4027)) + ((g827) & (g3427) & (!g4000) & (g4010) & (g4027)) + ((g827) & (g3427) & (g4000) & (!g4010) & (g4027)) + ((g827) & (g3427) & (g4000) & (g4010) & (!g4027)));
	assign g5573 = (((g827) & (!g3427) & (!g4000) & (!g4010) & (!g4027) & (g4036)) + ((g827) & (!g3427) & (!g4000) & (!g4010) & (g4027) & (g4036)) + ((g827) & (!g3427) & (!g4000) & (g4010) & (!g4027) & (g4036)) + ((g827) & (!g3427) & (!g4000) & (g4010) & (g4027) & (g4036)) + ((g827) & (!g3427) & (g4000) & (!g4010) & (!g4027) & (g4036)) + ((g827) & (!g3427) & (g4000) & (!g4010) & (g4027) & (g4036)) + ((g827) & (!g3427) & (g4000) & (g4010) & (!g4027) & (g4036)) + ((g827) & (!g3427) & (g4000) & (g4010) & (g4027) & (g4036)) + ((g827) & (g3427) & (!g4000) & (!g4010) & (!g4027) & (g4036)) + ((g827) & (g3427) & (!g4000) & (!g4010) & (g4027) & (g4036)) + ((g827) & (g3427) & (!g4000) & (g4010) & (!g4027) & (g4036)) + ((g827) & (g3427) & (!g4000) & (g4010) & (g4027) & (g4036)) + ((g827) & (g3427) & (g4000) & (!g4010) & (!g4027) & (g4036)) + ((g827) & (g3427) & (g4000) & (!g4010) & (g4027) & (g4036)) + ((g827) & (g3427) & (g4000) & (g4010) & (!g4027) & (g4036)) + ((g827) & (g3427) & (g4000) & (g4010) & (g4027) & (!g4036)));
	assign g5574 = (((g827) & (!g4046) & (g5561)) + ((g827) & (g4046) & (!g5561)));
	assign g5575 = (((g827) & (!g4046) & (g4053) & (!g5561)) + ((g827) & (!g4046) & (g4053) & (g5561)) + ((g827) & (g4046) & (!g4053) & (g5561)) + ((g827) & (g4046) & (g4053) & (!g5561)));
	assign g5576 = (((g827) & (!g4046) & (!g4053) & (g4060) & (!g5561)) + ((g827) & (!g4046) & (!g4053) & (g4060) & (g5561)) + ((g827) & (!g4046) & (g4053) & (g4060) & (!g5561)) + ((g827) & (!g4046) & (g4053) & (g4060) & (g5561)) + ((g827) & (g4046) & (!g4053) & (g4060) & (!g5561)) + ((g827) & (g4046) & (!g4053) & (g4060) & (g5561)) + ((g827) & (g4046) & (g4053) & (!g4060) & (g5561)) + ((g827) & (g4046) & (g4053) & (g4060) & (!g5561)));
	assign g5577 = (((g827) & (!g4068) & (g5562)) + ((g827) & (g4068) & (!g5562)));
	assign g5578 = (((g827) & (!g4068) & (g4075) & (!g5562)) + ((g827) & (!g4068) & (g4075) & (g5562)) + ((g827) & (g4068) & (!g4075) & (g5562)) + ((g827) & (g4068) & (g4075) & (!g5562)));
	assign g5579 = (((g827) & (!g4068) & (!g4075) & (g4083) & (!g5562)) + ((g827) & (!g4068) & (!g4075) & (g4083) & (g5562)) + ((g827) & (!g4068) & (g4075) & (g4083) & (!g5562)) + ((g827) & (!g4068) & (g4075) & (g4083) & (g5562)) + ((g827) & (g4068) & (!g4075) & (g4083) & (!g5562)) + ((g827) & (g4068) & (!g4075) & (g4083) & (g5562)) + ((g827) & (g4068) & (g4075) & (!g4083) & (g5562)) + ((g827) & (g4068) & (g4075) & (g4083) & (!g5562)));
	assign g5580 = (((g827) & (!g4091) & (g5563)) + ((g827) & (g4091) & (!g5563)));
	assign g5581 = (((g827) & (!g4091) & (g4098) & (!g5563)) + ((g827) & (!g4091) & (g4098) & (g5563)) + ((g827) & (g4091) & (!g4098) & (g5563)) + ((g827) & (g4091) & (g4098) & (!g5563)));
	assign g5582 = (((g827) & (!g4091) & (!g4098) & (g4104) & (!g5563)) + ((g827) & (!g4091) & (!g4098) & (g4104) & (g5563)) + ((g827) & (!g4091) & (g4098) & (g4104) & (!g5563)) + ((g827) & (!g4091) & (g4098) & (g4104) & (g5563)) + ((g827) & (g4091) & (!g4098) & (g4104) & (!g5563)) + ((g827) & (g4091) & (!g4098) & (g4104) & (g5563)) + ((g827) & (g4091) & (g4098) & (!g4104) & (g5563)) + ((g827) & (g4091) & (g4098) & (g4104) & (!g5563)));
	assign g5583 = (((g4091) & (g4098) & (g4104) & (g5563)));
	assign g5584 = (((g827) & (!g4110) & (g5583)) + ((g827) & (g4110) & (!g5583)));
	assign g5585 = (((g827) & (!g3687) & (g4127) & (!g5568)) + ((g827) & (!g3687) & (g4127) & (g5568)) + ((g827) & (g3687) & (!g4127) & (g5568)) + ((g827) & (g3687) & (g4127) & (!g5568)));
	assign g5586 = (((g827) & (!g4110) & (g4177) & (!g5583)) + ((g827) & (!g4110) & (g4177) & (g5583)) + ((g827) & (g4110) & (!g4177) & (g5583)) + ((g827) & (g4110) & (g4177) & (!g5583)));
	assign g5587 = (((g827) & (!g3687) & (!g4127) & (g4221) & (!g5568)) + ((g827) & (!g3687) & (!g4127) & (g4221) & (g5568)) + ((g827) & (!g3687) & (g4127) & (g4221) & (!g5568)) + ((g827) & (!g3687) & (g4127) & (g4221) & (g5568)) + ((g827) & (g3687) & (!g4127) & (g4221) & (!g5568)) + ((g827) & (g3687) & (!g4127) & (g4221) & (g5568)) + ((g827) & (g3687) & (g4127) & (!g4221) & (g5568)) + ((g827) & (g3687) & (g4127) & (g4221) & (!g5568)));
	assign g5588 = (((g827) & (!g4252) & (g5564)) + ((g827) & (g4252) & (!g5564)));
	assign g5589 = (((g827) & (!g3687) & (!g4127) & (!g4221) & (g4267) & (!g5568)) + ((g827) & (!g3687) & (!g4127) & (!g4221) & (g4267) & (g5568)) + ((g827) & (!g3687) & (!g4127) & (g4221) & (g4267) & (!g5568)) + ((g827) & (!g3687) & (!g4127) & (g4221) & (g4267) & (g5568)) + ((g827) & (!g3687) & (g4127) & (!g4221) & (g4267) & (!g5568)) + ((g827) & (!g3687) & (g4127) & (!g4221) & (g4267) & (g5568)) + ((g827) & (!g3687) & (g4127) & (g4221) & (g4267) & (!g5568)) + ((g827) & (!g3687) & (g4127) & (g4221) & (g4267) & (g5568)) + ((g827) & (g3687) & (!g4127) & (!g4221) & (g4267) & (!g5568)) + ((g827) & (g3687) & (!g4127) & (!g4221) & (g4267) & (g5568)) + ((g827) & (g3687) & (!g4127) & (g4221) & (g4267) & (!g5568)) + ((g827) & (g3687) & (!g4127) & (g4221) & (g4267) & (g5568)) + ((g827) & (g3687) & (g4127) & (!g4221) & (g4267) & (!g5568)) + ((g827) & (g3687) & (g4127) & (!g4221) & (g4267) & (g5568)) + ((g827) & (g3687) & (g4127) & (g4221) & (!g4267) & (g5568)) + ((g827) & (g3687) & (g4127) & (g4221) & (g4267) & (!g5568)));
	assign g5590 = (((g4252) & (g5564)));
	assign g5591 = (((g827) & (!g4315) & (g5590)) + ((g827) & (g4315) & (!g5590)));
	assign g5592 = (((g3687) & (g4127) & (g4221) & (g4267) & (g5033) & (g5567)));
	assign g5593 = (((g827) & (!g4342) & (g5592)) + ((g827) & (g4342) & (!g5592)));
	assign g5594 = (((g827) & (!g4315) & (g4377) & (!g5590)) + ((g827) & (!g4315) & (g4377) & (g5590)) + ((g827) & (g4315) & (!g4377) & (g5590)) + ((g827) & (g4315) & (g4377) & (!g5590)));
	assign g5595 = (((g827) & (!g4342) & (g4390) & (!g5592)) + ((g827) & (!g4342) & (g4390) & (g5592)) + ((g827) & (g4342) & (!g4390) & (g5592)) + ((g827) & (g4342) & (g4390) & (!g5592)));
	assign g5596 = (((g827) & (!g4315) & (!g4377) & (g4426) & (!g5590)) + ((g827) & (!g4315) & (!g4377) & (g4426) & (g5590)) + ((g827) & (!g4315) & (g4377) & (g4426) & (!g5590)) + ((g827) & (!g4315) & (g4377) & (g4426) & (g5590)) + ((g827) & (g4315) & (!g4377) & (g4426) & (!g5590)) + ((g827) & (g4315) & (!g4377) & (g4426) & (g5590)) + ((g827) & (g4315) & (g4377) & (!g4426) & (g5590)) + ((g827) & (g4315) & (g4377) & (g4426) & (!g5590)));
	assign g5597 = (((g4342) & (g4390) & (g5592)));
	assign g5598 = (((g827) & (!g4451) & (g5597)) + ((g827) & (g4451) & (!g5597)));
	assign g5599 = (((g827) & (!g4315) & (!g4377) & (!g4426) & (g4482) & (!g5590)) + ((g827) & (!g4315) & (!g4377) & (!g4426) & (g4482) & (g5590)) + ((g827) & (!g4315) & (!g4377) & (g4426) & (g4482) & (!g5590)) + ((g827) & (!g4315) & (!g4377) & (g4426) & (g4482) & (g5590)) + ((g827) & (!g4315) & (g4377) & (!g4426) & (g4482) & (!g5590)) + ((g827) & (!g4315) & (g4377) & (!g4426) & (g4482) & (g5590)) + ((g827) & (!g4315) & (g4377) & (g4426) & (g4482) & (!g5590)) + ((g827) & (!g4315) & (g4377) & (g4426) & (g4482) & (g5590)) + ((g827) & (g4315) & (!g4377) & (!g4426) & (g4482) & (!g5590)) + ((g827) & (g4315) & (!g4377) & (!g4426) & (g4482) & (g5590)) + ((g827) & (g4315) & (!g4377) & (g4426) & (g4482) & (!g5590)) + ((g827) & (g4315) & (!g4377) & (g4426) & (g4482) & (g5590)) + ((g827) & (g4315) & (g4377) & (!g4426) & (g4482) & (!g5590)) + ((g827) & (g4315) & (g4377) & (!g4426) & (g4482) & (g5590)) + ((g827) & (g4315) & (g4377) & (g4426) & (!g4482) & (g5590)) + ((g827) & (g4315) & (g4377) & (g4426) & (g4482) & (!g5590)));
	assign g5600 = (((g827) & (!g4451) & (g4501) & (!g5597)) + ((g827) & (!g4451) & (g4501) & (g5597)) + ((g827) & (g4451) & (!g4501) & (g5597)) + ((g827) & (g4451) & (g4501) & (!g5597)));
	assign g5601 = (((g827) & (!g4545) & (g5565)) + ((g827) & (g4545) & (!g5565)));
	assign g5602 = (((g827) & (!g4451) & (!g4501) & (g4572) & (!g5597)) + ((g827) & (!g4451) & (!g4501) & (g4572) & (g5597)) + ((g827) & (!g4451) & (g4501) & (g4572) & (!g5597)) + ((g827) & (!g4451) & (g4501) & (g4572) & (g5597)) + ((g827) & (g4451) & (!g4501) & (g4572) & (!g5597)) + ((g827) & (g4451) & (!g4501) & (g4572) & (g5597)) + ((g827) & (g4451) & (g4501) & (!g4572) & (g5597)) + ((g827) & (g4451) & (g4501) & (g4572) & (!g5597)));
	assign g5603 = (((g827) & (!g4545) & (g4596) & (!g5565)) + ((g827) & (!g4545) & (g4596) & (g5565)) + ((g827) & (g4545) & (!g4596) & (g5565)) + ((g827) & (g4545) & (g4596) & (!g5565)));
	assign g5604 = (((g4342) & (g4390) & (g4451) & (g4501) & (g4572) & (g5592)));
	assign g5605 = (((g827) & (!g4610) & (g5604)) + ((g827) & (g4610) & (!g5604)));
	assign g5606 = (((g4545) & (g4596) & (g5565)));
	assign g5607 = (((g827) & (!g4649) & (g5606)) + ((g827) & (g4649) & (!g5606)));
	assign g5608 = (((g827) & (!g4610) & (g4672) & (!g5604)) + ((g827) & (!g4610) & (g4672) & (g5604)) + ((g827) & (g4610) & (!g4672) & (g5604)) + ((g827) & (g4610) & (g4672) & (!g5604)));
	assign g5609 = (((g827) & (!g4649) & (g4696) & (!g5606)) + ((g827) & (!g4649) & (g4696) & (g5606)) + ((g827) & (g4649) & (!g4696) & (g5606)) + ((g827) & (g4649) & (g4696) & (!g5606)));
	assign g5610 = (((g827) & (!g4610) & (!g4672) & (g4709) & (!g5604)) + ((g827) & (!g4610) & (!g4672) & (g4709) & (g5604)) + ((g827) & (!g4610) & (g4672) & (g4709) & (!g5604)) + ((g827) & (!g4610) & (g4672) & (g4709) & (g5604)) + ((g827) & (g4610) & (!g4672) & (g4709) & (!g5604)) + ((g827) & (g4610) & (!g4672) & (g4709) & (g5604)) + ((g827) & (g4610) & (g4672) & (!g4709) & (g5604)) + ((g827) & (g4610) & (g4672) & (g4709) & (!g5604)));
	assign g5611 = (((g827) & (!g4649) & (!g4696) & (g4749) & (!g5606)) + ((g827) & (!g4649) & (!g4696) & (g4749) & (g5606)) + ((g827) & (!g4649) & (g4696) & (g4749) & (!g5606)) + ((g827) & (!g4649) & (g4696) & (g4749) & (g5606)) + ((g827) & (g4649) & (!g4696) & (g4749) & (!g5606)) + ((g827) & (g4649) & (!g4696) & (g4749) & (g5606)) + ((g827) & (g4649) & (g4696) & (!g4749) & (g5606)) + ((g827) & (g4649) & (g4696) & (g4749) & (!g5606)));
	assign g5612 = (((g4610) & (g4672) & (g4709) & (g5604)));
	assign g5613 = (((g827) & (!g4759) & (g5612)) + ((g827) & (g4759) & (!g5612)));
	assign g5614 = (((g827) & (!g4784) & (g5566)) + ((g827) & (g4784) & (!g5566)));
	assign g5615 = (((g827) & (!g4759) & (g4798) & (!g5612)) + ((g827) & (!g4759) & (g4798) & (g5612)) + ((g827) & (g4759) & (!g4798) & (g5612)) + ((g827) & (g4759) & (g4798) & (!g5612)));
	assign g5616 = (((g4784) & (g5566)));
	assign g5617 = (((g827) & (!g4835) & (g5616)) + ((g827) & (g4835) & (!g5616)));
	assign g5618 = (((g4610) & (g4672) & (g4709) & (g4759) & (g4798) & (g5604)));
	assign g5619 = (((g827) & (!g4850) & (g5618)) + ((g827) & (g4850) & (!g5618)));
	assign g5620 = (((g827) & (!g4835) & (g4877) & (!g5616)) + ((g827) & (!g4835) & (g4877) & (g5616)) + ((g827) & (g4835) & (!g4877) & (g5616)) + ((g827) & (g4835) & (g4877) & (!g5616)));
	assign g5621 = (((g4850) & (g5618)));
	assign g5622 = (((g827) & (!g4892) & (g5621)) + ((g827) & (g4892) & (!g5621)));
	assign g5623 = (((g4835) & (g4877) & (g5616)));
	assign g5624 = (((g827) & (!g4931) & (g5623)) + ((g827) & (g4931) & (!g5623)));
	assign g5625 = (((g827) & (!g4892) & (g4959) & (!g5621)) + ((g827) & (!g4892) & (g4959) & (g5621)) + ((g827) & (g4892) & (!g4959) & (g5621)) + ((g827) & (g4892) & (g4959) & (!g5621)));
	assign g5626 = (((g827) & (!g4931) & (g4987) & (!g5623)) + ((g827) & (!g4931) & (g4987) & (g5623)) + ((g827) & (g4931) & (!g4987) & (g5623)) + ((g827) & (g4931) & (g4987) & (!g5623)));
	assign g5627 = (((g827) & (!g4892) & (!g4959) & (g4999) & (!g5621)) + ((g827) & (!g4892) & (!g4959) & (g4999) & (g5621)) + ((g827) & (!g4892) & (g4959) & (g4999) & (!g5621)) + ((g827) & (!g4892) & (g4959) & (g4999) & (g5621)) + ((g827) & (g4892) & (!g4959) & (g4999) & (!g5621)) + ((g827) & (g4892) & (!g4959) & (g4999) & (g5621)) + ((g827) & (g4892) & (g4959) & (!g4999) & (g5621)) + ((g827) & (g4892) & (g4959) & (g4999) & (!g5621)));
	assign g5628 = (((g827) & (!g5033) & (g5567)) + ((g827) & (g5033) & (!g5567)));
	assign g5629 = (((g827) & (!g4892) & (!g4959) & (!g4999) & (g5057) & (!g5621)) + ((g827) & (!g4892) & (!g4959) & (!g4999) & (g5057) & (g5621)) + ((g827) & (!g4892) & (!g4959) & (g4999) & (g5057) & (!g5621)) + ((g827) & (!g4892) & (!g4959) & (g4999) & (g5057) & (g5621)) + ((g827) & (!g4892) & (g4959) & (!g4999) & (g5057) & (!g5621)) + ((g827) & (!g4892) & (g4959) & (!g4999) & (g5057) & (g5621)) + ((g827) & (!g4892) & (g4959) & (g4999) & (g5057) & (!g5621)) + ((g827) & (!g4892) & (g4959) & (g4999) & (g5057) & (g5621)) + ((g827) & (g4892) & (!g4959) & (!g4999) & (g5057) & (!g5621)) + ((g827) & (g4892) & (!g4959) & (!g4999) & (g5057) & (g5621)) + ((g827) & (g4892) & (!g4959) & (g4999) & (g5057) & (!g5621)) + ((g827) & (g4892) & (!g4959) & (g4999) & (g5057) & (g5621)) + ((g827) & (g4892) & (g4959) & (!g4999) & (g5057) & (!g5621)) + ((g827) & (g4892) & (g4959) & (!g4999) & (g5057) & (g5621)) + ((g827) & (g4892) & (g4959) & (g4999) & (!g5057) & (g5621)) + ((g827) & (g4892) & (g4959) & (g4999) & (g5057) & (!g5621)));
	assign g5630 = (((g4850) & (g4892) & (g4959) & (g4999) & (g5057) & (g5618)));
	assign g5631 = (((g827) & (!g5083) & (g5630)) + ((g827) & (g5083) & (!g5630)));
	assign g5632 = (((g827) & (!g5083) & (g5132) & (!g5630)) + ((g827) & (!g5083) & (g5132) & (g5630)) + ((g827) & (g5083) & (!g5132) & (g5630)) + ((g827) & (g5083) & (g5132) & (!g5630)));
	assign g5633 = (((g5083) & (g5132) & (g5630)));
	assign g5634 = (((g827) & (!g5165) & (g5633)) + ((g827) & (g5165) & (!g5633)));
	assign g5635 = (((g827) & (!g5165) & (g5210) & (!g5633)) + ((g827) & (!g5165) & (g5210) & (g5633)) + ((g827) & (g5165) & (!g5210) & (g5633)) + ((g827) & (g5165) & (g5210) & (!g5633)));
	assign g5636 = (((g827) & (!g5165) & (!g5210) & (g5241) & (!g5633)) + ((g827) & (!g5165) & (!g5210) & (g5241) & (g5633)) + ((g827) & (!g5165) & (g5210) & (g5241) & (!g5633)) + ((g827) & (!g5165) & (g5210) & (g5241) & (g5633)) + ((g827) & (g5165) & (!g5210) & (g5241) & (!g5633)) + ((g827) & (g5165) & (!g5210) & (g5241) & (g5633)) + ((g827) & (g5165) & (g5210) & (!g5241) & (g5633)) + ((g827) & (g5165) & (g5210) & (g5241) & (!g5633)));
	assign g5637 = (((g5083) & (g5132) & (g5165) & (g5210) & (g5241) & (g5630)));
	assign g5638 = (((g827) & (!g5294) & (g5637)) + ((g827) & (g5294) & (!g5637)));
	assign g5639 = (((g827) & (!g5294) & (g5323) & (!g5637)) + ((g827) & (!g5294) & (g5323) & (g5637)) + ((g827) & (g5294) & (!g5323) & (g5637)) + ((g827) & (g5294) & (g5323) & (!g5637)));
	assign g5640 = (((g827) & (!g5294) & (!g5323) & (g5373) & (!g5637)) + ((g827) & (!g5294) & (!g5323) & (g5373) & (g5637)) + ((g827) & (!g5294) & (g5323) & (g5373) & (!g5637)) + ((g827) & (!g5294) & (g5323) & (g5373) & (g5637)) + ((g827) & (g5294) & (!g5323) & (g5373) & (!g5637)) + ((g827) & (g5294) & (!g5323) & (g5373) & (g5637)) + ((g827) & (g5294) & (g5323) & (!g5373) & (g5637)) + ((g827) & (g5294) & (g5323) & (g5373) & (!g5637)));
	assign g5641 = (((g5294) & (g5323) & (g5373) & (g5637)));
	assign g5642 = (((g827) & (!g5393) & (g5294) & (g5323) & (g5373) & (g5637)) + ((g827) & (g5393) & (!g5294) & (!g5323) & (!g5373) & (!g5637)) + ((g827) & (g5393) & (!g5294) & (!g5323) & (!g5373) & (g5637)) + ((g827) & (g5393) & (!g5294) & (!g5323) & (g5373) & (!g5637)) + ((g827) & (g5393) & (!g5294) & (!g5323) & (g5373) & (g5637)) + ((g827) & (g5393) & (!g5294) & (g5323) & (!g5373) & (!g5637)) + ((g827) & (g5393) & (!g5294) & (g5323) & (!g5373) & (g5637)) + ((g827) & (g5393) & (!g5294) & (g5323) & (g5373) & (!g5637)) + ((g827) & (g5393) & (!g5294) & (g5323) & (g5373) & (g5637)) + ((g827) & (g5393) & (g5294) & (!g5323) & (!g5373) & (!g5637)) + ((g827) & (g5393) & (g5294) & (!g5323) & (!g5373) & (g5637)) + ((g827) & (g5393) & (g5294) & (!g5323) & (g5373) & (!g5637)) + ((g827) & (g5393) & (g5294) & (!g5323) & (g5373) & (g5637)) + ((g827) & (g5393) & (g5294) & (g5323) & (!g5373) & (!g5637)) + ((g827) & (g5393) & (g5294) & (g5323) & (!g5373) & (g5637)) + ((g827) & (g5393) & (g5294) & (g5323) & (g5373) & (!g5637)));
	assign g5643 = (((g827) & (!g5393) & (g5434) & (!g5641)) + ((g827) & (!g5393) & (g5434) & (g5641)) + ((g827) & (g5393) & (!g5434) & (g5641)) + ((g827) & (g5393) & (g5434) & (!g5641)));
	assign g5644 = (((g5294) & (g5323) & (g5373) & (g5393) & (g5434) & (g5637)));
	assign g5645 = (((g827) & (!g5463) & (g5644)) + ((g827) & (g5463) & (!g5644)));
	assign g5646 = (((g827) & (!g5463) & (g5510) & (!g5644)) + ((g827) & (!g5463) & (g5510) & (g5644)) + ((g827) & (g5463) & (!g5510) & (g5644)) + ((g827) & (g5463) & (g5510) & (!g5644)));
	assign g5647 = (((g827) & (!g5463) & (!g5510) & (g5533) & (!g5644)) + ((g827) & (!g5463) & (!g5510) & (g5533) & (g5644)) + ((g827) & (!g5463) & (g5510) & (g5533) & (!g5644)) + ((g827) & (!g5463) & (g5510) & (g5533) & (g5644)) + ((g827) & (g5463) & (!g5510) & (g5533) & (!g5644)) + ((g827) & (g5463) & (!g5510) & (g5533) & (g5644)) + ((g827) & (g5463) & (g5510) & (!g5533) & (g5644)) + ((g827) & (g5463) & (g5510) & (g5533) & (!g5644)));
	assign g5648 = (((!g827) & (!g731) & (g1814)) + ((!g827) & (g731) & (g1814)) + ((g827) & (!g731) & (!g1814)) + ((g827) & (g731) & (g1814)));
	assign g5649 = (((!g827) & (!g1784) & (g2678)) + ((!g827) & (g1784) & (g2678)) + ((g827) & (!g1784) & (!g2678)) + ((g827) & (g1784) & (g2678)));
	assign g5650 = (((!g827) & (!g1786) & (g3291)) + ((!g827) & (g1786) & (g3291)) + ((g827) & (!g1786) & (!g3291)) + ((g827) & (g1786) & (g3291)));
	assign g5651 = (((!g827) & (!g1788) & (g2679)) + ((!g827) & (g1788) & (g2679)) + ((g827) & (!g1788) & (!g2679)) + ((g827) & (g1788) & (g2679)));
	assign g5652 = (((!g827) & (!g1790) & (g2683)) + ((!g827) & (g1790) & (g2683)) + ((g827) & (!g1790) & (!g2683)) + ((g827) & (g1790) & (g2683)));
	assign g5653 = (((!g827) & (!g1792) & (g3295)) + ((!g827) & (g1792) & (g3295)) + ((g827) & (!g1792) & (!g3295)) + ((g827) & (g1792) & (g3295)));
	assign g5654 = (((!g827) & (!g1794) & (g3297)) + ((!g827) & (g1794) & (g3297)) + ((g827) & (!g1794) & (!g3297)) + ((g827) & (g1794) & (g3297)));
	assign g5655 = (((!g827) & (!g1796) & (g3299)) + ((!g827) & (g1796) & (g3299)) + ((g827) & (!g1796) & (!g3299)) + ((g827) & (g1796) & (g3299)));
	assign g5656 = (((!g827) & (!g1798) & (g3301)) + ((!g827) & (g1798) & (g3301)) + ((g827) & (!g1798) & (!g3301)) + ((g827) & (g1798) & (g3301)));
	assign g5657 = (((!g827) & (!g1800) & (g3303)) + ((!g827) & (g1800) & (g3303)) + ((g827) & (!g1800) & (!g3303)) + ((g827) & (g1800) & (g3303)));
	assign g5658 = (((!g827) & (!g1802) & (g3305)) + ((!g827) & (g1802) & (g3305)) + ((g827) & (!g1802) & (!g3305)) + ((g827) & (g1802) & (g3305)));
	assign g5659 = (((!g827) & (!g1804) & (g3307)) + ((!g827) & (g1804) & (g3307)) + ((g827) & (!g1804) & (!g3307)) + ((g827) & (g1804) & (g3307)));
	assign g5660 = (((!g827) & (!g1806) & (g2684)) + ((!g827) & (g1806) & (g2684)) + ((g827) & (!g1806) & (!g2684)) + ((g827) & (g1806) & (g2684)));
	assign g5661 = (((!g827) & (!g1808) & (g3310)) + ((!g827) & (g1808) & (g3310)) + ((g827) & (!g1808) & (!g3310)) + ((g827) & (g1808) & (g3310)));
	assign g5662 = (((!g827) & (!g1810) & (g3312)) + ((!g827) & (g1810) & (g3312)) + ((g827) & (!g1810) & (!g3312)) + ((g827) & (g1810) & (g3312)));
	assign g5663 = (((!g827) & (!g1812) & (g3314)) + ((!g827) & (g1812) & (g3314)) + ((g827) & (!g1812) & (!g3314)) + ((g827) & (g1812) & (g3314)));
	assign g5664 = (((!g2184) & (!g1914) & (!g2759) & (!g1847) & (!g3086) & (!g3090)) + ((!g2184) & (!g1914) & (!g2759) & (!g1847) & (g3086) & (g3090)) + ((!g2184) & (!g1914) & (!g2759) & (g1847) & (!g3086) & (!g3090)) + ((!g2184) & (!g1914) & (!g2759) & (g1847) & (g3086) & (g3090)) + ((!g2184) & (!g1914) & (g2759) & (!g1847) & (!g3086) & (!g3090)) + ((!g2184) & (!g1914) & (g2759) & (!g1847) & (g3086) & (g3090)) + ((!g2184) & (!g1914) & (g2759) & (g1847) & (!g3086) & (!g3090)) + ((!g2184) & (!g1914) & (g2759) & (g1847) & (g3086) & (g3090)) + ((!g2184) & (g1914) & (!g2759) & (!g1847) & (!g3086) & (!g3090)) + ((!g2184) & (g1914) & (!g2759) & (!g1847) & (!g3086) & (g3090)) + ((!g2184) & (g1914) & (!g2759) & (!g1847) & (g3086) & (!g3090)) + ((!g2184) & (g1914) & (!g2759) & (!g1847) & (g3086) & (g3090)) + ((!g2184) & (g1914) & (g2759) & (g1847) & (!g3086) & (!g3090)) + ((!g2184) & (g1914) & (g2759) & (g1847) & (!g3086) & (g3090)) + ((!g2184) & (g1914) & (g2759) & (g1847) & (g3086) & (!g3090)) + ((!g2184) & (g1914) & (g2759) & (g1847) & (g3086) & (g3090)) + ((g2184) & (!g1914) & (!g2759) & (!g1847) & (!g3086) & (g3090)) + ((g2184) & (!g1914) & (!g2759) & (!g1847) & (g3086) & (!g3090)) + ((g2184) & (!g1914) & (!g2759) & (g1847) & (!g3086) & (g3090)) + ((g2184) & (!g1914) & (!g2759) & (g1847) & (g3086) & (!g3090)) + ((g2184) & (!g1914) & (g2759) & (!g1847) & (!g3086) & (g3090)) + ((g2184) & (!g1914) & (g2759) & (!g1847) & (g3086) & (!g3090)) + ((g2184) & (!g1914) & (g2759) & (g1847) & (!g3086) & (g3090)) + ((g2184) & (!g1914) & (g2759) & (g1847) & (g3086) & (!g3090)) + ((g2184) & (g1914) & (!g2759) & (g1847) & (!g3086) & (!g3090)) + ((g2184) & (g1914) & (!g2759) & (g1847) & (!g3086) & (g3090)) + ((g2184) & (g1914) & (!g2759) & (g1847) & (g3086) & (!g3090)) + ((g2184) & (g1914) & (!g2759) & (g1847) & (g3086) & (g3090)) + ((g2184) & (g1914) & (g2759) & (!g1847) & (!g3086) & (!g3090)) + ((g2184) & (g1914) & (g2759) & (!g1847) & (!g3086) & (g3090)) + ((g2184) & (g1914) & (g2759) & (!g1847) & (g3086) & (!g3090)) + ((g2184) & (g1914) & (g2759) & (!g1847) & (g3086) & (g3090)));
	assign g5665 = (((!g1949) & (!g1914) & (!g3353) & (!g3359) & (!g2423) & (!g3084)) + ((!g1949) & (!g1914) & (!g3353) & (!g3359) & (!g2423) & (g3084)) + ((!g1949) & (!g1914) & (!g3353) & (!g3359) & (g2423) & (!g3084)) + ((!g1949) & (!g1914) & (!g3353) & (!g3359) & (g2423) & (g3084)) + ((!g1949) & (!g1914) & (g3353) & (g3359) & (!g2423) & (!g3084)) + ((!g1949) & (!g1914) & (g3353) & (g3359) & (!g2423) & (g3084)) + ((!g1949) & (!g1914) & (g3353) & (g3359) & (g2423) & (!g3084)) + ((!g1949) & (!g1914) & (g3353) & (g3359) & (g2423) & (g3084)) + ((!g1949) & (g1914) & (!g3353) & (!g3359) & (!g2423) & (!g3084)) + ((!g1949) & (g1914) & (!g3353) & (!g3359) & (g2423) & (g3084)) + ((!g1949) & (g1914) & (!g3353) & (g3359) & (!g2423) & (!g3084)) + ((!g1949) & (g1914) & (!g3353) & (g3359) & (g2423) & (g3084)) + ((!g1949) & (g1914) & (g3353) & (!g3359) & (!g2423) & (!g3084)) + ((!g1949) & (g1914) & (g3353) & (!g3359) & (g2423) & (g3084)) + ((!g1949) & (g1914) & (g3353) & (g3359) & (!g2423) & (!g3084)) + ((!g1949) & (g1914) & (g3353) & (g3359) & (g2423) & (g3084)) + ((g1949) & (!g1914) & (!g3353) & (g3359) & (!g2423) & (!g3084)) + ((g1949) & (!g1914) & (!g3353) & (g3359) & (!g2423) & (g3084)) + ((g1949) & (!g1914) & (!g3353) & (g3359) & (g2423) & (!g3084)) + ((g1949) & (!g1914) & (!g3353) & (g3359) & (g2423) & (g3084)) + ((g1949) & (!g1914) & (g3353) & (!g3359) & (!g2423) & (!g3084)) + ((g1949) & (!g1914) & (g3353) & (!g3359) & (!g2423) & (g3084)) + ((g1949) & (!g1914) & (g3353) & (!g3359) & (g2423) & (!g3084)) + ((g1949) & (!g1914) & (g3353) & (!g3359) & (g2423) & (g3084)) + ((g1949) & (g1914) & (!g3353) & (!g3359) & (!g2423) & (g3084)) + ((g1949) & (g1914) & (!g3353) & (!g3359) & (g2423) & (!g3084)) + ((g1949) & (g1914) & (!g3353) & (g3359) & (!g2423) & (g3084)) + ((g1949) & (g1914) & (!g3353) & (g3359) & (g2423) & (!g3084)) + ((g1949) & (g1914) & (g3353) & (!g3359) & (!g2423) & (g3084)) + ((g1949) & (g1914) & (g3353) & (!g3359) & (g2423) & (!g3084)) + ((g1949) & (g1914) & (g3353) & (g3359) & (!g2423) & (g3084)) + ((g1949) & (g1914) & (g3353) & (g3359) & (g2423) & (!g3084)));
	assign g5666 = (((!g2190) & (!g1914) & (!g3339) & (!g3345) & (!g2426) & (!g3093)) + ((!g2190) & (!g1914) & (!g3339) & (!g3345) & (!g2426) & (g3093)) + ((!g2190) & (!g1914) & (!g3339) & (!g3345) & (g2426) & (!g3093)) + ((!g2190) & (!g1914) & (!g3339) & (!g3345) & (g2426) & (g3093)) + ((!g2190) & (!g1914) & (g3339) & (g3345) & (!g2426) & (!g3093)) + ((!g2190) & (!g1914) & (g3339) & (g3345) & (!g2426) & (g3093)) + ((!g2190) & (!g1914) & (g3339) & (g3345) & (g2426) & (!g3093)) + ((!g2190) & (!g1914) & (g3339) & (g3345) & (g2426) & (g3093)) + ((!g2190) & (g1914) & (!g3339) & (!g3345) & (!g2426) & (!g3093)) + ((!g2190) & (g1914) & (!g3339) & (!g3345) & (g2426) & (g3093)) + ((!g2190) & (g1914) & (!g3339) & (g3345) & (!g2426) & (!g3093)) + ((!g2190) & (g1914) & (!g3339) & (g3345) & (g2426) & (g3093)) + ((!g2190) & (g1914) & (g3339) & (!g3345) & (!g2426) & (!g3093)) + ((!g2190) & (g1914) & (g3339) & (!g3345) & (g2426) & (g3093)) + ((!g2190) & (g1914) & (g3339) & (g3345) & (!g2426) & (!g3093)) + ((!g2190) & (g1914) & (g3339) & (g3345) & (g2426) & (g3093)) + ((g2190) & (!g1914) & (!g3339) & (g3345) & (!g2426) & (!g3093)) + ((g2190) & (!g1914) & (!g3339) & (g3345) & (!g2426) & (g3093)) + ((g2190) & (!g1914) & (!g3339) & (g3345) & (g2426) & (!g3093)) + ((g2190) & (!g1914) & (!g3339) & (g3345) & (g2426) & (g3093)) + ((g2190) & (!g1914) & (g3339) & (!g3345) & (!g2426) & (!g3093)) + ((g2190) & (!g1914) & (g3339) & (!g3345) & (!g2426) & (g3093)) + ((g2190) & (!g1914) & (g3339) & (!g3345) & (g2426) & (!g3093)) + ((g2190) & (!g1914) & (g3339) & (!g3345) & (g2426) & (g3093)) + ((g2190) & (g1914) & (!g3339) & (!g3345) & (!g2426) & (g3093)) + ((g2190) & (g1914) & (!g3339) & (!g3345) & (g2426) & (!g3093)) + ((g2190) & (g1914) & (!g3339) & (g3345) & (!g2426) & (g3093)) + ((g2190) & (g1914) & (!g3339) & (g3345) & (g2426) & (!g3093)) + ((g2190) & (g1914) & (g3339) & (!g3345) & (!g2426) & (g3093)) + ((g2190) & (g1914) & (g3339) & (!g3345) & (g2426) & (!g3093)) + ((g2190) & (g1914) & (g3339) & (g3345) & (!g2426) & (g3093)) + ((g2190) & (g1914) & (g3339) & (g3345) & (g2426) & (!g3093)));
	assign g5667 = (((!g2192) & (!g1914) & (!g3330) & (!g3342) & (!g2424) & (!g3095)) + ((!g2192) & (!g1914) & (!g3330) & (!g3342) & (g2424) & (g3095)) + ((!g2192) & (!g1914) & (!g3330) & (g3342) & (!g2424) & (!g3095)) + ((!g2192) & (!g1914) & (!g3330) & (g3342) & (g2424) & (g3095)) + ((!g2192) & (!g1914) & (g3330) & (!g3342) & (!g2424) & (!g3095)) + ((!g2192) & (!g1914) & (g3330) & (!g3342) & (g2424) & (g3095)) + ((!g2192) & (!g1914) & (g3330) & (g3342) & (!g2424) & (!g3095)) + ((!g2192) & (!g1914) & (g3330) & (g3342) & (g2424) & (g3095)) + ((!g2192) & (g1914) & (!g3330) & (!g3342) & (!g2424) & (!g3095)) + ((!g2192) & (g1914) & (!g3330) & (!g3342) & (!g2424) & (g3095)) + ((!g2192) & (g1914) & (!g3330) & (!g3342) & (g2424) & (!g3095)) + ((!g2192) & (g1914) & (!g3330) & (!g3342) & (g2424) & (g3095)) + ((!g2192) & (g1914) & (g3330) & (g3342) & (!g2424) & (!g3095)) + ((!g2192) & (g1914) & (g3330) & (g3342) & (!g2424) & (g3095)) + ((!g2192) & (g1914) & (g3330) & (g3342) & (g2424) & (!g3095)) + ((!g2192) & (g1914) & (g3330) & (g3342) & (g2424) & (g3095)) + ((g2192) & (!g1914) & (!g3330) & (!g3342) & (!g2424) & (g3095)) + ((g2192) & (!g1914) & (!g3330) & (!g3342) & (g2424) & (!g3095)) + ((g2192) & (!g1914) & (!g3330) & (g3342) & (!g2424) & (g3095)) + ((g2192) & (!g1914) & (!g3330) & (g3342) & (g2424) & (!g3095)) + ((g2192) & (!g1914) & (g3330) & (!g3342) & (!g2424) & (g3095)) + ((g2192) & (!g1914) & (g3330) & (!g3342) & (g2424) & (!g3095)) + ((g2192) & (!g1914) & (g3330) & (g3342) & (!g2424) & (g3095)) + ((g2192) & (!g1914) & (g3330) & (g3342) & (g2424) & (!g3095)) + ((g2192) & (g1914) & (!g3330) & (g3342) & (!g2424) & (!g3095)) + ((g2192) & (g1914) & (!g3330) & (g3342) & (!g2424) & (g3095)) + ((g2192) & (g1914) & (!g3330) & (g3342) & (g2424) & (!g3095)) + ((g2192) & (g1914) & (!g3330) & (g3342) & (g2424) & (g3095)) + ((g2192) & (g1914) & (g3330) & (!g3342) & (!g2424) & (!g3095)) + ((g2192) & (g1914) & (g3330) & (!g3342) & (!g2424) & (g3095)) + ((g2192) & (g1914) & (g3330) & (!g3342) & (g2424) & (!g3095)) + ((g2192) & (g1914) & (g3330) & (!g3342) & (g2424) & (g3095)));
	assign g5668 = (((!g2194) & (!g1914) & (!g2761) & (!g1847) & (!g3080) & (!g3095)) + ((!g2194) & (!g1914) & (!g2761) & (!g1847) & (!g3080) & (g3095)) + ((!g2194) & (!g1914) & (!g2761) & (!g1847) & (g3080) & (!g3095)) + ((!g2194) & (!g1914) & (!g2761) & (!g1847) & (g3080) & (g3095)) + ((!g2194) & (!g1914) & (g2761) & (g1847) & (!g3080) & (!g3095)) + ((!g2194) & (!g1914) & (g2761) & (g1847) & (!g3080) & (g3095)) + ((!g2194) & (!g1914) & (g2761) & (g1847) & (g3080) & (!g3095)) + ((!g2194) & (!g1914) & (g2761) & (g1847) & (g3080) & (g3095)) + ((!g2194) & (g1914) & (!g2761) & (!g1847) & (!g3080) & (!g3095)) + ((!g2194) & (g1914) & (!g2761) & (!g1847) & (g3080) & (g3095)) + ((!g2194) & (g1914) & (!g2761) & (g1847) & (!g3080) & (!g3095)) + ((!g2194) & (g1914) & (!g2761) & (g1847) & (g3080) & (g3095)) + ((!g2194) & (g1914) & (g2761) & (!g1847) & (!g3080) & (!g3095)) + ((!g2194) & (g1914) & (g2761) & (!g1847) & (g3080) & (g3095)) + ((!g2194) & (g1914) & (g2761) & (g1847) & (!g3080) & (!g3095)) + ((!g2194) & (g1914) & (g2761) & (g1847) & (g3080) & (g3095)) + ((g2194) & (!g1914) & (!g2761) & (g1847) & (!g3080) & (!g3095)) + ((g2194) & (!g1914) & (!g2761) & (g1847) & (!g3080) & (g3095)) + ((g2194) & (!g1914) & (!g2761) & (g1847) & (g3080) & (!g3095)) + ((g2194) & (!g1914) & (!g2761) & (g1847) & (g3080) & (g3095)) + ((g2194) & (!g1914) & (g2761) & (!g1847) & (!g3080) & (!g3095)) + ((g2194) & (!g1914) & (g2761) & (!g1847) & (!g3080) & (g3095)) + ((g2194) & (!g1914) & (g2761) & (!g1847) & (g3080) & (!g3095)) + ((g2194) & (!g1914) & (g2761) & (!g1847) & (g3080) & (g3095)) + ((g2194) & (g1914) & (!g2761) & (!g1847) & (!g3080) & (g3095)) + ((g2194) & (g1914) & (!g2761) & (!g1847) & (g3080) & (!g3095)) + ((g2194) & (g1914) & (!g2761) & (g1847) & (!g3080) & (g3095)) + ((g2194) & (g1914) & (!g2761) & (g1847) & (g3080) & (!g3095)) + ((g2194) & (g1914) & (g2761) & (!g1847) & (!g3080) & (g3095)) + ((g2194) & (g1914) & (g2761) & (!g1847) & (g3080) & (!g3095)) + ((g2194) & (g1914) & (g2761) & (g1847) & (!g3080) & (g3095)) + ((g2194) & (g1914) & (g2761) & (g1847) & (g3080) & (!g3095)));
	assign g5669 = (((!g2196) & (!g1914) & (!g3345) & (!g3323) & (!g2423) & (!g3082)) + ((!g2196) & (!g1914) & (!g3345) & (!g3323) & (g2423) & (g3082)) + ((!g2196) & (!g1914) & (!g3345) & (g3323) & (!g2423) & (!g3082)) + ((!g2196) & (!g1914) & (!g3345) & (g3323) & (g2423) & (g3082)) + ((!g2196) & (!g1914) & (g3345) & (!g3323) & (!g2423) & (!g3082)) + ((!g2196) & (!g1914) & (g3345) & (!g3323) & (g2423) & (g3082)) + ((!g2196) & (!g1914) & (g3345) & (g3323) & (!g2423) & (!g3082)) + ((!g2196) & (!g1914) & (g3345) & (g3323) & (g2423) & (g3082)) + ((!g2196) & (g1914) & (!g3345) & (!g3323) & (!g2423) & (!g3082)) + ((!g2196) & (g1914) & (!g3345) & (!g3323) & (!g2423) & (g3082)) + ((!g2196) & (g1914) & (!g3345) & (!g3323) & (g2423) & (!g3082)) + ((!g2196) & (g1914) & (!g3345) & (!g3323) & (g2423) & (g3082)) + ((!g2196) & (g1914) & (g3345) & (g3323) & (!g2423) & (!g3082)) + ((!g2196) & (g1914) & (g3345) & (g3323) & (!g2423) & (g3082)) + ((!g2196) & (g1914) & (g3345) & (g3323) & (g2423) & (!g3082)) + ((!g2196) & (g1914) & (g3345) & (g3323) & (g2423) & (g3082)) + ((g2196) & (!g1914) & (!g3345) & (!g3323) & (!g2423) & (g3082)) + ((g2196) & (!g1914) & (!g3345) & (!g3323) & (g2423) & (!g3082)) + ((g2196) & (!g1914) & (!g3345) & (g3323) & (!g2423) & (g3082)) + ((g2196) & (!g1914) & (!g3345) & (g3323) & (g2423) & (!g3082)) + ((g2196) & (!g1914) & (g3345) & (!g3323) & (!g2423) & (g3082)) + ((g2196) & (!g1914) & (g3345) & (!g3323) & (g2423) & (!g3082)) + ((g2196) & (!g1914) & (g3345) & (g3323) & (!g2423) & (g3082)) + ((g2196) & (!g1914) & (g3345) & (g3323) & (g2423) & (!g3082)) + ((g2196) & (g1914) & (!g3345) & (g3323) & (!g2423) & (!g3082)) + ((g2196) & (g1914) & (!g3345) & (g3323) & (!g2423) & (g3082)) + ((g2196) & (g1914) & (!g3345) & (g3323) & (g2423) & (!g3082)) + ((g2196) & (g1914) & (!g3345) & (g3323) & (g2423) & (g3082)) + ((g2196) & (g1914) & (g3345) & (!g3323) & (!g2423) & (!g3082)) + ((g2196) & (g1914) & (g3345) & (!g3323) & (!g2423) & (g3082)) + ((g2196) & (g1914) & (g3345) & (!g3323) & (g2423) & (!g3082)) + ((g2196) & (g1914) & (g3345) & (!g3323) & (g2423) & (g3082)));
	assign g5670 = (((!g1987) & (!g1914) & (!g3359) & (!g3336) & (!g2426) & (!g3074)) + ((!g1987) & (!g1914) & (!g3359) & (!g3336) & (g2426) & (g3074)) + ((!g1987) & (!g1914) & (!g3359) & (g3336) & (!g2426) & (!g3074)) + ((!g1987) & (!g1914) & (!g3359) & (g3336) & (g2426) & (g3074)) + ((!g1987) & (!g1914) & (g3359) & (!g3336) & (!g2426) & (!g3074)) + ((!g1987) & (!g1914) & (g3359) & (!g3336) & (g2426) & (g3074)) + ((!g1987) & (!g1914) & (g3359) & (g3336) & (!g2426) & (!g3074)) + ((!g1987) & (!g1914) & (g3359) & (g3336) & (g2426) & (g3074)) + ((!g1987) & (g1914) & (!g3359) & (!g3336) & (!g2426) & (!g3074)) + ((!g1987) & (g1914) & (!g3359) & (!g3336) & (!g2426) & (g3074)) + ((!g1987) & (g1914) & (!g3359) & (!g3336) & (g2426) & (!g3074)) + ((!g1987) & (g1914) & (!g3359) & (!g3336) & (g2426) & (g3074)) + ((!g1987) & (g1914) & (g3359) & (g3336) & (!g2426) & (!g3074)) + ((!g1987) & (g1914) & (g3359) & (g3336) & (!g2426) & (g3074)) + ((!g1987) & (g1914) & (g3359) & (g3336) & (g2426) & (!g3074)) + ((!g1987) & (g1914) & (g3359) & (g3336) & (g2426) & (g3074)) + ((g1987) & (!g1914) & (!g3359) & (!g3336) & (!g2426) & (g3074)) + ((g1987) & (!g1914) & (!g3359) & (!g3336) & (g2426) & (!g3074)) + ((g1987) & (!g1914) & (!g3359) & (g3336) & (!g2426) & (g3074)) + ((g1987) & (!g1914) & (!g3359) & (g3336) & (g2426) & (!g3074)) + ((g1987) & (!g1914) & (g3359) & (!g3336) & (!g2426) & (g3074)) + ((g1987) & (!g1914) & (g3359) & (!g3336) & (g2426) & (!g3074)) + ((g1987) & (!g1914) & (g3359) & (g3336) & (!g2426) & (g3074)) + ((g1987) & (!g1914) & (g3359) & (g3336) & (g2426) & (!g3074)) + ((g1987) & (g1914) & (!g3359) & (g3336) & (!g2426) & (!g3074)) + ((g1987) & (g1914) & (!g3359) & (g3336) & (!g2426) & (g3074)) + ((g1987) & (g1914) & (!g3359) & (g3336) & (g2426) & (!g3074)) + ((g1987) & (g1914) & (!g3359) & (g3336) & (g2426) & (g3074)) + ((g1987) & (g1914) & (g3359) & (!g3336) & (!g2426) & (!g3074)) + ((g1987) & (g1914) & (g3359) & (!g3336) & (!g2426) & (g3074)) + ((g1987) & (g1914) & (g3359) & (!g3336) & (g2426) & (!g3074)) + ((g1987) & (g1914) & (g3359) & (!g3336) & (g2426) & (g3074)));
	assign g5671 = (((!g2203) & (!g1914) & (!g3330) & (!g3333) & (!g2427) & (!g3090)) + ((!g2203) & (!g1914) & (!g3330) & (!g3333) & (!g2427) & (g3090)) + ((!g2203) & (!g1914) & (!g3330) & (!g3333) & (g2427) & (!g3090)) + ((!g2203) & (!g1914) & (!g3330) & (!g3333) & (g2427) & (g3090)) + ((!g2203) & (!g1914) & (g3330) & (g3333) & (!g2427) & (!g3090)) + ((!g2203) & (!g1914) & (g3330) & (g3333) & (!g2427) & (g3090)) + ((!g2203) & (!g1914) & (g3330) & (g3333) & (g2427) & (!g3090)) + ((!g2203) & (!g1914) & (g3330) & (g3333) & (g2427) & (g3090)) + ((!g2203) & (g1914) & (!g3330) & (!g3333) & (!g2427) & (!g3090)) + ((!g2203) & (g1914) & (!g3330) & (!g3333) & (g2427) & (g3090)) + ((!g2203) & (g1914) & (!g3330) & (g3333) & (!g2427) & (!g3090)) + ((!g2203) & (g1914) & (!g3330) & (g3333) & (g2427) & (g3090)) + ((!g2203) & (g1914) & (g3330) & (!g3333) & (!g2427) & (!g3090)) + ((!g2203) & (g1914) & (g3330) & (!g3333) & (g2427) & (g3090)) + ((!g2203) & (g1914) & (g3330) & (g3333) & (!g2427) & (!g3090)) + ((!g2203) & (g1914) & (g3330) & (g3333) & (g2427) & (g3090)) + ((g2203) & (!g1914) & (!g3330) & (g3333) & (!g2427) & (!g3090)) + ((g2203) & (!g1914) & (!g3330) & (g3333) & (!g2427) & (g3090)) + ((g2203) & (!g1914) & (!g3330) & (g3333) & (g2427) & (!g3090)) + ((g2203) & (!g1914) & (!g3330) & (g3333) & (g2427) & (g3090)) + ((g2203) & (!g1914) & (g3330) & (!g3333) & (!g2427) & (!g3090)) + ((g2203) & (!g1914) & (g3330) & (!g3333) & (!g2427) & (g3090)) + ((g2203) & (!g1914) & (g3330) & (!g3333) & (g2427) & (!g3090)) + ((g2203) & (!g1914) & (g3330) & (!g3333) & (g2427) & (g3090)) + ((g2203) & (g1914) & (!g3330) & (!g3333) & (!g2427) & (g3090)) + ((g2203) & (g1914) & (!g3330) & (!g3333) & (g2427) & (!g3090)) + ((g2203) & (g1914) & (!g3330) & (g3333) & (!g2427) & (g3090)) + ((g2203) & (g1914) & (!g3330) & (g3333) & (g2427) & (!g3090)) + ((g2203) & (g1914) & (g3330) & (!g3333) & (!g2427) & (g3090)) + ((g2203) & (g1914) & (g3330) & (!g3333) & (g2427) & (!g3090)) + ((g2203) & (g1914) & (g3330) & (g3333) & (!g2427) & (g3090)) + ((g2203) & (g1914) & (g3330) & (g3333) & (g2427) & (!g3090)));
	assign g5672 = (((!g1955) & (!g1914) & (!g1847) & (!g3339) & (!g3330) & (!g3336)) + ((!g1955) & (!g1914) & (!g1847) & (!g3339) & (g3330) & (g3336)) + ((!g1955) & (!g1914) & (!g1847) & (g3339) & (!g3330) & (!g3336)) + ((!g1955) & (!g1914) & (!g1847) & (g3339) & (g3330) & (g3336)) + ((!g1955) & (!g1914) & (g1847) & (!g3339) & (!g3330) & (!g3336)) + ((!g1955) & (!g1914) & (g1847) & (!g3339) & (g3330) & (g3336)) + ((!g1955) & (!g1914) & (g1847) & (g3339) & (!g3330) & (!g3336)) + ((!g1955) & (!g1914) & (g1847) & (g3339) & (g3330) & (g3336)) + ((!g1955) & (g1914) & (!g1847) & (!g3339) & (!g3330) & (!g3336)) + ((!g1955) & (g1914) & (!g1847) & (!g3339) & (!g3330) & (g3336)) + ((!g1955) & (g1914) & (!g1847) & (!g3339) & (g3330) & (!g3336)) + ((!g1955) & (g1914) & (!g1847) & (!g3339) & (g3330) & (g3336)) + ((!g1955) & (g1914) & (g1847) & (g3339) & (!g3330) & (!g3336)) + ((!g1955) & (g1914) & (g1847) & (g3339) & (!g3330) & (g3336)) + ((!g1955) & (g1914) & (g1847) & (g3339) & (g3330) & (!g3336)) + ((!g1955) & (g1914) & (g1847) & (g3339) & (g3330) & (g3336)) + ((g1955) & (!g1914) & (!g1847) & (!g3339) & (!g3330) & (g3336)) + ((g1955) & (!g1914) & (!g1847) & (!g3339) & (g3330) & (!g3336)) + ((g1955) & (!g1914) & (!g1847) & (g3339) & (!g3330) & (g3336)) + ((g1955) & (!g1914) & (!g1847) & (g3339) & (g3330) & (!g3336)) + ((g1955) & (!g1914) & (g1847) & (!g3339) & (!g3330) & (g3336)) + ((g1955) & (!g1914) & (g1847) & (!g3339) & (g3330) & (!g3336)) + ((g1955) & (!g1914) & (g1847) & (g3339) & (!g3330) & (g3336)) + ((g1955) & (!g1914) & (g1847) & (g3339) & (g3330) & (!g3336)) + ((g1955) & (g1914) & (!g1847) & (g3339) & (!g3330) & (!g3336)) + ((g1955) & (g1914) & (!g1847) & (g3339) & (!g3330) & (g3336)) + ((g1955) & (g1914) & (!g1847) & (g3339) & (g3330) & (!g3336)) + ((g1955) & (g1914) & (!g1847) & (g3339) & (g3330) & (g3336)) + ((g1955) & (g1914) & (g1847) & (!g3339) & (!g3330) & (!g3336)) + ((g1955) & (g1914) & (g1847) & (!g3339) & (!g3330) & (g3336)) + ((g1955) & (g1914) & (g1847) & (!g3339) & (g3330) & (!g3336)) + ((g1955) & (g1914) & (g1847) & (!g3339) & (g3330) & (g3336)));
	assign g5673 = (((!g1993) & (!g1914) & (!g3353) & (!g3330) & (!g1847) & (!g3323)) + ((!g1993) & (!g1914) & (!g3353) & (!g3330) & (g1847) & (g3323)) + ((!g1993) & (!g1914) & (!g3353) & (g3330) & (!g1847) & (!g3323)) + ((!g1993) & (!g1914) & (!g3353) & (g3330) & (g1847) & (g3323)) + ((!g1993) & (!g1914) & (g3353) & (!g3330) & (!g1847) & (!g3323)) + ((!g1993) & (!g1914) & (g3353) & (!g3330) & (g1847) & (g3323)) + ((!g1993) & (!g1914) & (g3353) & (g3330) & (!g1847) & (!g3323)) + ((!g1993) & (!g1914) & (g3353) & (g3330) & (g1847) & (g3323)) + ((!g1993) & (g1914) & (!g3353) & (!g3330) & (!g1847) & (!g3323)) + ((!g1993) & (g1914) & (!g3353) & (!g3330) & (!g1847) & (g3323)) + ((!g1993) & (g1914) & (!g3353) & (!g3330) & (g1847) & (!g3323)) + ((!g1993) & (g1914) & (!g3353) & (!g3330) & (g1847) & (g3323)) + ((!g1993) & (g1914) & (g3353) & (g3330) & (!g1847) & (!g3323)) + ((!g1993) & (g1914) & (g3353) & (g3330) & (!g1847) & (g3323)) + ((!g1993) & (g1914) & (g3353) & (g3330) & (g1847) & (!g3323)) + ((!g1993) & (g1914) & (g3353) & (g3330) & (g1847) & (g3323)) + ((g1993) & (!g1914) & (!g3353) & (!g3330) & (!g1847) & (g3323)) + ((g1993) & (!g1914) & (!g3353) & (!g3330) & (g1847) & (!g3323)) + ((g1993) & (!g1914) & (!g3353) & (g3330) & (!g1847) & (g3323)) + ((g1993) & (!g1914) & (!g3353) & (g3330) & (g1847) & (!g3323)) + ((g1993) & (!g1914) & (g3353) & (!g3330) & (!g1847) & (g3323)) + ((g1993) & (!g1914) & (g3353) & (!g3330) & (g1847) & (!g3323)) + ((g1993) & (!g1914) & (g3353) & (g3330) & (!g1847) & (g3323)) + ((g1993) & (!g1914) & (g3353) & (g3330) & (g1847) & (!g3323)) + ((g1993) & (g1914) & (!g3353) & (g3330) & (!g1847) & (!g3323)) + ((g1993) & (g1914) & (!g3353) & (g3330) & (!g1847) & (g3323)) + ((g1993) & (g1914) & (!g3353) & (g3330) & (g1847) & (!g3323)) + ((g1993) & (g1914) & (!g3353) & (g3330) & (g1847) & (g3323)) + ((g1993) & (g1914) & (g3353) & (!g3330) & (!g1847) & (!g3323)) + ((g1993) & (g1914) & (g3353) & (!g3330) & (!g1847) & (g3323)) + ((g1993) & (g1914) & (g3353) & (!g3330) & (g1847) & (!g3323)) + ((g1993) & (g1914) & (g3353) & (!g3330) & (g1847) & (g3323)));
	assign g5674 = (((!g2283) & (!g1914) & (!g3345) & (!g3333) & (!g2759) & (!g3359)) + ((!g2283) & (!g1914) & (!g3345) & (!g3333) & (g2759) & (g3359)) + ((!g2283) & (!g1914) & (!g3345) & (g3333) & (!g2759) & (!g3359)) + ((!g2283) & (!g1914) & (!g3345) & (g3333) & (g2759) & (g3359)) + ((!g2283) & (!g1914) & (g3345) & (!g3333) & (!g2759) & (!g3359)) + ((!g2283) & (!g1914) & (g3345) & (!g3333) & (g2759) & (g3359)) + ((!g2283) & (!g1914) & (g3345) & (g3333) & (!g2759) & (!g3359)) + ((!g2283) & (!g1914) & (g3345) & (g3333) & (g2759) & (g3359)) + ((!g2283) & (g1914) & (!g3345) & (!g3333) & (!g2759) & (!g3359)) + ((!g2283) & (g1914) & (!g3345) & (!g3333) & (!g2759) & (g3359)) + ((!g2283) & (g1914) & (!g3345) & (!g3333) & (g2759) & (!g3359)) + ((!g2283) & (g1914) & (!g3345) & (!g3333) & (g2759) & (g3359)) + ((!g2283) & (g1914) & (g3345) & (g3333) & (!g2759) & (!g3359)) + ((!g2283) & (g1914) & (g3345) & (g3333) & (!g2759) & (g3359)) + ((!g2283) & (g1914) & (g3345) & (g3333) & (g2759) & (!g3359)) + ((!g2283) & (g1914) & (g3345) & (g3333) & (g2759) & (g3359)) + ((g2283) & (!g1914) & (!g3345) & (!g3333) & (!g2759) & (g3359)) + ((g2283) & (!g1914) & (!g3345) & (!g3333) & (g2759) & (!g3359)) + ((g2283) & (!g1914) & (!g3345) & (g3333) & (!g2759) & (g3359)) + ((g2283) & (!g1914) & (!g3345) & (g3333) & (g2759) & (!g3359)) + ((g2283) & (!g1914) & (g3345) & (!g3333) & (!g2759) & (g3359)) + ((g2283) & (!g1914) & (g3345) & (!g3333) & (g2759) & (!g3359)) + ((g2283) & (!g1914) & (g3345) & (g3333) & (!g2759) & (g3359)) + ((g2283) & (!g1914) & (g3345) & (g3333) & (g2759) & (!g3359)) + ((g2283) & (g1914) & (!g3345) & (g3333) & (!g2759) & (!g3359)) + ((g2283) & (g1914) & (!g3345) & (g3333) & (!g2759) & (g3359)) + ((g2283) & (g1914) & (!g3345) & (g3333) & (g2759) & (!g3359)) + ((g2283) & (g1914) & (!g3345) & (g3333) & (g2759) & (g3359)) + ((g2283) & (g1914) & (g3345) & (!g3333) & (!g2759) & (!g3359)) + ((g2283) & (g1914) & (g3345) & (!g3333) & (!g2759) & (g3359)) + ((g2283) & (g1914) & (g3345) & (!g3333) & (g2759) & (!g3359)) + ((g2283) & (g1914) & (g3345) & (!g3333) & (g2759) & (g3359)));
	assign g5675 = (((!g2288) & (!g1914) & (!g2761) & (!g3359) & (!g3345) & (!g3342)) + ((!g2288) & (!g1914) & (!g2761) & (!g3359) & (g3345) & (g3342)) + ((!g2288) & (!g1914) & (!g2761) & (g3359) & (!g3345) & (!g3342)) + ((!g2288) & (!g1914) & (!g2761) & (g3359) & (g3345) & (g3342)) + ((!g2288) & (!g1914) & (g2761) & (!g3359) & (!g3345) & (!g3342)) + ((!g2288) & (!g1914) & (g2761) & (!g3359) & (g3345) & (g3342)) + ((!g2288) & (!g1914) & (g2761) & (g3359) & (!g3345) & (!g3342)) + ((!g2288) & (!g1914) & (g2761) & (g3359) & (g3345) & (g3342)) + ((!g2288) & (g1914) & (!g2761) & (!g3359) & (!g3345) & (!g3342)) + ((!g2288) & (g1914) & (!g2761) & (!g3359) & (!g3345) & (g3342)) + ((!g2288) & (g1914) & (!g2761) & (!g3359) & (g3345) & (!g3342)) + ((!g2288) & (g1914) & (!g2761) & (!g3359) & (g3345) & (g3342)) + ((!g2288) & (g1914) & (g2761) & (g3359) & (!g3345) & (!g3342)) + ((!g2288) & (g1914) & (g2761) & (g3359) & (!g3345) & (g3342)) + ((!g2288) & (g1914) & (g2761) & (g3359) & (g3345) & (!g3342)) + ((!g2288) & (g1914) & (g2761) & (g3359) & (g3345) & (g3342)) + ((g2288) & (!g1914) & (!g2761) & (!g3359) & (!g3345) & (g3342)) + ((g2288) & (!g1914) & (!g2761) & (!g3359) & (g3345) & (!g3342)) + ((g2288) & (!g1914) & (!g2761) & (g3359) & (!g3345) & (g3342)) + ((g2288) & (!g1914) & (!g2761) & (g3359) & (g3345) & (!g3342)) + ((g2288) & (!g1914) & (g2761) & (!g3359) & (!g3345) & (g3342)) + ((g2288) & (!g1914) & (g2761) & (!g3359) & (g3345) & (!g3342)) + ((g2288) & (!g1914) & (g2761) & (g3359) & (!g3345) & (g3342)) + ((g2288) & (!g1914) & (g2761) & (g3359) & (g3345) & (!g3342)) + ((g2288) & (g1914) & (!g2761) & (g3359) & (!g3345) & (!g3342)) + ((g2288) & (g1914) & (!g2761) & (g3359) & (!g3345) & (g3342)) + ((g2288) & (g1914) & (!g2761) & (g3359) & (g3345) & (!g3342)) + ((g2288) & (g1914) & (!g2761) & (g3359) & (g3345) & (g3342)) + ((g2288) & (g1914) & (g2761) & (!g3359) & (!g3345) & (!g3342)) + ((g2288) & (g1914) & (g2761) & (!g3359) & (!g3345) & (g3342)) + ((g2288) & (g1914) & (g2761) & (!g3359) & (g3345) & (!g3342)) + ((g2288) & (g1914) & (g2761) & (!g3359) & (g3345) & (g3342)));
	assign g5676 = (((!g2434) & (!g1914) & (!g3342) & (!g3348) & (!g964) & (!g4701)) + ((!g2434) & (!g1914) & (!g3342) & (!g3348) & (!g964) & (g4701)) + ((!g2434) & (!g1914) & (!g3342) & (!g3348) & (g964) & (!g4701)) + ((!g2434) & (!g1914) & (!g3342) & (!g3348) & (g964) & (g4701)) + ((!g2434) & (!g1914) & (g3342) & (g3348) & (!g964) & (!g4701)) + ((!g2434) & (!g1914) & (g3342) & (g3348) & (!g964) & (g4701)) + ((!g2434) & (!g1914) & (g3342) & (g3348) & (g964) & (!g4701)) + ((!g2434) & (!g1914) & (g3342) & (g3348) & (g964) & (g4701)) + ((!g2434) & (g1914) & (!g3342) & (!g3348) & (!g964) & (!g4701)) + ((!g2434) & (g1914) & (!g3342) & (!g3348) & (g964) & (g4701)) + ((!g2434) & (g1914) & (!g3342) & (g3348) & (!g964) & (!g4701)) + ((!g2434) & (g1914) & (!g3342) & (g3348) & (g964) & (g4701)) + ((!g2434) & (g1914) & (g3342) & (!g3348) & (!g964) & (!g4701)) + ((!g2434) & (g1914) & (g3342) & (!g3348) & (g964) & (g4701)) + ((!g2434) & (g1914) & (g3342) & (g3348) & (!g964) & (!g4701)) + ((!g2434) & (g1914) & (g3342) & (g3348) & (g964) & (g4701)) + ((g2434) & (!g1914) & (!g3342) & (g3348) & (!g964) & (!g4701)) + ((g2434) & (!g1914) & (!g3342) & (g3348) & (!g964) & (g4701)) + ((g2434) & (!g1914) & (!g3342) & (g3348) & (g964) & (!g4701)) + ((g2434) & (!g1914) & (!g3342) & (g3348) & (g964) & (g4701)) + ((g2434) & (!g1914) & (g3342) & (!g3348) & (!g964) & (!g4701)) + ((g2434) & (!g1914) & (g3342) & (!g3348) & (!g964) & (g4701)) + ((g2434) & (!g1914) & (g3342) & (!g3348) & (g964) & (!g4701)) + ((g2434) & (!g1914) & (g3342) & (!g3348) & (g964) & (g4701)) + ((g2434) & (g1914) & (!g3342) & (!g3348) & (!g964) & (g4701)) + ((g2434) & (g1914) & (!g3342) & (!g3348) & (g964) & (!g4701)) + ((g2434) & (g1914) & (!g3342) & (g3348) & (!g964) & (g4701)) + ((g2434) & (g1914) & (!g3342) & (g3348) & (g964) & (!g4701)) + ((g2434) & (g1914) & (g3342) & (!g3348) & (!g964) & (g4701)) + ((g2434) & (g1914) & (g3342) & (!g3348) & (g964) & (!g4701)) + ((g2434) & (g1914) & (g3342) & (g3348) & (!g964) & (g4701)) + ((g2434) & (g1914) & (g3342) & (g3348) & (g964) & (!g4701)));
	assign g5677 = (((!g1968) & (!g1914) & (!g2758) & (!g3339) & (!g2173) & (!g3980)) + ((!g1968) & (!g1914) & (!g2758) & (!g3339) & (g2173) & (g3980)) + ((!g1968) & (!g1914) & (!g2758) & (g3339) & (!g2173) & (!g3980)) + ((!g1968) & (!g1914) & (!g2758) & (g3339) & (g2173) & (g3980)) + ((!g1968) & (!g1914) & (g2758) & (!g3339) & (!g2173) & (!g3980)) + ((!g1968) & (!g1914) & (g2758) & (!g3339) & (g2173) & (g3980)) + ((!g1968) & (!g1914) & (g2758) & (g3339) & (!g2173) & (!g3980)) + ((!g1968) & (!g1914) & (g2758) & (g3339) & (g2173) & (g3980)) + ((!g1968) & (g1914) & (!g2758) & (!g3339) & (!g2173) & (!g3980)) + ((!g1968) & (g1914) & (!g2758) & (!g3339) & (!g2173) & (g3980)) + ((!g1968) & (g1914) & (!g2758) & (!g3339) & (g2173) & (!g3980)) + ((!g1968) & (g1914) & (!g2758) & (!g3339) & (g2173) & (g3980)) + ((!g1968) & (g1914) & (g2758) & (g3339) & (!g2173) & (!g3980)) + ((!g1968) & (g1914) & (g2758) & (g3339) & (!g2173) & (g3980)) + ((!g1968) & (g1914) & (g2758) & (g3339) & (g2173) & (!g3980)) + ((!g1968) & (g1914) & (g2758) & (g3339) & (g2173) & (g3980)) + ((g1968) & (!g1914) & (!g2758) & (!g3339) & (!g2173) & (g3980)) + ((g1968) & (!g1914) & (!g2758) & (!g3339) & (g2173) & (!g3980)) + ((g1968) & (!g1914) & (!g2758) & (g3339) & (!g2173) & (g3980)) + ((g1968) & (!g1914) & (!g2758) & (g3339) & (g2173) & (!g3980)) + ((g1968) & (!g1914) & (g2758) & (!g3339) & (!g2173) & (g3980)) + ((g1968) & (!g1914) & (g2758) & (!g3339) & (g2173) & (!g3980)) + ((g1968) & (!g1914) & (g2758) & (g3339) & (!g2173) & (g3980)) + ((g1968) & (!g1914) & (g2758) & (g3339) & (g2173) & (!g3980)) + ((g1968) & (g1914) & (!g2758) & (g3339) & (!g2173) & (!g3980)) + ((g1968) & (g1914) & (!g2758) & (g3339) & (!g2173) & (g3980)) + ((g1968) & (g1914) & (!g2758) & (g3339) & (g2173) & (!g3980)) + ((g1968) & (g1914) & (!g2758) & (g3339) & (g2173) & (g3980)) + ((g1968) & (g1914) & (g2758) & (!g3339) & (!g2173) & (!g3980)) + ((g1968) & (g1914) & (g2758) & (!g3339) & (!g2173) & (g3980)) + ((g1968) & (g1914) & (g2758) & (!g3339) & (g2173) & (!g3980)) + ((g1968) & (g1914) & (g2758) & (!g3339) & (g2173) & (g3980)));
	assign g5678 = (((!g2456) & (!g1914) & (!g2760) & (!g3353) & (!g2159) & (!g4708)) + ((!g2456) & (!g1914) & (!g2760) & (!g3353) & (g2159) & (g4708)) + ((!g2456) & (!g1914) & (!g2760) & (g3353) & (!g2159) & (!g4708)) + ((!g2456) & (!g1914) & (!g2760) & (g3353) & (g2159) & (g4708)) + ((!g2456) & (!g1914) & (g2760) & (!g3353) & (!g2159) & (!g4708)) + ((!g2456) & (!g1914) & (g2760) & (!g3353) & (g2159) & (g4708)) + ((!g2456) & (!g1914) & (g2760) & (g3353) & (!g2159) & (!g4708)) + ((!g2456) & (!g1914) & (g2760) & (g3353) & (g2159) & (g4708)) + ((!g2456) & (g1914) & (!g2760) & (!g3353) & (!g2159) & (!g4708)) + ((!g2456) & (g1914) & (!g2760) & (!g3353) & (!g2159) & (g4708)) + ((!g2456) & (g1914) & (!g2760) & (!g3353) & (g2159) & (!g4708)) + ((!g2456) & (g1914) & (!g2760) & (!g3353) & (g2159) & (g4708)) + ((!g2456) & (g1914) & (g2760) & (g3353) & (!g2159) & (!g4708)) + ((!g2456) & (g1914) & (g2760) & (g3353) & (!g2159) & (g4708)) + ((!g2456) & (g1914) & (g2760) & (g3353) & (g2159) & (!g4708)) + ((!g2456) & (g1914) & (g2760) & (g3353) & (g2159) & (g4708)) + ((g2456) & (!g1914) & (!g2760) & (!g3353) & (!g2159) & (g4708)) + ((g2456) & (!g1914) & (!g2760) & (!g3353) & (g2159) & (!g4708)) + ((g2456) & (!g1914) & (!g2760) & (g3353) & (!g2159) & (g4708)) + ((g2456) & (!g1914) & (!g2760) & (g3353) & (g2159) & (!g4708)) + ((g2456) & (!g1914) & (g2760) & (!g3353) & (!g2159) & (g4708)) + ((g2456) & (!g1914) & (g2760) & (!g3353) & (g2159) & (!g4708)) + ((g2456) & (!g1914) & (g2760) & (g3353) & (!g2159) & (g4708)) + ((g2456) & (!g1914) & (g2760) & (g3353) & (g2159) & (!g4708)) + ((g2456) & (g1914) & (!g2760) & (g3353) & (!g2159) & (!g4708)) + ((g2456) & (g1914) & (!g2760) & (g3353) & (!g2159) & (g4708)) + ((g2456) & (g1914) & (!g2760) & (g3353) & (g2159) & (!g4708)) + ((g2456) & (g1914) & (!g2760) & (g3353) & (g2159) & (g4708)) + ((g2456) & (g1914) & (g2760) & (!g3353) & (!g2159) & (!g4708)) + ((g2456) & (g1914) & (g2760) & (!g3353) & (!g2159) & (g4708)) + ((g2456) & (g1914) & (g2760) & (!g3353) & (g2159) & (!g4708)) + ((g2456) & (g1914) & (g2760) & (!g3353) & (g2159) & (g4708)));
	assign g5679 = (((!g2462) & (!g1914) & (!g2759) & (!g3356) & (!g2156) & (!g4711)) + ((!g2462) & (!g1914) & (!g2759) & (!g3356) & (!g2156) & (g4711)) + ((!g2462) & (!g1914) & (!g2759) & (!g3356) & (g2156) & (!g4711)) + ((!g2462) & (!g1914) & (!g2759) & (!g3356) & (g2156) & (g4711)) + ((!g2462) & (!g1914) & (g2759) & (g3356) & (!g2156) & (!g4711)) + ((!g2462) & (!g1914) & (g2759) & (g3356) & (!g2156) & (g4711)) + ((!g2462) & (!g1914) & (g2759) & (g3356) & (g2156) & (!g4711)) + ((!g2462) & (!g1914) & (g2759) & (g3356) & (g2156) & (g4711)) + ((!g2462) & (g1914) & (!g2759) & (!g3356) & (!g2156) & (!g4711)) + ((!g2462) & (g1914) & (!g2759) & (!g3356) & (g2156) & (g4711)) + ((!g2462) & (g1914) & (!g2759) & (g3356) & (!g2156) & (!g4711)) + ((!g2462) & (g1914) & (!g2759) & (g3356) & (g2156) & (g4711)) + ((!g2462) & (g1914) & (g2759) & (!g3356) & (!g2156) & (!g4711)) + ((!g2462) & (g1914) & (g2759) & (!g3356) & (g2156) & (g4711)) + ((!g2462) & (g1914) & (g2759) & (g3356) & (!g2156) & (!g4711)) + ((!g2462) & (g1914) & (g2759) & (g3356) & (g2156) & (g4711)) + ((g2462) & (!g1914) & (!g2759) & (g3356) & (!g2156) & (!g4711)) + ((g2462) & (!g1914) & (!g2759) & (g3356) & (!g2156) & (g4711)) + ((g2462) & (!g1914) & (!g2759) & (g3356) & (g2156) & (!g4711)) + ((g2462) & (!g1914) & (!g2759) & (g3356) & (g2156) & (g4711)) + ((g2462) & (!g1914) & (g2759) & (!g3356) & (!g2156) & (!g4711)) + ((g2462) & (!g1914) & (g2759) & (!g3356) & (!g2156) & (g4711)) + ((g2462) & (!g1914) & (g2759) & (!g3356) & (g2156) & (!g4711)) + ((g2462) & (!g1914) & (g2759) & (!g3356) & (g2156) & (g4711)) + ((g2462) & (g1914) & (!g2759) & (!g3356) & (!g2156) & (g4711)) + ((g2462) & (g1914) & (!g2759) & (!g3356) & (g2156) & (!g4711)) + ((g2462) & (g1914) & (!g2759) & (g3356) & (!g2156) & (g4711)) + ((g2462) & (g1914) & (!g2759) & (g3356) & (g2156) & (!g4711)) + ((g2462) & (g1914) & (g2759) & (!g3356) & (!g2156) & (g4711)) + ((g2462) & (g1914) & (g2759) & (!g3356) & (g2156) & (!g4711)) + ((g2462) & (g1914) & (g2759) & (g3356) & (!g2156) & (g4711)) + ((g2462) & (g1914) & (g2759) & (g3356) & (g2156) & (!g4711)));
	assign g5680 = (((!g2468) & (!g1914) & (!g3333) & (!g3356) & (!g964) & (!g4715)) + ((!g2468) & (!g1914) & (!g3333) & (!g3356) & (g964) & (g4715)) + ((!g2468) & (!g1914) & (!g3333) & (g3356) & (!g964) & (!g4715)) + ((!g2468) & (!g1914) & (!g3333) & (g3356) & (g964) & (g4715)) + ((!g2468) & (!g1914) & (g3333) & (!g3356) & (!g964) & (!g4715)) + ((!g2468) & (!g1914) & (g3333) & (!g3356) & (g964) & (g4715)) + ((!g2468) & (!g1914) & (g3333) & (g3356) & (!g964) & (!g4715)) + ((!g2468) & (!g1914) & (g3333) & (g3356) & (g964) & (g4715)) + ((!g2468) & (g1914) & (!g3333) & (!g3356) & (!g964) & (!g4715)) + ((!g2468) & (g1914) & (!g3333) & (!g3356) & (!g964) & (g4715)) + ((!g2468) & (g1914) & (!g3333) & (!g3356) & (g964) & (!g4715)) + ((!g2468) & (g1914) & (!g3333) & (!g3356) & (g964) & (g4715)) + ((!g2468) & (g1914) & (g3333) & (g3356) & (!g964) & (!g4715)) + ((!g2468) & (g1914) & (g3333) & (g3356) & (!g964) & (g4715)) + ((!g2468) & (g1914) & (g3333) & (g3356) & (g964) & (!g4715)) + ((!g2468) & (g1914) & (g3333) & (g3356) & (g964) & (g4715)) + ((g2468) & (!g1914) & (!g3333) & (!g3356) & (!g964) & (g4715)) + ((g2468) & (!g1914) & (!g3333) & (!g3356) & (g964) & (!g4715)) + ((g2468) & (!g1914) & (!g3333) & (g3356) & (!g964) & (g4715)) + ((g2468) & (!g1914) & (!g3333) & (g3356) & (g964) & (!g4715)) + ((g2468) & (!g1914) & (g3333) & (!g3356) & (!g964) & (g4715)) + ((g2468) & (!g1914) & (g3333) & (!g3356) & (g964) & (!g4715)) + ((g2468) & (!g1914) & (g3333) & (g3356) & (!g964) & (g4715)) + ((g2468) & (!g1914) & (g3333) & (g3356) & (g964) & (!g4715)) + ((g2468) & (g1914) & (!g3333) & (g3356) & (!g964) & (!g4715)) + ((g2468) & (g1914) & (!g3333) & (g3356) & (!g964) & (g4715)) + ((g2468) & (g1914) & (!g3333) & (g3356) & (g964) & (!g4715)) + ((g2468) & (g1914) & (!g3333) & (g3356) & (g964) & (g4715)) + ((g2468) & (g1914) & (g3333) & (!g3356) & (!g964) & (!g4715)) + ((g2468) & (g1914) & (g3333) & (!g3356) & (!g964) & (g4715)) + ((g2468) & (g1914) & (g3333) & (!g3356) & (g964) & (!g4715)) + ((g2468) & (g1914) & (g3333) & (!g3356) & (g964) & (g4715)));
	assign g5681 = (((!g2474) & (!g1914) & (!g2758) & (!g3336) & (!g4717) & (!g2159)) + ((!g2474) & (!g1914) & (!g2758) & (!g3336) & (!g4717) & (g2159)) + ((!g2474) & (!g1914) & (!g2758) & (!g3336) & (g4717) & (!g2159)) + ((!g2474) & (!g1914) & (!g2758) & (!g3336) & (g4717) & (g2159)) + ((!g2474) & (!g1914) & (g2758) & (g3336) & (!g4717) & (!g2159)) + ((!g2474) & (!g1914) & (g2758) & (g3336) & (!g4717) & (g2159)) + ((!g2474) & (!g1914) & (g2758) & (g3336) & (g4717) & (!g2159)) + ((!g2474) & (!g1914) & (g2758) & (g3336) & (g4717) & (g2159)) + ((!g2474) & (g1914) & (!g2758) & (!g3336) & (!g4717) & (!g2159)) + ((!g2474) & (g1914) & (!g2758) & (!g3336) & (g4717) & (g2159)) + ((!g2474) & (g1914) & (!g2758) & (g3336) & (!g4717) & (!g2159)) + ((!g2474) & (g1914) & (!g2758) & (g3336) & (g4717) & (g2159)) + ((!g2474) & (g1914) & (g2758) & (!g3336) & (!g4717) & (!g2159)) + ((!g2474) & (g1914) & (g2758) & (!g3336) & (g4717) & (g2159)) + ((!g2474) & (g1914) & (g2758) & (g3336) & (!g4717) & (!g2159)) + ((!g2474) & (g1914) & (g2758) & (g3336) & (g4717) & (g2159)) + ((g2474) & (!g1914) & (!g2758) & (g3336) & (!g4717) & (!g2159)) + ((g2474) & (!g1914) & (!g2758) & (g3336) & (!g4717) & (g2159)) + ((g2474) & (!g1914) & (!g2758) & (g3336) & (g4717) & (!g2159)) + ((g2474) & (!g1914) & (!g2758) & (g3336) & (g4717) & (g2159)) + ((g2474) & (!g1914) & (g2758) & (!g3336) & (!g4717) & (!g2159)) + ((g2474) & (!g1914) & (g2758) & (!g3336) & (!g4717) & (g2159)) + ((g2474) & (!g1914) & (g2758) & (!g3336) & (g4717) & (!g2159)) + ((g2474) & (!g1914) & (g2758) & (!g3336) & (g4717) & (g2159)) + ((g2474) & (g1914) & (!g2758) & (!g3336) & (!g4717) & (g2159)) + ((g2474) & (g1914) & (!g2758) & (!g3336) & (g4717) & (!g2159)) + ((g2474) & (g1914) & (!g2758) & (g3336) & (!g4717) & (g2159)) + ((g2474) & (g1914) & (!g2758) & (g3336) & (g4717) & (!g2159)) + ((g2474) & (g1914) & (g2758) & (!g3336) & (!g4717) & (g2159)) + ((g2474) & (g1914) & (g2758) & (!g3336) & (g4717) & (!g2159)) + ((g2474) & (g1914) & (g2758) & (g3336) & (!g4717) & (g2159)) + ((g2474) & (g1914) & (g2758) & (g3336) & (g4717) & (!g2159)));
	assign g5682 = (((!g2004) & (!g1914) & (!g2760) & (!g3323) & (!g2150) & (!g2173)) + ((!g2004) & (!g1914) & (!g2760) & (!g3323) & (!g2150) & (g2173)) + ((!g2004) & (!g1914) & (!g2760) & (!g3323) & (g2150) & (!g2173)) + ((!g2004) & (!g1914) & (!g2760) & (!g3323) & (g2150) & (g2173)) + ((!g2004) & (!g1914) & (g2760) & (g3323) & (!g2150) & (!g2173)) + ((!g2004) & (!g1914) & (g2760) & (g3323) & (!g2150) & (g2173)) + ((!g2004) & (!g1914) & (g2760) & (g3323) & (g2150) & (!g2173)) + ((!g2004) & (!g1914) & (g2760) & (g3323) & (g2150) & (g2173)) + ((!g2004) & (g1914) & (!g2760) & (!g3323) & (!g2150) & (!g2173)) + ((!g2004) & (g1914) & (!g2760) & (!g3323) & (g2150) & (g2173)) + ((!g2004) & (g1914) & (!g2760) & (g3323) & (!g2150) & (!g2173)) + ((!g2004) & (g1914) & (!g2760) & (g3323) & (g2150) & (g2173)) + ((!g2004) & (g1914) & (g2760) & (!g3323) & (!g2150) & (!g2173)) + ((!g2004) & (g1914) & (g2760) & (!g3323) & (g2150) & (g2173)) + ((!g2004) & (g1914) & (g2760) & (g3323) & (!g2150) & (!g2173)) + ((!g2004) & (g1914) & (g2760) & (g3323) & (g2150) & (g2173)) + ((g2004) & (!g1914) & (!g2760) & (g3323) & (!g2150) & (!g2173)) + ((g2004) & (!g1914) & (!g2760) & (g3323) & (!g2150) & (g2173)) + ((g2004) & (!g1914) & (!g2760) & (g3323) & (g2150) & (!g2173)) + ((g2004) & (!g1914) & (!g2760) & (g3323) & (g2150) & (g2173)) + ((g2004) & (!g1914) & (g2760) & (!g3323) & (!g2150) & (!g2173)) + ((g2004) & (!g1914) & (g2760) & (!g3323) & (!g2150) & (g2173)) + ((g2004) & (!g1914) & (g2760) & (!g3323) & (g2150) & (!g2173)) + ((g2004) & (!g1914) & (g2760) & (!g3323) & (g2150) & (g2173)) + ((g2004) & (g1914) & (!g2760) & (!g3323) & (!g2150) & (g2173)) + ((g2004) & (g1914) & (!g2760) & (!g3323) & (g2150) & (!g2173)) + ((g2004) & (g1914) & (!g2760) & (g3323) & (!g2150) & (g2173)) + ((g2004) & (g1914) & (!g2760) & (g3323) & (g2150) & (!g2173)) + ((g2004) & (g1914) & (g2760) & (!g3323) & (!g2150) & (g2173)) + ((g2004) & (g1914) & (g2760) & (!g3323) & (g2150) & (!g2173)) + ((g2004) & (g1914) & (g2760) & (g3323) & (!g2150) & (g2173)) + ((g2004) & (g1914) & (g2760) & (g3323) & (g2150) & (!g2173)));
	assign g5683 = (((!g2497) & (!g1914) & (!g2761) & (!g3348) & (!g2147) & (!g4729)) + ((!g2497) & (!g1914) & (!g2761) & (!g3348) & (g2147) & (g4729)) + ((!g2497) & (!g1914) & (!g2761) & (g3348) & (!g2147) & (!g4729)) + ((!g2497) & (!g1914) & (!g2761) & (g3348) & (g2147) & (g4729)) + ((!g2497) & (!g1914) & (g2761) & (!g3348) & (!g2147) & (!g4729)) + ((!g2497) & (!g1914) & (g2761) & (!g3348) & (g2147) & (g4729)) + ((!g2497) & (!g1914) & (g2761) & (g3348) & (!g2147) & (!g4729)) + ((!g2497) & (!g1914) & (g2761) & (g3348) & (g2147) & (g4729)) + ((!g2497) & (g1914) & (!g2761) & (!g3348) & (!g2147) & (!g4729)) + ((!g2497) & (g1914) & (!g2761) & (!g3348) & (!g2147) & (g4729)) + ((!g2497) & (g1914) & (!g2761) & (!g3348) & (g2147) & (!g4729)) + ((!g2497) & (g1914) & (!g2761) & (!g3348) & (g2147) & (g4729)) + ((!g2497) & (g1914) & (g2761) & (g3348) & (!g2147) & (!g4729)) + ((!g2497) & (g1914) & (g2761) & (g3348) & (!g2147) & (g4729)) + ((!g2497) & (g1914) & (g2761) & (g3348) & (g2147) & (!g4729)) + ((!g2497) & (g1914) & (g2761) & (g3348) & (g2147) & (g4729)) + ((g2497) & (!g1914) & (!g2761) & (!g3348) & (!g2147) & (g4729)) + ((g2497) & (!g1914) & (!g2761) & (!g3348) & (g2147) & (!g4729)) + ((g2497) & (!g1914) & (!g2761) & (g3348) & (!g2147) & (g4729)) + ((g2497) & (!g1914) & (!g2761) & (g3348) & (g2147) & (!g4729)) + ((g2497) & (!g1914) & (g2761) & (!g3348) & (!g2147) & (g4729)) + ((g2497) & (!g1914) & (g2761) & (!g3348) & (g2147) & (!g4729)) + ((g2497) & (!g1914) & (g2761) & (g3348) & (!g2147) & (g4729)) + ((g2497) & (!g1914) & (g2761) & (g3348) & (g2147) & (!g4729)) + ((g2497) & (g1914) & (!g2761) & (g3348) & (!g2147) & (!g4729)) + ((g2497) & (g1914) & (!g2761) & (g3348) & (!g2147) & (g4729)) + ((g2497) & (g1914) & (!g2761) & (g3348) & (g2147) & (!g4729)) + ((g2497) & (g1914) & (!g2761) & (g3348) & (g2147) & (g4729)) + ((g2497) & (g1914) & (g2761) & (!g3348) & (!g2147) & (!g4729)) + ((g2497) & (g1914) & (g2761) & (!g3348) & (!g2147) & (g4729)) + ((g2497) & (g1914) & (g2761) & (!g3348) & (g2147) & (!g4729)) + ((g2497) & (g1914) & (g2761) & (!g3348) & (g2147) & (g4729)));
	assign g5684 = (((!g2649) & (!g2650)) + ((g2649) & (g2650)));
	assign g5685 = (((!g2647) & (!g3240)) + ((g2647) & (g3240)));
	assign g5686 = (((!g3250) & (!g3265)) + ((g3250) & (g3265)));
	assign g5687 = (((!g3274) & (!g3279)) + ((g3274) & (g3279)));
	assign g5688 = (((!g1914) & (!g1337) & (!g2683) & (!g2684) & (!g2678) & (!g2679)) + ((!g1914) & (!g1337) & (!g2683) & (!g2684) & (!g2678) & (g2679)) + ((!g1914) & (!g1337) & (!g2683) & (!g2684) & (g2678) & (!g2679)) + ((!g1914) & (!g1337) & (!g2683) & (!g2684) & (g2678) & (g2679)) + ((!g1914) & (!g1337) & (g2683) & (g2684) & (!g2678) & (!g2679)) + ((!g1914) & (!g1337) & (g2683) & (g2684) & (!g2678) & (g2679)) + ((!g1914) & (!g1337) & (g2683) & (g2684) & (g2678) & (!g2679)) + ((!g1914) & (!g1337) & (g2683) & (g2684) & (g2678) & (g2679)) + ((!g1914) & (g1337) & (!g2683) & (g2684) & (!g2678) & (!g2679)) + ((!g1914) & (g1337) & (!g2683) & (g2684) & (!g2678) & (g2679)) + ((!g1914) & (g1337) & (!g2683) & (g2684) & (g2678) & (!g2679)) + ((!g1914) & (g1337) & (!g2683) & (g2684) & (g2678) & (g2679)) + ((!g1914) & (g1337) & (g2683) & (!g2684) & (!g2678) & (!g2679)) + ((!g1914) & (g1337) & (g2683) & (!g2684) & (!g2678) & (g2679)) + ((!g1914) & (g1337) & (g2683) & (!g2684) & (g2678) & (!g2679)) + ((!g1914) & (g1337) & (g2683) & (!g2684) & (g2678) & (g2679)) + ((g1914) & (!g1337) & (!g2683) & (!g2684) & (!g2678) & (!g2679)) + ((g1914) & (!g1337) & (!g2683) & (!g2684) & (g2678) & (g2679)) + ((g1914) & (!g1337) & (!g2683) & (g2684) & (!g2678) & (!g2679)) + ((g1914) & (!g1337) & (!g2683) & (g2684) & (g2678) & (g2679)) + ((g1914) & (!g1337) & (g2683) & (!g2684) & (!g2678) & (!g2679)) + ((g1914) & (!g1337) & (g2683) & (!g2684) & (g2678) & (g2679)) + ((g1914) & (!g1337) & (g2683) & (g2684) & (!g2678) & (!g2679)) + ((g1914) & (!g1337) & (g2683) & (g2684) & (g2678) & (g2679)) + ((g1914) & (g1337) & (!g2683) & (!g2684) & (!g2678) & (g2679)) + ((g1914) & (g1337) & (!g2683) & (!g2684) & (g2678) & (!g2679)) + ((g1914) & (g1337) & (!g2683) & (g2684) & (!g2678) & (g2679)) + ((g1914) & (g1337) & (!g2683) & (g2684) & (g2678) & (!g2679)) + ((g1914) & (g1337) & (g2683) & (!g2684) & (!g2678) & (g2679)) + ((g1914) & (g1337) & (g2683) & (!g2684) & (g2678) & (!g2679)) + ((g1914) & (g1337) & (g2683) & (g2684) & (!g2678) & (g2679)) + ((g1914) & (g1337) & (g2683) & (g2684) & (g2678) & (!g2679)));
	assign g5689 = (((!g1914) & (!g2682) & (!g2648) & (!g5688)) + ((!g1914) & (!g2682) & (g2648) & (!g5688)) + ((!g1914) & (g2682) & (!g2648) & (g5688)) + ((!g1914) & (g2682) & (g2648) & (g5688)) + ((g1914) & (!g2682) & (!g2648) & (!g5688)) + ((g1914) & (!g2682) & (g2648) & (g5688)) + ((g1914) & (g2682) & (!g2648) & (!g5688)) + ((g1914) & (g2682) & (g2648) & (g5688)));
	assign g5690 = (((!g2646) & (!g2647) & (!g5688) & (!g5689)) + ((!g2646) & (!g2647) & (!g5688) & (g5689)) + ((!g2646) & (g2647) & (!g5688) & (g5689)) + ((!g2646) & (g2647) & (g5688) & (g5689)) + ((g2646) & (!g2647) & (!g5688) & (g5689)) + ((g2646) & (!g2647) & (g5688) & (g5689)) + ((g2646) & (g2647) & (g5688) & (!g5689)) + ((g2646) & (g2647) & (g5688) & (g5689)));
	assign g5691 = (((!g1914) & (!g1370) & (!g2760) & (!g2761) & (!g2759)) + ((!g1914) & (!g1370) & (!g2760) & (!g2761) & (g2759)) + ((!g1914) & (!g1370) & (g2760) & (g2761) & (!g2759)) + ((!g1914) & (!g1370) & (g2760) & (g2761) & (g2759)) + ((!g1914) & (g1370) & (!g2760) & (g2761) & (!g2759)) + ((!g1914) & (g1370) & (!g2760) & (g2761) & (g2759)) + ((!g1914) & (g1370) & (g2760) & (!g2761) & (!g2759)) + ((!g1914) & (g1370) & (g2760) & (!g2761) & (g2759)) + ((g1914) & (!g1370) & (!g2760) & (!g2761) & (g2759)) + ((g1914) & (!g1370) & (!g2760) & (g2761) & (g2759)) + ((g1914) & (!g1370) & (g2760) & (!g2761) & (g2759)) + ((g1914) & (!g1370) & (g2760) & (g2761) & (g2759)) + ((g1914) & (g1370) & (!g2760) & (!g2761) & (!g2759)) + ((g1914) & (g1370) & (!g2760) & (g2761) & (!g2759)) + ((g1914) & (g1370) & (g2760) & (!g2761) & (!g2759)) + ((g1914) & (g1370) & (g2760) & (g2761) & (!g2759)));
	assign g5692 = (((!g1914) & (!g2682) & (!g2683) & (!g2684) & (!g2758) & (!g5691)) + ((!g1914) & (!g2682) & (!g2683) & (!g2684) & (g2758) & (!g5691)) + ((!g1914) & (!g2682) & (!g2683) & (g2684) & (!g2758) & (!g5691)) + ((!g1914) & (!g2682) & (!g2683) & (g2684) & (g2758) & (!g5691)) + ((!g1914) & (!g2682) & (g2683) & (!g2684) & (!g2758) & (!g5691)) + ((!g1914) & (!g2682) & (g2683) & (!g2684) & (g2758) & (!g5691)) + ((!g1914) & (!g2682) & (g2683) & (g2684) & (!g2758) & (g5691)) + ((!g1914) & (!g2682) & (g2683) & (g2684) & (g2758) & (g5691)) + ((!g1914) & (g2682) & (!g2683) & (!g2684) & (!g2758) & (!g5691)) + ((!g1914) & (g2682) & (!g2683) & (!g2684) & (g2758) & (!g5691)) + ((!g1914) & (g2682) & (!g2683) & (g2684) & (!g2758) & (g5691)) + ((!g1914) & (g2682) & (!g2683) & (g2684) & (g2758) & (g5691)) + ((!g1914) & (g2682) & (g2683) & (!g2684) & (!g2758) & (g5691)) + ((!g1914) & (g2682) & (g2683) & (!g2684) & (g2758) & (g5691)) + ((!g1914) & (g2682) & (g2683) & (g2684) & (!g2758) & (g5691)) + ((!g1914) & (g2682) & (g2683) & (g2684) & (g2758) & (g5691)) + ((g1914) & (!g2682) & (!g2683) & (!g2684) & (!g2758) & (!g5691)) + ((g1914) & (!g2682) & (!g2683) & (!g2684) & (g2758) & (g5691)) + ((g1914) & (!g2682) & (!g2683) & (g2684) & (!g2758) & (!g5691)) + ((g1914) & (!g2682) & (!g2683) & (g2684) & (g2758) & (g5691)) + ((g1914) & (!g2682) & (g2683) & (!g2684) & (!g2758) & (!g5691)) + ((g1914) & (!g2682) & (g2683) & (!g2684) & (g2758) & (g5691)) + ((g1914) & (!g2682) & (g2683) & (g2684) & (!g2758) & (!g5691)) + ((g1914) & (!g2682) & (g2683) & (g2684) & (g2758) & (g5691)) + ((g1914) & (g2682) & (!g2683) & (!g2684) & (!g2758) & (!g5691)) + ((g1914) & (g2682) & (!g2683) & (!g2684) & (g2758) & (g5691)) + ((g1914) & (g2682) & (!g2683) & (g2684) & (!g2758) & (!g5691)) + ((g1914) & (g2682) & (!g2683) & (g2684) & (g2758) & (g5691)) + ((g1914) & (g2682) & (g2683) & (!g2684) & (!g2758) & (!g5691)) + ((g1914) & (g2682) & (g2683) & (!g2684) & (g2758) & (g5691)) + ((g1914) & (g2682) & (g2683) & (g2684) & (!g2758) & (!g5691)) + ((g1914) & (g2682) & (g2683) & (g2684) & (g2758) & (g5691)));
	assign g5693 = (((!g2683) & (!g2684) & (!g5691) & (g5692)) + ((!g2683) & (!g2684) & (g5691) & (g5692)) + ((!g2683) & (g2684) & (g5691) & (!g5692)) + ((!g2683) & (g2684) & (g5691) & (g5692)) + ((g2683) & (!g2684) & (g5691) & (!g5692)) + ((g2683) & (!g2684) & (g5691) & (g5692)) + ((g2683) & (g2684) & (g5691) & (!g5692)) + ((g2683) & (g2684) & (g5691) & (g5692)));
	assign g5694 = (((!g1914) & (!g2523) & (!g3382) & (!g1985) & (g964) & (g4715)) + ((!g1914) & (!g2523) & (!g3382) & (g1985) & (!g964) & (g4715)) + ((!g1914) & (!g2523) & (!g3382) & (g1985) & (g964) & (!g4715)) + ((!g1914) & (!g2523) & (!g3382) & (g1985) & (g964) & (g4715)) + ((!g1914) & (!g2523) & (g3382) & (!g1985) & (g964) & (g4715)) + ((!g1914) & (!g2523) & (g3382) & (g1985) & (!g964) & (g4715)) + ((!g1914) & (!g2523) & (g3382) & (g1985) & (g964) & (!g4715)) + ((!g1914) & (!g2523) & (g3382) & (g1985) & (g964) & (g4715)) + ((!g1914) & (g2523) & (!g3382) & (!g1985) & (!g964) & (!g4715)) + ((!g1914) & (g2523) & (!g3382) & (!g1985) & (!g964) & (g4715)) + ((!g1914) & (g2523) & (!g3382) & (!g1985) & (g964) & (!g4715)) + ((!g1914) & (g2523) & (!g3382) & (g1985) & (!g964) & (!g4715)) + ((!g1914) & (g2523) & (g3382) & (!g1985) & (!g964) & (!g4715)) + ((!g1914) & (g2523) & (g3382) & (!g1985) & (!g964) & (g4715)) + ((!g1914) & (g2523) & (g3382) & (!g1985) & (g964) & (!g4715)) + ((!g1914) & (g2523) & (g3382) & (g1985) & (!g964) & (!g4715)) + ((g1914) & (!g2523) & (g3382) & (!g1985) & (!g964) & (!g4715)) + ((g1914) & (!g2523) & (g3382) & (!g1985) & (!g964) & (g4715)) + ((g1914) & (!g2523) & (g3382) & (!g1985) & (g964) & (!g4715)) + ((g1914) & (!g2523) & (g3382) & (!g1985) & (g964) & (g4715)) + ((g1914) & (!g2523) & (g3382) & (g1985) & (!g964) & (!g4715)) + ((g1914) & (!g2523) & (g3382) & (g1985) & (!g964) & (g4715)) + ((g1914) & (!g2523) & (g3382) & (g1985) & (g964) & (!g4715)) + ((g1914) & (!g2523) & (g3382) & (g1985) & (g964) & (g4715)) + ((g1914) & (g2523) & (!g3382) & (!g1985) & (!g964) & (!g4715)) + ((g1914) & (g2523) & (!g3382) & (!g1985) & (!g964) & (g4715)) + ((g1914) & (g2523) & (!g3382) & (!g1985) & (g964) & (!g4715)) + ((g1914) & (g2523) & (!g3382) & (!g1985) & (g964) & (g4715)) + ((g1914) & (g2523) & (!g3382) & (g1985) & (!g964) & (!g4715)) + ((g1914) & (g2523) & (!g3382) & (g1985) & (!g964) & (g4715)) + ((g1914) & (g2523) & (!g3382) & (g1985) & (g964) & (!g4715)) + ((g1914) & (g2523) & (!g3382) & (g1985) & (g964) & (g4715)));
	assign g5695 = (((!g1914) & (!g3378) & (!g1987) & (!g998) & (g5694)) + ((!g1914) & (!g3378) & (!g1987) & (g998) & (!g5694)) + ((!g1914) & (!g3378) & (g1987) & (!g998) & (!g5694)) + ((!g1914) & (!g3378) & (g1987) & (g998) & (g5694)) + ((!g1914) & (g3378) & (!g1987) & (!g998) & (g5694)) + ((!g1914) & (g3378) & (!g1987) & (g998) & (!g5694)) + ((!g1914) & (g3378) & (g1987) & (!g998) & (!g5694)) + ((!g1914) & (g3378) & (g1987) & (g998) & (g5694)) + ((g1914) & (!g3378) & (!g1987) & (!g998) & (!g5694)) + ((g1914) & (!g3378) & (!g1987) & (g998) & (!g5694)) + ((g1914) & (!g3378) & (g1987) & (!g998) & (!g5694)) + ((g1914) & (!g3378) & (g1987) & (g998) & (!g5694)) + ((g1914) & (g3378) & (!g1987) & (!g998) & (g5694)) + ((g1914) & (g3378) & (!g1987) & (g998) & (g5694)) + ((g1914) & (g3378) & (g1987) & (!g998) & (g5694)) + ((g1914) & (g3378) & (g1987) & (g998) & (g5694)));
	assign g5696 = (((!g1914) & (!g2006) & (g3376) & (!g4093) & (!g2150) & (!g2173)) + ((!g1914) & (!g2006) & (g3376) & (!g4093) & (!g2150) & (g2173)) + ((!g1914) & (!g2006) & (g3376) & (!g4093) & (g2150) & (!g2173)) + ((!g1914) & (!g2006) & (g3376) & (!g4093) & (g2150) & (g2173)) + ((!g1914) & (!g2006) & (g3376) & (g4093) & (!g2150) & (!g2173)) + ((!g1914) & (!g2006) & (g3376) & (g4093) & (!g2150) & (g2173)) + ((!g1914) & (!g2006) & (g3376) & (g4093) & (g2150) & (!g2173)) + ((!g1914) & (!g2006) & (g3376) & (g4093) & (g2150) & (g2173)) + ((!g1914) & (g2006) & (!g3376) & (!g4093) & (!g2150) & (!g2173)) + ((!g1914) & (g2006) & (!g3376) & (!g4093) & (!g2150) & (g2173)) + ((!g1914) & (g2006) & (!g3376) & (!g4093) & (g2150) & (!g2173)) + ((!g1914) & (g2006) & (!g3376) & (!g4093) & (g2150) & (g2173)) + ((!g1914) & (g2006) & (!g3376) & (g4093) & (!g2150) & (!g2173)) + ((!g1914) & (g2006) & (!g3376) & (g4093) & (!g2150) & (g2173)) + ((!g1914) & (g2006) & (!g3376) & (g4093) & (g2150) & (!g2173)) + ((!g1914) & (g2006) & (!g3376) & (g4093) & (g2150) & (g2173)) + ((g1914) & (!g2006) & (!g3376) & (!g4093) & (g2150) & (g2173)) + ((g1914) & (!g2006) & (!g3376) & (g4093) & (!g2150) & (g2173)) + ((g1914) & (!g2006) & (!g3376) & (g4093) & (g2150) & (!g2173)) + ((g1914) & (!g2006) & (!g3376) & (g4093) & (g2150) & (g2173)) + ((g1914) & (!g2006) & (g3376) & (!g4093) & (g2150) & (g2173)) + ((g1914) & (!g2006) & (g3376) & (g4093) & (!g2150) & (g2173)) + ((g1914) & (!g2006) & (g3376) & (g4093) & (g2150) & (!g2173)) + ((g1914) & (!g2006) & (g3376) & (g4093) & (g2150) & (g2173)) + ((g1914) & (g2006) & (!g3376) & (!g4093) & (!g2150) & (!g2173)) + ((g1914) & (g2006) & (!g3376) & (!g4093) & (!g2150) & (g2173)) + ((g1914) & (g2006) & (!g3376) & (!g4093) & (g2150) & (!g2173)) + ((g1914) & (g2006) & (!g3376) & (g4093) & (!g2150) & (!g2173)) + ((g1914) & (g2006) & (g3376) & (!g4093) & (!g2150) & (!g2173)) + ((g1914) & (g2006) & (g3376) & (!g4093) & (!g2150) & (g2173)) + ((g1914) & (g2006) & (g3376) & (!g4093) & (g2150) & (!g2173)) + ((g1914) & (g2006) & (g3376) & (g4093) & (!g2150) & (!g2173)));
	assign g5697 = (((!g1914) & (!g2793) & (!g2203) & (!g2207) & (!g5696)) + ((!g1914) & (!g2793) & (!g2203) & (g2207) & (!g5696)) + ((!g1914) & (!g2793) & (g2203) & (!g2207) & (!g5696)) + ((!g1914) & (!g2793) & (g2203) & (g2207) & (!g5696)) + ((!g1914) & (g2793) & (!g2203) & (!g2207) & (g5696)) + ((!g1914) & (g2793) & (!g2203) & (g2207) & (g5696)) + ((!g1914) & (g2793) & (g2203) & (!g2207) & (g5696)) + ((!g1914) & (g2793) & (g2203) & (g2207) & (g5696)) + ((g1914) & (!g2793) & (!g2203) & (!g2207) & (g5696)) + ((g1914) & (!g2793) & (!g2203) & (g2207) & (!g5696)) + ((g1914) & (!g2793) & (g2203) & (!g2207) & (!g5696)) + ((g1914) & (!g2793) & (g2203) & (g2207) & (g5696)) + ((g1914) & (g2793) & (!g2203) & (!g2207) & (g5696)) + ((g1914) & (g2793) & (!g2203) & (g2207) & (!g5696)) + ((g1914) & (g2793) & (g2203) & (!g2207) & (!g5696)) + ((g1914) & (g2793) & (g2203) & (g2207) & (g5696)));
	assign g5698 = (((!g1914) & (!g2529) & (g3385) & (!g2137) & (!g4717) & (!g2159)) + ((!g1914) & (!g2529) & (g3385) & (!g2137) & (!g4717) & (g2159)) + ((!g1914) & (!g2529) & (g3385) & (!g2137) & (g4717) & (!g2159)) + ((!g1914) & (!g2529) & (g3385) & (!g2137) & (g4717) & (g2159)) + ((!g1914) & (!g2529) & (g3385) & (g2137) & (!g4717) & (!g2159)) + ((!g1914) & (!g2529) & (g3385) & (g2137) & (!g4717) & (g2159)) + ((!g1914) & (!g2529) & (g3385) & (g2137) & (g4717) & (!g2159)) + ((!g1914) & (!g2529) & (g3385) & (g2137) & (g4717) & (g2159)) + ((!g1914) & (g2529) & (!g3385) & (!g2137) & (!g4717) & (!g2159)) + ((!g1914) & (g2529) & (!g3385) & (!g2137) & (!g4717) & (g2159)) + ((!g1914) & (g2529) & (!g3385) & (!g2137) & (g4717) & (!g2159)) + ((!g1914) & (g2529) & (!g3385) & (!g2137) & (g4717) & (g2159)) + ((!g1914) & (g2529) & (!g3385) & (g2137) & (!g4717) & (!g2159)) + ((!g1914) & (g2529) & (!g3385) & (g2137) & (!g4717) & (g2159)) + ((!g1914) & (g2529) & (!g3385) & (g2137) & (g4717) & (!g2159)) + ((!g1914) & (g2529) & (!g3385) & (g2137) & (g4717) & (g2159)) + ((g1914) & (!g2529) & (!g3385) & (!g2137) & (g4717) & (g2159)) + ((g1914) & (!g2529) & (!g3385) & (g2137) & (!g4717) & (g2159)) + ((g1914) & (!g2529) & (!g3385) & (g2137) & (g4717) & (!g2159)) + ((g1914) & (!g2529) & (!g3385) & (g2137) & (g4717) & (g2159)) + ((g1914) & (!g2529) & (g3385) & (!g2137) & (g4717) & (g2159)) + ((g1914) & (!g2529) & (g3385) & (g2137) & (!g4717) & (g2159)) + ((g1914) & (!g2529) & (g3385) & (g2137) & (g4717) & (!g2159)) + ((g1914) & (!g2529) & (g3385) & (g2137) & (g4717) & (g2159)) + ((g1914) & (g2529) & (!g3385) & (!g2137) & (!g4717) & (!g2159)) + ((g1914) & (g2529) & (!g3385) & (!g2137) & (!g4717) & (g2159)) + ((g1914) & (g2529) & (!g3385) & (!g2137) & (g4717) & (!g2159)) + ((g1914) & (g2529) & (!g3385) & (g2137) & (!g4717) & (!g2159)) + ((g1914) & (g2529) & (g3385) & (!g2137) & (!g4717) & (!g2159)) + ((g1914) & (g2529) & (g3385) & (!g2137) & (!g4717) & (g2159)) + ((g1914) & (g2529) & (g3385) & (!g2137) & (g4717) & (!g2159)) + ((g1914) & (g2529) & (g3385) & (g2137) & (!g4717) & (!g2159)));
	assign g5699 = (((!g1914) & (!g2789) & (!g2194) & (!g2198) & (!g5698)) + ((!g1914) & (!g2789) & (!g2194) & (g2198) & (!g5698)) + ((!g1914) & (!g2789) & (g2194) & (!g2198) & (!g5698)) + ((!g1914) & (!g2789) & (g2194) & (g2198) & (!g5698)) + ((!g1914) & (g2789) & (!g2194) & (!g2198) & (g5698)) + ((!g1914) & (g2789) & (!g2194) & (g2198) & (g5698)) + ((!g1914) & (g2789) & (g2194) & (!g2198) & (g5698)) + ((!g1914) & (g2789) & (g2194) & (g2198) & (g5698)) + ((g1914) & (!g2789) & (!g2194) & (!g2198) & (g5698)) + ((g1914) & (!g2789) & (!g2194) & (g2198) & (!g5698)) + ((g1914) & (!g2789) & (g2194) & (!g2198) & (!g5698)) + ((g1914) & (!g2789) & (g2194) & (g2198) & (g5698)) + ((g1914) & (g2789) & (!g2194) & (!g2198) & (g5698)) + ((g1914) & (g2789) & (!g2194) & (g2198) & (!g5698)) + ((g1914) & (g2789) & (g2194) & (!g2198) & (!g5698)) + ((g1914) & (g2789) & (g2194) & (g2198) & (g5698)));
	assign g5700 = (((!g1914) & (!g2531) & (!g3387) & (!g2144) & (g2147) & (g4729)) + ((!g1914) & (!g2531) & (!g3387) & (g2144) & (!g2147) & (g4729)) + ((!g1914) & (!g2531) & (!g3387) & (g2144) & (g2147) & (!g4729)) + ((!g1914) & (!g2531) & (!g3387) & (g2144) & (g2147) & (g4729)) + ((!g1914) & (!g2531) & (g3387) & (!g2144) & (g2147) & (g4729)) + ((!g1914) & (!g2531) & (g3387) & (g2144) & (!g2147) & (g4729)) + ((!g1914) & (!g2531) & (g3387) & (g2144) & (g2147) & (!g4729)) + ((!g1914) & (!g2531) & (g3387) & (g2144) & (g2147) & (g4729)) + ((!g1914) & (g2531) & (!g3387) & (!g2144) & (!g2147) & (!g4729)) + ((!g1914) & (g2531) & (!g3387) & (!g2144) & (!g2147) & (g4729)) + ((!g1914) & (g2531) & (!g3387) & (!g2144) & (g2147) & (!g4729)) + ((!g1914) & (g2531) & (!g3387) & (g2144) & (!g2147) & (!g4729)) + ((!g1914) & (g2531) & (g3387) & (!g2144) & (!g2147) & (!g4729)) + ((!g1914) & (g2531) & (g3387) & (!g2144) & (!g2147) & (g4729)) + ((!g1914) & (g2531) & (g3387) & (!g2144) & (g2147) & (!g4729)) + ((!g1914) & (g2531) & (g3387) & (g2144) & (!g2147) & (!g4729)) + ((g1914) & (!g2531) & (g3387) & (!g2144) & (!g2147) & (!g4729)) + ((g1914) & (!g2531) & (g3387) & (!g2144) & (!g2147) & (g4729)) + ((g1914) & (!g2531) & (g3387) & (!g2144) & (g2147) & (!g4729)) + ((g1914) & (!g2531) & (g3387) & (!g2144) & (g2147) & (g4729)) + ((g1914) & (!g2531) & (g3387) & (g2144) & (!g2147) & (!g4729)) + ((g1914) & (!g2531) & (g3387) & (g2144) & (!g2147) & (g4729)) + ((g1914) & (!g2531) & (g3387) & (g2144) & (g2147) & (!g4729)) + ((g1914) & (!g2531) & (g3387) & (g2144) & (g2147) & (g4729)) + ((g1914) & (g2531) & (!g3387) & (!g2144) & (!g2147) & (!g4729)) + ((g1914) & (g2531) & (!g3387) & (!g2144) & (!g2147) & (g4729)) + ((g1914) & (g2531) & (!g3387) & (!g2144) & (g2147) & (!g4729)) + ((g1914) & (g2531) & (!g3387) & (!g2144) & (g2147) & (g4729)) + ((g1914) & (g2531) & (!g3387) & (g2144) & (!g2147) & (!g4729)) + ((g1914) & (g2531) & (!g3387) & (g2144) & (!g2147) & (g4729)) + ((g1914) & (g2531) & (!g3387) & (g2144) & (g2147) & (!g4729)) + ((g1914) & (g2531) & (!g3387) & (g2144) & (g2147) & (g4729)));
	assign g5701 = (((!g1914) & (!g2794) & (!g2188) & (!g2196) & (g5700)) + ((!g1914) & (!g2794) & (!g2188) & (g2196) & (!g5700)) + ((!g1914) & (!g2794) & (g2188) & (!g2196) & (!g5700)) + ((!g1914) & (!g2794) & (g2188) & (g2196) & (g5700)) + ((!g1914) & (g2794) & (!g2188) & (!g2196) & (g5700)) + ((!g1914) & (g2794) & (!g2188) & (g2196) & (!g5700)) + ((!g1914) & (g2794) & (g2188) & (!g2196) & (!g5700)) + ((!g1914) & (g2794) & (g2188) & (g2196) & (g5700)) + ((g1914) & (!g2794) & (!g2188) & (!g2196) & (!g5700)) + ((g1914) & (!g2794) & (!g2188) & (g2196) & (!g5700)) + ((g1914) & (!g2794) & (g2188) & (!g2196) & (!g5700)) + ((g1914) & (!g2794) & (g2188) & (g2196) & (!g5700)) + ((g1914) & (g2794) & (!g2188) & (!g2196) & (g5700)) + ((g1914) & (g2794) & (!g2188) & (g2196) & (g5700)) + ((g1914) & (g2794) & (g2188) & (!g2196) & (g5700)) + ((g1914) & (g2794) & (g2188) & (g2196) & (g5700)));
	assign g5702 = (((!g1914) & (!g2533) & (g3387) & (!g1947) & (!g964) & (!g4701)) + ((!g1914) & (!g2533) & (g3387) & (!g1947) & (!g964) & (g4701)) + ((!g1914) & (!g2533) & (g3387) & (!g1947) & (g964) & (!g4701)) + ((!g1914) & (!g2533) & (g3387) & (!g1947) & (g964) & (g4701)) + ((!g1914) & (!g2533) & (g3387) & (g1947) & (!g964) & (!g4701)) + ((!g1914) & (!g2533) & (g3387) & (g1947) & (!g964) & (g4701)) + ((!g1914) & (!g2533) & (g3387) & (g1947) & (g964) & (!g4701)) + ((!g1914) & (!g2533) & (g3387) & (g1947) & (g964) & (g4701)) + ((!g1914) & (g2533) & (!g3387) & (!g1947) & (!g964) & (!g4701)) + ((!g1914) & (g2533) & (!g3387) & (!g1947) & (!g964) & (g4701)) + ((!g1914) & (g2533) & (!g3387) & (!g1947) & (g964) & (!g4701)) + ((!g1914) & (g2533) & (!g3387) & (!g1947) & (g964) & (g4701)) + ((!g1914) & (g2533) & (!g3387) & (g1947) & (!g964) & (!g4701)) + ((!g1914) & (g2533) & (!g3387) & (g1947) & (!g964) & (g4701)) + ((!g1914) & (g2533) & (!g3387) & (g1947) & (g964) & (!g4701)) + ((!g1914) & (g2533) & (!g3387) & (g1947) & (g964) & (g4701)) + ((g1914) & (!g2533) & (!g3387) & (!g1947) & (g964) & (g4701)) + ((g1914) & (!g2533) & (!g3387) & (g1947) & (!g964) & (g4701)) + ((g1914) & (!g2533) & (!g3387) & (g1947) & (g964) & (!g4701)) + ((g1914) & (!g2533) & (!g3387) & (g1947) & (g964) & (g4701)) + ((g1914) & (!g2533) & (g3387) & (!g1947) & (g964) & (g4701)) + ((g1914) & (!g2533) & (g3387) & (g1947) & (!g964) & (g4701)) + ((g1914) & (!g2533) & (g3387) & (g1947) & (g964) & (!g4701)) + ((g1914) & (!g2533) & (g3387) & (g1947) & (g964) & (g4701)) + ((g1914) & (g2533) & (!g3387) & (!g1947) & (!g964) & (!g4701)) + ((g1914) & (g2533) & (!g3387) & (!g1947) & (!g964) & (g4701)) + ((g1914) & (g2533) & (!g3387) & (!g1947) & (g964) & (!g4701)) + ((g1914) & (g2533) & (!g3387) & (g1947) & (!g964) & (!g4701)) + ((g1914) & (g2533) & (g3387) & (!g1947) & (!g964) & (!g4701)) + ((g1914) & (g2533) & (g3387) & (!g1947) & (!g964) & (g4701)) + ((g1914) & (g2533) & (g3387) & (!g1947) & (g964) & (!g4701)) + ((g1914) & (g2533) & (g3387) & (g1947) & (!g964) & (!g4701)));
	assign g5703 = (((!g1914) & (!g3372) & (!g1949) & (!g998) & (!g5702)) + ((!g1914) & (!g3372) & (!g1949) & (g998) & (!g5702)) + ((!g1914) & (!g3372) & (g1949) & (!g998) & (!g5702)) + ((!g1914) & (!g3372) & (g1949) & (g998) & (!g5702)) + ((!g1914) & (g3372) & (!g1949) & (!g998) & (g5702)) + ((!g1914) & (g3372) & (!g1949) & (g998) & (g5702)) + ((!g1914) & (g3372) & (g1949) & (!g998) & (g5702)) + ((!g1914) & (g3372) & (g1949) & (g998) & (g5702)) + ((g1914) & (!g3372) & (!g1949) & (!g998) & (g5702)) + ((g1914) & (!g3372) & (!g1949) & (g998) & (!g5702)) + ((g1914) & (!g3372) & (g1949) & (!g998) & (!g5702)) + ((g1914) & (!g3372) & (g1949) & (g998) & (g5702)) + ((g1914) & (g3372) & (!g1949) & (!g998) & (g5702)) + ((g1914) & (g3372) & (!g1949) & (g998) & (!g5702)) + ((g1914) & (g3372) & (g1949) & (!g998) & (!g5702)) + ((g1914) & (g3372) & (g1949) & (g998) & (g5702)));
	assign g5704 = (((!g1914) & (!g2535) & (!g3374) & (!g2153) & (g2159) & (g4708)) + ((!g1914) & (!g2535) & (!g3374) & (g2153) & (!g2159) & (g4708)) + ((!g1914) & (!g2535) & (!g3374) & (g2153) & (g2159) & (!g4708)) + ((!g1914) & (!g2535) & (!g3374) & (g2153) & (g2159) & (g4708)) + ((!g1914) & (!g2535) & (g3374) & (!g2153) & (g2159) & (g4708)) + ((!g1914) & (!g2535) & (g3374) & (g2153) & (!g2159) & (g4708)) + ((!g1914) & (!g2535) & (g3374) & (g2153) & (g2159) & (!g4708)) + ((!g1914) & (!g2535) & (g3374) & (g2153) & (g2159) & (g4708)) + ((!g1914) & (g2535) & (!g3374) & (!g2153) & (!g2159) & (!g4708)) + ((!g1914) & (g2535) & (!g3374) & (!g2153) & (!g2159) & (g4708)) + ((!g1914) & (g2535) & (!g3374) & (!g2153) & (g2159) & (!g4708)) + ((!g1914) & (g2535) & (!g3374) & (g2153) & (!g2159) & (!g4708)) + ((!g1914) & (g2535) & (g3374) & (!g2153) & (!g2159) & (!g4708)) + ((!g1914) & (g2535) & (g3374) & (!g2153) & (!g2159) & (g4708)) + ((!g1914) & (g2535) & (g3374) & (!g2153) & (g2159) & (!g4708)) + ((!g1914) & (g2535) & (g3374) & (g2153) & (!g2159) & (!g4708)) + ((g1914) & (!g2535) & (g3374) & (!g2153) & (!g2159) & (!g4708)) + ((g1914) & (!g2535) & (g3374) & (!g2153) & (!g2159) & (g4708)) + ((g1914) & (!g2535) & (g3374) & (!g2153) & (g2159) & (!g4708)) + ((g1914) & (!g2535) & (g3374) & (!g2153) & (g2159) & (g4708)) + ((g1914) & (!g2535) & (g3374) & (g2153) & (!g2159) & (!g4708)) + ((g1914) & (!g2535) & (g3374) & (g2153) & (!g2159) & (g4708)) + ((g1914) & (!g2535) & (g3374) & (g2153) & (g2159) & (!g4708)) + ((g1914) & (!g2535) & (g3374) & (g2153) & (g2159) & (g4708)) + ((g1914) & (g2535) & (!g3374) & (!g2153) & (!g2159) & (!g4708)) + ((g1914) & (g2535) & (!g3374) & (!g2153) & (!g2159) & (g4708)) + ((g1914) & (g2535) & (!g3374) & (!g2153) & (g2159) & (!g4708)) + ((g1914) & (g2535) & (!g3374) & (!g2153) & (g2159) & (g4708)) + ((g1914) & (g2535) & (!g3374) & (g2153) & (!g2159) & (!g4708)) + ((g1914) & (g2535) & (!g3374) & (g2153) & (!g2159) & (g4708)) + ((g1914) & (g2535) & (!g3374) & (g2153) & (g2159) & (!g4708)) + ((g1914) & (g2535) & (!g3374) & (g2153) & (g2159) & (g4708)));
	assign g5705 = (((!g1914) & (!g2793) & (!g2184) & (!g2198) & (g5704)) + ((!g1914) & (!g2793) & (!g2184) & (g2198) & (!g5704)) + ((!g1914) & (!g2793) & (g2184) & (!g2198) & (!g5704)) + ((!g1914) & (!g2793) & (g2184) & (g2198) & (g5704)) + ((!g1914) & (g2793) & (!g2184) & (!g2198) & (g5704)) + ((!g1914) & (g2793) & (!g2184) & (g2198) & (!g5704)) + ((!g1914) & (g2793) & (g2184) & (!g2198) & (!g5704)) + ((!g1914) & (g2793) & (g2184) & (g2198) & (g5704)) + ((g1914) & (!g2793) & (!g2184) & (!g2198) & (!g5704)) + ((g1914) & (!g2793) & (!g2184) & (g2198) & (!g5704)) + ((g1914) & (!g2793) & (g2184) & (!g2198) & (!g5704)) + ((g1914) & (!g2793) & (g2184) & (g2198) & (!g5704)) + ((g1914) & (g2793) & (!g2184) & (!g2198) & (g5704)) + ((g1914) & (g2793) & (!g2184) & (g2198) & (g5704)) + ((g1914) & (g2793) & (g2184) & (!g2198) & (g5704)) + ((g1914) & (g2793) & (g2184) & (g2198) & (g5704)));
	assign g5706 = (((!g1914) & (!g1970) & (!g3366) & (!g2167) & (g2173) & (g3980)) + ((!g1914) & (!g1970) & (!g3366) & (g2167) & (!g2173) & (g3980)) + ((!g1914) & (!g1970) & (!g3366) & (g2167) & (g2173) & (!g3980)) + ((!g1914) & (!g1970) & (!g3366) & (g2167) & (g2173) & (g3980)) + ((!g1914) & (!g1970) & (g3366) & (!g2167) & (g2173) & (g3980)) + ((!g1914) & (!g1970) & (g3366) & (g2167) & (!g2173) & (g3980)) + ((!g1914) & (!g1970) & (g3366) & (g2167) & (g2173) & (!g3980)) + ((!g1914) & (!g1970) & (g3366) & (g2167) & (g2173) & (g3980)) + ((!g1914) & (g1970) & (!g3366) & (!g2167) & (!g2173) & (!g3980)) + ((!g1914) & (g1970) & (!g3366) & (!g2167) & (!g2173) & (g3980)) + ((!g1914) & (g1970) & (!g3366) & (!g2167) & (g2173) & (!g3980)) + ((!g1914) & (g1970) & (!g3366) & (g2167) & (!g2173) & (!g3980)) + ((!g1914) & (g1970) & (g3366) & (!g2167) & (!g2173) & (!g3980)) + ((!g1914) & (g1970) & (g3366) & (!g2167) & (!g2173) & (g3980)) + ((!g1914) & (g1970) & (g3366) & (!g2167) & (g2173) & (!g3980)) + ((!g1914) & (g1970) & (g3366) & (g2167) & (!g2173) & (!g3980)) + ((g1914) & (!g1970) & (g3366) & (!g2167) & (!g2173) & (!g3980)) + ((g1914) & (!g1970) & (g3366) & (!g2167) & (!g2173) & (g3980)) + ((g1914) & (!g1970) & (g3366) & (!g2167) & (g2173) & (!g3980)) + ((g1914) & (!g1970) & (g3366) & (!g2167) & (g2173) & (g3980)) + ((g1914) & (!g1970) & (g3366) & (g2167) & (!g2173) & (!g3980)) + ((g1914) & (!g1970) & (g3366) & (g2167) & (!g2173) & (g3980)) + ((g1914) & (!g1970) & (g3366) & (g2167) & (g2173) & (!g3980)) + ((g1914) & (!g1970) & (g3366) & (g2167) & (g2173) & (g3980)) + ((g1914) & (g1970) & (!g3366) & (!g2167) & (!g2173) & (!g3980)) + ((g1914) & (g1970) & (!g3366) & (!g2167) & (!g2173) & (g3980)) + ((g1914) & (g1970) & (!g3366) & (!g2167) & (g2173) & (!g3980)) + ((g1914) & (g1970) & (!g3366) & (!g2167) & (g2173) & (g3980)) + ((g1914) & (g1970) & (!g3366) & (g2167) & (!g2173) & (!g3980)) + ((g1914) & (g1970) & (!g3366) & (g2167) & (!g2173) & (g3980)) + ((g1914) & (g1970) & (!g3366) & (g2167) & (g2173) & (!g3980)) + ((g1914) & (g1970) & (!g3366) & (g2167) & (g2173) & (g3980)));
	assign g5707 = (((!g1914) & (!g2789) & (!g2192) & (!g2207) & (g5706)) + ((!g1914) & (!g2789) & (!g2192) & (g2207) & (!g5706)) + ((!g1914) & (!g2789) & (g2192) & (!g2207) & (!g5706)) + ((!g1914) & (!g2789) & (g2192) & (g2207) & (g5706)) + ((!g1914) & (g2789) & (!g2192) & (!g2207) & (g5706)) + ((!g1914) & (g2789) & (!g2192) & (g2207) & (!g5706)) + ((!g1914) & (g2789) & (g2192) & (!g2207) & (!g5706)) + ((!g1914) & (g2789) & (g2192) & (g2207) & (g5706)) + ((g1914) & (!g2789) & (!g2192) & (!g2207) & (!g5706)) + ((g1914) & (!g2789) & (!g2192) & (g2207) & (!g5706)) + ((g1914) & (!g2789) & (g2192) & (!g2207) & (!g5706)) + ((g1914) & (!g2789) & (g2192) & (g2207) & (!g5706)) + ((g1914) & (g2789) & (!g2192) & (!g2207) & (g5706)) + ((g1914) & (g2789) & (!g2192) & (g2207) & (g5706)) + ((g1914) & (g2789) & (g2192) & (!g2207) & (g5706)) + ((g1914) & (g2789) & (g2192) & (g2207) & (g5706)));
	assign g5708 = (((!g1914) & (!g2542) & (g3382) & (!g2144) & (!g2156) & (!g4711)) + ((!g1914) & (!g2542) & (g3382) & (!g2144) & (!g2156) & (g4711)) + ((!g1914) & (!g2542) & (g3382) & (!g2144) & (g2156) & (!g4711)) + ((!g1914) & (!g2542) & (g3382) & (!g2144) & (g2156) & (g4711)) + ((!g1914) & (!g2542) & (g3382) & (g2144) & (!g2156) & (!g4711)) + ((!g1914) & (!g2542) & (g3382) & (g2144) & (!g2156) & (g4711)) + ((!g1914) & (!g2542) & (g3382) & (g2144) & (g2156) & (!g4711)) + ((!g1914) & (!g2542) & (g3382) & (g2144) & (g2156) & (g4711)) + ((!g1914) & (g2542) & (!g3382) & (!g2144) & (!g2156) & (!g4711)) + ((!g1914) & (g2542) & (!g3382) & (!g2144) & (!g2156) & (g4711)) + ((!g1914) & (g2542) & (!g3382) & (!g2144) & (g2156) & (!g4711)) + ((!g1914) & (g2542) & (!g3382) & (!g2144) & (g2156) & (g4711)) + ((!g1914) & (g2542) & (!g3382) & (g2144) & (!g2156) & (!g4711)) + ((!g1914) & (g2542) & (!g3382) & (g2144) & (!g2156) & (g4711)) + ((!g1914) & (g2542) & (!g3382) & (g2144) & (g2156) & (!g4711)) + ((!g1914) & (g2542) & (!g3382) & (g2144) & (g2156) & (g4711)) + ((g1914) & (!g2542) & (!g3382) & (!g2144) & (g2156) & (g4711)) + ((g1914) & (!g2542) & (!g3382) & (g2144) & (!g2156) & (g4711)) + ((g1914) & (!g2542) & (!g3382) & (g2144) & (g2156) & (!g4711)) + ((g1914) & (!g2542) & (!g3382) & (g2144) & (g2156) & (g4711)) + ((g1914) & (!g2542) & (g3382) & (!g2144) & (g2156) & (g4711)) + ((g1914) & (!g2542) & (g3382) & (g2144) & (!g2156) & (g4711)) + ((g1914) & (!g2542) & (g3382) & (g2144) & (g2156) & (!g4711)) + ((g1914) & (!g2542) & (g3382) & (g2144) & (g2156) & (g4711)) + ((g1914) & (g2542) & (!g3382) & (!g2144) & (!g2156) & (!g4711)) + ((g1914) & (g2542) & (!g3382) & (!g2144) & (!g2156) & (g4711)) + ((g1914) & (g2542) & (!g3382) & (!g2144) & (g2156) & (!g4711)) + ((g1914) & (g2542) & (!g3382) & (g2144) & (!g2156) & (!g4711)) + ((g1914) & (g2542) & (g3382) & (!g2144) & (!g2156) & (!g4711)) + ((g1914) & (g2542) & (g3382) & (!g2144) & (!g2156) & (g4711)) + ((g1914) & (g2542) & (g3382) & (!g2144) & (g2156) & (!g4711)) + ((g1914) & (g2542) & (g3382) & (g2144) & (!g2156) & (!g4711)));
	assign g5709 = (((!g1914) & (!g2790) & (!g2188) & (!g2190) & (!g5708)) + ((!g1914) & (!g2790) & (!g2188) & (g2190) & (!g5708)) + ((!g1914) & (!g2790) & (g2188) & (!g2190) & (!g5708)) + ((!g1914) & (!g2790) & (g2188) & (g2190) & (!g5708)) + ((!g1914) & (g2790) & (!g2188) & (!g2190) & (g5708)) + ((!g1914) & (g2790) & (!g2188) & (g2190) & (g5708)) + ((!g1914) & (g2790) & (g2188) & (!g2190) & (g5708)) + ((!g1914) & (g2790) & (g2188) & (g2190) & (g5708)) + ((g1914) & (!g2790) & (!g2188) & (!g2190) & (g5708)) + ((g1914) & (!g2790) & (!g2188) & (g2190) & (!g5708)) + ((g1914) & (!g2790) & (g2188) & (!g2190) & (!g5708)) + ((g1914) & (!g2790) & (g2188) & (g2190) & (g5708)) + ((g1914) & (g2790) & (!g2188) & (!g2190) & (g5708)) + ((g1914) & (g2790) & (!g2188) & (g2190) & (!g5708)) + ((g1914) & (g2790) & (g2188) & (!g2190) & (!g5708)) + ((g1914) & (g2790) & (g2188) & (g2190) & (g5708)));
	assign g5710 = (((!g1914) & (!g2657) & (!g2678) & (!g3303) & (!g2683) & (!g3297)) + ((!g1914) & (!g2657) & (!g2678) & (!g3303) & (!g2683) & (g3297)) + ((!g1914) & (!g2657) & (!g2678) & (!g3303) & (g2683) & (!g3297)) + ((!g1914) & (!g2657) & (!g2678) & (!g3303) & (g2683) & (g3297)) + ((!g1914) & (!g2657) & (g2678) & (g3303) & (!g2683) & (!g3297)) + ((!g1914) & (!g2657) & (g2678) & (g3303) & (!g2683) & (g3297)) + ((!g1914) & (!g2657) & (g2678) & (g3303) & (g2683) & (!g3297)) + ((!g1914) & (!g2657) & (g2678) & (g3303) & (g2683) & (g3297)) + ((!g1914) & (g2657) & (!g2678) & (g3303) & (!g2683) & (!g3297)) + ((!g1914) & (g2657) & (!g2678) & (g3303) & (!g2683) & (g3297)) + ((!g1914) & (g2657) & (!g2678) & (g3303) & (g2683) & (!g3297)) + ((!g1914) & (g2657) & (!g2678) & (g3303) & (g2683) & (g3297)) + ((!g1914) & (g2657) & (g2678) & (!g3303) & (!g2683) & (!g3297)) + ((!g1914) & (g2657) & (g2678) & (!g3303) & (!g2683) & (g3297)) + ((!g1914) & (g2657) & (g2678) & (!g3303) & (g2683) & (!g3297)) + ((!g1914) & (g2657) & (g2678) & (!g3303) & (g2683) & (g3297)) + ((g1914) & (!g2657) & (!g2678) & (!g3303) & (!g2683) & (!g3297)) + ((g1914) & (!g2657) & (!g2678) & (!g3303) & (g2683) & (g3297)) + ((g1914) & (!g2657) & (!g2678) & (g3303) & (!g2683) & (!g3297)) + ((g1914) & (!g2657) & (!g2678) & (g3303) & (g2683) & (g3297)) + ((g1914) & (!g2657) & (g2678) & (!g3303) & (!g2683) & (!g3297)) + ((g1914) & (!g2657) & (g2678) & (!g3303) & (g2683) & (g3297)) + ((g1914) & (!g2657) & (g2678) & (g3303) & (!g2683) & (!g3297)) + ((g1914) & (!g2657) & (g2678) & (g3303) & (g2683) & (g3297)) + ((g1914) & (g2657) & (!g2678) & (!g3303) & (!g2683) & (g3297)) + ((g1914) & (g2657) & (!g2678) & (!g3303) & (g2683) & (!g3297)) + ((g1914) & (g2657) & (!g2678) & (g3303) & (!g2683) & (g3297)) + ((g1914) & (g2657) & (!g2678) & (g3303) & (g2683) & (!g3297)) + ((g1914) & (g2657) & (g2678) & (!g3303) & (!g2683) & (g3297)) + ((g1914) & (g2657) & (g2678) & (!g3303) & (g2683) & (!g3297)) + ((g1914) & (g2657) & (g2678) & (g3303) & (!g2683) & (g3297)) + ((g1914) & (g2657) & (g2678) & (g3303) & (g2683) & (!g3297)));
	assign g5711 = (((!g3255) & (!g5710) & (!g2649) & (!g4841)) + ((!g3255) & (!g5710) & (!g2649) & (g4841)) + ((!g3255) & (!g5710) & (g2649) & (!g4841)) + ((!g3255) & (g5710) & (g2649) & (g4841)) + ((g3255) & (!g5710) & (!g2649) & (!g4841)) + ((g3255) & (g5710) & (!g2649) & (g4841)) + ((g3255) & (g5710) & (g2649) & (!g4841)) + ((g3255) & (g5710) & (g2649) & (g4841)));
	assign g5712 = (((!g1914) & (!g2667) & (!g3291) & (!g3312) & (!g3301) & (!g3307)) + ((!g1914) & (!g2667) & (!g3291) & (!g3312) & (!g3301) & (g3307)) + ((!g1914) & (!g2667) & (!g3291) & (!g3312) & (g3301) & (!g3307)) + ((!g1914) & (!g2667) & (!g3291) & (!g3312) & (g3301) & (g3307)) + ((!g1914) & (!g2667) & (g3291) & (g3312) & (!g3301) & (!g3307)) + ((!g1914) & (!g2667) & (g3291) & (g3312) & (!g3301) & (g3307)) + ((!g1914) & (!g2667) & (g3291) & (g3312) & (g3301) & (!g3307)) + ((!g1914) & (!g2667) & (g3291) & (g3312) & (g3301) & (g3307)) + ((!g1914) & (g2667) & (!g3291) & (g3312) & (!g3301) & (!g3307)) + ((!g1914) & (g2667) & (!g3291) & (g3312) & (!g3301) & (g3307)) + ((!g1914) & (g2667) & (!g3291) & (g3312) & (g3301) & (!g3307)) + ((!g1914) & (g2667) & (!g3291) & (g3312) & (g3301) & (g3307)) + ((!g1914) & (g2667) & (g3291) & (!g3312) & (!g3301) & (!g3307)) + ((!g1914) & (g2667) & (g3291) & (!g3312) & (!g3301) & (g3307)) + ((!g1914) & (g2667) & (g3291) & (!g3312) & (g3301) & (!g3307)) + ((!g1914) & (g2667) & (g3291) & (!g3312) & (g3301) & (g3307)) + ((g1914) & (!g2667) & (!g3291) & (!g3312) & (!g3301) & (!g3307)) + ((g1914) & (!g2667) & (!g3291) & (!g3312) & (g3301) & (g3307)) + ((g1914) & (!g2667) & (!g3291) & (g3312) & (!g3301) & (!g3307)) + ((g1914) & (!g2667) & (!g3291) & (g3312) & (g3301) & (g3307)) + ((g1914) & (!g2667) & (g3291) & (!g3312) & (!g3301) & (!g3307)) + ((g1914) & (!g2667) & (g3291) & (!g3312) & (g3301) & (g3307)) + ((g1914) & (!g2667) & (g3291) & (g3312) & (!g3301) & (!g3307)) + ((g1914) & (!g2667) & (g3291) & (g3312) & (g3301) & (g3307)) + ((g1914) & (g2667) & (!g3291) & (!g3312) & (!g3301) & (g3307)) + ((g1914) & (g2667) & (!g3291) & (!g3312) & (g3301) & (!g3307)) + ((g1914) & (g2667) & (!g3291) & (g3312) & (!g3301) & (g3307)) + ((g1914) & (g2667) & (!g3291) & (g3312) & (g3301) & (!g3307)) + ((g1914) & (g2667) & (g3291) & (!g3312) & (!g3301) & (g3307)) + ((g1914) & (g2667) & (g3291) & (!g3312) & (g3301) & (!g3307)) + ((g1914) & (g2667) & (g3291) & (g3312) & (!g3301) & (g3307)) + ((g1914) & (g2667) & (g3291) & (g3312) & (g3301) & (!g3307)));
	assign g5713 = (((!g3279) & (!g5712) & (!g3222) & (!g4852)) + ((!g3279) & (!g5712) & (!g3222) & (g4852)) + ((!g3279) & (!g5712) & (g3222) & (!g4852)) + ((!g3279) & (g5712) & (g3222) & (g4852)) + ((g3279) & (!g5712) & (!g3222) & (!g4852)) + ((g3279) & (g5712) & (!g3222) & (g4852)) + ((g3279) & (g5712) & (g3222) & (!g4852)) + ((g3279) & (g5712) & (g3222) & (g4852)));
	assign g5714 = (((!g1914) & (!g2676) & (!g3299) & (!g3307) & (!g3310) & (!g3312)) + ((!g1914) & (!g2676) & (!g3299) & (!g3307) & (!g3310) & (g3312)) + ((!g1914) & (!g2676) & (!g3299) & (!g3307) & (g3310) & (!g3312)) + ((!g1914) & (!g2676) & (!g3299) & (!g3307) & (g3310) & (g3312)) + ((!g1914) & (!g2676) & (g3299) & (g3307) & (!g3310) & (!g3312)) + ((!g1914) & (!g2676) & (g3299) & (g3307) & (!g3310) & (g3312)) + ((!g1914) & (!g2676) & (g3299) & (g3307) & (g3310) & (!g3312)) + ((!g1914) & (!g2676) & (g3299) & (g3307) & (g3310) & (g3312)) + ((!g1914) & (g2676) & (!g3299) & (g3307) & (!g3310) & (!g3312)) + ((!g1914) & (g2676) & (!g3299) & (g3307) & (!g3310) & (g3312)) + ((!g1914) & (g2676) & (!g3299) & (g3307) & (g3310) & (!g3312)) + ((!g1914) & (g2676) & (!g3299) & (g3307) & (g3310) & (g3312)) + ((!g1914) & (g2676) & (g3299) & (!g3307) & (!g3310) & (!g3312)) + ((!g1914) & (g2676) & (g3299) & (!g3307) & (!g3310) & (g3312)) + ((!g1914) & (g2676) & (g3299) & (!g3307) & (g3310) & (!g3312)) + ((!g1914) & (g2676) & (g3299) & (!g3307) & (g3310) & (g3312)) + ((g1914) & (!g2676) & (!g3299) & (!g3307) & (!g3310) & (!g3312)) + ((g1914) & (!g2676) & (!g3299) & (!g3307) & (g3310) & (g3312)) + ((g1914) & (!g2676) & (!g3299) & (g3307) & (!g3310) & (!g3312)) + ((g1914) & (!g2676) & (!g3299) & (g3307) & (g3310) & (g3312)) + ((g1914) & (!g2676) & (g3299) & (!g3307) & (!g3310) & (!g3312)) + ((g1914) & (!g2676) & (g3299) & (!g3307) & (g3310) & (g3312)) + ((g1914) & (!g2676) & (g3299) & (g3307) & (!g3310) & (!g3312)) + ((g1914) & (!g2676) & (g3299) & (g3307) & (g3310) & (g3312)) + ((g1914) & (g2676) & (!g3299) & (!g3307) & (!g3310) & (g3312)) + ((g1914) & (g2676) & (!g3299) & (!g3307) & (g3310) & (!g3312)) + ((g1914) & (g2676) & (!g3299) & (g3307) & (!g3310) & (g3312)) + ((g1914) & (g2676) & (!g3299) & (g3307) & (g3310) & (!g3312)) + ((g1914) & (g2676) & (g3299) & (!g3307) & (!g3310) & (g3312)) + ((g1914) & (g2676) & (g3299) & (!g3307) & (g3310) & (!g3312)) + ((g1914) & (g2676) & (g3299) & (g3307) & (!g3310) & (g3312)) + ((g1914) & (g2676) & (g3299) & (g3307) & (g3310) & (!g3312)));
	assign g5715 = (((!g3265) & (!g5714) & (!g3245) & (!g4862)) + ((!g3265) & (!g5714) & (!g3245) & (g4862)) + ((!g3265) & (!g5714) & (g3245) & (!g4862)) + ((!g3265) & (g5714) & (g3245) & (g4862)) + ((g3265) & (!g5714) & (!g3245) & (!g4862)) + ((g3265) & (g5714) & (!g3245) & (g4862)) + ((g3265) & (g5714) & (g3245) & (!g4862)) + ((g3265) & (g5714) & (g3245) & (g4862)));
	assign g5716 = (((g4053) & (g4060)));
	assign g5717 = (((!g2760) & (!g3342)) + ((g2760) & (g3342)));
	assign g5718 = (((!g3323) & (!g3356)) + ((g3323) & (g3356)));
	assign g5719 = (((!g3336) & (!g3348)) + ((g3336) & (g3348)));
	assign g5720 = (((!g363) & (!g386) & (g1269) & (g1303) & (!g409) & (g1337)) + ((!g363) & (!g386) & (g1269) & (g1303) & (g409) & (!g1337)) + ((!g363) & (g386) & (!g1269) & (g1303) & (!g409) & (g1337)) + ((!g363) & (g386) & (!g1269) & (g1303) & (g409) & (!g1337)) + ((!g363) & (g386) & (g1269) & (!g1303) & (!g409) & (g1337)) + ((!g363) & (g386) & (g1269) & (!g1303) & (g409) & (!g1337)) + ((!g363) & (g386) & (g1269) & (g1303) & (!g409) & (g1337)) + ((!g363) & (g386) & (g1269) & (g1303) & (g409) & (!g1337)) + ((g363) & (!g386) & (!g1269) & (g1303) & (!g409) & (g1337)) + ((g363) & (!g386) & (!g1269) & (g1303) & (g409) & (!g1337)) + ((g363) & (!g386) & (g1269) & (g1303) & (!g409) & (g1337)) + ((g363) & (!g386) & (g1269) & (g1303) & (g409) & (!g1337)) + ((g363) & (g386) & (!g1269) & (!g1303) & (!g409) & (g1337)) + ((g363) & (g386) & (!g1269) & (!g1303) & (g409) & (!g1337)) + ((g363) & (g386) & (!g1269) & (g1303) & (!g409) & (g1337)) + ((g363) & (g386) & (!g1269) & (g1303) & (g409) & (!g1337)) + ((g363) & (g386) & (g1269) & (!g1303) & (!g409) & (g1337)) + ((g363) & (g386) & (g1269) & (!g1303) & (g409) & (!g1337)) + ((g363) & (g386) & (g1269) & (g1303) & (!g409) & (g1337)) + ((g363) & (g386) & (g1269) & (g1303) & (g409) & (!g1337)));
	assign g5721 = (((!g363) & (!g386) & (!g1269) & (!g1303) & (!g340) & (!g1236)) + ((!g363) & (!g386) & (!g1269) & (!g1303) & (!g340) & (g1236)) + ((!g363) & (!g386) & (!g1269) & (!g1303) & (g340) & (!g1236)) + ((!g363) & (!g386) & (!g1269) & (g1303) & (!g340) & (!g1236)) + ((!g363) & (!g386) & (!g1269) & (g1303) & (!g340) & (g1236)) + ((!g363) & (!g386) & (!g1269) & (g1303) & (g340) & (!g1236)) + ((!g363) & (!g386) & (g1269) & (!g1303) & (!g340) & (!g1236)) + ((!g363) & (!g386) & (g1269) & (!g1303) & (!g340) & (g1236)) + ((!g363) & (!g386) & (g1269) & (!g1303) & (g340) & (!g1236)) + ((!g363) & (!g386) & (g1269) & (g1303) & (!g340) & (!g1236)) + ((!g363) & (!g386) & (g1269) & (g1303) & (!g340) & (g1236)) + ((!g363) & (!g386) & (g1269) & (g1303) & (g340) & (!g1236)) + ((!g363) & (g386) & (!g1269) & (!g1303) & (!g340) & (!g1236)) + ((!g363) & (g386) & (!g1269) & (!g1303) & (!g340) & (g1236)) + ((!g363) & (g386) & (!g1269) & (!g1303) & (g340) & (!g1236)) + ((!g363) & (g386) & (g1269) & (!g1303) & (!g340) & (!g1236)) + ((!g363) & (g386) & (g1269) & (!g1303) & (!g340) & (g1236)) + ((!g363) & (g386) & (g1269) & (!g1303) & (g340) & (!g1236)) + ((g363) & (!g386) & (!g1269) & (!g1303) & (!g340) & (!g1236)) + ((g363) & (!g386) & (!g1269) & (!g1303) & (!g340) & (g1236)) + ((g363) & (!g386) & (!g1269) & (!g1303) & (g340) & (!g1236)) + ((g363) & (!g386) & (!g1269) & (g1303) & (!g340) & (!g1236)) + ((g363) & (!g386) & (!g1269) & (g1303) & (!g340) & (g1236)) + ((g363) & (!g386) & (!g1269) & (g1303) & (g340) & (!g1236)) + ((g363) & (g386) & (!g1269) & (!g1303) & (!g340) & (!g1236)) + ((g363) & (g386) & (!g1269) & (!g1303) & (!g340) & (g1236)) + ((g363) & (g386) & (!g1269) & (!g1303) & (g340) & (!g1236)));
	assign g5722 = (((!g340) & (!g1236) & (g5720) & (!g5721)) + ((!g340) & (g1236) & (g5720) & (!g5721)) + ((!g340) & (g1236) & (g5720) & (g5721)) + ((g340) & (!g1236) & (g5720) & (!g5721)) + ((g340) & (!g1236) & (g5720) & (g5721)) + ((g340) & (g1236) & (g5720) & (!g5721)) + ((g340) & (g1236) & (g5720) & (g5721)));
	assign g5723 = (((!g2426) & (!g2427) & (!g2518) & (!g2519) & (!g2378) & (!g2379)) + ((!g2426) & (!g2427) & (!g2518) & (!g2519) & (!g2378) & (g2379)) + ((!g2426) & (!g2427) & (!g2518) & (!g2519) & (g2378) & (!g2379)) + ((!g2426) & (!g2427) & (!g2518) & (!g2519) & (g2378) & (g2379)) + ((!g2426) & (!g2427) & (!g2518) & (g2519) & (!g2378) & (!g2379)) + ((!g2426) & (!g2427) & (!g2518) & (g2519) & (!g2378) & (g2379)) + ((!g2426) & (!g2427) & (!g2518) & (g2519) & (g2378) & (!g2379)) + ((!g2426) & (!g2427) & (!g2518) & (g2519) & (g2378) & (g2379)) + ((!g2426) & (!g2427) & (g2518) & (!g2519) & (!g2378) & (!g2379)) + ((!g2426) & (!g2427) & (g2518) & (!g2519) & (!g2378) & (g2379)) + ((!g2426) & (!g2427) & (g2518) & (!g2519) & (g2378) & (!g2379)) + ((!g2426) & (!g2427) & (g2518) & (!g2519) & (g2378) & (g2379)) + ((!g2426) & (g2427) & (!g2518) & (!g2519) & (!g2378) & (!g2379)) + ((!g2426) & (g2427) & (!g2518) & (!g2519) & (!g2378) & (g2379)) + ((!g2426) & (g2427) & (!g2518) & (!g2519) & (g2378) & (!g2379)) + ((!g2426) & (g2427) & (!g2518) & (!g2519) & (g2378) & (g2379)) + ((!g2426) & (g2427) & (!g2518) & (g2519) & (!g2378) & (!g2379)) + ((!g2426) & (g2427) & (g2518) & (!g2519) & (!g2378) & (!g2379)) + ((g2426) & (!g2427) & (!g2518) & (!g2519) & (!g2378) & (!g2379)) + ((g2426) & (!g2427) & (!g2518) & (!g2519) & (!g2378) & (g2379)) + ((g2426) & (!g2427) & (!g2518) & (!g2519) & (g2378) & (!g2379)) + ((g2426) & (!g2427) & (!g2518) & (!g2519) & (g2378) & (g2379)) + ((g2426) & (!g2427) & (!g2518) & (g2519) & (!g2378) & (!g2379)) + ((g2426) & (!g2427) & (g2518) & (!g2519) & (!g2378) & (!g2379)) + ((g2426) & (g2427) & (!g2518) & (!g2519) & (!g2378) & (!g2379)) + ((g2426) & (g2427) & (!g2518) & (!g2519) & (!g2378) & (g2379)) + ((g2426) & (g2427) & (!g2518) & (!g2519) & (g2378) & (!g2379)) + ((g2426) & (g2427) & (!g2518) & (!g2519) & (g2378) & (g2379)));
	assign g5724 = (((!g2426) & (!g2427) & (!g2518) & (!g2519) & (!g2378) & (!g2379)) + ((!g2426) & (!g2427) & (!g2518) & (!g2519) & (!g2378) & (g2379)) + ((!g2426) & (!g2427) & (!g2518) & (!g2519) & (g2378) & (!g2379)) + ((!g2426) & (!g2427) & (!g2518) & (g2519) & (!g2378) & (!g2379)) + ((!g2426) & (!g2427) & (!g2518) & (g2519) & (!g2378) & (g2379)) + ((!g2426) & (!g2427) & (!g2518) & (g2519) & (g2378) & (!g2379)) + ((!g2426) & (!g2427) & (g2518) & (!g2519) & (!g2378) & (!g2379)) + ((!g2426) & (!g2427) & (g2518) & (!g2519) & (!g2378) & (g2379)) + ((!g2426) & (!g2427) & (g2518) & (!g2519) & (g2378) & (!g2379)) + ((!g2426) & (g2427) & (!g2518) & (!g2519) & (!g2378) & (!g2379)) + ((!g2426) & (g2427) & (!g2518) & (!g2519) & (!g2378) & (g2379)) + ((!g2426) & (g2427) & (!g2518) & (!g2519) & (g2378) & (!g2379)) + ((!g2426) & (g2427) & (!g2518) & (g2519) & (!g2378) & (!g2379)) + ((!g2426) & (g2427) & (!g2518) & (g2519) & (!g2378) & (g2379)) + ((!g2426) & (g2427) & (!g2518) & (g2519) & (g2378) & (!g2379)) + ((!g2426) & (g2427) & (g2518) & (!g2519) & (!g2378) & (!g2379)) + ((!g2426) & (g2427) & (g2518) & (!g2519) & (!g2378) & (g2379)) + ((!g2426) & (g2427) & (g2518) & (!g2519) & (g2378) & (!g2379)) + ((g2426) & (!g2427) & (!g2518) & (!g2519) & (!g2378) & (!g2379)) + ((g2426) & (!g2427) & (!g2518) & (!g2519) & (!g2378) & (g2379)) + ((g2426) & (!g2427) & (!g2518) & (!g2519) & (g2378) & (!g2379)) + ((g2426) & (!g2427) & (!g2518) & (g2519) & (!g2378) & (!g2379)) + ((g2426) & (!g2427) & (!g2518) & (g2519) & (!g2378) & (g2379)) + ((g2426) & (!g2427) & (!g2518) & (g2519) & (g2378) & (!g2379)) + ((g2426) & (!g2427) & (g2518) & (!g2519) & (!g2378) & (!g2379)) + ((g2426) & (!g2427) & (g2518) & (!g2519) & (!g2378) & (g2379)) + ((g2426) & (!g2427) & (g2518) & (!g2519) & (g2378) & (!g2379)));
	assign g5725 = (((!g1239) & (!g1279) & (g1972) & (g1975) & (!g1307) & (g2047)) + ((!g1239) & (!g1279) & (g1972) & (g1975) & (g1307) & (!g2047)) + ((!g1239) & (g1279) & (!g1972) & (g1975) & (!g1307) & (g2047)) + ((!g1239) & (g1279) & (!g1972) & (g1975) & (g1307) & (!g2047)) + ((!g1239) & (g1279) & (g1972) & (!g1975) & (!g1307) & (g2047)) + ((!g1239) & (g1279) & (g1972) & (!g1975) & (g1307) & (!g2047)) + ((!g1239) & (g1279) & (g1972) & (g1975) & (!g1307) & (g2047)) + ((!g1239) & (g1279) & (g1972) & (g1975) & (g1307) & (!g2047)) + ((g1239) & (!g1279) & (!g1972) & (g1975) & (!g1307) & (g2047)) + ((g1239) & (!g1279) & (!g1972) & (g1975) & (g1307) & (!g2047)) + ((g1239) & (!g1279) & (g1972) & (g1975) & (!g1307) & (g2047)) + ((g1239) & (!g1279) & (g1972) & (g1975) & (g1307) & (!g2047)) + ((g1239) & (g1279) & (!g1972) & (!g1975) & (!g1307) & (g2047)) + ((g1239) & (g1279) & (!g1972) & (!g1975) & (g1307) & (!g2047)) + ((g1239) & (g1279) & (!g1972) & (g1975) & (!g1307) & (g2047)) + ((g1239) & (g1279) & (!g1972) & (g1975) & (g1307) & (!g2047)) + ((g1239) & (g1279) & (g1972) & (!g1975) & (!g1307) & (g2047)) + ((g1239) & (g1279) & (g1972) & (!g1975) & (g1307) & (!g2047)) + ((g1239) & (g1279) & (g1972) & (g1975) & (!g1307) & (g2047)) + ((g1239) & (g1279) & (g1972) & (g1975) & (g1307) & (!g2047)));
	assign g5726 = (((!g1239) & (!g1279) & (!g1972) & (!g1975) & (!g1212) & (!g1969)) + ((!g1239) & (!g1279) & (!g1972) & (!g1975) & (!g1212) & (g1969)) + ((!g1239) & (!g1279) & (!g1972) & (!g1975) & (g1212) & (!g1969)) + ((!g1239) & (!g1279) & (!g1972) & (g1975) & (!g1212) & (!g1969)) + ((!g1239) & (!g1279) & (!g1972) & (g1975) & (!g1212) & (g1969)) + ((!g1239) & (!g1279) & (!g1972) & (g1975) & (g1212) & (!g1969)) + ((!g1239) & (!g1279) & (g1972) & (!g1975) & (!g1212) & (!g1969)) + ((!g1239) & (!g1279) & (g1972) & (!g1975) & (!g1212) & (g1969)) + ((!g1239) & (!g1279) & (g1972) & (!g1975) & (g1212) & (!g1969)) + ((!g1239) & (!g1279) & (g1972) & (g1975) & (!g1212) & (!g1969)) + ((!g1239) & (!g1279) & (g1972) & (g1975) & (!g1212) & (g1969)) + ((!g1239) & (!g1279) & (g1972) & (g1975) & (g1212) & (!g1969)) + ((!g1239) & (g1279) & (!g1972) & (!g1975) & (!g1212) & (!g1969)) + ((!g1239) & (g1279) & (!g1972) & (!g1975) & (!g1212) & (g1969)) + ((!g1239) & (g1279) & (!g1972) & (!g1975) & (g1212) & (!g1969)) + ((!g1239) & (g1279) & (g1972) & (!g1975) & (!g1212) & (!g1969)) + ((!g1239) & (g1279) & (g1972) & (!g1975) & (!g1212) & (g1969)) + ((!g1239) & (g1279) & (g1972) & (!g1975) & (g1212) & (!g1969)) + ((g1239) & (!g1279) & (!g1972) & (!g1975) & (!g1212) & (!g1969)) + ((g1239) & (!g1279) & (!g1972) & (!g1975) & (!g1212) & (g1969)) + ((g1239) & (!g1279) & (!g1972) & (!g1975) & (g1212) & (!g1969)) + ((g1239) & (!g1279) & (!g1972) & (g1975) & (!g1212) & (!g1969)) + ((g1239) & (!g1279) & (!g1972) & (g1975) & (!g1212) & (g1969)) + ((g1239) & (!g1279) & (!g1972) & (g1975) & (g1212) & (!g1969)) + ((g1239) & (g1279) & (!g1972) & (!g1975) & (!g1212) & (!g1969)) + ((g1239) & (g1279) & (!g1972) & (!g1975) & (!g1212) & (g1969)) + ((g1239) & (g1279) & (!g1972) & (!g1975) & (g1212) & (!g1969)));
	assign g5727 = (((!g1212) & (!g1969) & (g5725) & (!g5726)) + ((!g1212) & (g1969) & (g5725) & (!g5726)) + ((!g1212) & (g1969) & (g5725) & (g5726)) + ((g1212) & (!g1969) & (g5725) & (!g5726)) + ((g1212) & (!g1969) & (g5725) & (g5726)) + ((g1212) & (g1969) & (g5725) & (!g5726)) + ((g1212) & (g1969) & (g5725) & (g5726)));
	assign g5728 = (((!g1241) & (!g1287) & (g2559) & (g2623) & (!g1309) & (g2653)) + ((!g1241) & (!g1287) & (g2559) & (g2623) & (g1309) & (!g2653)) + ((!g1241) & (g1287) & (!g2559) & (g2623) & (!g1309) & (g2653)) + ((!g1241) & (g1287) & (!g2559) & (g2623) & (g1309) & (!g2653)) + ((!g1241) & (g1287) & (g2559) & (!g2623) & (!g1309) & (g2653)) + ((!g1241) & (g1287) & (g2559) & (!g2623) & (g1309) & (!g2653)) + ((!g1241) & (g1287) & (g2559) & (g2623) & (!g1309) & (g2653)) + ((!g1241) & (g1287) & (g2559) & (g2623) & (g1309) & (!g2653)) + ((g1241) & (!g1287) & (!g2559) & (g2623) & (!g1309) & (g2653)) + ((g1241) & (!g1287) & (!g2559) & (g2623) & (g1309) & (!g2653)) + ((g1241) & (!g1287) & (g2559) & (g2623) & (!g1309) & (g2653)) + ((g1241) & (!g1287) & (g2559) & (g2623) & (g1309) & (!g2653)) + ((g1241) & (g1287) & (!g2559) & (!g2623) & (!g1309) & (g2653)) + ((g1241) & (g1287) & (!g2559) & (!g2623) & (g1309) & (!g2653)) + ((g1241) & (g1287) & (!g2559) & (g2623) & (!g1309) & (g2653)) + ((g1241) & (g1287) & (!g2559) & (g2623) & (g1309) & (!g2653)) + ((g1241) & (g1287) & (g2559) & (!g2623) & (!g1309) & (g2653)) + ((g1241) & (g1287) & (g2559) & (!g2623) & (g1309) & (!g2653)) + ((g1241) & (g1287) & (g2559) & (g2623) & (!g1309) & (g2653)) + ((g1241) & (g1287) & (g2559) & (g2623) & (g1309) & (!g2653)));
	assign g5729 = (((!g1241) & (!g1287) & (!g2559) & (!g2623) & (!g1220) & (!g2533)) + ((!g1241) & (!g1287) & (!g2559) & (!g2623) & (!g1220) & (g2533)) + ((!g1241) & (!g1287) & (!g2559) & (!g2623) & (g1220) & (!g2533)) + ((!g1241) & (!g1287) & (!g2559) & (g2623) & (!g1220) & (!g2533)) + ((!g1241) & (!g1287) & (!g2559) & (g2623) & (!g1220) & (g2533)) + ((!g1241) & (!g1287) & (!g2559) & (g2623) & (g1220) & (!g2533)) + ((!g1241) & (!g1287) & (g2559) & (!g2623) & (!g1220) & (!g2533)) + ((!g1241) & (!g1287) & (g2559) & (!g2623) & (!g1220) & (g2533)) + ((!g1241) & (!g1287) & (g2559) & (!g2623) & (g1220) & (!g2533)) + ((!g1241) & (!g1287) & (g2559) & (g2623) & (!g1220) & (!g2533)) + ((!g1241) & (!g1287) & (g2559) & (g2623) & (!g1220) & (g2533)) + ((!g1241) & (!g1287) & (g2559) & (g2623) & (g1220) & (!g2533)) + ((!g1241) & (g1287) & (!g2559) & (!g2623) & (!g1220) & (!g2533)) + ((!g1241) & (g1287) & (!g2559) & (!g2623) & (!g1220) & (g2533)) + ((!g1241) & (g1287) & (!g2559) & (!g2623) & (g1220) & (!g2533)) + ((!g1241) & (g1287) & (g2559) & (!g2623) & (!g1220) & (!g2533)) + ((!g1241) & (g1287) & (g2559) & (!g2623) & (!g1220) & (g2533)) + ((!g1241) & (g1287) & (g2559) & (!g2623) & (g1220) & (!g2533)) + ((g1241) & (!g1287) & (!g2559) & (!g2623) & (!g1220) & (!g2533)) + ((g1241) & (!g1287) & (!g2559) & (!g2623) & (!g1220) & (g2533)) + ((g1241) & (!g1287) & (!g2559) & (!g2623) & (g1220) & (!g2533)) + ((g1241) & (!g1287) & (!g2559) & (g2623) & (!g1220) & (!g2533)) + ((g1241) & (!g1287) & (!g2559) & (g2623) & (!g1220) & (g2533)) + ((g1241) & (!g1287) & (!g2559) & (g2623) & (g1220) & (!g2533)) + ((g1241) & (g1287) & (!g2559) & (!g2623) & (!g1220) & (!g2533)) + ((g1241) & (g1287) & (!g2559) & (!g2623) & (!g1220) & (g2533)) + ((g1241) & (g1287) & (!g2559) & (!g2623) & (g1220) & (!g2533)));
	assign g5730 = (((!g1220) & (!g2533) & (g5728) & (!g5729)) + ((!g1220) & (g2533) & (g5728) & (!g5729)) + ((!g1220) & (g2533) & (g5728) & (g5729)) + ((g1220) & (!g2533) & (g5728) & (!g5729)) + ((g1220) & (!g2533) & (g5728) & (g5729)) + ((g1220) & (g2533) & (g5728) & (!g5729)) + ((g1220) & (g2533) & (g5728) & (g5729)));
	assign g5731 = (((!g1243) & (!g1295) & (g1973) & (g1976) & (!g1311) & (g2048)) + ((!g1243) & (!g1295) & (g1973) & (g1976) & (g1311) & (!g2048)) + ((!g1243) & (g1295) & (!g1973) & (g1976) & (!g1311) & (g2048)) + ((!g1243) & (g1295) & (!g1973) & (g1976) & (g1311) & (!g2048)) + ((!g1243) & (g1295) & (g1973) & (!g1976) & (!g1311) & (g2048)) + ((!g1243) & (g1295) & (g1973) & (!g1976) & (g1311) & (!g2048)) + ((!g1243) & (g1295) & (g1973) & (g1976) & (!g1311) & (g2048)) + ((!g1243) & (g1295) & (g1973) & (g1976) & (g1311) & (!g2048)) + ((g1243) & (!g1295) & (!g1973) & (g1976) & (!g1311) & (g2048)) + ((g1243) & (!g1295) & (!g1973) & (g1976) & (g1311) & (!g2048)) + ((g1243) & (!g1295) & (g1973) & (g1976) & (!g1311) & (g2048)) + ((g1243) & (!g1295) & (g1973) & (g1976) & (g1311) & (!g2048)) + ((g1243) & (g1295) & (!g1973) & (!g1976) & (!g1311) & (g2048)) + ((g1243) & (g1295) & (!g1973) & (!g1976) & (g1311) & (!g2048)) + ((g1243) & (g1295) & (!g1973) & (g1976) & (!g1311) & (g2048)) + ((g1243) & (g1295) & (!g1973) & (g1976) & (g1311) & (!g2048)) + ((g1243) & (g1295) & (g1973) & (!g1976) & (!g1311) & (g2048)) + ((g1243) & (g1295) & (g1973) & (!g1976) & (g1311) & (!g2048)) + ((g1243) & (g1295) & (g1973) & (g1976) & (!g1311) & (g2048)) + ((g1243) & (g1295) & (g1973) & (g1976) & (g1311) & (!g2048)));
	assign g5732 = (((!g1243) & (!g1295) & (!g1973) & (!g1976) & (!g1228) & (!g1970)) + ((!g1243) & (!g1295) & (!g1973) & (!g1976) & (!g1228) & (g1970)) + ((!g1243) & (!g1295) & (!g1973) & (!g1976) & (g1228) & (!g1970)) + ((!g1243) & (!g1295) & (!g1973) & (g1976) & (!g1228) & (!g1970)) + ((!g1243) & (!g1295) & (!g1973) & (g1976) & (!g1228) & (g1970)) + ((!g1243) & (!g1295) & (!g1973) & (g1976) & (g1228) & (!g1970)) + ((!g1243) & (!g1295) & (g1973) & (!g1976) & (!g1228) & (!g1970)) + ((!g1243) & (!g1295) & (g1973) & (!g1976) & (!g1228) & (g1970)) + ((!g1243) & (!g1295) & (g1973) & (!g1976) & (g1228) & (!g1970)) + ((!g1243) & (!g1295) & (g1973) & (g1976) & (!g1228) & (!g1970)) + ((!g1243) & (!g1295) & (g1973) & (g1976) & (!g1228) & (g1970)) + ((!g1243) & (!g1295) & (g1973) & (g1976) & (g1228) & (!g1970)) + ((!g1243) & (g1295) & (!g1973) & (!g1976) & (!g1228) & (!g1970)) + ((!g1243) & (g1295) & (!g1973) & (!g1976) & (!g1228) & (g1970)) + ((!g1243) & (g1295) & (!g1973) & (!g1976) & (g1228) & (!g1970)) + ((!g1243) & (g1295) & (g1973) & (!g1976) & (!g1228) & (!g1970)) + ((!g1243) & (g1295) & (g1973) & (!g1976) & (!g1228) & (g1970)) + ((!g1243) & (g1295) & (g1973) & (!g1976) & (g1228) & (!g1970)) + ((g1243) & (!g1295) & (!g1973) & (!g1976) & (!g1228) & (!g1970)) + ((g1243) & (!g1295) & (!g1973) & (!g1976) & (!g1228) & (g1970)) + ((g1243) & (!g1295) & (!g1973) & (!g1976) & (g1228) & (!g1970)) + ((g1243) & (!g1295) & (!g1973) & (g1976) & (!g1228) & (!g1970)) + ((g1243) & (!g1295) & (!g1973) & (g1976) & (!g1228) & (g1970)) + ((g1243) & (!g1295) & (!g1973) & (g1976) & (g1228) & (!g1970)) + ((g1243) & (g1295) & (!g1973) & (!g1976) & (!g1228) & (!g1970)) + ((g1243) & (g1295) & (!g1973) & (!g1976) & (!g1228) & (g1970)) + ((g1243) & (g1295) & (!g1973) & (!g1976) & (g1228) & (!g1970)));
	assign g5733 = (((!g1228) & (!g1970) & (g5731) & (!g5732)) + ((!g1228) & (g1970) & (g5731) & (!g5732)) + ((!g1228) & (g1970) & (g5731) & (g5732)) + ((g1228) & (!g1970) & (g5731) & (!g5732)) + ((g1228) & (!g1970) & (g5731) & (g5732)) + ((g1228) & (g1970) & (g5731) & (!g5732)) + ((g1228) & (g1970) & (g5731) & (g5732)));
	assign g5734 = (((!g1245) & (!g1273) & (g2011) & (g2013) & (!g1313) & (g2051)) + ((!g1245) & (!g1273) & (g2011) & (g2013) & (g1313) & (!g2051)) + ((!g1245) & (g1273) & (!g2011) & (g2013) & (!g1313) & (g2051)) + ((!g1245) & (g1273) & (!g2011) & (g2013) & (g1313) & (!g2051)) + ((!g1245) & (g1273) & (g2011) & (!g2013) & (!g1313) & (g2051)) + ((!g1245) & (g1273) & (g2011) & (!g2013) & (g1313) & (!g2051)) + ((!g1245) & (g1273) & (g2011) & (g2013) & (!g1313) & (g2051)) + ((!g1245) & (g1273) & (g2011) & (g2013) & (g1313) & (!g2051)) + ((g1245) & (!g1273) & (!g2011) & (g2013) & (!g1313) & (g2051)) + ((g1245) & (!g1273) & (!g2011) & (g2013) & (g1313) & (!g2051)) + ((g1245) & (!g1273) & (g2011) & (g2013) & (!g1313) & (g2051)) + ((g1245) & (!g1273) & (g2011) & (g2013) & (g1313) & (!g2051)) + ((g1245) & (g1273) & (!g2011) & (!g2013) & (!g1313) & (g2051)) + ((g1245) & (g1273) & (!g2011) & (!g2013) & (g1313) & (!g2051)) + ((g1245) & (g1273) & (!g2011) & (g2013) & (!g1313) & (g2051)) + ((g1245) & (g1273) & (!g2011) & (g2013) & (g1313) & (!g2051)) + ((g1245) & (g1273) & (g2011) & (!g2013) & (!g1313) & (g2051)) + ((g1245) & (g1273) & (g2011) & (!g2013) & (g1313) & (!g2051)) + ((g1245) & (g1273) & (g2011) & (g2013) & (!g1313) & (g2051)) + ((g1245) & (g1273) & (g2011) & (g2013) & (g1313) & (!g2051)));
	assign g5735 = (((!g1245) & (!g1273) & (!g2011) & (!g2013) & (!g1206) & (!g2005)) + ((!g1245) & (!g1273) & (!g2011) & (!g2013) & (!g1206) & (g2005)) + ((!g1245) & (!g1273) & (!g2011) & (!g2013) & (g1206) & (!g2005)) + ((!g1245) & (!g1273) & (!g2011) & (g2013) & (!g1206) & (!g2005)) + ((!g1245) & (!g1273) & (!g2011) & (g2013) & (!g1206) & (g2005)) + ((!g1245) & (!g1273) & (!g2011) & (g2013) & (g1206) & (!g2005)) + ((!g1245) & (!g1273) & (g2011) & (!g2013) & (!g1206) & (!g2005)) + ((!g1245) & (!g1273) & (g2011) & (!g2013) & (!g1206) & (g2005)) + ((!g1245) & (!g1273) & (g2011) & (!g2013) & (g1206) & (!g2005)) + ((!g1245) & (!g1273) & (g2011) & (g2013) & (!g1206) & (!g2005)) + ((!g1245) & (!g1273) & (g2011) & (g2013) & (!g1206) & (g2005)) + ((!g1245) & (!g1273) & (g2011) & (g2013) & (g1206) & (!g2005)) + ((!g1245) & (g1273) & (!g2011) & (!g2013) & (!g1206) & (!g2005)) + ((!g1245) & (g1273) & (!g2011) & (!g2013) & (!g1206) & (g2005)) + ((!g1245) & (g1273) & (!g2011) & (!g2013) & (g1206) & (!g2005)) + ((!g1245) & (g1273) & (g2011) & (!g2013) & (!g1206) & (!g2005)) + ((!g1245) & (g1273) & (g2011) & (!g2013) & (!g1206) & (g2005)) + ((!g1245) & (g1273) & (g2011) & (!g2013) & (g1206) & (!g2005)) + ((g1245) & (!g1273) & (!g2011) & (!g2013) & (!g1206) & (!g2005)) + ((g1245) & (!g1273) & (!g2011) & (!g2013) & (!g1206) & (g2005)) + ((g1245) & (!g1273) & (!g2011) & (!g2013) & (g1206) & (!g2005)) + ((g1245) & (!g1273) & (!g2011) & (g2013) & (!g1206) & (!g2005)) + ((g1245) & (!g1273) & (!g2011) & (g2013) & (!g1206) & (g2005)) + ((g1245) & (!g1273) & (!g2011) & (g2013) & (g1206) & (!g2005)) + ((g1245) & (g1273) & (!g2011) & (!g2013) & (!g1206) & (!g2005)) + ((g1245) & (g1273) & (!g2011) & (!g2013) & (!g1206) & (g2005)) + ((g1245) & (g1273) & (!g2011) & (!g2013) & (g1206) & (!g2005)));
	assign g5736 = (((!g1206) & (!g2005) & (g5734) & (!g5735)) + ((!g1206) & (g2005) & (g5734) & (!g5735)) + ((!g1206) & (g2005) & (g5734) & (g5735)) + ((g1206) & (!g2005) & (g5734) & (!g5735)) + ((g1206) & (!g2005) & (g5734) & (g5735)) + ((g1206) & (g2005) & (g5734) & (!g5735)) + ((g1206) & (g2005) & (g5734) & (g5735)));
	assign g5737 = (((!g1247) & (!g1281) & (g2566) & (g2614) & (!g1315) & (g2657)) + ((!g1247) & (!g1281) & (g2566) & (g2614) & (g1315) & (!g2657)) + ((!g1247) & (g1281) & (!g2566) & (g2614) & (!g1315) & (g2657)) + ((!g1247) & (g1281) & (!g2566) & (g2614) & (g1315) & (!g2657)) + ((!g1247) & (g1281) & (g2566) & (!g2614) & (!g1315) & (g2657)) + ((!g1247) & (g1281) & (g2566) & (!g2614) & (g1315) & (!g2657)) + ((!g1247) & (g1281) & (g2566) & (g2614) & (!g1315) & (g2657)) + ((!g1247) & (g1281) & (g2566) & (g2614) & (g1315) & (!g2657)) + ((g1247) & (!g1281) & (!g2566) & (g2614) & (!g1315) & (g2657)) + ((g1247) & (!g1281) & (!g2566) & (g2614) & (g1315) & (!g2657)) + ((g1247) & (!g1281) & (g2566) & (g2614) & (!g1315) & (g2657)) + ((g1247) & (!g1281) & (g2566) & (g2614) & (g1315) & (!g2657)) + ((g1247) & (g1281) & (!g2566) & (!g2614) & (!g1315) & (g2657)) + ((g1247) & (g1281) & (!g2566) & (!g2614) & (g1315) & (!g2657)) + ((g1247) & (g1281) & (!g2566) & (g2614) & (!g1315) & (g2657)) + ((g1247) & (g1281) & (!g2566) & (g2614) & (g1315) & (!g2657)) + ((g1247) & (g1281) & (g2566) & (!g2614) & (!g1315) & (g2657)) + ((g1247) & (g1281) & (g2566) & (!g2614) & (g1315) & (!g2657)) + ((g1247) & (g1281) & (g2566) & (g2614) & (!g1315) & (g2657)) + ((g1247) & (g1281) & (g2566) & (g2614) & (g1315) & (!g2657)));
	assign g5738 = (((!g1247) & (!g1281) & (!g2566) & (!g2614) & (!g1214) & (!g2527)) + ((!g1247) & (!g1281) & (!g2566) & (!g2614) & (!g1214) & (g2527)) + ((!g1247) & (!g1281) & (!g2566) & (!g2614) & (g1214) & (!g2527)) + ((!g1247) & (!g1281) & (!g2566) & (g2614) & (!g1214) & (!g2527)) + ((!g1247) & (!g1281) & (!g2566) & (g2614) & (!g1214) & (g2527)) + ((!g1247) & (!g1281) & (!g2566) & (g2614) & (g1214) & (!g2527)) + ((!g1247) & (!g1281) & (g2566) & (!g2614) & (!g1214) & (!g2527)) + ((!g1247) & (!g1281) & (g2566) & (!g2614) & (!g1214) & (g2527)) + ((!g1247) & (!g1281) & (g2566) & (!g2614) & (g1214) & (!g2527)) + ((!g1247) & (!g1281) & (g2566) & (g2614) & (!g1214) & (!g2527)) + ((!g1247) & (!g1281) & (g2566) & (g2614) & (!g1214) & (g2527)) + ((!g1247) & (!g1281) & (g2566) & (g2614) & (g1214) & (!g2527)) + ((!g1247) & (g1281) & (!g2566) & (!g2614) & (!g1214) & (!g2527)) + ((!g1247) & (g1281) & (!g2566) & (!g2614) & (!g1214) & (g2527)) + ((!g1247) & (g1281) & (!g2566) & (!g2614) & (g1214) & (!g2527)) + ((!g1247) & (g1281) & (g2566) & (!g2614) & (!g1214) & (!g2527)) + ((!g1247) & (g1281) & (g2566) & (!g2614) & (!g1214) & (g2527)) + ((!g1247) & (g1281) & (g2566) & (!g2614) & (g1214) & (!g2527)) + ((g1247) & (!g1281) & (!g2566) & (!g2614) & (!g1214) & (!g2527)) + ((g1247) & (!g1281) & (!g2566) & (!g2614) & (!g1214) & (g2527)) + ((g1247) & (!g1281) & (!g2566) & (!g2614) & (g1214) & (!g2527)) + ((g1247) & (!g1281) & (!g2566) & (g2614) & (!g1214) & (!g2527)) + ((g1247) & (!g1281) & (!g2566) & (g2614) & (!g1214) & (g2527)) + ((g1247) & (!g1281) & (!g2566) & (g2614) & (g1214) & (!g2527)) + ((g1247) & (g1281) & (!g2566) & (!g2614) & (!g1214) & (!g2527)) + ((g1247) & (g1281) & (!g2566) & (!g2614) & (!g1214) & (g2527)) + ((g1247) & (g1281) & (!g2566) & (!g2614) & (g1214) & (!g2527)));
	assign g5739 = (((!g1214) & (!g2527) & (g5737) & (!g5738)) + ((!g1214) & (g2527) & (g5737) & (!g5738)) + ((!g1214) & (g2527) & (g5737) & (g5738)) + ((g1214) & (!g2527) & (g5737) & (!g5738)) + ((g1214) & (!g2527) & (g5737) & (g5738)) + ((g1214) & (g2527) & (g5737) & (!g5738)) + ((g1214) & (g2527) & (g5737) & (g5738)));
	assign g5740 = (((!g1249) & (!g1289) & (g2569) & (g2626) & (!g1317) & (g2659)) + ((!g1249) & (!g1289) & (g2569) & (g2626) & (g1317) & (!g2659)) + ((!g1249) & (g1289) & (!g2569) & (g2626) & (!g1317) & (g2659)) + ((!g1249) & (g1289) & (!g2569) & (g2626) & (g1317) & (!g2659)) + ((!g1249) & (g1289) & (g2569) & (!g2626) & (!g1317) & (g2659)) + ((!g1249) & (g1289) & (g2569) & (!g2626) & (g1317) & (!g2659)) + ((!g1249) & (g1289) & (g2569) & (g2626) & (!g1317) & (g2659)) + ((!g1249) & (g1289) & (g2569) & (g2626) & (g1317) & (!g2659)) + ((g1249) & (!g1289) & (!g2569) & (g2626) & (!g1317) & (g2659)) + ((g1249) & (!g1289) & (!g2569) & (g2626) & (g1317) & (!g2659)) + ((g1249) & (!g1289) & (g2569) & (g2626) & (!g1317) & (g2659)) + ((g1249) & (!g1289) & (g2569) & (g2626) & (g1317) & (!g2659)) + ((g1249) & (g1289) & (!g2569) & (!g2626) & (!g1317) & (g2659)) + ((g1249) & (g1289) & (!g2569) & (!g2626) & (g1317) & (!g2659)) + ((g1249) & (g1289) & (!g2569) & (g2626) & (!g1317) & (g2659)) + ((g1249) & (g1289) & (!g2569) & (g2626) & (g1317) & (!g2659)) + ((g1249) & (g1289) & (g2569) & (!g2626) & (!g1317) & (g2659)) + ((g1249) & (g1289) & (g2569) & (!g2626) & (g1317) & (!g2659)) + ((g1249) & (g1289) & (g2569) & (g2626) & (!g1317) & (g2659)) + ((g1249) & (g1289) & (g2569) & (g2626) & (g1317) & (!g2659)));
	assign g5741 = (((!g1249) & (!g1289) & (!g2569) & (!g2626) & (!g1222) & (!g2535)) + ((!g1249) & (!g1289) & (!g2569) & (!g2626) & (!g1222) & (g2535)) + ((!g1249) & (!g1289) & (!g2569) & (!g2626) & (g1222) & (!g2535)) + ((!g1249) & (!g1289) & (!g2569) & (g2626) & (!g1222) & (!g2535)) + ((!g1249) & (!g1289) & (!g2569) & (g2626) & (!g1222) & (g2535)) + ((!g1249) & (!g1289) & (!g2569) & (g2626) & (g1222) & (!g2535)) + ((!g1249) & (!g1289) & (g2569) & (!g2626) & (!g1222) & (!g2535)) + ((!g1249) & (!g1289) & (g2569) & (!g2626) & (!g1222) & (g2535)) + ((!g1249) & (!g1289) & (g2569) & (!g2626) & (g1222) & (!g2535)) + ((!g1249) & (!g1289) & (g2569) & (g2626) & (!g1222) & (!g2535)) + ((!g1249) & (!g1289) & (g2569) & (g2626) & (!g1222) & (g2535)) + ((!g1249) & (!g1289) & (g2569) & (g2626) & (g1222) & (!g2535)) + ((!g1249) & (g1289) & (!g2569) & (!g2626) & (!g1222) & (!g2535)) + ((!g1249) & (g1289) & (!g2569) & (!g2626) & (!g1222) & (g2535)) + ((!g1249) & (g1289) & (!g2569) & (!g2626) & (g1222) & (!g2535)) + ((!g1249) & (g1289) & (g2569) & (!g2626) & (!g1222) & (!g2535)) + ((!g1249) & (g1289) & (g2569) & (!g2626) & (!g1222) & (g2535)) + ((!g1249) & (g1289) & (g2569) & (!g2626) & (g1222) & (!g2535)) + ((g1249) & (!g1289) & (!g2569) & (!g2626) & (!g1222) & (!g2535)) + ((g1249) & (!g1289) & (!g2569) & (!g2626) & (!g1222) & (g2535)) + ((g1249) & (!g1289) & (!g2569) & (!g2626) & (g1222) & (!g2535)) + ((g1249) & (!g1289) & (!g2569) & (g2626) & (!g1222) & (!g2535)) + ((g1249) & (!g1289) & (!g2569) & (g2626) & (!g1222) & (g2535)) + ((g1249) & (!g1289) & (!g2569) & (g2626) & (g1222) & (!g2535)) + ((g1249) & (g1289) & (!g2569) & (!g2626) & (!g1222) & (!g2535)) + ((g1249) & (g1289) & (!g2569) & (!g2626) & (!g1222) & (g2535)) + ((g1249) & (g1289) & (!g2569) & (!g2626) & (g1222) & (!g2535)));
	assign g5742 = (((!g1222) & (!g2535) & (g5740) & (!g5741)) + ((!g1222) & (g2535) & (g5740) & (!g5741)) + ((!g1222) & (g2535) & (g5740) & (g5741)) + ((g1222) & (!g2535) & (g5740) & (!g5741)) + ((g1222) & (!g2535) & (g5740) & (g5741)) + ((g1222) & (g2535) & (g5740) & (!g5741)) + ((g1222) & (g2535) & (g5740) & (g5741)));
	assign g5743 = (((!g1251) & (!g1297) & (g2572) & (g2637) & (!g1319) & (g2661)) + ((!g1251) & (!g1297) & (g2572) & (g2637) & (g1319) & (!g2661)) + ((!g1251) & (g1297) & (!g2572) & (g2637) & (!g1319) & (g2661)) + ((!g1251) & (g1297) & (!g2572) & (g2637) & (g1319) & (!g2661)) + ((!g1251) & (g1297) & (g2572) & (!g2637) & (!g1319) & (g2661)) + ((!g1251) & (g1297) & (g2572) & (!g2637) & (g1319) & (!g2661)) + ((!g1251) & (g1297) & (g2572) & (g2637) & (!g1319) & (g2661)) + ((!g1251) & (g1297) & (g2572) & (g2637) & (g1319) & (!g2661)) + ((g1251) & (!g1297) & (!g2572) & (g2637) & (!g1319) & (g2661)) + ((g1251) & (!g1297) & (!g2572) & (g2637) & (g1319) & (!g2661)) + ((g1251) & (!g1297) & (g2572) & (g2637) & (!g1319) & (g2661)) + ((g1251) & (!g1297) & (g2572) & (g2637) & (g1319) & (!g2661)) + ((g1251) & (g1297) & (!g2572) & (!g2637) & (!g1319) & (g2661)) + ((g1251) & (g1297) & (!g2572) & (!g2637) & (g1319) & (!g2661)) + ((g1251) & (g1297) & (!g2572) & (g2637) & (!g1319) & (g2661)) + ((g1251) & (g1297) & (!g2572) & (g2637) & (g1319) & (!g2661)) + ((g1251) & (g1297) & (g2572) & (!g2637) & (!g1319) & (g2661)) + ((g1251) & (g1297) & (g2572) & (!g2637) & (g1319) & (!g2661)) + ((g1251) & (g1297) & (g2572) & (g2637) & (!g1319) & (g2661)) + ((g1251) & (g1297) & (g2572) & (g2637) & (g1319) & (!g2661)));
	assign g5744 = (((!g1251) & (!g1297) & (!g2572) & (!g2637) & (!g1230) & (!g2542)) + ((!g1251) & (!g1297) & (!g2572) & (!g2637) & (!g1230) & (g2542)) + ((!g1251) & (!g1297) & (!g2572) & (!g2637) & (g1230) & (!g2542)) + ((!g1251) & (!g1297) & (!g2572) & (g2637) & (!g1230) & (!g2542)) + ((!g1251) & (!g1297) & (!g2572) & (g2637) & (!g1230) & (g2542)) + ((!g1251) & (!g1297) & (!g2572) & (g2637) & (g1230) & (!g2542)) + ((!g1251) & (!g1297) & (g2572) & (!g2637) & (!g1230) & (!g2542)) + ((!g1251) & (!g1297) & (g2572) & (!g2637) & (!g1230) & (g2542)) + ((!g1251) & (!g1297) & (g2572) & (!g2637) & (g1230) & (!g2542)) + ((!g1251) & (!g1297) & (g2572) & (g2637) & (!g1230) & (!g2542)) + ((!g1251) & (!g1297) & (g2572) & (g2637) & (!g1230) & (g2542)) + ((!g1251) & (!g1297) & (g2572) & (g2637) & (g1230) & (!g2542)) + ((!g1251) & (g1297) & (!g2572) & (!g2637) & (!g1230) & (!g2542)) + ((!g1251) & (g1297) & (!g2572) & (!g2637) & (!g1230) & (g2542)) + ((!g1251) & (g1297) & (!g2572) & (!g2637) & (g1230) & (!g2542)) + ((!g1251) & (g1297) & (g2572) & (!g2637) & (!g1230) & (!g2542)) + ((!g1251) & (g1297) & (g2572) & (!g2637) & (!g1230) & (g2542)) + ((!g1251) & (g1297) & (g2572) & (!g2637) & (g1230) & (!g2542)) + ((g1251) & (!g1297) & (!g2572) & (!g2637) & (!g1230) & (!g2542)) + ((g1251) & (!g1297) & (!g2572) & (!g2637) & (!g1230) & (g2542)) + ((g1251) & (!g1297) & (!g2572) & (!g2637) & (g1230) & (!g2542)) + ((g1251) & (!g1297) & (!g2572) & (g2637) & (!g1230) & (!g2542)) + ((g1251) & (!g1297) & (!g2572) & (g2637) & (!g1230) & (g2542)) + ((g1251) & (!g1297) & (!g2572) & (g2637) & (g1230) & (!g2542)) + ((g1251) & (g1297) & (!g2572) & (!g2637) & (!g1230) & (!g2542)) + ((g1251) & (g1297) & (!g2572) & (!g2637) & (!g1230) & (g2542)) + ((g1251) & (g1297) & (!g2572) & (!g2637) & (g1230) & (!g2542)));
	assign g5745 = (((!g1230) & (!g2542) & (g5743) & (!g5744)) + ((!g1230) & (g2542) & (g5743) & (!g5744)) + ((!g1230) & (g2542) & (g5743) & (g5744)) + ((g1230) & (!g2542) & (g5743) & (!g5744)) + ((g1230) & (!g2542) & (g5743) & (g5744)) + ((g1230) & (g2542) & (g5743) & (!g5744)) + ((g1230) & (g2542) & (g5743) & (g5744)));
	assign g5746 = (((!g1253) & (!g1275) & (g2575) & (g2607) & (!g1321) & (g2663)) + ((!g1253) & (!g1275) & (g2575) & (g2607) & (g1321) & (!g2663)) + ((!g1253) & (g1275) & (!g2575) & (g2607) & (!g1321) & (g2663)) + ((!g1253) & (g1275) & (!g2575) & (g2607) & (g1321) & (!g2663)) + ((!g1253) & (g1275) & (g2575) & (!g2607) & (!g1321) & (g2663)) + ((!g1253) & (g1275) & (g2575) & (!g2607) & (g1321) & (!g2663)) + ((!g1253) & (g1275) & (g2575) & (g2607) & (!g1321) & (g2663)) + ((!g1253) & (g1275) & (g2575) & (g2607) & (g1321) & (!g2663)) + ((g1253) & (!g1275) & (!g2575) & (g2607) & (!g1321) & (g2663)) + ((g1253) & (!g1275) & (!g2575) & (g2607) & (g1321) & (!g2663)) + ((g1253) & (!g1275) & (g2575) & (g2607) & (!g1321) & (g2663)) + ((g1253) & (!g1275) & (g2575) & (g2607) & (g1321) & (!g2663)) + ((g1253) & (g1275) & (!g2575) & (!g2607) & (!g1321) & (g2663)) + ((g1253) & (g1275) & (!g2575) & (!g2607) & (g1321) & (!g2663)) + ((g1253) & (g1275) & (!g2575) & (g2607) & (!g1321) & (g2663)) + ((g1253) & (g1275) & (!g2575) & (g2607) & (g1321) & (!g2663)) + ((g1253) & (g1275) & (g2575) & (!g2607) & (!g1321) & (g2663)) + ((g1253) & (g1275) & (g2575) & (!g2607) & (g1321) & (!g2663)) + ((g1253) & (g1275) & (g2575) & (g2607) & (!g1321) & (g2663)) + ((g1253) & (g1275) & (g2575) & (g2607) & (g1321) & (!g2663)));
	assign g5747 = (((!g1253) & (!g1275) & (!g2575) & (!g2607) & (!g1208) & (!g2523)) + ((!g1253) & (!g1275) & (!g2575) & (!g2607) & (!g1208) & (g2523)) + ((!g1253) & (!g1275) & (!g2575) & (!g2607) & (g1208) & (!g2523)) + ((!g1253) & (!g1275) & (!g2575) & (g2607) & (!g1208) & (!g2523)) + ((!g1253) & (!g1275) & (!g2575) & (g2607) & (!g1208) & (g2523)) + ((!g1253) & (!g1275) & (!g2575) & (g2607) & (g1208) & (!g2523)) + ((!g1253) & (!g1275) & (g2575) & (!g2607) & (!g1208) & (!g2523)) + ((!g1253) & (!g1275) & (g2575) & (!g2607) & (!g1208) & (g2523)) + ((!g1253) & (!g1275) & (g2575) & (!g2607) & (g1208) & (!g2523)) + ((!g1253) & (!g1275) & (g2575) & (g2607) & (!g1208) & (!g2523)) + ((!g1253) & (!g1275) & (g2575) & (g2607) & (!g1208) & (g2523)) + ((!g1253) & (!g1275) & (g2575) & (g2607) & (g1208) & (!g2523)) + ((!g1253) & (g1275) & (!g2575) & (!g2607) & (!g1208) & (!g2523)) + ((!g1253) & (g1275) & (!g2575) & (!g2607) & (!g1208) & (g2523)) + ((!g1253) & (g1275) & (!g2575) & (!g2607) & (g1208) & (!g2523)) + ((!g1253) & (g1275) & (g2575) & (!g2607) & (!g1208) & (!g2523)) + ((!g1253) & (g1275) & (g2575) & (!g2607) & (!g1208) & (g2523)) + ((!g1253) & (g1275) & (g2575) & (!g2607) & (g1208) & (!g2523)) + ((g1253) & (!g1275) & (!g2575) & (!g2607) & (!g1208) & (!g2523)) + ((g1253) & (!g1275) & (!g2575) & (!g2607) & (!g1208) & (g2523)) + ((g1253) & (!g1275) & (!g2575) & (!g2607) & (g1208) & (!g2523)) + ((g1253) & (!g1275) & (!g2575) & (g2607) & (!g1208) & (!g2523)) + ((g1253) & (!g1275) & (!g2575) & (g2607) & (!g1208) & (g2523)) + ((g1253) & (!g1275) & (!g2575) & (g2607) & (g1208) & (!g2523)) + ((g1253) & (g1275) & (!g2575) & (!g2607) & (!g1208) & (!g2523)) + ((g1253) & (g1275) & (!g2575) & (!g2607) & (!g1208) & (g2523)) + ((g1253) & (g1275) & (!g2575) & (!g2607) & (g1208) & (!g2523)));
	assign g5748 = (((!g1208) & (!g2523) & (g5746) & (!g5747)) + ((!g1208) & (g2523) & (g5746) & (!g5747)) + ((!g1208) & (g2523) & (g5746) & (g5747)) + ((g1208) & (!g2523) & (g5746) & (!g5747)) + ((g1208) & (!g2523) & (g5746) & (g5747)) + ((g1208) & (g2523) & (g5746) & (!g5747)) + ((g1208) & (g2523) & (g5746) & (g5747)));
	assign g5749 = (((!g1255) & (!g1283) & (g2578) & (g2617) & (!g1323) & (g2665)) + ((!g1255) & (!g1283) & (g2578) & (g2617) & (g1323) & (!g2665)) + ((!g1255) & (g1283) & (!g2578) & (g2617) & (!g1323) & (g2665)) + ((!g1255) & (g1283) & (!g2578) & (g2617) & (g1323) & (!g2665)) + ((!g1255) & (g1283) & (g2578) & (!g2617) & (!g1323) & (g2665)) + ((!g1255) & (g1283) & (g2578) & (!g2617) & (g1323) & (!g2665)) + ((!g1255) & (g1283) & (g2578) & (g2617) & (!g1323) & (g2665)) + ((!g1255) & (g1283) & (g2578) & (g2617) & (g1323) & (!g2665)) + ((g1255) & (!g1283) & (!g2578) & (g2617) & (!g1323) & (g2665)) + ((g1255) & (!g1283) & (!g2578) & (g2617) & (g1323) & (!g2665)) + ((g1255) & (!g1283) & (g2578) & (g2617) & (!g1323) & (g2665)) + ((g1255) & (!g1283) & (g2578) & (g2617) & (g1323) & (!g2665)) + ((g1255) & (g1283) & (!g2578) & (!g2617) & (!g1323) & (g2665)) + ((g1255) & (g1283) & (!g2578) & (!g2617) & (g1323) & (!g2665)) + ((g1255) & (g1283) & (!g2578) & (g2617) & (!g1323) & (g2665)) + ((g1255) & (g1283) & (!g2578) & (g2617) & (g1323) & (!g2665)) + ((g1255) & (g1283) & (g2578) & (!g2617) & (!g1323) & (g2665)) + ((g1255) & (g1283) & (g2578) & (!g2617) & (g1323) & (!g2665)) + ((g1255) & (g1283) & (g2578) & (g2617) & (!g1323) & (g2665)) + ((g1255) & (g1283) & (g2578) & (g2617) & (g1323) & (!g2665)));
	assign g5750 = (((!g1255) & (!g1283) & (!g2578) & (!g2617) & (!g1216) & (!g2529)) + ((!g1255) & (!g1283) & (!g2578) & (!g2617) & (!g1216) & (g2529)) + ((!g1255) & (!g1283) & (!g2578) & (!g2617) & (g1216) & (!g2529)) + ((!g1255) & (!g1283) & (!g2578) & (g2617) & (!g1216) & (!g2529)) + ((!g1255) & (!g1283) & (!g2578) & (g2617) & (!g1216) & (g2529)) + ((!g1255) & (!g1283) & (!g2578) & (g2617) & (g1216) & (!g2529)) + ((!g1255) & (!g1283) & (g2578) & (!g2617) & (!g1216) & (!g2529)) + ((!g1255) & (!g1283) & (g2578) & (!g2617) & (!g1216) & (g2529)) + ((!g1255) & (!g1283) & (g2578) & (!g2617) & (g1216) & (!g2529)) + ((!g1255) & (!g1283) & (g2578) & (g2617) & (!g1216) & (!g2529)) + ((!g1255) & (!g1283) & (g2578) & (g2617) & (!g1216) & (g2529)) + ((!g1255) & (!g1283) & (g2578) & (g2617) & (g1216) & (!g2529)) + ((!g1255) & (g1283) & (!g2578) & (!g2617) & (!g1216) & (!g2529)) + ((!g1255) & (g1283) & (!g2578) & (!g2617) & (!g1216) & (g2529)) + ((!g1255) & (g1283) & (!g2578) & (!g2617) & (g1216) & (!g2529)) + ((!g1255) & (g1283) & (g2578) & (!g2617) & (!g1216) & (!g2529)) + ((!g1255) & (g1283) & (g2578) & (!g2617) & (!g1216) & (g2529)) + ((!g1255) & (g1283) & (g2578) & (!g2617) & (g1216) & (!g2529)) + ((g1255) & (!g1283) & (!g2578) & (!g2617) & (!g1216) & (!g2529)) + ((g1255) & (!g1283) & (!g2578) & (!g2617) & (!g1216) & (g2529)) + ((g1255) & (!g1283) & (!g2578) & (!g2617) & (g1216) & (!g2529)) + ((g1255) & (!g1283) & (!g2578) & (g2617) & (!g1216) & (!g2529)) + ((g1255) & (!g1283) & (!g2578) & (g2617) & (!g1216) & (g2529)) + ((g1255) & (!g1283) & (!g2578) & (g2617) & (g1216) & (!g2529)) + ((g1255) & (g1283) & (!g2578) & (!g2617) & (!g1216) & (!g2529)) + ((g1255) & (g1283) & (!g2578) & (!g2617) & (!g1216) & (g2529)) + ((g1255) & (g1283) & (!g2578) & (!g2617) & (g1216) & (!g2529)));
	assign g5751 = (((!g1216) & (!g2529) & (g5749) & (!g5750)) + ((!g1216) & (g2529) & (g5749) & (!g5750)) + ((!g1216) & (g2529) & (g5749) & (g5750)) + ((g1216) & (!g2529) & (g5749) & (!g5750)) + ((g1216) & (!g2529) & (g5749) & (g5750)) + ((g1216) & (g2529) & (g5749) & (!g5750)) + ((g1216) & (g2529) & (g5749) & (g5750)));
	assign g5752 = (((!g1257) & (!g1291) & (g2581) & (g2629) & (!g1325) & (g2667)) + ((!g1257) & (!g1291) & (g2581) & (g2629) & (g1325) & (!g2667)) + ((!g1257) & (g1291) & (!g2581) & (g2629) & (!g1325) & (g2667)) + ((!g1257) & (g1291) & (!g2581) & (g2629) & (g1325) & (!g2667)) + ((!g1257) & (g1291) & (g2581) & (!g2629) & (!g1325) & (g2667)) + ((!g1257) & (g1291) & (g2581) & (!g2629) & (g1325) & (!g2667)) + ((!g1257) & (g1291) & (g2581) & (g2629) & (!g1325) & (g2667)) + ((!g1257) & (g1291) & (g2581) & (g2629) & (g1325) & (!g2667)) + ((g1257) & (!g1291) & (!g2581) & (g2629) & (!g1325) & (g2667)) + ((g1257) & (!g1291) & (!g2581) & (g2629) & (g1325) & (!g2667)) + ((g1257) & (!g1291) & (g2581) & (g2629) & (!g1325) & (g2667)) + ((g1257) & (!g1291) & (g2581) & (g2629) & (g1325) & (!g2667)) + ((g1257) & (g1291) & (!g2581) & (!g2629) & (!g1325) & (g2667)) + ((g1257) & (g1291) & (!g2581) & (!g2629) & (g1325) & (!g2667)) + ((g1257) & (g1291) & (!g2581) & (g2629) & (!g1325) & (g2667)) + ((g1257) & (g1291) & (!g2581) & (g2629) & (g1325) & (!g2667)) + ((g1257) & (g1291) & (g2581) & (!g2629) & (!g1325) & (g2667)) + ((g1257) & (g1291) & (g2581) & (!g2629) & (g1325) & (!g2667)) + ((g1257) & (g1291) & (g2581) & (g2629) & (!g1325) & (g2667)) + ((g1257) & (g1291) & (g2581) & (g2629) & (g1325) & (!g2667)));
	assign g5753 = (((!g1257) & (!g1291) & (!g2581) & (!g2629) & (!g1224) & (!g2537)) + ((!g1257) & (!g1291) & (!g2581) & (!g2629) & (!g1224) & (g2537)) + ((!g1257) & (!g1291) & (!g2581) & (!g2629) & (g1224) & (!g2537)) + ((!g1257) & (!g1291) & (!g2581) & (g2629) & (!g1224) & (!g2537)) + ((!g1257) & (!g1291) & (!g2581) & (g2629) & (!g1224) & (g2537)) + ((!g1257) & (!g1291) & (!g2581) & (g2629) & (g1224) & (!g2537)) + ((!g1257) & (!g1291) & (g2581) & (!g2629) & (!g1224) & (!g2537)) + ((!g1257) & (!g1291) & (g2581) & (!g2629) & (!g1224) & (g2537)) + ((!g1257) & (!g1291) & (g2581) & (!g2629) & (g1224) & (!g2537)) + ((!g1257) & (!g1291) & (g2581) & (g2629) & (!g1224) & (!g2537)) + ((!g1257) & (!g1291) & (g2581) & (g2629) & (!g1224) & (g2537)) + ((!g1257) & (!g1291) & (g2581) & (g2629) & (g1224) & (!g2537)) + ((!g1257) & (g1291) & (!g2581) & (!g2629) & (!g1224) & (!g2537)) + ((!g1257) & (g1291) & (!g2581) & (!g2629) & (!g1224) & (g2537)) + ((!g1257) & (g1291) & (!g2581) & (!g2629) & (g1224) & (!g2537)) + ((!g1257) & (g1291) & (g2581) & (!g2629) & (!g1224) & (!g2537)) + ((!g1257) & (g1291) & (g2581) & (!g2629) & (!g1224) & (g2537)) + ((!g1257) & (g1291) & (g2581) & (!g2629) & (g1224) & (!g2537)) + ((g1257) & (!g1291) & (!g2581) & (!g2629) & (!g1224) & (!g2537)) + ((g1257) & (!g1291) & (!g2581) & (!g2629) & (!g1224) & (g2537)) + ((g1257) & (!g1291) & (!g2581) & (!g2629) & (g1224) & (!g2537)) + ((g1257) & (!g1291) & (!g2581) & (g2629) & (!g1224) & (!g2537)) + ((g1257) & (!g1291) & (!g2581) & (g2629) & (!g1224) & (g2537)) + ((g1257) & (!g1291) & (!g2581) & (g2629) & (g1224) & (!g2537)) + ((g1257) & (g1291) & (!g2581) & (!g2629) & (!g1224) & (!g2537)) + ((g1257) & (g1291) & (!g2581) & (!g2629) & (!g1224) & (g2537)) + ((g1257) & (g1291) & (!g2581) & (!g2629) & (g1224) & (!g2537)));
	assign g5754 = (((!g1224) & (!g2537) & (g5752) & (!g5753)) + ((!g1224) & (g2537) & (g5752) & (!g5753)) + ((!g1224) & (g2537) & (g5752) & (g5753)) + ((g1224) & (!g2537) & (g5752) & (!g5753)) + ((g1224) & (!g2537) & (g5752) & (g5753)) + ((g1224) & (g2537) & (g5752) & (!g5753)) + ((g1224) & (g2537) & (g5752) & (g5753)));
	assign g5755 = (((!g1259) & (!g1299) & (g2584) & (g2640) & (!g1327) & (g2669)) + ((!g1259) & (!g1299) & (g2584) & (g2640) & (g1327) & (!g2669)) + ((!g1259) & (g1299) & (!g2584) & (g2640) & (!g1327) & (g2669)) + ((!g1259) & (g1299) & (!g2584) & (g2640) & (g1327) & (!g2669)) + ((!g1259) & (g1299) & (g2584) & (!g2640) & (!g1327) & (g2669)) + ((!g1259) & (g1299) & (g2584) & (!g2640) & (g1327) & (!g2669)) + ((!g1259) & (g1299) & (g2584) & (g2640) & (!g1327) & (g2669)) + ((!g1259) & (g1299) & (g2584) & (g2640) & (g1327) & (!g2669)) + ((g1259) & (!g1299) & (!g2584) & (g2640) & (!g1327) & (g2669)) + ((g1259) & (!g1299) & (!g2584) & (g2640) & (g1327) & (!g2669)) + ((g1259) & (!g1299) & (g2584) & (g2640) & (!g1327) & (g2669)) + ((g1259) & (!g1299) & (g2584) & (g2640) & (g1327) & (!g2669)) + ((g1259) & (g1299) & (!g2584) & (!g2640) & (!g1327) & (g2669)) + ((g1259) & (g1299) & (!g2584) & (!g2640) & (g1327) & (!g2669)) + ((g1259) & (g1299) & (!g2584) & (g2640) & (!g1327) & (g2669)) + ((g1259) & (g1299) & (!g2584) & (g2640) & (g1327) & (!g2669)) + ((g1259) & (g1299) & (g2584) & (!g2640) & (!g1327) & (g2669)) + ((g1259) & (g1299) & (g2584) & (!g2640) & (g1327) & (!g2669)) + ((g1259) & (g1299) & (g2584) & (g2640) & (!g1327) & (g2669)) + ((g1259) & (g1299) & (g2584) & (g2640) & (g1327) & (!g2669)));
	assign g5756 = (((!g1259) & (!g1299) & (!g2584) & (!g2640) & (!g1232) & (!g2544)) + ((!g1259) & (!g1299) & (!g2584) & (!g2640) & (!g1232) & (g2544)) + ((!g1259) & (!g1299) & (!g2584) & (!g2640) & (g1232) & (!g2544)) + ((!g1259) & (!g1299) & (!g2584) & (g2640) & (!g1232) & (!g2544)) + ((!g1259) & (!g1299) & (!g2584) & (g2640) & (!g1232) & (g2544)) + ((!g1259) & (!g1299) & (!g2584) & (g2640) & (g1232) & (!g2544)) + ((!g1259) & (!g1299) & (g2584) & (!g2640) & (!g1232) & (!g2544)) + ((!g1259) & (!g1299) & (g2584) & (!g2640) & (!g1232) & (g2544)) + ((!g1259) & (!g1299) & (g2584) & (!g2640) & (g1232) & (!g2544)) + ((!g1259) & (!g1299) & (g2584) & (g2640) & (!g1232) & (!g2544)) + ((!g1259) & (!g1299) & (g2584) & (g2640) & (!g1232) & (g2544)) + ((!g1259) & (!g1299) & (g2584) & (g2640) & (g1232) & (!g2544)) + ((!g1259) & (g1299) & (!g2584) & (!g2640) & (!g1232) & (!g2544)) + ((!g1259) & (g1299) & (!g2584) & (!g2640) & (!g1232) & (g2544)) + ((!g1259) & (g1299) & (!g2584) & (!g2640) & (g1232) & (!g2544)) + ((!g1259) & (g1299) & (g2584) & (!g2640) & (!g1232) & (!g2544)) + ((!g1259) & (g1299) & (g2584) & (!g2640) & (!g1232) & (g2544)) + ((!g1259) & (g1299) & (g2584) & (!g2640) & (g1232) & (!g2544)) + ((g1259) & (!g1299) & (!g2584) & (!g2640) & (!g1232) & (!g2544)) + ((g1259) & (!g1299) & (!g2584) & (!g2640) & (!g1232) & (g2544)) + ((g1259) & (!g1299) & (!g2584) & (!g2640) & (g1232) & (!g2544)) + ((g1259) & (!g1299) & (!g2584) & (g2640) & (!g1232) & (!g2544)) + ((g1259) & (!g1299) & (!g2584) & (g2640) & (!g1232) & (g2544)) + ((g1259) & (!g1299) & (!g2584) & (g2640) & (g1232) & (!g2544)) + ((g1259) & (g1299) & (!g2584) & (!g2640) & (!g1232) & (!g2544)) + ((g1259) & (g1299) & (!g2584) & (!g2640) & (!g1232) & (g2544)) + ((g1259) & (g1299) & (!g2584) & (!g2640) & (g1232) & (!g2544)));
	assign g5757 = (((!g1232) & (!g2544) & (g5755) & (!g5756)) + ((!g1232) & (g2544) & (g5755) & (!g5756)) + ((!g1232) & (g2544) & (g5755) & (g5756)) + ((g1232) & (!g2544) & (g5755) & (!g5756)) + ((g1232) & (!g2544) & (g5755) & (g5756)) + ((g1232) & (g2544) & (g5755) & (!g5756)) + ((g1232) & (g2544) & (g5755) & (g5756)));
	assign g5758 = (((!g1261) & (!g1277) & (g2012) & (g2014) & (!g1329) & (g2052)) + ((!g1261) & (!g1277) & (g2012) & (g2014) & (g1329) & (!g2052)) + ((!g1261) & (g1277) & (!g2012) & (g2014) & (!g1329) & (g2052)) + ((!g1261) & (g1277) & (!g2012) & (g2014) & (g1329) & (!g2052)) + ((!g1261) & (g1277) & (g2012) & (!g2014) & (!g1329) & (g2052)) + ((!g1261) & (g1277) & (g2012) & (!g2014) & (g1329) & (!g2052)) + ((!g1261) & (g1277) & (g2012) & (g2014) & (!g1329) & (g2052)) + ((!g1261) & (g1277) & (g2012) & (g2014) & (g1329) & (!g2052)) + ((g1261) & (!g1277) & (!g2012) & (g2014) & (!g1329) & (g2052)) + ((g1261) & (!g1277) & (!g2012) & (g2014) & (g1329) & (!g2052)) + ((g1261) & (!g1277) & (g2012) & (g2014) & (!g1329) & (g2052)) + ((g1261) & (!g1277) & (g2012) & (g2014) & (g1329) & (!g2052)) + ((g1261) & (g1277) & (!g2012) & (!g2014) & (!g1329) & (g2052)) + ((g1261) & (g1277) & (!g2012) & (!g2014) & (g1329) & (!g2052)) + ((g1261) & (g1277) & (!g2012) & (g2014) & (!g1329) & (g2052)) + ((g1261) & (g1277) & (!g2012) & (g2014) & (g1329) & (!g2052)) + ((g1261) & (g1277) & (g2012) & (!g2014) & (!g1329) & (g2052)) + ((g1261) & (g1277) & (g2012) & (!g2014) & (g1329) & (!g2052)) + ((g1261) & (g1277) & (g2012) & (g2014) & (!g1329) & (g2052)) + ((g1261) & (g1277) & (g2012) & (g2014) & (g1329) & (!g2052)));
	assign g5759 = (((!g1261) & (!g1277) & (!g2012) & (!g2014) & (!g1210) & (!g2006)) + ((!g1261) & (!g1277) & (!g2012) & (!g2014) & (!g1210) & (g2006)) + ((!g1261) & (!g1277) & (!g2012) & (!g2014) & (g1210) & (!g2006)) + ((!g1261) & (!g1277) & (!g2012) & (g2014) & (!g1210) & (!g2006)) + ((!g1261) & (!g1277) & (!g2012) & (g2014) & (!g1210) & (g2006)) + ((!g1261) & (!g1277) & (!g2012) & (g2014) & (g1210) & (!g2006)) + ((!g1261) & (!g1277) & (g2012) & (!g2014) & (!g1210) & (!g2006)) + ((!g1261) & (!g1277) & (g2012) & (!g2014) & (!g1210) & (g2006)) + ((!g1261) & (!g1277) & (g2012) & (!g2014) & (g1210) & (!g2006)) + ((!g1261) & (!g1277) & (g2012) & (g2014) & (!g1210) & (!g2006)) + ((!g1261) & (!g1277) & (g2012) & (g2014) & (!g1210) & (g2006)) + ((!g1261) & (!g1277) & (g2012) & (g2014) & (g1210) & (!g2006)) + ((!g1261) & (g1277) & (!g2012) & (!g2014) & (!g1210) & (!g2006)) + ((!g1261) & (g1277) & (!g2012) & (!g2014) & (!g1210) & (g2006)) + ((!g1261) & (g1277) & (!g2012) & (!g2014) & (g1210) & (!g2006)) + ((!g1261) & (g1277) & (g2012) & (!g2014) & (!g1210) & (!g2006)) + ((!g1261) & (g1277) & (g2012) & (!g2014) & (!g1210) & (g2006)) + ((!g1261) & (g1277) & (g2012) & (!g2014) & (g1210) & (!g2006)) + ((g1261) & (!g1277) & (!g2012) & (!g2014) & (!g1210) & (!g2006)) + ((g1261) & (!g1277) & (!g2012) & (!g2014) & (!g1210) & (g2006)) + ((g1261) & (!g1277) & (!g2012) & (!g2014) & (g1210) & (!g2006)) + ((g1261) & (!g1277) & (!g2012) & (g2014) & (!g1210) & (!g2006)) + ((g1261) & (!g1277) & (!g2012) & (g2014) & (!g1210) & (g2006)) + ((g1261) & (!g1277) & (!g2012) & (g2014) & (g1210) & (!g2006)) + ((g1261) & (g1277) & (!g2012) & (!g2014) & (!g1210) & (!g2006)) + ((g1261) & (g1277) & (!g2012) & (!g2014) & (!g1210) & (g2006)) + ((g1261) & (g1277) & (!g2012) & (!g2014) & (g1210) & (!g2006)));
	assign g5760 = (((!g1210) & (!g2006) & (g5758) & (!g5759)) + ((!g1210) & (g2006) & (g5758) & (!g5759)) + ((!g1210) & (g2006) & (g5758) & (g5759)) + ((g1210) & (!g2006) & (g5758) & (!g5759)) + ((g1210) & (!g2006) & (g5758) & (g5759)) + ((g1210) & (g2006) & (g5758) & (!g5759)) + ((g1210) & (g2006) & (g5758) & (g5759)));
	assign g5761 = (((!g1263) & (!g1285) & (g2589) & (g2620) & (!g1331) & (g2672)) + ((!g1263) & (!g1285) & (g2589) & (g2620) & (g1331) & (!g2672)) + ((!g1263) & (g1285) & (!g2589) & (g2620) & (!g1331) & (g2672)) + ((!g1263) & (g1285) & (!g2589) & (g2620) & (g1331) & (!g2672)) + ((!g1263) & (g1285) & (g2589) & (!g2620) & (!g1331) & (g2672)) + ((!g1263) & (g1285) & (g2589) & (!g2620) & (g1331) & (!g2672)) + ((!g1263) & (g1285) & (g2589) & (g2620) & (!g1331) & (g2672)) + ((!g1263) & (g1285) & (g2589) & (g2620) & (g1331) & (!g2672)) + ((g1263) & (!g1285) & (!g2589) & (g2620) & (!g1331) & (g2672)) + ((g1263) & (!g1285) & (!g2589) & (g2620) & (g1331) & (!g2672)) + ((g1263) & (!g1285) & (g2589) & (g2620) & (!g1331) & (g2672)) + ((g1263) & (!g1285) & (g2589) & (g2620) & (g1331) & (!g2672)) + ((g1263) & (g1285) & (!g2589) & (!g2620) & (!g1331) & (g2672)) + ((g1263) & (g1285) & (!g2589) & (!g2620) & (g1331) & (!g2672)) + ((g1263) & (g1285) & (!g2589) & (g2620) & (!g1331) & (g2672)) + ((g1263) & (g1285) & (!g2589) & (g2620) & (g1331) & (!g2672)) + ((g1263) & (g1285) & (g2589) & (!g2620) & (!g1331) & (g2672)) + ((g1263) & (g1285) & (g2589) & (!g2620) & (g1331) & (!g2672)) + ((g1263) & (g1285) & (g2589) & (g2620) & (!g1331) & (g2672)) + ((g1263) & (g1285) & (g2589) & (g2620) & (g1331) & (!g2672)));
	assign g5762 = (((!g1263) & (!g1285) & (!g2589) & (!g2620) & (!g1218) & (!g2531)) + ((!g1263) & (!g1285) & (!g2589) & (!g2620) & (!g1218) & (g2531)) + ((!g1263) & (!g1285) & (!g2589) & (!g2620) & (g1218) & (!g2531)) + ((!g1263) & (!g1285) & (!g2589) & (g2620) & (!g1218) & (!g2531)) + ((!g1263) & (!g1285) & (!g2589) & (g2620) & (!g1218) & (g2531)) + ((!g1263) & (!g1285) & (!g2589) & (g2620) & (g1218) & (!g2531)) + ((!g1263) & (!g1285) & (g2589) & (!g2620) & (!g1218) & (!g2531)) + ((!g1263) & (!g1285) & (g2589) & (!g2620) & (!g1218) & (g2531)) + ((!g1263) & (!g1285) & (g2589) & (!g2620) & (g1218) & (!g2531)) + ((!g1263) & (!g1285) & (g2589) & (g2620) & (!g1218) & (!g2531)) + ((!g1263) & (!g1285) & (g2589) & (g2620) & (!g1218) & (g2531)) + ((!g1263) & (!g1285) & (g2589) & (g2620) & (g1218) & (!g2531)) + ((!g1263) & (g1285) & (!g2589) & (!g2620) & (!g1218) & (!g2531)) + ((!g1263) & (g1285) & (!g2589) & (!g2620) & (!g1218) & (g2531)) + ((!g1263) & (g1285) & (!g2589) & (!g2620) & (g1218) & (!g2531)) + ((!g1263) & (g1285) & (g2589) & (!g2620) & (!g1218) & (!g2531)) + ((!g1263) & (g1285) & (g2589) & (!g2620) & (!g1218) & (g2531)) + ((!g1263) & (g1285) & (g2589) & (!g2620) & (g1218) & (!g2531)) + ((g1263) & (!g1285) & (!g2589) & (!g2620) & (!g1218) & (!g2531)) + ((g1263) & (!g1285) & (!g2589) & (!g2620) & (!g1218) & (g2531)) + ((g1263) & (!g1285) & (!g2589) & (!g2620) & (g1218) & (!g2531)) + ((g1263) & (!g1285) & (!g2589) & (g2620) & (!g1218) & (!g2531)) + ((g1263) & (!g1285) & (!g2589) & (g2620) & (!g1218) & (g2531)) + ((g1263) & (!g1285) & (!g2589) & (g2620) & (g1218) & (!g2531)) + ((g1263) & (g1285) & (!g2589) & (!g2620) & (!g1218) & (!g2531)) + ((g1263) & (g1285) & (!g2589) & (!g2620) & (!g1218) & (g2531)) + ((g1263) & (g1285) & (!g2589) & (!g2620) & (g1218) & (!g2531)));
	assign g5763 = (((!g1218) & (!g2531) & (g5761) & (!g5762)) + ((!g1218) & (g2531) & (g5761) & (!g5762)) + ((!g1218) & (g2531) & (g5761) & (g5762)) + ((g1218) & (!g2531) & (g5761) & (!g5762)) + ((g1218) & (!g2531) & (g5761) & (g5762)) + ((g1218) & (g2531) & (g5761) & (!g5762)) + ((g1218) & (g2531) & (g5761) & (g5762)));
	assign g5764 = (((!g1265) & (!g1293) & (g2592) & (g2632) & (!g1333) & (g2674)) + ((!g1265) & (!g1293) & (g2592) & (g2632) & (g1333) & (!g2674)) + ((!g1265) & (g1293) & (!g2592) & (g2632) & (!g1333) & (g2674)) + ((!g1265) & (g1293) & (!g2592) & (g2632) & (g1333) & (!g2674)) + ((!g1265) & (g1293) & (g2592) & (!g2632) & (!g1333) & (g2674)) + ((!g1265) & (g1293) & (g2592) & (!g2632) & (g1333) & (!g2674)) + ((!g1265) & (g1293) & (g2592) & (g2632) & (!g1333) & (g2674)) + ((!g1265) & (g1293) & (g2592) & (g2632) & (g1333) & (!g2674)) + ((g1265) & (!g1293) & (!g2592) & (g2632) & (!g1333) & (g2674)) + ((g1265) & (!g1293) & (!g2592) & (g2632) & (g1333) & (!g2674)) + ((g1265) & (!g1293) & (g2592) & (g2632) & (!g1333) & (g2674)) + ((g1265) & (!g1293) & (g2592) & (g2632) & (g1333) & (!g2674)) + ((g1265) & (g1293) & (!g2592) & (!g2632) & (!g1333) & (g2674)) + ((g1265) & (g1293) & (!g2592) & (!g2632) & (g1333) & (!g2674)) + ((g1265) & (g1293) & (!g2592) & (g2632) & (!g1333) & (g2674)) + ((g1265) & (g1293) & (!g2592) & (g2632) & (g1333) & (!g2674)) + ((g1265) & (g1293) & (g2592) & (!g2632) & (!g1333) & (g2674)) + ((g1265) & (g1293) & (g2592) & (!g2632) & (g1333) & (!g2674)) + ((g1265) & (g1293) & (g2592) & (g2632) & (!g1333) & (g2674)) + ((g1265) & (g1293) & (g2592) & (g2632) & (g1333) & (!g2674)));
	assign g5765 = (((!g1265) & (!g1293) & (!g2592) & (!g2632) & (!g1226) & (!g2539)) + ((!g1265) & (!g1293) & (!g2592) & (!g2632) & (!g1226) & (g2539)) + ((!g1265) & (!g1293) & (!g2592) & (!g2632) & (g1226) & (!g2539)) + ((!g1265) & (!g1293) & (!g2592) & (g2632) & (!g1226) & (!g2539)) + ((!g1265) & (!g1293) & (!g2592) & (g2632) & (!g1226) & (g2539)) + ((!g1265) & (!g1293) & (!g2592) & (g2632) & (g1226) & (!g2539)) + ((!g1265) & (!g1293) & (g2592) & (!g2632) & (!g1226) & (!g2539)) + ((!g1265) & (!g1293) & (g2592) & (!g2632) & (!g1226) & (g2539)) + ((!g1265) & (!g1293) & (g2592) & (!g2632) & (g1226) & (!g2539)) + ((!g1265) & (!g1293) & (g2592) & (g2632) & (!g1226) & (!g2539)) + ((!g1265) & (!g1293) & (g2592) & (g2632) & (!g1226) & (g2539)) + ((!g1265) & (!g1293) & (g2592) & (g2632) & (g1226) & (!g2539)) + ((!g1265) & (g1293) & (!g2592) & (!g2632) & (!g1226) & (!g2539)) + ((!g1265) & (g1293) & (!g2592) & (!g2632) & (!g1226) & (g2539)) + ((!g1265) & (g1293) & (!g2592) & (!g2632) & (g1226) & (!g2539)) + ((!g1265) & (g1293) & (g2592) & (!g2632) & (!g1226) & (!g2539)) + ((!g1265) & (g1293) & (g2592) & (!g2632) & (!g1226) & (g2539)) + ((!g1265) & (g1293) & (g2592) & (!g2632) & (g1226) & (!g2539)) + ((g1265) & (!g1293) & (!g2592) & (!g2632) & (!g1226) & (!g2539)) + ((g1265) & (!g1293) & (!g2592) & (!g2632) & (!g1226) & (g2539)) + ((g1265) & (!g1293) & (!g2592) & (!g2632) & (g1226) & (!g2539)) + ((g1265) & (!g1293) & (!g2592) & (g2632) & (!g1226) & (!g2539)) + ((g1265) & (!g1293) & (!g2592) & (g2632) & (!g1226) & (g2539)) + ((g1265) & (!g1293) & (!g2592) & (g2632) & (g1226) & (!g2539)) + ((g1265) & (g1293) & (!g2592) & (!g2632) & (!g1226) & (!g2539)) + ((g1265) & (g1293) & (!g2592) & (!g2632) & (!g1226) & (g2539)) + ((g1265) & (g1293) & (!g2592) & (!g2632) & (g1226) & (!g2539)));
	assign g5766 = (((!g1226) & (!g2539) & (g5764) & (!g5765)) + ((!g1226) & (g2539) & (g5764) & (!g5765)) + ((!g1226) & (g2539) & (g5764) & (g5765)) + ((g1226) & (!g2539) & (g5764) & (!g5765)) + ((g1226) & (!g2539) & (g5764) & (g5765)) + ((g1226) & (g2539) & (g5764) & (!g5765)) + ((g1226) & (g2539) & (g5764) & (g5765)));
	assign g5767 = (((!g1267) & (!g1301) & (g2595) & (g2643) & (!g1335) & (g2676)) + ((!g1267) & (!g1301) & (g2595) & (g2643) & (g1335) & (!g2676)) + ((!g1267) & (g1301) & (!g2595) & (g2643) & (!g1335) & (g2676)) + ((!g1267) & (g1301) & (!g2595) & (g2643) & (g1335) & (!g2676)) + ((!g1267) & (g1301) & (g2595) & (!g2643) & (!g1335) & (g2676)) + ((!g1267) & (g1301) & (g2595) & (!g2643) & (g1335) & (!g2676)) + ((!g1267) & (g1301) & (g2595) & (g2643) & (!g1335) & (g2676)) + ((!g1267) & (g1301) & (g2595) & (g2643) & (g1335) & (!g2676)) + ((g1267) & (!g1301) & (!g2595) & (g2643) & (!g1335) & (g2676)) + ((g1267) & (!g1301) & (!g2595) & (g2643) & (g1335) & (!g2676)) + ((g1267) & (!g1301) & (g2595) & (g2643) & (!g1335) & (g2676)) + ((g1267) & (!g1301) & (g2595) & (g2643) & (g1335) & (!g2676)) + ((g1267) & (g1301) & (!g2595) & (!g2643) & (!g1335) & (g2676)) + ((g1267) & (g1301) & (!g2595) & (!g2643) & (g1335) & (!g2676)) + ((g1267) & (g1301) & (!g2595) & (g2643) & (!g1335) & (g2676)) + ((g1267) & (g1301) & (!g2595) & (g2643) & (g1335) & (!g2676)) + ((g1267) & (g1301) & (g2595) & (!g2643) & (!g1335) & (g2676)) + ((g1267) & (g1301) & (g2595) & (!g2643) & (g1335) & (!g2676)) + ((g1267) & (g1301) & (g2595) & (g2643) & (!g1335) & (g2676)) + ((g1267) & (g1301) & (g2595) & (g2643) & (g1335) & (!g2676)));
	assign g5768 = (((!g1267) & (!g1301) & (!g2595) & (!g2643) & (!g1234) & (!g2546)) + ((!g1267) & (!g1301) & (!g2595) & (!g2643) & (!g1234) & (g2546)) + ((!g1267) & (!g1301) & (!g2595) & (!g2643) & (g1234) & (!g2546)) + ((!g1267) & (!g1301) & (!g2595) & (g2643) & (!g1234) & (!g2546)) + ((!g1267) & (!g1301) & (!g2595) & (g2643) & (!g1234) & (g2546)) + ((!g1267) & (!g1301) & (!g2595) & (g2643) & (g1234) & (!g2546)) + ((!g1267) & (!g1301) & (g2595) & (!g2643) & (!g1234) & (!g2546)) + ((!g1267) & (!g1301) & (g2595) & (!g2643) & (!g1234) & (g2546)) + ((!g1267) & (!g1301) & (g2595) & (!g2643) & (g1234) & (!g2546)) + ((!g1267) & (!g1301) & (g2595) & (g2643) & (!g1234) & (!g2546)) + ((!g1267) & (!g1301) & (g2595) & (g2643) & (!g1234) & (g2546)) + ((!g1267) & (!g1301) & (g2595) & (g2643) & (g1234) & (!g2546)) + ((!g1267) & (g1301) & (!g2595) & (!g2643) & (!g1234) & (!g2546)) + ((!g1267) & (g1301) & (!g2595) & (!g2643) & (!g1234) & (g2546)) + ((!g1267) & (g1301) & (!g2595) & (!g2643) & (g1234) & (!g2546)) + ((!g1267) & (g1301) & (g2595) & (!g2643) & (!g1234) & (!g2546)) + ((!g1267) & (g1301) & (g2595) & (!g2643) & (!g1234) & (g2546)) + ((!g1267) & (g1301) & (g2595) & (!g2643) & (g1234) & (!g2546)) + ((g1267) & (!g1301) & (!g2595) & (!g2643) & (!g1234) & (!g2546)) + ((g1267) & (!g1301) & (!g2595) & (!g2643) & (!g1234) & (g2546)) + ((g1267) & (!g1301) & (!g2595) & (!g2643) & (g1234) & (!g2546)) + ((g1267) & (!g1301) & (!g2595) & (g2643) & (!g1234) & (!g2546)) + ((g1267) & (!g1301) & (!g2595) & (g2643) & (!g1234) & (g2546)) + ((g1267) & (!g1301) & (!g2595) & (g2643) & (g1234) & (!g2546)) + ((g1267) & (g1301) & (!g2595) & (!g2643) & (!g1234) & (!g2546)) + ((g1267) & (g1301) & (!g2595) & (!g2643) & (!g1234) & (g2546)) + ((g1267) & (g1301) & (!g2595) & (!g2643) & (g1234) & (!g2546)));
	assign g5769 = (((!g1234) & (!g2546) & (g5767) & (!g5768)) + ((!g1234) & (g2546) & (g5767) & (!g5768)) + ((!g1234) & (g2546) & (g5767) & (g5768)) + ((g1234) & (!g2546) & (g5767) & (!g5768)) + ((g1234) & (!g2546) & (g5767) & (g5768)) + ((g1234) & (g2546) & (g5767) & (!g5768)) + ((g1234) & (g2546) & (g5767) & (g5768)));
	assign g5770 = (((!g2575) & (!g2607) & (g2584) & (g2640) & (!g2663) & (g2669)) + ((!g2575) & (!g2607) & (g2584) & (g2640) & (g2663) & (!g2669)) + ((!g2575) & (g2607) & (!g2584) & (g2640) & (!g2663) & (g2669)) + ((!g2575) & (g2607) & (!g2584) & (g2640) & (g2663) & (!g2669)) + ((!g2575) & (g2607) & (g2584) & (!g2640) & (!g2663) & (g2669)) + ((!g2575) & (g2607) & (g2584) & (!g2640) & (g2663) & (!g2669)) + ((!g2575) & (g2607) & (g2584) & (g2640) & (!g2663) & (g2669)) + ((!g2575) & (g2607) & (g2584) & (g2640) & (g2663) & (!g2669)) + ((g2575) & (!g2607) & (!g2584) & (g2640) & (!g2663) & (g2669)) + ((g2575) & (!g2607) & (!g2584) & (g2640) & (g2663) & (!g2669)) + ((g2575) & (!g2607) & (g2584) & (g2640) & (!g2663) & (g2669)) + ((g2575) & (!g2607) & (g2584) & (g2640) & (g2663) & (!g2669)) + ((g2575) & (g2607) & (!g2584) & (!g2640) & (!g2663) & (g2669)) + ((g2575) & (g2607) & (!g2584) & (!g2640) & (g2663) & (!g2669)) + ((g2575) & (g2607) & (!g2584) & (g2640) & (!g2663) & (g2669)) + ((g2575) & (g2607) & (!g2584) & (g2640) & (g2663) & (!g2669)) + ((g2575) & (g2607) & (g2584) & (!g2640) & (!g2663) & (g2669)) + ((g2575) & (g2607) & (g2584) & (!g2640) & (g2663) & (!g2669)) + ((g2575) & (g2607) & (g2584) & (g2640) & (!g2663) & (g2669)) + ((g2575) & (g2607) & (g2584) & (g2640) & (g2663) & (!g2669)));
	assign g5771 = (((!g2575) & (!g2607) & (!g2584) & (!g2640) & (!g2523) & (!g2544)) + ((!g2575) & (!g2607) & (!g2584) & (!g2640) & (!g2523) & (g2544)) + ((!g2575) & (!g2607) & (!g2584) & (!g2640) & (g2523) & (!g2544)) + ((!g2575) & (!g2607) & (!g2584) & (g2640) & (!g2523) & (!g2544)) + ((!g2575) & (!g2607) & (!g2584) & (g2640) & (!g2523) & (g2544)) + ((!g2575) & (!g2607) & (!g2584) & (g2640) & (g2523) & (!g2544)) + ((!g2575) & (!g2607) & (g2584) & (!g2640) & (!g2523) & (!g2544)) + ((!g2575) & (!g2607) & (g2584) & (!g2640) & (!g2523) & (g2544)) + ((!g2575) & (!g2607) & (g2584) & (!g2640) & (g2523) & (!g2544)) + ((!g2575) & (!g2607) & (g2584) & (g2640) & (!g2523) & (!g2544)) + ((!g2575) & (!g2607) & (g2584) & (g2640) & (!g2523) & (g2544)) + ((!g2575) & (!g2607) & (g2584) & (g2640) & (g2523) & (!g2544)) + ((!g2575) & (g2607) & (!g2584) & (!g2640) & (!g2523) & (!g2544)) + ((!g2575) & (g2607) & (!g2584) & (!g2640) & (!g2523) & (g2544)) + ((!g2575) & (g2607) & (!g2584) & (!g2640) & (g2523) & (!g2544)) + ((!g2575) & (g2607) & (g2584) & (!g2640) & (!g2523) & (!g2544)) + ((!g2575) & (g2607) & (g2584) & (!g2640) & (!g2523) & (g2544)) + ((!g2575) & (g2607) & (g2584) & (!g2640) & (g2523) & (!g2544)) + ((g2575) & (!g2607) & (!g2584) & (!g2640) & (!g2523) & (!g2544)) + ((g2575) & (!g2607) & (!g2584) & (!g2640) & (!g2523) & (g2544)) + ((g2575) & (!g2607) & (!g2584) & (!g2640) & (g2523) & (!g2544)) + ((g2575) & (!g2607) & (!g2584) & (g2640) & (!g2523) & (!g2544)) + ((g2575) & (!g2607) & (!g2584) & (g2640) & (!g2523) & (g2544)) + ((g2575) & (!g2607) & (!g2584) & (g2640) & (g2523) & (!g2544)) + ((g2575) & (g2607) & (!g2584) & (!g2640) & (!g2523) & (!g2544)) + ((g2575) & (g2607) & (!g2584) & (!g2640) & (!g2523) & (g2544)) + ((g2575) & (g2607) & (!g2584) & (!g2640) & (g2523) & (!g2544)));
	assign g5772 = (((!g2523) & (!g2544) & (g5770) & (!g5771)) + ((!g2523) & (g2544) & (g5770) & (!g5771)) + ((!g2523) & (g2544) & (g5770) & (g5771)) + ((g2523) & (!g2544) & (g5770) & (!g5771)) + ((g2523) & (!g2544) & (g5770) & (g5771)) + ((g2523) & (g2544) & (g5770) & (!g5771)) + ((g2523) & (g2544) & (g5770) & (g5771)));
	assign g5773 = (((!g2589) & (!g2620) & (g2592) & (g2632) & (!g2672) & (g2674)) + ((!g2589) & (!g2620) & (g2592) & (g2632) & (g2672) & (!g2674)) + ((!g2589) & (g2620) & (!g2592) & (g2632) & (!g2672) & (g2674)) + ((!g2589) & (g2620) & (!g2592) & (g2632) & (g2672) & (!g2674)) + ((!g2589) & (g2620) & (g2592) & (!g2632) & (!g2672) & (g2674)) + ((!g2589) & (g2620) & (g2592) & (!g2632) & (g2672) & (!g2674)) + ((!g2589) & (g2620) & (g2592) & (g2632) & (!g2672) & (g2674)) + ((!g2589) & (g2620) & (g2592) & (g2632) & (g2672) & (!g2674)) + ((g2589) & (!g2620) & (!g2592) & (g2632) & (!g2672) & (g2674)) + ((g2589) & (!g2620) & (!g2592) & (g2632) & (g2672) & (!g2674)) + ((g2589) & (!g2620) & (g2592) & (g2632) & (!g2672) & (g2674)) + ((g2589) & (!g2620) & (g2592) & (g2632) & (g2672) & (!g2674)) + ((g2589) & (g2620) & (!g2592) & (!g2632) & (!g2672) & (g2674)) + ((g2589) & (g2620) & (!g2592) & (!g2632) & (g2672) & (!g2674)) + ((g2589) & (g2620) & (!g2592) & (g2632) & (!g2672) & (g2674)) + ((g2589) & (g2620) & (!g2592) & (g2632) & (g2672) & (!g2674)) + ((g2589) & (g2620) & (g2592) & (!g2632) & (!g2672) & (g2674)) + ((g2589) & (g2620) & (g2592) & (!g2632) & (g2672) & (!g2674)) + ((g2589) & (g2620) & (g2592) & (g2632) & (!g2672) & (g2674)) + ((g2589) & (g2620) & (g2592) & (g2632) & (g2672) & (!g2674)));
	assign g5774 = (((!g2589) & (!g2620) & (!g2592) & (!g2632) & (!g2531) & (!g2539)) + ((!g2589) & (!g2620) & (!g2592) & (!g2632) & (!g2531) & (g2539)) + ((!g2589) & (!g2620) & (!g2592) & (!g2632) & (g2531) & (!g2539)) + ((!g2589) & (!g2620) & (!g2592) & (g2632) & (!g2531) & (!g2539)) + ((!g2589) & (!g2620) & (!g2592) & (g2632) & (!g2531) & (g2539)) + ((!g2589) & (!g2620) & (!g2592) & (g2632) & (g2531) & (!g2539)) + ((!g2589) & (!g2620) & (g2592) & (!g2632) & (!g2531) & (!g2539)) + ((!g2589) & (!g2620) & (g2592) & (!g2632) & (!g2531) & (g2539)) + ((!g2589) & (!g2620) & (g2592) & (!g2632) & (g2531) & (!g2539)) + ((!g2589) & (!g2620) & (g2592) & (g2632) & (!g2531) & (!g2539)) + ((!g2589) & (!g2620) & (g2592) & (g2632) & (!g2531) & (g2539)) + ((!g2589) & (!g2620) & (g2592) & (g2632) & (g2531) & (!g2539)) + ((!g2589) & (g2620) & (!g2592) & (!g2632) & (!g2531) & (!g2539)) + ((!g2589) & (g2620) & (!g2592) & (!g2632) & (!g2531) & (g2539)) + ((!g2589) & (g2620) & (!g2592) & (!g2632) & (g2531) & (!g2539)) + ((!g2589) & (g2620) & (g2592) & (!g2632) & (!g2531) & (!g2539)) + ((!g2589) & (g2620) & (g2592) & (!g2632) & (!g2531) & (g2539)) + ((!g2589) & (g2620) & (g2592) & (!g2632) & (g2531) & (!g2539)) + ((g2589) & (!g2620) & (!g2592) & (!g2632) & (!g2531) & (!g2539)) + ((g2589) & (!g2620) & (!g2592) & (!g2632) & (!g2531) & (g2539)) + ((g2589) & (!g2620) & (!g2592) & (!g2632) & (g2531) & (!g2539)) + ((g2589) & (!g2620) & (!g2592) & (g2632) & (!g2531) & (!g2539)) + ((g2589) & (!g2620) & (!g2592) & (g2632) & (!g2531) & (g2539)) + ((g2589) & (!g2620) & (!g2592) & (g2632) & (g2531) & (!g2539)) + ((g2589) & (g2620) & (!g2592) & (!g2632) & (!g2531) & (!g2539)) + ((g2589) & (g2620) & (!g2592) & (!g2632) & (!g2531) & (g2539)) + ((g2589) & (g2620) & (!g2592) & (!g2632) & (g2531) & (!g2539)));
	assign g5775 = (((!g2531) & (!g2539) & (g5773) & (!g5774)) + ((!g2531) & (g2539) & (g5773) & (!g5774)) + ((!g2531) & (g2539) & (g5773) & (g5774)) + ((g2531) & (!g2539) & (g5773) & (!g5774)) + ((g2531) & (!g2539) & (g5773) & (g5774)) + ((g2531) & (g2539) & (g5773) & (!g5774)) + ((g2531) & (g2539) & (g5773) & (g5774)));
	assign g5776 = (((!g3284) & (!g3245) & (!g3310) & (!g3314) & (!g3207) & (!g3213)) + ((!g3284) & (!g3245) & (!g3310) & (!g3314) & (!g3207) & (g3213)) + ((!g3284) & (!g3245) & (!g3310) & (!g3314) & (g3207) & (!g3213)) + ((!g3284) & (!g3245) & (!g3310) & (!g3314) & (g3207) & (g3213)) + ((!g3284) & (!g3245) & (!g3310) & (g3314) & (!g3207) & (!g3213)) + ((!g3284) & (!g3245) & (!g3310) & (g3314) & (!g3207) & (g3213)) + ((!g3284) & (!g3245) & (!g3310) & (g3314) & (g3207) & (!g3213)) + ((!g3284) & (!g3245) & (!g3310) & (g3314) & (g3207) & (g3213)) + ((!g3284) & (!g3245) & (g3310) & (!g3314) & (!g3207) & (!g3213)) + ((!g3284) & (!g3245) & (g3310) & (!g3314) & (!g3207) & (g3213)) + ((!g3284) & (!g3245) & (g3310) & (!g3314) & (g3207) & (!g3213)) + ((!g3284) & (!g3245) & (g3310) & (!g3314) & (g3207) & (g3213)) + ((!g3284) & (g3245) & (!g3310) & (!g3314) & (!g3207) & (!g3213)) + ((!g3284) & (g3245) & (!g3310) & (!g3314) & (!g3207) & (g3213)) + ((!g3284) & (g3245) & (!g3310) & (!g3314) & (g3207) & (!g3213)) + ((!g3284) & (g3245) & (!g3310) & (!g3314) & (g3207) & (g3213)) + ((!g3284) & (g3245) & (!g3310) & (g3314) & (!g3207) & (!g3213)) + ((!g3284) & (g3245) & (g3310) & (!g3314) & (!g3207) & (!g3213)) + ((g3284) & (!g3245) & (!g3310) & (!g3314) & (!g3207) & (!g3213)) + ((g3284) & (!g3245) & (!g3310) & (!g3314) & (!g3207) & (g3213)) + ((g3284) & (!g3245) & (!g3310) & (!g3314) & (g3207) & (!g3213)) + ((g3284) & (!g3245) & (!g3310) & (!g3314) & (g3207) & (g3213)) + ((g3284) & (!g3245) & (!g3310) & (g3314) & (!g3207) & (!g3213)) + ((g3284) & (!g3245) & (g3310) & (!g3314) & (!g3207) & (!g3213)) + ((g3284) & (g3245) & (!g3310) & (!g3314) & (!g3207) & (!g3213)) + ((g3284) & (g3245) & (!g3310) & (!g3314) & (!g3207) & (g3213)) + ((g3284) & (g3245) & (!g3310) & (!g3314) & (g3207) & (!g3213)) + ((g3284) & (g3245) & (!g3310) & (!g3314) & (g3207) & (g3213)));
	assign g5777 = (((!g3284) & (!g3245) & (!g3310) & (!g3314) & (!g3207) & (!g3213)) + ((!g3284) & (!g3245) & (!g3310) & (!g3314) & (!g3207) & (g3213)) + ((!g3284) & (!g3245) & (!g3310) & (!g3314) & (g3207) & (!g3213)) + ((!g3284) & (!g3245) & (!g3310) & (g3314) & (!g3207) & (!g3213)) + ((!g3284) & (!g3245) & (!g3310) & (g3314) & (!g3207) & (g3213)) + ((!g3284) & (!g3245) & (!g3310) & (g3314) & (g3207) & (!g3213)) + ((!g3284) & (!g3245) & (g3310) & (!g3314) & (!g3207) & (!g3213)) + ((!g3284) & (!g3245) & (g3310) & (!g3314) & (!g3207) & (g3213)) + ((!g3284) & (!g3245) & (g3310) & (!g3314) & (g3207) & (!g3213)) + ((!g3284) & (g3245) & (!g3310) & (!g3314) & (!g3207) & (!g3213)) + ((!g3284) & (g3245) & (!g3310) & (!g3314) & (!g3207) & (g3213)) + ((!g3284) & (g3245) & (!g3310) & (!g3314) & (g3207) & (!g3213)) + ((!g3284) & (g3245) & (!g3310) & (g3314) & (!g3207) & (!g3213)) + ((!g3284) & (g3245) & (!g3310) & (g3314) & (!g3207) & (g3213)) + ((!g3284) & (g3245) & (!g3310) & (g3314) & (g3207) & (!g3213)) + ((!g3284) & (g3245) & (g3310) & (!g3314) & (!g3207) & (!g3213)) + ((!g3284) & (g3245) & (g3310) & (!g3314) & (!g3207) & (g3213)) + ((!g3284) & (g3245) & (g3310) & (!g3314) & (g3207) & (!g3213)) + ((g3284) & (!g3245) & (!g3310) & (!g3314) & (!g3207) & (!g3213)) + ((g3284) & (!g3245) & (!g3310) & (!g3314) & (!g3207) & (g3213)) + ((g3284) & (!g3245) & (!g3310) & (!g3314) & (g3207) & (!g3213)) + ((g3284) & (!g3245) & (!g3310) & (g3314) & (!g3207) & (!g3213)) + ((g3284) & (!g3245) & (!g3310) & (g3314) & (!g3207) & (g3213)) + ((g3284) & (!g3245) & (!g3310) & (g3314) & (g3207) & (!g3213)) + ((g3284) & (!g3245) & (g3310) & (!g3314) & (!g3207) & (!g3213)) + ((g3284) & (!g3245) & (g3310) & (!g3314) & (!g3207) & (g3213)) + ((g3284) & (!g3245) & (g3310) & (!g3314) & (g3207) & (!g3213)));
	assign g5778 = (((!g2129) & (!g2177) & (g2776) & (g2807) & (!g2210) & (g2857)) + ((!g2129) & (!g2177) & (g2776) & (g2807) & (g2210) & (!g2857)) + ((!g2129) & (g2177) & (!g2776) & (g2807) & (!g2210) & (g2857)) + ((!g2129) & (g2177) & (!g2776) & (g2807) & (g2210) & (!g2857)) + ((!g2129) & (g2177) & (g2776) & (!g2807) & (!g2210) & (g2857)) + ((!g2129) & (g2177) & (g2776) & (!g2807) & (g2210) & (!g2857)) + ((!g2129) & (g2177) & (g2776) & (g2807) & (!g2210) & (g2857)) + ((!g2129) & (g2177) & (g2776) & (g2807) & (g2210) & (!g2857)) + ((g2129) & (!g2177) & (!g2776) & (g2807) & (!g2210) & (g2857)) + ((g2129) & (!g2177) & (!g2776) & (g2807) & (g2210) & (!g2857)) + ((g2129) & (!g2177) & (g2776) & (g2807) & (!g2210) & (g2857)) + ((g2129) & (!g2177) & (g2776) & (g2807) & (g2210) & (!g2857)) + ((g2129) & (g2177) & (!g2776) & (!g2807) & (!g2210) & (g2857)) + ((g2129) & (g2177) & (!g2776) & (!g2807) & (g2210) & (!g2857)) + ((g2129) & (g2177) & (!g2776) & (g2807) & (!g2210) & (g2857)) + ((g2129) & (g2177) & (!g2776) & (g2807) & (g2210) & (!g2857)) + ((g2129) & (g2177) & (g2776) & (!g2807) & (!g2210) & (g2857)) + ((g2129) & (g2177) & (g2776) & (!g2807) & (g2210) & (!g2857)) + ((g2129) & (g2177) & (g2776) & (g2807) & (!g2210) & (g2857)) + ((g2129) & (g2177) & (g2776) & (g2807) & (g2210) & (!g2857)));
	assign g5779 = (((!g2129) & (!g2177) & (!g2776) & (!g2807) & (!g2098) & (!g2708)) + ((!g2129) & (!g2177) & (!g2776) & (!g2807) & (!g2098) & (g2708)) + ((!g2129) & (!g2177) & (!g2776) & (!g2807) & (g2098) & (!g2708)) + ((!g2129) & (!g2177) & (!g2776) & (g2807) & (!g2098) & (!g2708)) + ((!g2129) & (!g2177) & (!g2776) & (g2807) & (!g2098) & (g2708)) + ((!g2129) & (!g2177) & (!g2776) & (g2807) & (g2098) & (!g2708)) + ((!g2129) & (!g2177) & (g2776) & (!g2807) & (!g2098) & (!g2708)) + ((!g2129) & (!g2177) & (g2776) & (!g2807) & (!g2098) & (g2708)) + ((!g2129) & (!g2177) & (g2776) & (!g2807) & (g2098) & (!g2708)) + ((!g2129) & (!g2177) & (g2776) & (g2807) & (!g2098) & (!g2708)) + ((!g2129) & (!g2177) & (g2776) & (g2807) & (!g2098) & (g2708)) + ((!g2129) & (!g2177) & (g2776) & (g2807) & (g2098) & (!g2708)) + ((!g2129) & (g2177) & (!g2776) & (!g2807) & (!g2098) & (!g2708)) + ((!g2129) & (g2177) & (!g2776) & (!g2807) & (!g2098) & (g2708)) + ((!g2129) & (g2177) & (!g2776) & (!g2807) & (g2098) & (!g2708)) + ((!g2129) & (g2177) & (g2776) & (!g2807) & (!g2098) & (!g2708)) + ((!g2129) & (g2177) & (g2776) & (!g2807) & (!g2098) & (g2708)) + ((!g2129) & (g2177) & (g2776) & (!g2807) & (g2098) & (!g2708)) + ((g2129) & (!g2177) & (!g2776) & (!g2807) & (!g2098) & (!g2708)) + ((g2129) & (!g2177) & (!g2776) & (!g2807) & (!g2098) & (g2708)) + ((g2129) & (!g2177) & (!g2776) & (!g2807) & (g2098) & (!g2708)) + ((g2129) & (!g2177) & (!g2776) & (g2807) & (!g2098) & (!g2708)) + ((g2129) & (!g2177) & (!g2776) & (g2807) & (!g2098) & (g2708)) + ((g2129) & (!g2177) & (!g2776) & (g2807) & (g2098) & (!g2708)) + ((g2129) & (g2177) & (!g2776) & (!g2807) & (!g2098) & (!g2708)) + ((g2129) & (g2177) & (!g2776) & (!g2807) & (!g2098) & (g2708)) + ((g2129) & (g2177) & (!g2776) & (!g2807) & (g2098) & (!g2708)));
	assign g5780 = (((!g2098) & (!g2708)));
	assign g5781 = (((!g2764) & (!g2813) & (g2785) & (g2822) & (!g2838) & (g2871)) + ((!g2764) & (!g2813) & (g2785) & (g2822) & (g2838) & (!g2871)) + ((!g2764) & (g2813) & (!g2785) & (g2822) & (!g2838) & (g2871)) + ((!g2764) & (g2813) & (!g2785) & (g2822) & (g2838) & (!g2871)) + ((!g2764) & (g2813) & (g2785) & (!g2822) & (!g2838) & (g2871)) + ((!g2764) & (g2813) & (g2785) & (!g2822) & (g2838) & (!g2871)) + ((!g2764) & (g2813) & (g2785) & (g2822) & (!g2838) & (g2871)) + ((!g2764) & (g2813) & (g2785) & (g2822) & (g2838) & (!g2871)) + ((g2764) & (!g2813) & (!g2785) & (g2822) & (!g2838) & (g2871)) + ((g2764) & (!g2813) & (!g2785) & (g2822) & (g2838) & (!g2871)) + ((g2764) & (!g2813) & (g2785) & (g2822) & (!g2838) & (g2871)) + ((g2764) & (!g2813) & (g2785) & (g2822) & (g2838) & (!g2871)) + ((g2764) & (g2813) & (!g2785) & (!g2822) & (!g2838) & (g2871)) + ((g2764) & (g2813) & (!g2785) & (!g2822) & (g2838) & (!g2871)) + ((g2764) & (g2813) & (!g2785) & (g2822) & (!g2838) & (g2871)) + ((g2764) & (g2813) & (!g2785) & (g2822) & (g2838) & (!g2871)) + ((g2764) & (g2813) & (g2785) & (!g2822) & (!g2838) & (g2871)) + ((g2764) & (g2813) & (g2785) & (!g2822) & (g2838) & (!g2871)) + ((g2764) & (g2813) & (g2785) & (g2822) & (!g2838) & (g2871)) + ((g2764) & (g2813) & (g2785) & (g2822) & (g2838) & (!g2871)));
	assign g5782 = (((!g2764) & (!g2813) & (!g2785) & (!g2822) & (!g2718) & (!g2733)) + ((!g2764) & (!g2813) & (!g2785) & (!g2822) & (!g2718) & (g2733)) + ((!g2764) & (!g2813) & (!g2785) & (!g2822) & (g2718) & (!g2733)) + ((!g2764) & (!g2813) & (!g2785) & (g2822) & (!g2718) & (!g2733)) + ((!g2764) & (!g2813) & (!g2785) & (g2822) & (!g2718) & (g2733)) + ((!g2764) & (!g2813) & (!g2785) & (g2822) & (g2718) & (!g2733)) + ((!g2764) & (!g2813) & (g2785) & (!g2822) & (!g2718) & (!g2733)) + ((!g2764) & (!g2813) & (g2785) & (!g2822) & (!g2718) & (g2733)) + ((!g2764) & (!g2813) & (g2785) & (!g2822) & (g2718) & (!g2733)) + ((!g2764) & (!g2813) & (g2785) & (g2822) & (!g2718) & (!g2733)) + ((!g2764) & (!g2813) & (g2785) & (g2822) & (!g2718) & (g2733)) + ((!g2764) & (!g2813) & (g2785) & (g2822) & (g2718) & (!g2733)) + ((!g2764) & (g2813) & (!g2785) & (!g2822) & (!g2718) & (!g2733)) + ((!g2764) & (g2813) & (!g2785) & (!g2822) & (!g2718) & (g2733)) + ((!g2764) & (g2813) & (!g2785) & (!g2822) & (g2718) & (!g2733)) + ((!g2764) & (g2813) & (g2785) & (!g2822) & (!g2718) & (!g2733)) + ((!g2764) & (g2813) & (g2785) & (!g2822) & (!g2718) & (g2733)) + ((!g2764) & (g2813) & (g2785) & (!g2822) & (g2718) & (!g2733)) + ((g2764) & (!g2813) & (!g2785) & (!g2822) & (!g2718) & (!g2733)) + ((g2764) & (!g2813) & (!g2785) & (!g2822) & (!g2718) & (g2733)) + ((g2764) & (!g2813) & (!g2785) & (!g2822) & (g2718) & (!g2733)) + ((g2764) & (!g2813) & (!g2785) & (g2822) & (!g2718) & (!g2733)) + ((g2764) & (!g2813) & (!g2785) & (g2822) & (!g2718) & (g2733)) + ((g2764) & (!g2813) & (!g2785) & (g2822) & (g2718) & (!g2733)) + ((g2764) & (g2813) & (!g2785) & (!g2822) & (!g2718) & (!g2733)) + ((g2764) & (g2813) & (!g2785) & (!g2822) & (!g2718) & (g2733)) + ((g2764) & (g2813) & (!g2785) & (!g2822) & (g2718) & (!g2733)));
	assign g5783 = (((!g2718) & (!g2733)));
	assign g5784 = (((!g2772) & (!g2827) & (g2780) & (g2830) & (!g2851) & (g2863)) + ((!g2772) & (!g2827) & (g2780) & (g2830) & (g2851) & (!g2863)) + ((!g2772) & (g2827) & (!g2780) & (g2830) & (!g2851) & (g2863)) + ((!g2772) & (g2827) & (!g2780) & (g2830) & (g2851) & (!g2863)) + ((!g2772) & (g2827) & (g2780) & (!g2830) & (!g2851) & (g2863)) + ((!g2772) & (g2827) & (g2780) & (!g2830) & (g2851) & (!g2863)) + ((!g2772) & (g2827) & (g2780) & (g2830) & (!g2851) & (g2863)) + ((!g2772) & (g2827) & (g2780) & (g2830) & (g2851) & (!g2863)) + ((g2772) & (!g2827) & (!g2780) & (g2830) & (!g2851) & (g2863)) + ((g2772) & (!g2827) & (!g2780) & (g2830) & (g2851) & (!g2863)) + ((g2772) & (!g2827) & (g2780) & (g2830) & (!g2851) & (g2863)) + ((g2772) & (!g2827) & (g2780) & (g2830) & (g2851) & (!g2863)) + ((g2772) & (g2827) & (!g2780) & (!g2830) & (!g2851) & (g2863)) + ((g2772) & (g2827) & (!g2780) & (!g2830) & (g2851) & (!g2863)) + ((g2772) & (g2827) & (!g2780) & (g2830) & (!g2851) & (g2863)) + ((g2772) & (g2827) & (!g2780) & (g2830) & (g2851) & (!g2863)) + ((g2772) & (g2827) & (g2780) & (!g2830) & (!g2851) & (g2863)) + ((g2772) & (g2827) & (g2780) & (!g2830) & (g2851) & (!g2863)) + ((g2772) & (g2827) & (g2780) & (g2830) & (!g2851) & (g2863)) + ((g2772) & (g2827) & (g2780) & (g2830) & (g2851) & (!g2863)));
	assign g5785 = (((!g2772) & (!g2827) & (!g2780) & (!g2830) & (!g2742) & (!g2747)) + ((!g2772) & (!g2827) & (!g2780) & (!g2830) & (!g2742) & (g2747)) + ((!g2772) & (!g2827) & (!g2780) & (!g2830) & (g2742) & (!g2747)) + ((!g2772) & (!g2827) & (!g2780) & (g2830) & (!g2742) & (!g2747)) + ((!g2772) & (!g2827) & (!g2780) & (g2830) & (!g2742) & (g2747)) + ((!g2772) & (!g2827) & (!g2780) & (g2830) & (g2742) & (!g2747)) + ((!g2772) & (!g2827) & (g2780) & (!g2830) & (!g2742) & (!g2747)) + ((!g2772) & (!g2827) & (g2780) & (!g2830) & (!g2742) & (g2747)) + ((!g2772) & (!g2827) & (g2780) & (!g2830) & (g2742) & (!g2747)) + ((!g2772) & (!g2827) & (g2780) & (g2830) & (!g2742) & (!g2747)) + ((!g2772) & (!g2827) & (g2780) & (g2830) & (!g2742) & (g2747)) + ((!g2772) & (!g2827) & (g2780) & (g2830) & (g2742) & (!g2747)) + ((!g2772) & (g2827) & (!g2780) & (!g2830) & (!g2742) & (!g2747)) + ((!g2772) & (g2827) & (!g2780) & (!g2830) & (!g2742) & (g2747)) + ((!g2772) & (g2827) & (!g2780) & (!g2830) & (g2742) & (!g2747)) + ((!g2772) & (g2827) & (g2780) & (!g2830) & (!g2742) & (!g2747)) + ((!g2772) & (g2827) & (g2780) & (!g2830) & (!g2742) & (g2747)) + ((!g2772) & (g2827) & (g2780) & (!g2830) & (g2742) & (!g2747)) + ((g2772) & (!g2827) & (!g2780) & (!g2830) & (!g2742) & (!g2747)) + ((g2772) & (!g2827) & (!g2780) & (!g2830) & (!g2742) & (g2747)) + ((g2772) & (!g2827) & (!g2780) & (!g2830) & (g2742) & (!g2747)) + ((g2772) & (!g2827) & (!g2780) & (g2830) & (!g2742) & (!g2747)) + ((g2772) & (!g2827) & (!g2780) & (g2830) & (!g2742) & (g2747)) + ((g2772) & (!g2827) & (!g2780) & (g2830) & (g2742) & (!g2747)) + ((g2772) & (g2827) & (!g2780) & (!g2830) & (!g2742) & (!g2747)) + ((g2772) & (g2827) & (!g2780) & (!g2830) & (!g2742) & (g2747)) + ((g2772) & (g2827) & (!g2780) & (!g2830) & (g2742) & (!g2747)));
	assign g5786 = (((!g2742) & (!g2747)));
	assign g5787 = (((!g2304) & (!g2360) & (g2326) & (g2364) & (!g2383) & (g2405)) + ((!g2304) & (!g2360) & (g2326) & (g2364) & (g2383) & (!g2405)) + ((!g2304) & (g2360) & (!g2326) & (g2364) & (!g2383) & (g2405)) + ((!g2304) & (g2360) & (!g2326) & (g2364) & (g2383) & (!g2405)) + ((!g2304) & (g2360) & (g2326) & (!g2364) & (!g2383) & (g2405)) + ((!g2304) & (g2360) & (g2326) & (!g2364) & (g2383) & (!g2405)) + ((!g2304) & (g2360) & (g2326) & (g2364) & (!g2383) & (g2405)) + ((!g2304) & (g2360) & (g2326) & (g2364) & (g2383) & (!g2405)) + ((g2304) & (!g2360) & (!g2326) & (g2364) & (!g2383) & (g2405)) + ((g2304) & (!g2360) & (!g2326) & (g2364) & (g2383) & (!g2405)) + ((g2304) & (!g2360) & (g2326) & (g2364) & (!g2383) & (g2405)) + ((g2304) & (!g2360) & (g2326) & (g2364) & (g2383) & (!g2405)) + ((g2304) & (g2360) & (!g2326) & (!g2364) & (!g2383) & (g2405)) + ((g2304) & (g2360) & (!g2326) & (!g2364) & (g2383) & (!g2405)) + ((g2304) & (g2360) & (!g2326) & (g2364) & (!g2383) & (g2405)) + ((g2304) & (g2360) & (!g2326) & (g2364) & (g2383) & (!g2405)) + ((g2304) & (g2360) & (g2326) & (!g2364) & (!g2383) & (g2405)) + ((g2304) & (g2360) & (g2326) & (!g2364) & (g2383) & (!g2405)) + ((g2304) & (g2360) & (g2326) & (g2364) & (!g2383) & (g2405)) + ((g2304) & (g2360) & (g2326) & (g2364) & (g2383) & (!g2405)));
	assign g5788 = (((!g2304) & (!g2360) & (!g2326) & (!g2364) & (!g2277) & (!g2281)) + ((!g2304) & (!g2360) & (!g2326) & (!g2364) & (!g2277) & (g2281)) + ((!g2304) & (!g2360) & (!g2326) & (!g2364) & (g2277) & (!g2281)) + ((!g2304) & (!g2360) & (!g2326) & (g2364) & (!g2277) & (!g2281)) + ((!g2304) & (!g2360) & (!g2326) & (g2364) & (!g2277) & (g2281)) + ((!g2304) & (!g2360) & (!g2326) & (g2364) & (g2277) & (!g2281)) + ((!g2304) & (!g2360) & (g2326) & (!g2364) & (!g2277) & (!g2281)) + ((!g2304) & (!g2360) & (g2326) & (!g2364) & (!g2277) & (g2281)) + ((!g2304) & (!g2360) & (g2326) & (!g2364) & (g2277) & (!g2281)) + ((!g2304) & (!g2360) & (g2326) & (g2364) & (!g2277) & (!g2281)) + ((!g2304) & (!g2360) & (g2326) & (g2364) & (!g2277) & (g2281)) + ((!g2304) & (!g2360) & (g2326) & (g2364) & (g2277) & (!g2281)) + ((!g2304) & (g2360) & (!g2326) & (!g2364) & (!g2277) & (!g2281)) + ((!g2304) & (g2360) & (!g2326) & (!g2364) & (!g2277) & (g2281)) + ((!g2304) & (g2360) & (!g2326) & (!g2364) & (g2277) & (!g2281)) + ((!g2304) & (g2360) & (g2326) & (!g2364) & (!g2277) & (!g2281)) + ((!g2304) & (g2360) & (g2326) & (!g2364) & (!g2277) & (g2281)) + ((!g2304) & (g2360) & (g2326) & (!g2364) & (g2277) & (!g2281)) + ((g2304) & (!g2360) & (!g2326) & (!g2364) & (!g2277) & (!g2281)) + ((g2304) & (!g2360) & (!g2326) & (!g2364) & (!g2277) & (g2281)) + ((g2304) & (!g2360) & (!g2326) & (!g2364) & (g2277) & (!g2281)) + ((g2304) & (!g2360) & (!g2326) & (g2364) & (!g2277) & (!g2281)) + ((g2304) & (!g2360) & (!g2326) & (g2364) & (!g2277) & (g2281)) + ((g2304) & (!g2360) & (!g2326) & (g2364) & (g2277) & (!g2281)) + ((g2304) & (g2360) & (!g2326) & (!g2364) & (!g2277) & (!g2281)) + ((g2304) & (g2360) & (!g2326) & (!g2364) & (!g2277) & (g2281)) + ((g2304) & (g2360) & (!g2326) & (!g2364) & (g2277) & (!g2281)));
	assign g5789 = (((!g2277) & (!g2281) & (g5787) & (!g5788)) + ((!g2277) & (g2281) & (g5787) & (!g5788)) + ((!g2277) & (g2281) & (g5787) & (g5788)) + ((g2277) & (!g2281) & (g5787) & (!g5788)) + ((g2277) & (!g2281) & (g5787) & (g5788)) + ((g2277) & (g2281) & (g5787) & (!g5788)) + ((g2277) & (g2281) & (g5787) & (g5788)));
	assign g5790 = (((!g1098) & (!g1132) & (g2320) & (g2350) & (!g1165) & (g2399)) + ((!g1098) & (!g1132) & (g2320) & (g2350) & (g1165) & (!g2399)) + ((!g1098) & (g1132) & (!g2320) & (g2350) & (!g1165) & (g2399)) + ((!g1098) & (g1132) & (!g2320) & (g2350) & (g1165) & (!g2399)) + ((!g1098) & (g1132) & (g2320) & (!g2350) & (!g1165) & (g2399)) + ((!g1098) & (g1132) & (g2320) & (!g2350) & (g1165) & (!g2399)) + ((!g1098) & (g1132) & (g2320) & (g2350) & (!g1165) & (g2399)) + ((!g1098) & (g1132) & (g2320) & (g2350) & (g1165) & (!g2399)) + ((g1098) & (!g1132) & (!g2320) & (g2350) & (!g1165) & (g2399)) + ((g1098) & (!g1132) & (!g2320) & (g2350) & (g1165) & (!g2399)) + ((g1098) & (!g1132) & (g2320) & (g2350) & (!g1165) & (g2399)) + ((g1098) & (!g1132) & (g2320) & (g2350) & (g1165) & (!g2399)) + ((g1098) & (g1132) & (!g2320) & (!g2350) & (!g1165) & (g2399)) + ((g1098) & (g1132) & (!g2320) & (!g2350) & (g1165) & (!g2399)) + ((g1098) & (g1132) & (!g2320) & (g2350) & (!g1165) & (g2399)) + ((g1098) & (g1132) & (!g2320) & (g2350) & (g1165) & (!g2399)) + ((g1098) & (g1132) & (g2320) & (!g2350) & (!g1165) & (g2399)) + ((g1098) & (g1132) & (g2320) & (!g2350) & (g1165) & (!g2399)) + ((g1098) & (g1132) & (g2320) & (g2350) & (!g1165) & (g2399)) + ((g1098) & (g1132) & (g2320) & (g2350) & (g1165) & (!g2399)));
	assign g5791 = (((!g1098) & (!g1132) & (!g2320) & (!g2350) & (!g1065) & (!g2267)) + ((!g1098) & (!g1132) & (!g2320) & (!g2350) & (!g1065) & (g2267)) + ((!g1098) & (!g1132) & (!g2320) & (!g2350) & (g1065) & (!g2267)) + ((!g1098) & (!g1132) & (!g2320) & (g2350) & (!g1065) & (!g2267)) + ((!g1098) & (!g1132) & (!g2320) & (g2350) & (!g1065) & (g2267)) + ((!g1098) & (!g1132) & (!g2320) & (g2350) & (g1065) & (!g2267)) + ((!g1098) & (!g1132) & (g2320) & (!g2350) & (!g1065) & (!g2267)) + ((!g1098) & (!g1132) & (g2320) & (!g2350) & (!g1065) & (g2267)) + ((!g1098) & (!g1132) & (g2320) & (!g2350) & (g1065) & (!g2267)) + ((!g1098) & (!g1132) & (g2320) & (g2350) & (!g1065) & (!g2267)) + ((!g1098) & (!g1132) & (g2320) & (g2350) & (!g1065) & (g2267)) + ((!g1098) & (!g1132) & (g2320) & (g2350) & (g1065) & (!g2267)) + ((!g1098) & (g1132) & (!g2320) & (!g2350) & (!g1065) & (!g2267)) + ((!g1098) & (g1132) & (!g2320) & (!g2350) & (!g1065) & (g2267)) + ((!g1098) & (g1132) & (!g2320) & (!g2350) & (g1065) & (!g2267)) + ((!g1098) & (g1132) & (g2320) & (!g2350) & (!g1065) & (!g2267)) + ((!g1098) & (g1132) & (g2320) & (!g2350) & (!g1065) & (g2267)) + ((!g1098) & (g1132) & (g2320) & (!g2350) & (g1065) & (!g2267)) + ((g1098) & (!g1132) & (!g2320) & (!g2350) & (!g1065) & (!g2267)) + ((g1098) & (!g1132) & (!g2320) & (!g2350) & (!g1065) & (g2267)) + ((g1098) & (!g1132) & (!g2320) & (!g2350) & (g1065) & (!g2267)) + ((g1098) & (!g1132) & (!g2320) & (g2350) & (!g1065) & (!g2267)) + ((g1098) & (!g1132) & (!g2320) & (g2350) & (!g1065) & (g2267)) + ((g1098) & (!g1132) & (!g2320) & (g2350) & (g1065) & (!g2267)) + ((g1098) & (g1132) & (!g2320) & (!g2350) & (!g1065) & (!g2267)) + ((g1098) & (g1132) & (!g2320) & (!g2350) & (!g1065) & (g2267)) + ((g1098) & (g1132) & (!g2320) & (!g2350) & (g1065) & (!g2267)));
	assign g5792 = (((!g1065) & (!g2267) & (g5790) & (!g5791)) + ((!g1065) & (g2267) & (g5790) & (!g5791)) + ((!g1065) & (g2267) & (g5790) & (g5791)) + ((g1065) & (!g2267) & (g5790) & (!g5791)) + ((g1065) & (!g2267) & (g5790) & (g5791)) + ((g1065) & (g2267) & (g5790) & (!g5791)) + ((g1065) & (g2267) & (g5790) & (g5791)));
	assign g5793 = (((!g1098) & (!g1132) & (g2304) & (g2360) & (!g1165) & (g2383)) + ((!g1098) & (!g1132) & (g2304) & (g2360) & (g1165) & (!g2383)) + ((!g1098) & (g1132) & (!g2304) & (g2360) & (!g1165) & (g2383)) + ((!g1098) & (g1132) & (!g2304) & (g2360) & (g1165) & (!g2383)) + ((!g1098) & (g1132) & (g2304) & (!g2360) & (!g1165) & (g2383)) + ((!g1098) & (g1132) & (g2304) & (!g2360) & (g1165) & (!g2383)) + ((!g1098) & (g1132) & (g2304) & (g2360) & (!g1165) & (g2383)) + ((!g1098) & (g1132) & (g2304) & (g2360) & (g1165) & (!g2383)) + ((g1098) & (!g1132) & (!g2304) & (g2360) & (!g1165) & (g2383)) + ((g1098) & (!g1132) & (!g2304) & (g2360) & (g1165) & (!g2383)) + ((g1098) & (!g1132) & (g2304) & (g2360) & (!g1165) & (g2383)) + ((g1098) & (!g1132) & (g2304) & (g2360) & (g1165) & (!g2383)) + ((g1098) & (g1132) & (!g2304) & (!g2360) & (!g1165) & (g2383)) + ((g1098) & (g1132) & (!g2304) & (!g2360) & (g1165) & (!g2383)) + ((g1098) & (g1132) & (!g2304) & (g2360) & (!g1165) & (g2383)) + ((g1098) & (g1132) & (!g2304) & (g2360) & (g1165) & (!g2383)) + ((g1098) & (g1132) & (g2304) & (!g2360) & (!g1165) & (g2383)) + ((g1098) & (g1132) & (g2304) & (!g2360) & (g1165) & (!g2383)) + ((g1098) & (g1132) & (g2304) & (g2360) & (!g1165) & (g2383)) + ((g1098) & (g1132) & (g2304) & (g2360) & (g1165) & (!g2383)));
	assign g5794 = (((!g1098) & (!g1132) & (!g2304) & (!g2360) & (!g1065) & (!g2277)) + ((!g1098) & (!g1132) & (!g2304) & (!g2360) & (!g1065) & (g2277)) + ((!g1098) & (!g1132) & (!g2304) & (!g2360) & (g1065) & (!g2277)) + ((!g1098) & (!g1132) & (!g2304) & (g2360) & (!g1065) & (!g2277)) + ((!g1098) & (!g1132) & (!g2304) & (g2360) & (!g1065) & (g2277)) + ((!g1098) & (!g1132) & (!g2304) & (g2360) & (g1065) & (!g2277)) + ((!g1098) & (!g1132) & (g2304) & (!g2360) & (!g1065) & (!g2277)) + ((!g1098) & (!g1132) & (g2304) & (!g2360) & (!g1065) & (g2277)) + ((!g1098) & (!g1132) & (g2304) & (!g2360) & (g1065) & (!g2277)) + ((!g1098) & (!g1132) & (g2304) & (g2360) & (!g1065) & (!g2277)) + ((!g1098) & (!g1132) & (g2304) & (g2360) & (!g1065) & (g2277)) + ((!g1098) & (!g1132) & (g2304) & (g2360) & (g1065) & (!g2277)) + ((!g1098) & (g1132) & (!g2304) & (!g2360) & (!g1065) & (!g2277)) + ((!g1098) & (g1132) & (!g2304) & (!g2360) & (!g1065) & (g2277)) + ((!g1098) & (g1132) & (!g2304) & (!g2360) & (g1065) & (!g2277)) + ((!g1098) & (g1132) & (g2304) & (!g2360) & (!g1065) & (!g2277)) + ((!g1098) & (g1132) & (g2304) & (!g2360) & (!g1065) & (g2277)) + ((!g1098) & (g1132) & (g2304) & (!g2360) & (g1065) & (!g2277)) + ((g1098) & (!g1132) & (!g2304) & (!g2360) & (!g1065) & (!g2277)) + ((g1098) & (!g1132) & (!g2304) & (!g2360) & (!g1065) & (g2277)) + ((g1098) & (!g1132) & (!g2304) & (!g2360) & (g1065) & (!g2277)) + ((g1098) & (!g1132) & (!g2304) & (g2360) & (!g1065) & (!g2277)) + ((g1098) & (!g1132) & (!g2304) & (g2360) & (!g1065) & (g2277)) + ((g1098) & (!g1132) & (!g2304) & (g2360) & (g1065) & (!g2277)) + ((g1098) & (g1132) & (!g2304) & (!g2360) & (!g1065) & (!g2277)) + ((g1098) & (g1132) & (!g2304) & (!g2360) & (!g1065) & (g2277)) + ((g1098) & (g1132) & (!g2304) & (!g2360) & (g1065) & (!g2277)));
	assign g5795 = (((!g1065) & (!g2277) & (g5793) & (!g5794)) + ((!g1065) & (g2277) & (g5793) & (!g5794)) + ((!g1065) & (g2277) & (g5793) & (g5794)) + ((g1065) & (!g2277) & (g5793) & (!g5794)) + ((g1065) & (!g2277) & (g5793) & (g5794)) + ((g1065) & (g2277) & (g5793) & (!g5794)) + ((g1065) & (g2277) & (g5793) & (g5794)));
	assign g5796 = (((!g2012) & (!g2014) & (g1269) & (g1303) & (!g2052) & (g1337)) + ((!g2012) & (!g2014) & (g1269) & (g1303) & (g2052) & (!g1337)) + ((!g2012) & (g2014) & (!g1269) & (g1303) & (!g2052) & (g1337)) + ((!g2012) & (g2014) & (!g1269) & (g1303) & (g2052) & (!g1337)) + ((!g2012) & (g2014) & (g1269) & (!g1303) & (!g2052) & (g1337)) + ((!g2012) & (g2014) & (g1269) & (!g1303) & (g2052) & (!g1337)) + ((!g2012) & (g2014) & (g1269) & (g1303) & (!g2052) & (g1337)) + ((!g2012) & (g2014) & (g1269) & (g1303) & (g2052) & (!g1337)) + ((g2012) & (!g2014) & (!g1269) & (g1303) & (!g2052) & (g1337)) + ((g2012) & (!g2014) & (!g1269) & (g1303) & (g2052) & (!g1337)) + ((g2012) & (!g2014) & (g1269) & (g1303) & (!g2052) & (g1337)) + ((g2012) & (!g2014) & (g1269) & (g1303) & (g2052) & (!g1337)) + ((g2012) & (g2014) & (!g1269) & (!g1303) & (!g2052) & (g1337)) + ((g2012) & (g2014) & (!g1269) & (!g1303) & (g2052) & (!g1337)) + ((g2012) & (g2014) & (!g1269) & (g1303) & (!g2052) & (g1337)) + ((g2012) & (g2014) & (!g1269) & (g1303) & (g2052) & (!g1337)) + ((g2012) & (g2014) & (g1269) & (!g1303) & (!g2052) & (g1337)) + ((g2012) & (g2014) & (g1269) & (!g1303) & (g2052) & (!g1337)) + ((g2012) & (g2014) & (g1269) & (g1303) & (!g2052) & (g1337)) + ((g2012) & (g2014) & (g1269) & (g1303) & (g2052) & (!g1337)));
	assign g5797 = (((!g2012) & (!g2014) & (!g1269) & (!g1303) & (!g2006) & (!g1236)) + ((!g2012) & (!g2014) & (!g1269) & (!g1303) & (!g2006) & (g1236)) + ((!g2012) & (!g2014) & (!g1269) & (!g1303) & (g2006) & (!g1236)) + ((!g2012) & (!g2014) & (!g1269) & (g1303) & (!g2006) & (!g1236)) + ((!g2012) & (!g2014) & (!g1269) & (g1303) & (!g2006) & (g1236)) + ((!g2012) & (!g2014) & (!g1269) & (g1303) & (g2006) & (!g1236)) + ((!g2012) & (!g2014) & (g1269) & (!g1303) & (!g2006) & (!g1236)) + ((!g2012) & (!g2014) & (g1269) & (!g1303) & (!g2006) & (g1236)) + ((!g2012) & (!g2014) & (g1269) & (!g1303) & (g2006) & (!g1236)) + ((!g2012) & (!g2014) & (g1269) & (g1303) & (!g2006) & (!g1236)) + ((!g2012) & (!g2014) & (g1269) & (g1303) & (!g2006) & (g1236)) + ((!g2012) & (!g2014) & (g1269) & (g1303) & (g2006) & (!g1236)) + ((!g2012) & (g2014) & (!g1269) & (!g1303) & (!g2006) & (!g1236)) + ((!g2012) & (g2014) & (!g1269) & (!g1303) & (!g2006) & (g1236)) + ((!g2012) & (g2014) & (!g1269) & (!g1303) & (g2006) & (!g1236)) + ((!g2012) & (g2014) & (g1269) & (!g1303) & (!g2006) & (!g1236)) + ((!g2012) & (g2014) & (g1269) & (!g1303) & (!g2006) & (g1236)) + ((!g2012) & (g2014) & (g1269) & (!g1303) & (g2006) & (!g1236)) + ((g2012) & (!g2014) & (!g1269) & (!g1303) & (!g2006) & (!g1236)) + ((g2012) & (!g2014) & (!g1269) & (!g1303) & (!g2006) & (g1236)) + ((g2012) & (!g2014) & (!g1269) & (!g1303) & (g2006) & (!g1236)) + ((g2012) & (!g2014) & (!g1269) & (g1303) & (!g2006) & (!g1236)) + ((g2012) & (!g2014) & (!g1269) & (g1303) & (!g2006) & (g1236)) + ((g2012) & (!g2014) & (!g1269) & (g1303) & (g2006) & (!g1236)) + ((g2012) & (g2014) & (!g1269) & (!g1303) & (!g2006) & (!g1236)) + ((g2012) & (g2014) & (!g1269) & (!g1303) & (!g2006) & (g1236)) + ((g2012) & (g2014) & (!g1269) & (!g1303) & (g2006) & (!g1236)));
	assign g5798 = (((!g2006) & (!g1236) & (g5796) & (!g5797)) + ((!g2006) & (g1236) & (g5796) & (!g5797)) + ((!g2006) & (g1236) & (g5796) & (g5797)) + ((g2006) & (!g1236) & (g5796) & (!g5797)) + ((g2006) & (!g1236) & (g5796) & (g5797)) + ((g2006) & (g1236) & (g5796) & (!g5797)) + ((g2006) & (g1236) & (g5796) & (g5797)));
	assign g5799 = (((!g2566) & (!g2614) & (g2578) & (g2617) & (!g2657) & (g2665)) + ((!g2566) & (!g2614) & (g2578) & (g2617) & (g2657) & (!g2665)) + ((!g2566) & (g2614) & (!g2578) & (g2617) & (!g2657) & (g2665)) + ((!g2566) & (g2614) & (!g2578) & (g2617) & (g2657) & (!g2665)) + ((!g2566) & (g2614) & (g2578) & (!g2617) & (!g2657) & (g2665)) + ((!g2566) & (g2614) & (g2578) & (!g2617) & (g2657) & (!g2665)) + ((!g2566) & (g2614) & (g2578) & (g2617) & (!g2657) & (g2665)) + ((!g2566) & (g2614) & (g2578) & (g2617) & (g2657) & (!g2665)) + ((g2566) & (!g2614) & (!g2578) & (g2617) & (!g2657) & (g2665)) + ((g2566) & (!g2614) & (!g2578) & (g2617) & (g2657) & (!g2665)) + ((g2566) & (!g2614) & (g2578) & (g2617) & (!g2657) & (g2665)) + ((g2566) & (!g2614) & (g2578) & (g2617) & (g2657) & (!g2665)) + ((g2566) & (g2614) & (!g2578) & (!g2617) & (!g2657) & (g2665)) + ((g2566) & (g2614) & (!g2578) & (!g2617) & (g2657) & (!g2665)) + ((g2566) & (g2614) & (!g2578) & (g2617) & (!g2657) & (g2665)) + ((g2566) & (g2614) & (!g2578) & (g2617) & (g2657) & (!g2665)) + ((g2566) & (g2614) & (g2578) & (!g2617) & (!g2657) & (g2665)) + ((g2566) & (g2614) & (g2578) & (!g2617) & (g2657) & (!g2665)) + ((g2566) & (g2614) & (g2578) & (g2617) & (!g2657) & (g2665)) + ((g2566) & (g2614) & (g2578) & (g2617) & (g2657) & (!g2665)));
	assign g5800 = (((!g2566) & (!g2614) & (!g2578) & (!g2617) & (!g2527) & (!g2529)) + ((!g2566) & (!g2614) & (!g2578) & (!g2617) & (!g2527) & (g2529)) + ((!g2566) & (!g2614) & (!g2578) & (!g2617) & (g2527) & (!g2529)) + ((!g2566) & (!g2614) & (!g2578) & (g2617) & (!g2527) & (!g2529)) + ((!g2566) & (!g2614) & (!g2578) & (g2617) & (!g2527) & (g2529)) + ((!g2566) & (!g2614) & (!g2578) & (g2617) & (g2527) & (!g2529)) + ((!g2566) & (!g2614) & (g2578) & (!g2617) & (!g2527) & (!g2529)) + ((!g2566) & (!g2614) & (g2578) & (!g2617) & (!g2527) & (g2529)) + ((!g2566) & (!g2614) & (g2578) & (!g2617) & (g2527) & (!g2529)) + ((!g2566) & (!g2614) & (g2578) & (g2617) & (!g2527) & (!g2529)) + ((!g2566) & (!g2614) & (g2578) & (g2617) & (!g2527) & (g2529)) + ((!g2566) & (!g2614) & (g2578) & (g2617) & (g2527) & (!g2529)) + ((!g2566) & (g2614) & (!g2578) & (!g2617) & (!g2527) & (!g2529)) + ((!g2566) & (g2614) & (!g2578) & (!g2617) & (!g2527) & (g2529)) + ((!g2566) & (g2614) & (!g2578) & (!g2617) & (g2527) & (!g2529)) + ((!g2566) & (g2614) & (g2578) & (!g2617) & (!g2527) & (!g2529)) + ((!g2566) & (g2614) & (g2578) & (!g2617) & (!g2527) & (g2529)) + ((!g2566) & (g2614) & (g2578) & (!g2617) & (g2527) & (!g2529)) + ((g2566) & (!g2614) & (!g2578) & (!g2617) & (!g2527) & (!g2529)) + ((g2566) & (!g2614) & (!g2578) & (!g2617) & (!g2527) & (g2529)) + ((g2566) & (!g2614) & (!g2578) & (!g2617) & (g2527) & (!g2529)) + ((g2566) & (!g2614) & (!g2578) & (g2617) & (!g2527) & (!g2529)) + ((g2566) & (!g2614) & (!g2578) & (g2617) & (!g2527) & (g2529)) + ((g2566) & (!g2614) & (!g2578) & (g2617) & (g2527) & (!g2529)) + ((g2566) & (g2614) & (!g2578) & (!g2617) & (!g2527) & (!g2529)) + ((g2566) & (g2614) & (!g2578) & (!g2617) & (!g2527) & (g2529)) + ((g2566) & (g2614) & (!g2578) & (!g2617) & (g2527) & (!g2529)));
	assign g5801 = (((!g2527) & (!g2529) & (g5799) & (!g5800)) + ((!g2527) & (g2529) & (g5799) & (!g5800)) + ((!g2527) & (g2529) & (g5799) & (g5800)) + ((g2527) & (!g2529) & (g5799) & (!g5800)) + ((g2527) & (!g2529) & (g5799) & (g5800)) + ((g2527) & (g2529) & (g5799) & (!g5800)) + ((g2527) & (g2529) & (g5799) & (g5800)));
	assign g5802 = (((!g1973) & (!g1976) & (g1269) & (g1303) & (!g2048) & (g1337)) + ((!g1973) & (!g1976) & (g1269) & (g1303) & (g2048) & (!g1337)) + ((!g1973) & (g1976) & (!g1269) & (g1303) & (!g2048) & (g1337)) + ((!g1973) & (g1976) & (!g1269) & (g1303) & (g2048) & (!g1337)) + ((!g1973) & (g1976) & (g1269) & (!g1303) & (!g2048) & (g1337)) + ((!g1973) & (g1976) & (g1269) & (!g1303) & (g2048) & (!g1337)) + ((!g1973) & (g1976) & (g1269) & (g1303) & (!g2048) & (g1337)) + ((!g1973) & (g1976) & (g1269) & (g1303) & (g2048) & (!g1337)) + ((g1973) & (!g1976) & (!g1269) & (g1303) & (!g2048) & (g1337)) + ((g1973) & (!g1976) & (!g1269) & (g1303) & (g2048) & (!g1337)) + ((g1973) & (!g1976) & (g1269) & (g1303) & (!g2048) & (g1337)) + ((g1973) & (!g1976) & (g1269) & (g1303) & (g2048) & (!g1337)) + ((g1973) & (g1976) & (!g1269) & (!g1303) & (!g2048) & (g1337)) + ((g1973) & (g1976) & (!g1269) & (!g1303) & (g2048) & (!g1337)) + ((g1973) & (g1976) & (!g1269) & (g1303) & (!g2048) & (g1337)) + ((g1973) & (g1976) & (!g1269) & (g1303) & (g2048) & (!g1337)) + ((g1973) & (g1976) & (g1269) & (!g1303) & (!g2048) & (g1337)) + ((g1973) & (g1976) & (g1269) & (!g1303) & (g2048) & (!g1337)) + ((g1973) & (g1976) & (g1269) & (g1303) & (!g2048) & (g1337)) + ((g1973) & (g1976) & (g1269) & (g1303) & (g2048) & (!g1337)));
	assign g5803 = (((!g1973) & (!g1976) & (!g1269) & (!g1303) & (!g1970) & (!g1236)) + ((!g1973) & (!g1976) & (!g1269) & (!g1303) & (!g1970) & (g1236)) + ((!g1973) & (!g1976) & (!g1269) & (!g1303) & (g1970) & (!g1236)) + ((!g1973) & (!g1976) & (!g1269) & (g1303) & (!g1970) & (!g1236)) + ((!g1973) & (!g1976) & (!g1269) & (g1303) & (!g1970) & (g1236)) + ((!g1973) & (!g1976) & (!g1269) & (g1303) & (g1970) & (!g1236)) + ((!g1973) & (!g1976) & (g1269) & (!g1303) & (!g1970) & (!g1236)) + ((!g1973) & (!g1976) & (g1269) & (!g1303) & (!g1970) & (g1236)) + ((!g1973) & (!g1976) & (g1269) & (!g1303) & (g1970) & (!g1236)) + ((!g1973) & (!g1976) & (g1269) & (g1303) & (!g1970) & (!g1236)) + ((!g1973) & (!g1976) & (g1269) & (g1303) & (!g1970) & (g1236)) + ((!g1973) & (!g1976) & (g1269) & (g1303) & (g1970) & (!g1236)) + ((!g1973) & (g1976) & (!g1269) & (!g1303) & (!g1970) & (!g1236)) + ((!g1973) & (g1976) & (!g1269) & (!g1303) & (!g1970) & (g1236)) + ((!g1973) & (g1976) & (!g1269) & (!g1303) & (g1970) & (!g1236)) + ((!g1973) & (g1976) & (g1269) & (!g1303) & (!g1970) & (!g1236)) + ((!g1973) & (g1976) & (g1269) & (!g1303) & (!g1970) & (g1236)) + ((!g1973) & (g1976) & (g1269) & (!g1303) & (g1970) & (!g1236)) + ((g1973) & (!g1976) & (!g1269) & (!g1303) & (!g1970) & (!g1236)) + ((g1973) & (!g1976) & (!g1269) & (!g1303) & (!g1970) & (g1236)) + ((g1973) & (!g1976) & (!g1269) & (!g1303) & (g1970) & (!g1236)) + ((g1973) & (!g1976) & (!g1269) & (g1303) & (!g1970) & (!g1236)) + ((g1973) & (!g1976) & (!g1269) & (g1303) & (!g1970) & (g1236)) + ((g1973) & (!g1976) & (!g1269) & (g1303) & (g1970) & (!g1236)) + ((g1973) & (g1976) & (!g1269) & (!g1303) & (!g1970) & (!g1236)) + ((g1973) & (g1976) & (!g1269) & (!g1303) & (!g1970) & (g1236)) + ((g1973) & (g1976) & (!g1269) & (!g1303) & (g1970) & (!g1236)));
	assign g5804 = (((!g1970) & (!g1236) & (g5802) & (!g5803)) + ((!g1970) & (g1236) & (g5802) & (!g5803)) + ((!g1970) & (g1236) & (g5802) & (g5803)) + ((g1970) & (!g1236) & (g5802) & (!g5803)) + ((g1970) & (!g1236) & (g5802) & (g5803)) + ((g1970) & (g1236) & (g5802) & (!g5803)) + ((g1970) & (g1236) & (g5802) & (g5803)));
	assign g5805 = (((!g2559) & (!g2623) & (g2581) & (g2629) & (!g2653) & (g2667)) + ((!g2559) & (!g2623) & (g2581) & (g2629) & (g2653) & (!g2667)) + ((!g2559) & (g2623) & (!g2581) & (g2629) & (!g2653) & (g2667)) + ((!g2559) & (g2623) & (!g2581) & (g2629) & (g2653) & (!g2667)) + ((!g2559) & (g2623) & (g2581) & (!g2629) & (!g2653) & (g2667)) + ((!g2559) & (g2623) & (g2581) & (!g2629) & (g2653) & (!g2667)) + ((!g2559) & (g2623) & (g2581) & (g2629) & (!g2653) & (g2667)) + ((!g2559) & (g2623) & (g2581) & (g2629) & (g2653) & (!g2667)) + ((g2559) & (!g2623) & (!g2581) & (g2629) & (!g2653) & (g2667)) + ((g2559) & (!g2623) & (!g2581) & (g2629) & (g2653) & (!g2667)) + ((g2559) & (!g2623) & (g2581) & (g2629) & (!g2653) & (g2667)) + ((g2559) & (!g2623) & (g2581) & (g2629) & (g2653) & (!g2667)) + ((g2559) & (g2623) & (!g2581) & (!g2629) & (!g2653) & (g2667)) + ((g2559) & (g2623) & (!g2581) & (!g2629) & (g2653) & (!g2667)) + ((g2559) & (g2623) & (!g2581) & (g2629) & (!g2653) & (g2667)) + ((g2559) & (g2623) & (!g2581) & (g2629) & (g2653) & (!g2667)) + ((g2559) & (g2623) & (g2581) & (!g2629) & (!g2653) & (g2667)) + ((g2559) & (g2623) & (g2581) & (!g2629) & (g2653) & (!g2667)) + ((g2559) & (g2623) & (g2581) & (g2629) & (!g2653) & (g2667)) + ((g2559) & (g2623) & (g2581) & (g2629) & (g2653) & (!g2667)));
	assign g5806 = (((!g2559) & (!g2623) & (!g2581) & (!g2629) & (!g2533) & (!g2537)) + ((!g2559) & (!g2623) & (!g2581) & (!g2629) & (!g2533) & (g2537)) + ((!g2559) & (!g2623) & (!g2581) & (!g2629) & (g2533) & (!g2537)) + ((!g2559) & (!g2623) & (!g2581) & (g2629) & (!g2533) & (!g2537)) + ((!g2559) & (!g2623) & (!g2581) & (g2629) & (!g2533) & (g2537)) + ((!g2559) & (!g2623) & (!g2581) & (g2629) & (g2533) & (!g2537)) + ((!g2559) & (!g2623) & (g2581) & (!g2629) & (!g2533) & (!g2537)) + ((!g2559) & (!g2623) & (g2581) & (!g2629) & (!g2533) & (g2537)) + ((!g2559) & (!g2623) & (g2581) & (!g2629) & (g2533) & (!g2537)) + ((!g2559) & (!g2623) & (g2581) & (g2629) & (!g2533) & (!g2537)) + ((!g2559) & (!g2623) & (g2581) & (g2629) & (!g2533) & (g2537)) + ((!g2559) & (!g2623) & (g2581) & (g2629) & (g2533) & (!g2537)) + ((!g2559) & (g2623) & (!g2581) & (!g2629) & (!g2533) & (!g2537)) + ((!g2559) & (g2623) & (!g2581) & (!g2629) & (!g2533) & (g2537)) + ((!g2559) & (g2623) & (!g2581) & (!g2629) & (g2533) & (!g2537)) + ((!g2559) & (g2623) & (g2581) & (!g2629) & (!g2533) & (!g2537)) + ((!g2559) & (g2623) & (g2581) & (!g2629) & (!g2533) & (g2537)) + ((!g2559) & (g2623) & (g2581) & (!g2629) & (g2533) & (!g2537)) + ((g2559) & (!g2623) & (!g2581) & (!g2629) & (!g2533) & (!g2537)) + ((g2559) & (!g2623) & (!g2581) & (!g2629) & (!g2533) & (g2537)) + ((g2559) & (!g2623) & (!g2581) & (!g2629) & (g2533) & (!g2537)) + ((g2559) & (!g2623) & (!g2581) & (g2629) & (!g2533) & (!g2537)) + ((g2559) & (!g2623) & (!g2581) & (g2629) & (!g2533) & (g2537)) + ((g2559) & (!g2623) & (!g2581) & (g2629) & (g2533) & (!g2537)) + ((g2559) & (g2623) & (!g2581) & (!g2629) & (!g2533) & (!g2537)) + ((g2559) & (g2623) & (!g2581) & (!g2629) & (!g2533) & (g2537)) + ((g2559) & (g2623) & (!g2581) & (!g2629) & (g2533) & (!g2537)));
	assign g5807 = (((!g2533) & (!g2537) & (g5805) & (!g5806)) + ((!g2533) & (g2537) & (g5805) & (!g5806)) + ((!g2533) & (g2537) & (g5805) & (g5806)) + ((g2533) & (!g2537) & (g5805) & (!g5806)) + ((g2533) & (!g2537) & (g5805) & (g5806)) + ((g2533) & (g2537) & (g5805) & (!g5806)) + ((g2533) & (g2537) & (g5805) & (g5806)));
	assign g5808 = (((!g2572) & (!g2637) & (g2595) & (g2643) & (!g2661) & (g2676)) + ((!g2572) & (!g2637) & (g2595) & (g2643) & (g2661) & (!g2676)) + ((!g2572) & (g2637) & (!g2595) & (g2643) & (!g2661) & (g2676)) + ((!g2572) & (g2637) & (!g2595) & (g2643) & (g2661) & (!g2676)) + ((!g2572) & (g2637) & (g2595) & (!g2643) & (!g2661) & (g2676)) + ((!g2572) & (g2637) & (g2595) & (!g2643) & (g2661) & (!g2676)) + ((!g2572) & (g2637) & (g2595) & (g2643) & (!g2661) & (g2676)) + ((!g2572) & (g2637) & (g2595) & (g2643) & (g2661) & (!g2676)) + ((g2572) & (!g2637) & (!g2595) & (g2643) & (!g2661) & (g2676)) + ((g2572) & (!g2637) & (!g2595) & (g2643) & (g2661) & (!g2676)) + ((g2572) & (!g2637) & (g2595) & (g2643) & (!g2661) & (g2676)) + ((g2572) & (!g2637) & (g2595) & (g2643) & (g2661) & (!g2676)) + ((g2572) & (g2637) & (!g2595) & (!g2643) & (!g2661) & (g2676)) + ((g2572) & (g2637) & (!g2595) & (!g2643) & (g2661) & (!g2676)) + ((g2572) & (g2637) & (!g2595) & (g2643) & (!g2661) & (g2676)) + ((g2572) & (g2637) & (!g2595) & (g2643) & (g2661) & (!g2676)) + ((g2572) & (g2637) & (g2595) & (!g2643) & (!g2661) & (g2676)) + ((g2572) & (g2637) & (g2595) & (!g2643) & (g2661) & (!g2676)) + ((g2572) & (g2637) & (g2595) & (g2643) & (!g2661) & (g2676)) + ((g2572) & (g2637) & (g2595) & (g2643) & (g2661) & (!g2676)));
	assign g5809 = (((!g2572) & (!g2637) & (!g2595) & (!g2643) & (!g2542) & (!g2546)) + ((!g2572) & (!g2637) & (!g2595) & (!g2643) & (!g2542) & (g2546)) + ((!g2572) & (!g2637) & (!g2595) & (!g2643) & (g2542) & (!g2546)) + ((!g2572) & (!g2637) & (!g2595) & (g2643) & (!g2542) & (!g2546)) + ((!g2572) & (!g2637) & (!g2595) & (g2643) & (!g2542) & (g2546)) + ((!g2572) & (!g2637) & (!g2595) & (g2643) & (g2542) & (!g2546)) + ((!g2572) & (!g2637) & (g2595) & (!g2643) & (!g2542) & (!g2546)) + ((!g2572) & (!g2637) & (g2595) & (!g2643) & (!g2542) & (g2546)) + ((!g2572) & (!g2637) & (g2595) & (!g2643) & (g2542) & (!g2546)) + ((!g2572) & (!g2637) & (g2595) & (g2643) & (!g2542) & (!g2546)) + ((!g2572) & (!g2637) & (g2595) & (g2643) & (!g2542) & (g2546)) + ((!g2572) & (!g2637) & (g2595) & (g2643) & (g2542) & (!g2546)) + ((!g2572) & (g2637) & (!g2595) & (!g2643) & (!g2542) & (!g2546)) + ((!g2572) & (g2637) & (!g2595) & (!g2643) & (!g2542) & (g2546)) + ((!g2572) & (g2637) & (!g2595) & (!g2643) & (g2542) & (!g2546)) + ((!g2572) & (g2637) & (g2595) & (!g2643) & (!g2542) & (!g2546)) + ((!g2572) & (g2637) & (g2595) & (!g2643) & (!g2542) & (g2546)) + ((!g2572) & (g2637) & (g2595) & (!g2643) & (g2542) & (!g2546)) + ((g2572) & (!g2637) & (!g2595) & (!g2643) & (!g2542) & (!g2546)) + ((g2572) & (!g2637) & (!g2595) & (!g2643) & (!g2542) & (g2546)) + ((g2572) & (!g2637) & (!g2595) & (!g2643) & (g2542) & (!g2546)) + ((g2572) & (!g2637) & (!g2595) & (g2643) & (!g2542) & (!g2546)) + ((g2572) & (!g2637) & (!g2595) & (g2643) & (!g2542) & (g2546)) + ((g2572) & (!g2637) & (!g2595) & (g2643) & (g2542) & (!g2546)) + ((g2572) & (g2637) & (!g2595) & (!g2643) & (!g2542) & (!g2546)) + ((g2572) & (g2637) & (!g2595) & (!g2643) & (!g2542) & (g2546)) + ((g2572) & (g2637) & (!g2595) & (!g2643) & (g2542) & (!g2546)));
	assign g5810 = (((!g2542) & (!g2546) & (g5808) & (!g5809)) + ((!g2542) & (g2546) & (g5808) & (!g5809)) + ((!g2542) & (g2546) & (g5808) & (g5809)) + ((g2542) & (!g2546) & (g5808) & (!g5809)) + ((g2542) & (!g2546) & (g5808) & (g5809)) + ((g2542) & (g2546) & (g5808) & (!g5809)) + ((g2542) & (g2546) & (g5808) & (g5809)));
	assign g5811 = (((!g2566) & (!g2614) & (g2569) & (g2626) & (!g2657) & (g2659)) + ((!g2566) & (!g2614) & (g2569) & (g2626) & (g2657) & (!g2659)) + ((!g2566) & (g2614) & (!g2569) & (g2626) & (!g2657) & (g2659)) + ((!g2566) & (g2614) & (!g2569) & (g2626) & (g2657) & (!g2659)) + ((!g2566) & (g2614) & (g2569) & (!g2626) & (!g2657) & (g2659)) + ((!g2566) & (g2614) & (g2569) & (!g2626) & (g2657) & (!g2659)) + ((!g2566) & (g2614) & (g2569) & (g2626) & (!g2657) & (g2659)) + ((!g2566) & (g2614) & (g2569) & (g2626) & (g2657) & (!g2659)) + ((g2566) & (!g2614) & (!g2569) & (g2626) & (!g2657) & (g2659)) + ((g2566) & (!g2614) & (!g2569) & (g2626) & (g2657) & (!g2659)) + ((g2566) & (!g2614) & (g2569) & (g2626) & (!g2657) & (g2659)) + ((g2566) & (!g2614) & (g2569) & (g2626) & (g2657) & (!g2659)) + ((g2566) & (g2614) & (!g2569) & (!g2626) & (!g2657) & (g2659)) + ((g2566) & (g2614) & (!g2569) & (!g2626) & (g2657) & (!g2659)) + ((g2566) & (g2614) & (!g2569) & (g2626) & (!g2657) & (g2659)) + ((g2566) & (g2614) & (!g2569) & (g2626) & (g2657) & (!g2659)) + ((g2566) & (g2614) & (g2569) & (!g2626) & (!g2657) & (g2659)) + ((g2566) & (g2614) & (g2569) & (!g2626) & (g2657) & (!g2659)) + ((g2566) & (g2614) & (g2569) & (g2626) & (!g2657) & (g2659)) + ((g2566) & (g2614) & (g2569) & (g2626) & (g2657) & (!g2659)));
	assign g5812 = (((!g2566) & (!g2614) & (!g2569) & (!g2626) & (!g2527) & (!g2535)) + ((!g2566) & (!g2614) & (!g2569) & (!g2626) & (!g2527) & (g2535)) + ((!g2566) & (!g2614) & (!g2569) & (!g2626) & (g2527) & (!g2535)) + ((!g2566) & (!g2614) & (!g2569) & (g2626) & (!g2527) & (!g2535)) + ((!g2566) & (!g2614) & (!g2569) & (g2626) & (!g2527) & (g2535)) + ((!g2566) & (!g2614) & (!g2569) & (g2626) & (g2527) & (!g2535)) + ((!g2566) & (!g2614) & (g2569) & (!g2626) & (!g2527) & (!g2535)) + ((!g2566) & (!g2614) & (g2569) & (!g2626) & (!g2527) & (g2535)) + ((!g2566) & (!g2614) & (g2569) & (!g2626) & (g2527) & (!g2535)) + ((!g2566) & (!g2614) & (g2569) & (g2626) & (!g2527) & (!g2535)) + ((!g2566) & (!g2614) & (g2569) & (g2626) & (!g2527) & (g2535)) + ((!g2566) & (!g2614) & (g2569) & (g2626) & (g2527) & (!g2535)) + ((!g2566) & (g2614) & (!g2569) & (!g2626) & (!g2527) & (!g2535)) + ((!g2566) & (g2614) & (!g2569) & (!g2626) & (!g2527) & (g2535)) + ((!g2566) & (g2614) & (!g2569) & (!g2626) & (g2527) & (!g2535)) + ((!g2566) & (g2614) & (g2569) & (!g2626) & (!g2527) & (!g2535)) + ((!g2566) & (g2614) & (g2569) & (!g2626) & (!g2527) & (g2535)) + ((!g2566) & (g2614) & (g2569) & (!g2626) & (g2527) & (!g2535)) + ((g2566) & (!g2614) & (!g2569) & (!g2626) & (!g2527) & (!g2535)) + ((g2566) & (!g2614) & (!g2569) & (!g2626) & (!g2527) & (g2535)) + ((g2566) & (!g2614) & (!g2569) & (!g2626) & (g2527) & (!g2535)) + ((g2566) & (!g2614) & (!g2569) & (g2626) & (!g2527) & (!g2535)) + ((g2566) & (!g2614) & (!g2569) & (g2626) & (!g2527) & (g2535)) + ((g2566) & (!g2614) & (!g2569) & (g2626) & (g2527) & (!g2535)) + ((g2566) & (g2614) & (!g2569) & (!g2626) & (!g2527) & (!g2535)) + ((g2566) & (g2614) & (!g2569) & (!g2626) & (!g2527) & (g2535)) + ((g2566) & (g2614) & (!g2569) & (!g2626) & (g2527) & (!g2535)));
	assign g5813 = (((!g2527) & (!g2535) & (g5811) & (!g5812)) + ((!g2527) & (g2535) & (g5811) & (!g5812)) + ((!g2527) & (g2535) & (g5811) & (g5812)) + ((g2527) & (!g2535) & (g5811) & (!g5812)) + ((g2527) & (!g2535) & (g5811) & (g5812)) + ((g2527) & (g2535) & (g5811) & (!g5812)) + ((g2527) & (g2535) & (g5811) & (g5812)));
	assign g5814 = (((!g2566) & (!g2614) & (g2589) & (g2620) & (!g2657) & (g2672)) + ((!g2566) & (!g2614) & (g2589) & (g2620) & (g2657) & (!g2672)) + ((!g2566) & (g2614) & (!g2589) & (g2620) & (!g2657) & (g2672)) + ((!g2566) & (g2614) & (!g2589) & (g2620) & (g2657) & (!g2672)) + ((!g2566) & (g2614) & (g2589) & (!g2620) & (!g2657) & (g2672)) + ((!g2566) & (g2614) & (g2589) & (!g2620) & (g2657) & (!g2672)) + ((!g2566) & (g2614) & (g2589) & (g2620) & (!g2657) & (g2672)) + ((!g2566) & (g2614) & (g2589) & (g2620) & (g2657) & (!g2672)) + ((g2566) & (!g2614) & (!g2589) & (g2620) & (!g2657) & (g2672)) + ((g2566) & (!g2614) & (!g2589) & (g2620) & (g2657) & (!g2672)) + ((g2566) & (!g2614) & (g2589) & (g2620) & (!g2657) & (g2672)) + ((g2566) & (!g2614) & (g2589) & (g2620) & (g2657) & (!g2672)) + ((g2566) & (g2614) & (!g2589) & (!g2620) & (!g2657) & (g2672)) + ((g2566) & (g2614) & (!g2589) & (!g2620) & (g2657) & (!g2672)) + ((g2566) & (g2614) & (!g2589) & (g2620) & (!g2657) & (g2672)) + ((g2566) & (g2614) & (!g2589) & (g2620) & (g2657) & (!g2672)) + ((g2566) & (g2614) & (g2589) & (!g2620) & (!g2657) & (g2672)) + ((g2566) & (g2614) & (g2589) & (!g2620) & (g2657) & (!g2672)) + ((g2566) & (g2614) & (g2589) & (g2620) & (!g2657) & (g2672)) + ((g2566) & (g2614) & (g2589) & (g2620) & (g2657) & (!g2672)));
	assign g5815 = (((!g2566) & (!g2614) & (!g2589) & (!g2620) & (!g2527) & (!g2531)) + ((!g2566) & (!g2614) & (!g2589) & (!g2620) & (!g2527) & (g2531)) + ((!g2566) & (!g2614) & (!g2589) & (!g2620) & (g2527) & (!g2531)) + ((!g2566) & (!g2614) & (!g2589) & (g2620) & (!g2527) & (!g2531)) + ((!g2566) & (!g2614) & (!g2589) & (g2620) & (!g2527) & (g2531)) + ((!g2566) & (!g2614) & (!g2589) & (g2620) & (g2527) & (!g2531)) + ((!g2566) & (!g2614) & (g2589) & (!g2620) & (!g2527) & (!g2531)) + ((!g2566) & (!g2614) & (g2589) & (!g2620) & (!g2527) & (g2531)) + ((!g2566) & (!g2614) & (g2589) & (!g2620) & (g2527) & (!g2531)) + ((!g2566) & (!g2614) & (g2589) & (g2620) & (!g2527) & (!g2531)) + ((!g2566) & (!g2614) & (g2589) & (g2620) & (!g2527) & (g2531)) + ((!g2566) & (!g2614) & (g2589) & (g2620) & (g2527) & (!g2531)) + ((!g2566) & (g2614) & (!g2589) & (!g2620) & (!g2527) & (!g2531)) + ((!g2566) & (g2614) & (!g2589) & (!g2620) & (!g2527) & (g2531)) + ((!g2566) & (g2614) & (!g2589) & (!g2620) & (g2527) & (!g2531)) + ((!g2566) & (g2614) & (g2589) & (!g2620) & (!g2527) & (!g2531)) + ((!g2566) & (g2614) & (g2589) & (!g2620) & (!g2527) & (g2531)) + ((!g2566) & (g2614) & (g2589) & (!g2620) & (g2527) & (!g2531)) + ((g2566) & (!g2614) & (!g2589) & (!g2620) & (!g2527) & (!g2531)) + ((g2566) & (!g2614) & (!g2589) & (!g2620) & (!g2527) & (g2531)) + ((g2566) & (!g2614) & (!g2589) & (!g2620) & (g2527) & (!g2531)) + ((g2566) & (!g2614) & (!g2589) & (g2620) & (!g2527) & (!g2531)) + ((g2566) & (!g2614) & (!g2589) & (g2620) & (!g2527) & (g2531)) + ((g2566) & (!g2614) & (!g2589) & (g2620) & (g2527) & (!g2531)) + ((g2566) & (g2614) & (!g2589) & (!g2620) & (!g2527) & (!g2531)) + ((g2566) & (g2614) & (!g2589) & (!g2620) & (!g2527) & (g2531)) + ((g2566) & (g2614) & (!g2589) & (!g2620) & (g2527) & (!g2531)));
	assign g5816 = (((!g2527) & (!g2531) & (g5814) & (!g5815)) + ((!g2527) & (g2531) & (g5814) & (!g5815)) + ((!g2527) & (g2531) & (g5814) & (g5815)) + ((g2527) & (!g2531) & (g5814) & (!g5815)) + ((g2527) & (!g2531) & (g5814) & (g5815)) + ((g2527) & (g2531) & (g5814) & (!g5815)) + ((g2527) & (g2531) & (g5814) & (g5815)));
	assign g5817 = (((!g2012) & (!g2014) & (g2595) & (g2643) & (!g2052) & (g2676)) + ((!g2012) & (!g2014) & (g2595) & (g2643) & (g2052) & (!g2676)) + ((!g2012) & (g2014) & (!g2595) & (g2643) & (!g2052) & (g2676)) + ((!g2012) & (g2014) & (!g2595) & (g2643) & (g2052) & (!g2676)) + ((!g2012) & (g2014) & (g2595) & (!g2643) & (!g2052) & (g2676)) + ((!g2012) & (g2014) & (g2595) & (!g2643) & (g2052) & (!g2676)) + ((!g2012) & (g2014) & (g2595) & (g2643) & (!g2052) & (g2676)) + ((!g2012) & (g2014) & (g2595) & (g2643) & (g2052) & (!g2676)) + ((g2012) & (!g2014) & (!g2595) & (g2643) & (!g2052) & (g2676)) + ((g2012) & (!g2014) & (!g2595) & (g2643) & (g2052) & (!g2676)) + ((g2012) & (!g2014) & (g2595) & (g2643) & (!g2052) & (g2676)) + ((g2012) & (!g2014) & (g2595) & (g2643) & (g2052) & (!g2676)) + ((g2012) & (g2014) & (!g2595) & (!g2643) & (!g2052) & (g2676)) + ((g2012) & (g2014) & (!g2595) & (!g2643) & (g2052) & (!g2676)) + ((g2012) & (g2014) & (!g2595) & (g2643) & (!g2052) & (g2676)) + ((g2012) & (g2014) & (!g2595) & (g2643) & (g2052) & (!g2676)) + ((g2012) & (g2014) & (g2595) & (!g2643) & (!g2052) & (g2676)) + ((g2012) & (g2014) & (g2595) & (!g2643) & (g2052) & (!g2676)) + ((g2012) & (g2014) & (g2595) & (g2643) & (!g2052) & (g2676)) + ((g2012) & (g2014) & (g2595) & (g2643) & (g2052) & (!g2676)));
	assign g5818 = (((!g2012) & (!g2014) & (!g2595) & (!g2643) & (!g2006) & (!g2546)) + ((!g2012) & (!g2014) & (!g2595) & (!g2643) & (!g2006) & (g2546)) + ((!g2012) & (!g2014) & (!g2595) & (!g2643) & (g2006) & (!g2546)) + ((!g2012) & (!g2014) & (!g2595) & (g2643) & (!g2006) & (!g2546)) + ((!g2012) & (!g2014) & (!g2595) & (g2643) & (!g2006) & (g2546)) + ((!g2012) & (!g2014) & (!g2595) & (g2643) & (g2006) & (!g2546)) + ((!g2012) & (!g2014) & (g2595) & (!g2643) & (!g2006) & (!g2546)) + ((!g2012) & (!g2014) & (g2595) & (!g2643) & (!g2006) & (g2546)) + ((!g2012) & (!g2014) & (g2595) & (!g2643) & (g2006) & (!g2546)) + ((!g2012) & (!g2014) & (g2595) & (g2643) & (!g2006) & (!g2546)) + ((!g2012) & (!g2014) & (g2595) & (g2643) & (!g2006) & (g2546)) + ((!g2012) & (!g2014) & (g2595) & (g2643) & (g2006) & (!g2546)) + ((!g2012) & (g2014) & (!g2595) & (!g2643) & (!g2006) & (!g2546)) + ((!g2012) & (g2014) & (!g2595) & (!g2643) & (!g2006) & (g2546)) + ((!g2012) & (g2014) & (!g2595) & (!g2643) & (g2006) & (!g2546)) + ((!g2012) & (g2014) & (g2595) & (!g2643) & (!g2006) & (!g2546)) + ((!g2012) & (g2014) & (g2595) & (!g2643) & (!g2006) & (g2546)) + ((!g2012) & (g2014) & (g2595) & (!g2643) & (g2006) & (!g2546)) + ((g2012) & (!g2014) & (!g2595) & (!g2643) & (!g2006) & (!g2546)) + ((g2012) & (!g2014) & (!g2595) & (!g2643) & (!g2006) & (g2546)) + ((g2012) & (!g2014) & (!g2595) & (!g2643) & (g2006) & (!g2546)) + ((g2012) & (!g2014) & (!g2595) & (g2643) & (!g2006) & (!g2546)) + ((g2012) & (!g2014) & (!g2595) & (g2643) & (!g2006) & (g2546)) + ((g2012) & (!g2014) & (!g2595) & (g2643) & (g2006) & (!g2546)) + ((g2012) & (g2014) & (!g2595) & (!g2643) & (!g2006) & (!g2546)) + ((g2012) & (g2014) & (!g2595) & (!g2643) & (!g2006) & (g2546)) + ((g2012) & (g2014) & (!g2595) & (!g2643) & (g2006) & (!g2546)));
	assign g5819 = (((!g2006) & (!g2546) & (g5817) & (!g5818)) + ((!g2006) & (g2546) & (g5817) & (!g5818)) + ((!g2006) & (g2546) & (g5817) & (g5818)) + ((g2006) & (!g2546) & (g5817) & (!g5818)) + ((g2006) & (!g2546) & (g5817) & (g5818)) + ((g2006) & (g2546) & (g5817) & (!g5818)) + ((g2006) & (g2546) & (g5817) & (g5818)));
	assign g5820 = (((!g2569) & (!g2626) & (g2581) & (g2629) & (!g2667) & (g2659)) + ((!g2569) & (!g2626) & (g2581) & (g2629) & (g2667) & (!g2659)) + ((!g2569) & (g2626) & (!g2581) & (g2629) & (!g2667) & (g2659)) + ((!g2569) & (g2626) & (!g2581) & (g2629) & (g2667) & (!g2659)) + ((!g2569) & (g2626) & (g2581) & (!g2629) & (!g2667) & (g2659)) + ((!g2569) & (g2626) & (g2581) & (!g2629) & (g2667) & (!g2659)) + ((!g2569) & (g2626) & (g2581) & (g2629) & (!g2667) & (g2659)) + ((!g2569) & (g2626) & (g2581) & (g2629) & (g2667) & (!g2659)) + ((g2569) & (!g2626) & (!g2581) & (g2629) & (!g2667) & (g2659)) + ((g2569) & (!g2626) & (!g2581) & (g2629) & (g2667) & (!g2659)) + ((g2569) & (!g2626) & (g2581) & (g2629) & (!g2667) & (g2659)) + ((g2569) & (!g2626) & (g2581) & (g2629) & (g2667) & (!g2659)) + ((g2569) & (g2626) & (!g2581) & (!g2629) & (!g2667) & (g2659)) + ((g2569) & (g2626) & (!g2581) & (!g2629) & (g2667) & (!g2659)) + ((g2569) & (g2626) & (!g2581) & (g2629) & (!g2667) & (g2659)) + ((g2569) & (g2626) & (!g2581) & (g2629) & (g2667) & (!g2659)) + ((g2569) & (g2626) & (g2581) & (!g2629) & (!g2667) & (g2659)) + ((g2569) & (g2626) & (g2581) & (!g2629) & (g2667) & (!g2659)) + ((g2569) & (g2626) & (g2581) & (g2629) & (!g2667) & (g2659)) + ((g2569) & (g2626) & (g2581) & (g2629) & (g2667) & (!g2659)));
	assign g5821 = (((!g2569) & (!g2626) & (!g2581) & (!g2629) & (!g2535) & (!g2537)) + ((!g2569) & (!g2626) & (!g2581) & (!g2629) & (!g2535) & (g2537)) + ((!g2569) & (!g2626) & (!g2581) & (!g2629) & (g2535) & (!g2537)) + ((!g2569) & (!g2626) & (!g2581) & (g2629) & (!g2535) & (!g2537)) + ((!g2569) & (!g2626) & (!g2581) & (g2629) & (!g2535) & (g2537)) + ((!g2569) & (!g2626) & (!g2581) & (g2629) & (g2535) & (!g2537)) + ((!g2569) & (!g2626) & (g2581) & (!g2629) & (!g2535) & (!g2537)) + ((!g2569) & (!g2626) & (g2581) & (!g2629) & (!g2535) & (g2537)) + ((!g2569) & (!g2626) & (g2581) & (!g2629) & (g2535) & (!g2537)) + ((!g2569) & (!g2626) & (g2581) & (g2629) & (!g2535) & (!g2537)) + ((!g2569) & (!g2626) & (g2581) & (g2629) & (!g2535) & (g2537)) + ((!g2569) & (!g2626) & (g2581) & (g2629) & (g2535) & (!g2537)) + ((!g2569) & (g2626) & (!g2581) & (!g2629) & (!g2535) & (!g2537)) + ((!g2569) & (g2626) & (!g2581) & (!g2629) & (!g2535) & (g2537)) + ((!g2569) & (g2626) & (!g2581) & (!g2629) & (g2535) & (!g2537)) + ((!g2569) & (g2626) & (g2581) & (!g2629) & (!g2535) & (!g2537)) + ((!g2569) & (g2626) & (g2581) & (!g2629) & (!g2535) & (g2537)) + ((!g2569) & (g2626) & (g2581) & (!g2629) & (g2535) & (!g2537)) + ((g2569) & (!g2626) & (!g2581) & (!g2629) & (!g2535) & (!g2537)) + ((g2569) & (!g2626) & (!g2581) & (!g2629) & (!g2535) & (g2537)) + ((g2569) & (!g2626) & (!g2581) & (!g2629) & (g2535) & (!g2537)) + ((g2569) & (!g2626) & (!g2581) & (g2629) & (!g2535) & (!g2537)) + ((g2569) & (!g2626) & (!g2581) & (g2629) & (!g2535) & (g2537)) + ((g2569) & (!g2626) & (!g2581) & (g2629) & (g2535) & (!g2537)) + ((g2569) & (g2626) & (!g2581) & (!g2629) & (!g2535) & (!g2537)) + ((g2569) & (g2626) & (!g2581) & (!g2629) & (!g2535) & (g2537)) + ((g2569) & (g2626) & (!g2581) & (!g2629) & (g2535) & (!g2537)));
	assign g5822 = (((!g2535) & (!g2537) & (g5820) & (!g5821)) + ((!g2535) & (g2537) & (g5820) & (!g5821)) + ((!g2535) & (g2537) & (g5820) & (g5821)) + ((g2535) & (!g2537) & (g5820) & (!g5821)) + ((g2535) & (!g2537) & (g5820) & (g5821)) + ((g2535) & (g2537) & (g5820) & (!g5821)) + ((g2535) & (g2537) & (g5820) & (g5821)));
	assign g5823 = (((!g2578) & (!g2617) & (g2581) & (g2629) & (!g2665) & (g2667)) + ((!g2578) & (!g2617) & (g2581) & (g2629) & (g2665) & (!g2667)) + ((!g2578) & (g2617) & (!g2581) & (g2629) & (!g2665) & (g2667)) + ((!g2578) & (g2617) & (!g2581) & (g2629) & (g2665) & (!g2667)) + ((!g2578) & (g2617) & (g2581) & (!g2629) & (!g2665) & (g2667)) + ((!g2578) & (g2617) & (g2581) & (!g2629) & (g2665) & (!g2667)) + ((!g2578) & (g2617) & (g2581) & (g2629) & (!g2665) & (g2667)) + ((!g2578) & (g2617) & (g2581) & (g2629) & (g2665) & (!g2667)) + ((g2578) & (!g2617) & (!g2581) & (g2629) & (!g2665) & (g2667)) + ((g2578) & (!g2617) & (!g2581) & (g2629) & (g2665) & (!g2667)) + ((g2578) & (!g2617) & (g2581) & (g2629) & (!g2665) & (g2667)) + ((g2578) & (!g2617) & (g2581) & (g2629) & (g2665) & (!g2667)) + ((g2578) & (g2617) & (!g2581) & (!g2629) & (!g2665) & (g2667)) + ((g2578) & (g2617) & (!g2581) & (!g2629) & (g2665) & (!g2667)) + ((g2578) & (g2617) & (!g2581) & (g2629) & (!g2665) & (g2667)) + ((g2578) & (g2617) & (!g2581) & (g2629) & (g2665) & (!g2667)) + ((g2578) & (g2617) & (g2581) & (!g2629) & (!g2665) & (g2667)) + ((g2578) & (g2617) & (g2581) & (!g2629) & (g2665) & (!g2667)) + ((g2578) & (g2617) & (g2581) & (g2629) & (!g2665) & (g2667)) + ((g2578) & (g2617) & (g2581) & (g2629) & (g2665) & (!g2667)));
	assign g5824 = (((!g2578) & (!g2617) & (!g2581) & (!g2629) & (!g2529) & (!g2537)) + ((!g2578) & (!g2617) & (!g2581) & (!g2629) & (!g2529) & (g2537)) + ((!g2578) & (!g2617) & (!g2581) & (!g2629) & (g2529) & (!g2537)) + ((!g2578) & (!g2617) & (!g2581) & (g2629) & (!g2529) & (!g2537)) + ((!g2578) & (!g2617) & (!g2581) & (g2629) & (!g2529) & (g2537)) + ((!g2578) & (!g2617) & (!g2581) & (g2629) & (g2529) & (!g2537)) + ((!g2578) & (!g2617) & (g2581) & (!g2629) & (!g2529) & (!g2537)) + ((!g2578) & (!g2617) & (g2581) & (!g2629) & (!g2529) & (g2537)) + ((!g2578) & (!g2617) & (g2581) & (!g2629) & (g2529) & (!g2537)) + ((!g2578) & (!g2617) & (g2581) & (g2629) & (!g2529) & (!g2537)) + ((!g2578) & (!g2617) & (g2581) & (g2629) & (!g2529) & (g2537)) + ((!g2578) & (!g2617) & (g2581) & (g2629) & (g2529) & (!g2537)) + ((!g2578) & (g2617) & (!g2581) & (!g2629) & (!g2529) & (!g2537)) + ((!g2578) & (g2617) & (!g2581) & (!g2629) & (!g2529) & (g2537)) + ((!g2578) & (g2617) & (!g2581) & (!g2629) & (g2529) & (!g2537)) + ((!g2578) & (g2617) & (g2581) & (!g2629) & (!g2529) & (!g2537)) + ((!g2578) & (g2617) & (g2581) & (!g2629) & (!g2529) & (g2537)) + ((!g2578) & (g2617) & (g2581) & (!g2629) & (g2529) & (!g2537)) + ((g2578) & (!g2617) & (!g2581) & (!g2629) & (!g2529) & (!g2537)) + ((g2578) & (!g2617) & (!g2581) & (!g2629) & (!g2529) & (g2537)) + ((g2578) & (!g2617) & (!g2581) & (!g2629) & (g2529) & (!g2537)) + ((g2578) & (!g2617) & (!g2581) & (g2629) & (!g2529) & (!g2537)) + ((g2578) & (!g2617) & (!g2581) & (g2629) & (!g2529) & (g2537)) + ((g2578) & (!g2617) & (!g2581) & (g2629) & (g2529) & (!g2537)) + ((g2578) & (g2617) & (!g2581) & (!g2629) & (!g2529) & (!g2537)) + ((g2578) & (g2617) & (!g2581) & (!g2629) & (!g2529) & (g2537)) + ((g2578) & (g2617) & (!g2581) & (!g2629) & (g2529) & (!g2537)));
	assign g5825 = (((!g2529) & (!g2537) & (g5823) & (!g5824)) + ((!g2529) & (g2537) & (g5823) & (!g5824)) + ((!g2529) & (g2537) & (g5823) & (g5824)) + ((g2529) & (!g2537) & (g5823) & (!g5824)) + ((g2529) & (!g2537) & (g5823) & (g5824)) + ((g2529) & (g2537) & (g5823) & (!g5824)) + ((g2529) & (g2537) & (g5823) & (g5824)));
	assign g5826 = (((!g1973) & (!g1976) & (g2595) & (g2643) & (!g2048) & (g2676)) + ((!g1973) & (!g1976) & (g2595) & (g2643) & (g2048) & (!g2676)) + ((!g1973) & (g1976) & (!g2595) & (g2643) & (!g2048) & (g2676)) + ((!g1973) & (g1976) & (!g2595) & (g2643) & (g2048) & (!g2676)) + ((!g1973) & (g1976) & (g2595) & (!g2643) & (!g2048) & (g2676)) + ((!g1973) & (g1976) & (g2595) & (!g2643) & (g2048) & (!g2676)) + ((!g1973) & (g1976) & (g2595) & (g2643) & (!g2048) & (g2676)) + ((!g1973) & (g1976) & (g2595) & (g2643) & (g2048) & (!g2676)) + ((g1973) & (!g1976) & (!g2595) & (g2643) & (!g2048) & (g2676)) + ((g1973) & (!g1976) & (!g2595) & (g2643) & (g2048) & (!g2676)) + ((g1973) & (!g1976) & (g2595) & (g2643) & (!g2048) & (g2676)) + ((g1973) & (!g1976) & (g2595) & (g2643) & (g2048) & (!g2676)) + ((g1973) & (g1976) & (!g2595) & (!g2643) & (!g2048) & (g2676)) + ((g1973) & (g1976) & (!g2595) & (!g2643) & (g2048) & (!g2676)) + ((g1973) & (g1976) & (!g2595) & (g2643) & (!g2048) & (g2676)) + ((g1973) & (g1976) & (!g2595) & (g2643) & (g2048) & (!g2676)) + ((g1973) & (g1976) & (g2595) & (!g2643) & (!g2048) & (g2676)) + ((g1973) & (g1976) & (g2595) & (!g2643) & (g2048) & (!g2676)) + ((g1973) & (g1976) & (g2595) & (g2643) & (!g2048) & (g2676)) + ((g1973) & (g1976) & (g2595) & (g2643) & (g2048) & (!g2676)));
	assign g5827 = (((!g1973) & (!g1976) & (!g2595) & (!g2643) & (!g1970) & (!g2546)) + ((!g1973) & (!g1976) & (!g2595) & (!g2643) & (!g1970) & (g2546)) + ((!g1973) & (!g1976) & (!g2595) & (!g2643) & (g1970) & (!g2546)) + ((!g1973) & (!g1976) & (!g2595) & (g2643) & (!g1970) & (!g2546)) + ((!g1973) & (!g1976) & (!g2595) & (g2643) & (!g1970) & (g2546)) + ((!g1973) & (!g1976) & (!g2595) & (g2643) & (g1970) & (!g2546)) + ((!g1973) & (!g1976) & (g2595) & (!g2643) & (!g1970) & (!g2546)) + ((!g1973) & (!g1976) & (g2595) & (!g2643) & (!g1970) & (g2546)) + ((!g1973) & (!g1976) & (g2595) & (!g2643) & (g1970) & (!g2546)) + ((!g1973) & (!g1976) & (g2595) & (g2643) & (!g1970) & (!g2546)) + ((!g1973) & (!g1976) & (g2595) & (g2643) & (!g1970) & (g2546)) + ((!g1973) & (!g1976) & (g2595) & (g2643) & (g1970) & (!g2546)) + ((!g1973) & (g1976) & (!g2595) & (!g2643) & (!g1970) & (!g2546)) + ((!g1973) & (g1976) & (!g2595) & (!g2643) & (!g1970) & (g2546)) + ((!g1973) & (g1976) & (!g2595) & (!g2643) & (g1970) & (!g2546)) + ((!g1973) & (g1976) & (g2595) & (!g2643) & (!g1970) & (!g2546)) + ((!g1973) & (g1976) & (g2595) & (!g2643) & (!g1970) & (g2546)) + ((!g1973) & (g1976) & (g2595) & (!g2643) & (g1970) & (!g2546)) + ((g1973) & (!g1976) & (!g2595) & (!g2643) & (!g1970) & (!g2546)) + ((g1973) & (!g1976) & (!g2595) & (!g2643) & (!g1970) & (g2546)) + ((g1973) & (!g1976) & (!g2595) & (!g2643) & (g1970) & (!g2546)) + ((g1973) & (!g1976) & (!g2595) & (g2643) & (!g1970) & (!g2546)) + ((g1973) & (!g1976) & (!g2595) & (g2643) & (!g1970) & (g2546)) + ((g1973) & (!g1976) & (!g2595) & (g2643) & (g1970) & (!g2546)) + ((g1973) & (g1976) & (!g2595) & (!g2643) & (!g1970) & (!g2546)) + ((g1973) & (g1976) & (!g2595) & (!g2643) & (!g1970) & (g2546)) + ((g1973) & (g1976) & (!g2595) & (!g2643) & (g1970) & (!g2546)));
	assign g5828 = (((!g1970) & (!g2546) & (g5826) & (!g5827)) + ((!g1970) & (g2546) & (g5826) & (!g5827)) + ((!g1970) & (g2546) & (g5826) & (g5827)) + ((g1970) & (!g2546) & (g5826) & (!g5827)) + ((g1970) & (!g2546) & (g5826) & (g5827)) + ((g1970) & (g2546) & (g5826) & (!g5827)) + ((g1970) & (g2546) & (g5826) & (g5827)));
	assign g5829 = (((!g1996) & (!g1998) & (g2323) & (g2356) & (!g2001) & (g2402)) + ((!g1996) & (!g1998) & (g2323) & (g2356) & (g2001) & (!g2402)) + ((!g1996) & (g1998) & (!g2323) & (g2356) & (!g2001) & (g2402)) + ((!g1996) & (g1998) & (!g2323) & (g2356) & (g2001) & (!g2402)) + ((!g1996) & (g1998) & (g2323) & (!g2356) & (!g2001) & (g2402)) + ((!g1996) & (g1998) & (g2323) & (!g2356) & (g2001) & (!g2402)) + ((!g1996) & (g1998) & (g2323) & (g2356) & (!g2001) & (g2402)) + ((!g1996) & (g1998) & (g2323) & (g2356) & (g2001) & (!g2402)) + ((g1996) & (!g1998) & (!g2323) & (g2356) & (!g2001) & (g2402)) + ((g1996) & (!g1998) & (!g2323) & (g2356) & (g2001) & (!g2402)) + ((g1996) & (!g1998) & (g2323) & (g2356) & (!g2001) & (g2402)) + ((g1996) & (!g1998) & (g2323) & (g2356) & (g2001) & (!g2402)) + ((g1996) & (g1998) & (!g2323) & (!g2356) & (!g2001) & (g2402)) + ((g1996) & (g1998) & (!g2323) & (!g2356) & (g2001) & (!g2402)) + ((g1996) & (g1998) & (!g2323) & (g2356) & (!g2001) & (g2402)) + ((g1996) & (g1998) & (!g2323) & (g2356) & (g2001) & (!g2402)) + ((g1996) & (g1998) & (g2323) & (!g2356) & (!g2001) & (g2402)) + ((g1996) & (g1998) & (g2323) & (!g2356) & (g2001) & (!g2402)) + ((g1996) & (g1998) & (g2323) & (g2356) & (!g2001) & (g2402)) + ((g1996) & (g1998) & (g2323) & (g2356) & (g2001) & (!g2402)));
	assign g5830 = (((!g1996) & (!g1998) & (!g2323) & (!g2356) & (!g1993) & (!g2273)) + ((!g1996) & (!g1998) & (!g2323) & (!g2356) & (!g1993) & (g2273)) + ((!g1996) & (!g1998) & (!g2323) & (!g2356) & (g1993) & (!g2273)) + ((!g1996) & (!g1998) & (!g2323) & (g2356) & (!g1993) & (!g2273)) + ((!g1996) & (!g1998) & (!g2323) & (g2356) & (!g1993) & (g2273)) + ((!g1996) & (!g1998) & (!g2323) & (g2356) & (g1993) & (!g2273)) + ((!g1996) & (!g1998) & (g2323) & (!g2356) & (!g1993) & (!g2273)) + ((!g1996) & (!g1998) & (g2323) & (!g2356) & (!g1993) & (g2273)) + ((!g1996) & (!g1998) & (g2323) & (!g2356) & (g1993) & (!g2273)) + ((!g1996) & (!g1998) & (g2323) & (g2356) & (!g1993) & (!g2273)) + ((!g1996) & (!g1998) & (g2323) & (g2356) & (!g1993) & (g2273)) + ((!g1996) & (!g1998) & (g2323) & (g2356) & (g1993) & (!g2273)) + ((!g1996) & (g1998) & (!g2323) & (!g2356) & (!g1993) & (!g2273)) + ((!g1996) & (g1998) & (!g2323) & (!g2356) & (!g1993) & (g2273)) + ((!g1996) & (g1998) & (!g2323) & (!g2356) & (g1993) & (!g2273)) + ((!g1996) & (g1998) & (g2323) & (!g2356) & (!g1993) & (!g2273)) + ((!g1996) & (g1998) & (g2323) & (!g2356) & (!g1993) & (g2273)) + ((!g1996) & (g1998) & (g2323) & (!g2356) & (g1993) & (!g2273)) + ((g1996) & (!g1998) & (!g2323) & (!g2356) & (!g1993) & (!g2273)) + ((g1996) & (!g1998) & (!g2323) & (!g2356) & (!g1993) & (g2273)) + ((g1996) & (!g1998) & (!g2323) & (!g2356) & (g1993) & (!g2273)) + ((g1996) & (!g1998) & (!g2323) & (g2356) & (!g1993) & (!g2273)) + ((g1996) & (!g1998) & (!g2323) & (g2356) & (!g1993) & (g2273)) + ((g1996) & (!g1998) & (!g2323) & (g2356) & (g1993) & (!g2273)) + ((g1996) & (g1998) & (!g2323) & (!g2356) & (!g1993) & (!g2273)) + ((g1996) & (g1998) & (!g2323) & (!g2356) & (!g1993) & (g2273)) + ((g1996) & (g1998) & (!g2323) & (!g2356) & (g1993) & (!g2273)));
	assign g5831 = (((!g1993) & (!g2273) & (g5829) & (!g5830)) + ((!g1993) & (g2273) & (g5829) & (!g5830)) + ((!g1993) & (g2273) & (g5829) & (g5830)) + ((g1993) & (!g2273) & (g5829) & (!g5830)) + ((g1993) & (!g2273) & (g5829) & (g5830)) + ((g1993) & (g2273) & (g5829) & (!g5830)) + ((g1993) & (g2273) & (g5829) & (g5830)));
	assign g5832 = (((g830) & (g5833)));
	assign g5833 = (((!g5834) & (!g5835)));
	assign g5834 = (((!g1914) & (g5836)));
	assign g5835 = (((g1914) & (g5837)));
	assign g5836 = (((!g5558) & (g3389)) + ((g5558) & (!g3389)));
	assign g5837 = (((!g3854) & (!g2592) & (!g2589) & (g3389)) + ((!g3854) & (!g2592) & (g2589) & (!g3389)) + ((!g3854) & (g2592) & (!g2589) & (!g3389)) + ((!g3854) & (g2592) & (g2589) & (g3389)) + ((g3854) & (!g2592) & (!g2589) & (!g3389)) + ((g3854) & (!g2592) & (g2589) & (g3389)) + ((g3854) & (g2592) & (!g2589) & (g3389)) + ((g3854) & (g2592) & (g2589) & (!g3389)));
	assign g5838 = (((g830) & (g5839)));
	assign g5839 = (((!g5840) & (!g5841)));
	assign g5840 = (((!g1914) & (g5842)));
	assign g5841 = (((g1914) & (g5843)));
	assign g5842 = (((!g5544) & (g3380)) + ((g5544) & (!g3380)));
	assign g5843 = (((!g3697) & (!g2584) & (!g2575) & (g3380)) + ((!g3697) & (!g2584) & (g2575) & (!g3380)) + ((!g3697) & (g2584) & (!g2575) & (!g3380)) + ((!g3697) & (g2584) & (g2575) & (g3380)) + ((g3697) & (!g2584) & (!g2575) & (!g3380)) + ((g3697) & (!g2584) & (g2575) & (g3380)) + ((g3697) & (g2584) & (!g2575) & (g3380)) + ((g3697) & (g2584) & (g2575) & (!g3380)));
	assign g5844 = (((g830) & (g5845)));
	assign g5845 = (((!g5846) & (!g5847)));
	assign g5846 = (((!g1914) & (g5848)));
	assign g5847 = (((g1914) & (g5849)));
	assign g5848 = (((!g5530) & (g3370)) + ((g5530) & (!g3370)));
	assign g5849 = (((!g2569) & (!g3542) & (!g2011) & (g3370)) + ((!g2569) & (!g3542) & (g2011) & (!g3370)) + ((!g2569) & (g3542) & (!g2011) & (!g3370)) + ((!g2569) & (g3542) & (g2011) & (g3370)) + ((g2569) & (!g3542) & (!g2011) & (!g3370)) + ((g2569) & (!g3542) & (g2011) & (g3370)) + ((g2569) & (g3542) & (!g2011) & (g3370)) + ((g2569) & (g3542) & (g2011) & (!g3370)));
	assign g5850 = (((!g5851) & (!g5852)));
	assign g5851 = (((!g3003) & (g5853)));
	assign g5852 = (((g3003) & (g5856)));
	assign g5853 = (((!g5854) & (!g5855)));
	assign g5854 = (((!g1914) & (g5859)));
	assign g5855 = (((g1914) & (g5860)));
	assign g5856 = (((!g5857) & (!g5858)));
	assign g5857 = (((!g1914) & (g5861)));
	assign g5858 = (((g1914) & (g5862)));
	assign g5859 = (((!g3005) & (g5482)) + ((g3005) & (!g5482)));
	assign g5860 = (((!g5483) & (!g2101) & (g2733)) + ((!g5483) & (g2101) & (!g2733)) + ((g5483) & (!g2101) & (!g2733)) + ((g5483) & (g2101) & (g2733)));
	assign g5861 = (((!g3005) & (!g5482)) + ((g3005) & (g5482)));
	assign g5862 = (((!g5483) & (!g2101) & (g2733)) + ((!g5483) & (g2101) & (!g2733)) + ((g5483) & (!g2101) & (!g2733)) + ((g5483) & (g2101) & (g2733)));
	assign g5863 = (((!g5864) & (!g5865)));
	assign g5864 = (((!g2999) & (g5866)));
	assign g5865 = (((g2999) & (g5869)));
	assign g5866 = (((!g5867) & (!g5868)));
	assign g5867 = (((!g1914) & (g5872)));
	assign g5868 = (((g1914) & (g5873)));
	assign g5869 = (((!g5870) & (!g5871)));
	assign g5870 = (((!g1914) & (g5874)));
	assign g5871 = (((g1914) & (g5875)));
	assign g5872 = (((!g2713) & (!g2098) & (g5472)) + ((!g2713) & (g2098) & (!g5472)) + ((g2713) & (!g2098) & (!g5472)) + ((g2713) & (g2098) & (g5472)));
	assign g5873 = (((!g3013) & (g5471)) + ((g3013) & (!g5471)));
	assign g5874 = (((!g2713) & (!g2098) & (g5472)) + ((!g2713) & (g2098) & (!g5472)) + ((g2713) & (!g2098) & (!g5472)) + ((g2713) & (g2098) & (g5472)));
	assign g5875 = (((!g3013) & (!g5471)) + ((g3013) & (g5471)));
	assign g5876 = (((!g5877) & (!g5878)));
	assign g5877 = (((!g2348) & (g5879)));
	assign g5878 = (((g2348) & (g5882)));
	assign g5879 = (((!g5880) & (!g5881)));
	assign g5880 = (((!g1914) & (g5885)));
	assign g5881 = (((g1914) & (g5886)));
	assign g5882 = (((!g5883) & (!g5884)));
	assign g5883 = (((!g1914) & (g5887)));
	assign g5884 = (((g1914) & (g5888)));
	assign g5885 = (((!g5468) & (g1577)) + ((g5468) & (!g1577)));
	assign g5886 = (((!g2708) & (!g5469) & (g2747)) + ((!g2708) & (g5469) & (!g2747)) + ((g2708) & (!g5469) & (!g2747)) + ((g2708) & (g5469) & (g2747)));
	assign g5887 = (((!g5468) & (!g1577)) + ((g5468) & (g1577)));
	assign g5888 = (((!g2708) & (!g5469) & (g2747)) + ((!g2708) & (g5469) & (!g2747)) + ((g2708) & (!g5469) & (!g2747)) + ((g2708) & (g5469) & (g2747)));
	assign g5889 = (((!g5890) & (!g5891)));
	assign g5890 = (((!g3003) & (g5892)));
	assign g5891 = (((g3003) & (g5895)));
	assign g5892 = (((!g5893) & (!g5894)));
	assign g5893 = (((!g1914) & (g5898)));
	assign g5894 = (((g1914) & (g5899)));
	assign g5895 = (((!g5896) & (!g5897)));
	assign g5896 = (((!g1914) & (g5900)));
	assign g5897 = (((g1914) & (g5901)));
	assign g5898 = (((!g2747) & (!g2099) & (g5466)) + ((!g2747) & (g2099) & (!g5466)) + ((g2747) & (!g2099) & (!g5466)) + ((g2747) & (g2099) & (g5466)));
	assign g5899 = (((!g5465) & (g3011)) + ((g5465) & (!g3011)));
	assign g5900 = (((!g2747) & (!g2099) & (g5466)) + ((!g2747) & (g2099) & (!g5466)) + ((g2747) & (!g2099) & (!g5466)) + ((g2747) & (g2099) & (g5466)));
	assign g5901 = (((!g5465) & (!g3011)) + ((g5465) & (g3011)));
	assign g5902 = (((!g5903) & (!g5904)));
	assign g5903 = (((!g2344) & (g5905)));
	assign g5904 = (((g2344) & (g5908)));
	assign g5905 = (((!g5906) & (!g5907)));
	assign g5906 = (((!g1914) & (g5911)));
	assign g5907 = (((g1914) & (g5912)));
	assign g5908 = (((!g5909) & (!g5910)));
	assign g5909 = (((!g1914) & (g5913)));
	assign g5910 = (((g1914) & (g5914)));
	assign g5911 = (((!g5453) & (!g2733) & (g2723)) + ((!g5453) & (g2733) & (!g2723)) + ((g5453) & (!g2733) & (!g2723)) + ((g5453) & (g2733) & (g2723)));
	assign g5912 = (((!g5452) & (g1577)) + ((g5452) & (!g1577)));
	assign g5913 = (((!g5453) & (!g2733) & (g2723)) + ((!g5453) & (g2733) & (!g2723)) + ((g5453) & (!g2733) & (!g2723)) + ((g5453) & (g2733) & (g2723)));
	assign g5914 = (((!g5452) & (!g1577)) + ((g5452) & (g1577)));
	assign g5915 = (((g830) & (g5916)));
	assign g5916 = (((!g5917) & (!g5918)));
	assign g5917 = (((!g1914) & (g5919)));
	assign g5918 = (((g1914) & (g5920)));
	assign g5919 = (((!g3861) & (!g2416) & (!g2413) & (g3284)) + ((!g3861) & (!g2416) & (g2413) & (!g3284)) + ((!g3861) & (g2416) & (!g2413) & (!g3284)) + ((!g3861) & (g2416) & (g2413) & (g3284)) + ((g3861) & (!g2416) & (!g2413) & (!g3284)) + ((g3861) & (!g2416) & (g2413) & (g3284)) + ((g3861) & (g2416) & (!g2413) & (g3284)) + ((g3861) & (g2416) & (g2413) & (!g3284)));
	assign g5920 = (((!g5451) & (g3284)) + ((g5451) & (!g3284)));
	assign g5921 = (((g830) & (!g5922)));
	assign g5922 = (((g830) & (g5923)));
	assign g5923 = (((!g5924) & (!g5925)));
	assign g5924 = (((!g1914) & (g5926)));
	assign g5925 = (((g1914) & (g5927)));
	assign g5926 = (((!g3704) & (!g2408) & (!g2399) & (g3260)) + ((!g3704) & (!g2408) & (g2399) & (!g3260)) + ((!g3704) & (g2408) & (!g2399) & (!g3260)) + ((!g3704) & (g2408) & (g2399) & (g3260)) + ((g3704) & (!g2408) & (!g2399) & (!g3260)) + ((g3704) & (!g2408) & (g2399) & (g3260)) + ((g3704) & (g2408) & (!g2399) & (g3260)) + ((g3704) & (g2408) & (g2399) & (!g3260)));
	assign g5927 = (((!g5436) & (g3260)) + ((g5436) & (!g3260)));
	assign g5928 = (((g830) & (!g5929)));
	assign g5929 = (((g830) & (g5930)));
	assign g5930 = (((!g5931) & (!g5932)));
	assign g5931 = (((!g1914) & (g5933)));
	assign g5932 = (((g1914) & (g5934)));
	assign g5933 = (((!g3549) & (!g2393) & (!g1962) & (g3235)) + ((!g3549) & (!g2393) & (g1962) & (!g3235)) + ((!g3549) & (g2393) & (!g1962) & (!g3235)) + ((!g3549) & (g2393) & (g1962) & (g3235)) + ((g3549) & (!g2393) & (!g1962) & (!g3235)) + ((g3549) & (!g2393) & (g1962) & (g3235)) + ((g3549) & (g2393) & (!g1962) & (g3235)) + ((g3549) & (g2393) & (g1962) & (!g3235)));
	assign g5934 = (((!g5417) & (g3235)) + ((g5417) & (!g3235)));
	assign g5935 = (((g830) & (!g5936)));
	assign g5936 = (((g830) & (g5937)));
	assign g5937 = (((!g5938) & (!g5939)));
	assign g5938 = (((!g1914) & (g5940)));
	assign g5939 = (((g1914) & (g5941)));
	assign g5940 = (((!g5412) & (g3213)) + ((g5412) & (!g3213)));
	assign g5941 = (((!g5411) & (!g2371) & (!g2369) & (g3213)) + ((!g5411) & (!g2371) & (g2369) & (!g3213)) + ((!g5411) & (g2371) & (!g2369) & (!g3213)) + ((!g5411) & (g2371) & (g2369) & (g3213)) + ((g5411) & (!g2371) & (!g2369) & (!g3213)) + ((g5411) & (!g2371) & (g2369) & (g3213)) + ((g5411) & (g2371) & (!g2369) & (g3213)) + ((g5411) & (g2371) & (g2369) & (!g3213)));
	assign g5942 = (((!g5943) & (!g5944)));
	assign g5943 = (((!g2885) & (g5945)));
	assign g5944 = (((g2885) & (g5948)));
	assign g5945 = (((!g5946) & (!g5947)));
	assign g5946 = (((!g1914) & (g5951)));
	assign g5947 = (((g1914) & (g5406)));
	assign g5948 = (((!g5949) & (!g5950)));
	assign g5949 = (((!g1914) & (g5952)));
	assign g5950 = (((g1914) & (g5406)));
	assign g5951 = (((!g2857) & (!g2845) & (!g5362) & (g2887)) + ((!g2857) & (!g2845) & (g5362) & (g2887)) + ((!g2857) & (g2845) & (!g5362) & (g2887)) + ((!g2857) & (g2845) & (g5362) & (!g2887)) + ((g2857) & (!g2845) & (!g5362) & (g2887)) + ((g2857) & (!g2845) & (g5362) & (!g2887)) + ((g2857) & (g2845) & (!g5362) & (!g2887)) + ((g2857) & (g2845) & (g5362) & (!g2887)));
	assign g5952 = (((!g2857) & (!g2845) & (!g5362) & (!g2887)) + ((!g2857) & (!g2845) & (g5362) & (!g2887)) + ((!g2857) & (g2845) & (!g5362) & (!g2887)) + ((!g2857) & (g2845) & (g5362) & (g2887)) + ((g2857) & (!g2845) & (!g5362) & (!g2887)) + ((g2857) & (!g2845) & (g5362) & (g2887)) + ((g2857) & (g2845) & (!g5362) & (g2887)) + ((g2857) & (g2845) & (g5362) & (g2887)));
	assign g5953 = (((g830) & (g5954)));
	assign g5954 = (((!g5955) & (!g5956)));
	assign g5955 = (((!g1914) & (g5957)));
	assign g5956 = (((g1914) & (g5958)));
	assign g5957 = (((!g5402) & (g3199)) + ((g5402) & (!g3199)));
	assign g5958 = (((!g5401) & (!g2366) & (!g2360) & (g3199)) + ((!g5401) & (!g2366) & (g2360) & (!g3199)) + ((!g5401) & (g2366) & (!g2360) & (!g3199)) + ((!g5401) & (g2366) & (g2360) & (g3199)) + ((g5401) & (!g2366) & (!g2360) & (!g3199)) + ((g5401) & (!g2366) & (g2360) & (g3199)) + ((g5401) & (g2366) & (!g2360) & (g3199)) + ((g5401) & (g2366) & (g2360) & (!g3199)));
	assign g5959 = (((!g5960) & (!g5961)));
	assign g5960 = (((!g2881) & (g5962)));
	assign g5961 = (((g2881) & (g5965)));
	assign g5962 = (((!g5963) & (!g5964)));
	assign g5963 = (((!g1914) & (g5399)));
	assign g5964 = (((g1914) & (g5968)));
	assign g5965 = (((!g5966) & (!g5967)));
	assign g5966 = (((!g1914) & (g5399)));
	assign g5967 = (((g1914) & (g5969)));
	assign g5968 = (((!g5358) & (!g2854) & (!g2860) & (g2895)) + ((!g5358) & (!g2854) & (g2860) & (g2895)) + ((!g5358) & (g2854) & (!g2860) & (g2895)) + ((!g5358) & (g2854) & (g2860) & (!g2895)) + ((g5358) & (!g2854) & (!g2860) & (g2895)) + ((g5358) & (!g2854) & (g2860) & (!g2895)) + ((g5358) & (g2854) & (!g2860) & (!g2895)) + ((g5358) & (g2854) & (g2860) & (!g2895)));
	assign g5969 = (((!g5358) & (!g2854) & (!g2860) & (!g2895)) + ((!g5358) & (!g2854) & (g2860) & (!g2895)) + ((!g5358) & (g2854) & (!g2860) & (!g2895)) + ((!g5358) & (g2854) & (g2860) & (g2895)) + ((g5358) & (!g2854) & (!g2860) & (!g2895)) + ((g5358) & (!g2854) & (g2860) & (g2895)) + ((g5358) & (g2854) & (!g2860) & (g2895)) + ((g5358) & (g2854) & (g2860) & (g2895)));
	assign g5970 = (((!g5971) & (!g5972)));
	assign g5971 = (((!g2263) & (g5973)));
	assign g5972 = (((g2263) & (g5976)));
	assign g5973 = (((!g5974) & (!g5975)));
	assign g5974 = (((!g1914) & (g5979)));
	assign g5975 = (((g1914) & (g5397)));
	assign g5976 = (((!g5977) & (!g5978)));
	assign g5977 = (((!g1914) & (g5980)));
	assign g5978 = (((g1914) & (g5397)));
	assign g5979 = (((!g1473) & (!g2213) & (!g5353) & (g1507)) + ((!g1473) & (!g2213) & (g5353) & (g1507)) + ((!g1473) & (g2213) & (!g5353) & (g1507)) + ((!g1473) & (g2213) & (g5353) & (!g1507)) + ((g1473) & (!g2213) & (!g5353) & (g1507)) + ((g1473) & (!g2213) & (g5353) & (!g1507)) + ((g1473) & (g2213) & (!g5353) & (!g1507)) + ((g1473) & (g2213) & (g5353) & (!g1507)));
	assign g5980 = (((!g1473) & (!g2213) & (!g5353) & (!g1507)) + ((!g1473) & (!g2213) & (g5353) & (!g1507)) + ((!g1473) & (g2213) & (!g5353) & (!g1507)) + ((!g1473) & (g2213) & (g5353) & (g1507)) + ((g1473) & (!g2213) & (!g5353) & (!g1507)) + ((g1473) & (!g2213) & (g5353) & (g1507)) + ((g1473) & (g2213) & (!g5353) & (g1507)) + ((g1473) & (g2213) & (g5353) & (g1507)));
	assign g5981 = (((!g5982) & (!g5983)));
	assign g5982 = (((!g2885) & (g5984)));
	assign g5983 = (((g2885) & (g5987)));
	assign g5984 = (((!g5985) & (!g5986)));
	assign g5985 = (((!g1914) & (g5395)));
	assign g5986 = (((g1914) & (g5990)));
	assign g5987 = (((!g5988) & (!g5989)));
	assign g5988 = (((!g1914) & (g5395)));
	assign g5989 = (((g1914) & (g5991)));
	assign g5990 = (((!g2848) & (!g2845) & (!g5379) & (g2893)) + ((!g2848) & (!g2845) & (g5379) & (g2893)) + ((!g2848) & (g2845) & (!g5379) & (g2893)) + ((!g2848) & (g2845) & (g5379) & (!g2893)) + ((g2848) & (!g2845) & (!g5379) & (g2893)) + ((g2848) & (!g2845) & (g5379) & (!g2893)) + ((g2848) & (g2845) & (!g5379) & (!g2893)) + ((g2848) & (g2845) & (g5379) & (!g2893)));
	assign g5991 = (((!g2848) & (!g2845) & (!g5379) & (!g2893)) + ((!g2848) & (!g2845) & (g5379) & (!g2893)) + ((!g2848) & (g2845) & (!g5379) & (!g2893)) + ((!g2848) & (g2845) & (g5379) & (g2893)) + ((g2848) & (!g2845) & (!g5379) & (!g2893)) + ((g2848) & (!g2845) & (g5379) & (g2893)) + ((g2848) & (g2845) & (!g5379) & (g2893)) + ((g2848) & (g2845) & (g5379) & (g2893)));
	assign g5992 = (((g830) & (!g5993)));
	assign g5993 = (((g830) & (g5994)));
	assign g5994 = (((!g5995) & (!g5996)));
	assign g5995 = (((!g1914) & (g5997)));
	assign g5996 = (((g1914) & (g5998)));
	assign g5997 = (((!g5390) & (g3184)) + ((g5390) & (!g3184)));
	assign g5998 = (((!g2356) & (!g5389) & (!g1998) & (g3184)) + ((!g2356) & (!g5389) & (g1998) & (!g3184)) + ((!g2356) & (g5389) & (!g1998) & (!g3184)) + ((!g2356) & (g5389) & (g1998) & (g3184)) + ((g2356) & (!g5389) & (!g1998) & (!g3184)) + ((g2356) & (!g5389) & (g1998) & (g3184)) + ((g2356) & (g5389) & (!g1998) & (g3184)) + ((g2356) & (g5389) & (g1998) & (!g3184)));
	assign g5999 = (((!g6000) & (!g6001)));
	assign g6000 = (((!g2257) & (g6002)));
	assign g6001 = (((g2257) & (g6005)));
	assign g6002 = (((!g6003) & (!g6004)));
	assign g6003 = (((!g1914) & (g5387)));
	assign g6004 = (((g1914) & (g6008)));
	assign g6005 = (((!g6006) & (!g6007)));
	assign g6006 = (((!g1914) & (g5387)));
	assign g6007 = (((g1914) & (g6009)));
	assign g6008 = (((!g1473) & (!g2211) & (!g5366) & (g1507)) + ((!g1473) & (!g2211) & (g5366) & (g1507)) + ((!g1473) & (g2211) & (!g5366) & (g1507)) + ((!g1473) & (g2211) & (g5366) & (!g1507)) + ((g1473) & (!g2211) & (!g5366) & (g1507)) + ((g1473) & (!g2211) & (g5366) & (!g1507)) + ((g1473) & (g2211) & (!g5366) & (!g1507)) + ((g1473) & (g2211) & (g5366) & (!g1507)));
	assign g6009 = (((!g1473) & (!g2211) & (!g5366) & (!g1507)) + ((!g1473) & (!g2211) & (g5366) & (!g1507)) + ((!g1473) & (g2211) & (!g5366) & (!g1507)) + ((!g1473) & (g2211) & (g5366) & (g1507)) + ((g1473) & (!g2211) & (!g5366) & (!g1507)) + ((g1473) & (!g2211) & (g5366) & (g1507)) + ((g1473) & (g2211) & (!g5366) & (g1507)) + ((g1473) & (g2211) & (g5366) & (g1507)));
	assign g6010 = (((g830) & (g6011)));
	assign g6011 = (((!g6012) & (!g6013)));
	assign g6012 = (((!g1914) & (g6014)));
	assign g6013 = (((g1914) & (g6015)));
	assign g6014 = (((!g5386) & (g3172)) + ((g5386) & (!g3172)));
	assign g6015 = (((!g3850) & (!g2329) & (!g2317) & (g3172)) + ((!g3850) & (!g2329) & (g2317) & (!g3172)) + ((!g3850) & (g2329) & (!g2317) & (!g3172)) + ((!g3850) & (g2329) & (g2317) & (g3172)) + ((g3850) & (!g2329) & (!g2317) & (!g3172)) + ((g3850) & (!g2329) & (g2317) & (g3172)) + ((g3850) & (g2329) & (!g2317) & (g3172)) + ((g3850) & (g2329) & (g2317) & (!g3172)));
	assign g6016 = (((g830) & (g6017)));
	assign g6017 = (((!g6018) & (!g6019)));
	assign g6018 = (((!g1914) & (g6020)));
	assign g6019 = (((g1914) & (g6021)));
	assign g6020 = (((!g5375) & (g3163)) + ((g5375) & (!g3163)));
	assign g6021 = (((!g3693) & (!g2337) & (!g2304) & (g3163)) + ((!g3693) & (!g2337) & (g2304) & (!g3163)) + ((!g3693) & (g2337) & (!g2304) & (!g3163)) + ((!g3693) & (g2337) & (g2304) & (g3163)) + ((g3693) & (!g2337) & (!g2304) & (!g3163)) + ((g3693) & (!g2337) & (g2304) & (g3163)) + ((g3693) & (g2337) & (!g2304) & (g3163)) + ((g3693) & (g2337) & (g2304) & (!g3163)));
	assign g6022 = (((g830) & (g6023)));
	assign g6023 = (((!g6024) & (!g6025)));
	assign g6024 = (((!g1914) & (g6026)));
	assign g6025 = (((g1914) & (g6027)));
	assign g6026 = (((!g5357) & (g3153)) + ((g5357) & (!g3153)));
	assign g6027 = (((!g2323) & (!g3539) & (!g1996) & (g3153)) + ((!g2323) & (!g3539) & (g1996) & (!g3153)) + ((!g2323) & (g3539) & (!g1996) & (!g3153)) + ((!g2323) & (g3539) & (g1996) & (g3153)) + ((g2323) & (!g3539) & (!g1996) & (!g3153)) + ((g2323) & (!g3539) & (g1996) & (g3153)) + ((g2323) & (g3539) & (!g1996) & (g3153)) + ((g2323) & (g3539) & (g1996) & (!g3153)));
	assign g6028 = (((!g6029) & (!g6030)));
	assign g6029 = (((!g2768) & (g6031)));
	assign g6030 = (((g2768) & (g6034)));
	assign g6031 = (((!g6032) & (!g6033)));
	assign g6032 = (((!g1914) & (g5305)));
	assign g6033 = (((g1914) & (g6037)));
	assign g6034 = (((!g6035) & (!g6036)));
	assign g6035 = (((!g1914) & (g5305)));
	assign g6036 = (((g1914) & (g6038)));
	assign g6037 = (((!g2723) & (!g2703) & (!g5243) & (g2770)) + ((!g2723) & (!g2703) & (g5243) & (g2770)) + ((!g2723) & (g2703) & (!g5243) & (g2770)) + ((!g2723) & (g2703) & (g5243) & (!g2770)) + ((g2723) & (!g2703) & (!g5243) & (g2770)) + ((g2723) & (!g2703) & (g5243) & (!g2770)) + ((g2723) & (g2703) & (!g5243) & (!g2770)) + ((g2723) & (g2703) & (g5243) & (!g2770)));
	assign g6038 = (((!g2723) & (!g2703) & (!g5243) & (!g2770)) + ((!g2723) & (!g2703) & (g5243) & (!g2770)) + ((!g2723) & (g2703) & (!g5243) & (!g2770)) + ((!g2723) & (g2703) & (g5243) & (g2770)) + ((g2723) & (!g2703) & (!g5243) & (!g2770)) + ((g2723) & (!g2703) & (g5243) & (g2770)) + ((g2723) & (g2703) & (!g5243) & (g2770)) + ((g2723) & (g2703) & (g5243) & (g2770)));
	assign g6039 = (((!g6040) & (!g6041)));
	assign g6040 = (((!g2764) & (g6042)));
	assign g6041 = (((g2764) & (g6045)));
	assign g6042 = (((!g6043) & (!g6044)));
	assign g6043 = (((!g1914) & (g6048)));
	assign g6044 = (((g1914) & (g5293)));
	assign g6045 = (((!g6046) & (!g6047)));
	assign g6046 = (((!g1914) & (g6049)));
	assign g6047 = (((g1914) & (g5293)));
	assign g6048 = (((!g2728) & (!g2718) & (!g5238) & (g2778)) + ((!g2728) & (!g2718) & (g5238) & (g2778)) + ((!g2728) & (g2718) & (!g5238) & (g2778)) + ((!g2728) & (g2718) & (g5238) & (!g2778)) + ((g2728) & (!g2718) & (!g5238) & (g2778)) + ((g2728) & (!g2718) & (g5238) & (!g2778)) + ((g2728) & (g2718) & (!g5238) & (!g2778)) + ((g2728) & (g2718) & (g5238) & (!g2778)));
	assign g6049 = (((!g2728) & (!g2718) & (!g5238) & (!g2778)) + ((!g2728) & (!g2718) & (g5238) & (!g2778)) + ((!g2728) & (g2718) & (!g5238) & (!g2778)) + ((!g2728) & (g2718) & (g5238) & (g2778)) + ((g2728) & (!g2718) & (!g5238) & (!g2778)) + ((g2728) & (!g2718) & (g5238) & (g2778)) + ((g2728) & (g2718) & (!g5238) & (g2778)) + ((g2728) & (g2718) & (g5238) & (g2778)));
	assign g6050 = (((!g6051) & (!g6052)));
	assign g6051 = (((!g2130) & (g6053)));
	assign g6052 = (((g2130) & (g6056)));
	assign g6053 = (((!g6054) & (!g6055)));
	assign g6054 = (((!g1914) & (g5290)));
	assign g6055 = (((g1914) & (g6059)));
	assign g6056 = (((!g6057) & (!g6058)));
	assign g6057 = (((!g1914) & (g5290)));
	assign g6058 = (((g1914) & (g6060)));
	assign g6059 = (((!g1370) & (!g2099) & (!g5231) & (g1406)) + ((!g1370) & (!g2099) & (g5231) & (g1406)) + ((!g1370) & (g2099) & (!g5231) & (g1406)) + ((!g1370) & (g2099) & (g5231) & (!g1406)) + ((g1370) & (!g2099) & (!g5231) & (g1406)) + ((g1370) & (!g2099) & (g5231) & (!g1406)) + ((g1370) & (g2099) & (!g5231) & (!g1406)) + ((g1370) & (g2099) & (g5231) & (!g1406)));
	assign g6060 = (((!g1370) & (!g2099) & (!g5231) & (!g1406)) + ((!g1370) & (!g2099) & (g5231) & (!g1406)) + ((!g1370) & (g2099) & (!g5231) & (!g1406)) + ((!g1370) & (g2099) & (g5231) & (g1406)) + ((g1370) & (!g2099) & (!g5231) & (!g1406)) + ((g1370) & (!g2099) & (g5231) & (g1406)) + ((g1370) & (g2099) & (!g5231) & (g1406)) + ((g1370) & (g2099) & (g5231) & (g1406)));
	assign g6061 = (((!g6062) & (!g6063)));
	assign g6062 = (((!g2768) & (g6064)));
	assign g6063 = (((g2768) & (g6067)));
	assign g6064 = (((!g6065) & (!g6066)));
	assign g6065 = (((!g1914) & (g6070)));
	assign g6066 = (((g1914) & (g5287)));
	assign g6067 = (((!g6068) & (!g6069)));
	assign g6068 = (((!g1914) & (g6071)));
	assign g6069 = (((g1914) & (g5287)));
	assign g6070 = (((!g2708) & (!g2703) & (!g5263) & (g2776)) + ((!g2708) & (!g2703) & (g5263) & (g2776)) + ((!g2708) & (g2703) & (!g5263) & (g2776)) + ((!g2708) & (g2703) & (g5263) & (!g2776)) + ((g2708) & (!g2703) & (!g5263) & (g2776)) + ((g2708) & (!g2703) & (g5263) & (!g2776)) + ((g2708) & (g2703) & (!g5263) & (!g2776)) + ((g2708) & (g2703) & (g5263) & (!g2776)));
	assign g6071 = (((!g2708) & (!g2703) & (!g5263) & (!g2776)) + ((!g2708) & (!g2703) & (g5263) & (!g2776)) + ((!g2708) & (g2703) & (!g5263) & (!g2776)) + ((!g2708) & (g2703) & (g5263) & (g2776)) + ((g2708) & (!g2703) & (!g5263) & (!g2776)) + ((g2708) & (!g2703) & (g5263) & (g2776)) + ((g2708) & (g2703) & (!g5263) & (g2776)) + ((g2708) & (g2703) & (g5263) & (g2776)));
	assign g6072 = (((!g6073) & (!g6074)));
	assign g6073 = (((!g2774) & (g6075)));
	assign g6074 = (((g2774) & (g6078)));
	assign g6075 = (((!g6076) & (!g6077)));
	assign g6076 = (((!g1914) & (g5284)));
	assign g6077 = (((g1914) & (g6081)));
	assign g6078 = (((!g6079) & (!g6080)));
	assign g6079 = (((!g1914) & (g5284)));
	assign g6080 = (((g1914) & (g6082)));
	assign g6081 = (((!g5251) & (!g2690) & (!g2728) & (g2778)) + ((!g5251) & (!g2690) & (g2728) & (g2778)) + ((!g5251) & (g2690) & (!g2728) & (g2778)) + ((!g5251) & (g2690) & (g2728) & (!g2778)) + ((g5251) & (!g2690) & (!g2728) & (g2778)) + ((g5251) & (!g2690) & (g2728) & (!g2778)) + ((g5251) & (g2690) & (!g2728) & (!g2778)) + ((g5251) & (g2690) & (g2728) & (!g2778)));
	assign g6082 = (((!g5251) & (!g2690) & (!g2728) & (!g2778)) + ((!g5251) & (!g2690) & (g2728) & (!g2778)) + ((!g5251) & (g2690) & (!g2728) & (!g2778)) + ((!g5251) & (g2690) & (g2728) & (g2778)) + ((g5251) & (!g2690) & (!g2728) & (!g2778)) + ((g5251) & (!g2690) & (g2728) & (g2778)) + ((g5251) & (g2690) & (!g2728) & (g2778)) + ((g5251) & (g2690) & (g2728) & (g2778)));
	assign g6083 = (((!g6084) & (!g6085)));
	assign g6084 = (((!g2134) & (g6086)));
	assign g6085 = (((g2134) & (g6089)));
	assign g6086 = (((!g6087) & (!g6088)));
	assign g6087 = (((!g1914) & (g6092)));
	assign g6088 = (((g1914) & (g5276)));
	assign g6089 = (((!g6090) & (!g6091)));
	assign g6090 = (((!g1914) & (g6093)));
	assign g6091 = (((g1914) & (g5276)));
	assign g6092 = (((!g1370) & (!g2101) & (!g5247) & (g1406)) + ((!g1370) & (!g2101) & (g5247) & (g1406)) + ((!g1370) & (g2101) & (!g5247) & (g1406)) + ((!g1370) & (g2101) & (g5247) & (!g1406)) + ((g1370) & (!g2101) & (!g5247) & (g1406)) + ((g1370) & (!g2101) & (g5247) & (!g1406)) + ((g1370) & (g2101) & (!g5247) & (!g1406)) + ((g1370) & (g2101) & (g5247) & (!g1406)));
	assign g6093 = (((!g1370) & (!g2101) & (!g5247) & (!g1406)) + ((!g1370) & (!g2101) & (g5247) & (!g1406)) + ((!g1370) & (g2101) & (!g5247) & (!g1406)) + ((!g1370) & (g2101) & (g5247) & (g1406)) + ((g1370) & (!g2101) & (!g5247) & (!g1406)) + ((g1370) & (!g2101) & (g5247) & (g1406)) + ((g1370) & (g2101) & (!g5247) & (g1406)) + ((g1370) & (g2101) & (g5247) & (g1406)));
	assign g6094 = (((!g6095) & (!g6096)));
	assign g6095 = (((!g2657) & (g6097)));
	assign g6096 = (((g2657) & (g6100)));
	assign g6097 = (((!g6098) & (!g6099)));
	assign g6098 = (((!g1914) & (g5221)));
	assign g6099 = (((g1914) & (g6103)));
	assign g6100 = (((!g6101) & (!g6102)));
	assign g6101 = (((!g1914) & (g5221)));
	assign g6102 = (((g1914) & (g6104)));
	assign g6103 = (((!g2626) & (!g2614) & (!g5167) & (g2659)) + ((!g2626) & (!g2614) & (g5167) & (g2659)) + ((!g2626) & (g2614) & (!g5167) & (g2659)) + ((!g2626) & (g2614) & (g5167) & (!g2659)) + ((g2626) & (!g2614) & (!g5167) & (g2659)) + ((g2626) & (!g2614) & (g5167) & (!g2659)) + ((g2626) & (g2614) & (!g5167) & (!g2659)) + ((g2626) & (g2614) & (g5167) & (!g2659)));
	assign g6104 = (((!g2626) & (!g2614) & (!g5167) & (!g2659)) + ((!g2626) & (!g2614) & (g5167) & (!g2659)) + ((!g2626) & (g2614) & (!g5167) & (!g2659)) + ((!g2626) & (g2614) & (g5167) & (g2659)) + ((g2626) & (!g2614) & (!g5167) & (!g2659)) + ((g2626) & (!g2614) & (g5167) & (g2659)) + ((g2626) & (g2614) & (!g5167) & (g2659)) + ((g2626) & (g2614) & (g5167) & (g2659)));
	assign g6105 = (((!g6106) & (!g6107)));
	assign g6106 = (((!g2653) & (g6108)));
	assign g6107 = (((g2653) & (g6111)));
	assign g6108 = (((!g6109) & (!g6110)));
	assign g6109 = (((!g1914) & (g6114)));
	assign g6110 = (((g1914) & (g5209)));
	assign g6111 = (((!g6112) & (!g6113)));
	assign g6112 = (((!g1914) & (g6115)));
	assign g6113 = (((g1914) & (g5209)));
	assign g6114 = (((!g2629) & (!g2623) & (!g5162) & (g2667)) + ((!g2629) & (!g2623) & (g5162) & (g2667)) + ((!g2629) & (g2623) & (!g5162) & (g2667)) + ((!g2629) & (g2623) & (g5162) & (!g2667)) + ((g2629) & (!g2623) & (!g5162) & (g2667)) + ((g2629) & (!g2623) & (g5162) & (!g2667)) + ((g2629) & (g2623) & (!g5162) & (!g2667)) + ((g2629) & (g2623) & (g5162) & (!g2667)));
	assign g6115 = (((!g2629) & (!g2623) & (!g5162) & (!g2667)) + ((!g2629) & (!g2623) & (g5162) & (!g2667)) + ((!g2629) & (g2623) & (!g5162) & (!g2667)) + ((!g2629) & (g2623) & (g5162) & (g2667)) + ((g2629) & (!g2623) & (!g5162) & (!g2667)) + ((g2629) & (!g2623) & (g5162) & (g2667)) + ((g2629) & (g2623) & (!g5162) & (g2667)) + ((g2629) & (g2623) & (g5162) & (g2667)));
	assign g6116 = (((!g6117) & (!g6118)));
	assign g6117 = (((!g2048) & (g6119)));
	assign g6118 = (((g2048) & (g6122)));
	assign g6119 = (((!g6120) & (!g6121)));
	assign g6120 = (((!g1914) & (g5206)));
	assign g6121 = (((g1914) & (g6125)));
	assign g6122 = (((!g6123) & (!g6124)));
	assign g6123 = (((!g1914) & (g5206)));
	assign g6124 = (((g1914) & (g6126)));
	assign g6125 = (((!g1303) & (!g1976) & (!g5157) & (g1337)) + ((!g1303) & (!g1976) & (g5157) & (g1337)) + ((!g1303) & (g1976) & (!g5157) & (g1337)) + ((!g1303) & (g1976) & (g5157) & (!g1337)) + ((g1303) & (!g1976) & (!g5157) & (g1337)) + ((g1303) & (!g1976) & (g5157) & (!g1337)) + ((g1303) & (g1976) & (!g5157) & (!g1337)) + ((g1303) & (g1976) & (g5157) & (!g1337)));
	assign g6126 = (((!g1303) & (!g1976) & (!g5157) & (!g1337)) + ((!g1303) & (!g1976) & (g5157) & (!g1337)) + ((!g1303) & (g1976) & (!g5157) & (!g1337)) + ((!g1303) & (g1976) & (g5157) & (g1337)) + ((g1303) & (!g1976) & (!g5157) & (!g1337)) + ((g1303) & (!g1976) & (g5157) & (g1337)) + ((g1303) & (g1976) & (!g5157) & (g1337)) + ((g1303) & (g1976) & (g5157) & (g1337)));
	assign g6127 = (((!g6128) & (!g6129)));
	assign g6128 = (((!g2657) & (g6130)));
	assign g6129 = (((g2657) & (g6133)));
	assign g6130 = (((!g6131) & (!g6132)));
	assign g6131 = (((!g1914) & (g6136)));
	assign g6132 = (((g1914) & (g5203)));
	assign g6133 = (((!g6134) & (!g6135)));
	assign g6134 = (((!g1914) & (g6137)));
	assign g6135 = (((g1914) & (g5203)));
	assign g6136 = (((!g2617) & (!g2614) & (!g5183) & (g2665)) + ((!g2617) & (!g2614) & (g5183) & (g2665)) + ((!g2617) & (g2614) & (!g5183) & (g2665)) + ((!g2617) & (g2614) & (g5183) & (!g2665)) + ((g2617) & (!g2614) & (!g5183) & (g2665)) + ((g2617) & (!g2614) & (g5183) & (!g2665)) + ((g2617) & (g2614) & (!g5183) & (!g2665)) + ((g2617) & (g2614) & (g5183) & (!g2665)));
	assign g6137 = (((!g2617) & (!g2614) & (!g5183) & (!g2665)) + ((!g2617) & (!g2614) & (g5183) & (!g2665)) + ((!g2617) & (g2614) & (!g5183) & (!g2665)) + ((!g2617) & (g2614) & (g5183) & (g2665)) + ((g2617) & (!g2614) & (!g5183) & (!g2665)) + ((g2617) & (!g2614) & (g5183) & (g2665)) + ((g2617) & (g2614) & (!g5183) & (g2665)) + ((g2617) & (g2614) & (g5183) & (g2665)));
	assign g6138 = (((!g6139) & (!g6140)));
	assign g6139 = (((!g2663) & (g6141)));
	assign g6140 = (((g2663) & (g6144)));
	assign g6141 = (((!g6142) & (!g6143)));
	assign g6142 = (((!g1914) & (g5200)));
	assign g6143 = (((g1914) & (g6147)));
	assign g6144 = (((!g6145) & (!g6146)));
	assign g6145 = (((!g1914) & (g5200)));
	assign g6146 = (((g1914) & (g6148)));
	assign g6147 = (((!g5175) & (!g2607) & (!g2629) & (g2667)) + ((!g5175) & (!g2607) & (g2629) & (g2667)) + ((!g5175) & (g2607) & (!g2629) & (g2667)) + ((!g5175) & (g2607) & (g2629) & (!g2667)) + ((g5175) & (!g2607) & (!g2629) & (g2667)) + ((g5175) & (!g2607) & (g2629) & (!g2667)) + ((g5175) & (g2607) & (!g2629) & (!g2667)) + ((g5175) & (g2607) & (g2629) & (!g2667)));
	assign g6148 = (((!g5175) & (!g2607) & (!g2629) & (!g2667)) + ((!g5175) & (!g2607) & (g2629) & (!g2667)) + ((!g5175) & (g2607) & (!g2629) & (!g2667)) + ((!g5175) & (g2607) & (g2629) & (g2667)) + ((g5175) & (!g2607) & (!g2629) & (!g2667)) + ((g5175) & (!g2607) & (g2629) & (g2667)) + ((g5175) & (g2607) & (!g2629) & (g2667)) + ((g5175) & (g2607) & (g2629) & (g2667)));
	assign g6149 = (((!g6150) & (!g6151)));
	assign g6150 = (((!g2052) & (g6152)));
	assign g6151 = (((g2052) & (g6155)));
	assign g6152 = (((!g6153) & (!g6154)));
	assign g6153 = (((!g1914) & (g6158)));
	assign g6154 = (((g1914) & (g5192)));
	assign g6155 = (((!g6156) & (!g6157)));
	assign g6156 = (((!g1914) & (g6159)));
	assign g6157 = (((g1914) & (g5192)));
	assign g6158 = (((!g1303) & (!g2014) & (!g5171) & (g1337)) + ((!g1303) & (!g2014) & (g5171) & (g1337)) + ((!g1303) & (g2014) & (!g5171) & (g1337)) + ((!g1303) & (g2014) & (g5171) & (!g1337)) + ((g1303) & (!g2014) & (!g5171) & (g1337)) + ((g1303) & (!g2014) & (g5171) & (!g1337)) + ((g1303) & (g2014) & (!g5171) & (!g1337)) + ((g1303) & (g2014) & (g5171) & (!g1337)));
	assign g6159 = (((!g1303) & (!g2014) & (!g5171) & (!g1337)) + ((!g1303) & (!g2014) & (g5171) & (!g1337)) + ((!g1303) & (g2014) & (!g5171) & (!g1337)) + ((!g1303) & (g2014) & (g5171) & (g1337)) + ((g1303) & (!g2014) & (!g5171) & (!g1337)) + ((g1303) & (!g2014) & (g5171) & (g1337)) + ((g1303) & (g2014) & (!g5171) & (g1337)) + ((g1303) & (g2014) & (g5171) & (g1337)));
	assign g6160 = (((g830) & (!g6161)));
	assign g6161 = (((g830) & (g6162)));
	assign g6162 = (((!g6163) & (!g6164)));
	assign g6163 = (((!g1914) & (g6165)));
	assign g6164 = (((g1914) & (g6166)));
	assign g6165 = (((!g5190) & (g2991)) + ((g5190) & (!g2991)));
	assign g6166 = (((!g3846) & (!g2125) & (!g2123) & (g2991)) + ((!g3846) & (!g2125) & (g2123) & (!g2991)) + ((!g3846) & (g2125) & (!g2123) & (!g2991)) + ((!g3846) & (g2125) & (g2123) & (g2991)) + ((g3846) & (!g2125) & (!g2123) & (!g2991)) + ((g3846) & (!g2125) & (g2123) & (g2991)) + ((g3846) & (g2125) & (!g2123) & (g2991)) + ((g3846) & (g2125) & (g2123) & (!g2991)));
	assign g6167 = (((g830) & (!g6168)));
	assign g6168 = (((g830) & (g6169)));
	assign g6169 = (((!g6170) & (!g6171)));
	assign g6170 = (((!g1914) & (g6172)));
	assign g6171 = (((g1914) & (g6173)));
	assign g6172 = (((!g5179) & (g2962)) + ((g5179) & (!g2962)));
	assign g6173 = (((!g3689) & (!g2120) & (!g2114) & (g2962)) + ((!g3689) & (!g2120) & (g2114) & (!g2962)) + ((!g3689) & (g2120) & (!g2114) & (!g2962)) + ((!g3689) & (g2120) & (g2114) & (g2962)) + ((g3689) & (!g2120) & (!g2114) & (!g2962)) + ((g3689) & (!g2120) & (g2114) & (g2962)) + ((g3689) & (g2120) & (!g2114) & (g2962)) + ((g3689) & (g2120) & (g2114) & (!g2962)));
	assign g6174 = (((g830) & (!g6175)));
	assign g6175 = (((g830) & (g6176)));
	assign g6176 = (((!g6177) & (!g6178)));
	assign g6177 = (((!g1914) & (g6179)));
	assign g6178 = (((g1914) & (g6180)));
	assign g6179 = (((!g5161) & (g2932)) + ((g5161) & (!g2932)));
	assign g6180 = (((!g2110) & (!g3535) & (!g1982) & (g2932)) + ((!g2110) & (!g3535) & (g1982) & (!g2932)) + ((!g2110) & (g3535) & (!g1982) & (!g2932)) + ((!g2110) & (g3535) & (g1982) & (g2932)) + ((g2110) & (!g3535) & (!g1982) & (!g2932)) + ((g2110) & (!g3535) & (g1982) & (g2932)) + ((g2110) & (g3535) & (!g1982) & (g2932)) + ((g2110) & (g3535) & (g1982) & (!g2932)));
	assign g6181 = (((g830) & (g6182)));
	assign g6182 = (((!g6183) & (!g6184)));
	assign g6183 = (((!g1914) & (g6185)));
	assign g6184 = (((g1914) & (g6186)));
	assign g6185 = (((!g1910) & (!g1908) & (g2833)) + ((!g1910) & (g1908) & (!g2833)) + ((g1910) & (!g1908) & (!g2833)) + ((g1910) & (g1908) & (g2833)));
	assign g6186 = (((!g1904) & (!g1896) & (g2833)) + ((!g1904) & (g1896) & (!g2833)) + ((g1904) & (!g1896) & (!g2833)) + ((g1904) & (g1896) & (g2833)));
	assign g6187 = (((g830) & (g6188)));
	assign g6188 = (((!g6189) & (!g6190)));
	assign g6189 = (((!g1914) & (g6191)));
	assign g6190 = (((g1914) & (g6192)));
	assign g6191 = (((!g1904) & (!g1898) & (g2819)) + ((!g1904) & (g1898) & (!g2819)) + ((g1904) & (!g1898) & (!g2819)) + ((g1904) & (g1898) & (g2819)));
	assign g6192 = (((!g1910) & (!g1886) & (g2819)) + ((!g1910) & (g1886) & (!g2819)) + ((g1910) & (!g1886) & (!g2819)) + ((g1910) & (g1886) & (g2819)));
	assign g6193 = (((g830) & (g6194)));
	assign g6194 = (((!g6195) & (!g6196)));
	assign g6195 = (((!g1914) & (g6197)));
	assign g6196 = (((g1914) & (g6198)));
	assign g6197 = (((!g1894) & (!g1890) & (g2804)) + ((!g1894) & (g1890) & (!g2804)) + ((g1894) & (!g1890) & (!g2804)) + ((g1894) & (g1890) & (g2804)));
	assign g6198 = (((!g1900) & (!g1884) & (g2804)) + ((!g1900) & (g1884) & (!g2804)) + ((g1900) & (!g1884) & (!g2804)) + ((g1900) & (g1884) & (g2804)));
	assign g6199 = (((g830) & (g6200)));
	assign g6200 = (((!g6201) & (!g6202)));
	assign g6201 = (((!g1914) & (g6203)));
	assign g6202 = (((g1914) & (g6204)));
	assign g6203 = (((!g3382) & (!g3374) & (!g5022) & (g2787)) + ((!g3382) & (!g3374) & (g5022) & (!g2787)) + ((!g3382) & (g3374) & (!g5022) & (!g2787)) + ((!g3382) & (g3374) & (g5022) & (g2787)) + ((g3382) & (!g3374) & (!g5022) & (!g2787)) + ((g3382) & (!g3374) & (g5022) & (g2787)) + ((g3382) & (g3374) & (!g5022) & (g2787)) + ((g3382) & (g3374) & (g5022) & (!g2787)));
	assign g6204 = (((!g5021) & (g2787)) + ((g5021) & (!g2787)));
	assign g6205 = (((!g6206) & (!g6207)));
	assign g6206 = (((!g2390) & (g6208)));
	assign g6207 = (((g2390) & (g6211)));
	assign g6208 = (((!g6209) & (!g6210)));
	assign g6209 = (((!g1914) & (g6214)));
	assign g6210 = (((g1914) & (g5016)));
	assign g6211 = (((!g6212) & (!g6213)));
	assign g6212 = (((!g1914) & (g6215)));
	assign g6213 = (((g1914) & (g5016)));
	assign g6214 = (((!g2362) & (!g2354) & (!g4948) & (g2393)) + ((!g2362) & (!g2354) & (g4948) & (g2393)) + ((!g2362) & (g2354) & (!g4948) & (g2393)) + ((!g2362) & (g2354) & (g4948) & (!g2393)) + ((g2362) & (!g2354) & (!g4948) & (g2393)) + ((g2362) & (!g2354) & (g4948) & (!g2393)) + ((g2362) & (g2354) & (!g4948) & (!g2393)) + ((g2362) & (g2354) & (g4948) & (!g2393)));
	assign g6215 = (((!g2362) & (!g2354) & (!g4948) & (!g2393)) + ((!g2362) & (!g2354) & (g4948) & (!g2393)) + ((!g2362) & (g2354) & (!g4948) & (!g2393)) + ((!g2362) & (g2354) & (g4948) & (g2393)) + ((g2362) & (!g2354) & (!g4948) & (!g2393)) + ((g2362) & (!g2354) & (g4948) & (g2393)) + ((g2362) & (g2354) & (!g4948) & (g2393)) + ((g2362) & (g2354) & (g4948) & (g2393)));
	assign g6216 = (((g830) & (g6217)));
	assign g6217 = (((!g6218) & (!g6219)));
	assign g6218 = (((!g1914) & (g6220)));
	assign g6219 = (((g1914) & (g6221)));
	assign g6220 = (((!g3387) & (!g3366) & (!g5011) & (g2778)) + ((!g3387) & (!g3366) & (g5011) & (!g2778)) + ((!g3387) & (g3366) & (!g5011) & (!g2778)) + ((!g3387) & (g3366) & (g5011) & (g2778)) + ((g3387) & (!g3366) & (!g5011) & (!g2778)) + ((g3387) & (!g3366) & (g5011) & (g2778)) + ((g3387) & (g3366) & (!g5011) & (g2778)) + ((g3387) & (g3366) & (g5011) & (!g2778)));
	assign g6221 = (((!g5010) & (g2778)) + ((g5010) & (!g2778)));
	assign g6222 = (((!g6223) & (!g6224)));
	assign g6223 = (((!g2383) & (g6225)));
	assign g6224 = (((g2383) & (g6228)));
	assign g6225 = (((!g6226) & (!g6227)));
	assign g6226 = (((!g1914) & (g5008)));
	assign g6227 = (((g1914) & (g6231)));
	assign g6228 = (((!g6229) & (!g6230)));
	assign g6229 = (((!g1914) & (g5008)));
	assign g6230 = (((g1914) & (g6232)));
	assign g6231 = (((!g4944) & (!g2360) & (!g2364) & (g2405)) + ((!g4944) & (!g2360) & (g2364) & (g2405)) + ((!g4944) & (g2360) & (!g2364) & (g2405)) + ((!g4944) & (g2360) & (g2364) & (!g2405)) + ((g4944) & (!g2360) & (!g2364) & (g2405)) + ((g4944) & (!g2360) & (g2364) & (!g2405)) + ((g4944) & (g2360) & (!g2364) & (!g2405)) + ((g4944) & (g2360) & (g2364) & (!g2405)));
	assign g6232 = (((!g4944) & (!g2360) & (!g2364) & (!g2405)) + ((!g4944) & (!g2360) & (g2364) & (!g2405)) + ((!g4944) & (g2360) & (!g2364) & (!g2405)) + ((!g4944) & (g2360) & (g2364) & (g2405)) + ((g4944) & (!g2360) & (!g2364) & (!g2405)) + ((g4944) & (!g2360) & (g2364) & (g2405)) + ((g4944) & (g2360) & (!g2364) & (g2405)) + ((g4944) & (g2360) & (g2364) & (g2405)));
	assign g6233 = (((!g6234) & (!g6235)));
	assign g6234 = (((!g2002) & (g6236)));
	assign g6235 = (((g2002) & (g6239)));
	assign g6236 = (((!g6237) & (!g6238)));
	assign g6237 = (((!g1914) & (g6242)));
	assign g6238 = (((g1914) & (g5005)));
	assign g6239 = (((!g6240) & (!g6241)));
	assign g6240 = (((!g1914) & (g6243)));
	assign g6241 = (((g1914) & (g5005)));
	assign g6242 = (((!g1132) & (!g1999) & (!g4936) & (g1165)) + ((!g1132) & (!g1999) & (g4936) & (g1165)) + ((!g1132) & (g1999) & (!g4936) & (g1165)) + ((!g1132) & (g1999) & (g4936) & (!g1165)) + ((g1132) & (!g1999) & (!g4936) & (g1165)) + ((g1132) & (!g1999) & (g4936) & (!g1165)) + ((g1132) & (g1999) & (!g4936) & (!g1165)) + ((g1132) & (g1999) & (g4936) & (!g1165)));
	assign g6243 = (((!g1132) & (!g1999) & (!g4936) & (!g1165)) + ((!g1132) & (!g1999) & (g4936) & (!g1165)) + ((!g1132) & (g1999) & (!g4936) & (!g1165)) + ((!g1132) & (g1999) & (g4936) & (g1165)) + ((g1132) & (!g1999) & (!g4936) & (!g1165)) + ((g1132) & (!g1999) & (g4936) & (g1165)) + ((g1132) & (g1999) & (!g4936) & (g1165)) + ((g1132) & (g1999) & (g4936) & (g1165)));
	assign g6244 = (((!g6245) & (!g6246)));
	assign g6245 = (((!g2390) & (g6247)));
	assign g6246 = (((g2390) & (g6250)));
	assign g6247 = (((!g6248) & (!g6249)));
	assign g6248 = (((!g1914) & (g5002)));
	assign g6249 = (((g1914) & (g6253)));
	assign g6250 = (((!g6251) & (!g6252)));
	assign g6251 = (((!g1914) & (g5002)));
	assign g6252 = (((g1914) & (g6254)));
	assign g6253 = (((!g2356) & (!g2354) & (!g4968) & (g2402)) + ((!g2356) & (!g2354) & (g4968) & (g2402)) + ((!g2356) & (g2354) & (!g4968) & (g2402)) + ((!g2356) & (g2354) & (g4968) & (!g2402)) + ((g2356) & (!g2354) & (!g4968) & (g2402)) + ((g2356) & (!g2354) & (g4968) & (!g2402)) + ((g2356) & (g2354) & (!g4968) & (!g2402)) + ((g2356) & (g2354) & (g4968) & (!g2402)));
	assign g6254 = (((!g2356) & (!g2354) & (!g4968) & (!g2402)) + ((!g2356) & (!g2354) & (g4968) & (!g2402)) + ((!g2356) & (g2354) & (!g4968) & (!g2402)) + ((!g2356) & (g2354) & (g4968) & (g2402)) + ((g2356) & (!g2354) & (!g4968) & (!g2402)) + ((g2356) & (!g2354) & (g4968) & (g2402)) + ((g2356) & (g2354) & (!g4968) & (g2402)) + ((g2356) & (g2354) & (g4968) & (g2402)));
	assign g6255 = (((!g6256) & (!g6257)));
	assign g6256 = (((!g2399) & (g6258)));
	assign g6257 = (((g2399) & (g6261)));
	assign g6258 = (((!g6259) & (!g6260)));
	assign g6259 = (((!g1914) & (g6264)));
	assign g6260 = (((g1914) & (g4998)));
	assign g6261 = (((!g6262) & (!g6263)));
	assign g6262 = (((!g1914) & (g6265)));
	assign g6263 = (((g1914) & (g4998)));
	assign g6264 = (((!g2364) & (!g2350) & (!g4956) & (g2405)) + ((!g2364) & (!g2350) & (g4956) & (g2405)) + ((!g2364) & (g2350) & (!g4956) & (g2405)) + ((!g2364) & (g2350) & (g4956) & (!g2405)) + ((g2364) & (!g2350) & (!g4956) & (g2405)) + ((g2364) & (!g2350) & (g4956) & (!g2405)) + ((g2364) & (g2350) & (!g4956) & (!g2405)) + ((g2364) & (g2350) & (g4956) & (!g2405)));
	assign g6265 = (((!g2364) & (!g2350) & (!g4956) & (!g2405)) + ((!g2364) & (!g2350) & (g4956) & (!g2405)) + ((!g2364) & (g2350) & (!g4956) & (!g2405)) + ((!g2364) & (g2350) & (g4956) & (g2405)) + ((g2364) & (!g2350) & (!g4956) & (!g2405)) + ((g2364) & (!g2350) & (g4956) & (g2405)) + ((g2364) & (g2350) & (!g4956) & (g2405)) + ((g2364) & (g2350) & (g4956) & (g2405)));
	assign g6266 = (((g830) & (!g6267)));
	assign g6267 = (((g830) & (g6268)));
	assign g6268 = (((!g6269) & (!g6270)));
	assign g6269 = (((!g1914) & (g6271)));
	assign g6270 = (((g1914) & (g6272)));
	assign g6271 = (((!g3378) & (!g2789) & (!g4996) & (g2768)) + ((!g3378) & (!g2789) & (g4996) & (!g2768)) + ((!g3378) & (g2789) & (!g4996) & (!g2768)) + ((!g3378) & (g2789) & (g4996) & (g2768)) + ((g3378) & (!g2789) & (!g4996) & (!g2768)) + ((g3378) & (!g2789) & (g4996) & (g2768)) + ((g3378) & (g2789) & (!g4996) & (g2768)) + ((g3378) & (g2789) & (g4996) & (!g2768)));
	assign g6272 = (((!g4995) & (g2768)) + ((g4995) & (!g2768)));
	assign g6273 = (((!g6274) & (!g6275)));
	assign g6274 = (((!g1963) & (g6276)));
	assign g6275 = (((g1963) & (g6279)));
	assign g6276 = (((!g6277) & (!g6278)));
	assign g6277 = (((!g1914) & (g4993)));
	assign g6278 = (((g1914) & (g6282)));
	assign g6279 = (((!g6280) & (!g6281)));
	assign g6280 = (((!g1914) & (g4993)));
	assign g6281 = (((g1914) & (g6283)));
	assign g6282 = (((!g1132) & (!g1961) & (!g4952) & (g1165)) + ((!g1132) & (!g1961) & (g4952) & (g1165)) + ((!g1132) & (g1961) & (!g4952) & (g1165)) + ((!g1132) & (g1961) & (g4952) & (!g1165)) + ((g1132) & (!g1961) & (!g4952) & (g1165)) + ((g1132) & (!g1961) & (g4952) & (!g1165)) + ((g1132) & (g1961) & (!g4952) & (!g1165)) + ((g1132) & (g1961) & (g4952) & (!g1165)));
	assign g6283 = (((!g1132) & (!g1961) & (!g4952) & (!g1165)) + ((!g1132) & (!g1961) & (g4952) & (!g1165)) + ((!g1132) & (g1961) & (!g4952) & (!g1165)) + ((!g1132) & (g1961) & (g4952) & (g1165)) + ((g1132) & (!g1961) & (!g4952) & (!g1165)) + ((g1132) & (!g1961) & (g4952) & (g1165)) + ((g1132) & (g1961) & (!g4952) & (g1165)) + ((g1132) & (g1961) & (g4952) & (g1165)));
	assign g6284 = (((!g6285) & (!g6286)));
	assign g6285 = (((!g1540) & (g6287)));
	assign g6286 = (((g1540) & (g6290)));
	assign g6287 = (((!g6288) & (!g6289)));
	assign g6288 = (((!g1914) & (g6293)));
	assign g6289 = (((g1914) & (g6294)));
	assign g6290 = (((!g6291) & (!g6292)));
	assign g6291 = (((!g1914) & (g6295)));
	assign g6292 = (((g1914) & (g6296)));
	assign g6293 = (((!g2950) & (g4985)) + ((g2950) & (!g4985)));
	assign g6294 = (((!g2932) & (!g4986) & (g2944)) + ((!g2932) & (g4986) & (!g2944)) + ((g2932) & (!g4986) & (!g2944)) + ((g2932) & (g4986) & (g2944)));
	assign g6295 = (((!g2950) & (!g4985)) + ((g2950) & (g4985)));
	assign g6296 = (((!g2932) & (!g4986) & (g2944)) + ((!g2932) & (g4986) & (!g2944)) + ((g2932) & (!g4986) & (!g2944)) + ((g2932) & (g4986) & (g2944)));
	assign g6297 = (((!g6298) & (!g6299)));
	assign g6298 = (((!g3018) & (g6300)));
	assign g6299 = (((g3018) & (g6303)));
	assign g6300 = (((!g6301) & (!g6302)));
	assign g6301 = (((!g1914) & (g6306)));
	assign g6302 = (((g1914) & (g6307)));
	assign g6303 = (((!g6304) & (!g6305)));
	assign g6304 = (((!g1914) & (g6308)));
	assign g6305 = (((g1914) & (g6309)));
	assign g6306 = (((!g4927) & (g3022)) + ((g4927) & (!g3022)));
	assign g6307 = (((!g2718) & (!g2098) & (g4928)) + ((!g2718) & (g2098) & (!g4928)) + ((g2718) & (!g2098) & (!g4928)) + ((g2718) & (g2098) & (g4928)));
	assign g6308 = (((!g4927) & (!g3022)) + ((g4927) & (g3022)));
	assign g6309 = (((!g2718) & (!g2098) & (g4928)) + ((!g2718) & (g2098) & (!g4928)) + ((g2718) & (!g2098) & (!g4928)) + ((g2718) & (g2098) & (g4928)));
	assign g6310 = (((!g6311) & (!g6312)));
	assign g6311 = (((!g4933) & (g6313)));
	assign g6312 = (((g4933) & (g6316)));
	assign g6313 = (((!g6314) & (!g6315)));
	assign g6314 = (((!g1914) & (g6319)));
	assign g6315 = (((g1914) & (g6320)));
	assign g6316 = (((!g6317) & (!g6318)));
	assign g6317 = (((!g1914) & (g6321)));
	assign g6318 = (((g1914) & (g6322)));
	assign g6319 = (((!g2690) & (!g2100) & (g4934)) + ((!g2690) & (g2100) & (!g4934)) + ((g2690) & (!g2100) & (!g4934)) + ((g2690) & (g2100) & (g4934)));
	assign g6320 = (((!g3022) & (g3007)) + ((g3022) & (!g3007)));
	assign g6321 = (((!g2690) & (!g2100) & (g4934)) + ((!g2690) & (g2100) & (!g4934)) + ((g2690) & (!g2100) & (!g4934)) + ((g2690) & (g2100) & (g4934)));
	assign g6322 = (((!g3022) & (!g3007)) + ((g3022) & (g3007)));
	assign g6323 = (((!g6324) & (!g6325)));
	assign g6324 = (((!g1507) & (g6326)));
	assign g6325 = (((g1507) & (g6329)));
	assign g6326 = (((!g6327) & (!g6328)));
	assign g6327 = (((!g1914) & (g6332)));
	assign g6328 = (((g1914) & (g4930)));
	assign g6329 = (((!g6330) & (!g6331)));
	assign g6330 = (((!g1914) & (g6333)));
	assign g6331 = (((g1914) & (g4930)));
	assign g6332 = (((!g4873) & (!g1473) & (!g2854) & (g2881)) + ((!g4873) & (!g1473) & (g2854) & (g2881)) + ((!g4873) & (g1473) & (!g2854) & (g2881)) + ((!g4873) & (g1473) & (g2854) & (!g2881)) + ((g4873) & (!g1473) & (!g2854) & (g2881)) + ((g4873) & (!g1473) & (g2854) & (!g2881)) + ((g4873) & (g1473) & (!g2854) & (!g2881)) + ((g4873) & (g1473) & (g2854) & (!g2881)));
	assign g6333 = (((!g4873) & (!g1473) & (!g2854) & (!g2881)) + ((!g4873) & (!g1473) & (g2854) & (!g2881)) + ((!g4873) & (g1473) & (!g2854) & (!g2881)) + ((!g4873) & (g1473) & (g2854) & (g2881)) + ((g4873) & (!g1473) & (!g2854) & (!g2881)) + ((g4873) & (!g1473) & (g2854) & (g2881)) + ((g4873) & (g1473) & (!g2854) & (g2881)) + ((g4873) & (g1473) & (g2854) & (g2881)));
	assign g6334 = (((g830) & (!g6335)));
	assign g6335 = (((g830) & (g6336)));
	assign g6336 = (((!g6337) & (!g6338)));
	assign g6337 = (((!g1914) & (g6339)));
	assign g6338 = (((g1914) & (g6340)));
	assign g6339 = (((!g4863) & (g2643)) + ((g4863) & (!g2643)));
	assign g6340 = (((!g4862) & (!g3265) & (!g3245) & (g2643)) + ((!g4862) & (!g3265) & (g3245) & (!g2643)) + ((!g4862) & (g3265) & (!g3245) & (!g2643)) + ((!g4862) & (g3265) & (g3245) & (g2643)) + ((g4862) & (!g3265) & (!g3245) & (!g2643)) + ((g4862) & (!g3265) & (g3245) & (g2643)) + ((g4862) & (g3265) & (!g3245) & (g2643)) + ((g4862) & (g3265) & (g3245) & (!g2643)));
	assign g6341 = (((!g6342) & (!g6343)));
	assign g6342 = (((!g2271) & (g6344)));
	assign g6343 = (((g2271) & (g6347)));
	assign g6344 = (((!g6345) & (!g6346)));
	assign g6345 = (((!g1914) & (g4857)));
	assign g6346 = (((g1914) & (g6350)));
	assign g6347 = (((!g6348) & (!g6349)));
	assign g6348 = (((!g1914) & (g4857)));
	assign g6349 = (((g1914) & (g6351)));
	assign g6350 = (((!g2236) & (!g2224) & (!g4800) & (g2273)) + ((!g2236) & (!g2224) & (g4800) & (g2273)) + ((!g2236) & (g2224) & (!g4800) & (g2273)) + ((!g2236) & (g2224) & (g4800) & (!g2273)) + ((g2236) & (!g2224) & (!g4800) & (g2273)) + ((g2236) & (!g2224) & (g4800) & (!g2273)) + ((g2236) & (g2224) & (!g4800) & (!g2273)) + ((g2236) & (g2224) & (g4800) & (!g2273)));
	assign g6351 = (((!g2236) & (!g2224) & (!g4800) & (!g2273)) + ((!g2236) & (!g2224) & (g4800) & (!g2273)) + ((!g2236) & (g2224) & (!g4800) & (!g2273)) + ((!g2236) & (g2224) & (g4800) & (g2273)) + ((g2236) & (!g2224) & (!g4800) & (!g2273)) + ((g2236) & (!g2224) & (g4800) & (g2273)) + ((g2236) & (g2224) & (!g4800) & (g2273)) + ((g2236) & (g2224) & (g4800) & (g2273)));
	assign g6352 = (((g830) & (!g6353)));
	assign g6353 = (((g830) & (g6354)));
	assign g6354 = (((!g6355) & (!g6356)));
	assign g6355 = (((!g1914) & (g6357)));
	assign g6356 = (((g1914) & (g6358)));
	assign g6357 = (((!g4853) & (g2629)) + ((g4853) & (!g2629)));
	assign g6358 = (((!g4852) & (!g3279) & (!g3222) & (g2629)) + ((!g4852) & (!g3279) & (g3222) & (!g2629)) + ((!g4852) & (g3279) & (!g3222) & (!g2629)) + ((!g4852) & (g3279) & (g3222) & (g2629)) + ((g4852) & (!g3279) & (!g3222) & (!g2629)) + ((g4852) & (!g3279) & (g3222) & (g2629)) + ((g4852) & (g3279) & (!g3222) & (g2629)) + ((g4852) & (g3279) & (g3222) & (!g2629)));
	assign g6359 = (((!g6360) & (!g6361)));
	assign g6360 = (((!g2267) & (g6362)));
	assign g6361 = (((g2267) & (g6365)));
	assign g6362 = (((!g6363) & (!g6364)));
	assign g6363 = (((!g1914) & (g6368)));
	assign g6364 = (((g1914) & (g4849)));
	assign g6365 = (((!g6366) & (!g6367)));
	assign g6366 = (((!g1914) & (g6369)));
	assign g6367 = (((g1914) & (g4849)));
	assign g6368 = (((!g2239) & (!g2233) & (!g4796) & (g2281)) + ((!g2239) & (!g2233) & (g4796) & (g2281)) + ((!g2239) & (g2233) & (!g4796) & (g2281)) + ((!g2239) & (g2233) & (g4796) & (!g2281)) + ((g2239) & (!g2233) & (!g4796) & (g2281)) + ((g2239) & (!g2233) & (g4796) & (!g2281)) + ((g2239) & (g2233) & (!g4796) & (!g2281)) + ((g2239) & (g2233) & (g4796) & (!g2281)));
	assign g6369 = (((!g2239) & (!g2233) & (!g4796) & (!g2281)) + ((!g2239) & (!g2233) & (g4796) & (!g2281)) + ((!g2239) & (g2233) & (!g4796) & (!g2281)) + ((!g2239) & (g2233) & (g4796) & (g2281)) + ((g2239) & (!g2233) & (!g4796) & (!g2281)) + ((g2239) & (!g2233) & (g4796) & (g2281)) + ((g2239) & (g2233) & (!g4796) & (g2281)) + ((g2239) & (g2233) & (g4796) & (g2281)));
	assign g6370 = (((!g6371) & (!g6372)));
	assign g6371 = (((!g1956) & (g6373)));
	assign g6372 = (((g1956) & (g6376)));
	assign g6373 = (((!g6374) & (!g6375)));
	assign g6374 = (((!g1914) & (g4847)));
	assign g6375 = (((g1914) & (g6379)));
	assign g6376 = (((!g6377) & (!g6378)));
	assign g6377 = (((!g1914) & (g4847)));
	assign g6378 = (((g1914) & (g6380)));
	assign g6379 = (((!g1031) & (!g1954) & (!g4790) & (g1065)) + ((!g1031) & (!g1954) & (g4790) & (g1065)) + ((!g1031) & (g1954) & (!g4790) & (g1065)) + ((!g1031) & (g1954) & (g4790) & (!g1065)) + ((g1031) & (!g1954) & (!g4790) & (g1065)) + ((g1031) & (!g1954) & (g4790) & (!g1065)) + ((g1031) & (g1954) & (!g4790) & (!g1065)) + ((g1031) & (g1954) & (g4790) & (!g1065)));
	assign g6380 = (((!g1031) & (!g1954) & (!g4790) & (!g1065)) + ((!g1031) & (!g1954) & (g4790) & (!g1065)) + ((!g1031) & (g1954) & (!g4790) & (!g1065)) + ((!g1031) & (g1954) & (g4790) & (g1065)) + ((g1031) & (!g1954) & (!g4790) & (!g1065)) + ((g1031) & (!g1954) & (g4790) & (g1065)) + ((g1031) & (g1954) & (!g4790) & (g1065)) + ((g1031) & (g1954) & (g4790) & (g1065)));
	assign g6381 = (((!g6382) & (!g6383)));
	assign g6382 = (((!g2271) & (g6384)));
	assign g6383 = (((g2271) & (g6387)));
	assign g6384 = (((!g6385) & (!g6386)));
	assign g6385 = (((!g1914) & (g6390)));
	assign g6386 = (((g1914) & (g4845)));
	assign g6387 = (((!g6388) & (!g6389)));
	assign g6388 = (((!g1914) & (g6391)));
	assign g6389 = (((g1914) & (g4845)));
	assign g6390 = (((!g2227) & (!g2224) & (!g4817) & (g2279)) + ((!g2227) & (!g2224) & (g4817) & (g2279)) + ((!g2227) & (g2224) & (!g4817) & (g2279)) + ((!g2227) & (g2224) & (g4817) & (!g2279)) + ((g2227) & (!g2224) & (!g4817) & (g2279)) + ((g2227) & (!g2224) & (g4817) & (!g2279)) + ((g2227) & (g2224) & (!g4817) & (!g2279)) + ((g2227) & (g2224) & (g4817) & (!g2279)));
	assign g6391 = (((!g2227) & (!g2224) & (!g4817) & (!g2279)) + ((!g2227) & (!g2224) & (g4817) & (!g2279)) + ((!g2227) & (g2224) & (!g4817) & (!g2279)) + ((!g2227) & (g2224) & (g4817) & (g2279)) + ((g2227) & (!g2224) & (!g4817) & (!g2279)) + ((g2227) & (!g2224) & (g4817) & (g2279)) + ((g2227) & (g2224) & (!g4817) & (g2279)) + ((g2227) & (g2224) & (g4817) & (g2279)));
	assign g6392 = (((!g6393) & (!g6394)));
	assign g6393 = (((!g2277) & (g6395)));
	assign g6394 = (((g2277) & (g6398)));
	assign g6395 = (((!g6396) & (!g6397)));
	assign g6396 = (((!g1914) & (g4843)));
	assign g6397 = (((g1914) & (g6401)));
	assign g6398 = (((!g6399) & (!g6400)));
	assign g6399 = (((!g1914) & (g4843)));
	assign g6400 = (((g1914) & (g6402)));
	assign g6401 = (((!g4806) & (!g2217) & (!g2239) & (g2281)) + ((!g4806) & (!g2217) & (g2239) & (g2281)) + ((!g4806) & (g2217) & (!g2239) & (g2281)) + ((!g4806) & (g2217) & (g2239) & (!g2281)) + ((g4806) & (!g2217) & (!g2239) & (g2281)) + ((g4806) & (!g2217) & (g2239) & (!g2281)) + ((g4806) & (g2217) & (!g2239) & (!g2281)) + ((g4806) & (g2217) & (g2239) & (!g2281)));
	assign g6402 = (((!g4806) & (!g2217) & (!g2239) & (!g2281)) + ((!g4806) & (!g2217) & (g2239) & (!g2281)) + ((!g4806) & (g2217) & (!g2239) & (!g2281)) + ((!g4806) & (g2217) & (g2239) & (g2281)) + ((g4806) & (!g2217) & (!g2239) & (!g2281)) + ((g4806) & (!g2217) & (g2239) & (g2281)) + ((g4806) & (g2217) & (!g2239) & (g2281)) + ((g4806) & (g2217) & (g2239) & (g2281)));
	assign g6403 = (((g830) & (g6404)));
	assign g6404 = (((!g6405) & (!g6406)));
	assign g6405 = (((!g1914) & (g6407)));
	assign g6406 = (((g1914) & (g6408)));
	assign g6407 = (((!g4842) & (g2614)) + ((g4842) & (!g2614)));
	assign g6408 = (((!g4841) & (!g3255) & (!g2649) & (g2614)) + ((!g4841) & (!g3255) & (g2649) & (!g2614)) + ((!g4841) & (g3255) & (!g2649) & (!g2614)) + ((!g4841) & (g3255) & (g2649) & (g2614)) + ((g4841) & (!g3255) & (!g2649) & (!g2614)) + ((g4841) & (!g3255) & (g2649) & (g2614)) + ((g4841) & (g3255) & (!g2649) & (g2614)) + ((g4841) & (g3255) & (g2649) & (!g2614)));
	assign g6409 = (((!g6410) & (!g6411)));
	assign g6410 = (((!g1994) & (g6412)));
	assign g6411 = (((g1994) & (g6415)));
	assign g6412 = (((!g6413) & (!g6414)));
	assign g6413 = (((!g1914) & (g6418)));
	assign g6414 = (((g1914) & (g4839)));
	assign g6415 = (((!g6416) & (!g6417)));
	assign g6416 = (((!g1914) & (g6419)));
	assign g6417 = (((g1914) & (g4839)));
	assign g6418 = (((!g1031) & (!g1992) & (!g4803) & (g1065)) + ((!g1031) & (!g1992) & (g4803) & (g1065)) + ((!g1031) & (g1992) & (!g4803) & (g1065)) + ((!g1031) & (g1992) & (g4803) & (!g1065)) + ((g1031) & (!g1992) & (!g4803) & (g1065)) + ((g1031) & (!g1992) & (g4803) & (!g1065)) + ((g1031) & (g1992) & (!g4803) & (!g1065)) + ((g1031) & (g1992) & (g4803) & (!g1065)));
	assign g6419 = (((!g1031) & (!g1992) & (!g4803) & (!g1065)) + ((!g1031) & (!g1992) & (g4803) & (!g1065)) + ((!g1031) & (g1992) & (!g4803) & (!g1065)) + ((!g1031) & (g1992) & (g4803) & (g1065)) + ((g1031) & (!g1992) & (!g4803) & (!g1065)) + ((g1031) & (!g1992) & (g4803) & (g1065)) + ((g1031) & (g1992) & (!g4803) & (g1065)) + ((g1031) & (g1992) & (g4803) & (g1065)));
	assign g6420 = (((!g6421) & (!g6422)));
	assign g6421 = (((!g2889) & (g6423)));
	assign g6422 = (((g2889) & (g6426)));
	assign g6423 = (((!g6424) & (!g6425)));
	assign g6424 = (((!g1914) & (g4837)));
	assign g6425 = (((g1914) & (g6429)));
	assign g6426 = (((!g6427) & (!g6428)));
	assign g6427 = (((!g1914) & (g4837)));
	assign g6428 = (((g1914) & (g6430)));
	assign g6429 = (((!g2868) & (!g4786) & (!g2874) & (g2904)) + ((!g2868) & (!g4786) & (g2874) & (g2904)) + ((!g2868) & (g4786) & (!g2874) & (g2904)) + ((!g2868) & (g4786) & (g2874) & (!g2904)) + ((g2868) & (!g4786) & (!g2874) & (g2904)) + ((g2868) & (!g4786) & (g2874) & (!g2904)) + ((g2868) & (g4786) & (!g2874) & (!g2904)) + ((g2868) & (g4786) & (g2874) & (!g2904)));
	assign g6430 = (((!g2868) & (!g4786) & (!g2874) & (!g2904)) + ((!g2868) & (!g4786) & (g2874) & (!g2904)) + ((!g2868) & (g4786) & (!g2874) & (!g2904)) + ((!g2868) & (g4786) & (g2874) & (g2904)) + ((g2868) & (!g4786) & (!g2874) & (!g2904)) + ((g2868) & (!g4786) & (g2874) & (g2904)) + ((g2868) & (g4786) & (!g2874) & (g2904)) + ((g2868) & (g4786) & (g2874) & (g2904)));
	assign g6431 = (((!g6432) & (!g6433)));
	assign g6432 = (((!g2900) & (g6434)));
	assign g6433 = (((g2900) & (g6437)));
	assign g6434 = (((!g6435) & (!g6436)));
	assign g6435 = (((!g1914) & (g6440)));
	assign g6436 = (((g1914) & (g4831)));
	assign g6437 = (((!g6438) & (!g6439)));
	assign g6438 = (((!g1914) & (g6441)));
	assign g6439 = (((g1914) & (g4831)));
	assign g6440 = (((!g2874) & (!g2851) & (!g4779) & (g2904)) + ((!g2874) & (!g2851) & (g4779) & (g2904)) + ((!g2874) & (g2851) & (!g4779) & (g2904)) + ((!g2874) & (g2851) & (g4779) & (!g2904)) + ((g2874) & (!g2851) & (!g4779) & (g2904)) + ((g2874) & (!g2851) & (g4779) & (!g2904)) + ((g2874) & (g2851) & (!g4779) & (!g2904)) + ((g2874) & (g2851) & (g4779) & (!g2904)));
	assign g6441 = (((!g2874) & (!g2851) & (!g4779) & (!g2904)) + ((!g2874) & (!g2851) & (g4779) & (!g2904)) + ((!g2874) & (g2851) & (!g4779) & (!g2904)) + ((!g2874) & (g2851) & (g4779) & (g2904)) + ((g2874) & (!g2851) & (!g4779) & (!g2904)) + ((g2874) & (!g2851) & (g4779) & (g2904)) + ((g2874) & (g2851) & (!g4779) & (g2904)) + ((g2874) & (g2851) & (g4779) & (g2904)));
	assign g6442 = (((!g6443) & (!g6444)));
	assign g6443 = (((!g1406) & (g6445)));
	assign g6444 = (((g1406) & (g6448)));
	assign g6445 = (((!g6446) & (!g6447)));
	assign g6446 = (((!g1914) & (g6451)));
	assign g6447 = (((g1914) & (g4783)));
	assign g6448 = (((!g6449) & (!g6450)));
	assign g6449 = (((!g1914) & (g6452)));
	assign g6450 = (((g1914) & (g4783)));
	assign g6451 = (((!g4747) & (!g1370) & (!g2690) & (g2774)) + ((!g4747) & (!g1370) & (g2690) & (g2774)) + ((!g4747) & (g1370) & (!g2690) & (g2774)) + ((!g4747) & (g1370) & (g2690) & (!g2774)) + ((g4747) & (!g1370) & (!g2690) & (g2774)) + ((g4747) & (!g1370) & (g2690) & (!g2774)) + ((g4747) & (g1370) & (!g2690) & (!g2774)) + ((g4747) & (g1370) & (g2690) & (!g2774)));
	assign g6452 = (((!g4747) & (!g1370) & (!g2690) & (!g2774)) + ((!g4747) & (!g1370) & (g2690) & (!g2774)) + ((!g4747) & (g1370) & (!g2690) & (!g2774)) + ((!g4747) & (g1370) & (g2690) & (g2774)) + ((g4747) & (!g1370) & (!g2690) & (!g2774)) + ((g4747) & (!g1370) & (g2690) & (g2774)) + ((g4747) & (g1370) & (!g2690) & (g2774)) + ((g4747) & (g1370) & (g2690) & (g2774)));
	assign g6453 = (((g830) & (g6454)));
	assign g6454 = (((!g6455) & (!g6456)));
	assign g6455 = (((!g1914) & (g6457)));
	assign g6456 = (((g1914) & (g6458)));
	assign g6457 = (((!g4775) & (!g3170) & (!g3168) & (g2546)) + ((!g4775) & (!g3170) & (g3168) & (!g2546)) + ((!g4775) & (g3170) & (!g3168) & (!g2546)) + ((!g4775) & (g3170) & (g3168) & (g2546)) + ((g4775) & (!g3170) & (!g3168) & (!g2546)) + ((g4775) & (!g3170) & (g3168) & (g2546)) + ((g4775) & (g3170) & (!g3168) & (g2546)) + ((g4775) & (g3170) & (g3168) & (!g2546)));
	assign g6458 = (((!g4774) & (g2546)) + ((g4774) & (!g2546)));
	assign g6459 = (((!g6460) & (!g6461)));
	assign g6460 = (((!g1914) & (g6462)));
	assign g6461 = (((g1914) & (g6465)));
	assign g6462 = (((!g6463) & (!g6464)));
	assign g6463 = (((!g830) & (key[140])));
	assign g6464 = (((g830) & (g6468)));
	assign g6465 = (((!g6466) & (!g6467)));
	assign g6466 = (((!g830) & (key[140])));
	assign g6467 = (((g830) & (g5709)));
	assign g6468 = (((!g5709) & (!g4712) & (!g3356) & (!g2759)) + ((!g5709) & (!g4712) & (!g3356) & (g2759)) + ((!g5709) & (!g4712) & (g3356) & (!g2759)) + ((!g5709) & (g4712) & (!g3356) & (!g2759)) + ((g5709) & (!g4712) & (g3356) & (g2759)) + ((g5709) & (g4712) & (!g3356) & (g2759)) + ((g5709) & (g4712) & (g3356) & (!g2759)) + ((g5709) & (g4712) & (g3356) & (g2759)));
	assign g6469 = (((g830) & (g6470)));
	assign g6470 = (((!g6471) & (!g6472)));
	assign g6471 = (((!g1914) & (g6473)));
	assign g6472 = (((g1914) & (g6474)));
	assign g6473 = (((!g4764) & (!g3165) & (!g3159) & (g2537)) + ((!g4764) & (!g3165) & (g3159) & (!g2537)) + ((!g4764) & (g3165) & (!g3159) & (!g2537)) + ((!g4764) & (g3165) & (g3159) & (g2537)) + ((g4764) & (!g3165) & (!g3159) & (!g2537)) + ((g4764) & (!g3165) & (g3159) & (g2537)) + ((g4764) & (g3165) & (!g3159) & (g2537)) + ((g4764) & (g3165) & (g3159) & (!g2537)));
	assign g6474 = (((!g4763) & (g2537)) + ((g4763) & (!g2537)));
	assign g6475 = (((!g6476) & (!g6477)));
	assign g6476 = (((!g1914) & (g6478)));
	assign g6477 = (((g1914) & (g6481)));
	assign g6478 = (((!g6479) & (!g6480)));
	assign g6479 = (((!g830) & (g4759)));
	assign g6480 = (((g830) & (g5705)));
	assign g6481 = (((!g6482) & (!g6483)));
	assign g6482 = (((!g830) & (g4759)));
	assign g6483 = (((g830) & (g6484)));
	assign g6484 = (((!g5705) & (!g4707) & (!g3353) & (!g2760)) + ((!g5705) & (!g4707) & (!g3353) & (g2760)) + ((!g5705) & (!g4707) & (g3353) & (!g2760)) + ((!g5705) & (g4707) & (!g3353) & (!g2760)) + ((g5705) & (!g4707) & (g3353) & (g2760)) + ((g5705) & (g4707) & (!g3353) & (g2760)) + ((g5705) & (g4707) & (g3353) & (!g2760)) + ((g5705) & (g4707) & (g3353) & (g2760)));
	assign g6485 = (((!g6486) & (!g6487)));
	assign g6486 = (((!g1914) & (g6488)));
	assign g6487 = (((g1914) & (g6491)));
	assign g6488 = (((!g6489) & (!g6490)));
	assign g6489 = (((!g830) & (key[12])));
	assign g6490 = (((g830) & (g6494)));
	assign g6491 = (((!g6492) & (!g6493)));
	assign g6492 = (((!g830) & (key[12])));
	assign g6493 = (((g830) & (g5703)));
	assign g6494 = (((!g5703) & (!g4702) & (!g3348) & (!g3342)) + ((!g5703) & (!g4702) & (!g3348) & (g3342)) + ((!g5703) & (!g4702) & (g3348) & (!g3342)) + ((!g5703) & (g4702) & (!g3348) & (!g3342)) + ((g5703) & (!g4702) & (g3348) & (g3342)) + ((g5703) & (g4702) & (!g3348) & (g3342)) + ((g5703) & (g4702) & (g3348) & (!g3342)) + ((g5703) & (g4702) & (g3348) & (g3342)));
	assign g6495 = (((!g6496) & (!g6497)));
	assign g6496 = (((!g1914) & (g6498)));
	assign g6497 = (((g1914) & (g6501)));
	assign g6498 = (((!g6499) & (!g6500)));
	assign g6499 = (((!g830) & (key[236])));
	assign g6500 = (((g830) & (g5701)));
	assign g6501 = (((!g6502) & (!g6503)));
	assign g6502 = (((!g830) & (key[236])));
	assign g6503 = (((g830) & (g6504)));
	assign g6504 = (((!g5701) & (!g4728) & (!g3348) & (!g2761)) + ((!g5701) & (!g4728) & (!g3348) & (g2761)) + ((!g5701) & (!g4728) & (g3348) & (!g2761)) + ((!g5701) & (g4728) & (!g3348) & (!g2761)) + ((g5701) & (!g4728) & (g3348) & (g2761)) + ((g5701) & (g4728) & (!g3348) & (g2761)) + ((g5701) & (g4728) & (g3348) & (!g2761)) + ((g5701) & (g4728) & (g3348) & (g2761)));
	assign g6505 = (((!g6506) & (!g6507)));
	assign g6506 = (((!g1914) & (g6508)));
	assign g6507 = (((g1914) & (g6511)));
	assign g6508 = (((!g6509) & (!g6510)));
	assign g6509 = (((!g830) & (nonce[12])));
	assign g6510 = (((g830) & (g6514)));
	assign g6511 = (((!g6512) & (!g6513)));
	assign g6512 = (((!g830) & (nonce[12])));
	assign g6513 = (((g830) & (g5699)));
	assign g6514 = (((!g5699) & (!g4718) & (!g3336) & (!g2758)) + ((!g5699) & (!g4718) & (!g3336) & (g2758)) + ((!g5699) & (!g4718) & (g3336) & (!g2758)) + ((!g5699) & (g4718) & (!g3336) & (!g2758)) + ((g5699) & (!g4718) & (g3336) & (g2758)) + ((g5699) & (g4718) & (!g3336) & (g2758)) + ((g5699) & (g4718) & (g3336) & (!g2758)) + ((g5699) & (g4718) & (g3336) & (g2758)));
	assign g6515 = (((g830) & (g6516)));
	assign g6516 = (((!g6517) & (!g6518)));
	assign g6517 = (((!g1914) & (g6519)));
	assign g6518 = (((g1914) & (g6520)));
	assign g6519 = (((!g4758) & (!g3155) & (!g2551) & (g2527)) + ((!g4758) & (!g3155) & (g2551) & (!g2527)) + ((!g4758) & (g3155) & (!g2551) & (!g2527)) + ((!g4758) & (g3155) & (g2551) & (g2527)) + ((g4758) & (!g3155) & (!g2551) & (!g2527)) + ((g4758) & (!g3155) & (g2551) & (g2527)) + ((g4758) & (g3155) & (!g2551) & (g2527)) + ((g4758) & (g3155) & (g2551) & (!g2527)));
	assign g6520 = (((!g4757) & (g2527)) + ((g4757) & (!g2527)));
	assign g6521 = (((!g6522) & (!g6523)));
	assign g6522 = (((!g1914) & (g6524)));
	assign g6523 = (((g1914) & (g6527)));
	assign g6524 = (((!g6525) & (!g6526)));
	assign g6525 = (((!g830) & (key[108])));
	assign g6526 = (((g830) & (g5695)));
	assign g6527 = (((!g6528) & (!g6529)));
	assign g6528 = (((!g830) & (key[108])));
	assign g6529 = (((g830) & (g6530)));
	assign g6530 = (((!g5695) & (!g4714) & (!g3356) & (!g3333)) + ((!g5695) & (!g4714) & (!g3356) & (g3333)) + ((!g5695) & (!g4714) & (g3356) & (!g3333)) + ((!g5695) & (g4714) & (!g3356) & (!g3333)) + ((g5695) & (!g4714) & (g3356) & (g3333)) + ((g5695) & (g4714) & (!g3356) & (g3333)) + ((g5695) & (g4714) & (g3356) & (!g3333)) + ((g5695) & (g4714) & (g3356) & (g3333)));
	assign g6531 = (((!g6532) & (!g6533)));
	assign g6532 = (((!g1370) & (g6534)));
	assign g6533 = (((g1370) & (g6537)));
	assign g6534 = (((!g6535) & (!g6536)));
	assign g6535 = (((!g1914) & (g6540)));
	assign g6536 = (((g1914) & (g6541)));
	assign g6537 = (((!g6538) & (!g6539)));
	assign g6538 = (((!g1914) & (g6542)));
	assign g6539 = (((g1914) & (g6543)));
	assign g6540 = (((!g2690) & (g4747)) + ((g2690) & (!g4747)));
	assign g6541 = (((!g2703) & (!g4748) & (g2742)) + ((!g2703) & (g4748) & (!g2742)) + ((g2703) & (!g4748) & (!g2742)) + ((g2703) & (g4748) & (g2742)));
	assign g6542 = (((!g2690) & (!g4747)) + ((g2690) & (g4747)));
	assign g6543 = (((!g2703) & (!g4748) & (g2742)) + ((!g2703) & (g4748) & (!g2742)) + ((g2703) & (!g4748) & (!g2742)) + ((g2703) & (g4748) & (g2742)));
	assign g6544 = (((!g6545) & (!g6546)));
	assign g6545 = (((!g2783) & (g6547)));
	assign g6546 = (((g2783) & (g6550)));
	assign g6547 = (((!g6548) & (!g6549)));
	assign g6548 = (((!g1914) & (g4699)));
	assign g6549 = (((g1914) & (g6553)));
	assign g6550 = (((!g6551) & (!g6552)));
	assign g6551 = (((!g1914) & (g4699)));
	assign g6552 = (((g1914) & (g6554)));
	assign g6553 = (((!g2713) & (!g4651) & (!g2752) & (g2787)) + ((!g2713) & (!g4651) & (g2752) & (g2787)) + ((!g2713) & (g4651) & (!g2752) & (g2787)) + ((!g2713) & (g4651) & (g2752) & (!g2787)) + ((g2713) & (!g4651) & (!g2752) & (g2787)) + ((g2713) & (!g4651) & (g2752) & (!g2787)) + ((g2713) & (g4651) & (!g2752) & (!g2787)) + ((g2713) & (g4651) & (g2752) & (!g2787)));
	assign g6554 = (((!g2713) & (!g4651) & (!g2752) & (!g2787)) + ((!g2713) & (!g4651) & (g2752) & (!g2787)) + ((!g2713) & (g4651) & (!g2752) & (!g2787)) + ((!g2713) & (g4651) & (g2752) & (g2787)) + ((g2713) & (!g4651) & (!g2752) & (!g2787)) + ((g2713) & (!g4651) & (g2752) & (g2787)) + ((g2713) & (g4651) & (!g2752) & (g2787)) + ((g2713) & (g4651) & (g2752) & (g2787)));
	assign g6555 = (((!g6556) & (!g6557)));
	assign g6556 = (((!g1337) & (g6558)));
	assign g6557 = (((g1337) & (g6561)));
	assign g6558 = (((!g6559) & (!g6560)));
	assign g6559 = (((!g1914) & (g6564)));
	assign g6560 = (((g1914) & (g4695)));
	assign g6561 = (((!g6562) & (!g6563)));
	assign g6562 = (((!g1914) & (g6565)));
	assign g6563 = (((g1914) & (g4695)));
	assign g6564 = (((!g4645) & (!g1303) & (!g2607) & (g2663)) + ((!g4645) & (!g1303) & (g2607) & (g2663)) + ((!g4645) & (g1303) & (!g2607) & (g2663)) + ((!g4645) & (g1303) & (g2607) & (!g2663)) + ((g4645) & (!g1303) & (!g2607) & (g2663)) + ((g4645) & (!g1303) & (g2607) & (!g2663)) + ((g4645) & (g1303) & (!g2607) & (!g2663)) + ((g4645) & (g1303) & (g2607) & (!g2663)));
	assign g6565 = (((!g4645) & (!g1303) & (!g2607) & (!g2663)) + ((!g4645) & (!g1303) & (g2607) & (!g2663)) + ((!g4645) & (g1303) & (!g2607) & (!g2663)) + ((!g4645) & (g1303) & (g2607) & (g2663)) + ((g4645) & (!g1303) & (!g2607) & (!g2663)) + ((g4645) & (!g1303) & (g2607) & (g2663)) + ((g4645) & (g1303) & (!g2607) & (g2663)) + ((g4645) & (g1303) & (g2607) & (g2663)));
	assign g6566 = (((!g6567) & (!g6568)));
	assign g6567 = (((!g2772) & (g6569)));
	assign g6568 = (((g2772) & (g6572)));
	assign g6569 = (((!g6570) & (!g6571)));
	assign g6570 = (((!g1914) & (g6575)));
	assign g6571 = (((g1914) & (g4693)));
	assign g6572 = (((!g6573) & (!g6574)));
	assign g6573 = (((!g1914) & (g6576)));
	assign g6574 = (((g1914) & (g4693)));
	assign g6575 = (((!g2752) & (!g2742) & (!g4641) & (g2787)) + ((!g2752) & (!g2742) & (g4641) & (g2787)) + ((!g2752) & (g2742) & (!g4641) & (g2787)) + ((!g2752) & (g2742) & (g4641) & (!g2787)) + ((g2752) & (!g2742) & (!g4641) & (g2787)) + ((g2752) & (!g2742) & (g4641) & (!g2787)) + ((g2752) & (g2742) & (!g4641) & (!g2787)) + ((g2752) & (g2742) & (g4641) & (!g2787)));
	assign g6576 = (((!g2752) & (!g2742) & (!g4641) & (!g2787)) + ((!g2752) & (!g2742) & (g4641) & (!g2787)) + ((!g2752) & (g2742) & (!g4641) & (!g2787)) + ((!g2752) & (g2742) & (g4641) & (g2787)) + ((g2752) & (!g2742) & (!g4641) & (!g2787)) + ((g2752) & (!g2742) & (g4641) & (g2787)) + ((g2752) & (g2742) & (!g4641) & (g2787)) + ((g2752) & (g2742) & (g4641) & (g2787)));
	assign g6577 = (((g830) & (!g6578)));
	assign g6578 = (((g830) & (g6579)));
	assign g6579 = (((!g6580) & (!g6581)));
	assign g6580 = (((!g1914) & (g6582)));
	assign g6581 = (((g1914) & (g6583)));
	assign g6582 = (((!g4688) & (g2419)) + ((g4688) & (!g2419)));
	assign g6583 = (((!g4686) & (!g3090) & (!g3082) & (g2419)) + ((!g4686) & (!g3090) & (g3082) & (!g2419)) + ((!g4686) & (g3090) & (!g3082) & (!g2419)) + ((!g4686) & (g3090) & (g3082) & (g2419)) + ((g4686) & (!g3090) & (!g3082) & (!g2419)) + ((g4686) & (!g3090) & (g3082) & (g2419)) + ((g4686) & (g3090) & (!g3082) & (g2419)) + ((g4686) & (g3090) & (g3082) & (!g2419)));
	assign g6584 = (((g830) & (!g6585)));
	assign g6585 = (((g830) & (g6586)));
	assign g6586 = (((!g6587) & (!g6588)));
	assign g6587 = (((!g1914) & (g6589)));
	assign g6588 = (((g1914) & (g6590)));
	assign g6589 = (((!g4676) & (g2405)) + ((g4676) & (!g2405)));
	assign g6590 = (((!g4674) & (!g3095) & (!g3074) & (g2405)) + ((!g4674) & (!g3095) & (g3074) & (!g2405)) + ((!g4674) & (g3095) & (!g3074) & (!g2405)) + ((!g4674) & (g3095) & (g3074) & (g2405)) + ((g4674) & (!g3095) & (!g3074) & (!g2405)) + ((g4674) & (!g3095) & (g3074) & (g2405)) + ((g4674) & (g3095) & (!g3074) & (g2405)) + ((g4674) & (g3095) & (g3074) & (!g2405)));
	assign g6591 = (((g830) & (!g6592)));
	assign g6592 = (((g830) & (g6593)));
	assign g6593 = (((!g6594) & (!g6595)));
	assign g6594 = (((!g1914) & (g6596)));
	assign g6595 = (((g1914) & (g6597)));
	assign g6596 = (((!g4660) & (g2390)) + ((g4660) & (!g2390)));
	assign g6597 = (((!g4658) & (!g3086) & (!g2426) & (g2390)) + ((!g4658) & (!g3086) & (g2426) & (!g2390)) + ((!g4658) & (g3086) & (!g2426) & (!g2390)) + ((!g4658) & (g3086) & (g2426) & (g2390)) + ((g4658) & (!g3086) & (!g2426) & (!g2390)) + ((g4658) & (!g3086) & (g2426) & (g2390)) + ((g4658) & (g3086) & (!g2426) & (g2390)) + ((g4658) & (g3086) & (g2426) & (!g2390)));
	assign g6598 = (((g830) & (g6599)));
	assign g6599 = (((!g6600) & (!g6601)));
	assign g6600 = (((!g1914) & (g6602)));
	assign g6601 = (((g1914) & (g6603)));
	assign g6602 = (((!g4635) & (g2373)) + ((g4635) & (!g2373)));
	assign g6603 = (((!g4634) & (!g3064) & (!g3061) & (g2373)) + ((!g4634) & (!g3064) & (g3061) & (!g2373)) + ((!g4634) & (g3064) & (!g3061) & (!g2373)) + ((!g4634) & (g3064) & (g3061) & (g2373)) + ((g4634) & (!g3064) & (!g3061) & (!g2373)) + ((g4634) & (!g3064) & (g3061) & (g2373)) + ((g4634) & (g3064) & (!g3061) & (g2373)) + ((g4634) & (g3064) & (g3061) & (!g2373)));
	assign g6604 = (((g830) & (g6605)));
	assign g6605 = (((!g6606) & (!g6607)));
	assign g6606 = (((!g1914) & (g6608)));
	assign g6607 = (((g1914) & (g6609)));
	assign g6608 = (((!g4625) & (g2364)) + ((g4625) & (!g2364)));
	assign g6609 = (((!g4624) & (!g3056) & (!g3047) & (g2364)) + ((!g4624) & (!g3056) & (g3047) & (!g2364)) + ((!g4624) & (g3056) & (!g3047) & (!g2364)) + ((!g4624) & (g3056) & (g3047) & (g2364)) + ((g4624) & (!g3056) & (!g3047) & (!g2364)) + ((g4624) & (!g3056) & (g3047) & (g2364)) + ((g4624) & (g3056) & (!g3047) & (g2364)) + ((g4624) & (g3056) & (g3047) & (!g2364)));
	assign g6610 = (((g830) & (g6611)));
	assign g6611 = (((!g6612) & (!g6613)));
	assign g6612 = (((!g1914) & (g6614)));
	assign g6613 = (((g1914) & (g6615)));
	assign g6614 = (((!g4606) & (g2354)) + ((g4606) & (!g2354)));
	assign g6615 = (((!g4605) & (!g3041) & (!g2378) & (g2354)) + ((!g4605) & (!g3041) & (g2378) & (!g2354)) + ((!g4605) & (g3041) & (!g2378) & (!g2354)) + ((!g4605) & (g3041) & (g2378) & (g2354)) + ((g4605) & (!g3041) & (!g2378) & (!g2354)) + ((g4605) & (!g3041) & (g2378) & (g2354)) + ((g4605) & (g3041) & (!g2378) & (g2354)) + ((g4605) & (g3041) & (g2378) & (!g2354)));
	assign g6616 = (((!g6617) & (!g6618)));
	assign g6617 = (((!g2672) & (g6619)));
	assign g6618 = (((g2672) & (g6622)));
	assign g6619 = (((!g6620) & (!g6621)));
	assign g6620 = (((!g1914) & (g4599)));
	assign g6621 = (((g1914) & (g6625)));
	assign g6622 = (((!g6623) & (!g6624)));
	assign g6623 = (((!g1914) & (g4599)));
	assign g6624 = (((g1914) & (g6626)));
	assign g6625 = (((!g2620) & (!g4547) & (!g2643) & (g2676)) + ((!g2620) & (!g4547) & (g2643) & (g2676)) + ((!g2620) & (g4547) & (!g2643) & (g2676)) + ((!g2620) & (g4547) & (g2643) & (!g2676)) + ((g2620) & (!g4547) & (!g2643) & (g2676)) + ((g2620) & (!g4547) & (g2643) & (!g2676)) + ((g2620) & (g4547) & (!g2643) & (!g2676)) + ((g2620) & (g4547) & (g2643) & (!g2676)));
	assign g6626 = (((!g2620) & (!g4547) & (!g2643) & (!g2676)) + ((!g2620) & (!g4547) & (g2643) & (!g2676)) + ((!g2620) & (g4547) & (!g2643) & (!g2676)) + ((!g2620) & (g4547) & (g2643) & (g2676)) + ((g2620) & (!g4547) & (!g2643) & (!g2676)) + ((g2620) & (!g4547) & (g2643) & (g2676)) + ((g2620) & (g4547) & (!g2643) & (g2676)) + ((g2620) & (g4547) & (g2643) & (g2676)));
	assign g6627 = (((!g6628) & (!g6629)));
	assign g6628 = (((!g2661) & (g6630)));
	assign g6629 = (((g2661) & (g6633)));
	assign g6630 = (((!g6631) & (!g6632)));
	assign g6631 = (((!g1914) & (g6636)));
	assign g6632 = (((g1914) & (g4592)));
	assign g6633 = (((!g6634) & (!g6635)));
	assign g6634 = (((!g1914) & (g6637)));
	assign g6635 = (((g1914) & (g4592)));
	assign g6636 = (((!g2643) & (!g2637) & (!g4539) & (g2676)) + ((!g2643) & (!g2637) & (g4539) & (g2676)) + ((!g2643) & (g2637) & (!g4539) & (g2676)) + ((!g2643) & (g2637) & (g4539) & (!g2676)) + ((g2643) & (!g2637) & (!g4539) & (g2676)) + ((g2643) & (!g2637) & (g4539) & (!g2676)) + ((g2643) & (g2637) & (!g4539) & (!g2676)) + ((g2643) & (g2637) & (g4539) & (!g2676)));
	assign g6637 = (((!g2643) & (!g2637) & (!g4539) & (!g2676)) + ((!g2643) & (!g2637) & (g4539) & (!g2676)) + ((!g2643) & (g2637) & (!g4539) & (!g2676)) + ((!g2643) & (g2637) & (g4539) & (g2676)) + ((g2643) & (!g2637) & (!g4539) & (!g2676)) + ((g2643) & (!g2637) & (g4539) & (g2676)) + ((g2643) & (g2637) & (!g4539) & (g2676)) + ((g2643) & (g2637) & (g4539) & (g2676)));
	assign g6638 = (((g830) & (!g6639)));
	assign g6639 = (((g830) & (g6640)));
	assign g6640 = (((!g6641) & (!g6642)));
	assign g6641 = (((!g1914) & (g6643)));
	assign g6642 = (((g1914) & (g6644)));
	assign g6643 = (((!g4587) & (!g3020) & (!g3018) & (g2340)) + ((!g4587) & (!g3020) & (g3018) & (!g2340)) + ((!g4587) & (g3020) & (!g3018) & (!g2340)) + ((!g4587) & (g3020) & (g3018) & (g2340)) + ((g4587) & (!g3020) & (!g3018) & (!g2340)) + ((g4587) & (!g3020) & (g3018) & (g2340)) + ((g4587) & (g3020) & (!g3018) & (g2340)) + ((g4587) & (g3020) & (g3018) & (!g2340)));
	assign g6644 = (((!g4586) & (g2340)) + ((g4586) & (!g2340)));
	assign g6645 = (((g830) & (g6646)));
	assign g6646 = (((!g6647) & (!g6648)));
	assign g6647 = (((!g1914) & (g6649)));
	assign g6648 = (((g1914) & (g6650)));
	assign g6649 = (((!g4575) & (!g3015) & (!g3009) & (g2326)) + ((!g4575) & (!g3015) & (g3009) & (!g2326)) + ((!g4575) & (g3015) & (!g3009) & (!g2326)) + ((!g4575) & (g3015) & (g3009) & (g2326)) + ((g4575) & (!g3015) & (!g3009) & (!g2326)) + ((g4575) & (!g3015) & (g3009) & (g2326)) + ((g4575) & (g3015) & (!g3009) & (g2326)) + ((g4575) & (g3015) & (g3009) & (!g2326)));
	assign g6650 = (((!g4574) & (g2326)) + ((g4574) & (!g2326)));
	assign g6651 = (((g830) & (!g6652)));
	assign g6652 = (((g830) & (g6653)));
	assign g6653 = (((!g6654) & (!g6655)));
	assign g6654 = (((!g1914) & (g6656)));
	assign g6655 = (((g1914) & (g6657)));
	assign g6656 = (((!g4556) & (!g3005) & (!g2343) & (g2311)) + ((!g4556) & (!g3005) & (g2343) & (!g2311)) + ((!g4556) & (g3005) & (!g2343) & (!g2311)) + ((!g4556) & (g3005) & (g2343) & (g2311)) + ((g4556) & (!g3005) & (!g2343) & (!g2311)) + ((g4556) & (!g3005) & (g2343) & (g2311)) + ((g4556) & (g3005) & (!g2343) & (g2311)) + ((g4556) & (g3005) & (g2343) & (!g2311)));
	assign g6657 = (((!g4555) & (g2311)) + ((g4555) & (!g2311)));
	assign g6658 = (((!g6659) & (!g6660)));
	assign g6659 = (((!g830) & (g6661)));
	assign g6660 = (((g830) & (g6664)));
	assign g6661 = (((!g6662) & (!g6663)));
	assign g6662 = (((!g1914) & (key[231])));
	assign g6663 = (((g1914) & (key[231])));
	assign g6664 = (((!g6665) & (!g6666)));
	assign g6665 = (((!g1914) & (g6667)));
	assign g6666 = (((g1914) & (g6668)));
	assign g6667 = (((!g1894) & (!g1892) & (g2286)) + ((!g1894) & (g1892) & (!g2286)) + ((g1894) & (!g1892) & (!g2286)) + ((g1894) & (g1892) & (g2286)));
	assign g6668 = (((!g4526) & (g2286)) + ((g4526) & (!g2286)));
	assign g6669 = (((!g6670) & (!g6671)));
	assign g6670 = (((!g830) & (g6672)));
	assign g6671 = (((g830) & (g6675)));
	assign g6672 = (((!g6673) & (!g6674)));
	assign g6673 = (((!g1914) & (nonce[7])));
	assign g6674 = (((g1914) & (nonce[7])));
	assign g6675 = (((!g6676) & (!g6677)));
	assign g6676 = (((!g1914) & (g6678)));
	assign g6677 = (((g1914) & (g6679)));
	assign g6678 = (((!g4513) & (g2279)) + ((g4513) & (!g2279)));
	assign g6679 = (((!g1902) & (!g1886) & (g2279)) + ((!g1902) & (g1886) & (!g2279)) + ((g1902) & (!g1886) & (!g2279)) + ((g1902) & (g1886) & (g2279)));
	assign g6680 = (((!g6681) & (!g6682)));
	assign g6681 = (((!g830) & (g6683)));
	assign g6682 = (((g830) & (g6686)));
	assign g6683 = (((!g6684) & (!g6685)));
	assign g6684 = (((!g1914) & (key[103])));
	assign g6685 = (((g1914) & (key[103])));
	assign g6686 = (((!g6687) & (!g6688)));
	assign g6687 = (((!g1914) & (g6689)));
	assign g6688 = (((g1914) & (g6690)));
	assign g6689 = (((!g828) & (!g1888) & (g2277)) + ((!g828) & (g1888) & (!g2277)) + ((g828) & (!g1888) & (!g2277)) + ((g828) & (g1888) & (g2277)));
	assign g6690 = (((!g4509) & (g2277)) + ((g4509) & (!g2277)));
	assign g6691 = (((!g6692) & (!g6693)));
	assign g6692 = (((!g830) & (g6694)));
	assign g6693 = (((g830) & (g6697)));
	assign g6694 = (((!g6695) & (!g6696)));
	assign g6695 = (((!g1914) & (key[135])));
	assign g6696 = (((g1914) & (key[135])));
	assign g6697 = (((!g6698) & (!g6699)));
	assign g6698 = (((!g1914) & (g6700)));
	assign g6699 = (((g1914) & (g6701)));
	assign g6700 = (((!g4505) & (g2275)) + ((g4505) & (!g2275)));
	assign g6701 = (((!g1900) & (!g1892) & (g2275)) + ((!g1900) & (g1892) & (!g2275)) + ((g1900) & (!g1892) & (!g2275)) + ((g1900) & (g1892) & (g2275)));
	assign g6702 = (((!g6703) & (!g6704)));
	assign g6703 = (((!g830) & (g6705)));
	assign g6704 = (((g830) & (g6708)));
	assign g6705 = (((!g6706) & (!g6707)));
	assign g6706 = (((!g1914) & (g4501)));
	assign g6707 = (((g1914) & (g4501)));
	assign g6708 = (((!g6709) & (!g6710)));
	assign g6709 = (((!g1914) & (g6711)));
	assign g6710 = (((g1914) & (g6712)));
	assign g6711 = (((!g1902) & (!g1898) & (g2273)) + ((!g1902) & (g1898) & (!g2273)) + ((g1902) & (!g1898) & (!g2273)) + ((g1902) & (g1898) & (g2273)));
	assign g6712 = (((!g4500) & (g2273)) + ((g4500) & (!g2273)));
	assign g6713 = (((!g6714) & (!g6715)));
	assign g6714 = (((!g830) & (g6716)));
	assign g6715 = (((g830) & (g6719)));
	assign g6716 = (((!g6717) & (!g6718)));
	assign g6717 = (((!g1914) & (key[7])));
	assign g6718 = (((g1914) & (key[7])));
	assign g6719 = (((!g6720) & (!g6721)));
	assign g6720 = (((!g1914) & (g6722)));
	assign g6721 = (((g1914) & (g6723)));
	assign g6722 = (((!g4490) & (g2267)) + ((g4490) & (!g2267)));
	assign g6723 = (((!g828) & (!g1906) & (g2267)) + ((!g828) & (g1906) & (!g2267)) + ((g828) & (!g1906) & (!g2267)) + ((g828) & (g1906) & (g2267)));
	assign g6724 = (((!g6725) & (!g6726)));
	assign g6725 = (((!g1199) & (g6727)));
	assign g6726 = (((g1199) & (g6730)));
	assign g6727 = (((!g6728) & (!g6729)));
	assign g6728 = (((!g1914) & (g6733)));
	assign g6729 = (((g1914) & (g6734)));
	assign g6730 = (((!g6731) & (!g6732)));
	assign g6731 = (((!g1914) & (g6735)));
	assign g6732 = (((g1914) & (g6736)));
	assign g6733 = (((!g2468) & (g4480)) + ((g2468) & (!g4480)));
	assign g6734 = (((!g2450) & (!g4481) & (g2462)) + ((!g2450) & (g4481) & (!g2462)) + ((g2450) & (!g4481) & (!g2462)) + ((g2450) & (g4481) & (g2462)));
	assign g6735 = (((!g2468) & (!g4480)) + ((g2468) & (g4480)));
	assign g6736 = (((!g2450) & (!g4481) & (g2462)) + ((!g2450) & (g4481) & (!g2462)) + ((g2450) & (!g4481) & (!g2462)) + ((g2450) & (g4481) & (g2462)));
	assign g6737 = (((!g6738) & (!g6739)));
	assign g6738 = (((!g1165) & (g6740)));
	assign g6739 = (((g1165) & (g6743)));
	assign g6740 = (((!g6741) & (!g6742)));
	assign g6741 = (((!g1914) & (g6746)));
	assign g6742 = (((g1914) & (g4425)));
	assign g6743 = (((!g6744) & (!g6745)));
	assign g6744 = (((!g1914) & (g6747)));
	assign g6745 = (((g1914) & (g4425)));
	assign g6746 = (((!g4373) & (!g1132) & (!g2360) & (g2383)) + ((!g4373) & (!g1132) & (g2360) & (g2383)) + ((!g4373) & (g1132) & (!g2360) & (g2383)) + ((!g4373) & (g1132) & (g2360) & (!g2383)) + ((g4373) & (!g1132) & (!g2360) & (g2383)) + ((g4373) & (!g1132) & (g2360) & (!g2383)) + ((g4373) & (g1132) & (!g2360) & (!g2383)) + ((g4373) & (g1132) & (g2360) & (!g2383)));
	assign g6747 = (((!g4373) & (!g1132) & (!g2360) & (!g2383)) + ((!g4373) & (!g1132) & (g2360) & (!g2383)) + ((!g4373) & (g1132) & (!g2360) & (!g2383)) + ((!g4373) & (g1132) & (g2360) & (g2383)) + ((g4373) & (!g1132) & (!g2360) & (!g2383)) + ((g4373) & (!g1132) & (g2360) & (g2383)) + ((g4373) & (g1132) & (!g2360) & (g2383)) + ((g4373) & (g1132) & (g2360) & (g2383)));
	assign g6748 = (((g830) & (!g6749)));
	assign g6749 = (((g830) & (g6750)));
	assign g6750 = (((!g6751) & (!g6752)));
	assign g6751 = (((!g1914) & (g6753)));
	assign g6752 = (((g1914) & (g6754)));
	assign g6753 = (((!g4417) & (g2207)) + ((g4417) & (!g2207)));
	assign g6754 = (((!g4416) & (!g2871) & (!g2868) & (g2207)) + ((!g4416) & (!g2871) & (g2868) & (!g2207)) + ((!g4416) & (g2871) & (!g2868) & (!g2207)) + ((!g4416) & (g2871) & (g2868) & (g2207)) + ((g4416) & (!g2871) & (!g2868) & (!g2207)) + ((g4416) & (!g2871) & (g2868) & (g2207)) + ((g4416) & (g2871) & (!g2868) & (g2207)) + ((g4416) & (g2871) & (g2868) & (!g2207)));
	assign g6755 = (((g830) & (!g6756)));
	assign g6756 = (((g830) & (g6757)));
	assign g6757 = (((!g6758) & (!g6759)));
	assign g6758 = (((!g1914) & (g6760)));
	assign g6759 = (((g1914) & (g6761)));
	assign g6760 = (((!g4402) & (g2198)) + ((g4402) & (!g2198)));
	assign g6761 = (((!g4401) & (!g2863) & (!g2854) & (g2198)) + ((!g4401) & (!g2863) & (g2854) & (!g2198)) + ((!g4401) & (g2863) & (!g2854) & (!g2198)) + ((!g4401) & (g2863) & (g2854) & (g2198)) + ((g4401) & (!g2863) & (!g2854) & (!g2198)) + ((g4401) & (!g2863) & (g2854) & (g2198)) + ((g4401) & (g2863) & (!g2854) & (g2198)) + ((g4401) & (g2863) & (g2854) & (!g2198)));
	assign g6762 = (((g830) & (!g6763)));
	assign g6763 = (((g830) & (g6764)));
	assign g6764 = (((!g6765) & (!g6766)));
	assign g6765 = (((!g1914) & (g6767)));
	assign g6766 = (((g1914) & (g6768)));
	assign g6767 = (((!g4387) & (g2188)) + ((g4387) & (!g2188)));
	assign g6768 = (((!g4386) & (!g2848) & (!g2212) & (g2188)) + ((!g4386) & (!g2848) & (g2212) & (!g2188)) + ((!g4386) & (g2848) & (!g2212) & (!g2188)) + ((!g4386) & (g2848) & (g2212) & (g2188)) + ((g4386) & (!g2848) & (!g2212) & (!g2188)) + ((g4386) & (!g2848) & (g2212) & (g2188)) + ((g4386) & (g2848) & (!g2212) & (g2188)) + ((g4386) & (g2848) & (g2212) & (!g2188)));
	assign g6769 = (((g830) & (!g6770)));
	assign g6770 = (((g830) & (g6771)));
	assign g6771 = (((!g6772) & (!g6773)));
	assign g6772 = (((!g1914) & (g6774)));
	assign g6773 = (((g1914) & (g6775)));
	assign g6774 = (((!g4363) & (g2173)) + ((g4363) & (!g2173)));
	assign g6775 = (((!g4361) & (!g2822) & (!g2810) & (g2173)) + ((!g4361) & (!g2822) & (g2810) & (!g2173)) + ((!g4361) & (g2822) & (!g2810) & (!g2173)) + ((!g4361) & (g2822) & (g2810) & (g2173)) + ((g4361) & (!g2822) & (!g2810) & (!g2173)) + ((g4361) & (!g2822) & (g2810) & (g2173)) + ((g4361) & (g2822) & (!g2810) & (g2173)) + ((g4361) & (g2822) & (g2810) & (!g2173)));
	assign g6776 = (((g830) & (g6777)));
	assign g6777 = (((!g6778) & (!g6779)));
	assign g6778 = (((!g1914) & (g6780)));
	assign g6779 = (((g1914) & (g6781)));
	assign g6780 = (((!g4346) & (g2159)) + ((g4346) & (!g2159)));
	assign g6781 = (((!g4344) & (!g2830) & (!g2797) & (g2159)) + ((!g4344) & (!g2830) & (g2797) & (!g2159)) + ((!g4344) & (g2830) & (!g2797) & (!g2159)) + ((!g4344) & (g2830) & (g2797) & (g2159)) + ((g4344) & (!g2830) & (!g2797) & (!g2159)) + ((g4344) & (!g2830) & (g2797) & (g2159)) + ((g4344) & (g2830) & (!g2797) & (g2159)) + ((g4344) & (g2830) & (g2797) & (!g2159)));
	assign g6782 = (((g830) & (!g6783)));
	assign g6783 = (((g830) & (g6784)));
	assign g6784 = (((!g6785) & (!g6786)));
	assign g6785 = (((!g1914) & (g6787)));
	assign g6786 = (((g1914) & (g6788)));
	assign g6787 = (((!g4326) & (g2144)) + ((g4326) & (!g2144)));
	assign g6788 = (((!g4324) & (!g2816) & (!g2180) & (g2144)) + ((!g4324) & (!g2816) & (g2180) & (!g2144)) + ((!g4324) & (g2816) & (!g2180) & (!g2144)) + ((!g4324) & (g2816) & (g2180) & (g2144)) + ((g4324) & (!g2816) & (!g2180) & (!g2144)) + ((g4324) & (!g2816) & (g2180) & (g2144)) + ((g4324) & (g2816) & (!g2180) & (g2144)) + ((g4324) & (g2816) & (g2180) & (!g2144)));
	assign g6789 = (((!g6790) & (!g6791)));
	assign g6790 = (((!g2396) & (g6792)));
	assign g6791 = (((g2396) & (g6795)));
	assign g6792 = (((!g6793) & (!g6794)));
	assign g6793 = (((!g1914) & (g4318)));
	assign g6794 = (((g1914) & (g6798)));
	assign g6795 = (((!g6796) & (!g6797)));
	assign g6796 = (((!g1914) & (g4318)));
	assign g6797 = (((g1914) & (g6799)));
	assign g6798 = (((!g2369) & (!g4254) & (!g2373) & (g2419)) + ((!g2369) & (!g4254) & (g2373) & (g2419)) + ((!g2369) & (g4254) & (!g2373) & (g2419)) + ((!g2369) & (g4254) & (g2373) & (!g2419)) + ((g2369) & (!g4254) & (!g2373) & (g2419)) + ((g2369) & (!g4254) & (g2373) & (!g2419)) + ((g2369) & (g4254) & (!g2373) & (!g2419)) + ((g2369) & (g4254) & (g2373) & (!g2419)));
	assign g6799 = (((!g2369) & (!g4254) & (!g2373) & (!g2419)) + ((!g2369) & (!g4254) & (g2373) & (!g2419)) + ((!g2369) & (g4254) & (!g2373) & (!g2419)) + ((!g2369) & (g4254) & (g2373) & (g2419)) + ((g2369) & (!g4254) & (!g2373) & (!g2419)) + ((g2369) & (!g4254) & (g2373) & (g2419)) + ((g2369) & (g4254) & (!g2373) & (g2419)) + ((g2369) & (g4254) & (g2373) & (g2419)));
	assign g6800 = (((!g6801) & (!g6802)));
	assign g6801 = (((!g2413) & (g6803)));
	assign g6802 = (((g2413) & (g6806)));
	assign g6803 = (((!g6804) & (!g6805)));
	assign g6804 = (((!g1914) & (g6809)));
	assign g6805 = (((g1914) & (g4311)));
	assign g6806 = (((!g6807) & (!g6808)));
	assign g6807 = (((!g1914) & (g6810)));
	assign g6808 = (((g1914) & (g4311)));
	assign g6809 = (((!g2373) & (!g2358) & (!g4247) & (g2419)) + ((!g2373) & (!g2358) & (g4247) & (g2419)) + ((!g2373) & (g2358) & (!g4247) & (g2419)) + ((!g2373) & (g2358) & (g4247) & (!g2419)) + ((g2373) & (!g2358) & (!g4247) & (g2419)) + ((g2373) & (!g2358) & (g4247) & (!g2419)) + ((g2373) & (g2358) & (!g4247) & (!g2419)) + ((g2373) & (g2358) & (g4247) & (!g2419)));
	assign g6810 = (((!g2373) & (!g2358) & (!g4247) & (!g2419)) + ((!g2373) & (!g2358) & (g4247) & (!g2419)) + ((!g2373) & (g2358) & (!g4247) & (!g2419)) + ((!g2373) & (g2358) & (g4247) & (g2419)) + ((g2373) & (!g2358) & (!g4247) & (!g2419)) + ((g2373) & (!g2358) & (g4247) & (g2419)) + ((g2373) & (g2358) & (!g4247) & (g2419)) + ((g2373) & (g2358) & (g4247) & (g2419)));
	assign g6811 = (((g830) & (g6812)));
	assign g6812 = (((!g6813) & (!g6814)));
	assign g6813 = (((!g1914) & (g6815)));
	assign g6814 = (((g1914) & (g6816)));
	assign g6815 = (((!g4306) & (!g2780) & (!g2772) & (g2127)) + ((!g4306) & (!g2780) & (g2772) & (!g2127)) + ((!g4306) & (g2780) & (!g2772) & (!g2127)) + ((!g4306) & (g2780) & (g2772) & (g2127)) + ((g4306) & (!g2780) & (!g2772) & (!g2127)) + ((g4306) & (!g2780) & (g2772) & (g2127)) + ((g4306) & (g2780) & (!g2772) & (g2127)) + ((g4306) & (g2780) & (g2772) & (!g2127)));
	assign g6816 = (((!g4305) & (g2127)) + ((g4305) & (!g2127)));
	assign g6817 = (((g830) & (!g6818)));
	assign g6818 = (((g830) & (g6819)));
	assign g6819 = (((!g6820) & (!g6821)));
	assign g6820 = (((!g1914) & (g6822)));
	assign g6821 = (((g1914) & (g6823)));
	assign g6822 = (((!g4282) & (!g2785) & (!g2764) & (g2118)) + ((!g4282) & (!g2785) & (g2764) & (!g2118)) + ((!g4282) & (g2785) & (!g2764) & (!g2118)) + ((!g4282) & (g2785) & (g2764) & (g2118)) + ((g4282) & (!g2785) & (!g2764) & (!g2118)) + ((g4282) & (!g2785) & (g2764) & (g2118)) + ((g4282) & (g2785) & (!g2764) & (g2118)) + ((g4282) & (g2785) & (g2764) & (!g2118)));
	assign g6823 = (((!g4281) & (g2118)) + ((g4281) & (!g2118)));
	assign g6824 = (((g830) & (g6825)));
	assign g6825 = (((!g6826) & (!g6827)));
	assign g6826 = (((!g1914) & (g6828)));
	assign g6827 = (((g1914) & (g6829)));
	assign g6828 = (((!g4263) & (!g2776) & (!g2129) & (g2108)) + ((!g4263) & (!g2776) & (g2129) & (!g2108)) + ((!g4263) & (g2776) & (!g2129) & (!g2108)) + ((!g4263) & (g2776) & (g2129) & (g2108)) + ((g4263) & (!g2776) & (!g2129) & (!g2108)) + ((g4263) & (!g2776) & (g2129) & (g2108)) + ((g4263) & (g2776) & (!g2129) & (g2108)) + ((g4263) & (g2776) & (g2129) & (!g2108)));
	assign g6829 = (((!g4262) & (g2108)) + ((g4262) & (!g2108)));
	assign g6830 = (((!g6831) & (!g6832)));
	assign g6831 = (((!g1065) & (g6833)));
	assign g6832 = (((g1065) & (g6836)));
	assign g6833 = (((!g6834) & (!g6835)));
	assign g6834 = (((!g1914) & (g6839)));
	assign g6835 = (((g1914) & (g4251)));
	assign g6836 = (((!g6837) & (!g6838)));
	assign g6837 = (((!g1914) & (g6840)));
	assign g6838 = (((g1914) & (g4251)));
	assign g6839 = (((!g4175) & (!g1031) & (!g2217) & (g2277)) + ((!g4175) & (!g1031) & (g2217) & (g2277)) + ((!g4175) & (g1031) & (!g2217) & (g2277)) + ((!g4175) & (g1031) & (g2217) & (!g2277)) + ((g4175) & (!g1031) & (!g2217) & (g2277)) + ((g4175) & (!g1031) & (g2217) & (!g2277)) + ((g4175) & (g1031) & (!g2217) & (!g2277)) + ((g4175) & (g1031) & (g2217) & (!g2277)));
	assign g6840 = (((!g4175) & (!g1031) & (!g2217) & (!g2277)) + ((!g4175) & (!g1031) & (g2217) & (!g2277)) + ((!g4175) & (g1031) & (!g2217) & (!g2277)) + ((!g4175) & (g1031) & (g2217) & (g2277)) + ((g4175) & (!g1031) & (!g2217) & (!g2277)) + ((g4175) & (!g1031) & (g2217) & (g2277)) + ((g4175) & (g1031) & (!g2217) & (g2277)) + ((g4175) & (g1031) & (g2217) & (g2277)));
	assign g6841 = (((g830) & (!g6842)));
	assign g6842 = (((g830) & (g6843)));
	assign g6843 = (((!g6844) & (!g6845)));
	assign g6844 = (((!g1914) & (g6846)));
	assign g6845 = (((g1914) & (g6847)));
	assign g6846 = (((!g4243) & (g2091)) + ((g4243) & (!g2091)));
	assign g6847 = (((!g4242) & (!g2733) & (!g2713) & (g2091)) + ((!g4242) & (!g2733) & (g2713) & (!g2091)) + ((!g4242) & (g2733) & (!g2713) & (!g2091)) + ((!g4242) & (g2733) & (g2713) & (g2091)) + ((g4242) & (!g2733) & (!g2713) & (!g2091)) + ((g4242) & (!g2733) & (g2713) & (g2091)) + ((g4242) & (g2733) & (!g2713) & (g2091)) + ((g4242) & (g2733) & (g2713) & (!g2091)));
	assign g6848 = (((g830) & (!g6849)));
	assign g6849 = (((g830) & (g6850)));
	assign g6850 = (((!g6851) & (!g6852)));
	assign g6851 = (((!g1914) & (g6853)));
	assign g6852 = (((g1914) & (g6854)));
	assign g6853 = (((!g4226) & (g2077)) + ((g4226) & (!g2077)));
	assign g6854 = (((!g4225) & (!g2747) & (!g2690) & (g2077)) + ((!g4225) & (!g2747) & (g2690) & (!g2077)) + ((!g4225) & (g2747) & (!g2690) & (!g2077)) + ((!g4225) & (g2747) & (g2690) & (g2077)) + ((g4225) & (!g2747) & (!g2690) & (!g2077)) + ((g4225) & (!g2747) & (g2690) & (g2077)) + ((g4225) & (g2747) & (!g2690) & (g2077)) + ((g4225) & (g2747) & (g2690) & (!g2077)));
	assign g6855 = (((g830) & (g6856)));
	assign g6856 = (((!g6857) & (!g6858)));
	assign g6857 = (((!g1914) & (g6859)));
	assign g6858 = (((g1914) & (g6860)));
	assign g6859 = (((!g4193) & (g2062)) + ((g4193) & (!g2062)));
	assign g6860 = (((!g4192) & (!g2723) & (!g2100) & (g2062)) + ((!g4192) & (!g2723) & (g2100) & (!g2062)) + ((!g4192) & (g2723) & (!g2100) & (!g2062)) + ((!g4192) & (g2723) & (g2100) & (g2062)) + ((g4192) & (!g2723) & (!g2100) & (!g2062)) + ((g4192) & (!g2723) & (g2100) & (g2062)) + ((g4192) & (g2723) & (!g2100) & (g2062)) + ((g4192) & (g2723) & (g2100) & (!g2062)));
	assign g6861 = (((!g6862) & (!g6863)));
	assign g6862 = (((!g1031) & (g6864)));
	assign g6863 = (((g1031) & (g6867)));
	assign g6864 = (((!g6865) & (!g6866)));
	assign g6865 = (((!g1914) & (g6870)));
	assign g6866 = (((g1914) & (g6871)));
	assign g6867 = (((!g6868) & (!g6869)));
	assign g6868 = (((!g1914) & (g6872)));
	assign g6869 = (((g1914) & (g6873)));
	assign g6870 = (((!g2217) & (g4175)) + ((g2217) & (!g4175)));
	assign g6871 = (((!g2224) & (!g4176) & (g2247)) + ((!g2224) & (g4176) & (!g2247)) + ((g2224) & (!g4176) & (!g2247)) + ((g2224) & (g4176) & (g2247)));
	assign g6872 = (((!g2217) & (!g4175)) + ((g2217) & (g4175)));
	assign g6873 = (((!g2224) & (!g4176) & (g2247)) + ((!g2224) & (g4176) & (!g2247)) + ((g2224) & (!g4176) & (!g2247)) + ((g2224) & (g4176) & (g2247)));
	assign g6874 = (((g830) & (g6875)));
	assign g6875 = (((!g6876) & (!g6877)));
	assign g6876 = (((!g1914) & (g6878)));
	assign g6877 = (((g1914) & (g6879)));
	assign g6878 = (((!g4166) & (!g2669) & (!g2661) & (g2045)) + ((!g4166) & (!g2669) & (g2661) & (!g2045)) + ((!g4166) & (g2669) & (!g2661) & (!g2045)) + ((!g4166) & (g2669) & (g2661) & (g2045)) + ((g4166) & (!g2669) & (!g2661) & (!g2045)) + ((g4166) & (!g2669) & (g2661) & (g2045)) + ((g4166) & (g2669) & (!g2661) & (g2045)) + ((g4166) & (g2669) & (g2661) & (!g2045)));
	assign g6879 = (((!g4165) & (g2045)) + ((g4165) & (!g2045)));
	assign g6880 = (((g830) & (!g6881)));
	assign g6881 = (((g830) & (g6882)));
	assign g6882 = (((!g6883) & (!g6884)));
	assign g6883 = (((!g1914) & (g6885)));
	assign g6884 = (((g1914) & (g6886)));
	assign g6885 = (((!g4148) & (!g2674) & (!g2653) & (g2036)) + ((!g4148) & (!g2674) & (g2653) & (!g2036)) + ((!g4148) & (g2674) & (!g2653) & (!g2036)) + ((!g4148) & (g2674) & (g2653) & (g2036)) + ((g4148) & (!g2674) & (!g2653) & (!g2036)) + ((g4148) & (!g2674) & (g2653) & (g2036)) + ((g4148) & (g2674) & (!g2653) & (g2036)) + ((g4148) & (g2674) & (g2653) & (!g2036)));
	assign g6886 = (((!g4147) & (g2036)) + ((g4147) & (!g2036)));
	assign g6887 = (((g830) & (!g6888)));
	assign g6888 = (((g830) & (g6889)));
	assign g6889 = (((!g6890) & (!g6891)));
	assign g6890 = (((!g1914) & (g6892)));
	assign g6891 = (((g1914) & (g6893)));
	assign g6892 = (((!g4121) & (!g2665) & (!g2047) & (g2026)) + ((!g4121) & (!g2665) & (g2047) & (!g2026)) + ((!g4121) & (g2665) & (!g2047) & (!g2026)) + ((!g4121) & (g2665) & (g2047) & (g2026)) + ((g4121) & (!g2665) & (!g2047) & (!g2026)) + ((g4121) & (!g2665) & (g2047) & (g2026)) + ((g4121) & (g2665) & (!g2047) & (g2026)) + ((g4121) & (g2665) & (g2047) & (!g2026)));
	assign g6893 = (((!g4120) & (g2026)) + ((g4120) & (!g2026)));
	assign g6894 = (((!g6895) & (!g6896)));
	assign g6895 = (((!g2286) & (g6897)));
	assign g6896 = (((g2286) & (g6900)));
	assign g6897 = (((!g6898) & (!g6899)));
	assign g6898 = (((!g1914) & (g4112)));
	assign g6899 = (((g1914) & (g6903)));
	assign g6900 = (((!g6901) & (!g6902)));
	assign g6901 = (((!g1914) & (g4112)));
	assign g6902 = (((g1914) & (g6904)));
	assign g6903 = (((!g2230) & (!g4106) & (!g2253) & (g2290)) + ((!g2230) & (!g4106) & (g2253) & (g2290)) + ((!g2230) & (g4106) & (!g2253) & (g2290)) + ((!g2230) & (g4106) & (g2253) & (!g2290)) + ((g2230) & (!g4106) & (!g2253) & (g2290)) + ((g2230) & (!g4106) & (g2253) & (!g2290)) + ((g2230) & (g4106) & (!g2253) & (!g2290)) + ((g2230) & (g4106) & (g2253) & (!g2290)));
	assign g6904 = (((!g2230) & (!g4106) & (!g2253) & (!g2290)) + ((!g2230) & (!g4106) & (g2253) & (!g2290)) + ((!g2230) & (g4106) & (!g2253) & (!g2290)) + ((!g2230) & (g4106) & (g2253) & (g2290)) + ((g2230) & (!g4106) & (!g2253) & (!g2290)) + ((g2230) & (!g4106) & (g2253) & (g2290)) + ((g2230) & (g4106) & (!g2253) & (g2290)) + ((g2230) & (g4106) & (g2253) & (g2290)));
	assign g6905 = (((!g6906) & (!g6907)));
	assign g6906 = (((!g998) & (g6908)));
	assign g6907 = (((g998) & (g6911)));
	assign g6908 = (((!g6909) & (!g6910)));
	assign g6909 = (((!g1914) & (g6914)));
	assign g6910 = (((g1914) & (g4109)));
	assign g6911 = (((!g6912) & (!g6913)));
	assign g6912 = (((!g1914) & (g6915)));
	assign g6913 = (((g1914) & (g4109)));
	assign g6914 = (((!g4100) & (!g964) & (!g2137) & (g2194)) + ((!g4100) & (!g964) & (g2137) & (g2194)) + ((!g4100) & (g964) & (!g2137) & (g2194)) + ((!g4100) & (g964) & (g2137) & (!g2194)) + ((g4100) & (!g964) & (!g2137) & (g2194)) + ((g4100) & (!g964) & (g2137) & (!g2194)) + ((g4100) & (g964) & (!g2137) & (!g2194)) + ((g4100) & (g964) & (g2137) & (!g2194)));
	assign g6915 = (((!g4100) & (!g964) & (!g2137) & (!g2194)) + ((!g4100) & (!g964) & (g2137) & (!g2194)) + ((!g4100) & (g964) & (!g2137) & (!g2194)) + ((!g4100) & (g964) & (g2137) & (g2194)) + ((g4100) & (!g964) & (!g2137) & (!g2194)) + ((g4100) & (!g964) & (g2137) & (g2194)) + ((g4100) & (g964) & (!g2137) & (g2194)) + ((g4100) & (g964) & (g2137) & (g2194)));
	assign g6916 = (((!g6917) & (!g6918)));
	assign g6917 = (((!g1914) & (g6919)));
	assign g6918 = (((g1914) & (g6922)));
	assign g6919 = (((!g6920) & (!g6921)));
	assign g6920 = (((!g830) & (key[172])));
	assign g6921 = (((g830) & (g6925)));
	assign g6922 = (((!g6923) & (!g6924)));
	assign g6923 = (((!g830) & (key[172])));
	assign g6924 = (((g830) & (g5697)));
	assign g6925 = (((!g5697) & (!g4094) & (!g3323) & (!g2760)) + ((!g5697) & (!g4094) & (!g3323) & (g2760)) + ((!g5697) & (!g4094) & (g3323) & (!g2760)) + ((!g5697) & (g4094) & (!g3323) & (!g2760)) + ((g5697) & (!g4094) & (g3323) & (g2760)) + ((g5697) & (g4094) & (!g3323) & (g2760)) + ((g5697) & (g4094) & (g3323) & (!g2760)) + ((g5697) & (g4094) & (g3323) & (g2760)));
	assign g6926 = (((!g6927) & (!g6928)));
	assign g6927 = (((!g830) & (g6929)));
	assign g6928 = (((g830) & (g6932)));
	assign g6929 = (((!g6930) & (!g6931)));
	assign g6930 = (((!g1914) & (key[167])));
	assign g6931 = (((g1914) & (key[167])));
	assign g6932 = (((!g6933) & (!g6934)));
	assign g6933 = (((!g1914) & (g6935)));
	assign g6934 = (((g1914) & (g6936)));
	assign g6935 = (((!g4065) & (g1994)) + ((g4065) & (!g1994)));
	assign g6936 = (((!g1912) & (!g1896) & (g1994)) + ((!g1912) & (g1896) & (!g1994)) + ((g1912) & (!g1896) & (!g1994)) + ((g1912) & (g1896) & (g1994)));
	assign g6937 = (((!g6938) & (!g6939)));
	assign g6938 = (((!g1644) & (g6940)));
	assign g6939 = (((g1644) & (g6943)));
	assign g6940 = (((!g6941) & (!g6942)));
	assign g6941 = (((!g1914) & (g6946)));
	assign g6942 = (((g1914) & (g6947)));
	assign g6943 = (((!g6944) & (!g6945)));
	assign g6944 = (((!g1914) & (g6948)));
	assign g6945 = (((g1914) & (g6949)));
	assign g6946 = (((!g3999) & (g3074)) + ((g3999) & (!g3074)));
	assign g6947 = (((!g3093) & (!g3078) & (g3998)) + ((!g3093) & (g3078) & (!g3998)) + ((g3093) & (!g3078) & (!g3998)) + ((g3093) & (g3078) & (g3998)));
	assign g6948 = (((!g3999) & (!g3074)) + ((g3999) & (g3074)));
	assign g6949 = (((!g3093) & (!g3078) & (g3998)) + ((!g3093) & (g3078) & (!g3998)) + ((g3093) & (!g3078) & (!g3998)) + ((g3093) & (g3078) & (g3998)));
	assign g6950 = (((!g6951) & (!g6952)));
	assign g6951 = (((!g2275) & (g6953)));
	assign g6952 = (((g2275) & (g6956)));
	assign g6953 = (((!g6954) & (!g6955)));
	assign g6954 = (((!g1914) & (g6959)));
	assign g6955 = (((g1914) & (g3996)));
	assign g6956 = (((!g6957) & (!g6958)));
	assign g6957 = (((!g1914) & (g6960)));
	assign g6958 = (((g1914) & (g3996)));
	assign g6959 = (((!g2253) & (!g2247) & (!g3990) & (g2290)) + ((!g2253) & (!g2247) & (g3990) & (g2290)) + ((!g2253) & (g2247) & (!g3990) & (g2290)) + ((!g2253) & (g2247) & (g3990) & (!g2290)) + ((g2253) & (!g2247) & (!g3990) & (g2290)) + ((g2253) & (!g2247) & (g3990) & (!g2290)) + ((g2253) & (g2247) & (!g3990) & (!g2290)) + ((g2253) & (g2247) & (g3990) & (!g2290)));
	assign g6960 = (((!g2253) & (!g2247) & (!g3990) & (!g2290)) + ((!g2253) & (!g2247) & (g3990) & (!g2290)) + ((!g2253) & (g2247) & (!g3990) & (!g2290)) + ((!g2253) & (g2247) & (g3990) & (g2290)) + ((g2253) & (!g2247) & (!g3990) & (!g2290)) + ((g2253) & (!g2247) & (g3990) & (g2290)) + ((g2253) & (g2247) & (!g3990) & (g2290)) + ((g2253) & (g2247) & (g3990) & (g2290)));
	assign g6961 = (((!g6962) & (!g6963)));
	assign g6962 = (((!g1914) & (g6964)));
	assign g6963 = (((g1914) & (g6967)));
	assign g6964 = (((!g6965) & (!g6966)));
	assign g6965 = (((!g830) & (key[76])));
	assign g6966 = (((g830) & (g5707)));
	assign g6967 = (((!g6968) & (!g6969)));
	assign g6968 = (((!g830) & (key[76])));
	assign g6969 = (((g830) & (g6970)));
	assign g6970 = (((!g5707) & (!g3979) & (!g3339) & (!g2758)) + ((!g5707) & (!g3979) & (!g3339) & (g2758)) + ((!g5707) & (!g3979) & (g3339) & (!g2758)) + ((!g5707) & (g3979) & (!g3339) & (!g2758)) + ((g5707) & (!g3979) & (g3339) & (g2758)) + ((g5707) & (g3979) & (!g3339) & (g2758)) + ((g5707) & (g3979) & (g3339) & (!g2758)) + ((g5707) & (g3979) & (g3339) & (g2758)));
	assign g6971 = (((!g6972) & (!g6973)));
	assign g6972 = (((!g830) & (g6974)));
	assign g6973 = (((g830) & (g6977)));
	assign g6974 = (((!g6975) & (!g6976)));
	assign g6975 = (((!g1914) & (key[71])));
	assign g6976 = (((g1914) & (key[71])));
	assign g6977 = (((!g6978) & (!g6979)));
	assign g6978 = (((!g1914) & (g6980)));
	assign g6979 = (((g1914) & (g6981)));
	assign g6980 = (((!g1912) & (!g1908) & (g1956)) + ((!g1912) & (g1908) & (!g1956)) + ((g1912) & (!g1908) & (!g1956)) + ((g1912) & (g1908) & (g1956)));
	assign g6981 = (((!g3954) & (g1956)) + ((g3954) & (!g1956)));
	assign g6982 = (((g830) & (g6983)));
	assign g6983 = (((!g6984) & (!g6985)));
	assign g6984 = (((!g1914) & (g6986)));
	assign g6985 = (((g1914) & (g6987)));
	assign g6986 = (((!g3866) & (g1912)) + ((g3866) & (!g1912)));
	assign g6987 = (((!g3855) & (!g2632) & (!g2620) & (g1912)) + ((!g3855) & (!g2632) & (g2620) & (!g1912)) + ((!g3855) & (g2632) & (!g2620) & (!g1912)) + ((!g3855) & (g2632) & (g2620) & (g1912)) + ((g3855) & (!g2632) & (!g2620) & (!g1912)) + ((g3855) & (!g2632) & (g2620) & (g1912)) + ((g3855) & (g2632) & (!g2620) & (g1912)) + ((g3855) & (g2632) & (g2620) & (!g1912)));
	assign g6988 = (((!g6989) & (!g6990)));
	assign g6989 = (((!g3113) & (g6991)));
	assign g6990 = (((g3113) & (g6994)));
	assign g6991 = (((!g6992) & (!g6993)));
	assign g6992 = (((!g1914) & (g3809)));
	assign g6993 = (((g1914) & (g6997)));
	assign g6994 = (((!g6995) & (!g6996)));
	assign g6995 = (((!g1914) & (g3809)));
	assign g6996 = (((g1914) & (g6998)));
	assign g6997 = (((!g3794) & (!g3078) & (!g3086) & (g3116)) + ((!g3794) & (!g3078) & (g3086) & (g3116)) + ((!g3794) & (g3078) & (!g3086) & (g3116)) + ((!g3794) & (g3078) & (g3086) & (!g3116)) + ((g3794) & (!g3078) & (!g3086) & (g3116)) + ((g3794) & (!g3078) & (g3086) & (!g3116)) + ((g3794) & (g3078) & (!g3086) & (!g3116)) + ((g3794) & (g3078) & (g3086) & (!g3116)));
	assign g6998 = (((!g3794) & (!g3078) & (!g3086) & (!g3116)) + ((!g3794) & (!g3078) & (g3086) & (!g3116)) + ((!g3794) & (g3078) & (!g3086) & (!g3116)) + ((!g3794) & (g3078) & (g3086) & (g3116)) + ((g3794) & (!g3078) & (!g3086) & (!g3116)) + ((g3794) & (!g3078) & (g3086) & (g3116)) + ((g3794) & (g3078) & (!g3086) & (g3116)) + ((g3794) & (g3078) & (g3086) & (g3116)));
	assign g6999 = (((!g7000) & (!g7001)));
	assign g7000 = (((!g3142) & (g7002)));
	assign g7001 = (((g3142) & (g7005)));
	assign g7002 = (((!g7003) & (!g7004)));
	assign g7003 = (((!g1914) & (g7008)));
	assign g7004 = (((g1914) & (g7009)));
	assign g7005 = (((!g7006) & (!g7007)));
	assign g7006 = (((!g1914) & (g7010)));
	assign g7007 = (((g1914) & (g7011)));
	assign g7008 = (((!g3119) & (g3776)) + ((g3119) & (!g3776)));
	assign g7009 = (((!g2838) & (!g2210) & (g3758)) + ((!g2838) & (g2210) & (!g3758)) + ((g2838) & (!g2210) & (!g3758)) + ((g2838) & (g2210) & (g3758)));
	assign g7010 = (((!g3119) & (!g3776)) + ((g3119) & (g3776)));
	assign g7011 = (((!g2838) & (!g2210) & (g3758)) + ((!g2838) & (g2210) & (!g3758)) + ((g2838) & (!g2210) & (!g3758)) + ((g2838) & (g2210) & (g3758)));
	assign g7012 = (((g830) & (g7013)));
	assign g7013 = (((!g7014) & (!g7015)));
	assign g7014 = (((!g1914) & (g7016)));
	assign g7015 = (((g1914) & (g7017)));
	assign g7016 = (((!g3709) & (g1902)) + ((g3709) & (!g1902)));
	assign g7017 = (((!g3698) & (!g2640) & (!g2607) & (g1902)) + ((!g3698) & (!g2640) & (g2607) & (!g1902)) + ((!g3698) & (g2640) & (!g2607) & (!g1902)) + ((!g3698) & (g2640) & (g2607) & (g1902)) + ((g3698) & (!g2640) & (!g2607) & (!g1902)) + ((g3698) & (!g2640) & (g2607) & (g1902)) + ((g3698) & (g2640) & (!g2607) & (g1902)) + ((g3698) & (g2640) & (g2607) & (!g1902)));
	assign g7018 = (((!g7019) & (!g7020)));
	assign g7019 = (((!g2516) & (g7021)));
	assign g7020 = (((g2516) & (g7024)));
	assign g7021 = (((!g7022) & (!g7023)));
	assign g7022 = (((!g1914) & (g3652)));
	assign g7023 = (((g1914) & (g7027)));
	assign g7024 = (((!g7025) & (!g7026)));
	assign g7025 = (((!g1914) & (g3652)));
	assign g7026 = (((g1914) & (g7028)));
	assign g7027 = (((!g1644) & (!g2424) & (!g3637) & (g1677)) + ((!g1644) & (!g2424) & (g3637) & (g1677)) + ((!g1644) & (g2424) & (!g3637) & (g1677)) + ((!g1644) & (g2424) & (g3637) & (!g1677)) + ((g1644) & (!g2424) & (!g3637) & (g1677)) + ((g1644) & (!g2424) & (g3637) & (!g1677)) + ((g1644) & (g2424) & (!g3637) & (!g1677)) + ((g1644) & (g2424) & (g3637) & (!g1677)));
	assign g7028 = (((!g1644) & (!g2424) & (!g3637) & (!g1677)) + ((!g1644) & (!g2424) & (g3637) & (!g1677)) + ((!g1644) & (g2424) & (!g3637) & (!g1677)) + ((!g1644) & (g2424) & (g3637) & (g1677)) + ((g1644) & (!g2424) & (!g3637) & (!g1677)) + ((g1644) & (!g2424) & (g3637) & (g1677)) + ((g1644) & (g2424) & (!g3637) & (g1677)) + ((g1644) & (g2424) & (g3637) & (g1677)));
	assign g7029 = (((!g7030) & (!g7031)));
	assign g7030 = (((!g3619) & (g7032)));
	assign g7031 = (((g3619) & (g7035)));
	assign g7032 = (((!g7033) & (!g7034)));
	assign g7033 = (((!g1914) & (g7038)));
	assign g7034 = (((g1914) & (g7039)));
	assign g7035 = (((!g7036) & (!g7037)));
	assign g7036 = (((!g1914) & (g7040)));
	assign g7037 = (((g1914) & (g7041)));
	assign g7038 = (((!g3125) & (g3113)) + ((g3125) & (!g3113)));
	assign g7039 = (((!g3601) & (!g2213) & (g2871)) + ((!g3601) & (g2213) & (!g2871)) + ((g3601) & (!g2213) & (!g2871)) + ((g3601) & (g2213) & (g2871)));
	assign g7040 = (((!g3125) & (!g3113)) + ((g3125) & (g3113)));
	assign g7041 = (((!g3601) & (!g2213) & (g2871)) + ((!g3601) & (g2213) & (!g2871)) + ((g3601) & (!g2213) & (!g2871)) + ((g3601) & (g2213) & (g2871)));
	assign g7042 = (((!g7043) & (!g7044)));
	assign g7043 = (((!g3122) & (g7045)));
	assign g7044 = (((g3122) & (g7048)));
	assign g7045 = (((!g7046) & (!g7047)));
	assign g7046 = (((!g1914) & (g3586)));
	assign g7047 = (((g1914) & (g7051)));
	assign g7048 = (((!g7049) & (!g7050)));
	assign g7049 = (((!g1914) & (g3586)));
	assign g7050 = (((g1914) & (g7052)));
	assign g7051 = (((!g3074) & (!g3571) & (!g3088) & (g3128)) + ((!g3074) & (!g3571) & (g3088) & (g3128)) + ((!g3074) & (g3571) & (!g3088) & (g3128)) + ((!g3074) & (g3571) & (g3088) & (!g3128)) + ((g3074) & (!g3571) & (!g3088) & (g3128)) + ((g3074) & (!g3571) & (g3088) & (!g3128)) + ((g3074) & (g3571) & (!g3088) & (!g3128)) + ((g3074) & (g3571) & (g3088) & (!g3128)));
	assign g7052 = (((!g3074) & (!g3571) & (!g3088) & (!g3128)) + ((!g3074) & (!g3571) & (g3088) & (!g3128)) + ((!g3074) & (g3571) & (!g3088) & (!g3128)) + ((!g3074) & (g3571) & (g3088) & (g3128)) + ((g3074) & (!g3571) & (!g3088) & (!g3128)) + ((g3074) & (!g3571) & (g3088) & (g3128)) + ((g3074) & (g3571) & (!g3088) & (g3128)) + ((g3074) & (g3571) & (g3088) & (g3128)));
	assign g7053 = (((g830) & (g7054)));
	assign g7054 = (((!g7055) & (!g7056)));
	assign g7055 = (((!g1914) & (g7057)));
	assign g7056 = (((g1914) & (g7058)));
	assign g7057 = (((!g3554) & (g1892)) + ((g3554) & (!g1892)));
	assign g7058 = (((!g2626) & (!g3543) & (!g2013) & (g1892)) + ((!g2626) & (!g3543) & (g2013) & (!g1892)) + ((!g2626) & (g3543) & (!g2013) & (!g1892)) + ((!g2626) & (g3543) & (g2013) & (g1892)) + ((g2626) & (!g3543) & (!g2013) & (!g1892)) + ((g2626) & (!g3543) & (g2013) & (g1892)) + ((g2626) & (g3543) & (!g2013) & (g1892)) + ((g2626) & (g3543) & (g2013) & (!g1892)));
	assign g7059 = (((!g7060) & (!g7061)));
	assign g7060 = (((!g3136) & (g7062)));
	assign g7061 = (((g3136) & (g7065)));
	assign g7062 = (((!g7063) & (!g7064)));
	assign g7063 = (((!g1914) & (g3497)));
	assign g7064 = (((g1914) & (g7068)));
	assign g7065 = (((!g7066) & (!g7067)));
	assign g7066 = (((!g1914) & (g3497)));
	assign g7067 = (((g1914) & (g7069)));
	assign g7068 = (((!g3082) & (!g3482) & (!g3097) & (g3142)) + ((!g3082) & (!g3482) & (g3097) & (g3142)) + ((!g3082) & (g3482) & (!g3097) & (g3142)) + ((!g3082) & (g3482) & (g3097) & (!g3142)) + ((g3082) & (!g3482) & (!g3097) & (g3142)) + ((g3082) & (!g3482) & (g3097) & (!g3142)) + ((g3082) & (g3482) & (!g3097) & (!g3142)) + ((g3082) & (g3482) & (g3097) & (!g3142)));
	assign g7069 = (((!g3082) & (!g3482) & (!g3097) & (!g3142)) + ((!g3082) & (!g3482) & (g3097) & (!g3142)) + ((!g3082) & (g3482) & (!g3097) & (!g3142)) + ((!g3082) & (g3482) & (g3097) & (g3142)) + ((g3082) & (!g3482) & (!g3097) & (!g3142)) + ((g3082) & (!g3482) & (g3097) & (g3142)) + ((g3082) & (g3482) & (!g3097) & (g3142)) + ((g3082) & (g3482) & (g3097) & (g3142)));
	assign g7070 = (((!g7071) & (!g7072)));
	assign g7071 = (((!g2519) & (g7073)));
	assign g7072 = (((g2519) & (g7076)));
	assign g7073 = (((!g7074) & (!g7075)));
	assign g7074 = (((!g1914) & (g7079)));
	assign g7075 = (((g1914) & (g7080)));
	assign g7076 = (((!g7077) & (!g7078)));
	assign g7077 = (((!g1914) & (g7081)));
	assign g7078 = (((g1914) & (g7082)));
	assign g7079 = (((!g3461) & (g1677)) + ((g3461) & (!g1677)));
	assign g7080 = (((!g2857) & (!g3443) & (g2863)) + ((!g2857) & (g3443) & (!g2863)) + ((g2857) & (!g3443) & (!g2863)) + ((g2857) & (g3443) & (g2863)));
	assign g7081 = (((!g3461) & (!g1677)) + ((g3461) & (g1677)));
	assign g7082 = (((!g2857) & (!g3443) & (g2863)) + ((!g2857) & (g3443) & (!g2863)) + ((g2857) & (!g3443) & (!g2863)) + ((g2857) & (g3443) & (g2863)));
	assign g7083 = (((g830) & (g7084)));
	assign g7084 = (((!g7085) & (!g7086)));
	assign g7085 = (((!g1914) & (g7087)));
	assign g7086 = (((g1914) & (g7088)));
	assign g7087 = (((!g3391) & (g1881)) + ((g3391) & (!g1881)));
	assign g7088 = (((!g1973) & (!g1972) & (!g1971) & (g1881)) + ((!g1973) & (!g1972) & (g1971) & (!g1881)) + ((!g1973) & (g1972) & (!g1971) & (!g1881)) + ((!g1973) & (g1972) & (g1971) & (g1881)) + ((g1973) & (!g1972) & (!g1971) & (!g1881)) + ((g1973) & (!g1972) & (g1971) & (g1881)) + ((g1973) & (g1972) & (!g1971) & (g1881)) + ((g1973) & (g1972) & (g1971) & (!g1881)));
	assign g7089 = (((g830) & (g7090)));
	assign g7090 = (((!g7091) & (!g7092)));
	assign g7091 = (((!g1914) & (g7093)));
	assign g7092 = (((g1914) & (g7094)));
	assign g7093 = (((!g2002) & (!g2001) & (!g2000) & (g1778)) + ((!g2002) & (!g2001) & (g2000) & (!g1778)) + ((!g2002) & (g2001) & (!g2000) & (!g1778)) + ((!g2002) & (g2001) & (g2000) & (g1778)) + ((g2002) & (!g2001) & (!g2000) & (!g1778)) + ((g2002) & (!g2001) & (g2000) & (g1778)) + ((g2002) & (g2001) & (!g2000) & (g1778)) + ((g2002) & (g2001) & (g2000) & (!g1778)));
	assign g7094 = (((!g3289) & (g1778)) + ((g3289) & (!g1778)));
	assign g7095 = (((g830) & (g7096)));
	assign g7096 = (((!g7097) & (!g7098)));
	assign g7097 = (((!g1914) & (g7099)));
	assign g7098 = (((g1914) & (g7100)));
	assign g7099 = (((!g3217) & (g1744)) + ((g3217) & (!g1744)));
	assign g7100 = (((!g1961) & (!g1960) & (!g3216) & (g1744)) + ((!g1961) & (!g1960) & (g3216) & (!g1744)) + ((!g1961) & (g1960) & (!g3216) & (!g1744)) + ((!g1961) & (g1960) & (g3216) & (g1744)) + ((g1961) & (!g1960) & (!g3216) & (!g1744)) + ((g1961) & (!g1960) & (g3216) & (g1744)) + ((g1961) & (g1960) & (!g3216) & (g1744)) + ((g1961) & (g1960) & (g3216) & (!g1744)));
	assign g7101 = (((g830) & (g7102)));
	assign g7102 = (((!g7103) & (!g7104)));
	assign g7103 = (((!g1914) & (g7105)));
	assign g7104 = (((g1914) & (g7106)));
	assign g7105 = (((!g3174) & (g1711)) + ((g3174) & (!g1711)));
	assign g7106 = (((!g1959) & (!g1958) & (!g1957) & (g1711)) + ((!g1959) & (!g1958) & (g1957) & (!g1711)) + ((!g1959) & (g1958) & (!g1957) & (!g1711)) + ((!g1959) & (g1958) & (g1957) & (g1711)) + ((g1959) & (!g1958) & (!g1957) & (!g1711)) + ((g1959) & (!g1958) & (g1957) & (g1711)) + ((g1959) & (g1958) & (!g1957) & (g1711)) + ((g1959) & (g1958) & (g1957) & (!g1711)));
	assign g7107 = (((g830) & (!g7108)));
	assign g7108 = (((g830) & (g7109)));
	assign g7109 = (((!g7110) & (!g7111)));
	assign g7110 = (((!g1914) & (g7112)));
	assign g7111 = (((g1914) & (g7113)));
	assign g7112 = (((!g2997) & (g1540)) + ((g2997) & (!g1540)));
	assign g7113 = (((!g1945) & (!g1944) & (!g1943) & (g1540)) + ((!g1945) & (!g1944) & (g1943) & (!g1540)) + ((!g1945) & (g1944) & (!g1943) & (!g1540)) + ((!g1945) & (g1944) & (g1943) & (g1540)) + ((g1945) & (!g1944) & (!g1943) & (!g1540)) + ((g1945) & (!g1944) & (g1943) & (g1540)) + ((g1945) & (g1944) & (!g1943) & (g1540)) + ((g1945) & (g1944) & (g1943) & (!g1540)));
	assign g7114 = (((g830) & (g7115)));
	assign g7115 = (((!g7116) & (!g7117)));
	assign g7116 = (((!g1914) & (g7118)));
	assign g7117 = (((g1914) & (g7119)));
	assign g7118 = (((!g1888) & (!g1884) & (g1439)) + ((!g1888) & (g1884) & (!g1439)) + ((g1888) & (!g1884) & (!g1439)) + ((g1888) & (g1884) & (g1439)));
	assign g7119 = (((!g1906) & (!g1890) & (g1439)) + ((!g1906) & (g1890) & (!g1439)) + ((g1906) & (!g1890) & (!g1439)) + ((g1906) & (g1890) & (g1439)));
	assign g7120 = (((g830) & (g7121)));
	assign g7121 = (((!g7122) & (!g7123)));
	assign g7122 = (((!g1914) & (g7124)));
	assign g7123 = (((g1914) & (g7125)));
	assign g7124 = (((!g2794) & (!g2793) & (!g2792) & (g1406)) + ((!g2794) & (!g2793) & (g2792) & (!g1406)) + ((!g2794) & (g2793) & (!g2792) & (!g1406)) + ((!g2794) & (g2793) & (g2792) & (g1406)) + ((g2794) & (!g2793) & (!g2792) & (!g1406)) + ((g2794) & (!g2793) & (g2792) & (g1406)) + ((g2794) & (g2793) & (!g2792) & (g1406)) + ((g2794) & (g2793) & (g2792) & (!g1406)));
	assign g7125 = (((!g2791) & (g1406)) + ((g2791) & (!g1406)));
	assign g7126 = (((g830) & (!g7127)));
	assign g7127 = (((g830) & (g7128)));
	assign g7128 = (((!g7129) & (!g7130)));
	assign g7129 = (((!g1914) & (g7131)));
	assign g7130 = (((g1914) & (g7132)));
	assign g7131 = (((!g2651) & (g1303)) + ((g2651) & (!g1303)));
	assign g7132 = (((!g2648) & (!g2647) & (!g2646) & (g1303)) + ((!g2648) & (!g2647) & (g2646) & (!g1303)) + ((!g2648) & (g2647) & (!g2646) & (!g1303)) + ((!g2648) & (g2647) & (g2646) & (g1303)) + ((g2648) & (!g2647) & (!g2646) & (!g1303)) + ((g2648) & (!g2647) & (g2646) & (g1303)) + ((g2648) & (g2647) & (!g2646) & (g1303)) + ((g2648) & (g2647) & (g2646) & (!g1303)));
	assign g7133 = (((g830) & (!g7134)));
	assign g7134 = (((g830) & (g7135)));
	assign g7135 = (((!g7136) & (!g7137)));
	assign g7136 = (((!g1914) & (g7138)));
	assign g7137 = (((g1914) & (g7139)));
	assign g7138 = (((!g2556) & (!g2555) & (!g2554) & (g1236)) + ((!g2556) & (!g2555) & (g2554) & (!g1236)) + ((!g2556) & (g2555) & (!g2554) & (!g1236)) + ((!g2556) & (g2555) & (g2554) & (g1236)) + ((g2556) & (!g2555) & (!g2554) & (!g1236)) + ((g2556) & (!g2555) & (g2554) & (g1236)) + ((g2556) & (g2555) & (!g2554) & (g1236)) + ((g2556) & (g2555) & (g2554) & (!g1236)));
	assign g7139 = (((!g2553) & (g1236)) + ((g2553) & (!g1236)));
	assign g7140 = (((g830) & (g7141)));
	assign g7141 = (((!g7142) & (!g7143)));
	assign g7142 = (((!g1914) & (g7144)));
	assign g7143 = (((g1914) & (g7145)));
	assign g7144 = (((!g2428) & (g1165)) + ((g2428) & (!g1165)));
	assign g7145 = (((!g2424) & (!g2423) & (!g2422) & (g1165)) + ((!g2424) & (!g2423) & (g2422) & (!g1165)) + ((!g2424) & (g2423) & (!g2422) & (!g1165)) + ((!g2424) & (g2423) & (g2422) & (g1165)) + ((g2424) & (!g2423) & (!g2422) & (!g1165)) + ((g2424) & (!g2423) & (g2422) & (g1165)) + ((g2424) & (g2423) & (!g2422) & (g1165)) + ((g2424) & (g2423) & (g2422) & (!g1165)));
	assign g7146 = (((g830) & (g7147)));
	assign g7147 = (((!g7148) & (!g7149)));
	assign g7148 = (((!g1914) & (g7150)));
	assign g7149 = (((g1914) & (g7151)));
	assign g7150 = (((!g2380) & (g1132)) + ((g2380) & (!g1132)));
	assign g7151 = (((!g2377) & (!g2376) & (!g2375) & (g1132)) + ((!g2377) & (!g2376) & (g2375) & (!g1132)) + ((!g2377) & (g2376) & (!g2375) & (!g1132)) + ((!g2377) & (g2376) & (g2375) & (g1132)) + ((g2377) & (!g2376) & (!g2375) & (!g1132)) + ((g2377) & (!g2376) & (g2375) & (g1132)) + ((g2377) & (g2376) & (!g2375) & (g1132)) + ((g2377) & (g2376) & (g2375) & (!g1132)));
	assign g7152 = (((g830) & (g7153)));
	assign g7153 = (((!g7154) & (!g7155)));
	assign g7154 = (((!g1914) & (g7156)));
	assign g7155 = (((g1914) & (g7157)));
	assign g7156 = (((!g2348) & (!g2347) & (!g2346) & (g1098)) + ((!g2348) & (!g2347) & (g2346) & (!g1098)) + ((!g2348) & (g2347) & (!g2346) & (!g1098)) + ((!g2348) & (g2347) & (g2346) & (g1098)) + ((g2348) & (!g2347) & (!g2346) & (!g1098)) + ((g2348) & (!g2347) & (g2346) & (g1098)) + ((g2348) & (g2347) & (!g2346) & (g1098)) + ((g2348) & (g2347) & (g2346) & (!g1098)));
	assign g7157 = (((!g2345) & (g1098)) + ((g2345) & (!g1098)));
	assign g7158 = (((g830) & (!g7159)));
	assign g7159 = (((g830) & (g7160)));
	assign g7160 = (((!g7161) & (!g7162)));
	assign g7161 = (((!g1914) & (g7163)));
	assign g7162 = (((g1914) & (g7164)));
	assign g7163 = (((!g2214) & (g998)) + ((g2214) & (!g998)));
	assign g7164 = (((!g2211) & (!g2210) & (!g2209) & (g998)) + ((!g2211) & (!g2210) & (g2209) & (!g998)) + ((!g2211) & (g2210) & (!g2209) & (!g998)) + ((!g2211) & (g2210) & (g2209) & (g998)) + ((g2211) & (!g2210) & (!g2209) & (!g998)) + ((g2211) & (!g2210) & (g2209) & (g998)) + ((g2211) & (g2210) & (!g2209) & (g998)) + ((g2211) & (g2210) & (g2209) & (!g998)));
	assign g7165 = (((g830) & (g7166)));
	assign g7166 = (((!g7167) & (!g7168)));
	assign g7167 = (((!g1914) & (g7169)));
	assign g7168 = (((g1914) & (g7170)));
	assign g7169 = (((!g2182) & (g964)) + ((g2182) & (!g964)));
	assign g7170 = (((!g2178) & (!g2177) & (!g2176) & (g964)) + ((!g2178) & (!g2177) & (g2176) & (!g964)) + ((!g2178) & (g2177) & (!g2176) & (!g964)) + ((!g2178) & (g2177) & (g2176) & (g964)) + ((g2178) & (!g2177) & (!g2176) & (!g964)) + ((g2178) & (!g2177) & (g2176) & (g964)) + ((g2178) & (g2177) & (!g2176) & (g964)) + ((g2178) & (g2177) & (g2176) & (!g964)));
	assign g7171 = (((g830) & (g7172)));
	assign g7172 = (((!g7173) & (!g7174)));
	assign g7173 = (((!g1914) & (g7175)));
	assign g7174 = (((g1914) & (g7176)));
	assign g7175 = (((!g2134) & (!g2133) & (!g2132) & (g931)) + ((!g2134) & (!g2133) & (g2132) & (!g931)) + ((!g2134) & (g2133) & (!g2132) & (!g931)) + ((!g2134) & (g2133) & (g2132) & (g931)) + ((g2134) & (!g2133) & (!g2132) & (!g931)) + ((g2134) & (!g2133) & (g2132) & (g931)) + ((g2134) & (g2133) & (!g2132) & (g931)) + ((g2134) & (g2133) & (g2132) & (!g931)));
	assign g7176 = (((!g2131) & (g931)) + ((g2131) & (!g931)));
	assign g7177 = (((g830) & (!g7178)));
	assign g7178 = (((g830) & (g7179)));
	assign g7179 = (((!g7180) & (!g7181)));
	assign g7180 = (((!g1914) & (g7182)));
	assign g7181 = (((g1914) & (g7183)));
	assign g7182 = (((!g2102) & (g897)) + ((g2102) & (!g897)));
	assign g7183 = (((!g2099) & (!g2098) & (!g2097) & (g897)) + ((!g2099) & (!g2098) & (g2097) & (!g897)) + ((!g2099) & (g2098) & (!g2097) & (!g897)) + ((!g2099) & (g2098) & (g2097) & (g897)) + ((g2099) & (!g2098) & (!g2097) & (!g897)) + ((g2099) & (!g2098) & (g2097) & (g897)) + ((g2099) & (g2098) & (!g2097) & (g897)) + ((g2099) & (g2098) & (g2097) & (!g897)));
	assign g7184 = (((g830) & (g7185)));
	assign g7185 = (((!g7186) & (!g7187)));
	assign g7186 = (((!g1914) & (g7188)));
	assign g7187 = (((g1914) & (g7189)));
	assign g7188 = (((!g2052) & (!g2051) & (!g2050) & (g864)) + ((!g2052) & (!g2051) & (g2050) & (!g864)) + ((!g2052) & (g2051) & (!g2050) & (!g864)) + ((!g2052) & (g2051) & (g2050) & (g864)) + ((g2052) & (!g2051) & (!g2050) & (!g864)) + ((g2052) & (!g2051) & (g2050) & (g864)) + ((g2052) & (g2051) & (!g2050) & (g864)) + ((g2052) & (g2051) & (g2050) & (!g864)));
	assign g7189 = (((!g2049) & (g864)) + ((g2049) & (!g864)));
	assign g7190 = (((g830) & (!g7191)));
	assign g7191 = (((g830) & (g7192)));
	assign g7192 = (((!g7193) & (!g7194)));
	assign g7193 = (((!g1914) & (g7195)));
	assign g7194 = (((g1914) & (g7196)));
	assign g7195 = (((!g2015) & (g828)) + ((g2015) & (!g828)));
	assign g7196 = (((!g1976) & (!g1975) & (!g1974) & (g828)) + ((!g1976) & (!g1975) & (g1974) & (!g828)) + ((!g1976) & (g1975) & (!g1974) & (!g828)) + ((!g1976) & (g1975) & (g1974) & (g828)) + ((g1976) & (!g1975) & (!g1974) & (!g828)) + ((g1976) & (!g1975) & (g1974) & (g828)) + ((g1976) & (g1975) & (!g1974) & (g828)) + ((g1976) & (g1975) & (g1974) & (!g828)));

endmodule