module misex3 (
	a, b, c, d, e, f, g, h, 
	i, j, k, l, m, n, r2, s2, t2, u2, 
	n2, o2, p2, q2, h2, i2, j2, k2, m2, l2);

input a, b, c, d, e, f, g, h, i, j, k, l, m, n;

output r2, s2, t2, u2, n2, o2, p2, q2, h2, i2, j2, k2, m2, l2;

wire n1, n917, n3, n4, n8, n10, n11, n12, n9, n14, n15, n16, n17, n13, n18, n23, n24, n25, n26, n27, n19, n29, n32, n33, n34, n35, n28, n40, n41, n42, n43, n44, n36, n46, n45, n49, n47, n52, n53, n54, n51, n58, n57, n55, n61, n62, n60, n59, n66, n64, n65, n63, n68, n69, n70, n67, n73, n72, n71, n75, n76, n77, n74, n79, n80, n78, n82, n81, n84, n83, n88, n86, n87, n85, n91, n90, n89, n93, n94, n92, n96, n95, n100, n101, n98, n99, n97, n103, n102, n106, n107, n105, n104, n109, n110, n108, n111, n115, n119, n123, n130, n131, n132, n133, n134, n135, n128, n138, n139, n137, n136, n142, n141, n140, n144, n145, n143, n149, n150, n147, n148, n146, n152, n151, n156, n154, n155, n153, n159, n160, n157, n163, n162, n161, n165, n164, n167, n168, n169, n170, n166, n172, n173, n171, n174, n182, n181, n180, n179, n186, n184, n185, n183, n187, n189, n190, n188, n192, n193, n191, n195, n194, n196, n200, n198, n199, n197, n201, n206, n207, n208, n209, n210, n211, n212, n205, n214, n215, n213, n219, n218, n216, n222, n223, n221, n227, n228, n226, n225, n230, n229, n231, n238, n236, n235, n241, n239, n242, n247, n246, n250, n249, n248, n251, n253, n254, n252, n256, n255, n258, n259, n260, n261, n257, n262, n265, n266, n264, n263, n268, n267, n269, n274, n275, n278, n281, n288, n287, n286, n290, n289, n293, n292, n295, n296, n294, n299, n300, n298, n297, n301, n303, n302, n307, n305, n306, n304, n309, n310, n311, n312, n308, n313, n315, n314, n316, n320, n323, n324, n322, n327, n325, n330, n329, n328, n331, n332, n338, n339, n337, n336, n341, n342, n343, n340, n345, n346, n344, n349, n350, n348, n347, n352, n351, n355, n354, n353, n357, n356, n360, n359, n358, n363, n362, n361, n364, n369, n372, n371, n373, n379, n380, n381, n382, n383, n384, n385, n378, n388, n387, n390, n391, n389, n395, n393, n394, n392, n399, n398, n397, n400, n401, n402, n406, n405, n410, n409, n408, n407, n412, n413, n411, n417, n416, n415, n414, n419, n418, n421, n422, n423, n424, n425, n426, n427, n428, n420, n429, n434, n435, n433, n437, n436, n439, n440, n441, n438, n443, n442, n446, n445, n449, n447, n452, n453, n451, n450, n454, n455, n457, n461, n459, n462, n465, n468, n472, n476, n479, n482, n485, n484, n488, n489, n487, n491, n492, n490, n494, n495, n493, n497, n498, n496, n500, n501, n499, n504, n503, n505, n506, n507, n508, n512, n510, n511, n509, n514, n513, n516, n517, n515, n519, n520, n521, n518, n522, n523, n526, n527, n525, n532, n530, n529, n534, n533, n535, n536, n542, n543, n541, n539, n545, n544, n546, n548, n552, n551, n554, n553, n556, n558, n559, n560, n561, n555, n562, n564, n563, n566, n565, n568, n572, n573, n571, n574, n576, n575, n578, n579, n580, n581, n577, n582, n585, n587, n588, n589, n590, n592, n586, n596, n597, n595, n593, n598, n600, n599, n603, n601, n605, n604, n606, n609, n608, n610, n612, n611, n615, n616, n617, n618, n614, n621, n619, n624, n627, n628, n629, n633, n634, n637, n640, n641, n644, n642, n645, n648, n651, n652, n653, n654, n655, n657, n656, n660, n659, n658, n661, n665, n663, n667, n668, n669, n670, n671, n672, n673, n666, n675, n674, n676, n677, n678, n679, n680, n681, n682, n683, n685, n686, n687, n688, n689, n690, n684, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n721, n722, n723, n724, n725, n726, n727, n728, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n758, n759, n760, n761, n762, n763, n764, n765, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n782, n783, n784, n785, n786, n788, n789, n790, n792, n794, n796, n799, n798, n797, n801, n800, n802, n803, n806, n808, n809, n810, n811, n813, n815, n816, n817, n818, n819, n820, n821, n823, n824, n827, n831, n833, n834, n836, n837, n838, n839, n840, n842, n843, n844, n845, n847, n848, n849, n850, n852, n851, n854, n856, n857, n860, n861, n859, n862, n864, n865, n867, n871, n872, n870, n869, n874, n875, n876, n878, n880, n882, n883, n886, n888, n892, n893, n894, n895, n896, n897, n899, n898, n900, n902, n903, n904, n905, n906, n908, n911, n912, n914;

assign r2 = ( (~ n308) ) ;
 assign s2 = ( (~ n36) ) ;
 assign t2 = ( (~ n205) ) ;
 assign u2 = ( (~ n128) ) ;
 assign n2 = ( (~ n28) ) ;
 assign o2 = ( (~ n19) ) ;
 assign p2 = ( (~ n420) ) ;
 assign q2 = ( (~ n378) ) ;
 assign h2 = ( (~ n18) ) ;
 assign i2 = ( (~ n666) ) ;
 assign j2 = ( (~ n13) ) ;
 assign k2 = ( (~ n9) ) ;
 assign m2 = ( (~ n518) ) ;
 assign l2 = ( n1 ) | ( n917 ) | ( n3 ) | ( n4 ) | ( n8 ) | ( (~ n894) ) | ( (~ n905) ) | ( (~ n908) ) ;
 assign n1 = ( f  &  (~ n796) ) | ( f  &  (~ n878) ) | ( f  &  (~ n880) ) ;
 assign n917 = ( (~ f)  &  n546 ) | ( (~ f)  &  n548 ) | ( (~ f)  &  (~ n869) ) ;
 assign n3 = ( (~ n)  &  (~ n854) ) | ( (~ n)  &  (~ n857) ) | ( (~ n)  &  (~ n862) ) ;
 assign n4 = ( n  &  (~ n599) ) | ( n  &  (~ n865) ) | ( n  &  (~ n867) ) ;
 assign n8 = ( (~ n633) ) | ( n634 ) | ( n637 ) | ( (~ n640) ) | ( n641 ) | ( n645 ) | ( n648 ) | ( (~ n888) ) ;
 assign n10 = ( i ) | ( l ) | ( n413 ) | ( n788 ) | ( n789 ) ;
 assign n11 = ( n651 ) | ( n180 ) | ( n504 ) ;
 assign n12 = ( n499  &  n503  &  n14  &  n772  &  n773  &  n496 ) ;
 assign n9 = ( n10  &  n11  &  n12 ) ;
 assign n14 = ( n487  &  n490  &  n493  &  n767  &  n677  &  n768 ) ;
 assign n15 = ( n505  &  n506  &  n507  &  n508 ) ;
 assign n16 = ( n180 ) | ( n504 ) | ( n788 ) ;
 assign n17 = ( n652 ) | ( n653 ) | ( n168 ) | ( n553 ) ;
 assign n13 = ( n14  &  n15  &  n16  &  n17 ) ;
 assign n18 = ( n676  &  n677  &  n678  &  n679  &  n680  &  n681  &  n682  &  n683 ) ;
 assign n23 = ( n454  &  n69 ) | ( n60  &  n69 ) | ( n454  &  n450 ) | ( n60  &  n450 ) ;
 assign n24 = ( n70 ) | ( n92 ) ;
 assign n25 = ( n397  &  n445  &  (~ n447)  &  n758 ) ;
 assign n26 = ( n58 ) | ( n345 ) ;
 assign n27 = ( n401  &  n400 ) | ( n491  &  n400 ) | ( n401  &  n324 ) | ( n491  &  n324 ) ;
 assign n19 = ( n23  &  n24  &  n25  &  n26  &  n27  &  (~ n462)  &  (~ n465)  &  (~ n468) ) ;
 assign n29 = ( n93 ) | ( n696 ) | ( j ) | ( n249 ) ;
 assign n32 = ( n801  &  n164 ) | ( n454  &  n164 ) | ( n801  &  n400 ) | ( n454  &  n400 ) ;
 assign n33 = ( n69  &  (~ n316) ) | ( n260  &  (~ n316) ) | ( (~ n316)  &  n320 ) ;
 assign n34 = ( n678  &  n207  &  n40  &  n723  &  n724  &  n676  &  n725  &  n726 ) ;
 assign n35 = ( (~ n484)  &  n696 ) | ( (~ n484)  &  n839  &  n840 ) ;
 assign n28 = ( n25  &  n29  &  n32  &  n33  &  n34  &  n35  &  (~ n479)  &  (~ n482) ) ;
 assign n40 = ( n451 ) | ( n64 ) | ( n65 ) ;
 assign n41 = ( n700 ) | ( n65 ) ;
 assign n42 = ( (~ d) ) | ( n252 ) | ( n274 ) ;
 assign n43 = ( n823  &  n235 ) | ( n823  &  n52 ) ;
 assign n44 = ( n229  &  n136 ) | ( n229  &  n739 ) ;
 assign n36 = ( n40  &  n41  &  n42  &  n43  &  n44  &  (~ n275)  &  (~ n278)  &  (~ n281) ) ;
 assign n46 = ( (~ h) ) | ( (~ k) ) ;
 assign n45 = ( n46 ) | ( l ) ;
 assign n49 = ( n730 ) | ( (~ n769) ) ;
 assign n47 = ( n49  &  (~ n154) ) | ( (~ n154)  &  (~ n684) ) ;
 assign n52 = ( (~ c) ) | ( n526 ) ;
 assign n53 = ( e ) | ( n605 ) ;
 assign n54 = ( n717  &  n327 ) ;
 assign n51 = ( n52  &  n53  &  n54 ) ;
 assign n58 = ( (~ k) ) | ( n192 ) ;
 assign n57 = ( j ) | ( (~ l) ) | ( m ) ;
 assign n55 = ( (~ n)  &  n58 ) | ( n58  &  n57 ) ;
 assign n61 = ( n801 ) | ( n58 ) ;
 assign n62 = ( n198  &  n184 ) | ( n709  &  n184 ) | ( n198  &  n710 ) | ( n709  &  n710 ) ;
 assign n60 = ( (~ g) ) | ( n708 ) ;
 assign n59 = ( n61  &  n62  &  n55 ) | ( n61  &  n62  &  n60 ) ;
 assign n66 = ( n86  &  n84 ) | ( n295  &  n84 ) | ( n86  &  n144 ) | ( n295  &  n144 ) ;
 assign n64 = ( (~ i) ) | ( n628 ) ;
 assign n65 = ( (~ a) ) | ( n605 ) ;
 assign n63 = ( n66  &  n64 ) | ( n66  &  n65 ) ;
 assign n68 = ( (~ g) ) | ( n705 ) ;
 assign n69 = ( n307  &  n441 ) ;
 assign n70 = ( (~ k) ) | ( n154 ) ;
 assign n67 = ( n68 ) | ( n69 ) | ( n70 ) ;
 assign n73 = ( n706 ) | ( n192 ) ;
 assign n72 = ( (~ i) ) | ( n409 ) ;
 assign n71 = ( (~ n)  &  n73 ) | ( n73  &  n72 ) ;
 assign n75 = ( (~ h) ) | ( n628 ) ;
 assign n76 = ( (~ n) ) | ( n103 ) ;
 assign n77 = ( h ) | ( n628 ) ;
 assign n74 = ( n75  &  n71 ) | ( n76  &  n71 ) | ( n75  &  n77 ) | ( n76  &  n77 ) ;
 assign n79 = ( (~ g) ) | ( n256 ) ;
 assign n80 = ( h ) | ( n190 ) ;
 assign n78 = ( n76  &  n71 ) | ( n79  &  n71 ) | ( n76  &  n80 ) | ( n79  &  n80 ) ;
 assign n82 = ( (~ k) ) | ( n168 ) ;
 assign n81 = ( n82  &  n ) | ( n82  &  n57 ) ;
 assign n84 = ( n306  &  n712  &  n713 ) ;
 assign n83 = ( n84  &  n75 ) | ( n79  &  n75 ) | ( n84  &  n65 ) | ( n79  &  n65 ) ;
 assign n88 = ( n109 ) | ( n93 ) ;
 assign n86 = ( n214  &  n315 ) ;
 assign n87 = ( (~ g) ) | ( n437 ) ;
 assign n85 = ( n88  &  n83  &  n86 ) | ( n88  &  n83  &  n87 ) ;
 assign n91 = ( n86  &  n84 ) | ( n180  &  n84 ) | ( n86  &  n152 ) | ( n180  &  n152 ) ;
 assign n90 = ( e ) | ( n714 ) ;
 assign n89 = ( n91  &  n65 ) | ( n91  &  n90 ) ;
 assign n93 = ( (~ a) ) | ( n290 ) ;
 assign n94 = ( (~ e) ) | ( n714 ) ;
 assign n92 = ( n89  &  n93 ) | ( n89  &  n94 ) ;
 assign n96 = ( n86  &  n84 ) | ( n195  &  n84 ) | ( n86  &  n80 ) | ( n195  &  n80 ) ;
 assign n95 = ( n96  &  n65 ) | ( n96  &  n77 ) ;
 assign n100 = ( n142 ) | ( n443 ) ;
 assign n101 = ( (~ g) ) | ( n241 ) | ( (~ n715) ) ;
 assign n98 = ( j ) | ( n141 ) ;
 assign n99 = ( (~ i) ) | ( n714 ) ;
 assign n97 = ( n100  &  n101  &  n98 ) | ( n100  &  n101  &  n99 ) ;
 assign n103 = ( n612  &  n911  &  n596  &  n446 ) ;
 assign n102 = ( n103  &  n80 ) | ( n79  &  n80 ) | ( n103  &  n72 ) | ( n79  &  n72 ) ;
 assign n106 = ( (~ i) ) | ( n92 ) | ( n603 ) ;
 assign n107 = ( n69  &  n95 ) | ( n97  &  n95 ) | ( n69  &  n693 ) | ( n97  &  n693 ) ;
 assign n105 = ( (~ e) ) | ( n290 ) ;
 assign n104 = ( n106  &  n107  &  n102 ) | ( n106  &  n107  &  n105 ) ;
 assign n109 = ( (~ h) ) | ( n249 ) ;
 assign n110 = ( h ) | ( n249 ) ;
 assign n108 = ( n109  &  n71 ) | ( n76  &  n71 ) | ( n109  &  n110 ) | ( n76  &  n110 ) ;
 assign n111 = ( (~ n108)  &  (~ n732) ) | ( b  &  (~ n108)  &  (~ n554) ) ;
 assign n115 = ( (~ n59)  &  (~ n351) ) | ( (~ n59)  &  (~ n711) ) ;
 assign n119 = ( (~ n154)  &  (~ n797) ) | ( (~ n92)  &  (~ n154)  &  (~ n706) ) ;
 assign n123 = ( (~ n69)  &  (~ n803) ) | ( (~ n69)  &  (~ n70)  &  (~ n99) ) ;
 assign n130 = ( n168 ) | ( n80 ) | ( n105 ) | ( n706 ) ;
 assign n131 = ( n695 ) | ( n696 ) ;
 assign n132 = ( n692 ) | ( n693 ) | ( n110 ) ;
 assign n133 = ( n  &  (~ n115)  &  (~ n119) ) | ( n104  &  (~ n115)  &  (~ n119) ) ;
 assign n134 = ( n74  &  n63 ) | ( n722  &  n63 ) | ( n74  &  n696 ) | ( n722  &  n696 ) ;
 assign n135 = ( n806  &  n78 ) | ( n806  &  n287 ) ;
 assign n128 = ( n34  &  (~ n111)  &  n130  &  n131  &  n132  &  n133  &  n134  &  n135 ) ;
 assign n138 = ( n808 ) | ( n82 ) ;
 assign n139 = ( n718  &  n413 ) | ( n731  &  n413 ) | ( n718  &  n185 ) | ( n731  &  n185 ) ;
 assign n137 = ( (~ f) ) | ( n708 ) ;
 assign n136 = ( n138  &  n139  &  n81 ) | ( n138  &  n139  &  n137 ) ;
 assign n142 = ( (~ m) ) | ( n716 ) ;
 assign n141 = ( (~ l) ) | ( (~ m) ) ;
 assign n140 = ( n142  &  i ) | ( n142  &  n141 ) ;
 assign n144 = ( (~ i) ) | ( n190 ) ;
 assign n145 = ( j ) | ( n190 ) ;
 assign n143 = ( n144  &  n145 ) ;
 assign n149 = ( n143  &  n140 ) | ( n694  &  n140 ) | ( n143  &  n79 ) | ( n694  &  n79 ) ;
 assign n150 = ( n809  &  n152 ) | ( n809  &  n98 ) ;
 assign n147 = ( n752  &  n755 ) ;
 assign n148 = ( i ) | ( n190 ) ;
 assign n146 = ( n149  &  n150  &  n147 ) | ( n149  &  n150  &  n148 ) ;
 assign n152 = ( g ) | ( n256 ) ;
 assign n151 = ( n  &  n152 ) | ( n146  &  n152 ) | ( n  &  n70 ) | ( n146  &  n70 ) ;
 assign n156 = ( (~ m) ) | ( n ) | ( n46 ) ;
 assign n154 = ( (~ m) ) | ( n ) ;
 assign n155 = ( (~ h) ) | ( j ) | ( (~ l) ) ;
 assign n153 = ( n156  &  n154 ) | ( n156  &  n155 ) ;
 assign n159 = ( (~ f) ) | ( n249 ) ;
 assign n160 = ( (~ e) ) | ( n189 ) ;
 assign n157 = ( (~ n47)  &  n153 ) | ( n153  &  n159 ) | ( (~ n47)  &  n160 ) | ( n159  &  n160 ) ;
 assign n163 = ( d ) | ( n153 ) | ( n189 ) ;
 assign n162 = ( d ) | ( n190 ) ;
 assign n161 = ( (~ n47)  &  n163 ) | ( n163  &  n162 ) ;
 assign n165 = ( j ) | ( n46 ) ;
 assign n164 = ( n165  &  i ) | ( n165  &  n46 ) ;
 assign n167 = ( n45  &  n164  &  n324  &  n323 ) ;
 assign n168 = ( m ) | ( n ) ;
 assign n169 = ( j ) | ( n708 ) ;
 assign n170 = ( (~ l) ) | ( n168 ) ;
 assign n166 = ( n167  &  n169 ) | ( n168  &  n169 ) | ( n167  &  n170 ) | ( n168  &  n170 ) ;
 assign n172 = ( (~ e) ) | ( n721 ) ;
 assign n173 = ( (~ n) ) | ( n172 ) ;
 assign n171 = ( n73  &  n72 ) | ( n172  &  n72 ) | ( n73  &  n173 ) | ( n172  &  n173 ) ;
 assign n174 = ( (~ n87)  &  (~ n173)  &  (~ n912) ) | ( (~ n173)  &  (~ n180)  &  (~ n912) ) ;
 assign n182 = ( n171  &  (~ n174) ) | ( (~ n174)  &  n195  &  n789 ) ;
 assign n181 = ( n172 ) | ( n435 ) ;
 assign n180 = ( g ) | ( n437 ) ;
 assign n179 = ( n182  &  n181 ) | ( n182  &  n87  &  n180 ) ;
 assign n186 = ( n808  &  n198 ) | ( n58  &  n198 ) | ( n808  &  n731 ) | ( n58  &  n731 ) ;
 assign n184 = ( k ) | ( n192 ) ;
 assign n185 = ( (~ j) ) | ( n256 ) ;
 assign n183 = ( n186  &  n184 ) | ( n186  &  n185 ) ;
 assign n187 = ( n183  &  n55 ) | ( n183  &  n137 ) ;
 assign n189 = ( (~ f) ) | ( g ) ;
 assign n190 = ( (~ f) ) | ( (~ g) ) ;
 assign n188 = ( (~ n47)  &  n153 ) | ( (~ n47)  &  n189 ) | ( n153  &  n190 ) | ( n189  &  n190 ) ;
 assign n192 = ( m ) | ( (~ n) ) ;
 assign n193 = ( (~ l) ) | ( n192 ) ;
 assign n191 = ( n167  &  n169 ) | ( n192  &  n169 ) | ( n167  &  n193 ) | ( n192  &  n193 ) ;
 assign n195 = ( h ) | ( n675 ) ;
 assign n194 = ( n76  &  n71 ) | ( n87  &  n71 ) | ( n76  &  n195 ) | ( n87  &  n195 ) ;
 assign n196 = ( n194  &  n191 ) | ( n194  &  n159  &  n160 ) ;
 assign n200 = ( n810  &  n811  &  n55 ) | ( n810  &  n811  &  n342 ) ;
 assign n198 = ( l ) | ( n192 ) ;
 assign n199 = ( (~ k) ) | ( n437 ) ;
 assign n197 = ( n59  &  n200  &  n198 ) | ( n59  &  n200  &  n199 ) ;
 assign n201 = ( (~ n105)  &  (~ n136) ) | ( (~ n136)  &  (~ n495) ) ;
 assign n206 = ( n700 ) | ( n704 ) ;
 assign n207 = ( n700 ) | ( n391 ) ;
 assign n208 = ( (~ e)  &  n813 ) | ( n187  &  n813 ) | ( n352  &  n813 ) ;
 assign n209 = ( (~ n201)  &  n307 ) | ( n151  &  (~ n201)  &  n700 ) ;
 assign n210 = ( n197 ) | ( n343 ) ;
 assign n211 = ( n161  &  n157 ) | ( n306  &  n157 ) | ( n161  &  n93 ) | ( n306  &  n93 ) ;
 assign n212 = ( n815  &  n166 ) | ( n815  &  n327 ) ;
 assign n205 = ( n206  &  n207  &  n208  &  n209  &  n210  &  n211  &  n179  &  n212 ) ;
 assign n214 = ( (~ a) ) | ( n665 ) ;
 assign n215 = ( n154 ) | ( n214 ) ;
 assign n213 = ( n214  &  n155 ) | ( n156  &  n155 ) | ( n214  &  n215 ) | ( n156  &  n215 ) ;
 assign n219 = ( (~ n684) ) | ( n730 ) | ( (~ n769) ) ;
 assign n218 = ( (~ f)  &  (~ n628) ) ;
 assign n216 = ( (~ n215)  &  n219  &  n218 ) | ( (~ n215)  &  n219  &  (~ n268) ) ;
 assign n222 = ( e ) | ( n564 ) ;
 assign n223 = ( e ) | ( n189 ) ;
 assign n221 = ( n213  &  (~ n216) ) | ( (~ n216)  &  n222  &  n223 ) ;
 assign n227 = ( (~ j) ) | ( n413 ) | ( n437 ) ;
 assign n228 = ( n81  &  n718 ) | ( n342  &  n718 ) | ( n81  &  n199 ) | ( n342  &  n199 ) ;
 assign n226 = ( n748  &  n751 ) ;
 assign n225 = ( n227  &  n228  &  n226 ) | ( n227  &  n228  &  n82 ) ;
 assign n230 = ( (~ e) ) | ( n733 ) ;
 assign n229 = ( n179  &  n221  &  n225 ) | ( n179  &  n221  &  n230 ) ;
 assign n231 = ( (~ n58)  &  (~ n259) ) | ( (~ n58)  &  (~ n747) ) ;
 assign n238 = ( n262  &  n184 ) | ( n198  &  n184 ) | ( n262  &  n348 ) | ( n198  &  n348 ) ;
 assign n236 = ( g ) | ( n708 ) ;
 assign n235 = ( n55  &  (~ n231)  &  n238 ) | ( (~ n231)  &  n238  &  n236 ) ;
 assign n241 = ( k ) | ( n141 ) ;
 assign n239 = ( i  &  (~ j) ) | ( (~ j)  &  n147 ) | ( i  &  n241 ) | ( n147  &  n241 ) ;
 assign n242 = ( (~ n64)  &  (~ n696) ) | ( (~ j)  &  (~ n628)  &  (~ n696) ) ;
 assign n247 = ( n  &  (~ n242) ) | ( (~ n242)  &  n820  &  n821 ) ;
 assign n246 = ( n151  &  n247  &  n70 ) | ( n151  &  n247  &  n90 ) ;
 assign n250 = ( (~ i) ) | ( n249 ) ;
 assign n249 = ( (~ e) ) | ( (~ g) ) ;
 assign n248 = ( n250  &  j ) | ( n250  &  n249 ) ;
 assign n251 = ( n70 ) | ( n94 ) ;
 assign n253 = ( n818  &  n94 ) | ( n818  &  n98 ) ;
 assign n254 = ( n817  &  n816  &  n248 ) | ( n817  &  n816  &  n694 ) ;
 assign n252 = ( n251  &  n ) | ( n251  &  n253  &  n254 ) ;
 assign n256 = ( (~ f) ) | ( (~ h) ) ;
 assign n255 = ( n76 ) | ( e ) | ( n256 ) ;
 assign n258 = ( n736  &  n60 ) ;
 assign n259 = ( j ) | ( n714 ) ;
 assign n260 = ( i ) | ( n707 ) ;
 assign n261 = ( (~ g) ) | ( n398 ) ;
 assign n257 = ( n258  &  n259  &  n260  &  n261 ) ;
 assign n262 = ( g ) | ( n46 ) ;
 assign n265 = ( n819  &  n415 ) | ( n819  &  n735  &  n759 ) ;
 assign n266 = ( n736  &  n68 ) | ( n737  &  n68 ) | ( n736  &  n70 ) | ( n737  &  n70 ) ;
 assign n264 = ( (~ l) ) | ( n154 ) ;
 assign n263 = ( n265  &  n266  &  n257 ) | ( n265  &  n266  &  n264 ) ;
 assign n268 = ( (~ f) ) | ( n628 ) ;
 assign n267 = ( (~ n47)  &  n153 ) | ( (~ n47)  &  n223 ) | ( n153  &  n268 ) | ( n223  &  n268 ) ;
 assign n269 = ( (~ n263)  &  (~ n765) ) | ( d  &  (~ n263)  &  (~ n609) ) ;
 assign n274 = ( a ) | ( (~ b) ) ;
 assign n275 = ( (~ n191)  &  (~ n351) ) | ( (~ n191)  &  (~ n268)  &  (~ n722) ) ;
 assign n278 = ( (~ n267)  &  (~ n390) ) | ( n269  &  (~ n390) ) ;
 assign n281 = ( (~ n255)  &  (~ n610) ) | ( (~ n71)  &  (~ n610)  &  (~ n738) ) ;
 assign n288 = ( n381  &  n58 ) | ( n381  &  n740 ) ;
 assign n287 = ( (~ b) ) | ( n703 ) ;
 assign n286 = ( n288  &  n183 ) | ( n288  &  n287 ) ;
 assign n290 = ( (~ c) ) | ( d ) ;
 assign n289 = ( (~ f)  &  n52 ) | ( n52  &  n290 ) ;
 assign n293 = ( n152  &  n71 ) | ( n76  &  n71 ) | ( n152  &  n742 ) | ( n76  &  n742 ) ;
 assign n292 = ( n293  &  n78 ) ;
 assign n295 = ( (~ i) ) | ( n675 ) ;
 assign n296 = ( j ) | ( n675 ) ;
 assign n294 = ( n295  &  n296 ) ;
 assign n299 = ( n294  &  n140 ) | ( n694  &  n140 ) | ( n294  &  n87 ) | ( n694  &  n87 ) ;
 assign n300 = ( n896  &  n180 ) | ( n896  &  n98 ) ;
 assign n298 = ( i ) | ( n675 ) ;
 assign n297 = ( n299  &  n300  &  n147 ) | ( n299  &  n300  &  n298 ) ;
 assign n301 = ( n  &  n70 ) | ( n297  &  n70 ) | ( n  &  n180 ) | ( n297  &  n180 ) ;
 assign n303 = ( g ) | ( n153 ) | ( n305 ) ;
 assign n302 = ( d  &  n303 ) | ( (~ n47)  &  n303 ) | ( n249  &  n303 ) ;
 assign n307 = ( (~ e) ) | ( n274 ) ;
 assign n305 = ( d ) | ( (~ e) ) ;
 assign n306 = ( (~ a) ) | ( (~ b) ) | ( c ) ;
 assign n304 = ( n307  &  n305 ) | ( n307  &  n306 ) ;
 assign n309 = ( n74  &  n235 ) | ( n722  &  n235 ) | ( n74  &  n743 ) | ( n722  &  n743 ) ;
 assign n310 = ( n263  &  n302 ) | ( n302  &  n304 ) | ( n263  &  (~ n644) ) | ( n304  &  (~ n644) ) ;
 assign n311 = ( n78 ) | ( n343 ) ;
 assign n312 = ( n292  &  n166 ) | ( n732  &  n166 ) | ( n292  &  n289 ) | ( n732  &  n289 ) ;
 assign n308 = ( n286  &  n229  &  n309  &  n310  &  n311  &  n312 ) ;
 assign n313 = ( n95  &  n93 ) | ( n95  &  n110 ) ;
 assign n315 = ( n701  &  n699 ) ;
 assign n314 = ( n88  &  n83  &  n315 ) | ( n88  &  n83  &  n87 ) ;
 assign n316 = ( (~ n395)  &  (~ n744) ) | ( (~ n154)  &  (~ n314)  &  (~ n744) ) ;
 assign n320 = ( n ) | ( n98 ) ;
 assign n323 = ( (~ h) ) | ( n398 ) ;
 assign n324 = ( (~ k) ) | ( n708 ) ;
 assign n322 = ( n323  &  n165  &  n324  &  n169 ) ;
 assign n327 = ( (~ c) ) | ( n609 ) ;
 assign n325 = ( (~ c)  &  n327 ) | ( n189  &  n327 ) ;
 assign n330 = ( (~ j)  &  n86 ) | ( n86  &  n753 ) | ( (~ j)  &  n754 ) | ( n753  &  n754 ) ;
 assign n329 = ( (~ j) ) | ( n190 ) ;
 assign n328 = ( n330  &  n84 ) | ( n330  &  n329 ) ;
 assign n331 = ( n92  &  n69 ) | ( n92  &  n68 ) ;
 assign n332 = ( (~ n60)  &  (~ n69)  &  (~ n752) ) | ( (~ n69)  &  (~ n752)  &  (~ n771) ) ;
 assign n338 = ( (~ n332)  &  n357 ) | ( (~ n332)  &  n372 ) | ( (~ n332)  &  n500 ) ;
 assign n339 = ( n328  &  n89 ) | ( n241  &  n89 ) | ( n328  &  n98 ) | ( n241  &  n98 ) ;
 assign n337 = ( (~ l) ) | ( n603 ) ;
 assign n336 = ( n338  &  n339  &  n331 ) | ( n338  &  n339  &  n337 ) ;
 assign n341 = ( n172  &  n434 ) ;
 assign n342 = ( f ) | ( n708 ) ;
 assign n343 = ( (~ b) ) | ( n305 ) ;
 assign n340 = ( n341  &  n342 ) | ( n236  &  n342 ) | ( n341  &  n343 ) | ( n236  &  n343 ) ;
 assign n345 = ( n740  &  n340 ) ;
 assign n346 = ( (~ n)  &  n53 ) | ( n  &  n412 ) | ( n53  &  n412 ) ;
 assign n344 = ( (~ n)  &  n60 ) | ( n60  &  n345 ) | ( (~ n)  &  n346 ) | ( n345  &  n346 ) ;
 assign n349 = ( (~ j) ) | ( n343 ) | ( n437 ) ;
 assign n350 = ( n287 ) | ( n185 ) ;
 assign n348 = ( (~ j) ) | ( n714 ) ;
 assign n347 = ( n349  &  n350  &  n341 ) | ( n349  &  n350  &  n348 ) ;
 assign n352 = ( b ) | ( (~ c) ) ;
 assign n351 = ( (~ f) ) | ( n352 ) ;
 assign n355 = ( n341  &  n343 ) | ( n259  &  n343 ) | ( n341  &  n751 ) | ( n259  &  n751 ) ;
 assign n354 = ( j ) | ( n256 ) ;
 assign n353 = ( n355  &  n287 ) | ( n355  &  n354 ) ;
 assign n357 = ( (~ h) ) | ( n727 ) ;
 assign n356 = ( n353  &  n351 ) | ( n353  &  n357 ) ;
 assign n360 = ( n356  &  n340 ) | ( n500  &  n340 ) | ( n356  &  n57 ) | ( n500  &  n57 ) ;
 assign n359 = ( k ) | ( (~ l) ) | ( m ) ;
 assign n358 = ( n360  &  n347 ) | ( n360  &  n359 ) ;
 assign n363 = ( n341  &  n343 ) | ( n747  &  n343 ) | ( n341  &  n748 ) | ( n747  &  n748 ) ;
 assign n362 = ( i ) | ( n256 ) ;
 assign n361 = ( n363  &  n287 ) | ( n363  &  n362 ) ;
 assign n364 = ( (~ n192)  &  (~ n361) ) | ( (~ n192)  &  (~ n260)  &  (~ n412) ) ;
 assign n369 = ( n53  &  (~ n364) ) | ( n168  &  (~ n364) ) | ( n260  &  (~ n364) ) ;
 assign n372 = ( n325  &  n745 ) ;
 assign n371 = ( n351  &  n372 ) | ( n193  &  n372 ) | ( n351  &  n170 ) | ( n193  &  n170 ) ;
 assign n373 = ( (~ n346)  &  (~ n831) ) | ( (~ n346)  &  (~ n359)  &  (~ n710) ) ;
 assign n379 = ( (~ j) ) | ( n93 ) | ( n249 ) | ( n566 ) ;
 assign n380 = ( n93 ) | ( n94 ) | ( n320 ) ;
 assign n381 = ( (~ n) ) | ( n57 ) | ( n740 ) ;
 assign n382 = ( n833  &  n322 ) | ( n833  &  n371 ) ;
 assign n383 = ( n33  &  n344 ) | ( n33  &  n500 ) ;
 assign n384 = ( (~ n)  &  n336 ) | ( n  &  n358 ) | ( n336  &  n358 ) ;
 assign n385 = ( n369  &  n798 ) | ( n498  &  n798 ) | ( n369  &  n749 ) | ( n498  &  n749 ) ;
 assign n378 = ( (~ n373)  &  n379  &  n380  &  n381  &  n382  &  n383  &  n384  &  n385 ) ;
 assign n388 = ( i  &  n86 ) | ( n753  &  n86 ) | ( i  &  n298 ) | ( n753  &  n298 ) ;
 assign n387 = ( n388  &  n84 ) | ( n388  &  n148 ) ;
 assign n390 = ( (~ a) ) | ( n352 ) ;
 assign n391 = ( (~ b) ) | ( n702 ) ;
 assign n389 = ( n306  &  n390  &  n391 ) ;
 assign n395 = ( n87 ) | ( n215 ) ;
 assign n393 = ( n315  &  n704 ) | ( n87  &  n704 ) | ( n315  &  n79 ) | ( n87  &  n79 ) ;
 assign n394 = ( n88  &  n65 ) | ( n88  &  n79  &  n75 ) ;
 assign n392 = ( n395  &  n154 ) | ( n395  &  n393  &  n394 ) ;
 assign n399 = ( n836  &  n307 ) | ( n836  &  n737 ) | ( n836  &  n710 ) ;
 assign n398 = ( (~ j) ) | ( k ) ;
 assign n397 = ( n399  &  n392 ) | ( n399  &  n398 ) ;
 assign n400 = ( n351  &  n372 ) | ( n192  &  n372 ) | ( n351  &  n168 ) | ( n192  &  n168 ) ;
 assign n401 = ( n351  &  n372 ) | ( n58  &  n372 ) | ( n351  &  n82 ) | ( n58  &  n82 ) ;
 assign n402 = ( (~ n60)  &  (~ n834) ) | ( (~ n60)  &  (~ n154)  &  (~ n498) ) ;
 assign n406 = ( (~ n402)  &  n736 ) | ( n264  &  (~ n402)  &  n737 ) ;
 assign n405 = ( n406  &  n70 ) | ( n406  &  n348 ) ;
 assign n410 = ( n ) | ( n92 ) | ( n603 ) ;
 assign n409 = ( (~ k) ) | ( m ) ;
 assign n408 = ( (~ n)  &  n260 ) | ( (~ n)  &  n346 ) | ( n260  &  n361 ) | ( n346  &  n361 ) ;
 assign n407 = ( n410  &  n409 ) | ( n410  &  n408  &  n344 ) ;
 assign n412 = ( n343  &  n711  &  n439 ) ;
 assign n413 = ( k ) | ( n168 ) ;
 assign n411 = ( n412  &  n413 ) | ( n184  &  n413 ) | ( n412  &  n53 ) | ( n184  &  n53 ) ;
 assign n417 = ( (~ i) ) | ( k ) | ( (~ l) ) | ( n154 ) ;
 assign n416 = ( (~ k) ) | ( (~ n715) ) ;
 assign n415 = ( l ) | ( n154 ) ;
 assign n414 = ( n417  &  n416 ) | ( n417  &  n415  &  n264 ) ;
 assign n419 = ( (~ j) ) | ( n708 ) ;
 assign n418 = ( n419  &  n357 ) ;
 assign n421 = ( n692 ) | ( n734 ) | ( n752 ) ;
 assign n422 = ( n692 ) | ( n734 ) | ( n755 ) ;
 assign n423 = ( n ) | ( n147 ) | ( n387 ) ;
 assign n424 = ( n401  &  n313 ) | ( n418  &  n313 ) | ( n401  &  n414 ) | ( n418  &  n414 ) ;
 assign n425 = ( n411 ) | ( n710 ) ;
 assign n426 = ( (~ j)  &  n69 ) | ( (~ j)  &  n405 ) | ( n69  &  n407 ) | ( n405  &  n407 ) ;
 assign n427 = ( n400 ) | ( n323 ) ;
 assign n428 = ( n397  &  n347 ) | ( n397  &  n184 ) ;
 assign n420 = ( n421  &  n422  &  n423  &  n424  &  n425  &  n426  &  n427  &  n428 ) ;
 assign n429 = ( (~ n325)  &  (~ n413) ) | ( (~ n413)  &  (~ n745) ) ;
 assign n434 = ( n743  &  n746 ) ;
 assign n435 = ( (~ n) ) | ( n446 ) ;
 assign n433 = ( n181  &  n434 ) | ( n181  &  n435 ) ;
 assign n437 = ( f ) | ( (~ h) ) ;
 assign n436 = ( n256  &  n437 ) | ( n287  &  n437 ) | ( n256  &  n343 ) | ( n287  &  n343 ) ;
 assign n439 = ( n722  &  n732 ) ;
 assign n440 = ( e ) | ( n352 ) ;
 assign n441 = ( (~ b) ) | ( n609 ) ;
 assign n438 = ( n439  &  n343  &  n440  &  n441 ) ;
 assign n443 = ( (~ i) ) | ( n707 ) ;
 assign n442 = ( (~ i)  &  n438 ) | ( n436  &  n438 ) | ( (~ i)  &  n443 ) | ( n436  &  n443 ) ;
 assign n446 = ( m ) | ( n398 ) ;
 assign n445 = ( n53 ) | ( n446 ) | ( n443 ) | ( n ) ;
 assign n449 = ( h  &  n715 ) ;
 assign n447 = ( n429  &  n449 ) | ( (~ n184)  &  (~ n351)  &  n449 ) ;
 assign n452 = ( n260 ) | ( n749 ) ;
 assign n453 = ( n415  &  n262 ) | ( n165  &  n262 ) | ( n415  &  n154 ) | ( n165  &  n154 ) ;
 assign n451 = ( n ) | ( n697 ) ;
 assign n450 = ( n452  &  n453  &  n451 ) | ( n452  &  n453  &  n443 ) ;
 assign n454 = ( n412  &  n82 ) | ( n58  &  n82 ) | ( n412  &  n53 ) | ( n58  &  n53 ) ;
 assign n455 = ( i  &  (~ n436) ) ;
 assign n457 = ( n  &  n455 ) | ( n  &  (~ n99)  &  (~ n341) ) ;
 assign n461 = ( j ) | ( i ) ;
 assign n459 = ( (~ k) ) | ( n264 ) | ( n461 ) ;
 assign n462 = ( (~ n85)  &  (~ n459) ) | ( n49  &  (~ n85)  &  (~ n154) ) ;
 assign n465 = ( n457  &  (~ n612) ) | ( (~ n346)  &  (~ n443)  &  (~ n612) ) ;
 assign n468 = ( (~ n696)  &  (~ n838) ) | ( (~ n84)  &  (~ n354)  &  (~ n696) ) ;
 assign n472 = ( (~ n387)  &  (~ n498) ) | ( (~ n93)  &  (~ n498)  &  (~ n734) ) ;
 assign n476 = ( (~ n)  &  (~ n258)  &  (~ n337) ) ;
 assign n479 = ( (~ n69)  &  n476 ) | ( (~ n69)  &  (~ n415)  &  (~ n759) ) ;
 assign n482 = ( (~ n58)  &  (~ n353) ) | ( (~ n58)  &  (~ n361) ) ;
 assign n485 = ( i  &  k ) ;
 assign n484 = ( (~ n154)  &  n472 ) | ( (~ n154)  &  (~ n313)  &  n485 ) ;
 assign n488 = ( (~ f) ) | ( n703 ) | ( n764 ) ;
 assign n489 = ( j ) | ( k ) ;
 assign n487 = ( n488 ) | ( n489 ) | ( n264 ) | ( n443 ) ;
 assign n491 = ( (~ h) ) | ( n705 ) ;
 assign n492 = ( (~ n) ) | ( n659 ) | ( n761 ) ;
 assign n490 = ( n491 ) | ( n359 ) | ( n492 ) ;
 assign n494 = ( n87 ) | ( n170 ) | ( n760 ) ;
 assign n495 = ( (~ e) ) | ( n605 ) ;
 assign n493 = ( n494 ) | ( n495 ) ;
 assign n497 = ( (~ n644) ) | ( n765 ) ;
 assign n498 = ( (~ j) ) | ( (~ k) ) | ( (~ l) ) ;
 assign n496 = ( n497 ) | ( n498 ) | ( n443 ) | ( n154 ) ;
 assign n500 = ( (~ l) ) | ( n409 ) ;
 assign n501 = ( n159 ) | ( n610 ) ;
 assign n499 = ( (~ n449) ) | ( n500 ) | ( n501 ) ;
 assign n504 = ( n170 ) | ( n416 ) ;
 assign n503 = ( n230 ) | ( n79 ) | ( n504 ) ;
 assign n505 = ( n195 ) | ( n739 ) | ( n762 ) ;
 assign n506 = ( n500 ) | ( n510 ) | ( (~ n763) ) ;
 assign n507 = ( n170 ) | ( n195 ) | ( n495 ) | ( (~ n545) ) ;
 assign n508 = ( n842  &  n359 ) | ( n842  &  n492 ) | ( n842  &  n419 ) ;
 assign n512 = ( n230 ) | ( n769 ) | ( n80 ) | ( n718 ) ;
 assign n510 = ( h ) | ( n727 ) ;
 assign n511 = ( k ) | ( l ) | ( m ) ;
 assign n509 = ( n512  &  n501 ) | ( n512  &  n510 ) | ( n512  &  n511 ) ;
 assign n514 = ( n ) | ( n511 ) | ( n653 ) ;
 assign n513 = ( n514  &  n168 ) | ( n514  &  n99 ) | ( n514  &  n498 ) ;
 assign n516 = ( n170 ) | ( n739 ) | ( k ) | ( n180 ) ;
 assign n517 = ( (~ h) ) | ( n222 ) | ( n359 ) | ( n761 ) ;
 assign n515 = ( n516  &  n517 ) ;
 assign n519 = ( n771 ) | ( n552 ) | ( n749 ) | ( n764 ) ;
 assign n520 = ( n651 ) | ( n760 ) | ( n79 ) | ( n170 ) ;
 assign n521 = ( n515  &  n513 ) | ( n461  &  n513 ) | ( n515  &  n553 ) | ( n461  &  n553 ) ;
 assign n518 = ( n15  &  n509  &  n12  &  n519  &  n520  &  n521 ) ;
 assign n522 = ( i ) | ( n168 ) ;
 assign n523 = ( (~ k)  &  n168 ) | ( (~ k)  &  (~ n461) ) | ( n168  &  n522 ) | ( (~ n461)  &  n522 ) ;
 assign n526 = ( e ) | ( (~ f) ) ;
 assign n527 = ( a ) | ( n610 ) ;
 assign n525 = ( j  &  n526  &  (~ n737) ) | ( j  &  n527  &  (~ n737) ) ;
 assign n532 = ( (~ h)  &  (~ n906) ) | ( n504  &  (~ n906) ) | ( (~ n554)  &  (~ n906) ) ;
 assign n530 = ( (~ c) ) | ( e ) | ( f ) ;
 assign n529 = ( n523  &  (~ n525)  &  n532 ) | ( (~ n525)  &  n532  &  n530 ) ;
 assign n534 = ( b ) | ( n192 ) ;
 assign n533 = ( n534  &  n320  &  n58  &  n193 ) ;
 assign n535 = ( c  &  b ) | ( n170  &  b ) | ( c  &  n193 ) | ( n170  &  n193 ) ;
 assign n536 = ( (~ n154)  &  (~ n875) ) | ( (~ b)  &  (~ n154)  &  (~ n554) ) ;
 assign n542 = ( j ) | ( n192 ) | ( h ) ;
 assign n543 = ( (~ i)  &  j ) | ( (~ i)  &  n58 ) | ( j  &  n774 ) | ( n58  &  n774 ) ;
 assign n541 = ( (~ j) ) | ( n192 ) ;
 assign n539 = ( (~ h)  &  n542  &  n543 ) | ( n542  &  n543  &  n541 ) ;
 assign n545 = ( (~ k)  &  n715 ) ;
 assign n544 = ( b  &  (~ n192)  &  n545 ) ;
 assign n546 = ( (~ h)  &  n544 ) | ( (~ h)  &  (~ i)  &  (~ n198) ) ;
 assign n548 = ( (~ n605)  &  (~ n785) ) | ( (~ e)  &  n352  &  (~ n785) ) ;
 assign n552 = ( f ) | ( n770 ) ;
 assign n551 = ( n552  &  f ) | ( n552  &  a ) | ( n552  &  e ) ;
 assign n554 = ( c ) | ( d ) ;
 assign n553 = ( f ) | ( n554 ) ;
 assign n556 = ( c ) | ( e ) | ( n780 ) ;
 assign n558 = ( b ) | ( e ) | ( (~ n) ) | ( n780 ) ;
 assign n559 = ( (~ h) ) | ( n264 ) | ( n416 ) | ( (~ n721) ) ;
 assign n560 = ( n522  &  d ) | ( n553  &  d ) | ( n522  &  n870 ) | ( n553  &  n870 ) ;
 assign n561 = ( n192 ) | ( n788 ) ;
 assign n555 = ( n556  &  n558  &  n559  &  n560  &  n561  &  (~ n914) ) ;
 assign n562 = ( c  &  (~ n765) ) ;
 assign n564 = ( f ) | ( g ) ;
 assign n563 = ( b ) | ( n564 ) ;
 assign n566 = ( n ) | ( n241 ) ;
 assign n565 = ( j  &  n192 ) | ( n192  &  n566 ) | ( j  &  (~ n733) ) | ( n566  &  (~ n733) ) ;
 assign n568 = ( (~ n192)  &  (~ n882) ) | ( (~ j)  &  (~ n192)  &  (~ n608) ) ;
 assign n572 = ( n883  &  n782 ) | ( n883  &  n783 ) ;
 assign n573 = ( i  &  (~ n568)  &  (~ n904) ) | ( n565  &  (~ n568)  &  (~ n904) ) ;
 assign n571 = ( n572  &  n573  &  n522 ) | ( n572  &  n573  &  n290 ) ;
 assign n574 = ( c ) | ( n564 ) ;
 assign n576 = ( n775  &  n530 ) ;
 assign n575 = ( (~ j)  &  n80 ) | ( (~ j)  &  n230 ) | ( n80  &  n576 ) | ( n230  &  n576 ) ;
 assign n578 = ( n575  &  n847 ) | ( n168  &  n847 ) | ( n575  &  n154 ) | ( n168  &  n154 ) ;
 assign n579 = ( n574 ) | ( n413 ) ;
 assign n580 = ( n850  &  n612 ) | ( n718  &  n612 ) | ( n850  &  n783 ) | ( n718  &  n783 ) ;
 assign n581 = ( n849  &  n501 ) | ( n849  &  n198  &  n184 ) ;
 assign n577 = ( n578  &  n579  &  n580  &  n581 ) ;
 assign n582 = ( (~ j)  &  (~ n290)  &  (~ n413) ) | ( (~ j)  &  (~ n327)  &  (~ n413) ) ;
 assign n585 = ( c  &  b ) | ( n168  &  b ) | ( c  &  n192 ) | ( n168  &  n192 ) ;
 assign n587 = ( (~ b) ) | ( (~ e) ) | ( (~ n) ) | ( n777 ) ;
 assign n588 = ( n585 ) | ( n760 ) | ( e ) ;
 assign n589 = ( n522  &  n608 ) | ( n554  &  n608 ) | ( n522  &  n541 ) | ( n554  &  n541 ) ;
 assign n590 = ( n551 ) | ( n154 ) ;
 assign n592 = ( j ) | ( n184 ) | ( (~ n733) ) ;
 assign n586 = ( (~ n582)  &  n587  &  n588  &  n589  &  n590  &  n592 ) ;
 assign n596 = ( i ) | ( n409 ) ;
 assign n597 = ( m ) | ( n708 ) ;
 assign n595 = ( i ) | ( m ) ;
 assign n593 = ( (~ l)  &  n596  &  n597 ) | ( n596  &  n597  &  n595 ) ;
 assign n598 = ( n260  &  n99 ) ;
 assign n600 = ( n598  &  n491 ) | ( n777  &  n491 ) | ( n598  &  n511 ) | ( n777  &  n511 ) ;
 assign n599 = ( n600  &  n446 ) | ( n600  &  n137 ) ;
 assign n603 = ( (~ k) ) | ( (~ m) ) ;
 assign n601 = ( j  &  n603 ) | ( (~ m)  &  n603 ) ;
 assign n605 = ( c ) | ( (~ d) ) ;
 assign n604 = ( n54  &  g ) | ( n54  &  n605 ) ;
 assign n606 = ( (~ n162)  &  (~ n337)  &  n449 ) | ( (~ n268)  &  (~ n337)  &  n449 ) ;
 assign n609 = ( (~ e) ) | ( f ) ;
 assign n608 = ( b ) | ( n609 ) ;
 assign n610 = ( (~ d) ) | ( n721 ) ;
 assign n612 = ( j ) | ( n409 ) ;
 assign n611 = ( n72  &  n612 ) ;
 assign n615 = ( n848  &  h ) | ( n848  &  n609 ) | ( n848  &  n744 ) ;
 assign n616 = ( (~ j)  &  n605 ) | ( (~ j)  &  n608 ) | ( n605  &  n847 ) | ( n608  &  n847 ) ;
 assign n617 = ( n261  &  i ) | ( n776  &  i ) | ( n261  &  n497 ) | ( n776  &  n497 ) ;
 assign n618 = ( n742  &  n652  &  n109 ) | ( n742  &  n652  &  n760 ) ;
 assign n614 = ( n615  &  n616  &  n617  &  n618 ) ;
 assign n621 = ( (~ c)  &  (~ n609) ) ;
 assign n619 = ( (~ n169)  &  (~ n530) ) | ( (~ n169)  &  n621 ) | ( (~ n530)  &  (~ n735) ) | ( n621  &  (~ n735) ) ;
 assign n624 = ( (~ j)  &  (~ n771) ) | ( (~ j)  &  (~ n144)  &  (~ n230) ) ;
 assign n627 = ( n440  &  a ) | ( n440  &  c ) | ( n440  &  e ) ;
 assign n628 = ( e ) | ( (~ g) ) ;
 assign n629 = ( (~ n82)  &  (~ n148) ) | ( (~ n148)  &  (~ n170) ) ;
 assign n633 = ( n264 ) | ( n87 ) | ( n416 ) ;
 assign n634 = ( (~ n198)  &  (~ n563) ) | ( (~ n563)  &  (~ n774) ) ;
 assign n637 = ( (~ n576)  &  (~ n718) ) | ( (~ c)  &  (~ n718)  &  (~ n771) ) ;
 assign n640 = ( n504 ) | ( n75 ) ;
 assign n641 = ( (~ n230)  &  n629 ) | ( (~ n144)  &  (~ n230)  &  (~ n718) ) ;
 assign n644 = ( a  &  (~ n721) ) ;
 assign n642 = ( n644  &  (~ n737)  &  (~ n765) ) | ( n644  &  (~ n765)  &  (~ n784) ) ;
 assign n645 = ( (~ n522)  &  (~ n738) ) | ( (~ n79)  &  (~ n230)  &  (~ n522) ) ;
 assign n648 = ( (~ n168)  &  n619 ) | ( (~ n168)  &  n624 ) | ( (~ n168)  &  (~ n845) ) ;
 assign n651 = ( (~ e) ) | ( n554 ) ;
 assign n652 = ( l ) | ( n489 ) ;
 assign n653 = ( g ) | ( h ) | ( i ) ;
 assign n654 = ( n140 ) | ( n ) | ( n88 ) ;
 assign n655 = ( n93 ) | ( n251 ) ;
 assign n657 = ( f ) | ( n154 ) ;
 assign n656 = ( f  &  n155 ) | ( n156  &  n155 ) | ( f  &  n657 ) | ( n156  &  n657 ) ;
 assign n660 = ( (~ e) ) | ( g ) | ( n656 ) ;
 assign n659 = ( f ) | ( n249 ) ;
 assign n658 = ( (~ n47)  &  n660 ) | ( n660  &  n659 ) ;
 assign n661 = ( (~ g)  &  n  &  (~ n72) ) ;
 assign n665 = ( (~ b) ) | ( (~ d) ) ;
 assign n663 = ( n194  &  n610 ) | ( n610  &  n665 ) | ( n194  &  (~ n895) ) | ( n665  &  (~ n895) ) ;
 assign n667 = ( n301  &  n161 ) | ( n699  &  n161 ) | ( n301  &  n306 ) | ( n699  &  n306 ) ;
 assign n668 = ( n235 ) | ( n746 ) ;
 assign n669 = ( (~ e)  &  n390 ) | ( (~ e)  &  n658 ) | ( n390  &  n663 ) | ( n658  &  n663 ) ;
 assign n670 = ( n713 ) | ( n157 ) ;
 assign n671 = ( n131  &  n29  &  n379  &  n654  &  n655  &  n790 ) ;
 assign n672 = ( n221  &  n286  &  n59 ) | ( n221  &  n286  &  n732 ) ;
 assign n673 = ( n505  &  n773  &  n768  &  n506  &  n772  &  n767  &  n898  &  n897 ) ;
 assign n666 = ( n667  &  n668  &  n669  &  n670  &  n671  &  n509  &  n672  &  n673 ) ;
 assign n675 = ( f ) | ( (~ g) ) ;
 assign n674 = ( g  &  (~ n47) ) | ( (~ n47)  &  n656 ) | ( g  &  n675 ) | ( n656  &  n675 ) ;
 assign n676 = ( n700 ) | ( n390 ) ;
 assign n677 = ( n80 ) | ( n651 ) | ( n762 ) ;
 assign n678 = ( n698 ) | ( n701 ) ;
 assign n679 = ( (~ a) ) | ( n267 ) | ( n733 ) ;
 assign n680 = ( (~ d) ) | ( (~ n644) ) | ( n674 ) ;
 assign n681 = ( n900  &  n764 ) | ( n900  &  n161  &  n252 ) ;
 assign n682 = ( n301 ) | ( n701 ) ;
 assign n683 = ( n671  &  n151 ) | ( n671  &  n390 ) ;
 assign n685 = ( l ) | ( (~ n485) ) ;
 assign n686 = ( (~ h) ) | ( i ) | ( (~ l) ) ;
 assign n687 = ( l  &  n708 ) | ( (~ l)  &  n728 ) | ( n708  &  n728 ) ;
 assign n688 = ( (~ h) ) | ( n716 ) ;
 assign n689 = ( (~ l) ) | ( n398 ) ;
 assign n690 = ( (~ l) ) | ( n727 ) ;
 assign n684 = ( n685  &  n686  &  n687  &  n688  &  n689  &  n690 ) ;
 assign n692 = ( n ) | ( n93 ) ;
 assign n693 = ( (~ i) ) | ( n141 ) ;
 assign n694 = ( l ) | ( n603 ) ;
 assign n695 = ( n93 ) | ( n250 ) ;
 assign n696 = ( n ) | ( n694 ) ;
 assign n697 = ( j ) | ( n603 ) ;
 assign n698 = ( n451 ) | ( n295 ) ;
 assign n699 = ( (~ a) ) | ( n305 ) ;
 assign n700 = ( n144 ) | ( n451 ) ;
 assign n701 = ( (~ a) ) | ( (~ c) ) | ( (~ e) ) ;
 assign n702 = ( d ) | ( a ) ;
 assign n703 = ( (~ d) ) | ( e ) ;
 assign n704 = ( (~ a) ) | ( n703 ) ;
 assign n705 = ( (~ i) ) | ( j ) ;
 assign n706 = ( (~ l) ) | ( n705 ) ;
 assign n707 = ( (~ g) ) | ( (~ h) ) ;
 assign n708 = ( h ) | ( (~ i) ) ;
 assign n709 = ( (~ g) ) | ( n46 ) ;
 assign n710 = ( (~ j) ) | ( n707 ) ;
 assign n711 = ( n440  &  n441 ) ;
 assign n712 = ( n704  &  n391 ) ;
 assign n713 = ( n65  &  n390 ) ;
 assign n714 = ( g ) | ( (~ h) ) ;
 assign n715 = ( i  &  j ) ;
 assign n716 = ( (~ j) ) | ( l ) ;
 assign n717 = ( (~ f) ) | ( n605 ) ;
 assign n718 = ( l ) | ( n168 ) ;
 assign n719 = ( (~ g) ) | ( (~ n485) ) ;
 assign n721 = ( (~ b) ) | ( (~ c) ) ;
 assign n722 = ( d ) | ( n721 ) ;
 assign n723 = ( n695 ) | ( n451 ) ;
 assign n724 = ( n698 ) | ( n699 ) ;
 assign n725 = ( n41  &  n206  &  n67 ) ;
 assign n726 = ( n698  &  n700 ) | ( n214  &  n700 ) | ( n698  &  n306 ) | ( n214  &  n306 ) ;
 assign n727 = ( i ) | ( (~ j) ) ;
 assign n728 = ( j ) | ( (~ k) ) ;
 assign n730 = ( k  &  (~ n705) ) ;
 assign n731 = ( (~ k) ) | ( n256 ) ;
 assign n732 = ( (~ b) ) | ( n605 ) ;
 assign n733 = ( (~ c) ) | ( (~ d) ) ;
 assign n734 = ( i ) | ( n249 ) ;
 assign n735 = ( n719  &  n710 ) ;
 assign n736 = ( (~ g) ) | ( n727 ) ;
 assign n737 = ( k ) | ( n154 ) ;
 assign n738 = ( h ) | ( n526 ) ;
 assign n739 = ( e ) | ( n733 ) ;
 assign n740 = ( n287 ) | ( n137 ) ;
 assign n742 = ( h ) | ( n189 ) ;
 assign n743 = ( (~ b) ) | ( n526 ) ;
 assign n744 = ( (~ l) ) | ( n461 ) ;
 assign n745 = ( n717  &  n289 ) ;
 assign n746 = ( (~ f) ) | ( n665 ) ;
 assign n747 = ( i ) | ( n714 ) ;
 assign n748 = ( i ) | ( n437 ) ;
 assign n749 = ( (~ l) ) | ( n154 ) | ( n728 ) ;
 assign n750 = ( j ) | ( n707 ) ;
 assign n751 = ( j ) | ( n437 ) ;
 assign n752 = ( (~ j) ) | ( n141 ) ;
 assign n753 = ( n628 ) | ( n65 ) ;
 assign n754 = ( (~ j) ) | ( n675 ) ;
 assign n755 = ( (~ m) ) | ( n398 ) ;
 assign n758 = ( n442  &  n433 ) | ( n435  &  n433 ) | ( n442  &  n99 ) | ( n435  &  n99 ) ;
 assign n759 = ( (~ g) ) | ( n728 ) ;
 assign n760 = ( k ) | ( n705 ) ;
 assign n761 = ( b ) | ( n733 ) ;
 assign n762 = ( (~ k) ) | ( n170 ) | ( n727 ) ;
 assign n763 = ( n218  &  (~ n610) ) ;
 assign n764 = ( a ) | ( n721 ) ;
 assign n765 = ( (~ d) ) | ( (~ e) ) | ( (~ f) ) ;
 assign n767 = ( n359 ) | ( n491 ) | ( (~ n763) ) ;
 assign n768 = ( n739 ) | ( n494 ) ;
 assign n769 = ( k ) | ( n727 ) ;
 assign n770 = ( d ) | ( e ) ;
 assign n771 = ( (~ g) ) | ( h ) | ( i ) ;
 assign n772 = ( n500 ) | ( n492 ) | ( n510 ) ;
 assign n773 = ( n195 ) | ( n762 ) | ( n495 ) ;
 assign n774 = ( n58  &  n541 ) ;
 assign n775 = ( (~ g) ) | ( n554 ) ;
 assign n776 = ( a ) | ( n703 ) ;
 assign n777 = ( m ) | ( n489 ) ;
 assign n778 = ( (~ h) ) | ( n595 ) ;
 assign n779 = ( k ) | ( n595 ) ;
 assign n780 = ( h ) | ( n595 ) ;
 assign n782 = ( m ) | ( n705 ) ;
 assign n783 = ( n ) | ( n554 ) ;
 assign n784 = ( h ) | ( n154 ) ;
 assign n785 = ( g ) | ( n192 ) ;
 assign n786 = ( h  &  (~ n760) ) ;
 assign n788 = ( e ) | ( n554 ) ;
 assign n789 = ( h ) | ( n564 ) ;
 assign n790 = ( n422  &  n421  &  n723  &  n520  &  n132  &  n380 ) ;
 assign n792 = ( (~ e)  &  (~ n65) ) | ( e  &  (~ n93) ) | ( (~ n65)  &  (~ n93) ) ;
 assign n794 = ( (~ g)  &  (~ n554) ) | ( (~ g)  &  n786 ) | ( n554  &  n786 ) ;
 assign n796 = ( n903  &  i ) | ( n903  &  n533 ) | ( n903  &  h ) ;
 assign n799 = ( l ) | ( n85 ) | ( (~ n715) ) ;
 assign n798 = ( n695  &  n63 ) ;
 assign n797 = ( n799  &  n798 ) | ( n799  &  n689 ) ;
 assign n801 = ( n750  &  n260 ) ;
 assign n800 = ( n81  &  n801 ) | ( n60  &  n801 ) | ( n81  &  n82 ) | ( n60  &  n82 ) ;
 assign n802 = ( n709  &  n710 ) | ( n718  &  n710 ) | ( n709  &  n413 ) | ( n718  &  n413 ) ;
 assign n803 = ( n60  &  n719 ) | ( n264  &  n719 ) | ( n60  &  n415 ) | ( n264  &  n415 ) ;
 assign n806 = ( n51  &  (~ n123) ) | ( (~ n123)  &  n800  &  n802 ) ;
 assign n808 = ( n362  &  n354 ) ;
 assign n809 = ( n241  &  n693 ) | ( n329  &  n693 ) | ( n241  &  n80 ) | ( n329  &  n80 ) ;
 assign n810 = ( n226 ) | ( n58 ) ;
 assign n811 = ( (~ j) ) | ( n184 ) | ( n437 ) ;
 assign n813 = ( (~ a) ) | ( b ) | ( (~ d) ) | ( n188 ) ;
 assign n815 = ( n196  &  n712 ) | ( n732  &  n712 ) | ( n196  &  n151 ) | ( n732  &  n151 ) ;
 assign n816 = ( n140  &  n147 ) | ( n109  &  n147 ) | ( n140  &  n734 ) | ( n109  &  n734 ) ;
 assign n817 = ( (~ j) ) | ( n241 ) | ( n249 ) ;
 assign n818 = ( n250  &  n693 ) | ( n697  &  n693 ) | ( n250  &  n110 ) | ( n697  &  n110 ) ;
 assign n819 = ( n262 ) | ( n154 ) ;
 assign n820 = ( n239  &  n140 ) | ( n628  &  n140 ) | ( n239  &  n75 ) | ( n628  &  n75 ) ;
 assign n821 = ( n90  &  n693 ) | ( n98  &  n693 ) | ( n90  &  n77 ) | ( n98  &  n77 ) ;
 assign n823 = ( n246  &  n166 ) | ( n65  &  n166 ) | ( n246  &  n717 ) | ( n65  &  n717 ) ;
 assign n824 = ( (~ n313)  &  (~ n690) ) | ( l  &  (~ n313)  &  n715 ) ;
 assign n827 = ( (~ n69)  &  (~ n259) ) | ( (~ n69)  &  (~ n261) ) | ( (~ n69)  &  (~ n262) ) ;
 assign n831 = ( n750  &  n57 ) | ( n500  &  n57 ) | ( n750  &  n60 ) | ( n500  &  n60 ) ;
 assign n833 = ( n154  &  n264 ) | ( n264  &  (~ n824) ) | ( n154  &  (~ n827) ) | ( (~ n824)  &  (~ n827) ) ;
 assign n834 = ( n566  &  n70 ) | ( n566  &  n716 ) ;
 assign n836 = ( n154 ) | ( n79 ) | ( n389 ) | ( n398 ) ;
 assign n837 = ( (~ h) ) | ( j ) ;
 assign n838 = ( n86  &  (~ n792) ) | ( n751  &  (~ n792) ) | ( n86  &  n837 ) | ( n751  &  n837 ) ;
 assign n839 = ( j  &  n69 ) | ( n753  &  n69 ) | ( j  &  n60 ) | ( n753  &  n60 ) ;
 assign n840 = ( n86  &  n84 ) | ( n296  &  n84 ) | ( n86  &  n145 ) | ( n296  &  n145 ) ;
 assign n842 = ( n689 ) | ( n488 ) | ( n154 ) | ( n99 ) ;
 assign n843 = ( j  &  d ) | ( n501  &  d ) | ( j  &  n608 ) | ( n501  &  n608 ) ;
 assign n844 = ( n99  &  b ) | ( n498  &  b ) | ( n99  &  c ) | ( n498  &  c ) ;
 assign n845 = ( n77  &  n260 ) | ( n77  &  n530 ) | ( n260  &  (~ n545) ) | ( n530  &  (~ n545) ) ;
 assign n847 = ( n789  &  n551 ) ;
 assign n848 = ( a ) | ( b ) ;
 assign n849 = ( (~ h) ) | ( n192 ) | ( n498 ) | ( n562 ) ;
 assign n850 = ( n574  &  (~ n621) ) ;
 assign n852 = ( n776  &  n497  &  n551 ) ;
 assign n851 = ( g  &  (~ n606) ) | ( n601  &  (~ n606) ) | ( (~ n606)  &  n852 ) ;
 assign n854 = ( n851  &  n782 ) | ( n851  &  n574  &  n553 ) ;
 assign n856 = ( n152  &  n604 ) | ( n777  &  n604 ) | ( n152  &  n780 ) | ( n777  &  n780 ) ;
 assign n857 = ( n856  &  n779 ) | ( n856  &  n195  &  n775 ) ;
 assign n860 = ( n144 ) | ( n446 ) | ( n230 ) ;
 assign n861 = ( n697 ) | ( n497 ) ;
 assign n859 = ( n860  &  n861  &  n850 ) | ( n860  &  n861  &  n778 ) ;
 assign n862 = ( n599  &  n859  &  n574 ) | ( n599  &  n859  &  n593 ) ;
 assign n864 = ( n608  &  n501 ) | ( n611  &  n501 ) | ( n608  &  n778 ) | ( n611  &  n778 ) ;
 assign n865 = ( n864  &  n593 ) | ( n864  &  n501 ) ;
 assign n867 = ( n608  &  n780 ) | ( n779  &  n780 ) | ( n608  &  n441 ) | ( n779  &  n441 ) ;
 assign n871 = ( e ) | ( n539 ) | ( n610 ) ;
 assign n872 = ( (~ n702) ) | ( n744 ) | ( n784 ) ;
 assign n870 = ( (~ h)  &  n902 ) | ( n504  &  n902 ) ;
 assign n869 = ( (~ c)  &  n871  &  n872 ) | ( n871  &  n872  &  n870 ) ;
 assign n874 = ( a ) | ( (~ g) ) | ( n ) ;
 assign n875 = ( i  &  (~ n644) ) | ( i  &  n770 ) | ( (~ n644)  &  n776 ) | ( n770  &  n776 ) ;
 assign n876 = ( n337  &  (~ n536) ) | ( (~ n449)  &  (~ n536) ) | ( (~ n536)  &  n874 ) ;
 assign n878 = ( n876  &  n776 ) | ( n876  &  n784  &  n70 ) ;
 assign n880 = ( n168  &  n651 ) | ( n168  &  n785 ) | ( n651  &  (~ n794) ) | ( n785  &  (~ n794) ) ;
 assign n882 = ( n563  &  e ) | ( n563  &  n261 ) ;
 assign n883 = ( k ) | ( n198 ) | ( (~ n736) ) ;
 assign n886 = ( n627  &  (~ n642) ) | ( (~ n642)  &  n657 ) ;
 assign n888 = ( n886  &  n192 ) | ( n886  &  n844  &  n843 ) ;
 assign n892 = ( n614  &  n852 ) | ( n154  &  n852 ) | ( n614  &  n415 ) | ( n154  &  n415 ) ;
 assign n893 = ( (~ i)  &  n184 ) | ( (~ i)  &  n354 ) | ( n184  &  n577 ) | ( n354  &  n577 ) ;
 assign n894 = ( n892  &  n893  &  n696 ) | ( n892  &  n893  &  n510 ) ;
 assign n895 = ( (~ h)  &  n661 ) | ( (~ h)  &  (~ n706)  &  (~ n785) ) ;
 assign n896 = ( n241  &  n693 ) | ( n754  &  n693 ) | ( n241  &  n195 ) | ( n754  &  n195 ) ;
 assign n897 = ( n10  &  n724  &  n16 ) ;
 assign n899 = ( n76 ) | ( n94 ) | ( n610 ) ;
 assign n898 = ( n899  &  n761 ) | ( n899  &  n74  &  n187 ) ;
 assign n900 = ( n513 ) | ( n553 ) ;
 assign n902 = ( h ) | ( n168 ) | ( (~ n545) ) ;
 assign n903 = ( (~ h) ) | ( n416 ) | ( n535 ) ;
 assign n904 = ( i  &  (~ k)  &  (~ n415) ) | ( i  &  (~ k)  &  (~ n718) ) ;
 assign n905 = ( (~ h)  &  n571 ) | ( h  &  n586 ) | ( n571  &  n586 ) ;
 assign n906 = ( (~ h)  &  (~ n70) ) | ( c  &  (~ h)  &  (~ n522) ) ;
 assign n908 = ( (~ g)  &  n529 ) | ( g  &  n555 ) | ( n529  &  n555 ) ;
 assign n911 = ( l ) | ( n409 ) ;
 assign n912 = ( n596  &  n612  &  n911 ) ;
 assign n914 = ( (~ n154)  &  n527  &  n786 ) ;


endmodule

