module adder_qmap_map (sk, ax0x, bx0x, ax1x, bx1x, ax2x, bx2x, ax3x, bx3x, ax4x, bx4x, ax5x, bx5x, ax6x, bx6x, ax7x, bx7x, ax8x, bx8x, ax9x, bx9x, ax10x, bx10x, ax11x, bx11x, ax12x, bx12x, ax13x, bx13x, ax14x, bx14x, ax15x, bx15x, ax16x, bx16x, ax17x, bx17x, ax18x, bx18x, ax19x, bx19x, ax20x, bx20x, ax21x, bx21x, ax22x, bx22x, ax23x, bx23x, ax24x, bx24x, ax25x, bx25x, ax26x, bx26x, ax27x, bx27x, ax28x, bx28x, ax29x, bx29x, ax30x, bx30x, ax31x, bx31x, ax32x, bx32x, ax33x, bx33x, ax34x, bx34x, ax35x, bx35x, ax36x, bx36x, ax37x, bx37x, ax38x, bx38x, ax39x, bx39x, ax40x, bx40x, ax41x, bx41x, ax42x, bx42x, ax43x, bx43x, ax44x, bx44x, ax45x, bx45x, ax46x, bx46x, ax47x, bx47x, ax48x, bx48x, ax49x, bx49x, ax50x, bx50x, ax51x, bx51x, ax52x, bx52x, ax53x, bx53x, ax54x, bx54x, ax55x, bx55x, ax56x, bx56x, ax57x, bx57x, ax58x, bx58x, ax59x, bx59x, ax60x, bx60x, ax61x, bx61x, ax62x, bx62x, ax63x, bx63x, ax64x, bx64x, ax65x, bx65x, ax66x, bx66x, ax67x, bx67x, ax68x, bx68x, ax69x, bx69x, ax70x, bx70x, ax71x, bx71x, ax72x, bx72x, ax73x, bx73x, ax74x, bx74x, ax75x, bx75x, ax76x, bx76x, ax77x, bx77x, ax78x, bx78x, ax79x, bx79x, ax80x, bx80x, ax81x, bx81x, ax82x, bx82x, ax83x, bx83x, ax84x, bx84x, ax85x, bx85x, ax86x, bx86x, ax87x, bx87x, ax88x, bx88x, ax89x, bx89x, ax90x, bx90x, ax91x, bx91x, ax92x, bx92x, ax93x, bx93x, ax94x, bx94x, ax95x, bx95x, ax96x, bx96x, ax97x, bx97x, ax98x, bx98x, ax99x, bx99x, ax100x, bx100x, ax101x, bx101x, ax102x, bx102x, ax103x, bx103x, ax104x, bx104x, ax105x, bx105x, ax106x, bx106x, ax107x, bx107x, ax108x, bx108x, ax109x, bx109x, ax110x, bx110x, ax111x, bx111x, ax112x, bx112x, ax113x, bx113x, ax114x, bx114x, ax115x, bx115x, ax116x, bx116x, ax117x, bx117x, ax118x, bx118x, ax119x, bx119x, ax120x, bx120x, ax121x, bx121x, ax122x, bx122x, ax123x, bx123x, ax124x, bx124x, ax125x, bx125x, ax126x, bx126x, ax127x, bx127x, fx0x, fx1x, fx2x, fx3x, fx4x, fx5x, fx6x, fx7x, fx8x, fx9x, fx10x, fx11x, fx12x, fx13x, fx14x, fx15x, fx16x, fx17x, fx18x, fx19x, fx20x, fx21x, fx22x, fx23x, fx24x, fx25x, fx26x, fx27x, fx28x, fx29x, fx30x, fx31x, fx32x, fx33x, fx34x, fx35x, fx36x, fx37x, fx38x, fx39x, fx40x, fx41x, fx42x, fx43x, fx44x, fx45x, fx46x, fx47x, fx48x, fx49x, fx50x, fx51x, fx52x, fx53x, fx54x, fx55x, fx56x, fx57x, fx58x, fx59x, fx60x, fx61x, fx62x, fx63x, fx64x, fx65x, fx66x, fx67x, fx68x, fx69x, fx70x, fx71x, fx72x, fx73x, fx74x, fx75x, fx76x, fx77x, fx78x, fx79x, fx80x, fx81x, fx82x, fx83x, fx84x, fx85x, fx86x, fx87x, fx88x, fx89x, fx90x, fx91x, fx92x, fx93x, fx94x, fx95x, fx96x, fx97x, fx98x, fx99x, fx100x, fx101x, fx102x, fx103x, fx104x, fx105x, fx106x, fx107x, fx108x, fx109x, fx110x, fx111x, fx112x, fx113x, fx114x, fx115x, fx116x, fx117x, fx118x, fx119x, fx120x, fx121x, fx122x, fx123x, fx124x, fx125x, fx126x, fx127x, cOut);

	input ax0x;
	input bx0x;
	input ax1x;
	input bx1x;
	input ax2x;
	input bx2x;
	input ax3x;
	input bx3x;
	input ax4x;
	input bx4x;
	input ax5x;
	input bx5x;
	input ax6x;
	input bx6x;
	input ax7x;
	input bx7x;
	input ax8x;
	input bx8x;
	input ax9x;
	input bx9x;
	input ax10x;
	input bx10x;
	input ax11x;
	input bx11x;
	input ax12x;
	input bx12x;
	input ax13x;
	input bx13x;
	input ax14x;
	input bx14x;
	input ax15x;
	input bx15x;
	input ax16x;
	input bx16x;
	input ax17x;
	input bx17x;
	input ax18x;
	input bx18x;
	input ax19x;
	input bx19x;
	input ax20x;
	input bx20x;
	input ax21x;
	input bx21x;
	input ax22x;
	input bx22x;
	input ax23x;
	input bx23x;
	input ax24x;
	input bx24x;
	input ax25x;
	input bx25x;
	input ax26x;
	input bx26x;
	input ax27x;
	input bx27x;
	input ax28x;
	input bx28x;
	input ax29x;
	input bx29x;
	input ax30x;
	input bx30x;
	input ax31x;
	input bx31x;
	input ax32x;
	input bx32x;
	input ax33x;
	input bx33x;
	input ax34x;
	input bx34x;
	input ax35x;
	input bx35x;
	input ax36x;
	input bx36x;
	input ax37x;
	input bx37x;
	input ax38x;
	input bx38x;
	input ax39x;
	input bx39x;
	input ax40x;
	input bx40x;
	input ax41x;
	input bx41x;
	input ax42x;
	input bx42x;
	input ax43x;
	input bx43x;
	input ax44x;
	input bx44x;
	input ax45x;
	input bx45x;
	input ax46x;
	input bx46x;
	input ax47x;
	input bx47x;
	input ax48x;
	input bx48x;
	input ax49x;
	input bx49x;
	input ax50x;
	input bx50x;
	input ax51x;
	input bx51x;
	input ax52x;
	input bx52x;
	input ax53x;
	input bx53x;
	input ax54x;
	input bx54x;
	input ax55x;
	input bx55x;
	input ax56x;
	input bx56x;
	input ax57x;
	input bx57x;
	input ax58x;
	input bx58x;
	input ax59x;
	input bx59x;
	input ax60x;
	input bx60x;
	input ax61x;
	input bx61x;
	input ax62x;
	input bx62x;
	input ax63x;
	input bx63x;
	input ax64x;
	input bx64x;
	input ax65x;
	input bx65x;
	input ax66x;
	input bx66x;
	input ax67x;
	input bx67x;
	input ax68x;
	input bx68x;
	input ax69x;
	input bx69x;
	input ax70x;
	input bx70x;
	input ax71x;
	input bx71x;
	input ax72x;
	input bx72x;
	input ax73x;
	input bx73x;
	input ax74x;
	input bx74x;
	input ax75x;
	input bx75x;
	input ax76x;
	input bx76x;
	input ax77x;
	input bx77x;
	input ax78x;
	input bx78x;
	input ax79x;
	input bx79x;
	input ax80x;
	input bx80x;
	input ax81x;
	input bx81x;
	input ax82x;
	input bx82x;
	input ax83x;
	input bx83x;
	input ax84x;
	input bx84x;
	input ax85x;
	input bx85x;
	input ax86x;
	input bx86x;
	input ax87x;
	input bx87x;
	input ax88x;
	input bx88x;
	input ax89x;
	input bx89x;
	input ax90x;
	input bx90x;
	input ax91x;
	input bx91x;
	input ax92x;
	input bx92x;
	input ax93x;
	input bx93x;
	input ax94x;
	input bx94x;
	input ax95x;
	input bx95x;
	input ax96x;
	input bx96x;
	input ax97x;
	input bx97x;
	input ax98x;
	input bx98x;
	input ax99x;
	input bx99x;
	input ax100x;
	input bx100x;
	input ax101x;
	input bx101x;
	input ax102x;
	input bx102x;
	input ax103x;
	input bx103x;
	input ax104x;
	input bx104x;
	input ax105x;
	input bx105x;
	input ax106x;
	input bx106x;
	input ax107x;
	input bx107x;
	input ax108x;
	input bx108x;
	input ax109x;
	input bx109x;
	input ax110x;
	input bx110x;
	input ax111x;
	input bx111x;
	input ax112x;
	input bx112x;
	input ax113x;
	input bx113x;
	input ax114x;
	input bx114x;
	input ax115x;
	input bx115x;
	input ax116x;
	input bx116x;
	input ax117x;
	input bx117x;
	input ax118x;
	input bx118x;
	input ax119x;
	input bx119x;
	input ax120x;
	input bx120x;
	input ax121x;
	input bx121x;
	input ax122x;
	input bx122x;
	input ax123x;
	input bx123x;
	input ax124x;
	input bx124x;
	input ax125x;
	input bx125x;
	input ax126x;
	input bx126x;
	input ax127x;
	input bx127x;
	output fx0x;
	output fx1x;
	output fx2x;
	output fx3x;
	output fx4x;
	output fx5x;
	output fx6x;
	output fx7x;
	output fx8x;
	output fx9x;
	output fx10x;
	output fx11x;
	output fx12x;
	output fx13x;
	output fx14x;
	output fx15x;
	output fx16x;
	output fx17x;
	output fx18x;
	output fx19x;
	output fx20x;
	output fx21x;
	output fx22x;
	output fx23x;
	output fx24x;
	output fx25x;
	output fx26x;
	output fx27x;
	output fx28x;
	output fx29x;
	output fx30x;
	output fx31x;
	output fx32x;
	output fx33x;
	output fx34x;
	output fx35x;
	output fx36x;
	output fx37x;
	output fx38x;
	output fx39x;
	output fx40x;
	output fx41x;
	output fx42x;
	output fx43x;
	output fx44x;
	output fx45x;
	output fx46x;
	output fx47x;
	output fx48x;
	output fx49x;
	output fx50x;
	output fx51x;
	output fx52x;
	output fx53x;
	output fx54x;
	output fx55x;
	output fx56x;
	output fx57x;
	output fx58x;
	output fx59x;
	output fx60x;
	output fx61x;
	output fx62x;
	output fx63x;
	output fx64x;
	output fx65x;
	output fx66x;
	output fx67x;
	output fx68x;
	output fx69x;
	output fx70x;
	output fx71x;
	output fx72x;
	output fx73x;
	output fx74x;
	output fx75x;
	output fx76x;
	output fx77x;
	output fx78x;
	output fx79x;
	output fx80x;
	output fx81x;
	output fx82x;
	output fx83x;
	output fx84x;
	output fx85x;
	output fx86x;
	output fx87x;
	output fx88x;
	output fx89x;
	output fx90x;
	output fx91x;
	output fx92x;
	output fx93x;
	output fx94x;
	output fx95x;
	output fx96x;
	output fx97x;
	output fx98x;
	output fx99x;
	output fx100x;
	output fx101x;
	output fx102x;
	output fx103x;
	output fx104x;
	output fx105x;
	output fx106x;
	output fx107x;
	output fx108x;
	output fx109x;
	output fx110x;
	output fx111x;
	output fx112x;
	output fx113x;
	output fx114x;
	output fx115x;
	output fx116x;
	output fx117x;
	output fx118x;
	output fx119x;
	output fx120x;
	output fx121x;
	output fx122x;
	output fx123x;
	output fx124x;
	output fx125x;
	output fx126x;
	output fx127x;
	output cOut;



	wire g4, g6, g9, g10, g11, g12, g15, g17, g20, g21, g22, g23, g26, g28, g31, g32, g33, g34, g37, g39, g42;
	wire g43, g44, g45, g48, g50, g53, g54, g55, g56, g59, g61, g64, g65, g66, g67, g70, g72, g75, g76, g77, g78;
	wire g81, g83, g86, g87, g88, g89, g92, g94, g97, g98, g99, g100, g103, g105, g108, g109, g110, g113, g115, g118, g119;
	wire g120, g121, g124, g126, g129, g130, g131, g132, g135, g137, g140, g141, g142, g143, g146, g148, g151, g152, g153, g154, g157;
	wire g159, g162, g163, g164, g165, g168, g170, g173, g174, g175, g178, g180, g183, g184, g185, g186, g189, g191, g194, g195, g196;
	wire g199, g201, g204, g205, g206, g207, g210, g212, g215, g216, g217, g218, g221, g223, g226, g227, g228, g231, g234, g236, g237;
	wire g238, g241, g244, g246, g247, g248, g251, g254, g256, g257, g258, g261, g264, g266, g267, g268;

	assign fx0x = (((!ax0x) & (bx0x)) + ((ax0x) & (!bx0x)));
	assign fx1x = (((!ax0x) & (!bx0x) & (!ax1x) & (bx1x)) + ((!ax0x) & (!bx0x) & (ax1x) & (!bx1x)) + ((!ax0x) & (bx0x) & (!ax1x) & (bx1x)) + ((!ax0x) & (bx0x) & (ax1x) & (!bx1x)) + ((ax0x) & (!bx0x) & (!ax1x) & (bx1x)) + ((ax0x) & (!bx0x) & (ax1x) & (!bx1x)) + ((ax0x) & (bx0x) & (!ax1x) & (!bx1x)) + ((ax0x) & (bx0x) & (ax1x) & (bx1x)));
	assign fx2x = (((!ax0x) & (!bx0x) & (!ax1x) & (!bx1x) & (!ax2x) & (bx2x)) + ((!ax0x) & (!bx0x) & (!ax1x) & (!bx1x) & (ax2x) & (!bx2x)) + ((!ax0x) & (!bx0x) & (!ax1x) & (bx1x) & (!ax2x) & (bx2x)) + ((!ax0x) & (!bx0x) & (!ax1x) & (bx1x) & (ax2x) & (!bx2x)) + ((!ax0x) & (!bx0x) & (ax1x) & (!bx1x) & (!ax2x) & (bx2x)) + ((!ax0x) & (!bx0x) & (ax1x) & (!bx1x) & (ax2x) & (!bx2x)) + ((!ax0x) & (!bx0x) & (ax1x) & (bx1x) & (!ax2x) & (!bx2x)) + ((!ax0x) & (!bx0x) & (ax1x) & (bx1x) & (ax2x) & (bx2x)) + ((!ax0x) & (bx0x) & (!ax1x) & (!bx1x) & (!ax2x) & (bx2x)) + ((!ax0x) & (bx0x) & (!ax1x) & (!bx1x) & (ax2x) & (!bx2x)) + ((!ax0x) & (bx0x) & (!ax1x) & (bx1x) & (!ax2x) & (bx2x)) + ((!ax0x) & (bx0x) & (!ax1x) & (bx1x) & (ax2x) & (!bx2x)) + ((!ax0x) & (bx0x) & (ax1x) & (!bx1x) & (!ax2x) & (bx2x)) + ((!ax0x) & (bx0x) & (ax1x) & (!bx1x) & (ax2x) & (!bx2x)) + ((!ax0x) & (bx0x) & (ax1x) & (bx1x) & (!ax2x) & (!bx2x)) + ((!ax0x) & (bx0x) & (ax1x) & (bx1x) & (ax2x) & (bx2x)) + ((ax0x) & (!bx0x) & (!ax1x) & (!bx1x) & (!ax2x) & (bx2x)) + ((ax0x) & (!bx0x) & (!ax1x) & (!bx1x) & (ax2x) & (!bx2x)) + ((ax0x) & (!bx0x) & (!ax1x) & (bx1x) & (!ax2x) & (bx2x)) + ((ax0x) & (!bx0x) & (!ax1x) & (bx1x) & (ax2x) & (!bx2x)) + ((ax0x) & (!bx0x) & (ax1x) & (!bx1x) & (!ax2x) & (bx2x)) + ((ax0x) & (!bx0x) & (ax1x) & (!bx1x) & (ax2x) & (!bx2x)) + ((ax0x) & (!bx0x) & (ax1x) & (bx1x) & (!ax2x) & (!bx2x)) + ((ax0x) & (!bx0x) & (ax1x) & (bx1x) & (ax2x) & (bx2x)) + ((ax0x) & (bx0x) & (!ax1x) & (!bx1x) & (!ax2x) & (bx2x)) + ((ax0x) & (bx0x) & (!ax1x) & (!bx1x) & (ax2x) & (!bx2x)) + ((ax0x) & (bx0x) & (!ax1x) & (bx1x) & (!ax2x) & (!bx2x)) + ((ax0x) & (bx0x) & (!ax1x) & (bx1x) & (ax2x) & (bx2x)) + ((ax0x) & (bx0x) & (ax1x) & (!bx1x) & (!ax2x) & (!bx2x)) + ((ax0x) & (bx0x) & (ax1x) & (!bx1x) & (ax2x) & (bx2x)) + ((ax0x) & (bx0x) & (ax1x) & (bx1x) & (!ax2x) & (!bx2x)) + ((ax0x) & (bx0x) & (ax1x) & (bx1x) & (ax2x) & (bx2x)));
	assign g4 = (((!ax0x) & (!bx0x) & (!ax1x) & (!bx1x) & (ax2x) & (bx2x)) + ((!ax0x) & (!bx0x) & (!ax1x) & (bx1x) & (ax2x) & (bx2x)) + ((!ax0x) & (!bx0x) & (ax1x) & (!bx1x) & (ax2x) & (bx2x)) + ((!ax0x) & (!bx0x) & (ax1x) & (bx1x) & (!ax2x) & (bx2x)) + ((!ax0x) & (!bx0x) & (ax1x) & (bx1x) & (ax2x) & (!bx2x)) + ((!ax0x) & (!bx0x) & (ax1x) & (bx1x) & (ax2x) & (bx2x)) + ((!ax0x) & (bx0x) & (!ax1x) & (!bx1x) & (ax2x) & (bx2x)) + ((!ax0x) & (bx0x) & (!ax1x) & (bx1x) & (ax2x) & (bx2x)) + ((!ax0x) & (bx0x) & (ax1x) & (!bx1x) & (ax2x) & (bx2x)) + ((!ax0x) & (bx0x) & (ax1x) & (bx1x) & (!ax2x) & (bx2x)) + ((!ax0x) & (bx0x) & (ax1x) & (bx1x) & (ax2x) & (!bx2x)) + ((!ax0x) & (bx0x) & (ax1x) & (bx1x) & (ax2x) & (bx2x)) + ((ax0x) & (!bx0x) & (!ax1x) & (!bx1x) & (ax2x) & (bx2x)) + ((ax0x) & (!bx0x) & (!ax1x) & (bx1x) & (ax2x) & (bx2x)) + ((ax0x) & (!bx0x) & (ax1x) & (!bx1x) & (ax2x) & (bx2x)) + ((ax0x) & (!bx0x) & (ax1x) & (bx1x) & (!ax2x) & (bx2x)) + ((ax0x) & (!bx0x) & (ax1x) & (bx1x) & (ax2x) & (!bx2x)) + ((ax0x) & (!bx0x) & (ax1x) & (bx1x) & (ax2x) & (bx2x)) + ((ax0x) & (bx0x) & (!ax1x) & (!bx1x) & (ax2x) & (bx2x)) + ((ax0x) & (bx0x) & (!ax1x) & (bx1x) & (!ax2x) & (bx2x)) + ((ax0x) & (bx0x) & (!ax1x) & (bx1x) & (ax2x) & (!bx2x)) + ((ax0x) & (bx0x) & (!ax1x) & (bx1x) & (ax2x) & (bx2x)) + ((ax0x) & (bx0x) & (ax1x) & (!bx1x) & (!ax2x) & (bx2x)) + ((ax0x) & (bx0x) & (ax1x) & (!bx1x) & (ax2x) & (!bx2x)) + ((ax0x) & (bx0x) & (ax1x) & (!bx1x) & (ax2x) & (bx2x)) + ((ax0x) & (bx0x) & (ax1x) & (bx1x) & (!ax2x) & (bx2x)) + ((ax0x) & (bx0x) & (ax1x) & (bx1x) & (ax2x) & (!bx2x)) + ((ax0x) & (bx0x) & (ax1x) & (bx1x) & (ax2x) & (bx2x)));
	assign fx3x = (((!ax3x) & (!bx3x) & (g4)) + ((!ax3x) & (bx3x) & (!g4)) + ((ax3x) & (!bx3x) & (!g4)) + ((ax3x) & (bx3x) & (g4)));
	assign g6 = (((!ax3x) & (bx3x) & (g4)) + ((ax3x) & (!bx3x) & (g4)) + ((ax3x) & (bx3x) & (!g4)) + ((ax3x) & (bx3x) & (g4)));
	assign fx4x = (((!ax4x) & (!bx4x) & (g6)) + ((!ax4x) & (bx4x) & (!g6)) + ((ax4x) & (!bx4x) & (!g6)) + ((ax4x) & (bx4x) & (g6)));
	assign fx5x = (((!ax4x) & (!bx4x) & (!g6) & (!ax5x) & (bx5x)) + ((!ax4x) & (!bx4x) & (!g6) & (ax5x) & (!bx5x)) + ((!ax4x) & (!bx4x) & (g6) & (!ax5x) & (bx5x)) + ((!ax4x) & (!bx4x) & (g6) & (ax5x) & (!bx5x)) + ((!ax4x) & (bx4x) & (!g6) & (!ax5x) & (bx5x)) + ((!ax4x) & (bx4x) & (!g6) & (ax5x) & (!bx5x)) + ((!ax4x) & (bx4x) & (g6) & (!ax5x) & (!bx5x)) + ((!ax4x) & (bx4x) & (g6) & (ax5x) & (bx5x)) + ((ax4x) & (!bx4x) & (!g6) & (!ax5x) & (bx5x)) + ((ax4x) & (!bx4x) & (!g6) & (ax5x) & (!bx5x)) + ((ax4x) & (!bx4x) & (g6) & (!ax5x) & (!bx5x)) + ((ax4x) & (!bx4x) & (g6) & (ax5x) & (bx5x)) + ((ax4x) & (bx4x) & (!g6) & (!ax5x) & (!bx5x)) + ((ax4x) & (bx4x) & (!g6) & (ax5x) & (bx5x)) + ((ax4x) & (bx4x) & (g6) & (!ax5x) & (!bx5x)) + ((ax4x) & (bx4x) & (g6) & (ax5x) & (bx5x)));
	assign g9 = (((ax5x) & (bx5x)));
	assign g10 = (((!ax5x) & (!bx5x)));
	assign g11 = (((!ax3x) & (!bx3x) & (!g4) & (ax4x) & (bx4x) & (!g10)) + ((!ax3x) & (!bx3x) & (g4) & (ax4x) & (bx4x) & (!g10)) + ((!ax3x) & (bx3x) & (!g4) & (ax4x) & (bx4x) & (!g10)) + ((!ax3x) & (bx3x) & (g4) & (!ax4x) & (bx4x) & (!g10)) + ((!ax3x) & (bx3x) & (g4) & (ax4x) & (!bx4x) & (!g10)) + ((!ax3x) & (bx3x) & (g4) & (ax4x) & (bx4x) & (!g10)) + ((ax3x) & (!bx3x) & (!g4) & (ax4x) & (bx4x) & (!g10)) + ((ax3x) & (!bx3x) & (g4) & (!ax4x) & (bx4x) & (!g10)) + ((ax3x) & (!bx3x) & (g4) & (ax4x) & (!bx4x) & (!g10)) + ((ax3x) & (!bx3x) & (g4) & (ax4x) & (bx4x) & (!g10)) + ((ax3x) & (bx3x) & (!g4) & (!ax4x) & (bx4x) & (!g10)) + ((ax3x) & (bx3x) & (!g4) & (ax4x) & (!bx4x) & (!g10)) + ((ax3x) & (bx3x) & (!g4) & (ax4x) & (bx4x) & (!g10)) + ((ax3x) & (bx3x) & (g4) & (!ax4x) & (bx4x) & (!g10)) + ((ax3x) & (bx3x) & (g4) & (ax4x) & (!bx4x) & (!g10)) + ((ax3x) & (bx3x) & (g4) & (ax4x) & (bx4x) & (!g10)));
	assign g12 = (((!g9) & (!g11)));
	assign fx6x = (((!ax6x) & (!bx6x) & (!g12)) + ((!ax6x) & (bx6x) & (g12)) + ((ax6x) & (!bx6x) & (g12)) + ((ax6x) & (bx6x) & (!g12)));
	assign fx7x = (((!ax6x) & (!bx6x) & (!g12) & (!ax7x) & (bx7x)) + ((!ax6x) & (!bx6x) & (!g12) & (ax7x) & (!bx7x)) + ((!ax6x) & (!bx6x) & (g12) & (!ax7x) & (bx7x)) + ((!ax6x) & (!bx6x) & (g12) & (ax7x) & (!bx7x)) + ((!ax6x) & (bx6x) & (!g12) & (!ax7x) & (!bx7x)) + ((!ax6x) & (bx6x) & (!g12) & (ax7x) & (bx7x)) + ((!ax6x) & (bx6x) & (g12) & (!ax7x) & (bx7x)) + ((!ax6x) & (bx6x) & (g12) & (ax7x) & (!bx7x)) + ((ax6x) & (!bx6x) & (!g12) & (!ax7x) & (!bx7x)) + ((ax6x) & (!bx6x) & (!g12) & (ax7x) & (bx7x)) + ((ax6x) & (!bx6x) & (g12) & (!ax7x) & (bx7x)) + ((ax6x) & (!bx6x) & (g12) & (ax7x) & (!bx7x)) + ((ax6x) & (bx6x) & (!g12) & (!ax7x) & (!bx7x)) + ((ax6x) & (bx6x) & (!g12) & (ax7x) & (bx7x)) + ((ax6x) & (bx6x) & (g12) & (!ax7x) & (!bx7x)) + ((ax6x) & (bx6x) & (g12) & (ax7x) & (bx7x)));
	assign g15 = (((!ax6x) & (!bx6x) & (!g9) & (!g11) & (!ax7x) & (!bx7x)) + ((!ax6x) & (!bx6x) & (!g9) & (!g11) & (!ax7x) & (bx7x)) + ((!ax6x) & (!bx6x) & (!g9) & (!g11) & (ax7x) & (!bx7x)) + ((!ax6x) & (!bx6x) & (!g9) & (g11) & (!ax7x) & (!bx7x)) + ((!ax6x) & (!bx6x) & (!g9) & (g11) & (!ax7x) & (bx7x)) + ((!ax6x) & (!bx6x) & (!g9) & (g11) & (ax7x) & (!bx7x)) + ((!ax6x) & (!bx6x) & (g9) & (!g11) & (!ax7x) & (!bx7x)) + ((!ax6x) & (!bx6x) & (g9) & (!g11) & (!ax7x) & (bx7x)) + ((!ax6x) & (!bx6x) & (g9) & (!g11) & (ax7x) & (!bx7x)) + ((!ax6x) & (!bx6x) & (g9) & (g11) & (!ax7x) & (!bx7x)) + ((!ax6x) & (!bx6x) & (g9) & (g11) & (!ax7x) & (bx7x)) + ((!ax6x) & (!bx6x) & (g9) & (g11) & (ax7x) & (!bx7x)) + ((!ax6x) & (bx6x) & (!g9) & (!g11) & (!ax7x) & (!bx7x)) + ((!ax6x) & (bx6x) & (!g9) & (!g11) & (!ax7x) & (bx7x)) + ((!ax6x) & (bx6x) & (!g9) & (!g11) & (ax7x) & (!bx7x)) + ((!ax6x) & (bx6x) & (!g9) & (g11) & (!ax7x) & (!bx7x)) + ((!ax6x) & (bx6x) & (g9) & (!g11) & (!ax7x) & (!bx7x)) + ((!ax6x) & (bx6x) & (g9) & (g11) & (!ax7x) & (!bx7x)) + ((ax6x) & (!bx6x) & (!g9) & (!g11) & (!ax7x) & (!bx7x)) + ((ax6x) & (!bx6x) & (!g9) & (!g11) & (!ax7x) & (bx7x)) + ((ax6x) & (!bx6x) & (!g9) & (!g11) & (ax7x) & (!bx7x)) + ((ax6x) & (!bx6x) & (!g9) & (g11) & (!ax7x) & (!bx7x)) + ((ax6x) & (!bx6x) & (g9) & (!g11) & (!ax7x) & (!bx7x)) + ((ax6x) & (!bx6x) & (g9) & (g11) & (!ax7x) & (!bx7x)) + ((ax6x) & (bx6x) & (!g9) & (!g11) & (!ax7x) & (!bx7x)) + ((ax6x) & (bx6x) & (!g9) & (g11) & (!ax7x) & (!bx7x)) + ((ax6x) & (bx6x) & (g9) & (!g11) & (!ax7x) & (!bx7x)) + ((ax6x) & (bx6x) & (g9) & (g11) & (!ax7x) & (!bx7x)));
	assign fx8x = (((!ax8x) & (!bx8x) & (!g15)) + ((!ax8x) & (bx8x) & (g15)) + ((ax8x) & (!bx8x) & (g15)) + ((ax8x) & (bx8x) & (!g15)));
	assign g17 = (((!ax8x) & (bx8x) & (!g15)) + ((ax8x) & (!bx8x) & (!g15)) + ((ax8x) & (bx8x) & (!g15)) + ((ax8x) & (bx8x) & (g15)));
	assign fx9x = (((!ax9x) & (!bx9x) & (g17)) + ((!ax9x) & (bx9x) & (!g17)) + ((ax9x) & (!bx9x) & (!g17)) + ((ax9x) & (bx9x) & (g17)));
	assign fx10x = (((!ax9x) & (!bx9x) & (!g17) & (!ax10x) & (bx10x)) + ((!ax9x) & (!bx9x) & (!g17) & (ax10x) & (!bx10x)) + ((!ax9x) & (!bx9x) & (g17) & (!ax10x) & (bx10x)) + ((!ax9x) & (!bx9x) & (g17) & (ax10x) & (!bx10x)) + ((!ax9x) & (bx9x) & (!g17) & (!ax10x) & (bx10x)) + ((!ax9x) & (bx9x) & (!g17) & (ax10x) & (!bx10x)) + ((!ax9x) & (bx9x) & (g17) & (!ax10x) & (!bx10x)) + ((!ax9x) & (bx9x) & (g17) & (ax10x) & (bx10x)) + ((ax9x) & (!bx9x) & (!g17) & (!ax10x) & (bx10x)) + ((ax9x) & (!bx9x) & (!g17) & (ax10x) & (!bx10x)) + ((ax9x) & (!bx9x) & (g17) & (!ax10x) & (!bx10x)) + ((ax9x) & (!bx9x) & (g17) & (ax10x) & (bx10x)) + ((ax9x) & (bx9x) & (!g17) & (!ax10x) & (!bx10x)) + ((ax9x) & (bx9x) & (!g17) & (ax10x) & (bx10x)) + ((ax9x) & (bx9x) & (g17) & (!ax10x) & (!bx10x)) + ((ax9x) & (bx9x) & (g17) & (ax10x) & (bx10x)));
	assign g20 = (((ax10x) & (bx10x)));
	assign g21 = (((!ax10x) & (!bx10x)));
	assign g22 = (((!ax8x) & (!bx8x) & (!g15) & (ax9x) & (bx9x) & (!g21)) + ((!ax8x) & (!bx8x) & (g15) & (ax9x) & (bx9x) & (!g21)) + ((!ax8x) & (bx8x) & (!g15) & (!ax9x) & (bx9x) & (!g21)) + ((!ax8x) & (bx8x) & (!g15) & (ax9x) & (!bx9x) & (!g21)) + ((!ax8x) & (bx8x) & (!g15) & (ax9x) & (bx9x) & (!g21)) + ((!ax8x) & (bx8x) & (g15) & (ax9x) & (bx9x) & (!g21)) + ((ax8x) & (!bx8x) & (!g15) & (!ax9x) & (bx9x) & (!g21)) + ((ax8x) & (!bx8x) & (!g15) & (ax9x) & (!bx9x) & (!g21)) + ((ax8x) & (!bx8x) & (!g15) & (ax9x) & (bx9x) & (!g21)) + ((ax8x) & (!bx8x) & (g15) & (ax9x) & (bx9x) & (!g21)) + ((ax8x) & (bx8x) & (!g15) & (!ax9x) & (bx9x) & (!g21)) + ((ax8x) & (bx8x) & (!g15) & (ax9x) & (!bx9x) & (!g21)) + ((ax8x) & (bx8x) & (!g15) & (ax9x) & (bx9x) & (!g21)) + ((ax8x) & (bx8x) & (g15) & (!ax9x) & (bx9x) & (!g21)) + ((ax8x) & (bx8x) & (g15) & (ax9x) & (!bx9x) & (!g21)) + ((ax8x) & (bx8x) & (g15) & (ax9x) & (bx9x) & (!g21)));
	assign g23 = (((!g20) & (!g22)));
	assign fx11x = (((!ax11x) & (!bx11x) & (!g23)) + ((!ax11x) & (bx11x) & (g23)) + ((ax11x) & (!bx11x) & (g23)) + ((ax11x) & (bx11x) & (!g23)));
	assign fx12x = (((!ax11x) & (!bx11x) & (!g23) & (!ax12x) & (bx12x)) + ((!ax11x) & (!bx11x) & (!g23) & (ax12x) & (!bx12x)) + ((!ax11x) & (!bx11x) & (g23) & (!ax12x) & (bx12x)) + ((!ax11x) & (!bx11x) & (g23) & (ax12x) & (!bx12x)) + ((!ax11x) & (bx11x) & (!g23) & (!ax12x) & (!bx12x)) + ((!ax11x) & (bx11x) & (!g23) & (ax12x) & (bx12x)) + ((!ax11x) & (bx11x) & (g23) & (!ax12x) & (bx12x)) + ((!ax11x) & (bx11x) & (g23) & (ax12x) & (!bx12x)) + ((ax11x) & (!bx11x) & (!g23) & (!ax12x) & (!bx12x)) + ((ax11x) & (!bx11x) & (!g23) & (ax12x) & (bx12x)) + ((ax11x) & (!bx11x) & (g23) & (!ax12x) & (bx12x)) + ((ax11x) & (!bx11x) & (g23) & (ax12x) & (!bx12x)) + ((ax11x) & (bx11x) & (!g23) & (!ax12x) & (!bx12x)) + ((ax11x) & (bx11x) & (!g23) & (ax12x) & (bx12x)) + ((ax11x) & (bx11x) & (g23) & (!ax12x) & (!bx12x)) + ((ax11x) & (bx11x) & (g23) & (ax12x) & (bx12x)));
	assign g26 = (((!ax11x) & (!bx11x) & (!g20) & (!g22) & (!ax12x) & (!bx12x)) + ((!ax11x) & (!bx11x) & (!g20) & (!g22) & (!ax12x) & (bx12x)) + ((!ax11x) & (!bx11x) & (!g20) & (!g22) & (ax12x) & (!bx12x)) + ((!ax11x) & (!bx11x) & (!g20) & (g22) & (!ax12x) & (!bx12x)) + ((!ax11x) & (!bx11x) & (!g20) & (g22) & (!ax12x) & (bx12x)) + ((!ax11x) & (!bx11x) & (!g20) & (g22) & (ax12x) & (!bx12x)) + ((!ax11x) & (!bx11x) & (g20) & (!g22) & (!ax12x) & (!bx12x)) + ((!ax11x) & (!bx11x) & (g20) & (!g22) & (!ax12x) & (bx12x)) + ((!ax11x) & (!bx11x) & (g20) & (!g22) & (ax12x) & (!bx12x)) + ((!ax11x) & (!bx11x) & (g20) & (g22) & (!ax12x) & (!bx12x)) + ((!ax11x) & (!bx11x) & (g20) & (g22) & (!ax12x) & (bx12x)) + ((!ax11x) & (!bx11x) & (g20) & (g22) & (ax12x) & (!bx12x)) + ((!ax11x) & (bx11x) & (!g20) & (!g22) & (!ax12x) & (!bx12x)) + ((!ax11x) & (bx11x) & (!g20) & (!g22) & (!ax12x) & (bx12x)) + ((!ax11x) & (bx11x) & (!g20) & (!g22) & (ax12x) & (!bx12x)) + ((!ax11x) & (bx11x) & (!g20) & (g22) & (!ax12x) & (!bx12x)) + ((!ax11x) & (bx11x) & (g20) & (!g22) & (!ax12x) & (!bx12x)) + ((!ax11x) & (bx11x) & (g20) & (g22) & (!ax12x) & (!bx12x)) + ((ax11x) & (!bx11x) & (!g20) & (!g22) & (!ax12x) & (!bx12x)) + ((ax11x) & (!bx11x) & (!g20) & (!g22) & (!ax12x) & (bx12x)) + ((ax11x) & (!bx11x) & (!g20) & (!g22) & (ax12x) & (!bx12x)) + ((ax11x) & (!bx11x) & (!g20) & (g22) & (!ax12x) & (!bx12x)) + ((ax11x) & (!bx11x) & (g20) & (!g22) & (!ax12x) & (!bx12x)) + ((ax11x) & (!bx11x) & (g20) & (g22) & (!ax12x) & (!bx12x)) + ((ax11x) & (bx11x) & (!g20) & (!g22) & (!ax12x) & (!bx12x)) + ((ax11x) & (bx11x) & (!g20) & (g22) & (!ax12x) & (!bx12x)) + ((ax11x) & (bx11x) & (g20) & (!g22) & (!ax12x) & (!bx12x)) + ((ax11x) & (bx11x) & (g20) & (g22) & (!ax12x) & (!bx12x)));
	assign fx13x = (((!ax13x) & (!bx13x) & (!g26)) + ((!ax13x) & (bx13x) & (g26)) + ((ax13x) & (!bx13x) & (g26)) + ((ax13x) & (bx13x) & (!g26)));
	assign g28 = (((!ax13x) & (bx13x) & (!g26)) + ((ax13x) & (!bx13x) & (!g26)) + ((ax13x) & (bx13x) & (!g26)) + ((ax13x) & (bx13x) & (g26)));
	assign fx14x = (((!ax14x) & (!bx14x) & (g28)) + ((!ax14x) & (bx14x) & (!g28)) + ((ax14x) & (!bx14x) & (!g28)) + ((ax14x) & (bx14x) & (g28)));
	assign fx15x = (((!ax14x) & (!bx14x) & (!g28) & (!ax15x) & (bx15x)) + ((!ax14x) & (!bx14x) & (!g28) & (ax15x) & (!bx15x)) + ((!ax14x) & (!bx14x) & (g28) & (!ax15x) & (bx15x)) + ((!ax14x) & (!bx14x) & (g28) & (ax15x) & (!bx15x)) + ((!ax14x) & (bx14x) & (!g28) & (!ax15x) & (bx15x)) + ((!ax14x) & (bx14x) & (!g28) & (ax15x) & (!bx15x)) + ((!ax14x) & (bx14x) & (g28) & (!ax15x) & (!bx15x)) + ((!ax14x) & (bx14x) & (g28) & (ax15x) & (bx15x)) + ((ax14x) & (!bx14x) & (!g28) & (!ax15x) & (bx15x)) + ((ax14x) & (!bx14x) & (!g28) & (ax15x) & (!bx15x)) + ((ax14x) & (!bx14x) & (g28) & (!ax15x) & (!bx15x)) + ((ax14x) & (!bx14x) & (g28) & (ax15x) & (bx15x)) + ((ax14x) & (bx14x) & (!g28) & (!ax15x) & (!bx15x)) + ((ax14x) & (bx14x) & (!g28) & (ax15x) & (bx15x)) + ((ax14x) & (bx14x) & (g28) & (!ax15x) & (!bx15x)) + ((ax14x) & (bx14x) & (g28) & (ax15x) & (bx15x)));
	assign g31 = (((ax15x) & (bx15x)));
	assign g32 = (((!ax15x) & (!bx15x)));
	assign g33 = (((!ax13x) & (!bx13x) & (!g26) & (ax14x) & (bx14x) & (!g32)) + ((!ax13x) & (!bx13x) & (g26) & (ax14x) & (bx14x) & (!g32)) + ((!ax13x) & (bx13x) & (!g26) & (!ax14x) & (bx14x) & (!g32)) + ((!ax13x) & (bx13x) & (!g26) & (ax14x) & (!bx14x) & (!g32)) + ((!ax13x) & (bx13x) & (!g26) & (ax14x) & (bx14x) & (!g32)) + ((!ax13x) & (bx13x) & (g26) & (ax14x) & (bx14x) & (!g32)) + ((ax13x) & (!bx13x) & (!g26) & (!ax14x) & (bx14x) & (!g32)) + ((ax13x) & (!bx13x) & (!g26) & (ax14x) & (!bx14x) & (!g32)) + ((ax13x) & (!bx13x) & (!g26) & (ax14x) & (bx14x) & (!g32)) + ((ax13x) & (!bx13x) & (g26) & (ax14x) & (bx14x) & (!g32)) + ((ax13x) & (bx13x) & (!g26) & (!ax14x) & (bx14x) & (!g32)) + ((ax13x) & (bx13x) & (!g26) & (ax14x) & (!bx14x) & (!g32)) + ((ax13x) & (bx13x) & (!g26) & (ax14x) & (bx14x) & (!g32)) + ((ax13x) & (bx13x) & (g26) & (!ax14x) & (bx14x) & (!g32)) + ((ax13x) & (bx13x) & (g26) & (ax14x) & (!bx14x) & (!g32)) + ((ax13x) & (bx13x) & (g26) & (ax14x) & (bx14x) & (!g32)));
	assign g34 = (((!g31) & (!g33)));
	assign fx16x = (((!ax16x) & (!bx16x) & (!g34)) + ((!ax16x) & (bx16x) & (g34)) + ((ax16x) & (!bx16x) & (g34)) + ((ax16x) & (bx16x) & (!g34)));
	assign fx17x = (((!ax16x) & (!bx16x) & (!g34) & (!ax17x) & (bx17x)) + ((!ax16x) & (!bx16x) & (!g34) & (ax17x) & (!bx17x)) + ((!ax16x) & (!bx16x) & (g34) & (!ax17x) & (bx17x)) + ((!ax16x) & (!bx16x) & (g34) & (ax17x) & (!bx17x)) + ((!ax16x) & (bx16x) & (!g34) & (!ax17x) & (!bx17x)) + ((!ax16x) & (bx16x) & (!g34) & (ax17x) & (bx17x)) + ((!ax16x) & (bx16x) & (g34) & (!ax17x) & (bx17x)) + ((!ax16x) & (bx16x) & (g34) & (ax17x) & (!bx17x)) + ((ax16x) & (!bx16x) & (!g34) & (!ax17x) & (!bx17x)) + ((ax16x) & (!bx16x) & (!g34) & (ax17x) & (bx17x)) + ((ax16x) & (!bx16x) & (g34) & (!ax17x) & (bx17x)) + ((ax16x) & (!bx16x) & (g34) & (ax17x) & (!bx17x)) + ((ax16x) & (bx16x) & (!g34) & (!ax17x) & (!bx17x)) + ((ax16x) & (bx16x) & (!g34) & (ax17x) & (bx17x)) + ((ax16x) & (bx16x) & (g34) & (!ax17x) & (!bx17x)) + ((ax16x) & (bx16x) & (g34) & (ax17x) & (bx17x)));
	assign g37 = (((!ax16x) & (!bx16x) & (!g31) & (!g33) & (!ax17x) & (!bx17x)) + ((!ax16x) & (!bx16x) & (!g31) & (!g33) & (!ax17x) & (bx17x)) + ((!ax16x) & (!bx16x) & (!g31) & (!g33) & (ax17x) & (!bx17x)) + ((!ax16x) & (!bx16x) & (!g31) & (g33) & (!ax17x) & (!bx17x)) + ((!ax16x) & (!bx16x) & (!g31) & (g33) & (!ax17x) & (bx17x)) + ((!ax16x) & (!bx16x) & (!g31) & (g33) & (ax17x) & (!bx17x)) + ((!ax16x) & (!bx16x) & (g31) & (!g33) & (!ax17x) & (!bx17x)) + ((!ax16x) & (!bx16x) & (g31) & (!g33) & (!ax17x) & (bx17x)) + ((!ax16x) & (!bx16x) & (g31) & (!g33) & (ax17x) & (!bx17x)) + ((!ax16x) & (!bx16x) & (g31) & (g33) & (!ax17x) & (!bx17x)) + ((!ax16x) & (!bx16x) & (g31) & (g33) & (!ax17x) & (bx17x)) + ((!ax16x) & (!bx16x) & (g31) & (g33) & (ax17x) & (!bx17x)) + ((!ax16x) & (bx16x) & (!g31) & (!g33) & (!ax17x) & (!bx17x)) + ((!ax16x) & (bx16x) & (!g31) & (!g33) & (!ax17x) & (bx17x)) + ((!ax16x) & (bx16x) & (!g31) & (!g33) & (ax17x) & (!bx17x)) + ((!ax16x) & (bx16x) & (!g31) & (g33) & (!ax17x) & (!bx17x)) + ((!ax16x) & (bx16x) & (g31) & (!g33) & (!ax17x) & (!bx17x)) + ((!ax16x) & (bx16x) & (g31) & (g33) & (!ax17x) & (!bx17x)) + ((ax16x) & (!bx16x) & (!g31) & (!g33) & (!ax17x) & (!bx17x)) + ((ax16x) & (!bx16x) & (!g31) & (!g33) & (!ax17x) & (bx17x)) + ((ax16x) & (!bx16x) & (!g31) & (!g33) & (ax17x) & (!bx17x)) + ((ax16x) & (!bx16x) & (!g31) & (g33) & (!ax17x) & (!bx17x)) + ((ax16x) & (!bx16x) & (g31) & (!g33) & (!ax17x) & (!bx17x)) + ((ax16x) & (!bx16x) & (g31) & (g33) & (!ax17x) & (!bx17x)) + ((ax16x) & (bx16x) & (!g31) & (!g33) & (!ax17x) & (!bx17x)) + ((ax16x) & (bx16x) & (!g31) & (g33) & (!ax17x) & (!bx17x)) + ((ax16x) & (bx16x) & (g31) & (!g33) & (!ax17x) & (!bx17x)) + ((ax16x) & (bx16x) & (g31) & (g33) & (!ax17x) & (!bx17x)));
	assign fx18x = (((!ax18x) & (!bx18x) & (!g37)) + ((!ax18x) & (bx18x) & (g37)) + ((ax18x) & (!bx18x) & (g37)) + ((ax18x) & (bx18x) & (!g37)));
	assign g39 = (((!ax18x) & (bx18x) & (!g37)) + ((ax18x) & (!bx18x) & (!g37)) + ((ax18x) & (bx18x) & (!g37)) + ((ax18x) & (bx18x) & (g37)));
	assign fx19x = (((!ax19x) & (!bx19x) & (g39)) + ((!ax19x) & (bx19x) & (!g39)) + ((ax19x) & (!bx19x) & (!g39)) + ((ax19x) & (bx19x) & (g39)));
	assign fx20x = (((!ax19x) & (!bx19x) & (!g39) & (!ax20x) & (bx20x)) + ((!ax19x) & (!bx19x) & (!g39) & (ax20x) & (!bx20x)) + ((!ax19x) & (!bx19x) & (g39) & (!ax20x) & (bx20x)) + ((!ax19x) & (!bx19x) & (g39) & (ax20x) & (!bx20x)) + ((!ax19x) & (bx19x) & (!g39) & (!ax20x) & (bx20x)) + ((!ax19x) & (bx19x) & (!g39) & (ax20x) & (!bx20x)) + ((!ax19x) & (bx19x) & (g39) & (!ax20x) & (!bx20x)) + ((!ax19x) & (bx19x) & (g39) & (ax20x) & (bx20x)) + ((ax19x) & (!bx19x) & (!g39) & (!ax20x) & (bx20x)) + ((ax19x) & (!bx19x) & (!g39) & (ax20x) & (!bx20x)) + ((ax19x) & (!bx19x) & (g39) & (!ax20x) & (!bx20x)) + ((ax19x) & (!bx19x) & (g39) & (ax20x) & (bx20x)) + ((ax19x) & (bx19x) & (!g39) & (!ax20x) & (!bx20x)) + ((ax19x) & (bx19x) & (!g39) & (ax20x) & (bx20x)) + ((ax19x) & (bx19x) & (g39) & (!ax20x) & (!bx20x)) + ((ax19x) & (bx19x) & (g39) & (ax20x) & (bx20x)));
	assign g42 = (((ax20x) & (bx20x)));
	assign g43 = (((!ax20x) & (!bx20x)));
	assign g44 = (((!ax18x) & (!bx18x) & (!g37) & (ax19x) & (bx19x) & (!g43)) + ((!ax18x) & (!bx18x) & (g37) & (ax19x) & (bx19x) & (!g43)) + ((!ax18x) & (bx18x) & (!g37) & (!ax19x) & (bx19x) & (!g43)) + ((!ax18x) & (bx18x) & (!g37) & (ax19x) & (!bx19x) & (!g43)) + ((!ax18x) & (bx18x) & (!g37) & (ax19x) & (bx19x) & (!g43)) + ((!ax18x) & (bx18x) & (g37) & (ax19x) & (bx19x) & (!g43)) + ((ax18x) & (!bx18x) & (!g37) & (!ax19x) & (bx19x) & (!g43)) + ((ax18x) & (!bx18x) & (!g37) & (ax19x) & (!bx19x) & (!g43)) + ((ax18x) & (!bx18x) & (!g37) & (ax19x) & (bx19x) & (!g43)) + ((ax18x) & (!bx18x) & (g37) & (ax19x) & (bx19x) & (!g43)) + ((ax18x) & (bx18x) & (!g37) & (!ax19x) & (bx19x) & (!g43)) + ((ax18x) & (bx18x) & (!g37) & (ax19x) & (!bx19x) & (!g43)) + ((ax18x) & (bx18x) & (!g37) & (ax19x) & (bx19x) & (!g43)) + ((ax18x) & (bx18x) & (g37) & (!ax19x) & (bx19x) & (!g43)) + ((ax18x) & (bx18x) & (g37) & (ax19x) & (!bx19x) & (!g43)) + ((ax18x) & (bx18x) & (g37) & (ax19x) & (bx19x) & (!g43)));
	assign g45 = (((!g42) & (!g44)));
	assign fx21x = (((!ax21x) & (!bx21x) & (!g45)) + ((!ax21x) & (bx21x) & (g45)) + ((ax21x) & (!bx21x) & (g45)) + ((ax21x) & (bx21x) & (!g45)));
	assign fx22x = (((!ax21x) & (!bx21x) & (!g45) & (!ax22x) & (bx22x)) + ((!ax21x) & (!bx21x) & (!g45) & (ax22x) & (!bx22x)) + ((!ax21x) & (!bx21x) & (g45) & (!ax22x) & (bx22x)) + ((!ax21x) & (!bx21x) & (g45) & (ax22x) & (!bx22x)) + ((!ax21x) & (bx21x) & (!g45) & (!ax22x) & (!bx22x)) + ((!ax21x) & (bx21x) & (!g45) & (ax22x) & (bx22x)) + ((!ax21x) & (bx21x) & (g45) & (!ax22x) & (bx22x)) + ((!ax21x) & (bx21x) & (g45) & (ax22x) & (!bx22x)) + ((ax21x) & (!bx21x) & (!g45) & (!ax22x) & (!bx22x)) + ((ax21x) & (!bx21x) & (!g45) & (ax22x) & (bx22x)) + ((ax21x) & (!bx21x) & (g45) & (!ax22x) & (bx22x)) + ((ax21x) & (!bx21x) & (g45) & (ax22x) & (!bx22x)) + ((ax21x) & (bx21x) & (!g45) & (!ax22x) & (!bx22x)) + ((ax21x) & (bx21x) & (!g45) & (ax22x) & (bx22x)) + ((ax21x) & (bx21x) & (g45) & (!ax22x) & (!bx22x)) + ((ax21x) & (bx21x) & (g45) & (ax22x) & (bx22x)));
	assign g48 = (((!ax21x) & (!bx21x) & (!g42) & (!g44) & (!ax22x) & (!bx22x)) + ((!ax21x) & (!bx21x) & (!g42) & (!g44) & (!ax22x) & (bx22x)) + ((!ax21x) & (!bx21x) & (!g42) & (!g44) & (ax22x) & (!bx22x)) + ((!ax21x) & (!bx21x) & (!g42) & (g44) & (!ax22x) & (!bx22x)) + ((!ax21x) & (!bx21x) & (!g42) & (g44) & (!ax22x) & (bx22x)) + ((!ax21x) & (!bx21x) & (!g42) & (g44) & (ax22x) & (!bx22x)) + ((!ax21x) & (!bx21x) & (g42) & (!g44) & (!ax22x) & (!bx22x)) + ((!ax21x) & (!bx21x) & (g42) & (!g44) & (!ax22x) & (bx22x)) + ((!ax21x) & (!bx21x) & (g42) & (!g44) & (ax22x) & (!bx22x)) + ((!ax21x) & (!bx21x) & (g42) & (g44) & (!ax22x) & (!bx22x)) + ((!ax21x) & (!bx21x) & (g42) & (g44) & (!ax22x) & (bx22x)) + ((!ax21x) & (!bx21x) & (g42) & (g44) & (ax22x) & (!bx22x)) + ((!ax21x) & (bx21x) & (!g42) & (!g44) & (!ax22x) & (!bx22x)) + ((!ax21x) & (bx21x) & (!g42) & (!g44) & (!ax22x) & (bx22x)) + ((!ax21x) & (bx21x) & (!g42) & (!g44) & (ax22x) & (!bx22x)) + ((!ax21x) & (bx21x) & (!g42) & (g44) & (!ax22x) & (!bx22x)) + ((!ax21x) & (bx21x) & (g42) & (!g44) & (!ax22x) & (!bx22x)) + ((!ax21x) & (bx21x) & (g42) & (g44) & (!ax22x) & (!bx22x)) + ((ax21x) & (!bx21x) & (!g42) & (!g44) & (!ax22x) & (!bx22x)) + ((ax21x) & (!bx21x) & (!g42) & (!g44) & (!ax22x) & (bx22x)) + ((ax21x) & (!bx21x) & (!g42) & (!g44) & (ax22x) & (!bx22x)) + ((ax21x) & (!bx21x) & (!g42) & (g44) & (!ax22x) & (!bx22x)) + ((ax21x) & (!bx21x) & (g42) & (!g44) & (!ax22x) & (!bx22x)) + ((ax21x) & (!bx21x) & (g42) & (g44) & (!ax22x) & (!bx22x)) + ((ax21x) & (bx21x) & (!g42) & (!g44) & (!ax22x) & (!bx22x)) + ((ax21x) & (bx21x) & (!g42) & (g44) & (!ax22x) & (!bx22x)) + ((ax21x) & (bx21x) & (g42) & (!g44) & (!ax22x) & (!bx22x)) + ((ax21x) & (bx21x) & (g42) & (g44) & (!ax22x) & (!bx22x)));
	assign fx23x = (((!ax23x) & (!bx23x) & (!g48)) + ((!ax23x) & (bx23x) & (g48)) + ((ax23x) & (!bx23x) & (g48)) + ((ax23x) & (bx23x) & (!g48)));
	assign g50 = (((!ax23x) & (bx23x) & (!g48)) + ((ax23x) & (!bx23x) & (!g48)) + ((ax23x) & (bx23x) & (!g48)) + ((ax23x) & (bx23x) & (g48)));
	assign fx24x = (((!ax24x) & (!bx24x) & (g50)) + ((!ax24x) & (bx24x) & (!g50)) + ((ax24x) & (!bx24x) & (!g50)) + ((ax24x) & (bx24x) & (g50)));
	assign fx25x = (((!ax24x) & (!bx24x) & (!g50) & (!ax25x) & (bx25x)) + ((!ax24x) & (!bx24x) & (!g50) & (ax25x) & (!bx25x)) + ((!ax24x) & (!bx24x) & (g50) & (!ax25x) & (bx25x)) + ((!ax24x) & (!bx24x) & (g50) & (ax25x) & (!bx25x)) + ((!ax24x) & (bx24x) & (!g50) & (!ax25x) & (bx25x)) + ((!ax24x) & (bx24x) & (!g50) & (ax25x) & (!bx25x)) + ((!ax24x) & (bx24x) & (g50) & (!ax25x) & (!bx25x)) + ((!ax24x) & (bx24x) & (g50) & (ax25x) & (bx25x)) + ((ax24x) & (!bx24x) & (!g50) & (!ax25x) & (bx25x)) + ((ax24x) & (!bx24x) & (!g50) & (ax25x) & (!bx25x)) + ((ax24x) & (!bx24x) & (g50) & (!ax25x) & (!bx25x)) + ((ax24x) & (!bx24x) & (g50) & (ax25x) & (bx25x)) + ((ax24x) & (bx24x) & (!g50) & (!ax25x) & (!bx25x)) + ((ax24x) & (bx24x) & (!g50) & (ax25x) & (bx25x)) + ((ax24x) & (bx24x) & (g50) & (!ax25x) & (!bx25x)) + ((ax24x) & (bx24x) & (g50) & (ax25x) & (bx25x)));
	assign g53 = (((ax25x) & (bx25x)));
	assign g54 = (((!ax25x) & (!bx25x)));
	assign g55 = (((!ax23x) & (!bx23x) & (!g48) & (ax24x) & (bx24x) & (!g54)) + ((!ax23x) & (!bx23x) & (g48) & (ax24x) & (bx24x) & (!g54)) + ((!ax23x) & (bx23x) & (!g48) & (!ax24x) & (bx24x) & (!g54)) + ((!ax23x) & (bx23x) & (!g48) & (ax24x) & (!bx24x) & (!g54)) + ((!ax23x) & (bx23x) & (!g48) & (ax24x) & (bx24x) & (!g54)) + ((!ax23x) & (bx23x) & (g48) & (ax24x) & (bx24x) & (!g54)) + ((ax23x) & (!bx23x) & (!g48) & (!ax24x) & (bx24x) & (!g54)) + ((ax23x) & (!bx23x) & (!g48) & (ax24x) & (!bx24x) & (!g54)) + ((ax23x) & (!bx23x) & (!g48) & (ax24x) & (bx24x) & (!g54)) + ((ax23x) & (!bx23x) & (g48) & (ax24x) & (bx24x) & (!g54)) + ((ax23x) & (bx23x) & (!g48) & (!ax24x) & (bx24x) & (!g54)) + ((ax23x) & (bx23x) & (!g48) & (ax24x) & (!bx24x) & (!g54)) + ((ax23x) & (bx23x) & (!g48) & (ax24x) & (bx24x) & (!g54)) + ((ax23x) & (bx23x) & (g48) & (!ax24x) & (bx24x) & (!g54)) + ((ax23x) & (bx23x) & (g48) & (ax24x) & (!bx24x) & (!g54)) + ((ax23x) & (bx23x) & (g48) & (ax24x) & (bx24x) & (!g54)));
	assign g56 = (((!g53) & (!g55)));
	assign fx26x = (((!ax26x) & (!bx26x) & (!g56)) + ((!ax26x) & (bx26x) & (g56)) + ((ax26x) & (!bx26x) & (g56)) + ((ax26x) & (bx26x) & (!g56)));
	assign fx27x = (((!ax26x) & (!bx26x) & (!g56) & (!ax27x) & (bx27x)) + ((!ax26x) & (!bx26x) & (!g56) & (ax27x) & (!bx27x)) + ((!ax26x) & (!bx26x) & (g56) & (!ax27x) & (bx27x)) + ((!ax26x) & (!bx26x) & (g56) & (ax27x) & (!bx27x)) + ((!ax26x) & (bx26x) & (!g56) & (!ax27x) & (!bx27x)) + ((!ax26x) & (bx26x) & (!g56) & (ax27x) & (bx27x)) + ((!ax26x) & (bx26x) & (g56) & (!ax27x) & (bx27x)) + ((!ax26x) & (bx26x) & (g56) & (ax27x) & (!bx27x)) + ((ax26x) & (!bx26x) & (!g56) & (!ax27x) & (!bx27x)) + ((ax26x) & (!bx26x) & (!g56) & (ax27x) & (bx27x)) + ((ax26x) & (!bx26x) & (g56) & (!ax27x) & (bx27x)) + ((ax26x) & (!bx26x) & (g56) & (ax27x) & (!bx27x)) + ((ax26x) & (bx26x) & (!g56) & (!ax27x) & (!bx27x)) + ((ax26x) & (bx26x) & (!g56) & (ax27x) & (bx27x)) + ((ax26x) & (bx26x) & (g56) & (!ax27x) & (!bx27x)) + ((ax26x) & (bx26x) & (g56) & (ax27x) & (bx27x)));
	assign g59 = (((!ax26x) & (!bx26x) & (!g53) & (!g55) & (!ax27x) & (!bx27x)) + ((!ax26x) & (!bx26x) & (!g53) & (!g55) & (!ax27x) & (bx27x)) + ((!ax26x) & (!bx26x) & (!g53) & (!g55) & (ax27x) & (!bx27x)) + ((!ax26x) & (!bx26x) & (!g53) & (g55) & (!ax27x) & (!bx27x)) + ((!ax26x) & (!bx26x) & (!g53) & (g55) & (!ax27x) & (bx27x)) + ((!ax26x) & (!bx26x) & (!g53) & (g55) & (ax27x) & (!bx27x)) + ((!ax26x) & (!bx26x) & (g53) & (!g55) & (!ax27x) & (!bx27x)) + ((!ax26x) & (!bx26x) & (g53) & (!g55) & (!ax27x) & (bx27x)) + ((!ax26x) & (!bx26x) & (g53) & (!g55) & (ax27x) & (!bx27x)) + ((!ax26x) & (!bx26x) & (g53) & (g55) & (!ax27x) & (!bx27x)) + ((!ax26x) & (!bx26x) & (g53) & (g55) & (!ax27x) & (bx27x)) + ((!ax26x) & (!bx26x) & (g53) & (g55) & (ax27x) & (!bx27x)) + ((!ax26x) & (bx26x) & (!g53) & (!g55) & (!ax27x) & (!bx27x)) + ((!ax26x) & (bx26x) & (!g53) & (!g55) & (!ax27x) & (bx27x)) + ((!ax26x) & (bx26x) & (!g53) & (!g55) & (ax27x) & (!bx27x)) + ((!ax26x) & (bx26x) & (!g53) & (g55) & (!ax27x) & (!bx27x)) + ((!ax26x) & (bx26x) & (g53) & (!g55) & (!ax27x) & (!bx27x)) + ((!ax26x) & (bx26x) & (g53) & (g55) & (!ax27x) & (!bx27x)) + ((ax26x) & (!bx26x) & (!g53) & (!g55) & (!ax27x) & (!bx27x)) + ((ax26x) & (!bx26x) & (!g53) & (!g55) & (!ax27x) & (bx27x)) + ((ax26x) & (!bx26x) & (!g53) & (!g55) & (ax27x) & (!bx27x)) + ((ax26x) & (!bx26x) & (!g53) & (g55) & (!ax27x) & (!bx27x)) + ((ax26x) & (!bx26x) & (g53) & (!g55) & (!ax27x) & (!bx27x)) + ((ax26x) & (!bx26x) & (g53) & (g55) & (!ax27x) & (!bx27x)) + ((ax26x) & (bx26x) & (!g53) & (!g55) & (!ax27x) & (!bx27x)) + ((ax26x) & (bx26x) & (!g53) & (g55) & (!ax27x) & (!bx27x)) + ((ax26x) & (bx26x) & (g53) & (!g55) & (!ax27x) & (!bx27x)) + ((ax26x) & (bx26x) & (g53) & (g55) & (!ax27x) & (!bx27x)));
	assign fx28x = (((!ax28x) & (!bx28x) & (!g59)) + ((!ax28x) & (bx28x) & (g59)) + ((ax28x) & (!bx28x) & (g59)) + ((ax28x) & (bx28x) & (!g59)));
	assign g61 = (((!ax28x) & (bx28x) & (!g59)) + ((ax28x) & (!bx28x) & (!g59)) + ((ax28x) & (bx28x) & (!g59)) + ((ax28x) & (bx28x) & (g59)));
	assign fx29x = (((!ax29x) & (!bx29x) & (g61)) + ((!ax29x) & (bx29x) & (!g61)) + ((ax29x) & (!bx29x) & (!g61)) + ((ax29x) & (bx29x) & (g61)));
	assign fx30x = (((!ax29x) & (!bx29x) & (!g61) & (!ax30x) & (bx30x)) + ((!ax29x) & (!bx29x) & (!g61) & (ax30x) & (!bx30x)) + ((!ax29x) & (!bx29x) & (g61) & (!ax30x) & (bx30x)) + ((!ax29x) & (!bx29x) & (g61) & (ax30x) & (!bx30x)) + ((!ax29x) & (bx29x) & (!g61) & (!ax30x) & (bx30x)) + ((!ax29x) & (bx29x) & (!g61) & (ax30x) & (!bx30x)) + ((!ax29x) & (bx29x) & (g61) & (!ax30x) & (!bx30x)) + ((!ax29x) & (bx29x) & (g61) & (ax30x) & (bx30x)) + ((ax29x) & (!bx29x) & (!g61) & (!ax30x) & (bx30x)) + ((ax29x) & (!bx29x) & (!g61) & (ax30x) & (!bx30x)) + ((ax29x) & (!bx29x) & (g61) & (!ax30x) & (!bx30x)) + ((ax29x) & (!bx29x) & (g61) & (ax30x) & (bx30x)) + ((ax29x) & (bx29x) & (!g61) & (!ax30x) & (!bx30x)) + ((ax29x) & (bx29x) & (!g61) & (ax30x) & (bx30x)) + ((ax29x) & (bx29x) & (g61) & (!ax30x) & (!bx30x)) + ((ax29x) & (bx29x) & (g61) & (ax30x) & (bx30x)));
	assign g64 = (((ax30x) & (bx30x)));
	assign g65 = (((!ax30x) & (!bx30x)));
	assign g66 = (((!ax28x) & (!bx28x) & (!g59) & (ax29x) & (bx29x) & (!g65)) + ((!ax28x) & (!bx28x) & (g59) & (ax29x) & (bx29x) & (!g65)) + ((!ax28x) & (bx28x) & (!g59) & (!ax29x) & (bx29x) & (!g65)) + ((!ax28x) & (bx28x) & (!g59) & (ax29x) & (!bx29x) & (!g65)) + ((!ax28x) & (bx28x) & (!g59) & (ax29x) & (bx29x) & (!g65)) + ((!ax28x) & (bx28x) & (g59) & (ax29x) & (bx29x) & (!g65)) + ((ax28x) & (!bx28x) & (!g59) & (!ax29x) & (bx29x) & (!g65)) + ((ax28x) & (!bx28x) & (!g59) & (ax29x) & (!bx29x) & (!g65)) + ((ax28x) & (!bx28x) & (!g59) & (ax29x) & (bx29x) & (!g65)) + ((ax28x) & (!bx28x) & (g59) & (ax29x) & (bx29x) & (!g65)) + ((ax28x) & (bx28x) & (!g59) & (!ax29x) & (bx29x) & (!g65)) + ((ax28x) & (bx28x) & (!g59) & (ax29x) & (!bx29x) & (!g65)) + ((ax28x) & (bx28x) & (!g59) & (ax29x) & (bx29x) & (!g65)) + ((ax28x) & (bx28x) & (g59) & (!ax29x) & (bx29x) & (!g65)) + ((ax28x) & (bx28x) & (g59) & (ax29x) & (!bx29x) & (!g65)) + ((ax28x) & (bx28x) & (g59) & (ax29x) & (bx29x) & (!g65)));
	assign g67 = (((!g64) & (!g66)));
	assign fx31x = (((!ax31x) & (!bx31x) & (!g67)) + ((!ax31x) & (bx31x) & (g67)) + ((ax31x) & (!bx31x) & (g67)) + ((ax31x) & (bx31x) & (!g67)));
	assign fx32x = (((!ax31x) & (!bx31x) & (!g67) & (!ax32x) & (bx32x)) + ((!ax31x) & (!bx31x) & (!g67) & (ax32x) & (!bx32x)) + ((!ax31x) & (!bx31x) & (g67) & (!ax32x) & (bx32x)) + ((!ax31x) & (!bx31x) & (g67) & (ax32x) & (!bx32x)) + ((!ax31x) & (bx31x) & (!g67) & (!ax32x) & (!bx32x)) + ((!ax31x) & (bx31x) & (!g67) & (ax32x) & (bx32x)) + ((!ax31x) & (bx31x) & (g67) & (!ax32x) & (bx32x)) + ((!ax31x) & (bx31x) & (g67) & (ax32x) & (!bx32x)) + ((ax31x) & (!bx31x) & (!g67) & (!ax32x) & (!bx32x)) + ((ax31x) & (!bx31x) & (!g67) & (ax32x) & (bx32x)) + ((ax31x) & (!bx31x) & (g67) & (!ax32x) & (bx32x)) + ((ax31x) & (!bx31x) & (g67) & (ax32x) & (!bx32x)) + ((ax31x) & (bx31x) & (!g67) & (!ax32x) & (!bx32x)) + ((ax31x) & (bx31x) & (!g67) & (ax32x) & (bx32x)) + ((ax31x) & (bx31x) & (g67) & (!ax32x) & (!bx32x)) + ((ax31x) & (bx31x) & (g67) & (ax32x) & (bx32x)));
	assign g70 = (((!ax31x) & (!bx31x) & (!g64) & (!g66) & (!ax32x) & (!bx32x)) + ((!ax31x) & (!bx31x) & (!g64) & (!g66) & (!ax32x) & (bx32x)) + ((!ax31x) & (!bx31x) & (!g64) & (!g66) & (ax32x) & (!bx32x)) + ((!ax31x) & (!bx31x) & (!g64) & (g66) & (!ax32x) & (!bx32x)) + ((!ax31x) & (!bx31x) & (!g64) & (g66) & (!ax32x) & (bx32x)) + ((!ax31x) & (!bx31x) & (!g64) & (g66) & (ax32x) & (!bx32x)) + ((!ax31x) & (!bx31x) & (g64) & (!g66) & (!ax32x) & (!bx32x)) + ((!ax31x) & (!bx31x) & (g64) & (!g66) & (!ax32x) & (bx32x)) + ((!ax31x) & (!bx31x) & (g64) & (!g66) & (ax32x) & (!bx32x)) + ((!ax31x) & (!bx31x) & (g64) & (g66) & (!ax32x) & (!bx32x)) + ((!ax31x) & (!bx31x) & (g64) & (g66) & (!ax32x) & (bx32x)) + ((!ax31x) & (!bx31x) & (g64) & (g66) & (ax32x) & (!bx32x)) + ((!ax31x) & (bx31x) & (!g64) & (!g66) & (!ax32x) & (!bx32x)) + ((!ax31x) & (bx31x) & (!g64) & (!g66) & (!ax32x) & (bx32x)) + ((!ax31x) & (bx31x) & (!g64) & (!g66) & (ax32x) & (!bx32x)) + ((!ax31x) & (bx31x) & (!g64) & (g66) & (!ax32x) & (!bx32x)) + ((!ax31x) & (bx31x) & (g64) & (!g66) & (!ax32x) & (!bx32x)) + ((!ax31x) & (bx31x) & (g64) & (g66) & (!ax32x) & (!bx32x)) + ((ax31x) & (!bx31x) & (!g64) & (!g66) & (!ax32x) & (!bx32x)) + ((ax31x) & (!bx31x) & (!g64) & (!g66) & (!ax32x) & (bx32x)) + ((ax31x) & (!bx31x) & (!g64) & (!g66) & (ax32x) & (!bx32x)) + ((ax31x) & (!bx31x) & (!g64) & (g66) & (!ax32x) & (!bx32x)) + ((ax31x) & (!bx31x) & (g64) & (!g66) & (!ax32x) & (!bx32x)) + ((ax31x) & (!bx31x) & (g64) & (g66) & (!ax32x) & (!bx32x)) + ((ax31x) & (bx31x) & (!g64) & (!g66) & (!ax32x) & (!bx32x)) + ((ax31x) & (bx31x) & (!g64) & (g66) & (!ax32x) & (!bx32x)) + ((ax31x) & (bx31x) & (g64) & (!g66) & (!ax32x) & (!bx32x)) + ((ax31x) & (bx31x) & (g64) & (g66) & (!ax32x) & (!bx32x)));
	assign fx33x = (((!ax33x) & (!bx33x) & (!g70)) + ((!ax33x) & (bx33x) & (g70)) + ((ax33x) & (!bx33x) & (g70)) + ((ax33x) & (bx33x) & (!g70)));
	assign g72 = (((!ax33x) & (bx33x) & (!g70)) + ((ax33x) & (!bx33x) & (!g70)) + ((ax33x) & (bx33x) & (!g70)) + ((ax33x) & (bx33x) & (g70)));
	assign fx34x = (((!ax34x) & (!bx34x) & (g72)) + ((!ax34x) & (bx34x) & (!g72)) + ((ax34x) & (!bx34x) & (!g72)) + ((ax34x) & (bx34x) & (g72)));
	assign fx35x = (((!ax34x) & (!bx34x) & (!g72) & (!ax35x) & (bx35x)) + ((!ax34x) & (!bx34x) & (!g72) & (ax35x) & (!bx35x)) + ((!ax34x) & (!bx34x) & (g72) & (!ax35x) & (bx35x)) + ((!ax34x) & (!bx34x) & (g72) & (ax35x) & (!bx35x)) + ((!ax34x) & (bx34x) & (!g72) & (!ax35x) & (bx35x)) + ((!ax34x) & (bx34x) & (!g72) & (ax35x) & (!bx35x)) + ((!ax34x) & (bx34x) & (g72) & (!ax35x) & (!bx35x)) + ((!ax34x) & (bx34x) & (g72) & (ax35x) & (bx35x)) + ((ax34x) & (!bx34x) & (!g72) & (!ax35x) & (bx35x)) + ((ax34x) & (!bx34x) & (!g72) & (ax35x) & (!bx35x)) + ((ax34x) & (!bx34x) & (g72) & (!ax35x) & (!bx35x)) + ((ax34x) & (!bx34x) & (g72) & (ax35x) & (bx35x)) + ((ax34x) & (bx34x) & (!g72) & (!ax35x) & (!bx35x)) + ((ax34x) & (bx34x) & (!g72) & (ax35x) & (bx35x)) + ((ax34x) & (bx34x) & (g72) & (!ax35x) & (!bx35x)) + ((ax34x) & (bx34x) & (g72) & (ax35x) & (bx35x)));
	assign g75 = (((ax35x) & (bx35x)));
	assign g76 = (((!ax35x) & (!bx35x)));
	assign g77 = (((!ax33x) & (!bx33x) & (!g70) & (ax34x) & (bx34x) & (!g76)) + ((!ax33x) & (!bx33x) & (g70) & (ax34x) & (bx34x) & (!g76)) + ((!ax33x) & (bx33x) & (!g70) & (!ax34x) & (bx34x) & (!g76)) + ((!ax33x) & (bx33x) & (!g70) & (ax34x) & (!bx34x) & (!g76)) + ((!ax33x) & (bx33x) & (!g70) & (ax34x) & (bx34x) & (!g76)) + ((!ax33x) & (bx33x) & (g70) & (ax34x) & (bx34x) & (!g76)) + ((ax33x) & (!bx33x) & (!g70) & (!ax34x) & (bx34x) & (!g76)) + ((ax33x) & (!bx33x) & (!g70) & (ax34x) & (!bx34x) & (!g76)) + ((ax33x) & (!bx33x) & (!g70) & (ax34x) & (bx34x) & (!g76)) + ((ax33x) & (!bx33x) & (g70) & (ax34x) & (bx34x) & (!g76)) + ((ax33x) & (bx33x) & (!g70) & (!ax34x) & (bx34x) & (!g76)) + ((ax33x) & (bx33x) & (!g70) & (ax34x) & (!bx34x) & (!g76)) + ((ax33x) & (bx33x) & (!g70) & (ax34x) & (bx34x) & (!g76)) + ((ax33x) & (bx33x) & (g70) & (!ax34x) & (bx34x) & (!g76)) + ((ax33x) & (bx33x) & (g70) & (ax34x) & (!bx34x) & (!g76)) + ((ax33x) & (bx33x) & (g70) & (ax34x) & (bx34x) & (!g76)));
	assign g78 = (((!g75) & (!g77)));
	assign fx36x = (((!ax36x) & (!bx36x) & (!g78)) + ((!ax36x) & (bx36x) & (g78)) + ((ax36x) & (!bx36x) & (g78)) + ((ax36x) & (bx36x) & (!g78)));
	assign fx37x = (((!ax36x) & (!bx36x) & (!g78) & (!ax37x) & (bx37x)) + ((!ax36x) & (!bx36x) & (!g78) & (ax37x) & (!bx37x)) + ((!ax36x) & (!bx36x) & (g78) & (!ax37x) & (bx37x)) + ((!ax36x) & (!bx36x) & (g78) & (ax37x) & (!bx37x)) + ((!ax36x) & (bx36x) & (!g78) & (!ax37x) & (!bx37x)) + ((!ax36x) & (bx36x) & (!g78) & (ax37x) & (bx37x)) + ((!ax36x) & (bx36x) & (g78) & (!ax37x) & (bx37x)) + ((!ax36x) & (bx36x) & (g78) & (ax37x) & (!bx37x)) + ((ax36x) & (!bx36x) & (!g78) & (!ax37x) & (!bx37x)) + ((ax36x) & (!bx36x) & (!g78) & (ax37x) & (bx37x)) + ((ax36x) & (!bx36x) & (g78) & (!ax37x) & (bx37x)) + ((ax36x) & (!bx36x) & (g78) & (ax37x) & (!bx37x)) + ((ax36x) & (bx36x) & (!g78) & (!ax37x) & (!bx37x)) + ((ax36x) & (bx36x) & (!g78) & (ax37x) & (bx37x)) + ((ax36x) & (bx36x) & (g78) & (!ax37x) & (!bx37x)) + ((ax36x) & (bx36x) & (g78) & (ax37x) & (bx37x)));
	assign g81 = (((!ax36x) & (!bx36x) & (!g75) & (!g77) & (!ax37x) & (!bx37x)) + ((!ax36x) & (!bx36x) & (!g75) & (!g77) & (!ax37x) & (bx37x)) + ((!ax36x) & (!bx36x) & (!g75) & (!g77) & (ax37x) & (!bx37x)) + ((!ax36x) & (!bx36x) & (!g75) & (g77) & (!ax37x) & (!bx37x)) + ((!ax36x) & (!bx36x) & (!g75) & (g77) & (!ax37x) & (bx37x)) + ((!ax36x) & (!bx36x) & (!g75) & (g77) & (ax37x) & (!bx37x)) + ((!ax36x) & (!bx36x) & (g75) & (!g77) & (!ax37x) & (!bx37x)) + ((!ax36x) & (!bx36x) & (g75) & (!g77) & (!ax37x) & (bx37x)) + ((!ax36x) & (!bx36x) & (g75) & (!g77) & (ax37x) & (!bx37x)) + ((!ax36x) & (!bx36x) & (g75) & (g77) & (!ax37x) & (!bx37x)) + ((!ax36x) & (!bx36x) & (g75) & (g77) & (!ax37x) & (bx37x)) + ((!ax36x) & (!bx36x) & (g75) & (g77) & (ax37x) & (!bx37x)) + ((!ax36x) & (bx36x) & (!g75) & (!g77) & (!ax37x) & (!bx37x)) + ((!ax36x) & (bx36x) & (!g75) & (!g77) & (!ax37x) & (bx37x)) + ((!ax36x) & (bx36x) & (!g75) & (!g77) & (ax37x) & (!bx37x)) + ((!ax36x) & (bx36x) & (!g75) & (g77) & (!ax37x) & (!bx37x)) + ((!ax36x) & (bx36x) & (g75) & (!g77) & (!ax37x) & (!bx37x)) + ((!ax36x) & (bx36x) & (g75) & (g77) & (!ax37x) & (!bx37x)) + ((ax36x) & (!bx36x) & (!g75) & (!g77) & (!ax37x) & (!bx37x)) + ((ax36x) & (!bx36x) & (!g75) & (!g77) & (!ax37x) & (bx37x)) + ((ax36x) & (!bx36x) & (!g75) & (!g77) & (ax37x) & (!bx37x)) + ((ax36x) & (!bx36x) & (!g75) & (g77) & (!ax37x) & (!bx37x)) + ((ax36x) & (!bx36x) & (g75) & (!g77) & (!ax37x) & (!bx37x)) + ((ax36x) & (!bx36x) & (g75) & (g77) & (!ax37x) & (!bx37x)) + ((ax36x) & (bx36x) & (!g75) & (!g77) & (!ax37x) & (!bx37x)) + ((ax36x) & (bx36x) & (!g75) & (g77) & (!ax37x) & (!bx37x)) + ((ax36x) & (bx36x) & (g75) & (!g77) & (!ax37x) & (!bx37x)) + ((ax36x) & (bx36x) & (g75) & (g77) & (!ax37x) & (!bx37x)));
	assign fx38x = (((!ax38x) & (!bx38x) & (!g81)) + ((!ax38x) & (bx38x) & (g81)) + ((ax38x) & (!bx38x) & (g81)) + ((ax38x) & (bx38x) & (!g81)));
	assign g83 = (((!ax38x) & (bx38x) & (!g81)) + ((ax38x) & (!bx38x) & (!g81)) + ((ax38x) & (bx38x) & (!g81)) + ((ax38x) & (bx38x) & (g81)));
	assign fx39x = (((!ax39x) & (!bx39x) & (g83)) + ((!ax39x) & (bx39x) & (!g83)) + ((ax39x) & (!bx39x) & (!g83)) + ((ax39x) & (bx39x) & (g83)));
	assign fx40x = (((!ax39x) & (!bx39x) & (!g83) & (!ax40x) & (bx40x)) + ((!ax39x) & (!bx39x) & (!g83) & (ax40x) & (!bx40x)) + ((!ax39x) & (!bx39x) & (g83) & (!ax40x) & (bx40x)) + ((!ax39x) & (!bx39x) & (g83) & (ax40x) & (!bx40x)) + ((!ax39x) & (bx39x) & (!g83) & (!ax40x) & (bx40x)) + ((!ax39x) & (bx39x) & (!g83) & (ax40x) & (!bx40x)) + ((!ax39x) & (bx39x) & (g83) & (!ax40x) & (!bx40x)) + ((!ax39x) & (bx39x) & (g83) & (ax40x) & (bx40x)) + ((ax39x) & (!bx39x) & (!g83) & (!ax40x) & (bx40x)) + ((ax39x) & (!bx39x) & (!g83) & (ax40x) & (!bx40x)) + ((ax39x) & (!bx39x) & (g83) & (!ax40x) & (!bx40x)) + ((ax39x) & (!bx39x) & (g83) & (ax40x) & (bx40x)) + ((ax39x) & (bx39x) & (!g83) & (!ax40x) & (!bx40x)) + ((ax39x) & (bx39x) & (!g83) & (ax40x) & (bx40x)) + ((ax39x) & (bx39x) & (g83) & (!ax40x) & (!bx40x)) + ((ax39x) & (bx39x) & (g83) & (ax40x) & (bx40x)));
	assign g86 = (((ax40x) & (bx40x)));
	assign g87 = (((!ax40x) & (!bx40x)));
	assign g88 = (((!ax38x) & (!bx38x) & (!g81) & (ax39x) & (bx39x) & (!g87)) + ((!ax38x) & (!bx38x) & (g81) & (ax39x) & (bx39x) & (!g87)) + ((!ax38x) & (bx38x) & (!g81) & (!ax39x) & (bx39x) & (!g87)) + ((!ax38x) & (bx38x) & (!g81) & (ax39x) & (!bx39x) & (!g87)) + ((!ax38x) & (bx38x) & (!g81) & (ax39x) & (bx39x) & (!g87)) + ((!ax38x) & (bx38x) & (g81) & (ax39x) & (bx39x) & (!g87)) + ((ax38x) & (!bx38x) & (!g81) & (!ax39x) & (bx39x) & (!g87)) + ((ax38x) & (!bx38x) & (!g81) & (ax39x) & (!bx39x) & (!g87)) + ((ax38x) & (!bx38x) & (!g81) & (ax39x) & (bx39x) & (!g87)) + ((ax38x) & (!bx38x) & (g81) & (ax39x) & (bx39x) & (!g87)) + ((ax38x) & (bx38x) & (!g81) & (!ax39x) & (bx39x) & (!g87)) + ((ax38x) & (bx38x) & (!g81) & (ax39x) & (!bx39x) & (!g87)) + ((ax38x) & (bx38x) & (!g81) & (ax39x) & (bx39x) & (!g87)) + ((ax38x) & (bx38x) & (g81) & (!ax39x) & (bx39x) & (!g87)) + ((ax38x) & (bx38x) & (g81) & (ax39x) & (!bx39x) & (!g87)) + ((ax38x) & (bx38x) & (g81) & (ax39x) & (bx39x) & (!g87)));
	assign g89 = (((!g86) & (!g88)));
	assign fx41x = (((!ax41x) & (!bx41x) & (!g89)) + ((!ax41x) & (bx41x) & (g89)) + ((ax41x) & (!bx41x) & (g89)) + ((ax41x) & (bx41x) & (!g89)));
	assign fx42x = (((!ax41x) & (!bx41x) & (!g89) & (!ax42x) & (bx42x)) + ((!ax41x) & (!bx41x) & (!g89) & (ax42x) & (!bx42x)) + ((!ax41x) & (!bx41x) & (g89) & (!ax42x) & (bx42x)) + ((!ax41x) & (!bx41x) & (g89) & (ax42x) & (!bx42x)) + ((!ax41x) & (bx41x) & (!g89) & (!ax42x) & (!bx42x)) + ((!ax41x) & (bx41x) & (!g89) & (ax42x) & (bx42x)) + ((!ax41x) & (bx41x) & (g89) & (!ax42x) & (bx42x)) + ((!ax41x) & (bx41x) & (g89) & (ax42x) & (!bx42x)) + ((ax41x) & (!bx41x) & (!g89) & (!ax42x) & (!bx42x)) + ((ax41x) & (!bx41x) & (!g89) & (ax42x) & (bx42x)) + ((ax41x) & (!bx41x) & (g89) & (!ax42x) & (bx42x)) + ((ax41x) & (!bx41x) & (g89) & (ax42x) & (!bx42x)) + ((ax41x) & (bx41x) & (!g89) & (!ax42x) & (!bx42x)) + ((ax41x) & (bx41x) & (!g89) & (ax42x) & (bx42x)) + ((ax41x) & (bx41x) & (g89) & (!ax42x) & (!bx42x)) + ((ax41x) & (bx41x) & (g89) & (ax42x) & (bx42x)));
	assign g92 = (((!ax41x) & (!bx41x) & (!g86) & (!g88) & (!ax42x) & (!bx42x)) + ((!ax41x) & (!bx41x) & (!g86) & (!g88) & (!ax42x) & (bx42x)) + ((!ax41x) & (!bx41x) & (!g86) & (!g88) & (ax42x) & (!bx42x)) + ((!ax41x) & (!bx41x) & (!g86) & (g88) & (!ax42x) & (!bx42x)) + ((!ax41x) & (!bx41x) & (!g86) & (g88) & (!ax42x) & (bx42x)) + ((!ax41x) & (!bx41x) & (!g86) & (g88) & (ax42x) & (!bx42x)) + ((!ax41x) & (!bx41x) & (g86) & (!g88) & (!ax42x) & (!bx42x)) + ((!ax41x) & (!bx41x) & (g86) & (!g88) & (!ax42x) & (bx42x)) + ((!ax41x) & (!bx41x) & (g86) & (!g88) & (ax42x) & (!bx42x)) + ((!ax41x) & (!bx41x) & (g86) & (g88) & (!ax42x) & (!bx42x)) + ((!ax41x) & (!bx41x) & (g86) & (g88) & (!ax42x) & (bx42x)) + ((!ax41x) & (!bx41x) & (g86) & (g88) & (ax42x) & (!bx42x)) + ((!ax41x) & (bx41x) & (!g86) & (!g88) & (!ax42x) & (!bx42x)) + ((!ax41x) & (bx41x) & (!g86) & (!g88) & (!ax42x) & (bx42x)) + ((!ax41x) & (bx41x) & (!g86) & (!g88) & (ax42x) & (!bx42x)) + ((!ax41x) & (bx41x) & (!g86) & (g88) & (!ax42x) & (!bx42x)) + ((!ax41x) & (bx41x) & (g86) & (!g88) & (!ax42x) & (!bx42x)) + ((!ax41x) & (bx41x) & (g86) & (g88) & (!ax42x) & (!bx42x)) + ((ax41x) & (!bx41x) & (!g86) & (!g88) & (!ax42x) & (!bx42x)) + ((ax41x) & (!bx41x) & (!g86) & (!g88) & (!ax42x) & (bx42x)) + ((ax41x) & (!bx41x) & (!g86) & (!g88) & (ax42x) & (!bx42x)) + ((ax41x) & (!bx41x) & (!g86) & (g88) & (!ax42x) & (!bx42x)) + ((ax41x) & (!bx41x) & (g86) & (!g88) & (!ax42x) & (!bx42x)) + ((ax41x) & (!bx41x) & (g86) & (g88) & (!ax42x) & (!bx42x)) + ((ax41x) & (bx41x) & (!g86) & (!g88) & (!ax42x) & (!bx42x)) + ((ax41x) & (bx41x) & (!g86) & (g88) & (!ax42x) & (!bx42x)) + ((ax41x) & (bx41x) & (g86) & (!g88) & (!ax42x) & (!bx42x)) + ((ax41x) & (bx41x) & (g86) & (g88) & (!ax42x) & (!bx42x)));
	assign fx43x = (((!ax43x) & (!bx43x) & (!g92)) + ((!ax43x) & (bx43x) & (g92)) + ((ax43x) & (!bx43x) & (g92)) + ((ax43x) & (bx43x) & (!g92)));
	assign g94 = (((!ax43x) & (bx43x) & (!g92)) + ((ax43x) & (!bx43x) & (!g92)) + ((ax43x) & (bx43x) & (!g92)) + ((ax43x) & (bx43x) & (g92)));
	assign fx44x = (((!ax44x) & (!bx44x) & (g94)) + ((!ax44x) & (bx44x) & (!g94)) + ((ax44x) & (!bx44x) & (!g94)) + ((ax44x) & (bx44x) & (g94)));
	assign fx45x = (((!ax44x) & (!bx44x) & (!g94) & (!ax45x) & (bx45x)) + ((!ax44x) & (!bx44x) & (!g94) & (ax45x) & (!bx45x)) + ((!ax44x) & (!bx44x) & (g94) & (!ax45x) & (bx45x)) + ((!ax44x) & (!bx44x) & (g94) & (ax45x) & (!bx45x)) + ((!ax44x) & (bx44x) & (!g94) & (!ax45x) & (bx45x)) + ((!ax44x) & (bx44x) & (!g94) & (ax45x) & (!bx45x)) + ((!ax44x) & (bx44x) & (g94) & (!ax45x) & (!bx45x)) + ((!ax44x) & (bx44x) & (g94) & (ax45x) & (bx45x)) + ((ax44x) & (!bx44x) & (!g94) & (!ax45x) & (bx45x)) + ((ax44x) & (!bx44x) & (!g94) & (ax45x) & (!bx45x)) + ((ax44x) & (!bx44x) & (g94) & (!ax45x) & (!bx45x)) + ((ax44x) & (!bx44x) & (g94) & (ax45x) & (bx45x)) + ((ax44x) & (bx44x) & (!g94) & (!ax45x) & (!bx45x)) + ((ax44x) & (bx44x) & (!g94) & (ax45x) & (bx45x)) + ((ax44x) & (bx44x) & (g94) & (!ax45x) & (!bx45x)) + ((ax44x) & (bx44x) & (g94) & (ax45x) & (bx45x)));
	assign g97 = (((ax45x) & (bx45x)));
	assign g98 = (((!ax45x) & (!bx45x)));
	assign g99 = (((!ax43x) & (!bx43x) & (!g92) & (ax44x) & (bx44x) & (!g98)) + ((!ax43x) & (!bx43x) & (g92) & (ax44x) & (bx44x) & (!g98)) + ((!ax43x) & (bx43x) & (!g92) & (!ax44x) & (bx44x) & (!g98)) + ((!ax43x) & (bx43x) & (!g92) & (ax44x) & (!bx44x) & (!g98)) + ((!ax43x) & (bx43x) & (!g92) & (ax44x) & (bx44x) & (!g98)) + ((!ax43x) & (bx43x) & (g92) & (ax44x) & (bx44x) & (!g98)) + ((ax43x) & (!bx43x) & (!g92) & (!ax44x) & (bx44x) & (!g98)) + ((ax43x) & (!bx43x) & (!g92) & (ax44x) & (!bx44x) & (!g98)) + ((ax43x) & (!bx43x) & (!g92) & (ax44x) & (bx44x) & (!g98)) + ((ax43x) & (!bx43x) & (g92) & (ax44x) & (bx44x) & (!g98)) + ((ax43x) & (bx43x) & (!g92) & (!ax44x) & (bx44x) & (!g98)) + ((ax43x) & (bx43x) & (!g92) & (ax44x) & (!bx44x) & (!g98)) + ((ax43x) & (bx43x) & (!g92) & (ax44x) & (bx44x) & (!g98)) + ((ax43x) & (bx43x) & (g92) & (!ax44x) & (bx44x) & (!g98)) + ((ax43x) & (bx43x) & (g92) & (ax44x) & (!bx44x) & (!g98)) + ((ax43x) & (bx43x) & (g92) & (ax44x) & (bx44x) & (!g98)));
	assign g100 = (((!g97) & (!g99)));
	assign fx46x = (((!ax46x) & (!bx46x) & (!g100)) + ((!ax46x) & (bx46x) & (g100)) + ((ax46x) & (!bx46x) & (g100)) + ((ax46x) & (bx46x) & (!g100)));
	assign fx47x = (((!ax46x) & (!bx46x) & (!g100) & (!ax47x) & (bx47x)) + ((!ax46x) & (!bx46x) & (!g100) & (ax47x) & (!bx47x)) + ((!ax46x) & (!bx46x) & (g100) & (!ax47x) & (bx47x)) + ((!ax46x) & (!bx46x) & (g100) & (ax47x) & (!bx47x)) + ((!ax46x) & (bx46x) & (!g100) & (!ax47x) & (!bx47x)) + ((!ax46x) & (bx46x) & (!g100) & (ax47x) & (bx47x)) + ((!ax46x) & (bx46x) & (g100) & (!ax47x) & (bx47x)) + ((!ax46x) & (bx46x) & (g100) & (ax47x) & (!bx47x)) + ((ax46x) & (!bx46x) & (!g100) & (!ax47x) & (!bx47x)) + ((ax46x) & (!bx46x) & (!g100) & (ax47x) & (bx47x)) + ((ax46x) & (!bx46x) & (g100) & (!ax47x) & (bx47x)) + ((ax46x) & (!bx46x) & (g100) & (ax47x) & (!bx47x)) + ((ax46x) & (bx46x) & (!g100) & (!ax47x) & (!bx47x)) + ((ax46x) & (bx46x) & (!g100) & (ax47x) & (bx47x)) + ((ax46x) & (bx46x) & (g100) & (!ax47x) & (!bx47x)) + ((ax46x) & (bx46x) & (g100) & (ax47x) & (bx47x)));
	assign g103 = (((!ax46x) & (!bx46x) & (!g97) & (!g99) & (!ax47x) & (!bx47x)) + ((!ax46x) & (!bx46x) & (!g97) & (!g99) & (!ax47x) & (bx47x)) + ((!ax46x) & (!bx46x) & (!g97) & (!g99) & (ax47x) & (!bx47x)) + ((!ax46x) & (!bx46x) & (!g97) & (g99) & (!ax47x) & (!bx47x)) + ((!ax46x) & (!bx46x) & (!g97) & (g99) & (!ax47x) & (bx47x)) + ((!ax46x) & (!bx46x) & (!g97) & (g99) & (ax47x) & (!bx47x)) + ((!ax46x) & (!bx46x) & (g97) & (!g99) & (!ax47x) & (!bx47x)) + ((!ax46x) & (!bx46x) & (g97) & (!g99) & (!ax47x) & (bx47x)) + ((!ax46x) & (!bx46x) & (g97) & (!g99) & (ax47x) & (!bx47x)) + ((!ax46x) & (!bx46x) & (g97) & (g99) & (!ax47x) & (!bx47x)) + ((!ax46x) & (!bx46x) & (g97) & (g99) & (!ax47x) & (bx47x)) + ((!ax46x) & (!bx46x) & (g97) & (g99) & (ax47x) & (!bx47x)) + ((!ax46x) & (bx46x) & (!g97) & (!g99) & (!ax47x) & (!bx47x)) + ((!ax46x) & (bx46x) & (!g97) & (!g99) & (!ax47x) & (bx47x)) + ((!ax46x) & (bx46x) & (!g97) & (!g99) & (ax47x) & (!bx47x)) + ((!ax46x) & (bx46x) & (!g97) & (g99) & (!ax47x) & (!bx47x)) + ((!ax46x) & (bx46x) & (g97) & (!g99) & (!ax47x) & (!bx47x)) + ((!ax46x) & (bx46x) & (g97) & (g99) & (!ax47x) & (!bx47x)) + ((ax46x) & (!bx46x) & (!g97) & (!g99) & (!ax47x) & (!bx47x)) + ((ax46x) & (!bx46x) & (!g97) & (!g99) & (!ax47x) & (bx47x)) + ((ax46x) & (!bx46x) & (!g97) & (!g99) & (ax47x) & (!bx47x)) + ((ax46x) & (!bx46x) & (!g97) & (g99) & (!ax47x) & (!bx47x)) + ((ax46x) & (!bx46x) & (g97) & (!g99) & (!ax47x) & (!bx47x)) + ((ax46x) & (!bx46x) & (g97) & (g99) & (!ax47x) & (!bx47x)) + ((ax46x) & (bx46x) & (!g97) & (!g99) & (!ax47x) & (!bx47x)) + ((ax46x) & (bx46x) & (!g97) & (g99) & (!ax47x) & (!bx47x)) + ((ax46x) & (bx46x) & (g97) & (!g99) & (!ax47x) & (!bx47x)) + ((ax46x) & (bx46x) & (g97) & (g99) & (!ax47x) & (!bx47x)));
	assign fx48x = (((!ax48x) & (!bx48x) & (!g103)) + ((!ax48x) & (bx48x) & (g103)) + ((ax48x) & (!bx48x) & (g103)) + ((ax48x) & (bx48x) & (!g103)));
	assign g105 = (((!ax48x) & (bx48x) & (!g103)) + ((ax48x) & (!bx48x) & (!g103)) + ((ax48x) & (bx48x) & (!g103)) + ((ax48x) & (bx48x) & (g103)));
	assign fx49x = (((!ax49x) & (!bx49x) & (g105)) + ((!ax49x) & (bx49x) & (!g105)) + ((ax49x) & (!bx49x) & (!g105)) + ((ax49x) & (bx49x) & (g105)));
	assign fx50x = (((!ax49x) & (!bx49x) & (!g105) & (!ax50x) & (bx50x)) + ((!ax49x) & (!bx49x) & (!g105) & (ax50x) & (!bx50x)) + ((!ax49x) & (!bx49x) & (g105) & (!ax50x) & (bx50x)) + ((!ax49x) & (!bx49x) & (g105) & (ax50x) & (!bx50x)) + ((!ax49x) & (bx49x) & (!g105) & (!ax50x) & (bx50x)) + ((!ax49x) & (bx49x) & (!g105) & (ax50x) & (!bx50x)) + ((!ax49x) & (bx49x) & (g105) & (!ax50x) & (!bx50x)) + ((!ax49x) & (bx49x) & (g105) & (ax50x) & (bx50x)) + ((ax49x) & (!bx49x) & (!g105) & (!ax50x) & (bx50x)) + ((ax49x) & (!bx49x) & (!g105) & (ax50x) & (!bx50x)) + ((ax49x) & (!bx49x) & (g105) & (!ax50x) & (!bx50x)) + ((ax49x) & (!bx49x) & (g105) & (ax50x) & (bx50x)) + ((ax49x) & (bx49x) & (!g105) & (!ax50x) & (!bx50x)) + ((ax49x) & (bx49x) & (!g105) & (ax50x) & (bx50x)) + ((ax49x) & (bx49x) & (g105) & (!ax50x) & (!bx50x)) + ((ax49x) & (bx49x) & (g105) & (ax50x) & (bx50x)));
	assign g108 = (((ax50x) & (bx50x)));
	assign g109 = (((!ax50x) & (!bx50x)));
	assign g110 = (((!ax48x) & (!bx48x) & (!g103) & (ax49x) & (bx49x) & (!g109)) + ((!ax48x) & (!bx48x) & (g103) & (ax49x) & (bx49x) & (!g109)) + ((!ax48x) & (bx48x) & (!g103) & (!ax49x) & (bx49x) & (!g109)) + ((!ax48x) & (bx48x) & (!g103) & (ax49x) & (!bx49x) & (!g109)) + ((!ax48x) & (bx48x) & (!g103) & (ax49x) & (bx49x) & (!g109)) + ((!ax48x) & (bx48x) & (g103) & (ax49x) & (bx49x) & (!g109)) + ((ax48x) & (!bx48x) & (!g103) & (!ax49x) & (bx49x) & (!g109)) + ((ax48x) & (!bx48x) & (!g103) & (ax49x) & (!bx49x) & (!g109)) + ((ax48x) & (!bx48x) & (!g103) & (ax49x) & (bx49x) & (!g109)) + ((ax48x) & (!bx48x) & (g103) & (ax49x) & (bx49x) & (!g109)) + ((ax48x) & (bx48x) & (!g103) & (!ax49x) & (bx49x) & (!g109)) + ((ax48x) & (bx48x) & (!g103) & (ax49x) & (!bx49x) & (!g109)) + ((ax48x) & (bx48x) & (!g103) & (ax49x) & (bx49x) & (!g109)) + ((ax48x) & (bx48x) & (g103) & (!ax49x) & (bx49x) & (!g109)) + ((ax48x) & (bx48x) & (g103) & (ax49x) & (!bx49x) & (!g109)) + ((ax48x) & (bx48x) & (g103) & (ax49x) & (bx49x) & (!g109)));
	assign fx51x = (((!ax51x) & (!bx51x) & (!g108) & (g110)) + ((!ax51x) & (!bx51x) & (g108) & (!g110)) + ((!ax51x) & (!bx51x) & (g108) & (g110)) + ((!ax51x) & (bx51x) & (!g108) & (!g110)) + ((ax51x) & (!bx51x) & (!g108) & (!g110)) + ((ax51x) & (bx51x) & (!g108) & (g110)) + ((ax51x) & (bx51x) & (g108) & (!g110)) + ((ax51x) & (bx51x) & (g108) & (g110)));
	assign fx52x = (((!ax51x) & (!bx51x) & (!g108) & (!g110) & (!ax52x) & (bx52x)) + ((!ax51x) & (!bx51x) & (!g108) & (!g110) & (ax52x) & (!bx52x)) + ((!ax51x) & (!bx51x) & (!g108) & (g110) & (!ax52x) & (bx52x)) + ((!ax51x) & (!bx51x) & (!g108) & (g110) & (ax52x) & (!bx52x)) + ((!ax51x) & (!bx51x) & (g108) & (!g110) & (!ax52x) & (bx52x)) + ((!ax51x) & (!bx51x) & (g108) & (!g110) & (ax52x) & (!bx52x)) + ((!ax51x) & (!bx51x) & (g108) & (g110) & (!ax52x) & (bx52x)) + ((!ax51x) & (!bx51x) & (g108) & (g110) & (ax52x) & (!bx52x)) + ((!ax51x) & (bx51x) & (!g108) & (!g110) & (!ax52x) & (bx52x)) + ((!ax51x) & (bx51x) & (!g108) & (!g110) & (ax52x) & (!bx52x)) + ((!ax51x) & (bx51x) & (!g108) & (g110) & (!ax52x) & (!bx52x)) + ((!ax51x) & (bx51x) & (!g108) & (g110) & (ax52x) & (bx52x)) + ((!ax51x) & (bx51x) & (g108) & (!g110) & (!ax52x) & (!bx52x)) + ((!ax51x) & (bx51x) & (g108) & (!g110) & (ax52x) & (bx52x)) + ((!ax51x) & (bx51x) & (g108) & (g110) & (!ax52x) & (!bx52x)) + ((!ax51x) & (bx51x) & (g108) & (g110) & (ax52x) & (bx52x)) + ((ax51x) & (!bx51x) & (!g108) & (!g110) & (!ax52x) & (bx52x)) + ((ax51x) & (!bx51x) & (!g108) & (!g110) & (ax52x) & (!bx52x)) + ((ax51x) & (!bx51x) & (!g108) & (g110) & (!ax52x) & (!bx52x)) + ((ax51x) & (!bx51x) & (!g108) & (g110) & (ax52x) & (bx52x)) + ((ax51x) & (!bx51x) & (g108) & (!g110) & (!ax52x) & (!bx52x)) + ((ax51x) & (!bx51x) & (g108) & (!g110) & (ax52x) & (bx52x)) + ((ax51x) & (!bx51x) & (g108) & (g110) & (!ax52x) & (!bx52x)) + ((ax51x) & (!bx51x) & (g108) & (g110) & (ax52x) & (bx52x)) + ((ax51x) & (bx51x) & (!g108) & (!g110) & (!ax52x) & (!bx52x)) + ((ax51x) & (bx51x) & (!g108) & (!g110) & (ax52x) & (bx52x)) + ((ax51x) & (bx51x) & (!g108) & (g110) & (!ax52x) & (!bx52x)) + ((ax51x) & (bx51x) & (!g108) & (g110) & (ax52x) & (bx52x)) + ((ax51x) & (bx51x) & (g108) & (!g110) & (!ax52x) & (!bx52x)) + ((ax51x) & (bx51x) & (g108) & (!g110) & (ax52x) & (bx52x)) + ((ax51x) & (bx51x) & (g108) & (g110) & (!ax52x) & (!bx52x)) + ((ax51x) & (bx51x) & (g108) & (g110) & (ax52x) & (bx52x)));
	assign g113 = (((!ax51x) & (!bx51x) & (!g108) & (!g110) & (!ax52x) & (!bx52x)) + ((!ax51x) & (!bx51x) & (!g108) & (!g110) & (!ax52x) & (bx52x)) + ((!ax51x) & (!bx51x) & (!g108) & (!g110) & (ax52x) & (!bx52x)) + ((!ax51x) & (!bx51x) & (!g108) & (g110) & (!ax52x) & (!bx52x)) + ((!ax51x) & (!bx51x) & (!g108) & (g110) & (!ax52x) & (bx52x)) + ((!ax51x) & (!bx51x) & (!g108) & (g110) & (ax52x) & (!bx52x)) + ((!ax51x) & (!bx51x) & (g108) & (!g110) & (!ax52x) & (!bx52x)) + ((!ax51x) & (!bx51x) & (g108) & (!g110) & (!ax52x) & (bx52x)) + ((!ax51x) & (!bx51x) & (g108) & (!g110) & (ax52x) & (!bx52x)) + ((!ax51x) & (!bx51x) & (g108) & (g110) & (!ax52x) & (!bx52x)) + ((!ax51x) & (!bx51x) & (g108) & (g110) & (!ax52x) & (bx52x)) + ((!ax51x) & (!bx51x) & (g108) & (g110) & (ax52x) & (!bx52x)) + ((!ax51x) & (bx51x) & (!g108) & (!g110) & (!ax52x) & (!bx52x)) + ((!ax51x) & (bx51x) & (!g108) & (!g110) & (!ax52x) & (bx52x)) + ((!ax51x) & (bx51x) & (!g108) & (!g110) & (ax52x) & (!bx52x)) + ((!ax51x) & (bx51x) & (!g108) & (g110) & (!ax52x) & (!bx52x)) + ((!ax51x) & (bx51x) & (g108) & (!g110) & (!ax52x) & (!bx52x)) + ((!ax51x) & (bx51x) & (g108) & (g110) & (!ax52x) & (!bx52x)) + ((ax51x) & (!bx51x) & (!g108) & (!g110) & (!ax52x) & (!bx52x)) + ((ax51x) & (!bx51x) & (!g108) & (!g110) & (!ax52x) & (bx52x)) + ((ax51x) & (!bx51x) & (!g108) & (!g110) & (ax52x) & (!bx52x)) + ((ax51x) & (!bx51x) & (!g108) & (g110) & (!ax52x) & (!bx52x)) + ((ax51x) & (!bx51x) & (g108) & (!g110) & (!ax52x) & (!bx52x)) + ((ax51x) & (!bx51x) & (g108) & (g110) & (!ax52x) & (!bx52x)) + ((ax51x) & (bx51x) & (!g108) & (!g110) & (!ax52x) & (!bx52x)) + ((ax51x) & (bx51x) & (!g108) & (g110) & (!ax52x) & (!bx52x)) + ((ax51x) & (bx51x) & (g108) & (!g110) & (!ax52x) & (!bx52x)) + ((ax51x) & (bx51x) & (g108) & (g110) & (!ax52x) & (!bx52x)));
	assign fx53x = (((!ax53x) & (!bx53x) & (!g113)) + ((!ax53x) & (bx53x) & (g113)) + ((ax53x) & (!bx53x) & (g113)) + ((ax53x) & (bx53x) & (!g113)));
	assign g115 = (((!ax53x) & (bx53x) & (!g113)) + ((ax53x) & (!bx53x) & (!g113)) + ((ax53x) & (bx53x) & (!g113)) + ((ax53x) & (bx53x) & (g113)));
	assign fx54x = (((!ax54x) & (!bx54x) & (g115)) + ((!ax54x) & (bx54x) & (!g115)) + ((ax54x) & (!bx54x) & (!g115)) + ((ax54x) & (bx54x) & (g115)));
	assign fx55x = (((!ax54x) & (!bx54x) & (!g115) & (!ax55x) & (bx55x)) + ((!ax54x) & (!bx54x) & (!g115) & (ax55x) & (!bx55x)) + ((!ax54x) & (!bx54x) & (g115) & (!ax55x) & (bx55x)) + ((!ax54x) & (!bx54x) & (g115) & (ax55x) & (!bx55x)) + ((!ax54x) & (bx54x) & (!g115) & (!ax55x) & (bx55x)) + ((!ax54x) & (bx54x) & (!g115) & (ax55x) & (!bx55x)) + ((!ax54x) & (bx54x) & (g115) & (!ax55x) & (!bx55x)) + ((!ax54x) & (bx54x) & (g115) & (ax55x) & (bx55x)) + ((ax54x) & (!bx54x) & (!g115) & (!ax55x) & (bx55x)) + ((ax54x) & (!bx54x) & (!g115) & (ax55x) & (!bx55x)) + ((ax54x) & (!bx54x) & (g115) & (!ax55x) & (!bx55x)) + ((ax54x) & (!bx54x) & (g115) & (ax55x) & (bx55x)) + ((ax54x) & (bx54x) & (!g115) & (!ax55x) & (!bx55x)) + ((ax54x) & (bx54x) & (!g115) & (ax55x) & (bx55x)) + ((ax54x) & (bx54x) & (g115) & (!ax55x) & (!bx55x)) + ((ax54x) & (bx54x) & (g115) & (ax55x) & (bx55x)));
	assign g118 = (((ax55x) & (bx55x)));
	assign g119 = (((!ax55x) & (!bx55x)));
	assign g120 = (((!ax53x) & (!bx53x) & (!g113) & (ax54x) & (bx54x) & (!g119)) + ((!ax53x) & (!bx53x) & (g113) & (ax54x) & (bx54x) & (!g119)) + ((!ax53x) & (bx53x) & (!g113) & (!ax54x) & (bx54x) & (!g119)) + ((!ax53x) & (bx53x) & (!g113) & (ax54x) & (!bx54x) & (!g119)) + ((!ax53x) & (bx53x) & (!g113) & (ax54x) & (bx54x) & (!g119)) + ((!ax53x) & (bx53x) & (g113) & (ax54x) & (bx54x) & (!g119)) + ((ax53x) & (!bx53x) & (!g113) & (!ax54x) & (bx54x) & (!g119)) + ((ax53x) & (!bx53x) & (!g113) & (ax54x) & (!bx54x) & (!g119)) + ((ax53x) & (!bx53x) & (!g113) & (ax54x) & (bx54x) & (!g119)) + ((ax53x) & (!bx53x) & (g113) & (ax54x) & (bx54x) & (!g119)) + ((ax53x) & (bx53x) & (!g113) & (!ax54x) & (bx54x) & (!g119)) + ((ax53x) & (bx53x) & (!g113) & (ax54x) & (!bx54x) & (!g119)) + ((ax53x) & (bx53x) & (!g113) & (ax54x) & (bx54x) & (!g119)) + ((ax53x) & (bx53x) & (g113) & (!ax54x) & (bx54x) & (!g119)) + ((ax53x) & (bx53x) & (g113) & (ax54x) & (!bx54x) & (!g119)) + ((ax53x) & (bx53x) & (g113) & (ax54x) & (bx54x) & (!g119)));
	assign g121 = (((!g118) & (!g120)));
	assign fx56x = (((!ax56x) & (!bx56x) & (!g121)) + ((!ax56x) & (bx56x) & (g121)) + ((ax56x) & (!bx56x) & (g121)) + ((ax56x) & (bx56x) & (!g121)));
	assign fx57x = (((!ax56x) & (!bx56x) & (!g121) & (!ax57x) & (bx57x)) + ((!ax56x) & (!bx56x) & (!g121) & (ax57x) & (!bx57x)) + ((!ax56x) & (!bx56x) & (g121) & (!ax57x) & (bx57x)) + ((!ax56x) & (!bx56x) & (g121) & (ax57x) & (!bx57x)) + ((!ax56x) & (bx56x) & (!g121) & (!ax57x) & (!bx57x)) + ((!ax56x) & (bx56x) & (!g121) & (ax57x) & (bx57x)) + ((!ax56x) & (bx56x) & (g121) & (!ax57x) & (bx57x)) + ((!ax56x) & (bx56x) & (g121) & (ax57x) & (!bx57x)) + ((ax56x) & (!bx56x) & (!g121) & (!ax57x) & (!bx57x)) + ((ax56x) & (!bx56x) & (!g121) & (ax57x) & (bx57x)) + ((ax56x) & (!bx56x) & (g121) & (!ax57x) & (bx57x)) + ((ax56x) & (!bx56x) & (g121) & (ax57x) & (!bx57x)) + ((ax56x) & (bx56x) & (!g121) & (!ax57x) & (!bx57x)) + ((ax56x) & (bx56x) & (!g121) & (ax57x) & (bx57x)) + ((ax56x) & (bx56x) & (g121) & (!ax57x) & (!bx57x)) + ((ax56x) & (bx56x) & (g121) & (ax57x) & (bx57x)));
	assign g124 = (((!ax56x) & (!bx56x) & (!g118) & (!g120) & (!ax57x) & (!bx57x)) + ((!ax56x) & (!bx56x) & (!g118) & (!g120) & (!ax57x) & (bx57x)) + ((!ax56x) & (!bx56x) & (!g118) & (!g120) & (ax57x) & (!bx57x)) + ((!ax56x) & (!bx56x) & (!g118) & (g120) & (!ax57x) & (!bx57x)) + ((!ax56x) & (!bx56x) & (!g118) & (g120) & (!ax57x) & (bx57x)) + ((!ax56x) & (!bx56x) & (!g118) & (g120) & (ax57x) & (!bx57x)) + ((!ax56x) & (!bx56x) & (g118) & (!g120) & (!ax57x) & (!bx57x)) + ((!ax56x) & (!bx56x) & (g118) & (!g120) & (!ax57x) & (bx57x)) + ((!ax56x) & (!bx56x) & (g118) & (!g120) & (ax57x) & (!bx57x)) + ((!ax56x) & (!bx56x) & (g118) & (g120) & (!ax57x) & (!bx57x)) + ((!ax56x) & (!bx56x) & (g118) & (g120) & (!ax57x) & (bx57x)) + ((!ax56x) & (!bx56x) & (g118) & (g120) & (ax57x) & (!bx57x)) + ((!ax56x) & (bx56x) & (!g118) & (!g120) & (!ax57x) & (!bx57x)) + ((!ax56x) & (bx56x) & (!g118) & (!g120) & (!ax57x) & (bx57x)) + ((!ax56x) & (bx56x) & (!g118) & (!g120) & (ax57x) & (!bx57x)) + ((!ax56x) & (bx56x) & (!g118) & (g120) & (!ax57x) & (!bx57x)) + ((!ax56x) & (bx56x) & (g118) & (!g120) & (!ax57x) & (!bx57x)) + ((!ax56x) & (bx56x) & (g118) & (g120) & (!ax57x) & (!bx57x)) + ((ax56x) & (!bx56x) & (!g118) & (!g120) & (!ax57x) & (!bx57x)) + ((ax56x) & (!bx56x) & (!g118) & (!g120) & (!ax57x) & (bx57x)) + ((ax56x) & (!bx56x) & (!g118) & (!g120) & (ax57x) & (!bx57x)) + ((ax56x) & (!bx56x) & (!g118) & (g120) & (!ax57x) & (!bx57x)) + ((ax56x) & (!bx56x) & (g118) & (!g120) & (!ax57x) & (!bx57x)) + ((ax56x) & (!bx56x) & (g118) & (g120) & (!ax57x) & (!bx57x)) + ((ax56x) & (bx56x) & (!g118) & (!g120) & (!ax57x) & (!bx57x)) + ((ax56x) & (bx56x) & (!g118) & (g120) & (!ax57x) & (!bx57x)) + ((ax56x) & (bx56x) & (g118) & (!g120) & (!ax57x) & (!bx57x)) + ((ax56x) & (bx56x) & (g118) & (g120) & (!ax57x) & (!bx57x)));
	assign fx58x = (((!ax58x) & (!bx58x) & (!g124)) + ((!ax58x) & (bx58x) & (g124)) + ((ax58x) & (!bx58x) & (g124)) + ((ax58x) & (bx58x) & (!g124)));
	assign g126 = (((!ax58x) & (bx58x) & (!g124)) + ((ax58x) & (!bx58x) & (!g124)) + ((ax58x) & (bx58x) & (!g124)) + ((ax58x) & (bx58x) & (g124)));
	assign fx59x = (((!ax59x) & (!bx59x) & (g126)) + ((!ax59x) & (bx59x) & (!g126)) + ((ax59x) & (!bx59x) & (!g126)) + ((ax59x) & (bx59x) & (g126)));
	assign fx60x = (((!ax59x) & (!bx59x) & (!g126) & (!ax60x) & (bx60x)) + ((!ax59x) & (!bx59x) & (!g126) & (ax60x) & (!bx60x)) + ((!ax59x) & (!bx59x) & (g126) & (!ax60x) & (bx60x)) + ((!ax59x) & (!bx59x) & (g126) & (ax60x) & (!bx60x)) + ((!ax59x) & (bx59x) & (!g126) & (!ax60x) & (bx60x)) + ((!ax59x) & (bx59x) & (!g126) & (ax60x) & (!bx60x)) + ((!ax59x) & (bx59x) & (g126) & (!ax60x) & (!bx60x)) + ((!ax59x) & (bx59x) & (g126) & (ax60x) & (bx60x)) + ((ax59x) & (!bx59x) & (!g126) & (!ax60x) & (bx60x)) + ((ax59x) & (!bx59x) & (!g126) & (ax60x) & (!bx60x)) + ((ax59x) & (!bx59x) & (g126) & (!ax60x) & (!bx60x)) + ((ax59x) & (!bx59x) & (g126) & (ax60x) & (bx60x)) + ((ax59x) & (bx59x) & (!g126) & (!ax60x) & (!bx60x)) + ((ax59x) & (bx59x) & (!g126) & (ax60x) & (bx60x)) + ((ax59x) & (bx59x) & (g126) & (!ax60x) & (!bx60x)) + ((ax59x) & (bx59x) & (g126) & (ax60x) & (bx60x)));
	assign g129 = (((ax60x) & (bx60x)));
	assign g130 = (((!ax60x) & (!bx60x)));
	assign g131 = (((!ax58x) & (!bx58x) & (!g124) & (ax59x) & (bx59x) & (!g130)) + ((!ax58x) & (!bx58x) & (g124) & (ax59x) & (bx59x) & (!g130)) + ((!ax58x) & (bx58x) & (!g124) & (!ax59x) & (bx59x) & (!g130)) + ((!ax58x) & (bx58x) & (!g124) & (ax59x) & (!bx59x) & (!g130)) + ((!ax58x) & (bx58x) & (!g124) & (ax59x) & (bx59x) & (!g130)) + ((!ax58x) & (bx58x) & (g124) & (ax59x) & (bx59x) & (!g130)) + ((ax58x) & (!bx58x) & (!g124) & (!ax59x) & (bx59x) & (!g130)) + ((ax58x) & (!bx58x) & (!g124) & (ax59x) & (!bx59x) & (!g130)) + ((ax58x) & (!bx58x) & (!g124) & (ax59x) & (bx59x) & (!g130)) + ((ax58x) & (!bx58x) & (g124) & (ax59x) & (bx59x) & (!g130)) + ((ax58x) & (bx58x) & (!g124) & (!ax59x) & (bx59x) & (!g130)) + ((ax58x) & (bx58x) & (!g124) & (ax59x) & (!bx59x) & (!g130)) + ((ax58x) & (bx58x) & (!g124) & (ax59x) & (bx59x) & (!g130)) + ((ax58x) & (bx58x) & (g124) & (!ax59x) & (bx59x) & (!g130)) + ((ax58x) & (bx58x) & (g124) & (ax59x) & (!bx59x) & (!g130)) + ((ax58x) & (bx58x) & (g124) & (ax59x) & (bx59x) & (!g130)));
	assign g132 = (((!g129) & (!g131)));
	assign fx61x = (((!ax61x) & (!bx61x) & (!g132)) + ((!ax61x) & (bx61x) & (g132)) + ((ax61x) & (!bx61x) & (g132)) + ((ax61x) & (bx61x) & (!g132)));
	assign fx62x = (((!ax61x) & (!bx61x) & (!g132) & (!ax62x) & (bx62x)) + ((!ax61x) & (!bx61x) & (!g132) & (ax62x) & (!bx62x)) + ((!ax61x) & (!bx61x) & (g132) & (!ax62x) & (bx62x)) + ((!ax61x) & (!bx61x) & (g132) & (ax62x) & (!bx62x)) + ((!ax61x) & (bx61x) & (!g132) & (!ax62x) & (!bx62x)) + ((!ax61x) & (bx61x) & (!g132) & (ax62x) & (bx62x)) + ((!ax61x) & (bx61x) & (g132) & (!ax62x) & (bx62x)) + ((!ax61x) & (bx61x) & (g132) & (ax62x) & (!bx62x)) + ((ax61x) & (!bx61x) & (!g132) & (!ax62x) & (!bx62x)) + ((ax61x) & (!bx61x) & (!g132) & (ax62x) & (bx62x)) + ((ax61x) & (!bx61x) & (g132) & (!ax62x) & (bx62x)) + ((ax61x) & (!bx61x) & (g132) & (ax62x) & (!bx62x)) + ((ax61x) & (bx61x) & (!g132) & (!ax62x) & (!bx62x)) + ((ax61x) & (bx61x) & (!g132) & (ax62x) & (bx62x)) + ((ax61x) & (bx61x) & (g132) & (!ax62x) & (!bx62x)) + ((ax61x) & (bx61x) & (g132) & (ax62x) & (bx62x)));
	assign g135 = (((!ax61x) & (!bx61x) & (!g129) & (!g131) & (!ax62x) & (!bx62x)) + ((!ax61x) & (!bx61x) & (!g129) & (!g131) & (!ax62x) & (bx62x)) + ((!ax61x) & (!bx61x) & (!g129) & (!g131) & (ax62x) & (!bx62x)) + ((!ax61x) & (!bx61x) & (!g129) & (g131) & (!ax62x) & (!bx62x)) + ((!ax61x) & (!bx61x) & (!g129) & (g131) & (!ax62x) & (bx62x)) + ((!ax61x) & (!bx61x) & (!g129) & (g131) & (ax62x) & (!bx62x)) + ((!ax61x) & (!bx61x) & (g129) & (!g131) & (!ax62x) & (!bx62x)) + ((!ax61x) & (!bx61x) & (g129) & (!g131) & (!ax62x) & (bx62x)) + ((!ax61x) & (!bx61x) & (g129) & (!g131) & (ax62x) & (!bx62x)) + ((!ax61x) & (!bx61x) & (g129) & (g131) & (!ax62x) & (!bx62x)) + ((!ax61x) & (!bx61x) & (g129) & (g131) & (!ax62x) & (bx62x)) + ((!ax61x) & (!bx61x) & (g129) & (g131) & (ax62x) & (!bx62x)) + ((!ax61x) & (bx61x) & (!g129) & (!g131) & (!ax62x) & (!bx62x)) + ((!ax61x) & (bx61x) & (!g129) & (!g131) & (!ax62x) & (bx62x)) + ((!ax61x) & (bx61x) & (!g129) & (!g131) & (ax62x) & (!bx62x)) + ((!ax61x) & (bx61x) & (!g129) & (g131) & (!ax62x) & (!bx62x)) + ((!ax61x) & (bx61x) & (g129) & (!g131) & (!ax62x) & (!bx62x)) + ((!ax61x) & (bx61x) & (g129) & (g131) & (!ax62x) & (!bx62x)) + ((ax61x) & (!bx61x) & (!g129) & (!g131) & (!ax62x) & (!bx62x)) + ((ax61x) & (!bx61x) & (!g129) & (!g131) & (!ax62x) & (bx62x)) + ((ax61x) & (!bx61x) & (!g129) & (!g131) & (ax62x) & (!bx62x)) + ((ax61x) & (!bx61x) & (!g129) & (g131) & (!ax62x) & (!bx62x)) + ((ax61x) & (!bx61x) & (g129) & (!g131) & (!ax62x) & (!bx62x)) + ((ax61x) & (!bx61x) & (g129) & (g131) & (!ax62x) & (!bx62x)) + ((ax61x) & (bx61x) & (!g129) & (!g131) & (!ax62x) & (!bx62x)) + ((ax61x) & (bx61x) & (!g129) & (g131) & (!ax62x) & (!bx62x)) + ((ax61x) & (bx61x) & (g129) & (!g131) & (!ax62x) & (!bx62x)) + ((ax61x) & (bx61x) & (g129) & (g131) & (!ax62x) & (!bx62x)));
	assign fx63x = (((!ax63x) & (!bx63x) & (!g135)) + ((!ax63x) & (bx63x) & (g135)) + ((ax63x) & (!bx63x) & (g135)) + ((ax63x) & (bx63x) & (!g135)));
	assign g137 = (((!ax63x) & (bx63x) & (!g135)) + ((ax63x) & (!bx63x) & (!g135)) + ((ax63x) & (bx63x) & (!g135)) + ((ax63x) & (bx63x) & (g135)));
	assign fx64x = (((!ax64x) & (!bx64x) & (g137)) + ((!ax64x) & (bx64x) & (!g137)) + ((ax64x) & (!bx64x) & (!g137)) + ((ax64x) & (bx64x) & (g137)));
	assign fx65x = (((!ax64x) & (!bx64x) & (!g137) & (!ax65x) & (bx65x)) + ((!ax64x) & (!bx64x) & (!g137) & (ax65x) & (!bx65x)) + ((!ax64x) & (!bx64x) & (g137) & (!ax65x) & (bx65x)) + ((!ax64x) & (!bx64x) & (g137) & (ax65x) & (!bx65x)) + ((!ax64x) & (bx64x) & (!g137) & (!ax65x) & (bx65x)) + ((!ax64x) & (bx64x) & (!g137) & (ax65x) & (!bx65x)) + ((!ax64x) & (bx64x) & (g137) & (!ax65x) & (!bx65x)) + ((!ax64x) & (bx64x) & (g137) & (ax65x) & (bx65x)) + ((ax64x) & (!bx64x) & (!g137) & (!ax65x) & (bx65x)) + ((ax64x) & (!bx64x) & (!g137) & (ax65x) & (!bx65x)) + ((ax64x) & (!bx64x) & (g137) & (!ax65x) & (!bx65x)) + ((ax64x) & (!bx64x) & (g137) & (ax65x) & (bx65x)) + ((ax64x) & (bx64x) & (!g137) & (!ax65x) & (!bx65x)) + ((ax64x) & (bx64x) & (!g137) & (ax65x) & (bx65x)) + ((ax64x) & (bx64x) & (g137) & (!ax65x) & (!bx65x)) + ((ax64x) & (bx64x) & (g137) & (ax65x) & (bx65x)));
	assign g140 = (((ax65x) & (bx65x)));
	assign g141 = (((!ax65x) & (!bx65x)));
	assign g142 = (((!ax63x) & (!bx63x) & (!g135) & (ax64x) & (bx64x) & (!g141)) + ((!ax63x) & (!bx63x) & (g135) & (ax64x) & (bx64x) & (!g141)) + ((!ax63x) & (bx63x) & (!g135) & (!ax64x) & (bx64x) & (!g141)) + ((!ax63x) & (bx63x) & (!g135) & (ax64x) & (!bx64x) & (!g141)) + ((!ax63x) & (bx63x) & (!g135) & (ax64x) & (bx64x) & (!g141)) + ((!ax63x) & (bx63x) & (g135) & (ax64x) & (bx64x) & (!g141)) + ((ax63x) & (!bx63x) & (!g135) & (!ax64x) & (bx64x) & (!g141)) + ((ax63x) & (!bx63x) & (!g135) & (ax64x) & (!bx64x) & (!g141)) + ((ax63x) & (!bx63x) & (!g135) & (ax64x) & (bx64x) & (!g141)) + ((ax63x) & (!bx63x) & (g135) & (ax64x) & (bx64x) & (!g141)) + ((ax63x) & (bx63x) & (!g135) & (!ax64x) & (bx64x) & (!g141)) + ((ax63x) & (bx63x) & (!g135) & (ax64x) & (!bx64x) & (!g141)) + ((ax63x) & (bx63x) & (!g135) & (ax64x) & (bx64x) & (!g141)) + ((ax63x) & (bx63x) & (g135) & (!ax64x) & (bx64x) & (!g141)) + ((ax63x) & (bx63x) & (g135) & (ax64x) & (!bx64x) & (!g141)) + ((ax63x) & (bx63x) & (g135) & (ax64x) & (bx64x) & (!g141)));
	assign g143 = (((!g140) & (!g142)));
	assign fx66x = (((!ax66x) & (!bx66x) & (!g143)) + ((!ax66x) & (bx66x) & (g143)) + ((ax66x) & (!bx66x) & (g143)) + ((ax66x) & (bx66x) & (!g143)));
	assign fx67x = (((!ax66x) & (!bx66x) & (!g143) & (!ax67x) & (bx67x)) + ((!ax66x) & (!bx66x) & (!g143) & (ax67x) & (!bx67x)) + ((!ax66x) & (!bx66x) & (g143) & (!ax67x) & (bx67x)) + ((!ax66x) & (!bx66x) & (g143) & (ax67x) & (!bx67x)) + ((!ax66x) & (bx66x) & (!g143) & (!ax67x) & (!bx67x)) + ((!ax66x) & (bx66x) & (!g143) & (ax67x) & (bx67x)) + ((!ax66x) & (bx66x) & (g143) & (!ax67x) & (bx67x)) + ((!ax66x) & (bx66x) & (g143) & (ax67x) & (!bx67x)) + ((ax66x) & (!bx66x) & (!g143) & (!ax67x) & (!bx67x)) + ((ax66x) & (!bx66x) & (!g143) & (ax67x) & (bx67x)) + ((ax66x) & (!bx66x) & (g143) & (!ax67x) & (bx67x)) + ((ax66x) & (!bx66x) & (g143) & (ax67x) & (!bx67x)) + ((ax66x) & (bx66x) & (!g143) & (!ax67x) & (!bx67x)) + ((ax66x) & (bx66x) & (!g143) & (ax67x) & (bx67x)) + ((ax66x) & (bx66x) & (g143) & (!ax67x) & (!bx67x)) + ((ax66x) & (bx66x) & (g143) & (ax67x) & (bx67x)));
	assign g146 = (((!ax66x) & (!bx66x) & (!g140) & (!g142) & (!ax67x) & (!bx67x)) + ((!ax66x) & (!bx66x) & (!g140) & (!g142) & (!ax67x) & (bx67x)) + ((!ax66x) & (!bx66x) & (!g140) & (!g142) & (ax67x) & (!bx67x)) + ((!ax66x) & (!bx66x) & (!g140) & (g142) & (!ax67x) & (!bx67x)) + ((!ax66x) & (!bx66x) & (!g140) & (g142) & (!ax67x) & (bx67x)) + ((!ax66x) & (!bx66x) & (!g140) & (g142) & (ax67x) & (!bx67x)) + ((!ax66x) & (!bx66x) & (g140) & (!g142) & (!ax67x) & (!bx67x)) + ((!ax66x) & (!bx66x) & (g140) & (!g142) & (!ax67x) & (bx67x)) + ((!ax66x) & (!bx66x) & (g140) & (!g142) & (ax67x) & (!bx67x)) + ((!ax66x) & (!bx66x) & (g140) & (g142) & (!ax67x) & (!bx67x)) + ((!ax66x) & (!bx66x) & (g140) & (g142) & (!ax67x) & (bx67x)) + ((!ax66x) & (!bx66x) & (g140) & (g142) & (ax67x) & (!bx67x)) + ((!ax66x) & (bx66x) & (!g140) & (!g142) & (!ax67x) & (!bx67x)) + ((!ax66x) & (bx66x) & (!g140) & (!g142) & (!ax67x) & (bx67x)) + ((!ax66x) & (bx66x) & (!g140) & (!g142) & (ax67x) & (!bx67x)) + ((!ax66x) & (bx66x) & (!g140) & (g142) & (!ax67x) & (!bx67x)) + ((!ax66x) & (bx66x) & (g140) & (!g142) & (!ax67x) & (!bx67x)) + ((!ax66x) & (bx66x) & (g140) & (g142) & (!ax67x) & (!bx67x)) + ((ax66x) & (!bx66x) & (!g140) & (!g142) & (!ax67x) & (!bx67x)) + ((ax66x) & (!bx66x) & (!g140) & (!g142) & (!ax67x) & (bx67x)) + ((ax66x) & (!bx66x) & (!g140) & (!g142) & (ax67x) & (!bx67x)) + ((ax66x) & (!bx66x) & (!g140) & (g142) & (!ax67x) & (!bx67x)) + ((ax66x) & (!bx66x) & (g140) & (!g142) & (!ax67x) & (!bx67x)) + ((ax66x) & (!bx66x) & (g140) & (g142) & (!ax67x) & (!bx67x)) + ((ax66x) & (bx66x) & (!g140) & (!g142) & (!ax67x) & (!bx67x)) + ((ax66x) & (bx66x) & (!g140) & (g142) & (!ax67x) & (!bx67x)) + ((ax66x) & (bx66x) & (g140) & (!g142) & (!ax67x) & (!bx67x)) + ((ax66x) & (bx66x) & (g140) & (g142) & (!ax67x) & (!bx67x)));
	assign fx68x = (((!ax68x) & (!bx68x) & (!g146)) + ((!ax68x) & (bx68x) & (g146)) + ((ax68x) & (!bx68x) & (g146)) + ((ax68x) & (bx68x) & (!g146)));
	assign g148 = (((!ax68x) & (bx68x) & (!g146)) + ((ax68x) & (!bx68x) & (!g146)) + ((ax68x) & (bx68x) & (!g146)) + ((ax68x) & (bx68x) & (g146)));
	assign fx69x = (((!ax69x) & (!bx69x) & (g148)) + ((!ax69x) & (bx69x) & (!g148)) + ((ax69x) & (!bx69x) & (!g148)) + ((ax69x) & (bx69x) & (g148)));
	assign fx70x = (((!ax69x) & (!bx69x) & (!g148) & (!ax70x) & (bx70x)) + ((!ax69x) & (!bx69x) & (!g148) & (ax70x) & (!bx70x)) + ((!ax69x) & (!bx69x) & (g148) & (!ax70x) & (bx70x)) + ((!ax69x) & (!bx69x) & (g148) & (ax70x) & (!bx70x)) + ((!ax69x) & (bx69x) & (!g148) & (!ax70x) & (bx70x)) + ((!ax69x) & (bx69x) & (!g148) & (ax70x) & (!bx70x)) + ((!ax69x) & (bx69x) & (g148) & (!ax70x) & (!bx70x)) + ((!ax69x) & (bx69x) & (g148) & (ax70x) & (bx70x)) + ((ax69x) & (!bx69x) & (!g148) & (!ax70x) & (bx70x)) + ((ax69x) & (!bx69x) & (!g148) & (ax70x) & (!bx70x)) + ((ax69x) & (!bx69x) & (g148) & (!ax70x) & (!bx70x)) + ((ax69x) & (!bx69x) & (g148) & (ax70x) & (bx70x)) + ((ax69x) & (bx69x) & (!g148) & (!ax70x) & (!bx70x)) + ((ax69x) & (bx69x) & (!g148) & (ax70x) & (bx70x)) + ((ax69x) & (bx69x) & (g148) & (!ax70x) & (!bx70x)) + ((ax69x) & (bx69x) & (g148) & (ax70x) & (bx70x)));
	assign g151 = (((ax70x) & (bx70x)));
	assign g152 = (((!ax70x) & (!bx70x)));
	assign g153 = (((!ax68x) & (!bx68x) & (!g146) & (ax69x) & (bx69x) & (!g152)) + ((!ax68x) & (!bx68x) & (g146) & (ax69x) & (bx69x) & (!g152)) + ((!ax68x) & (bx68x) & (!g146) & (!ax69x) & (bx69x) & (!g152)) + ((!ax68x) & (bx68x) & (!g146) & (ax69x) & (!bx69x) & (!g152)) + ((!ax68x) & (bx68x) & (!g146) & (ax69x) & (bx69x) & (!g152)) + ((!ax68x) & (bx68x) & (g146) & (ax69x) & (bx69x) & (!g152)) + ((ax68x) & (!bx68x) & (!g146) & (!ax69x) & (bx69x) & (!g152)) + ((ax68x) & (!bx68x) & (!g146) & (ax69x) & (!bx69x) & (!g152)) + ((ax68x) & (!bx68x) & (!g146) & (ax69x) & (bx69x) & (!g152)) + ((ax68x) & (!bx68x) & (g146) & (ax69x) & (bx69x) & (!g152)) + ((ax68x) & (bx68x) & (!g146) & (!ax69x) & (bx69x) & (!g152)) + ((ax68x) & (bx68x) & (!g146) & (ax69x) & (!bx69x) & (!g152)) + ((ax68x) & (bx68x) & (!g146) & (ax69x) & (bx69x) & (!g152)) + ((ax68x) & (bx68x) & (g146) & (!ax69x) & (bx69x) & (!g152)) + ((ax68x) & (bx68x) & (g146) & (ax69x) & (!bx69x) & (!g152)) + ((ax68x) & (bx68x) & (g146) & (ax69x) & (bx69x) & (!g152)));
	assign g154 = (((!g151) & (!g153)));
	assign fx71x = (((!ax71x) & (!bx71x) & (!g154)) + ((!ax71x) & (bx71x) & (g154)) + ((ax71x) & (!bx71x) & (g154)) + ((ax71x) & (bx71x) & (!g154)));
	assign fx72x = (((!ax71x) & (!bx71x) & (!g154) & (!ax72x) & (bx72x)) + ((!ax71x) & (!bx71x) & (!g154) & (ax72x) & (!bx72x)) + ((!ax71x) & (!bx71x) & (g154) & (!ax72x) & (bx72x)) + ((!ax71x) & (!bx71x) & (g154) & (ax72x) & (!bx72x)) + ((!ax71x) & (bx71x) & (!g154) & (!ax72x) & (!bx72x)) + ((!ax71x) & (bx71x) & (!g154) & (ax72x) & (bx72x)) + ((!ax71x) & (bx71x) & (g154) & (!ax72x) & (bx72x)) + ((!ax71x) & (bx71x) & (g154) & (ax72x) & (!bx72x)) + ((ax71x) & (!bx71x) & (!g154) & (!ax72x) & (!bx72x)) + ((ax71x) & (!bx71x) & (!g154) & (ax72x) & (bx72x)) + ((ax71x) & (!bx71x) & (g154) & (!ax72x) & (bx72x)) + ((ax71x) & (!bx71x) & (g154) & (ax72x) & (!bx72x)) + ((ax71x) & (bx71x) & (!g154) & (!ax72x) & (!bx72x)) + ((ax71x) & (bx71x) & (!g154) & (ax72x) & (bx72x)) + ((ax71x) & (bx71x) & (g154) & (!ax72x) & (!bx72x)) + ((ax71x) & (bx71x) & (g154) & (ax72x) & (bx72x)));
	assign g157 = (((!ax71x) & (!bx71x) & (!g151) & (!g153) & (!ax72x) & (!bx72x)) + ((!ax71x) & (!bx71x) & (!g151) & (!g153) & (!ax72x) & (bx72x)) + ((!ax71x) & (!bx71x) & (!g151) & (!g153) & (ax72x) & (!bx72x)) + ((!ax71x) & (!bx71x) & (!g151) & (g153) & (!ax72x) & (!bx72x)) + ((!ax71x) & (!bx71x) & (!g151) & (g153) & (!ax72x) & (bx72x)) + ((!ax71x) & (!bx71x) & (!g151) & (g153) & (ax72x) & (!bx72x)) + ((!ax71x) & (!bx71x) & (g151) & (!g153) & (!ax72x) & (!bx72x)) + ((!ax71x) & (!bx71x) & (g151) & (!g153) & (!ax72x) & (bx72x)) + ((!ax71x) & (!bx71x) & (g151) & (!g153) & (ax72x) & (!bx72x)) + ((!ax71x) & (!bx71x) & (g151) & (g153) & (!ax72x) & (!bx72x)) + ((!ax71x) & (!bx71x) & (g151) & (g153) & (!ax72x) & (bx72x)) + ((!ax71x) & (!bx71x) & (g151) & (g153) & (ax72x) & (!bx72x)) + ((!ax71x) & (bx71x) & (!g151) & (!g153) & (!ax72x) & (!bx72x)) + ((!ax71x) & (bx71x) & (!g151) & (!g153) & (!ax72x) & (bx72x)) + ((!ax71x) & (bx71x) & (!g151) & (!g153) & (ax72x) & (!bx72x)) + ((!ax71x) & (bx71x) & (!g151) & (g153) & (!ax72x) & (!bx72x)) + ((!ax71x) & (bx71x) & (g151) & (!g153) & (!ax72x) & (!bx72x)) + ((!ax71x) & (bx71x) & (g151) & (g153) & (!ax72x) & (!bx72x)) + ((ax71x) & (!bx71x) & (!g151) & (!g153) & (!ax72x) & (!bx72x)) + ((ax71x) & (!bx71x) & (!g151) & (!g153) & (!ax72x) & (bx72x)) + ((ax71x) & (!bx71x) & (!g151) & (!g153) & (ax72x) & (!bx72x)) + ((ax71x) & (!bx71x) & (!g151) & (g153) & (!ax72x) & (!bx72x)) + ((ax71x) & (!bx71x) & (g151) & (!g153) & (!ax72x) & (!bx72x)) + ((ax71x) & (!bx71x) & (g151) & (g153) & (!ax72x) & (!bx72x)) + ((ax71x) & (bx71x) & (!g151) & (!g153) & (!ax72x) & (!bx72x)) + ((ax71x) & (bx71x) & (!g151) & (g153) & (!ax72x) & (!bx72x)) + ((ax71x) & (bx71x) & (g151) & (!g153) & (!ax72x) & (!bx72x)) + ((ax71x) & (bx71x) & (g151) & (g153) & (!ax72x) & (!bx72x)));
	assign fx73x = (((!ax73x) & (!bx73x) & (!g157)) + ((!ax73x) & (bx73x) & (g157)) + ((ax73x) & (!bx73x) & (g157)) + ((ax73x) & (bx73x) & (!g157)));
	assign g159 = (((!ax73x) & (bx73x) & (!g157)) + ((ax73x) & (!bx73x) & (!g157)) + ((ax73x) & (bx73x) & (!g157)) + ((ax73x) & (bx73x) & (g157)));
	assign fx74x = (((!ax74x) & (!bx74x) & (g159)) + ((!ax74x) & (bx74x) & (!g159)) + ((ax74x) & (!bx74x) & (!g159)) + ((ax74x) & (bx74x) & (g159)));
	assign fx75x = (((!ax74x) & (!bx74x) & (!g159) & (!ax75x) & (bx75x)) + ((!ax74x) & (!bx74x) & (!g159) & (ax75x) & (!bx75x)) + ((!ax74x) & (!bx74x) & (g159) & (!ax75x) & (bx75x)) + ((!ax74x) & (!bx74x) & (g159) & (ax75x) & (!bx75x)) + ((!ax74x) & (bx74x) & (!g159) & (!ax75x) & (bx75x)) + ((!ax74x) & (bx74x) & (!g159) & (ax75x) & (!bx75x)) + ((!ax74x) & (bx74x) & (g159) & (!ax75x) & (!bx75x)) + ((!ax74x) & (bx74x) & (g159) & (ax75x) & (bx75x)) + ((ax74x) & (!bx74x) & (!g159) & (!ax75x) & (bx75x)) + ((ax74x) & (!bx74x) & (!g159) & (ax75x) & (!bx75x)) + ((ax74x) & (!bx74x) & (g159) & (!ax75x) & (!bx75x)) + ((ax74x) & (!bx74x) & (g159) & (ax75x) & (bx75x)) + ((ax74x) & (bx74x) & (!g159) & (!ax75x) & (!bx75x)) + ((ax74x) & (bx74x) & (!g159) & (ax75x) & (bx75x)) + ((ax74x) & (bx74x) & (g159) & (!ax75x) & (!bx75x)) + ((ax74x) & (bx74x) & (g159) & (ax75x) & (bx75x)));
	assign g162 = (((ax75x) & (bx75x)));
	assign g163 = (((!ax75x) & (!bx75x)));
	assign g164 = (((!ax73x) & (!bx73x) & (!g157) & (ax74x) & (bx74x) & (!g163)) + ((!ax73x) & (!bx73x) & (g157) & (ax74x) & (bx74x) & (!g163)) + ((!ax73x) & (bx73x) & (!g157) & (!ax74x) & (bx74x) & (!g163)) + ((!ax73x) & (bx73x) & (!g157) & (ax74x) & (!bx74x) & (!g163)) + ((!ax73x) & (bx73x) & (!g157) & (ax74x) & (bx74x) & (!g163)) + ((!ax73x) & (bx73x) & (g157) & (ax74x) & (bx74x) & (!g163)) + ((ax73x) & (!bx73x) & (!g157) & (!ax74x) & (bx74x) & (!g163)) + ((ax73x) & (!bx73x) & (!g157) & (ax74x) & (!bx74x) & (!g163)) + ((ax73x) & (!bx73x) & (!g157) & (ax74x) & (bx74x) & (!g163)) + ((ax73x) & (!bx73x) & (g157) & (ax74x) & (bx74x) & (!g163)) + ((ax73x) & (bx73x) & (!g157) & (!ax74x) & (bx74x) & (!g163)) + ((ax73x) & (bx73x) & (!g157) & (ax74x) & (!bx74x) & (!g163)) + ((ax73x) & (bx73x) & (!g157) & (ax74x) & (bx74x) & (!g163)) + ((ax73x) & (bx73x) & (g157) & (!ax74x) & (bx74x) & (!g163)) + ((ax73x) & (bx73x) & (g157) & (ax74x) & (!bx74x) & (!g163)) + ((ax73x) & (bx73x) & (g157) & (ax74x) & (bx74x) & (!g163)));
	assign g165 = (((!g162) & (!g164)));
	assign fx76x = (((!ax76x) & (!bx76x) & (!g165)) + ((!ax76x) & (bx76x) & (g165)) + ((ax76x) & (!bx76x) & (g165)) + ((ax76x) & (bx76x) & (!g165)));
	assign fx77x = (((!ax76x) & (!bx76x) & (!g165) & (!ax77x) & (bx77x)) + ((!ax76x) & (!bx76x) & (!g165) & (ax77x) & (!bx77x)) + ((!ax76x) & (!bx76x) & (g165) & (!ax77x) & (bx77x)) + ((!ax76x) & (!bx76x) & (g165) & (ax77x) & (!bx77x)) + ((!ax76x) & (bx76x) & (!g165) & (!ax77x) & (!bx77x)) + ((!ax76x) & (bx76x) & (!g165) & (ax77x) & (bx77x)) + ((!ax76x) & (bx76x) & (g165) & (!ax77x) & (bx77x)) + ((!ax76x) & (bx76x) & (g165) & (ax77x) & (!bx77x)) + ((ax76x) & (!bx76x) & (!g165) & (!ax77x) & (!bx77x)) + ((ax76x) & (!bx76x) & (!g165) & (ax77x) & (bx77x)) + ((ax76x) & (!bx76x) & (g165) & (!ax77x) & (bx77x)) + ((ax76x) & (!bx76x) & (g165) & (ax77x) & (!bx77x)) + ((ax76x) & (bx76x) & (!g165) & (!ax77x) & (!bx77x)) + ((ax76x) & (bx76x) & (!g165) & (ax77x) & (bx77x)) + ((ax76x) & (bx76x) & (g165) & (!ax77x) & (!bx77x)) + ((ax76x) & (bx76x) & (g165) & (ax77x) & (bx77x)));
	assign g168 = (((!ax76x) & (!bx76x) & (!g162) & (!g164) & (!ax77x) & (!bx77x)) + ((!ax76x) & (!bx76x) & (!g162) & (!g164) & (!ax77x) & (bx77x)) + ((!ax76x) & (!bx76x) & (!g162) & (!g164) & (ax77x) & (!bx77x)) + ((!ax76x) & (!bx76x) & (!g162) & (g164) & (!ax77x) & (!bx77x)) + ((!ax76x) & (!bx76x) & (!g162) & (g164) & (!ax77x) & (bx77x)) + ((!ax76x) & (!bx76x) & (!g162) & (g164) & (ax77x) & (!bx77x)) + ((!ax76x) & (!bx76x) & (g162) & (!g164) & (!ax77x) & (!bx77x)) + ((!ax76x) & (!bx76x) & (g162) & (!g164) & (!ax77x) & (bx77x)) + ((!ax76x) & (!bx76x) & (g162) & (!g164) & (ax77x) & (!bx77x)) + ((!ax76x) & (!bx76x) & (g162) & (g164) & (!ax77x) & (!bx77x)) + ((!ax76x) & (!bx76x) & (g162) & (g164) & (!ax77x) & (bx77x)) + ((!ax76x) & (!bx76x) & (g162) & (g164) & (ax77x) & (!bx77x)) + ((!ax76x) & (bx76x) & (!g162) & (!g164) & (!ax77x) & (!bx77x)) + ((!ax76x) & (bx76x) & (!g162) & (!g164) & (!ax77x) & (bx77x)) + ((!ax76x) & (bx76x) & (!g162) & (!g164) & (ax77x) & (!bx77x)) + ((!ax76x) & (bx76x) & (!g162) & (g164) & (!ax77x) & (!bx77x)) + ((!ax76x) & (bx76x) & (g162) & (!g164) & (!ax77x) & (!bx77x)) + ((!ax76x) & (bx76x) & (g162) & (g164) & (!ax77x) & (!bx77x)) + ((ax76x) & (!bx76x) & (!g162) & (!g164) & (!ax77x) & (!bx77x)) + ((ax76x) & (!bx76x) & (!g162) & (!g164) & (!ax77x) & (bx77x)) + ((ax76x) & (!bx76x) & (!g162) & (!g164) & (ax77x) & (!bx77x)) + ((ax76x) & (!bx76x) & (!g162) & (g164) & (!ax77x) & (!bx77x)) + ((ax76x) & (!bx76x) & (g162) & (!g164) & (!ax77x) & (!bx77x)) + ((ax76x) & (!bx76x) & (g162) & (g164) & (!ax77x) & (!bx77x)) + ((ax76x) & (bx76x) & (!g162) & (!g164) & (!ax77x) & (!bx77x)) + ((ax76x) & (bx76x) & (!g162) & (g164) & (!ax77x) & (!bx77x)) + ((ax76x) & (bx76x) & (g162) & (!g164) & (!ax77x) & (!bx77x)) + ((ax76x) & (bx76x) & (g162) & (g164) & (!ax77x) & (!bx77x)));
	assign fx78x = (((!ax78x) & (!bx78x) & (!g168)) + ((!ax78x) & (bx78x) & (g168)) + ((ax78x) & (!bx78x) & (g168)) + ((ax78x) & (bx78x) & (!g168)));
	assign g170 = (((!ax78x) & (bx78x) & (!g168)) + ((ax78x) & (!bx78x) & (!g168)) + ((ax78x) & (bx78x) & (!g168)) + ((ax78x) & (bx78x) & (g168)));
	assign fx79x = (((!ax79x) & (!bx79x) & (g170)) + ((!ax79x) & (bx79x) & (!g170)) + ((ax79x) & (!bx79x) & (!g170)) + ((ax79x) & (bx79x) & (g170)));
	assign fx80x = (((!ax79x) & (!bx79x) & (!g170) & (!ax80x) & (bx80x)) + ((!ax79x) & (!bx79x) & (!g170) & (ax80x) & (!bx80x)) + ((!ax79x) & (!bx79x) & (g170) & (!ax80x) & (bx80x)) + ((!ax79x) & (!bx79x) & (g170) & (ax80x) & (!bx80x)) + ((!ax79x) & (bx79x) & (!g170) & (!ax80x) & (bx80x)) + ((!ax79x) & (bx79x) & (!g170) & (ax80x) & (!bx80x)) + ((!ax79x) & (bx79x) & (g170) & (!ax80x) & (!bx80x)) + ((!ax79x) & (bx79x) & (g170) & (ax80x) & (bx80x)) + ((ax79x) & (!bx79x) & (!g170) & (!ax80x) & (bx80x)) + ((ax79x) & (!bx79x) & (!g170) & (ax80x) & (!bx80x)) + ((ax79x) & (!bx79x) & (g170) & (!ax80x) & (!bx80x)) + ((ax79x) & (!bx79x) & (g170) & (ax80x) & (bx80x)) + ((ax79x) & (bx79x) & (!g170) & (!ax80x) & (!bx80x)) + ((ax79x) & (bx79x) & (!g170) & (ax80x) & (bx80x)) + ((ax79x) & (bx79x) & (g170) & (!ax80x) & (!bx80x)) + ((ax79x) & (bx79x) & (g170) & (ax80x) & (bx80x)));
	assign g173 = (((ax80x) & (bx80x)));
	assign g174 = (((!ax80x) & (!bx80x)));
	assign g175 = (((!ax78x) & (!bx78x) & (!g168) & (ax79x) & (bx79x) & (!g174)) + ((!ax78x) & (!bx78x) & (g168) & (ax79x) & (bx79x) & (!g174)) + ((!ax78x) & (bx78x) & (!g168) & (!ax79x) & (bx79x) & (!g174)) + ((!ax78x) & (bx78x) & (!g168) & (ax79x) & (!bx79x) & (!g174)) + ((!ax78x) & (bx78x) & (!g168) & (ax79x) & (bx79x) & (!g174)) + ((!ax78x) & (bx78x) & (g168) & (ax79x) & (bx79x) & (!g174)) + ((ax78x) & (!bx78x) & (!g168) & (!ax79x) & (bx79x) & (!g174)) + ((ax78x) & (!bx78x) & (!g168) & (ax79x) & (!bx79x) & (!g174)) + ((ax78x) & (!bx78x) & (!g168) & (ax79x) & (bx79x) & (!g174)) + ((ax78x) & (!bx78x) & (g168) & (ax79x) & (bx79x) & (!g174)) + ((ax78x) & (bx78x) & (!g168) & (!ax79x) & (bx79x) & (!g174)) + ((ax78x) & (bx78x) & (!g168) & (ax79x) & (!bx79x) & (!g174)) + ((ax78x) & (bx78x) & (!g168) & (ax79x) & (bx79x) & (!g174)) + ((ax78x) & (bx78x) & (g168) & (!ax79x) & (bx79x) & (!g174)) + ((ax78x) & (bx78x) & (g168) & (ax79x) & (!bx79x) & (!g174)) + ((ax78x) & (bx78x) & (g168) & (ax79x) & (bx79x) & (!g174)));
	assign fx81x = (((!ax81x) & (!bx81x) & (!g173) & (g175)) + ((!ax81x) & (!bx81x) & (g173) & (!g175)) + ((!ax81x) & (!bx81x) & (g173) & (g175)) + ((!ax81x) & (bx81x) & (!g173) & (!g175)) + ((ax81x) & (!bx81x) & (!g173) & (!g175)) + ((ax81x) & (bx81x) & (!g173) & (g175)) + ((ax81x) & (bx81x) & (g173) & (!g175)) + ((ax81x) & (bx81x) & (g173) & (g175)));
	assign fx82x = (((!ax81x) & (!bx81x) & (!g173) & (!g175) & (!ax82x) & (bx82x)) + ((!ax81x) & (!bx81x) & (!g173) & (!g175) & (ax82x) & (!bx82x)) + ((!ax81x) & (!bx81x) & (!g173) & (g175) & (!ax82x) & (bx82x)) + ((!ax81x) & (!bx81x) & (!g173) & (g175) & (ax82x) & (!bx82x)) + ((!ax81x) & (!bx81x) & (g173) & (!g175) & (!ax82x) & (bx82x)) + ((!ax81x) & (!bx81x) & (g173) & (!g175) & (ax82x) & (!bx82x)) + ((!ax81x) & (!bx81x) & (g173) & (g175) & (!ax82x) & (bx82x)) + ((!ax81x) & (!bx81x) & (g173) & (g175) & (ax82x) & (!bx82x)) + ((!ax81x) & (bx81x) & (!g173) & (!g175) & (!ax82x) & (bx82x)) + ((!ax81x) & (bx81x) & (!g173) & (!g175) & (ax82x) & (!bx82x)) + ((!ax81x) & (bx81x) & (!g173) & (g175) & (!ax82x) & (!bx82x)) + ((!ax81x) & (bx81x) & (!g173) & (g175) & (ax82x) & (bx82x)) + ((!ax81x) & (bx81x) & (g173) & (!g175) & (!ax82x) & (!bx82x)) + ((!ax81x) & (bx81x) & (g173) & (!g175) & (ax82x) & (bx82x)) + ((!ax81x) & (bx81x) & (g173) & (g175) & (!ax82x) & (!bx82x)) + ((!ax81x) & (bx81x) & (g173) & (g175) & (ax82x) & (bx82x)) + ((ax81x) & (!bx81x) & (!g173) & (!g175) & (!ax82x) & (bx82x)) + ((ax81x) & (!bx81x) & (!g173) & (!g175) & (ax82x) & (!bx82x)) + ((ax81x) & (!bx81x) & (!g173) & (g175) & (!ax82x) & (!bx82x)) + ((ax81x) & (!bx81x) & (!g173) & (g175) & (ax82x) & (bx82x)) + ((ax81x) & (!bx81x) & (g173) & (!g175) & (!ax82x) & (!bx82x)) + ((ax81x) & (!bx81x) & (g173) & (!g175) & (ax82x) & (bx82x)) + ((ax81x) & (!bx81x) & (g173) & (g175) & (!ax82x) & (!bx82x)) + ((ax81x) & (!bx81x) & (g173) & (g175) & (ax82x) & (bx82x)) + ((ax81x) & (bx81x) & (!g173) & (!g175) & (!ax82x) & (!bx82x)) + ((ax81x) & (bx81x) & (!g173) & (!g175) & (ax82x) & (bx82x)) + ((ax81x) & (bx81x) & (!g173) & (g175) & (!ax82x) & (!bx82x)) + ((ax81x) & (bx81x) & (!g173) & (g175) & (ax82x) & (bx82x)) + ((ax81x) & (bx81x) & (g173) & (!g175) & (!ax82x) & (!bx82x)) + ((ax81x) & (bx81x) & (g173) & (!g175) & (ax82x) & (bx82x)) + ((ax81x) & (bx81x) & (g173) & (g175) & (!ax82x) & (!bx82x)) + ((ax81x) & (bx81x) & (g173) & (g175) & (ax82x) & (bx82x)));
	assign g178 = (((!ax81x) & (!bx81x) & (!g173) & (!g175) & (!ax82x) & (!bx82x)) + ((!ax81x) & (!bx81x) & (!g173) & (!g175) & (!ax82x) & (bx82x)) + ((!ax81x) & (!bx81x) & (!g173) & (!g175) & (ax82x) & (!bx82x)) + ((!ax81x) & (!bx81x) & (!g173) & (g175) & (!ax82x) & (!bx82x)) + ((!ax81x) & (!bx81x) & (!g173) & (g175) & (!ax82x) & (bx82x)) + ((!ax81x) & (!bx81x) & (!g173) & (g175) & (ax82x) & (!bx82x)) + ((!ax81x) & (!bx81x) & (g173) & (!g175) & (!ax82x) & (!bx82x)) + ((!ax81x) & (!bx81x) & (g173) & (!g175) & (!ax82x) & (bx82x)) + ((!ax81x) & (!bx81x) & (g173) & (!g175) & (ax82x) & (!bx82x)) + ((!ax81x) & (!bx81x) & (g173) & (g175) & (!ax82x) & (!bx82x)) + ((!ax81x) & (!bx81x) & (g173) & (g175) & (!ax82x) & (bx82x)) + ((!ax81x) & (!bx81x) & (g173) & (g175) & (ax82x) & (!bx82x)) + ((!ax81x) & (bx81x) & (!g173) & (!g175) & (!ax82x) & (!bx82x)) + ((!ax81x) & (bx81x) & (!g173) & (!g175) & (!ax82x) & (bx82x)) + ((!ax81x) & (bx81x) & (!g173) & (!g175) & (ax82x) & (!bx82x)) + ((!ax81x) & (bx81x) & (!g173) & (g175) & (!ax82x) & (!bx82x)) + ((!ax81x) & (bx81x) & (g173) & (!g175) & (!ax82x) & (!bx82x)) + ((!ax81x) & (bx81x) & (g173) & (g175) & (!ax82x) & (!bx82x)) + ((ax81x) & (!bx81x) & (!g173) & (!g175) & (!ax82x) & (!bx82x)) + ((ax81x) & (!bx81x) & (!g173) & (!g175) & (!ax82x) & (bx82x)) + ((ax81x) & (!bx81x) & (!g173) & (!g175) & (ax82x) & (!bx82x)) + ((ax81x) & (!bx81x) & (!g173) & (g175) & (!ax82x) & (!bx82x)) + ((ax81x) & (!bx81x) & (g173) & (!g175) & (!ax82x) & (!bx82x)) + ((ax81x) & (!bx81x) & (g173) & (g175) & (!ax82x) & (!bx82x)) + ((ax81x) & (bx81x) & (!g173) & (!g175) & (!ax82x) & (!bx82x)) + ((ax81x) & (bx81x) & (!g173) & (g175) & (!ax82x) & (!bx82x)) + ((ax81x) & (bx81x) & (g173) & (!g175) & (!ax82x) & (!bx82x)) + ((ax81x) & (bx81x) & (g173) & (g175) & (!ax82x) & (!bx82x)));
	assign fx83x = (((!ax83x) & (!bx83x) & (!g178)) + ((!ax83x) & (bx83x) & (g178)) + ((ax83x) & (!bx83x) & (g178)) + ((ax83x) & (bx83x) & (!g178)));
	assign g180 = (((!ax83x) & (bx83x) & (!g178)) + ((ax83x) & (!bx83x) & (!g178)) + ((ax83x) & (bx83x) & (!g178)) + ((ax83x) & (bx83x) & (g178)));
	assign fx84x = (((!ax84x) & (!bx84x) & (g180)) + ((!ax84x) & (bx84x) & (!g180)) + ((ax84x) & (!bx84x) & (!g180)) + ((ax84x) & (bx84x) & (g180)));
	assign fx85x = (((!ax84x) & (!bx84x) & (!g180) & (!ax85x) & (bx85x)) + ((!ax84x) & (!bx84x) & (!g180) & (ax85x) & (!bx85x)) + ((!ax84x) & (!bx84x) & (g180) & (!ax85x) & (bx85x)) + ((!ax84x) & (!bx84x) & (g180) & (ax85x) & (!bx85x)) + ((!ax84x) & (bx84x) & (!g180) & (!ax85x) & (bx85x)) + ((!ax84x) & (bx84x) & (!g180) & (ax85x) & (!bx85x)) + ((!ax84x) & (bx84x) & (g180) & (!ax85x) & (!bx85x)) + ((!ax84x) & (bx84x) & (g180) & (ax85x) & (bx85x)) + ((ax84x) & (!bx84x) & (!g180) & (!ax85x) & (bx85x)) + ((ax84x) & (!bx84x) & (!g180) & (ax85x) & (!bx85x)) + ((ax84x) & (!bx84x) & (g180) & (!ax85x) & (!bx85x)) + ((ax84x) & (!bx84x) & (g180) & (ax85x) & (bx85x)) + ((ax84x) & (bx84x) & (!g180) & (!ax85x) & (!bx85x)) + ((ax84x) & (bx84x) & (!g180) & (ax85x) & (bx85x)) + ((ax84x) & (bx84x) & (g180) & (!ax85x) & (!bx85x)) + ((ax84x) & (bx84x) & (g180) & (ax85x) & (bx85x)));
	assign g183 = (((ax85x) & (bx85x)));
	assign g184 = (((!ax85x) & (!bx85x)));
	assign g185 = (((!ax83x) & (!bx83x) & (!g178) & (ax84x) & (bx84x) & (!g184)) + ((!ax83x) & (!bx83x) & (g178) & (ax84x) & (bx84x) & (!g184)) + ((!ax83x) & (bx83x) & (!g178) & (!ax84x) & (bx84x) & (!g184)) + ((!ax83x) & (bx83x) & (!g178) & (ax84x) & (!bx84x) & (!g184)) + ((!ax83x) & (bx83x) & (!g178) & (ax84x) & (bx84x) & (!g184)) + ((!ax83x) & (bx83x) & (g178) & (ax84x) & (bx84x) & (!g184)) + ((ax83x) & (!bx83x) & (!g178) & (!ax84x) & (bx84x) & (!g184)) + ((ax83x) & (!bx83x) & (!g178) & (ax84x) & (!bx84x) & (!g184)) + ((ax83x) & (!bx83x) & (!g178) & (ax84x) & (bx84x) & (!g184)) + ((ax83x) & (!bx83x) & (g178) & (ax84x) & (bx84x) & (!g184)) + ((ax83x) & (bx83x) & (!g178) & (!ax84x) & (bx84x) & (!g184)) + ((ax83x) & (bx83x) & (!g178) & (ax84x) & (!bx84x) & (!g184)) + ((ax83x) & (bx83x) & (!g178) & (ax84x) & (bx84x) & (!g184)) + ((ax83x) & (bx83x) & (g178) & (!ax84x) & (bx84x) & (!g184)) + ((ax83x) & (bx83x) & (g178) & (ax84x) & (!bx84x) & (!g184)) + ((ax83x) & (bx83x) & (g178) & (ax84x) & (bx84x) & (!g184)));
	assign g186 = (((!g183) & (!g185)));
	assign fx86x = (((!ax86x) & (!bx86x) & (!g186)) + ((!ax86x) & (bx86x) & (g186)) + ((ax86x) & (!bx86x) & (g186)) + ((ax86x) & (bx86x) & (!g186)));
	assign fx87x = (((!ax86x) & (!bx86x) & (!g186) & (!ax87x) & (bx87x)) + ((!ax86x) & (!bx86x) & (!g186) & (ax87x) & (!bx87x)) + ((!ax86x) & (!bx86x) & (g186) & (!ax87x) & (bx87x)) + ((!ax86x) & (!bx86x) & (g186) & (ax87x) & (!bx87x)) + ((!ax86x) & (bx86x) & (!g186) & (!ax87x) & (!bx87x)) + ((!ax86x) & (bx86x) & (!g186) & (ax87x) & (bx87x)) + ((!ax86x) & (bx86x) & (g186) & (!ax87x) & (bx87x)) + ((!ax86x) & (bx86x) & (g186) & (ax87x) & (!bx87x)) + ((ax86x) & (!bx86x) & (!g186) & (!ax87x) & (!bx87x)) + ((ax86x) & (!bx86x) & (!g186) & (ax87x) & (bx87x)) + ((ax86x) & (!bx86x) & (g186) & (!ax87x) & (bx87x)) + ((ax86x) & (!bx86x) & (g186) & (ax87x) & (!bx87x)) + ((ax86x) & (bx86x) & (!g186) & (!ax87x) & (!bx87x)) + ((ax86x) & (bx86x) & (!g186) & (ax87x) & (bx87x)) + ((ax86x) & (bx86x) & (g186) & (!ax87x) & (!bx87x)) + ((ax86x) & (bx86x) & (g186) & (ax87x) & (bx87x)));
	assign g189 = (((!ax86x) & (!bx86x) & (!g183) & (!g185) & (!ax87x) & (!bx87x)) + ((!ax86x) & (!bx86x) & (!g183) & (!g185) & (!ax87x) & (bx87x)) + ((!ax86x) & (!bx86x) & (!g183) & (!g185) & (ax87x) & (!bx87x)) + ((!ax86x) & (!bx86x) & (!g183) & (g185) & (!ax87x) & (!bx87x)) + ((!ax86x) & (!bx86x) & (!g183) & (g185) & (!ax87x) & (bx87x)) + ((!ax86x) & (!bx86x) & (!g183) & (g185) & (ax87x) & (!bx87x)) + ((!ax86x) & (!bx86x) & (g183) & (!g185) & (!ax87x) & (!bx87x)) + ((!ax86x) & (!bx86x) & (g183) & (!g185) & (!ax87x) & (bx87x)) + ((!ax86x) & (!bx86x) & (g183) & (!g185) & (ax87x) & (!bx87x)) + ((!ax86x) & (!bx86x) & (g183) & (g185) & (!ax87x) & (!bx87x)) + ((!ax86x) & (!bx86x) & (g183) & (g185) & (!ax87x) & (bx87x)) + ((!ax86x) & (!bx86x) & (g183) & (g185) & (ax87x) & (!bx87x)) + ((!ax86x) & (bx86x) & (!g183) & (!g185) & (!ax87x) & (!bx87x)) + ((!ax86x) & (bx86x) & (!g183) & (!g185) & (!ax87x) & (bx87x)) + ((!ax86x) & (bx86x) & (!g183) & (!g185) & (ax87x) & (!bx87x)) + ((!ax86x) & (bx86x) & (!g183) & (g185) & (!ax87x) & (!bx87x)) + ((!ax86x) & (bx86x) & (g183) & (!g185) & (!ax87x) & (!bx87x)) + ((!ax86x) & (bx86x) & (g183) & (g185) & (!ax87x) & (!bx87x)) + ((ax86x) & (!bx86x) & (!g183) & (!g185) & (!ax87x) & (!bx87x)) + ((ax86x) & (!bx86x) & (!g183) & (!g185) & (!ax87x) & (bx87x)) + ((ax86x) & (!bx86x) & (!g183) & (!g185) & (ax87x) & (!bx87x)) + ((ax86x) & (!bx86x) & (!g183) & (g185) & (!ax87x) & (!bx87x)) + ((ax86x) & (!bx86x) & (g183) & (!g185) & (!ax87x) & (!bx87x)) + ((ax86x) & (!bx86x) & (g183) & (g185) & (!ax87x) & (!bx87x)) + ((ax86x) & (bx86x) & (!g183) & (!g185) & (!ax87x) & (!bx87x)) + ((ax86x) & (bx86x) & (!g183) & (g185) & (!ax87x) & (!bx87x)) + ((ax86x) & (bx86x) & (g183) & (!g185) & (!ax87x) & (!bx87x)) + ((ax86x) & (bx86x) & (g183) & (g185) & (!ax87x) & (!bx87x)));
	assign fx88x = (((!ax88x) & (!bx88x) & (!g189)) + ((!ax88x) & (bx88x) & (g189)) + ((ax88x) & (!bx88x) & (g189)) + ((ax88x) & (bx88x) & (!g189)));
	assign g191 = (((!ax88x) & (bx88x) & (!g189)) + ((ax88x) & (!bx88x) & (!g189)) + ((ax88x) & (bx88x) & (!g189)) + ((ax88x) & (bx88x) & (g189)));
	assign fx89x = (((!ax89x) & (!bx89x) & (g191)) + ((!ax89x) & (bx89x) & (!g191)) + ((ax89x) & (!bx89x) & (!g191)) + ((ax89x) & (bx89x) & (g191)));
	assign fx90x = (((!ax89x) & (!bx89x) & (!g191) & (!ax90x) & (bx90x)) + ((!ax89x) & (!bx89x) & (!g191) & (ax90x) & (!bx90x)) + ((!ax89x) & (!bx89x) & (g191) & (!ax90x) & (bx90x)) + ((!ax89x) & (!bx89x) & (g191) & (ax90x) & (!bx90x)) + ((!ax89x) & (bx89x) & (!g191) & (!ax90x) & (bx90x)) + ((!ax89x) & (bx89x) & (!g191) & (ax90x) & (!bx90x)) + ((!ax89x) & (bx89x) & (g191) & (!ax90x) & (!bx90x)) + ((!ax89x) & (bx89x) & (g191) & (ax90x) & (bx90x)) + ((ax89x) & (!bx89x) & (!g191) & (!ax90x) & (bx90x)) + ((ax89x) & (!bx89x) & (!g191) & (ax90x) & (!bx90x)) + ((ax89x) & (!bx89x) & (g191) & (!ax90x) & (!bx90x)) + ((ax89x) & (!bx89x) & (g191) & (ax90x) & (bx90x)) + ((ax89x) & (bx89x) & (!g191) & (!ax90x) & (!bx90x)) + ((ax89x) & (bx89x) & (!g191) & (ax90x) & (bx90x)) + ((ax89x) & (bx89x) & (g191) & (!ax90x) & (!bx90x)) + ((ax89x) & (bx89x) & (g191) & (ax90x) & (bx90x)));
	assign g194 = (((ax90x) & (bx90x)));
	assign g195 = (((!ax90x) & (!bx90x)));
	assign g196 = (((!ax88x) & (!bx88x) & (!g189) & (ax89x) & (bx89x) & (!g195)) + ((!ax88x) & (!bx88x) & (g189) & (ax89x) & (bx89x) & (!g195)) + ((!ax88x) & (bx88x) & (!g189) & (!ax89x) & (bx89x) & (!g195)) + ((!ax88x) & (bx88x) & (!g189) & (ax89x) & (!bx89x) & (!g195)) + ((!ax88x) & (bx88x) & (!g189) & (ax89x) & (bx89x) & (!g195)) + ((!ax88x) & (bx88x) & (g189) & (ax89x) & (bx89x) & (!g195)) + ((ax88x) & (!bx88x) & (!g189) & (!ax89x) & (bx89x) & (!g195)) + ((ax88x) & (!bx88x) & (!g189) & (ax89x) & (!bx89x) & (!g195)) + ((ax88x) & (!bx88x) & (!g189) & (ax89x) & (bx89x) & (!g195)) + ((ax88x) & (!bx88x) & (g189) & (ax89x) & (bx89x) & (!g195)) + ((ax88x) & (bx88x) & (!g189) & (!ax89x) & (bx89x) & (!g195)) + ((ax88x) & (bx88x) & (!g189) & (ax89x) & (!bx89x) & (!g195)) + ((ax88x) & (bx88x) & (!g189) & (ax89x) & (bx89x) & (!g195)) + ((ax88x) & (bx88x) & (g189) & (!ax89x) & (bx89x) & (!g195)) + ((ax88x) & (bx88x) & (g189) & (ax89x) & (!bx89x) & (!g195)) + ((ax88x) & (bx88x) & (g189) & (ax89x) & (bx89x) & (!g195)));
	assign fx91x = (((!ax91x) & (!bx91x) & (!g194) & (g196)) + ((!ax91x) & (!bx91x) & (g194) & (!g196)) + ((!ax91x) & (!bx91x) & (g194) & (g196)) + ((!ax91x) & (bx91x) & (!g194) & (!g196)) + ((ax91x) & (!bx91x) & (!g194) & (!g196)) + ((ax91x) & (bx91x) & (!g194) & (g196)) + ((ax91x) & (bx91x) & (g194) & (!g196)) + ((ax91x) & (bx91x) & (g194) & (g196)));
	assign fx92x = (((!ax91x) & (!bx91x) & (!g194) & (!g196) & (!ax92x) & (bx92x)) + ((!ax91x) & (!bx91x) & (!g194) & (!g196) & (ax92x) & (!bx92x)) + ((!ax91x) & (!bx91x) & (!g194) & (g196) & (!ax92x) & (bx92x)) + ((!ax91x) & (!bx91x) & (!g194) & (g196) & (ax92x) & (!bx92x)) + ((!ax91x) & (!bx91x) & (g194) & (!g196) & (!ax92x) & (bx92x)) + ((!ax91x) & (!bx91x) & (g194) & (!g196) & (ax92x) & (!bx92x)) + ((!ax91x) & (!bx91x) & (g194) & (g196) & (!ax92x) & (bx92x)) + ((!ax91x) & (!bx91x) & (g194) & (g196) & (ax92x) & (!bx92x)) + ((!ax91x) & (bx91x) & (!g194) & (!g196) & (!ax92x) & (bx92x)) + ((!ax91x) & (bx91x) & (!g194) & (!g196) & (ax92x) & (!bx92x)) + ((!ax91x) & (bx91x) & (!g194) & (g196) & (!ax92x) & (!bx92x)) + ((!ax91x) & (bx91x) & (!g194) & (g196) & (ax92x) & (bx92x)) + ((!ax91x) & (bx91x) & (g194) & (!g196) & (!ax92x) & (!bx92x)) + ((!ax91x) & (bx91x) & (g194) & (!g196) & (ax92x) & (bx92x)) + ((!ax91x) & (bx91x) & (g194) & (g196) & (!ax92x) & (!bx92x)) + ((!ax91x) & (bx91x) & (g194) & (g196) & (ax92x) & (bx92x)) + ((ax91x) & (!bx91x) & (!g194) & (!g196) & (!ax92x) & (bx92x)) + ((ax91x) & (!bx91x) & (!g194) & (!g196) & (ax92x) & (!bx92x)) + ((ax91x) & (!bx91x) & (!g194) & (g196) & (!ax92x) & (!bx92x)) + ((ax91x) & (!bx91x) & (!g194) & (g196) & (ax92x) & (bx92x)) + ((ax91x) & (!bx91x) & (g194) & (!g196) & (!ax92x) & (!bx92x)) + ((ax91x) & (!bx91x) & (g194) & (!g196) & (ax92x) & (bx92x)) + ((ax91x) & (!bx91x) & (g194) & (g196) & (!ax92x) & (!bx92x)) + ((ax91x) & (!bx91x) & (g194) & (g196) & (ax92x) & (bx92x)) + ((ax91x) & (bx91x) & (!g194) & (!g196) & (!ax92x) & (!bx92x)) + ((ax91x) & (bx91x) & (!g194) & (!g196) & (ax92x) & (bx92x)) + ((ax91x) & (bx91x) & (!g194) & (g196) & (!ax92x) & (!bx92x)) + ((ax91x) & (bx91x) & (!g194) & (g196) & (ax92x) & (bx92x)) + ((ax91x) & (bx91x) & (g194) & (!g196) & (!ax92x) & (!bx92x)) + ((ax91x) & (bx91x) & (g194) & (!g196) & (ax92x) & (bx92x)) + ((ax91x) & (bx91x) & (g194) & (g196) & (!ax92x) & (!bx92x)) + ((ax91x) & (bx91x) & (g194) & (g196) & (ax92x) & (bx92x)));
	assign g199 = (((!ax91x) & (!bx91x) & (!g194) & (!g196) & (!ax92x) & (!bx92x)) + ((!ax91x) & (!bx91x) & (!g194) & (!g196) & (!ax92x) & (bx92x)) + ((!ax91x) & (!bx91x) & (!g194) & (!g196) & (ax92x) & (!bx92x)) + ((!ax91x) & (!bx91x) & (!g194) & (g196) & (!ax92x) & (!bx92x)) + ((!ax91x) & (!bx91x) & (!g194) & (g196) & (!ax92x) & (bx92x)) + ((!ax91x) & (!bx91x) & (!g194) & (g196) & (ax92x) & (!bx92x)) + ((!ax91x) & (!bx91x) & (g194) & (!g196) & (!ax92x) & (!bx92x)) + ((!ax91x) & (!bx91x) & (g194) & (!g196) & (!ax92x) & (bx92x)) + ((!ax91x) & (!bx91x) & (g194) & (!g196) & (ax92x) & (!bx92x)) + ((!ax91x) & (!bx91x) & (g194) & (g196) & (!ax92x) & (!bx92x)) + ((!ax91x) & (!bx91x) & (g194) & (g196) & (!ax92x) & (bx92x)) + ((!ax91x) & (!bx91x) & (g194) & (g196) & (ax92x) & (!bx92x)) + ((!ax91x) & (bx91x) & (!g194) & (!g196) & (!ax92x) & (!bx92x)) + ((!ax91x) & (bx91x) & (!g194) & (!g196) & (!ax92x) & (bx92x)) + ((!ax91x) & (bx91x) & (!g194) & (!g196) & (ax92x) & (!bx92x)) + ((!ax91x) & (bx91x) & (!g194) & (g196) & (!ax92x) & (!bx92x)) + ((!ax91x) & (bx91x) & (g194) & (!g196) & (!ax92x) & (!bx92x)) + ((!ax91x) & (bx91x) & (g194) & (g196) & (!ax92x) & (!bx92x)) + ((ax91x) & (!bx91x) & (!g194) & (!g196) & (!ax92x) & (!bx92x)) + ((ax91x) & (!bx91x) & (!g194) & (!g196) & (!ax92x) & (bx92x)) + ((ax91x) & (!bx91x) & (!g194) & (!g196) & (ax92x) & (!bx92x)) + ((ax91x) & (!bx91x) & (!g194) & (g196) & (!ax92x) & (!bx92x)) + ((ax91x) & (!bx91x) & (g194) & (!g196) & (!ax92x) & (!bx92x)) + ((ax91x) & (!bx91x) & (g194) & (g196) & (!ax92x) & (!bx92x)) + ((ax91x) & (bx91x) & (!g194) & (!g196) & (!ax92x) & (!bx92x)) + ((ax91x) & (bx91x) & (!g194) & (g196) & (!ax92x) & (!bx92x)) + ((ax91x) & (bx91x) & (g194) & (!g196) & (!ax92x) & (!bx92x)) + ((ax91x) & (bx91x) & (g194) & (g196) & (!ax92x) & (!bx92x)));
	assign fx93x = (((!ax93x) & (!bx93x) & (!g199)) + ((!ax93x) & (bx93x) & (g199)) + ((ax93x) & (!bx93x) & (g199)) + ((ax93x) & (bx93x) & (!g199)));
	assign g201 = (((!ax93x) & (bx93x) & (!g199)) + ((ax93x) & (!bx93x) & (!g199)) + ((ax93x) & (bx93x) & (!g199)) + ((ax93x) & (bx93x) & (g199)));
	assign fx94x = (((!ax94x) & (!bx94x) & (g201)) + ((!ax94x) & (bx94x) & (!g201)) + ((ax94x) & (!bx94x) & (!g201)) + ((ax94x) & (bx94x) & (g201)));
	assign fx95x = (((!ax94x) & (!bx94x) & (!g201) & (!ax95x) & (bx95x)) + ((!ax94x) & (!bx94x) & (!g201) & (ax95x) & (!bx95x)) + ((!ax94x) & (!bx94x) & (g201) & (!ax95x) & (bx95x)) + ((!ax94x) & (!bx94x) & (g201) & (ax95x) & (!bx95x)) + ((!ax94x) & (bx94x) & (!g201) & (!ax95x) & (bx95x)) + ((!ax94x) & (bx94x) & (!g201) & (ax95x) & (!bx95x)) + ((!ax94x) & (bx94x) & (g201) & (!ax95x) & (!bx95x)) + ((!ax94x) & (bx94x) & (g201) & (ax95x) & (bx95x)) + ((ax94x) & (!bx94x) & (!g201) & (!ax95x) & (bx95x)) + ((ax94x) & (!bx94x) & (!g201) & (ax95x) & (!bx95x)) + ((ax94x) & (!bx94x) & (g201) & (!ax95x) & (!bx95x)) + ((ax94x) & (!bx94x) & (g201) & (ax95x) & (bx95x)) + ((ax94x) & (bx94x) & (!g201) & (!ax95x) & (!bx95x)) + ((ax94x) & (bx94x) & (!g201) & (ax95x) & (bx95x)) + ((ax94x) & (bx94x) & (g201) & (!ax95x) & (!bx95x)) + ((ax94x) & (bx94x) & (g201) & (ax95x) & (bx95x)));
	assign g204 = (((ax95x) & (bx95x)));
	assign g205 = (((!ax95x) & (!bx95x)));
	assign g206 = (((!ax93x) & (!bx93x) & (!g199) & (ax94x) & (bx94x) & (!g205)) + ((!ax93x) & (!bx93x) & (g199) & (ax94x) & (bx94x) & (!g205)) + ((!ax93x) & (bx93x) & (!g199) & (!ax94x) & (bx94x) & (!g205)) + ((!ax93x) & (bx93x) & (!g199) & (ax94x) & (!bx94x) & (!g205)) + ((!ax93x) & (bx93x) & (!g199) & (ax94x) & (bx94x) & (!g205)) + ((!ax93x) & (bx93x) & (g199) & (ax94x) & (bx94x) & (!g205)) + ((ax93x) & (!bx93x) & (!g199) & (!ax94x) & (bx94x) & (!g205)) + ((ax93x) & (!bx93x) & (!g199) & (ax94x) & (!bx94x) & (!g205)) + ((ax93x) & (!bx93x) & (!g199) & (ax94x) & (bx94x) & (!g205)) + ((ax93x) & (!bx93x) & (g199) & (ax94x) & (bx94x) & (!g205)) + ((ax93x) & (bx93x) & (!g199) & (!ax94x) & (bx94x) & (!g205)) + ((ax93x) & (bx93x) & (!g199) & (ax94x) & (!bx94x) & (!g205)) + ((ax93x) & (bx93x) & (!g199) & (ax94x) & (bx94x) & (!g205)) + ((ax93x) & (bx93x) & (g199) & (!ax94x) & (bx94x) & (!g205)) + ((ax93x) & (bx93x) & (g199) & (ax94x) & (!bx94x) & (!g205)) + ((ax93x) & (bx93x) & (g199) & (ax94x) & (bx94x) & (!g205)));
	assign g207 = (((!g204) & (!g206)));
	assign fx96x = (((!ax96x) & (!bx96x) & (!g207)) + ((!ax96x) & (bx96x) & (g207)) + ((ax96x) & (!bx96x) & (g207)) + ((ax96x) & (bx96x) & (!g207)));
	assign fx97x = (((!ax96x) & (!bx96x) & (!g207) & (!ax97x) & (bx97x)) + ((!ax96x) & (!bx96x) & (!g207) & (ax97x) & (!bx97x)) + ((!ax96x) & (!bx96x) & (g207) & (!ax97x) & (bx97x)) + ((!ax96x) & (!bx96x) & (g207) & (ax97x) & (!bx97x)) + ((!ax96x) & (bx96x) & (!g207) & (!ax97x) & (!bx97x)) + ((!ax96x) & (bx96x) & (!g207) & (ax97x) & (bx97x)) + ((!ax96x) & (bx96x) & (g207) & (!ax97x) & (bx97x)) + ((!ax96x) & (bx96x) & (g207) & (ax97x) & (!bx97x)) + ((ax96x) & (!bx96x) & (!g207) & (!ax97x) & (!bx97x)) + ((ax96x) & (!bx96x) & (!g207) & (ax97x) & (bx97x)) + ((ax96x) & (!bx96x) & (g207) & (!ax97x) & (bx97x)) + ((ax96x) & (!bx96x) & (g207) & (ax97x) & (!bx97x)) + ((ax96x) & (bx96x) & (!g207) & (!ax97x) & (!bx97x)) + ((ax96x) & (bx96x) & (!g207) & (ax97x) & (bx97x)) + ((ax96x) & (bx96x) & (g207) & (!ax97x) & (!bx97x)) + ((ax96x) & (bx96x) & (g207) & (ax97x) & (bx97x)));
	assign g210 = (((!ax96x) & (!bx96x) & (!g204) & (!g206) & (!ax97x) & (!bx97x)) + ((!ax96x) & (!bx96x) & (!g204) & (!g206) & (!ax97x) & (bx97x)) + ((!ax96x) & (!bx96x) & (!g204) & (!g206) & (ax97x) & (!bx97x)) + ((!ax96x) & (!bx96x) & (!g204) & (g206) & (!ax97x) & (!bx97x)) + ((!ax96x) & (!bx96x) & (!g204) & (g206) & (!ax97x) & (bx97x)) + ((!ax96x) & (!bx96x) & (!g204) & (g206) & (ax97x) & (!bx97x)) + ((!ax96x) & (!bx96x) & (g204) & (!g206) & (!ax97x) & (!bx97x)) + ((!ax96x) & (!bx96x) & (g204) & (!g206) & (!ax97x) & (bx97x)) + ((!ax96x) & (!bx96x) & (g204) & (!g206) & (ax97x) & (!bx97x)) + ((!ax96x) & (!bx96x) & (g204) & (g206) & (!ax97x) & (!bx97x)) + ((!ax96x) & (!bx96x) & (g204) & (g206) & (!ax97x) & (bx97x)) + ((!ax96x) & (!bx96x) & (g204) & (g206) & (ax97x) & (!bx97x)) + ((!ax96x) & (bx96x) & (!g204) & (!g206) & (!ax97x) & (!bx97x)) + ((!ax96x) & (bx96x) & (!g204) & (!g206) & (!ax97x) & (bx97x)) + ((!ax96x) & (bx96x) & (!g204) & (!g206) & (ax97x) & (!bx97x)) + ((!ax96x) & (bx96x) & (!g204) & (g206) & (!ax97x) & (!bx97x)) + ((!ax96x) & (bx96x) & (g204) & (!g206) & (!ax97x) & (!bx97x)) + ((!ax96x) & (bx96x) & (g204) & (g206) & (!ax97x) & (!bx97x)) + ((ax96x) & (!bx96x) & (!g204) & (!g206) & (!ax97x) & (!bx97x)) + ((ax96x) & (!bx96x) & (!g204) & (!g206) & (!ax97x) & (bx97x)) + ((ax96x) & (!bx96x) & (!g204) & (!g206) & (ax97x) & (!bx97x)) + ((ax96x) & (!bx96x) & (!g204) & (g206) & (!ax97x) & (!bx97x)) + ((ax96x) & (!bx96x) & (g204) & (!g206) & (!ax97x) & (!bx97x)) + ((ax96x) & (!bx96x) & (g204) & (g206) & (!ax97x) & (!bx97x)) + ((ax96x) & (bx96x) & (!g204) & (!g206) & (!ax97x) & (!bx97x)) + ((ax96x) & (bx96x) & (!g204) & (g206) & (!ax97x) & (!bx97x)) + ((ax96x) & (bx96x) & (g204) & (!g206) & (!ax97x) & (!bx97x)) + ((ax96x) & (bx96x) & (g204) & (g206) & (!ax97x) & (!bx97x)));
	assign fx98x = (((!ax98x) & (!bx98x) & (!g210)) + ((!ax98x) & (bx98x) & (g210)) + ((ax98x) & (!bx98x) & (g210)) + ((ax98x) & (bx98x) & (!g210)));
	assign g212 = (((!ax98x) & (bx98x) & (!g210)) + ((ax98x) & (!bx98x) & (!g210)) + ((ax98x) & (bx98x) & (!g210)) + ((ax98x) & (bx98x) & (g210)));
	assign fx99x = (((!ax99x) & (!bx99x) & (g212)) + ((!ax99x) & (bx99x) & (!g212)) + ((ax99x) & (!bx99x) & (!g212)) + ((ax99x) & (bx99x) & (g212)));
	assign fx100x = (((!ax99x) & (!bx99x) & (!g212) & (!ax100x) & (bx100x)) + ((!ax99x) & (!bx99x) & (!g212) & (ax100x) & (!bx100x)) + ((!ax99x) & (!bx99x) & (g212) & (!ax100x) & (bx100x)) + ((!ax99x) & (!bx99x) & (g212) & (ax100x) & (!bx100x)) + ((!ax99x) & (bx99x) & (!g212) & (!ax100x) & (bx100x)) + ((!ax99x) & (bx99x) & (!g212) & (ax100x) & (!bx100x)) + ((!ax99x) & (bx99x) & (g212) & (!ax100x) & (!bx100x)) + ((!ax99x) & (bx99x) & (g212) & (ax100x) & (bx100x)) + ((ax99x) & (!bx99x) & (!g212) & (!ax100x) & (bx100x)) + ((ax99x) & (!bx99x) & (!g212) & (ax100x) & (!bx100x)) + ((ax99x) & (!bx99x) & (g212) & (!ax100x) & (!bx100x)) + ((ax99x) & (!bx99x) & (g212) & (ax100x) & (bx100x)) + ((ax99x) & (bx99x) & (!g212) & (!ax100x) & (!bx100x)) + ((ax99x) & (bx99x) & (!g212) & (ax100x) & (bx100x)) + ((ax99x) & (bx99x) & (g212) & (!ax100x) & (!bx100x)) + ((ax99x) & (bx99x) & (g212) & (ax100x) & (bx100x)));
	assign g215 = (((ax100x) & (bx100x)));
	assign g216 = (((!ax100x) & (!bx100x)));
	assign g217 = (((!ax98x) & (!bx98x) & (!g210) & (ax99x) & (bx99x) & (!g216)) + ((!ax98x) & (!bx98x) & (g210) & (ax99x) & (bx99x) & (!g216)) + ((!ax98x) & (bx98x) & (!g210) & (!ax99x) & (bx99x) & (!g216)) + ((!ax98x) & (bx98x) & (!g210) & (ax99x) & (!bx99x) & (!g216)) + ((!ax98x) & (bx98x) & (!g210) & (ax99x) & (bx99x) & (!g216)) + ((!ax98x) & (bx98x) & (g210) & (ax99x) & (bx99x) & (!g216)) + ((ax98x) & (!bx98x) & (!g210) & (!ax99x) & (bx99x) & (!g216)) + ((ax98x) & (!bx98x) & (!g210) & (ax99x) & (!bx99x) & (!g216)) + ((ax98x) & (!bx98x) & (!g210) & (ax99x) & (bx99x) & (!g216)) + ((ax98x) & (!bx98x) & (g210) & (ax99x) & (bx99x) & (!g216)) + ((ax98x) & (bx98x) & (!g210) & (!ax99x) & (bx99x) & (!g216)) + ((ax98x) & (bx98x) & (!g210) & (ax99x) & (!bx99x) & (!g216)) + ((ax98x) & (bx98x) & (!g210) & (ax99x) & (bx99x) & (!g216)) + ((ax98x) & (bx98x) & (g210) & (!ax99x) & (bx99x) & (!g216)) + ((ax98x) & (bx98x) & (g210) & (ax99x) & (!bx99x) & (!g216)) + ((ax98x) & (bx98x) & (g210) & (ax99x) & (bx99x) & (!g216)));
	assign g218 = (((!g215) & (!g217)));
	assign fx101x = (((!ax101x) & (!bx101x) & (!g218)) + ((!ax101x) & (bx101x) & (g218)) + ((ax101x) & (!bx101x) & (g218)) + ((ax101x) & (bx101x) & (!g218)));
	assign fx102x = (((!ax101x) & (!bx101x) & (!g218) & (!ax102x) & (bx102x)) + ((!ax101x) & (!bx101x) & (!g218) & (ax102x) & (!bx102x)) + ((!ax101x) & (!bx101x) & (g218) & (!ax102x) & (bx102x)) + ((!ax101x) & (!bx101x) & (g218) & (ax102x) & (!bx102x)) + ((!ax101x) & (bx101x) & (!g218) & (!ax102x) & (!bx102x)) + ((!ax101x) & (bx101x) & (!g218) & (ax102x) & (bx102x)) + ((!ax101x) & (bx101x) & (g218) & (!ax102x) & (bx102x)) + ((!ax101x) & (bx101x) & (g218) & (ax102x) & (!bx102x)) + ((ax101x) & (!bx101x) & (!g218) & (!ax102x) & (!bx102x)) + ((ax101x) & (!bx101x) & (!g218) & (ax102x) & (bx102x)) + ((ax101x) & (!bx101x) & (g218) & (!ax102x) & (bx102x)) + ((ax101x) & (!bx101x) & (g218) & (ax102x) & (!bx102x)) + ((ax101x) & (bx101x) & (!g218) & (!ax102x) & (!bx102x)) + ((ax101x) & (bx101x) & (!g218) & (ax102x) & (bx102x)) + ((ax101x) & (bx101x) & (g218) & (!ax102x) & (!bx102x)) + ((ax101x) & (bx101x) & (g218) & (ax102x) & (bx102x)));
	assign g221 = (((!ax101x) & (!bx101x) & (!g215) & (!g217) & (!ax102x) & (!bx102x)) + ((!ax101x) & (!bx101x) & (!g215) & (!g217) & (!ax102x) & (bx102x)) + ((!ax101x) & (!bx101x) & (!g215) & (!g217) & (ax102x) & (!bx102x)) + ((!ax101x) & (!bx101x) & (!g215) & (g217) & (!ax102x) & (!bx102x)) + ((!ax101x) & (!bx101x) & (!g215) & (g217) & (!ax102x) & (bx102x)) + ((!ax101x) & (!bx101x) & (!g215) & (g217) & (ax102x) & (!bx102x)) + ((!ax101x) & (!bx101x) & (g215) & (!g217) & (!ax102x) & (!bx102x)) + ((!ax101x) & (!bx101x) & (g215) & (!g217) & (!ax102x) & (bx102x)) + ((!ax101x) & (!bx101x) & (g215) & (!g217) & (ax102x) & (!bx102x)) + ((!ax101x) & (!bx101x) & (g215) & (g217) & (!ax102x) & (!bx102x)) + ((!ax101x) & (!bx101x) & (g215) & (g217) & (!ax102x) & (bx102x)) + ((!ax101x) & (!bx101x) & (g215) & (g217) & (ax102x) & (!bx102x)) + ((!ax101x) & (bx101x) & (!g215) & (!g217) & (!ax102x) & (!bx102x)) + ((!ax101x) & (bx101x) & (!g215) & (!g217) & (!ax102x) & (bx102x)) + ((!ax101x) & (bx101x) & (!g215) & (!g217) & (ax102x) & (!bx102x)) + ((!ax101x) & (bx101x) & (!g215) & (g217) & (!ax102x) & (!bx102x)) + ((!ax101x) & (bx101x) & (g215) & (!g217) & (!ax102x) & (!bx102x)) + ((!ax101x) & (bx101x) & (g215) & (g217) & (!ax102x) & (!bx102x)) + ((ax101x) & (!bx101x) & (!g215) & (!g217) & (!ax102x) & (!bx102x)) + ((ax101x) & (!bx101x) & (!g215) & (!g217) & (!ax102x) & (bx102x)) + ((ax101x) & (!bx101x) & (!g215) & (!g217) & (ax102x) & (!bx102x)) + ((ax101x) & (!bx101x) & (!g215) & (g217) & (!ax102x) & (!bx102x)) + ((ax101x) & (!bx101x) & (g215) & (!g217) & (!ax102x) & (!bx102x)) + ((ax101x) & (!bx101x) & (g215) & (g217) & (!ax102x) & (!bx102x)) + ((ax101x) & (bx101x) & (!g215) & (!g217) & (!ax102x) & (!bx102x)) + ((ax101x) & (bx101x) & (!g215) & (g217) & (!ax102x) & (!bx102x)) + ((ax101x) & (bx101x) & (g215) & (!g217) & (!ax102x) & (!bx102x)) + ((ax101x) & (bx101x) & (g215) & (g217) & (!ax102x) & (!bx102x)));
	assign fx103x = (((!ax103x) & (!bx103x) & (!g221)) + ((!ax103x) & (bx103x) & (g221)) + ((ax103x) & (!bx103x) & (g221)) + ((ax103x) & (bx103x) & (!g221)));
	assign g223 = (((!ax103x) & (bx103x) & (!g221)) + ((ax103x) & (!bx103x) & (!g221)) + ((ax103x) & (bx103x) & (!g221)) + ((ax103x) & (bx103x) & (g221)));
	assign fx104x = (((!ax104x) & (!bx104x) & (g223)) + ((!ax104x) & (bx104x) & (!g223)) + ((ax104x) & (!bx104x) & (!g223)) + ((ax104x) & (bx104x) & (g223)));
	assign fx105x = (((!ax104x) & (!bx104x) & (!g223) & (!ax105x) & (bx105x)) + ((!ax104x) & (!bx104x) & (!g223) & (ax105x) & (!bx105x)) + ((!ax104x) & (!bx104x) & (g223) & (!ax105x) & (bx105x)) + ((!ax104x) & (!bx104x) & (g223) & (ax105x) & (!bx105x)) + ((!ax104x) & (bx104x) & (!g223) & (!ax105x) & (bx105x)) + ((!ax104x) & (bx104x) & (!g223) & (ax105x) & (!bx105x)) + ((!ax104x) & (bx104x) & (g223) & (!ax105x) & (!bx105x)) + ((!ax104x) & (bx104x) & (g223) & (ax105x) & (bx105x)) + ((ax104x) & (!bx104x) & (!g223) & (!ax105x) & (bx105x)) + ((ax104x) & (!bx104x) & (!g223) & (ax105x) & (!bx105x)) + ((ax104x) & (!bx104x) & (g223) & (!ax105x) & (!bx105x)) + ((ax104x) & (!bx104x) & (g223) & (ax105x) & (bx105x)) + ((ax104x) & (bx104x) & (!g223) & (!ax105x) & (!bx105x)) + ((ax104x) & (bx104x) & (!g223) & (ax105x) & (bx105x)) + ((ax104x) & (bx104x) & (g223) & (!ax105x) & (!bx105x)) + ((ax104x) & (bx104x) & (g223) & (ax105x) & (bx105x)));
	assign g226 = (((ax105x) & (bx105x)));
	assign g227 = (((!ax105x) & (!bx105x)));
	assign g228 = (((!ax103x) & (!bx103x) & (!g221) & (ax104x) & (bx104x) & (!g227)) + ((!ax103x) & (!bx103x) & (g221) & (ax104x) & (bx104x) & (!g227)) + ((!ax103x) & (bx103x) & (!g221) & (!ax104x) & (bx104x) & (!g227)) + ((!ax103x) & (bx103x) & (!g221) & (ax104x) & (!bx104x) & (!g227)) + ((!ax103x) & (bx103x) & (!g221) & (ax104x) & (bx104x) & (!g227)) + ((!ax103x) & (bx103x) & (g221) & (ax104x) & (bx104x) & (!g227)) + ((ax103x) & (!bx103x) & (!g221) & (!ax104x) & (bx104x) & (!g227)) + ((ax103x) & (!bx103x) & (!g221) & (ax104x) & (!bx104x) & (!g227)) + ((ax103x) & (!bx103x) & (!g221) & (ax104x) & (bx104x) & (!g227)) + ((ax103x) & (!bx103x) & (g221) & (ax104x) & (bx104x) & (!g227)) + ((ax103x) & (bx103x) & (!g221) & (!ax104x) & (bx104x) & (!g227)) + ((ax103x) & (bx103x) & (!g221) & (ax104x) & (!bx104x) & (!g227)) + ((ax103x) & (bx103x) & (!g221) & (ax104x) & (bx104x) & (!g227)) + ((ax103x) & (bx103x) & (g221) & (!ax104x) & (bx104x) & (!g227)) + ((ax103x) & (bx103x) & (g221) & (ax104x) & (!bx104x) & (!g227)) + ((ax103x) & (bx103x) & (g221) & (ax104x) & (bx104x) & (!g227)));
	assign fx106x = (((!ax106x) & (!bx106x) & (!g226) & (g228)) + ((!ax106x) & (!bx106x) & (g226) & (!g228)) + ((!ax106x) & (!bx106x) & (g226) & (g228)) + ((!ax106x) & (bx106x) & (!g226) & (!g228)) + ((ax106x) & (!bx106x) & (!g226) & (!g228)) + ((ax106x) & (bx106x) & (!g226) & (g228)) + ((ax106x) & (bx106x) & (g226) & (!g228)) + ((ax106x) & (bx106x) & (g226) & (g228)));
	assign fx107x = (((!ax106x) & (!bx106x) & (!g226) & (!g228) & (!ax107x) & (bx107x)) + ((!ax106x) & (!bx106x) & (!g226) & (!g228) & (ax107x) & (!bx107x)) + ((!ax106x) & (!bx106x) & (!g226) & (g228) & (!ax107x) & (bx107x)) + ((!ax106x) & (!bx106x) & (!g226) & (g228) & (ax107x) & (!bx107x)) + ((!ax106x) & (!bx106x) & (g226) & (!g228) & (!ax107x) & (bx107x)) + ((!ax106x) & (!bx106x) & (g226) & (!g228) & (ax107x) & (!bx107x)) + ((!ax106x) & (!bx106x) & (g226) & (g228) & (!ax107x) & (bx107x)) + ((!ax106x) & (!bx106x) & (g226) & (g228) & (ax107x) & (!bx107x)) + ((!ax106x) & (bx106x) & (!g226) & (!g228) & (!ax107x) & (bx107x)) + ((!ax106x) & (bx106x) & (!g226) & (!g228) & (ax107x) & (!bx107x)) + ((!ax106x) & (bx106x) & (!g226) & (g228) & (!ax107x) & (!bx107x)) + ((!ax106x) & (bx106x) & (!g226) & (g228) & (ax107x) & (bx107x)) + ((!ax106x) & (bx106x) & (g226) & (!g228) & (!ax107x) & (!bx107x)) + ((!ax106x) & (bx106x) & (g226) & (!g228) & (ax107x) & (bx107x)) + ((!ax106x) & (bx106x) & (g226) & (g228) & (!ax107x) & (!bx107x)) + ((!ax106x) & (bx106x) & (g226) & (g228) & (ax107x) & (bx107x)) + ((ax106x) & (!bx106x) & (!g226) & (!g228) & (!ax107x) & (bx107x)) + ((ax106x) & (!bx106x) & (!g226) & (!g228) & (ax107x) & (!bx107x)) + ((ax106x) & (!bx106x) & (!g226) & (g228) & (!ax107x) & (!bx107x)) + ((ax106x) & (!bx106x) & (!g226) & (g228) & (ax107x) & (bx107x)) + ((ax106x) & (!bx106x) & (g226) & (!g228) & (!ax107x) & (!bx107x)) + ((ax106x) & (!bx106x) & (g226) & (!g228) & (ax107x) & (bx107x)) + ((ax106x) & (!bx106x) & (g226) & (g228) & (!ax107x) & (!bx107x)) + ((ax106x) & (!bx106x) & (g226) & (g228) & (ax107x) & (bx107x)) + ((ax106x) & (bx106x) & (!g226) & (!g228) & (!ax107x) & (!bx107x)) + ((ax106x) & (bx106x) & (!g226) & (!g228) & (ax107x) & (bx107x)) + ((ax106x) & (bx106x) & (!g226) & (g228) & (!ax107x) & (!bx107x)) + ((ax106x) & (bx106x) & (!g226) & (g228) & (ax107x) & (bx107x)) + ((ax106x) & (bx106x) & (g226) & (!g228) & (!ax107x) & (!bx107x)) + ((ax106x) & (bx106x) & (g226) & (!g228) & (ax107x) & (bx107x)) + ((ax106x) & (bx106x) & (g226) & (g228) & (!ax107x) & (!bx107x)) + ((ax106x) & (bx106x) & (g226) & (g228) & (ax107x) & (bx107x)));
	assign g231 = (((!ax106x) & (!bx106x) & (!g226) & (!g228) & (!ax107x) & (!bx107x)) + ((!ax106x) & (!bx106x) & (!g226) & (!g228) & (!ax107x) & (bx107x)) + ((!ax106x) & (!bx106x) & (!g226) & (!g228) & (ax107x) & (!bx107x)) + ((!ax106x) & (!bx106x) & (!g226) & (g228) & (!ax107x) & (!bx107x)) + ((!ax106x) & (!bx106x) & (!g226) & (g228) & (!ax107x) & (bx107x)) + ((!ax106x) & (!bx106x) & (!g226) & (g228) & (ax107x) & (!bx107x)) + ((!ax106x) & (!bx106x) & (g226) & (!g228) & (!ax107x) & (!bx107x)) + ((!ax106x) & (!bx106x) & (g226) & (!g228) & (!ax107x) & (bx107x)) + ((!ax106x) & (!bx106x) & (g226) & (!g228) & (ax107x) & (!bx107x)) + ((!ax106x) & (!bx106x) & (g226) & (g228) & (!ax107x) & (!bx107x)) + ((!ax106x) & (!bx106x) & (g226) & (g228) & (!ax107x) & (bx107x)) + ((!ax106x) & (!bx106x) & (g226) & (g228) & (ax107x) & (!bx107x)) + ((!ax106x) & (bx106x) & (!g226) & (!g228) & (!ax107x) & (!bx107x)) + ((!ax106x) & (bx106x) & (!g226) & (!g228) & (!ax107x) & (bx107x)) + ((!ax106x) & (bx106x) & (!g226) & (!g228) & (ax107x) & (!bx107x)) + ((!ax106x) & (bx106x) & (!g226) & (g228) & (!ax107x) & (!bx107x)) + ((!ax106x) & (bx106x) & (g226) & (!g228) & (!ax107x) & (!bx107x)) + ((!ax106x) & (bx106x) & (g226) & (g228) & (!ax107x) & (!bx107x)) + ((ax106x) & (!bx106x) & (!g226) & (!g228) & (!ax107x) & (!bx107x)) + ((ax106x) & (!bx106x) & (!g226) & (!g228) & (!ax107x) & (bx107x)) + ((ax106x) & (!bx106x) & (!g226) & (!g228) & (ax107x) & (!bx107x)) + ((ax106x) & (!bx106x) & (!g226) & (g228) & (!ax107x) & (!bx107x)) + ((ax106x) & (!bx106x) & (g226) & (!g228) & (!ax107x) & (!bx107x)) + ((ax106x) & (!bx106x) & (g226) & (g228) & (!ax107x) & (!bx107x)) + ((ax106x) & (bx106x) & (!g226) & (!g228) & (!ax107x) & (!bx107x)) + ((ax106x) & (bx106x) & (!g226) & (g228) & (!ax107x) & (!bx107x)) + ((ax106x) & (bx106x) & (g226) & (!g228) & (!ax107x) & (!bx107x)) + ((ax106x) & (bx106x) & (g226) & (g228) & (!ax107x) & (!bx107x)));
	assign fx108x = (((!ax108x) & (!bx108x) & (!g231)) + ((!ax108x) & (bx108x) & (g231)) + ((ax108x) & (!bx108x) & (g231)) + ((ax108x) & (bx108x) & (!g231)));
	assign fx109x = (((!ax108x) & (!bx108x) & (!g231) & (!ax109x) & (bx109x)) + ((!ax108x) & (!bx108x) & (!g231) & (ax109x) & (!bx109x)) + ((!ax108x) & (!bx108x) & (g231) & (!ax109x) & (bx109x)) + ((!ax108x) & (!bx108x) & (g231) & (ax109x) & (!bx109x)) + ((!ax108x) & (bx108x) & (!g231) & (!ax109x) & (!bx109x)) + ((!ax108x) & (bx108x) & (!g231) & (ax109x) & (bx109x)) + ((!ax108x) & (bx108x) & (g231) & (!ax109x) & (bx109x)) + ((!ax108x) & (bx108x) & (g231) & (ax109x) & (!bx109x)) + ((ax108x) & (!bx108x) & (!g231) & (!ax109x) & (!bx109x)) + ((ax108x) & (!bx108x) & (!g231) & (ax109x) & (bx109x)) + ((ax108x) & (!bx108x) & (g231) & (!ax109x) & (bx109x)) + ((ax108x) & (!bx108x) & (g231) & (ax109x) & (!bx109x)) + ((ax108x) & (bx108x) & (!g231) & (!ax109x) & (!bx109x)) + ((ax108x) & (bx108x) & (!g231) & (ax109x) & (bx109x)) + ((ax108x) & (bx108x) & (g231) & (!ax109x) & (!bx109x)) + ((ax108x) & (bx108x) & (g231) & (ax109x) & (bx109x)));
	assign g234 = (((!ax110x) & (bx110x)) + ((ax110x) & (!bx110x)));
	assign fx110x = (((!ax108x) & (!bx108x) & (!g231) & (!ax109x) & (!bx109x) & (g234)) + ((!ax108x) & (!bx108x) & (!g231) & (!ax109x) & (bx109x) & (g234)) + ((!ax108x) & (!bx108x) & (!g231) & (ax109x) & (!bx109x) & (g234)) + ((!ax108x) & (!bx108x) & (!g231) & (ax109x) & (bx109x) & (!g234)) + ((!ax108x) & (!bx108x) & (g231) & (!ax109x) & (!bx109x) & (g234)) + ((!ax108x) & (!bx108x) & (g231) & (!ax109x) & (bx109x) & (g234)) + ((!ax108x) & (!bx108x) & (g231) & (ax109x) & (!bx109x) & (g234)) + ((!ax108x) & (!bx108x) & (g231) & (ax109x) & (bx109x) & (!g234)) + ((!ax108x) & (bx108x) & (!g231) & (!ax109x) & (!bx109x) & (g234)) + ((!ax108x) & (bx108x) & (!g231) & (!ax109x) & (bx109x) & (!g234)) + ((!ax108x) & (bx108x) & (!g231) & (ax109x) & (!bx109x) & (!g234)) + ((!ax108x) & (bx108x) & (!g231) & (ax109x) & (bx109x) & (!g234)) + ((!ax108x) & (bx108x) & (g231) & (!ax109x) & (!bx109x) & (g234)) + ((!ax108x) & (bx108x) & (g231) & (!ax109x) & (bx109x) & (g234)) + ((!ax108x) & (bx108x) & (g231) & (ax109x) & (!bx109x) & (g234)) + ((!ax108x) & (bx108x) & (g231) & (ax109x) & (bx109x) & (!g234)) + ((ax108x) & (!bx108x) & (!g231) & (!ax109x) & (!bx109x) & (g234)) + ((ax108x) & (!bx108x) & (!g231) & (!ax109x) & (bx109x) & (!g234)) + ((ax108x) & (!bx108x) & (!g231) & (ax109x) & (!bx109x) & (!g234)) + ((ax108x) & (!bx108x) & (!g231) & (ax109x) & (bx109x) & (!g234)) + ((ax108x) & (!bx108x) & (g231) & (!ax109x) & (!bx109x) & (g234)) + ((ax108x) & (!bx108x) & (g231) & (!ax109x) & (bx109x) & (g234)) + ((ax108x) & (!bx108x) & (g231) & (ax109x) & (!bx109x) & (g234)) + ((ax108x) & (!bx108x) & (g231) & (ax109x) & (bx109x) & (!g234)) + ((ax108x) & (bx108x) & (!g231) & (!ax109x) & (!bx109x) & (g234)) + ((ax108x) & (bx108x) & (!g231) & (!ax109x) & (bx109x) & (!g234)) + ((ax108x) & (bx108x) & (!g231) & (ax109x) & (!bx109x) & (!g234)) + ((ax108x) & (bx108x) & (!g231) & (ax109x) & (bx109x) & (!g234)) + ((ax108x) & (bx108x) & (g231) & (!ax109x) & (!bx109x) & (g234)) + ((ax108x) & (bx108x) & (g231) & (!ax109x) & (bx109x) & (!g234)) + ((ax108x) & (bx108x) & (g231) & (ax109x) & (!bx109x) & (!g234)) + ((ax108x) & (bx108x) & (g231) & (ax109x) & (bx109x) & (!g234)));
	assign g236 = (((ax110x) & (bx110x)));
	assign g237 = (((!ax110x) & (!bx110x)));
	assign g238 = (((!ax108x) & (!bx108x) & (!g231) & (ax109x) & (bx109x) & (!g237)) + ((!ax108x) & (!bx108x) & (g231) & (ax109x) & (bx109x) & (!g237)) + ((!ax108x) & (bx108x) & (!g231) & (!ax109x) & (bx109x) & (!g237)) + ((!ax108x) & (bx108x) & (!g231) & (ax109x) & (!bx109x) & (!g237)) + ((!ax108x) & (bx108x) & (!g231) & (ax109x) & (bx109x) & (!g237)) + ((!ax108x) & (bx108x) & (g231) & (ax109x) & (bx109x) & (!g237)) + ((ax108x) & (!bx108x) & (!g231) & (!ax109x) & (bx109x) & (!g237)) + ((ax108x) & (!bx108x) & (!g231) & (ax109x) & (!bx109x) & (!g237)) + ((ax108x) & (!bx108x) & (!g231) & (ax109x) & (bx109x) & (!g237)) + ((ax108x) & (!bx108x) & (g231) & (ax109x) & (bx109x) & (!g237)) + ((ax108x) & (bx108x) & (!g231) & (!ax109x) & (bx109x) & (!g237)) + ((ax108x) & (bx108x) & (!g231) & (ax109x) & (!bx109x) & (!g237)) + ((ax108x) & (bx108x) & (!g231) & (ax109x) & (bx109x) & (!g237)) + ((ax108x) & (bx108x) & (g231) & (!ax109x) & (bx109x) & (!g237)) + ((ax108x) & (bx108x) & (g231) & (ax109x) & (!bx109x) & (!g237)) + ((ax108x) & (bx108x) & (g231) & (ax109x) & (bx109x) & (!g237)));
	assign fx111x = (((!ax111x) & (!bx111x) & (!g236) & (g238)) + ((!ax111x) & (!bx111x) & (g236) & (!g238)) + ((!ax111x) & (!bx111x) & (g236) & (g238)) + ((!ax111x) & (bx111x) & (!g236) & (!g238)) + ((ax111x) & (!bx111x) & (!g236) & (!g238)) + ((ax111x) & (bx111x) & (!g236) & (g238)) + ((ax111x) & (bx111x) & (g236) & (!g238)) + ((ax111x) & (bx111x) & (g236) & (g238)));
	assign fx112x = (((!ax111x) & (!bx111x) & (!g236) & (!g238) & (!ax112x) & (bx112x)) + ((!ax111x) & (!bx111x) & (!g236) & (!g238) & (ax112x) & (!bx112x)) + ((!ax111x) & (!bx111x) & (!g236) & (g238) & (!ax112x) & (bx112x)) + ((!ax111x) & (!bx111x) & (!g236) & (g238) & (ax112x) & (!bx112x)) + ((!ax111x) & (!bx111x) & (g236) & (!g238) & (!ax112x) & (bx112x)) + ((!ax111x) & (!bx111x) & (g236) & (!g238) & (ax112x) & (!bx112x)) + ((!ax111x) & (!bx111x) & (g236) & (g238) & (!ax112x) & (bx112x)) + ((!ax111x) & (!bx111x) & (g236) & (g238) & (ax112x) & (!bx112x)) + ((!ax111x) & (bx111x) & (!g236) & (!g238) & (!ax112x) & (bx112x)) + ((!ax111x) & (bx111x) & (!g236) & (!g238) & (ax112x) & (!bx112x)) + ((!ax111x) & (bx111x) & (!g236) & (g238) & (!ax112x) & (!bx112x)) + ((!ax111x) & (bx111x) & (!g236) & (g238) & (ax112x) & (bx112x)) + ((!ax111x) & (bx111x) & (g236) & (!g238) & (!ax112x) & (!bx112x)) + ((!ax111x) & (bx111x) & (g236) & (!g238) & (ax112x) & (bx112x)) + ((!ax111x) & (bx111x) & (g236) & (g238) & (!ax112x) & (!bx112x)) + ((!ax111x) & (bx111x) & (g236) & (g238) & (ax112x) & (bx112x)) + ((ax111x) & (!bx111x) & (!g236) & (!g238) & (!ax112x) & (bx112x)) + ((ax111x) & (!bx111x) & (!g236) & (!g238) & (ax112x) & (!bx112x)) + ((ax111x) & (!bx111x) & (!g236) & (g238) & (!ax112x) & (!bx112x)) + ((ax111x) & (!bx111x) & (!g236) & (g238) & (ax112x) & (bx112x)) + ((ax111x) & (!bx111x) & (g236) & (!g238) & (!ax112x) & (!bx112x)) + ((ax111x) & (!bx111x) & (g236) & (!g238) & (ax112x) & (bx112x)) + ((ax111x) & (!bx111x) & (g236) & (g238) & (!ax112x) & (!bx112x)) + ((ax111x) & (!bx111x) & (g236) & (g238) & (ax112x) & (bx112x)) + ((ax111x) & (bx111x) & (!g236) & (!g238) & (!ax112x) & (!bx112x)) + ((ax111x) & (bx111x) & (!g236) & (!g238) & (ax112x) & (bx112x)) + ((ax111x) & (bx111x) & (!g236) & (g238) & (!ax112x) & (!bx112x)) + ((ax111x) & (bx111x) & (!g236) & (g238) & (ax112x) & (bx112x)) + ((ax111x) & (bx111x) & (g236) & (!g238) & (!ax112x) & (!bx112x)) + ((ax111x) & (bx111x) & (g236) & (!g238) & (ax112x) & (bx112x)) + ((ax111x) & (bx111x) & (g236) & (g238) & (!ax112x) & (!bx112x)) + ((ax111x) & (bx111x) & (g236) & (g238) & (ax112x) & (bx112x)));
	assign g241 = (((!ax111x) & (!bx111x) & (!g236) & (!g238) & (!ax112x) & (!bx112x)) + ((!ax111x) & (!bx111x) & (!g236) & (!g238) & (!ax112x) & (bx112x)) + ((!ax111x) & (!bx111x) & (!g236) & (!g238) & (ax112x) & (!bx112x)) + ((!ax111x) & (!bx111x) & (!g236) & (g238) & (!ax112x) & (!bx112x)) + ((!ax111x) & (!bx111x) & (!g236) & (g238) & (!ax112x) & (bx112x)) + ((!ax111x) & (!bx111x) & (!g236) & (g238) & (ax112x) & (!bx112x)) + ((!ax111x) & (!bx111x) & (g236) & (!g238) & (!ax112x) & (!bx112x)) + ((!ax111x) & (!bx111x) & (g236) & (!g238) & (!ax112x) & (bx112x)) + ((!ax111x) & (!bx111x) & (g236) & (!g238) & (ax112x) & (!bx112x)) + ((!ax111x) & (!bx111x) & (g236) & (g238) & (!ax112x) & (!bx112x)) + ((!ax111x) & (!bx111x) & (g236) & (g238) & (!ax112x) & (bx112x)) + ((!ax111x) & (!bx111x) & (g236) & (g238) & (ax112x) & (!bx112x)) + ((!ax111x) & (bx111x) & (!g236) & (!g238) & (!ax112x) & (!bx112x)) + ((!ax111x) & (bx111x) & (!g236) & (!g238) & (!ax112x) & (bx112x)) + ((!ax111x) & (bx111x) & (!g236) & (!g238) & (ax112x) & (!bx112x)) + ((!ax111x) & (bx111x) & (!g236) & (g238) & (!ax112x) & (!bx112x)) + ((!ax111x) & (bx111x) & (g236) & (!g238) & (!ax112x) & (!bx112x)) + ((!ax111x) & (bx111x) & (g236) & (g238) & (!ax112x) & (!bx112x)) + ((ax111x) & (!bx111x) & (!g236) & (!g238) & (!ax112x) & (!bx112x)) + ((ax111x) & (!bx111x) & (!g236) & (!g238) & (!ax112x) & (bx112x)) + ((ax111x) & (!bx111x) & (!g236) & (!g238) & (ax112x) & (!bx112x)) + ((ax111x) & (!bx111x) & (!g236) & (g238) & (!ax112x) & (!bx112x)) + ((ax111x) & (!bx111x) & (g236) & (!g238) & (!ax112x) & (!bx112x)) + ((ax111x) & (!bx111x) & (g236) & (g238) & (!ax112x) & (!bx112x)) + ((ax111x) & (bx111x) & (!g236) & (!g238) & (!ax112x) & (!bx112x)) + ((ax111x) & (bx111x) & (!g236) & (g238) & (!ax112x) & (!bx112x)) + ((ax111x) & (bx111x) & (g236) & (!g238) & (!ax112x) & (!bx112x)) + ((ax111x) & (bx111x) & (g236) & (g238) & (!ax112x) & (!bx112x)));
	assign fx113x = (((!ax113x) & (!bx113x) & (!g241)) + ((!ax113x) & (bx113x) & (g241)) + ((ax113x) & (!bx113x) & (g241)) + ((ax113x) & (bx113x) & (!g241)));
	assign fx114x = (((!ax113x) & (!bx113x) & (!g241) & (!ax114x) & (bx114x)) + ((!ax113x) & (!bx113x) & (!g241) & (ax114x) & (!bx114x)) + ((!ax113x) & (!bx113x) & (g241) & (!ax114x) & (bx114x)) + ((!ax113x) & (!bx113x) & (g241) & (ax114x) & (!bx114x)) + ((!ax113x) & (bx113x) & (!g241) & (!ax114x) & (!bx114x)) + ((!ax113x) & (bx113x) & (!g241) & (ax114x) & (bx114x)) + ((!ax113x) & (bx113x) & (g241) & (!ax114x) & (bx114x)) + ((!ax113x) & (bx113x) & (g241) & (ax114x) & (!bx114x)) + ((ax113x) & (!bx113x) & (!g241) & (!ax114x) & (!bx114x)) + ((ax113x) & (!bx113x) & (!g241) & (ax114x) & (bx114x)) + ((ax113x) & (!bx113x) & (g241) & (!ax114x) & (bx114x)) + ((ax113x) & (!bx113x) & (g241) & (ax114x) & (!bx114x)) + ((ax113x) & (bx113x) & (!g241) & (!ax114x) & (!bx114x)) + ((ax113x) & (bx113x) & (!g241) & (ax114x) & (bx114x)) + ((ax113x) & (bx113x) & (g241) & (!ax114x) & (!bx114x)) + ((ax113x) & (bx113x) & (g241) & (ax114x) & (bx114x)));
	assign g244 = (((!ax115x) & (bx115x)) + ((ax115x) & (!bx115x)));
	assign fx115x = (((!ax113x) & (!bx113x) & (!g241) & (!ax114x) & (!bx114x) & (g244)) + ((!ax113x) & (!bx113x) & (!g241) & (!ax114x) & (bx114x) & (g244)) + ((!ax113x) & (!bx113x) & (!g241) & (ax114x) & (!bx114x) & (g244)) + ((!ax113x) & (!bx113x) & (!g241) & (ax114x) & (bx114x) & (!g244)) + ((!ax113x) & (!bx113x) & (g241) & (!ax114x) & (!bx114x) & (g244)) + ((!ax113x) & (!bx113x) & (g241) & (!ax114x) & (bx114x) & (g244)) + ((!ax113x) & (!bx113x) & (g241) & (ax114x) & (!bx114x) & (g244)) + ((!ax113x) & (!bx113x) & (g241) & (ax114x) & (bx114x) & (!g244)) + ((!ax113x) & (bx113x) & (!g241) & (!ax114x) & (!bx114x) & (g244)) + ((!ax113x) & (bx113x) & (!g241) & (!ax114x) & (bx114x) & (!g244)) + ((!ax113x) & (bx113x) & (!g241) & (ax114x) & (!bx114x) & (!g244)) + ((!ax113x) & (bx113x) & (!g241) & (ax114x) & (bx114x) & (!g244)) + ((!ax113x) & (bx113x) & (g241) & (!ax114x) & (!bx114x) & (g244)) + ((!ax113x) & (bx113x) & (g241) & (!ax114x) & (bx114x) & (g244)) + ((!ax113x) & (bx113x) & (g241) & (ax114x) & (!bx114x) & (g244)) + ((!ax113x) & (bx113x) & (g241) & (ax114x) & (bx114x) & (!g244)) + ((ax113x) & (!bx113x) & (!g241) & (!ax114x) & (!bx114x) & (g244)) + ((ax113x) & (!bx113x) & (!g241) & (!ax114x) & (bx114x) & (!g244)) + ((ax113x) & (!bx113x) & (!g241) & (ax114x) & (!bx114x) & (!g244)) + ((ax113x) & (!bx113x) & (!g241) & (ax114x) & (bx114x) & (!g244)) + ((ax113x) & (!bx113x) & (g241) & (!ax114x) & (!bx114x) & (g244)) + ((ax113x) & (!bx113x) & (g241) & (!ax114x) & (bx114x) & (g244)) + ((ax113x) & (!bx113x) & (g241) & (ax114x) & (!bx114x) & (g244)) + ((ax113x) & (!bx113x) & (g241) & (ax114x) & (bx114x) & (!g244)) + ((ax113x) & (bx113x) & (!g241) & (!ax114x) & (!bx114x) & (g244)) + ((ax113x) & (bx113x) & (!g241) & (!ax114x) & (bx114x) & (!g244)) + ((ax113x) & (bx113x) & (!g241) & (ax114x) & (!bx114x) & (!g244)) + ((ax113x) & (bx113x) & (!g241) & (ax114x) & (bx114x) & (!g244)) + ((ax113x) & (bx113x) & (g241) & (!ax114x) & (!bx114x) & (g244)) + ((ax113x) & (bx113x) & (g241) & (!ax114x) & (bx114x) & (!g244)) + ((ax113x) & (bx113x) & (g241) & (ax114x) & (!bx114x) & (!g244)) + ((ax113x) & (bx113x) & (g241) & (ax114x) & (bx114x) & (!g244)));
	assign g246 = (((ax115x) & (bx115x)));
	assign g247 = (((!ax115x) & (!bx115x)));
	assign g248 = (((!ax113x) & (!bx113x) & (!g241) & (ax114x) & (bx114x) & (!g247)) + ((!ax113x) & (!bx113x) & (g241) & (ax114x) & (bx114x) & (!g247)) + ((!ax113x) & (bx113x) & (!g241) & (!ax114x) & (bx114x) & (!g247)) + ((!ax113x) & (bx113x) & (!g241) & (ax114x) & (!bx114x) & (!g247)) + ((!ax113x) & (bx113x) & (!g241) & (ax114x) & (bx114x) & (!g247)) + ((!ax113x) & (bx113x) & (g241) & (ax114x) & (bx114x) & (!g247)) + ((ax113x) & (!bx113x) & (!g241) & (!ax114x) & (bx114x) & (!g247)) + ((ax113x) & (!bx113x) & (!g241) & (ax114x) & (!bx114x) & (!g247)) + ((ax113x) & (!bx113x) & (!g241) & (ax114x) & (bx114x) & (!g247)) + ((ax113x) & (!bx113x) & (g241) & (ax114x) & (bx114x) & (!g247)) + ((ax113x) & (bx113x) & (!g241) & (!ax114x) & (bx114x) & (!g247)) + ((ax113x) & (bx113x) & (!g241) & (ax114x) & (!bx114x) & (!g247)) + ((ax113x) & (bx113x) & (!g241) & (ax114x) & (bx114x) & (!g247)) + ((ax113x) & (bx113x) & (g241) & (!ax114x) & (bx114x) & (!g247)) + ((ax113x) & (bx113x) & (g241) & (ax114x) & (!bx114x) & (!g247)) + ((ax113x) & (bx113x) & (g241) & (ax114x) & (bx114x) & (!g247)));
	assign fx116x = (((!ax116x) & (!bx116x) & (!g246) & (g248)) + ((!ax116x) & (!bx116x) & (g246) & (!g248)) + ((!ax116x) & (!bx116x) & (g246) & (g248)) + ((!ax116x) & (bx116x) & (!g246) & (!g248)) + ((ax116x) & (!bx116x) & (!g246) & (!g248)) + ((ax116x) & (bx116x) & (!g246) & (g248)) + ((ax116x) & (bx116x) & (g246) & (!g248)) + ((ax116x) & (bx116x) & (g246) & (g248)));
	assign fx117x = (((!ax116x) & (!bx116x) & (!g246) & (!g248) & (!ax117x) & (bx117x)) + ((!ax116x) & (!bx116x) & (!g246) & (!g248) & (ax117x) & (!bx117x)) + ((!ax116x) & (!bx116x) & (!g246) & (g248) & (!ax117x) & (bx117x)) + ((!ax116x) & (!bx116x) & (!g246) & (g248) & (ax117x) & (!bx117x)) + ((!ax116x) & (!bx116x) & (g246) & (!g248) & (!ax117x) & (bx117x)) + ((!ax116x) & (!bx116x) & (g246) & (!g248) & (ax117x) & (!bx117x)) + ((!ax116x) & (!bx116x) & (g246) & (g248) & (!ax117x) & (bx117x)) + ((!ax116x) & (!bx116x) & (g246) & (g248) & (ax117x) & (!bx117x)) + ((!ax116x) & (bx116x) & (!g246) & (!g248) & (!ax117x) & (bx117x)) + ((!ax116x) & (bx116x) & (!g246) & (!g248) & (ax117x) & (!bx117x)) + ((!ax116x) & (bx116x) & (!g246) & (g248) & (!ax117x) & (!bx117x)) + ((!ax116x) & (bx116x) & (!g246) & (g248) & (ax117x) & (bx117x)) + ((!ax116x) & (bx116x) & (g246) & (!g248) & (!ax117x) & (!bx117x)) + ((!ax116x) & (bx116x) & (g246) & (!g248) & (ax117x) & (bx117x)) + ((!ax116x) & (bx116x) & (g246) & (g248) & (!ax117x) & (!bx117x)) + ((!ax116x) & (bx116x) & (g246) & (g248) & (ax117x) & (bx117x)) + ((ax116x) & (!bx116x) & (!g246) & (!g248) & (!ax117x) & (bx117x)) + ((ax116x) & (!bx116x) & (!g246) & (!g248) & (ax117x) & (!bx117x)) + ((ax116x) & (!bx116x) & (!g246) & (g248) & (!ax117x) & (!bx117x)) + ((ax116x) & (!bx116x) & (!g246) & (g248) & (ax117x) & (bx117x)) + ((ax116x) & (!bx116x) & (g246) & (!g248) & (!ax117x) & (!bx117x)) + ((ax116x) & (!bx116x) & (g246) & (!g248) & (ax117x) & (bx117x)) + ((ax116x) & (!bx116x) & (g246) & (g248) & (!ax117x) & (!bx117x)) + ((ax116x) & (!bx116x) & (g246) & (g248) & (ax117x) & (bx117x)) + ((ax116x) & (bx116x) & (!g246) & (!g248) & (!ax117x) & (!bx117x)) + ((ax116x) & (bx116x) & (!g246) & (!g248) & (ax117x) & (bx117x)) + ((ax116x) & (bx116x) & (!g246) & (g248) & (!ax117x) & (!bx117x)) + ((ax116x) & (bx116x) & (!g246) & (g248) & (ax117x) & (bx117x)) + ((ax116x) & (bx116x) & (g246) & (!g248) & (!ax117x) & (!bx117x)) + ((ax116x) & (bx116x) & (g246) & (!g248) & (ax117x) & (bx117x)) + ((ax116x) & (bx116x) & (g246) & (g248) & (!ax117x) & (!bx117x)) + ((ax116x) & (bx116x) & (g246) & (g248) & (ax117x) & (bx117x)));
	assign g251 = (((!ax116x) & (!bx116x) & (!g246) & (!g248) & (!ax117x) & (!bx117x)) + ((!ax116x) & (!bx116x) & (!g246) & (!g248) & (!ax117x) & (bx117x)) + ((!ax116x) & (!bx116x) & (!g246) & (!g248) & (ax117x) & (!bx117x)) + ((!ax116x) & (!bx116x) & (!g246) & (g248) & (!ax117x) & (!bx117x)) + ((!ax116x) & (!bx116x) & (!g246) & (g248) & (!ax117x) & (bx117x)) + ((!ax116x) & (!bx116x) & (!g246) & (g248) & (ax117x) & (!bx117x)) + ((!ax116x) & (!bx116x) & (g246) & (!g248) & (!ax117x) & (!bx117x)) + ((!ax116x) & (!bx116x) & (g246) & (!g248) & (!ax117x) & (bx117x)) + ((!ax116x) & (!bx116x) & (g246) & (!g248) & (ax117x) & (!bx117x)) + ((!ax116x) & (!bx116x) & (g246) & (g248) & (!ax117x) & (!bx117x)) + ((!ax116x) & (!bx116x) & (g246) & (g248) & (!ax117x) & (bx117x)) + ((!ax116x) & (!bx116x) & (g246) & (g248) & (ax117x) & (!bx117x)) + ((!ax116x) & (bx116x) & (!g246) & (!g248) & (!ax117x) & (!bx117x)) + ((!ax116x) & (bx116x) & (!g246) & (!g248) & (!ax117x) & (bx117x)) + ((!ax116x) & (bx116x) & (!g246) & (!g248) & (ax117x) & (!bx117x)) + ((!ax116x) & (bx116x) & (!g246) & (g248) & (!ax117x) & (!bx117x)) + ((!ax116x) & (bx116x) & (g246) & (!g248) & (!ax117x) & (!bx117x)) + ((!ax116x) & (bx116x) & (g246) & (g248) & (!ax117x) & (!bx117x)) + ((ax116x) & (!bx116x) & (!g246) & (!g248) & (!ax117x) & (!bx117x)) + ((ax116x) & (!bx116x) & (!g246) & (!g248) & (!ax117x) & (bx117x)) + ((ax116x) & (!bx116x) & (!g246) & (!g248) & (ax117x) & (!bx117x)) + ((ax116x) & (!bx116x) & (!g246) & (g248) & (!ax117x) & (!bx117x)) + ((ax116x) & (!bx116x) & (g246) & (!g248) & (!ax117x) & (!bx117x)) + ((ax116x) & (!bx116x) & (g246) & (g248) & (!ax117x) & (!bx117x)) + ((ax116x) & (bx116x) & (!g246) & (!g248) & (!ax117x) & (!bx117x)) + ((ax116x) & (bx116x) & (!g246) & (g248) & (!ax117x) & (!bx117x)) + ((ax116x) & (bx116x) & (g246) & (!g248) & (!ax117x) & (!bx117x)) + ((ax116x) & (bx116x) & (g246) & (g248) & (!ax117x) & (!bx117x)));
	assign fx118x = (((!ax118x) & (!bx118x) & (!g251)) + ((!ax118x) & (bx118x) & (g251)) + ((ax118x) & (!bx118x) & (g251)) + ((ax118x) & (bx118x) & (!g251)));
	assign fx119x = (((!ax118x) & (!bx118x) & (!g251) & (!ax119x) & (bx119x)) + ((!ax118x) & (!bx118x) & (!g251) & (ax119x) & (!bx119x)) + ((!ax118x) & (!bx118x) & (g251) & (!ax119x) & (bx119x)) + ((!ax118x) & (!bx118x) & (g251) & (ax119x) & (!bx119x)) + ((!ax118x) & (bx118x) & (!g251) & (!ax119x) & (!bx119x)) + ((!ax118x) & (bx118x) & (!g251) & (ax119x) & (bx119x)) + ((!ax118x) & (bx118x) & (g251) & (!ax119x) & (bx119x)) + ((!ax118x) & (bx118x) & (g251) & (ax119x) & (!bx119x)) + ((ax118x) & (!bx118x) & (!g251) & (!ax119x) & (!bx119x)) + ((ax118x) & (!bx118x) & (!g251) & (ax119x) & (bx119x)) + ((ax118x) & (!bx118x) & (g251) & (!ax119x) & (bx119x)) + ((ax118x) & (!bx118x) & (g251) & (ax119x) & (!bx119x)) + ((ax118x) & (bx118x) & (!g251) & (!ax119x) & (!bx119x)) + ((ax118x) & (bx118x) & (!g251) & (ax119x) & (bx119x)) + ((ax118x) & (bx118x) & (g251) & (!ax119x) & (!bx119x)) + ((ax118x) & (bx118x) & (g251) & (ax119x) & (bx119x)));
	assign g254 = (((!ax120x) & (bx120x)) + ((ax120x) & (!bx120x)));
	assign fx120x = (((!ax118x) & (!bx118x) & (!g251) & (!ax119x) & (!bx119x) & (g254)) + ((!ax118x) & (!bx118x) & (!g251) & (!ax119x) & (bx119x) & (g254)) + ((!ax118x) & (!bx118x) & (!g251) & (ax119x) & (!bx119x) & (g254)) + ((!ax118x) & (!bx118x) & (!g251) & (ax119x) & (bx119x) & (!g254)) + ((!ax118x) & (!bx118x) & (g251) & (!ax119x) & (!bx119x) & (g254)) + ((!ax118x) & (!bx118x) & (g251) & (!ax119x) & (bx119x) & (g254)) + ((!ax118x) & (!bx118x) & (g251) & (ax119x) & (!bx119x) & (g254)) + ((!ax118x) & (!bx118x) & (g251) & (ax119x) & (bx119x) & (!g254)) + ((!ax118x) & (bx118x) & (!g251) & (!ax119x) & (!bx119x) & (g254)) + ((!ax118x) & (bx118x) & (!g251) & (!ax119x) & (bx119x) & (!g254)) + ((!ax118x) & (bx118x) & (!g251) & (ax119x) & (!bx119x) & (!g254)) + ((!ax118x) & (bx118x) & (!g251) & (ax119x) & (bx119x) & (!g254)) + ((!ax118x) & (bx118x) & (g251) & (!ax119x) & (!bx119x) & (g254)) + ((!ax118x) & (bx118x) & (g251) & (!ax119x) & (bx119x) & (g254)) + ((!ax118x) & (bx118x) & (g251) & (ax119x) & (!bx119x) & (g254)) + ((!ax118x) & (bx118x) & (g251) & (ax119x) & (bx119x) & (!g254)) + ((ax118x) & (!bx118x) & (!g251) & (!ax119x) & (!bx119x) & (g254)) + ((ax118x) & (!bx118x) & (!g251) & (!ax119x) & (bx119x) & (!g254)) + ((ax118x) & (!bx118x) & (!g251) & (ax119x) & (!bx119x) & (!g254)) + ((ax118x) & (!bx118x) & (!g251) & (ax119x) & (bx119x) & (!g254)) + ((ax118x) & (!bx118x) & (g251) & (!ax119x) & (!bx119x) & (g254)) + ((ax118x) & (!bx118x) & (g251) & (!ax119x) & (bx119x) & (g254)) + ((ax118x) & (!bx118x) & (g251) & (ax119x) & (!bx119x) & (g254)) + ((ax118x) & (!bx118x) & (g251) & (ax119x) & (bx119x) & (!g254)) + ((ax118x) & (bx118x) & (!g251) & (!ax119x) & (!bx119x) & (g254)) + ((ax118x) & (bx118x) & (!g251) & (!ax119x) & (bx119x) & (!g254)) + ((ax118x) & (bx118x) & (!g251) & (ax119x) & (!bx119x) & (!g254)) + ((ax118x) & (bx118x) & (!g251) & (ax119x) & (bx119x) & (!g254)) + ((ax118x) & (bx118x) & (g251) & (!ax119x) & (!bx119x) & (g254)) + ((ax118x) & (bx118x) & (g251) & (!ax119x) & (bx119x) & (!g254)) + ((ax118x) & (bx118x) & (g251) & (ax119x) & (!bx119x) & (!g254)) + ((ax118x) & (bx118x) & (g251) & (ax119x) & (bx119x) & (!g254)));
	assign g256 = (((ax120x) & (bx120x)));
	assign g257 = (((!ax120x) & (!bx120x)));
	assign g258 = (((!ax118x) & (!bx118x) & (!g251) & (ax119x) & (bx119x) & (!g257)) + ((!ax118x) & (!bx118x) & (g251) & (ax119x) & (bx119x) & (!g257)) + ((!ax118x) & (bx118x) & (!g251) & (!ax119x) & (bx119x) & (!g257)) + ((!ax118x) & (bx118x) & (!g251) & (ax119x) & (!bx119x) & (!g257)) + ((!ax118x) & (bx118x) & (!g251) & (ax119x) & (bx119x) & (!g257)) + ((!ax118x) & (bx118x) & (g251) & (ax119x) & (bx119x) & (!g257)) + ((ax118x) & (!bx118x) & (!g251) & (!ax119x) & (bx119x) & (!g257)) + ((ax118x) & (!bx118x) & (!g251) & (ax119x) & (!bx119x) & (!g257)) + ((ax118x) & (!bx118x) & (!g251) & (ax119x) & (bx119x) & (!g257)) + ((ax118x) & (!bx118x) & (g251) & (ax119x) & (bx119x) & (!g257)) + ((ax118x) & (bx118x) & (!g251) & (!ax119x) & (bx119x) & (!g257)) + ((ax118x) & (bx118x) & (!g251) & (ax119x) & (!bx119x) & (!g257)) + ((ax118x) & (bx118x) & (!g251) & (ax119x) & (bx119x) & (!g257)) + ((ax118x) & (bx118x) & (g251) & (!ax119x) & (bx119x) & (!g257)) + ((ax118x) & (bx118x) & (g251) & (ax119x) & (!bx119x) & (!g257)) + ((ax118x) & (bx118x) & (g251) & (ax119x) & (bx119x) & (!g257)));
	assign fx121x = (((!ax121x) & (!bx121x) & (!g256) & (g258)) + ((!ax121x) & (!bx121x) & (g256) & (!g258)) + ((!ax121x) & (!bx121x) & (g256) & (g258)) + ((!ax121x) & (bx121x) & (!g256) & (!g258)) + ((ax121x) & (!bx121x) & (!g256) & (!g258)) + ((ax121x) & (bx121x) & (!g256) & (g258)) + ((ax121x) & (bx121x) & (g256) & (!g258)) + ((ax121x) & (bx121x) & (g256) & (g258)));
	assign fx122x = (((!ax121x) & (!bx121x) & (!g256) & (!g258) & (!ax122x) & (bx122x)) + ((!ax121x) & (!bx121x) & (!g256) & (!g258) & (ax122x) & (!bx122x)) + ((!ax121x) & (!bx121x) & (!g256) & (g258) & (!ax122x) & (bx122x)) + ((!ax121x) & (!bx121x) & (!g256) & (g258) & (ax122x) & (!bx122x)) + ((!ax121x) & (!bx121x) & (g256) & (!g258) & (!ax122x) & (bx122x)) + ((!ax121x) & (!bx121x) & (g256) & (!g258) & (ax122x) & (!bx122x)) + ((!ax121x) & (!bx121x) & (g256) & (g258) & (!ax122x) & (bx122x)) + ((!ax121x) & (!bx121x) & (g256) & (g258) & (ax122x) & (!bx122x)) + ((!ax121x) & (bx121x) & (!g256) & (!g258) & (!ax122x) & (bx122x)) + ((!ax121x) & (bx121x) & (!g256) & (!g258) & (ax122x) & (!bx122x)) + ((!ax121x) & (bx121x) & (!g256) & (g258) & (!ax122x) & (!bx122x)) + ((!ax121x) & (bx121x) & (!g256) & (g258) & (ax122x) & (bx122x)) + ((!ax121x) & (bx121x) & (g256) & (!g258) & (!ax122x) & (!bx122x)) + ((!ax121x) & (bx121x) & (g256) & (!g258) & (ax122x) & (bx122x)) + ((!ax121x) & (bx121x) & (g256) & (g258) & (!ax122x) & (!bx122x)) + ((!ax121x) & (bx121x) & (g256) & (g258) & (ax122x) & (bx122x)) + ((ax121x) & (!bx121x) & (!g256) & (!g258) & (!ax122x) & (bx122x)) + ((ax121x) & (!bx121x) & (!g256) & (!g258) & (ax122x) & (!bx122x)) + ((ax121x) & (!bx121x) & (!g256) & (g258) & (!ax122x) & (!bx122x)) + ((ax121x) & (!bx121x) & (!g256) & (g258) & (ax122x) & (bx122x)) + ((ax121x) & (!bx121x) & (g256) & (!g258) & (!ax122x) & (!bx122x)) + ((ax121x) & (!bx121x) & (g256) & (!g258) & (ax122x) & (bx122x)) + ((ax121x) & (!bx121x) & (g256) & (g258) & (!ax122x) & (!bx122x)) + ((ax121x) & (!bx121x) & (g256) & (g258) & (ax122x) & (bx122x)) + ((ax121x) & (bx121x) & (!g256) & (!g258) & (!ax122x) & (!bx122x)) + ((ax121x) & (bx121x) & (!g256) & (!g258) & (ax122x) & (bx122x)) + ((ax121x) & (bx121x) & (!g256) & (g258) & (!ax122x) & (!bx122x)) + ((ax121x) & (bx121x) & (!g256) & (g258) & (ax122x) & (bx122x)) + ((ax121x) & (bx121x) & (g256) & (!g258) & (!ax122x) & (!bx122x)) + ((ax121x) & (bx121x) & (g256) & (!g258) & (ax122x) & (bx122x)) + ((ax121x) & (bx121x) & (g256) & (g258) & (!ax122x) & (!bx122x)) + ((ax121x) & (bx121x) & (g256) & (g258) & (ax122x) & (bx122x)));
	assign g261 = (((!ax121x) & (!bx121x) & (!g256) & (!g258) & (!ax122x) & (!bx122x)) + ((!ax121x) & (!bx121x) & (!g256) & (!g258) & (!ax122x) & (bx122x)) + ((!ax121x) & (!bx121x) & (!g256) & (!g258) & (ax122x) & (!bx122x)) + ((!ax121x) & (!bx121x) & (!g256) & (g258) & (!ax122x) & (!bx122x)) + ((!ax121x) & (!bx121x) & (!g256) & (g258) & (!ax122x) & (bx122x)) + ((!ax121x) & (!bx121x) & (!g256) & (g258) & (ax122x) & (!bx122x)) + ((!ax121x) & (!bx121x) & (g256) & (!g258) & (!ax122x) & (!bx122x)) + ((!ax121x) & (!bx121x) & (g256) & (!g258) & (!ax122x) & (bx122x)) + ((!ax121x) & (!bx121x) & (g256) & (!g258) & (ax122x) & (!bx122x)) + ((!ax121x) & (!bx121x) & (g256) & (g258) & (!ax122x) & (!bx122x)) + ((!ax121x) & (!bx121x) & (g256) & (g258) & (!ax122x) & (bx122x)) + ((!ax121x) & (!bx121x) & (g256) & (g258) & (ax122x) & (!bx122x)) + ((!ax121x) & (bx121x) & (!g256) & (!g258) & (!ax122x) & (!bx122x)) + ((!ax121x) & (bx121x) & (!g256) & (!g258) & (!ax122x) & (bx122x)) + ((!ax121x) & (bx121x) & (!g256) & (!g258) & (ax122x) & (!bx122x)) + ((!ax121x) & (bx121x) & (!g256) & (g258) & (!ax122x) & (!bx122x)) + ((!ax121x) & (bx121x) & (g256) & (!g258) & (!ax122x) & (!bx122x)) + ((!ax121x) & (bx121x) & (g256) & (g258) & (!ax122x) & (!bx122x)) + ((ax121x) & (!bx121x) & (!g256) & (!g258) & (!ax122x) & (!bx122x)) + ((ax121x) & (!bx121x) & (!g256) & (!g258) & (!ax122x) & (bx122x)) + ((ax121x) & (!bx121x) & (!g256) & (!g258) & (ax122x) & (!bx122x)) + ((ax121x) & (!bx121x) & (!g256) & (g258) & (!ax122x) & (!bx122x)) + ((ax121x) & (!bx121x) & (g256) & (!g258) & (!ax122x) & (!bx122x)) + ((ax121x) & (!bx121x) & (g256) & (g258) & (!ax122x) & (!bx122x)) + ((ax121x) & (bx121x) & (!g256) & (!g258) & (!ax122x) & (!bx122x)) + ((ax121x) & (bx121x) & (!g256) & (g258) & (!ax122x) & (!bx122x)) + ((ax121x) & (bx121x) & (g256) & (!g258) & (!ax122x) & (!bx122x)) + ((ax121x) & (bx121x) & (g256) & (g258) & (!ax122x) & (!bx122x)));
	assign fx123x = (((!ax123x) & (!bx123x) & (!g261)) + ((!ax123x) & (bx123x) & (g261)) + ((ax123x) & (!bx123x) & (g261)) + ((ax123x) & (bx123x) & (!g261)));
	assign fx124x = (((!ax123x) & (!bx123x) & (!g261) & (!ax124x) & (bx124x)) + ((!ax123x) & (!bx123x) & (!g261) & (ax124x) & (!bx124x)) + ((!ax123x) & (!bx123x) & (g261) & (!ax124x) & (bx124x)) + ((!ax123x) & (!bx123x) & (g261) & (ax124x) & (!bx124x)) + ((!ax123x) & (bx123x) & (!g261) & (!ax124x) & (!bx124x)) + ((!ax123x) & (bx123x) & (!g261) & (ax124x) & (bx124x)) + ((!ax123x) & (bx123x) & (g261) & (!ax124x) & (bx124x)) + ((!ax123x) & (bx123x) & (g261) & (ax124x) & (!bx124x)) + ((ax123x) & (!bx123x) & (!g261) & (!ax124x) & (!bx124x)) + ((ax123x) & (!bx123x) & (!g261) & (ax124x) & (bx124x)) + ((ax123x) & (!bx123x) & (g261) & (!ax124x) & (bx124x)) + ((ax123x) & (!bx123x) & (g261) & (ax124x) & (!bx124x)) + ((ax123x) & (bx123x) & (!g261) & (!ax124x) & (!bx124x)) + ((ax123x) & (bx123x) & (!g261) & (ax124x) & (bx124x)) + ((ax123x) & (bx123x) & (g261) & (!ax124x) & (!bx124x)) + ((ax123x) & (bx123x) & (g261) & (ax124x) & (bx124x)));
	assign g264 = (((!ax125x) & (bx125x)) + ((ax125x) & (!bx125x)));
	assign fx125x = (((!ax123x) & (!bx123x) & (!g261) & (!ax124x) & (!bx124x) & (g264)) + ((!ax123x) & (!bx123x) & (!g261) & (!ax124x) & (bx124x) & (g264)) + ((!ax123x) & (!bx123x) & (!g261) & (ax124x) & (!bx124x) & (g264)) + ((!ax123x) & (!bx123x) & (!g261) & (ax124x) & (bx124x) & (!g264)) + ((!ax123x) & (!bx123x) & (g261) & (!ax124x) & (!bx124x) & (g264)) + ((!ax123x) & (!bx123x) & (g261) & (!ax124x) & (bx124x) & (g264)) + ((!ax123x) & (!bx123x) & (g261) & (ax124x) & (!bx124x) & (g264)) + ((!ax123x) & (!bx123x) & (g261) & (ax124x) & (bx124x) & (!g264)) + ((!ax123x) & (bx123x) & (!g261) & (!ax124x) & (!bx124x) & (g264)) + ((!ax123x) & (bx123x) & (!g261) & (!ax124x) & (bx124x) & (!g264)) + ((!ax123x) & (bx123x) & (!g261) & (ax124x) & (!bx124x) & (!g264)) + ((!ax123x) & (bx123x) & (!g261) & (ax124x) & (bx124x) & (!g264)) + ((!ax123x) & (bx123x) & (g261) & (!ax124x) & (!bx124x) & (g264)) + ((!ax123x) & (bx123x) & (g261) & (!ax124x) & (bx124x) & (g264)) + ((!ax123x) & (bx123x) & (g261) & (ax124x) & (!bx124x) & (g264)) + ((!ax123x) & (bx123x) & (g261) & (ax124x) & (bx124x) & (!g264)) + ((ax123x) & (!bx123x) & (!g261) & (!ax124x) & (!bx124x) & (g264)) + ((ax123x) & (!bx123x) & (!g261) & (!ax124x) & (bx124x) & (!g264)) + ((ax123x) & (!bx123x) & (!g261) & (ax124x) & (!bx124x) & (!g264)) + ((ax123x) & (!bx123x) & (!g261) & (ax124x) & (bx124x) & (!g264)) + ((ax123x) & (!bx123x) & (g261) & (!ax124x) & (!bx124x) & (g264)) + ((ax123x) & (!bx123x) & (g261) & (!ax124x) & (bx124x) & (g264)) + ((ax123x) & (!bx123x) & (g261) & (ax124x) & (!bx124x) & (g264)) + ((ax123x) & (!bx123x) & (g261) & (ax124x) & (bx124x) & (!g264)) + ((ax123x) & (bx123x) & (!g261) & (!ax124x) & (!bx124x) & (g264)) + ((ax123x) & (bx123x) & (!g261) & (!ax124x) & (bx124x) & (!g264)) + ((ax123x) & (bx123x) & (!g261) & (ax124x) & (!bx124x) & (!g264)) + ((ax123x) & (bx123x) & (!g261) & (ax124x) & (bx124x) & (!g264)) + ((ax123x) & (bx123x) & (g261) & (!ax124x) & (!bx124x) & (g264)) + ((ax123x) & (bx123x) & (g261) & (!ax124x) & (bx124x) & (!g264)) + ((ax123x) & (bx123x) & (g261) & (ax124x) & (!bx124x) & (!g264)) + ((ax123x) & (bx123x) & (g261) & (ax124x) & (bx124x) & (!g264)));
	assign g266 = (((ax125x) & (bx125x)));
	assign g267 = (((!ax125x) & (!bx125x)));
	assign g268 = (((!ax123x) & (!bx123x) & (!g261) & (ax124x) & (bx124x) & (!g267)) + ((!ax123x) & (!bx123x) & (g261) & (ax124x) & (bx124x) & (!g267)) + ((!ax123x) & (bx123x) & (!g261) & (!ax124x) & (bx124x) & (!g267)) + ((!ax123x) & (bx123x) & (!g261) & (ax124x) & (!bx124x) & (!g267)) + ((!ax123x) & (bx123x) & (!g261) & (ax124x) & (bx124x) & (!g267)) + ((!ax123x) & (bx123x) & (g261) & (ax124x) & (bx124x) & (!g267)) + ((ax123x) & (!bx123x) & (!g261) & (!ax124x) & (bx124x) & (!g267)) + ((ax123x) & (!bx123x) & (!g261) & (ax124x) & (!bx124x) & (!g267)) + ((ax123x) & (!bx123x) & (!g261) & (ax124x) & (bx124x) & (!g267)) + ((ax123x) & (!bx123x) & (g261) & (ax124x) & (bx124x) & (!g267)) + ((ax123x) & (bx123x) & (!g261) & (!ax124x) & (bx124x) & (!g267)) + ((ax123x) & (bx123x) & (!g261) & (ax124x) & (!bx124x) & (!g267)) + ((ax123x) & (bx123x) & (!g261) & (ax124x) & (bx124x) & (!g267)) + ((ax123x) & (bx123x) & (g261) & (!ax124x) & (bx124x) & (!g267)) + ((ax123x) & (bx123x) & (g261) & (ax124x) & (!bx124x) & (!g267)) + ((ax123x) & (bx123x) & (g261) & (ax124x) & (bx124x) & (!g267)));
	assign fx126x = (((!ax126x) & (!bx126x) & (!g266) & (g268)) + ((!ax126x) & (!bx126x) & (g266) & (!g268)) + ((!ax126x) & (!bx126x) & (g266) & (g268)) + ((!ax126x) & (bx126x) & (!g266) & (!g268)) + ((ax126x) & (!bx126x) & (!g266) & (!g268)) + ((ax126x) & (bx126x) & (!g266) & (g268)) + ((ax126x) & (bx126x) & (g266) & (!g268)) + ((ax126x) & (bx126x) & (g266) & (g268)));
	assign fx127x = (((!ax126x) & (!bx126x) & (!g266) & (!g268) & (!ax127x) & (bx127x)) + ((!ax126x) & (!bx126x) & (!g266) & (!g268) & (ax127x) & (!bx127x)) + ((!ax126x) & (!bx126x) & (!g266) & (g268) & (!ax127x) & (bx127x)) + ((!ax126x) & (!bx126x) & (!g266) & (g268) & (ax127x) & (!bx127x)) + ((!ax126x) & (!bx126x) & (g266) & (!g268) & (!ax127x) & (bx127x)) + ((!ax126x) & (!bx126x) & (g266) & (!g268) & (ax127x) & (!bx127x)) + ((!ax126x) & (!bx126x) & (g266) & (g268) & (!ax127x) & (bx127x)) + ((!ax126x) & (!bx126x) & (g266) & (g268) & (ax127x) & (!bx127x)) + ((!ax126x) & (bx126x) & (!g266) & (!g268) & (!ax127x) & (bx127x)) + ((!ax126x) & (bx126x) & (!g266) & (!g268) & (ax127x) & (!bx127x)) + ((!ax126x) & (bx126x) & (!g266) & (g268) & (!ax127x) & (!bx127x)) + ((!ax126x) & (bx126x) & (!g266) & (g268) & (ax127x) & (bx127x)) + ((!ax126x) & (bx126x) & (g266) & (!g268) & (!ax127x) & (!bx127x)) + ((!ax126x) & (bx126x) & (g266) & (!g268) & (ax127x) & (bx127x)) + ((!ax126x) & (bx126x) & (g266) & (g268) & (!ax127x) & (!bx127x)) + ((!ax126x) & (bx126x) & (g266) & (g268) & (ax127x) & (bx127x)) + ((ax126x) & (!bx126x) & (!g266) & (!g268) & (!ax127x) & (bx127x)) + ((ax126x) & (!bx126x) & (!g266) & (!g268) & (ax127x) & (!bx127x)) + ((ax126x) & (!bx126x) & (!g266) & (g268) & (!ax127x) & (!bx127x)) + ((ax126x) & (!bx126x) & (!g266) & (g268) & (ax127x) & (bx127x)) + ((ax126x) & (!bx126x) & (g266) & (!g268) & (!ax127x) & (!bx127x)) + ((ax126x) & (!bx126x) & (g266) & (!g268) & (ax127x) & (bx127x)) + ((ax126x) & (!bx126x) & (g266) & (g268) & (!ax127x) & (!bx127x)) + ((ax126x) & (!bx126x) & (g266) & (g268) & (ax127x) & (bx127x)) + ((ax126x) & (bx126x) & (!g266) & (!g268) & (!ax127x) & (!bx127x)) + ((ax126x) & (bx126x) & (!g266) & (!g268) & (ax127x) & (bx127x)) + ((ax126x) & (bx126x) & (!g266) & (g268) & (!ax127x) & (!bx127x)) + ((ax126x) & (bx126x) & (!g266) & (g268) & (ax127x) & (bx127x)) + ((ax126x) & (bx126x) & (g266) & (!g268) & (!ax127x) & (!bx127x)) + ((ax126x) & (bx126x) & (g266) & (!g268) & (ax127x) & (bx127x)) + ((ax126x) & (bx126x) & (g266) & (g268) & (!ax127x) & (!bx127x)) + ((ax126x) & (bx126x) & (g266) & (g268) & (ax127x) & (bx127x)));
	assign cOut = (((!ax126x) & (!bx126x) & (!g266) & (!g268) & (ax127x) & (bx127x)) + ((!ax126x) & (!bx126x) & (!g266) & (g268) & (ax127x) & (bx127x)) + ((!ax126x) & (!bx126x) & (g266) & (!g268) & (ax127x) & (bx127x)) + ((!ax126x) & (!bx126x) & (g266) & (g268) & (ax127x) & (bx127x)) + ((!ax126x) & (bx126x) & (!g266) & (!g268) & (ax127x) & (bx127x)) + ((!ax126x) & (bx126x) & (!g266) & (g268) & (!ax127x) & (bx127x)) + ((!ax126x) & (bx126x) & (!g266) & (g268) & (ax127x) & (!bx127x)) + ((!ax126x) & (bx126x) & (!g266) & (g268) & (ax127x) & (bx127x)) + ((!ax126x) & (bx126x) & (g266) & (!g268) & (!ax127x) & (bx127x)) + ((!ax126x) & (bx126x) & (g266) & (!g268) & (ax127x) & (!bx127x)) + ((!ax126x) & (bx126x) & (g266) & (!g268) & (ax127x) & (bx127x)) + ((!ax126x) & (bx126x) & (g266) & (g268) & (!ax127x) & (bx127x)) + ((!ax126x) & (bx126x) & (g266) & (g268) & (ax127x) & (!bx127x)) + ((!ax126x) & (bx126x) & (g266) & (g268) & (ax127x) & (bx127x)) + ((ax126x) & (!bx126x) & (!g266) & (!g268) & (ax127x) & (bx127x)) + ((ax126x) & (!bx126x) & (!g266) & (g268) & (!ax127x) & (bx127x)) + ((ax126x) & (!bx126x) & (!g266) & (g268) & (ax127x) & (!bx127x)) + ((ax126x) & (!bx126x) & (!g266) & (g268) & (ax127x) & (bx127x)) + ((ax126x) & (!bx126x) & (g266) & (!g268) & (!ax127x) & (bx127x)) + ((ax126x) & (!bx126x) & (g266) & (!g268) & (ax127x) & (!bx127x)) + ((ax126x) & (!bx126x) & (g266) & (!g268) & (ax127x) & (bx127x)) + ((ax126x) & (!bx126x) & (g266) & (g268) & (!ax127x) & (bx127x)) + ((ax126x) & (!bx126x) & (g266) & (g268) & (ax127x) & (!bx127x)) + ((ax126x) & (!bx126x) & (g266) & (g268) & (ax127x) & (bx127x)) + ((ax126x) & (bx126x) & (!g266) & (!g268) & (!ax127x) & (bx127x)) + ((ax126x) & (bx126x) & (!g266) & (!g268) & (ax127x) & (!bx127x)) + ((ax126x) & (bx126x) & (!g266) & (!g268) & (ax127x) & (bx127x)) + ((ax126x) & (bx126x) & (!g266) & (g268) & (!ax127x) & (bx127x)) + ((ax126x) & (bx126x) & (!g266) & (g268) & (ax127x) & (!bx127x)) + ((ax126x) & (bx126x) & (!g266) & (g268) & (ax127x) & (bx127x)) + ((ax126x) & (bx126x) & (g266) & (!g268) & (!ax127x) & (bx127x)) + ((ax126x) & (bx126x) & (g266) & (!g268) & (ax127x) & (!bx127x)) + ((ax126x) & (bx126x) & (g266) & (!g268) & (ax127x) & (bx127x)) + ((ax126x) & (bx126x) & (g266) & (g268) & (!ax127x) & (bx127x)) + ((ax126x) & (bx126x) & (g266) & (g268) & (ax127x) & (!bx127x)) + ((ax126x) & (bx126x) & (g266) & (g268) & (ax127x) & (bx127x)));

endmodule