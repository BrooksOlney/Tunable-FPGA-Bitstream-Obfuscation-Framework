module ks_ex5p_qmap_map (sk, i_4_, i_5_, i_6_, i_7_, i_3_, i_1_, i_0_, i_2_, o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_, o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_, o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_, o_41_, o_42_, o_43_, o_44_, o_45_, o_46_, o_47_, o_48_, o_49_, o_50_, o_51_, o_52_, o_53_, o_54_, o_55_, o_56_, o_57_, o_58_, o_59_, o_60_, o_61_, o_62_);

	input i_4_;
	input i_5_;
	input i_6_;
	input i_7_;
	input i_3_;
	input i_1_;
	input i_0_;
	input i_2_;
	output o_0_;
	output o_1_;
	output o_2_;
	output o_3_;
	output o_4_;
	output o_5_;
	output o_6_;
	output o_7_;
	output o_8_;
	output o_9_;
	output o_10_;
	output o_11_;
	output o_12_;
	output o_13_;
	output o_14_;
	output o_15_;
	output o_16_;
	output o_17_;
	output o_18_;
	output o_19_;
	output o_20_;
	output o_21_;
	output o_22_;
	output o_23_;
	output o_24_;
	output o_25_;
	output o_26_;
	output o_27_;
	output o_28_;
	output o_29_;
	output o_30_;
	output o_31_;
	output o_32_;
	output o_33_;
	output o_34_;
	output o_35_;
	output o_36_;
	output o_37_;
	output o_38_;
	output o_39_;
	output o_40_;
	output o_41_;
	output o_42_;
	output o_43_;
	output o_44_;
	output o_45_;
	output o_46_;
	output o_47_;
	output o_48_;
	output o_49_;
	output o_50_;
	output o_51_;
	output o_52_;
	output o_53_;
	output o_54_;
	output o_55_;
	output o_56_;
	output o_57_;
	output o_58_;
	output o_59_;
	output o_60_;
	output o_61_;
	output o_62_;

	input [127 : 0] sk /* synthesis noprune */;


	wire g1, g3, g5, g7, g10, g14, g18, g20, g22, g24, g26, g28, g30, g32, g33, g34, g35, g37, g40, g41, g42;
	wire g45, g46, g47, g48, g49, g51, g52, g53, g365, g92, g94, g121, g122, g124, g152, g165, g175, g188, g194, g207, g214;
	wire g215, g223, g224, g235, g236, g237, g239, g247, g257, g262, g270, g276, g281, g288, g291, g298, g300, g303, g307, g2, g4;
	wire g6, g8, g9, g12, g13, g15, g16, g17, g19, g21, g23, g25, g27, g29, g31, g36, g38, g39, g44, g50, g54;
	wire g55, g56, g57, g58, g59, g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g70, g71, g72, g73, g74, g75;
	wire g76, g77, g78, g79, g80, g81, g82, g83, g354, g84, g85, g86, g87, g88, g89, g90, g91, g93, g95, g96, g97;
	wire g98, g99, g100, g101, g102, g103, g104, g105, g106, g107, g108, g109, g110, g111, g112, g113, g114, g115, g116, g117, g118;
	wire g119, g120, g123, g125, g126, g127, g128, g129, g130, g131, g132, g133, g134, g135, g310, g136, g137, g138, g139, g140, g141;
	wire g142, g143, g144, g145, g146, g147, g148, g149, g150, g343, g333, g151, g153, g154, g155, g156, g157, g158, g159, g160, g161;
	wire g162, g163, g164, g166, g167, g168, g169, g170, g171, g172, g173, g174, g176, g177, g178, g179, g180, g181, g182, g183, g184;
	wire g185, g186, g187, g189, g190, g191, g192, g193, g322, g195, g196, g197, g198, g199, g200, g201, g202, g203, g204, g205, g206;
	wire g311, g208, g209, g210, g211, g212, g213, g216, g217, g218, g219, g220, g221, g222, g225, g226, g227, g228, g229, g230, g231;
	wire g232, g233, g234, g238, g240, g241, g242, g243, g244, g245, g246, g309, g248, g249, g250, g251, g252, g253, g254, g255, g256;
	wire g258, g259, g260, g261, g263, g264, g265, g266, g267, g268, g269, g271, g272, g273, g274, g275, g277, g278, g279, g280, g282;
	wire g283, g284, g285, g286, g287, g289, g290, g292, g293, g294, g295, g296, g297, g299, g308, g301, g302, g304, g305, g306, g312;
	wire g313, g314, g317, g315, g316, g319, g320, g318, g321, g323, g324, g325, g328, g326, g327, g330, g331, g329, g332, g334, g335;
	wire g336, g339, g337, g338, g340, g341, g342, g344, g345, g346, g349, g347, g348, g352, g350, g351, g353, g355, g356, g357, g360;
	wire g358, g359, g362, g363, g361, g364, g366, g367, g368, g369, g370;

	assign o_0_ = (((sk[0]) & (g1)));
	assign o_1_ = (((sk[1]) & (!g3)));
	assign o_2_ = (((sk[2]) & (!g5)));
	assign o_3_ = (((sk[3]) & (!g7)));
	assign o_4_ = (((sk[4]) & (!g10)));
	assign o_6_ = (((sk[5]) & (!g14)));
	assign o_7_ = (((sk[6]) & (!g18)));
	assign o_8_ = (((sk[7]) & (!g20)));
	assign o_9_ = (((sk[8]) & (!g22)));
	assign o_10_ = (((sk[9]) & (g24)));
	assign o_11_ = (((sk[10]) & (!g26)));
	assign o_12_ = (((sk[11]) & (!g28)));
	assign o_13_ = (((sk[12]) & (!g30)));
	assign o_14_ = (((sk[13]) & (!g32)));
	assign o_15_ = (((sk[14]) & (!g33)));
	assign o_16_ = (((sk[15]) & (!g34)));
	assign o_17_ = (((sk[16]) & (g35)));
	assign o_18_ = (((sk[17]) & (!g37)));
	assign o_19_ = (((sk[18]) & (!g40)));
	assign o_20_ = (((sk[19]) & (!g41)));
	assign o_21_ = (((sk[20]) & (!g42)));
	assign o_23_ = (((sk[21]) & (!g45)));
	assign o_24_ = (((sk[22]) & (!g46)));
	assign o_25_ = (((sk[23]) & (!g47)));
	assign o_26_ = (((sk[24]) & (g48)));
	assign o_27_ = (((sk[25]) & (!g49)));
	assign o_28_ = (((sk[26]) & (!g51)));
	assign o_29_ = (((sk[27]) & (!g52)));
	assign o_30_ = (((sk[28]) & (!g53)));
	assign o_31_ = (((sk[29]) & (!g365)));
	assign o_32_ = (((sk[30]) & (!g92)));
	assign o_33_ = (((sk[31]) & (!g94)));
	assign o_34_ = (((sk[32]) & (!g121)));
	assign o_35_ = (((sk[33]) & (!g122)));
	assign o_36_ = (((sk[34]) & (!g124)));
	assign o_37_ = (((sk[35]) & (!g152)));
	assign o_38_ = (((sk[36]) & (!g165)));
	assign o_39_ = (((sk[37]) & (!g175)));
	assign o_40_ = (((sk[38]) & (!g188)));
	assign o_41_ = (((sk[39]) & (!g194)));
	assign o_42_ = (((sk[40]) & (!g207)));
	assign o_43_ = (((sk[41]) & (!g214)));
	assign o_44_ = (((sk[42]) & (!g215)));
	assign o_45_ = (((sk[43]) & (!g223)));
	assign o_46_ = (((sk[44]) & (!g224)));
	assign o_47_ = (((sk[45]) & (!g235)));
	assign o_48_ = (((sk[46]) & (!g236)));
	assign o_49_ = (((sk[47]) & (!g237)));
	assign o_50_ = (((sk[48]) & (!g239)));
	assign o_51_ = (((sk[49]) & (!g247)));
	assign o_52_ = (((sk[50]) & (!g257)));
	assign o_53_ = (((sk[51]) & (!g262)));
	assign o_54_ = (((sk[52]) & (!g270)));
	assign o_55_ = (((sk[53]) & (!g276)));
	assign o_56_ = (((sk[54]) & (!g281)));
	assign o_57_ = (((sk[55]) & (!g288)));
	assign o_58_ = (((sk[56]) & (!g291)));
	assign o_59_ = (((sk[57]) & (!g298)));
	assign o_60_ = (((sk[58]) & (!g300)));
	assign o_61_ = (((sk[59]) & (!g303)));
	assign o_62_ = (((sk[60]) & (!g307)));
	assign g1 = (((!sk[61]) & (!i_4_) & (i_5_) & (!i_6_)) + ((!sk[61]) & (!i_4_) & (!i_5_) & (i_6_)) + ((sk[61]) & (!i_4_) & (!i_5_) & (!i_6_)));
	assign g2 = (((!sk[62]) & (i_6_) & (!i_7_)) + ((sk[62]) & (!i_6_) & (!i_7_)));
	assign g3 = (((i_5_) & (!sk[63]) & (!g2)) + ((!i_5_) & (sk[63]) & (!g2)));
	assign g4 = (((!i_4_) & (i_5_) & (!sk[64]) & (!i_3_)) + ((!i_4_) & (!i_5_) & (!sk[64]) & (i_3_)) + ((!i_4_) & (i_5_) & (!sk[64]) & (!i_3_)));
	assign g5 = (((!g2) & (sk[65]) & (!g4)) + ((g2) & (!sk[65]) & (!g4)) + ((!g2) & (sk[65]) & (!g4)));
	assign g6 = (((!i_4_) & (i_5_) & (!sk[66]) & (!i_3_)) + ((!i_4_) & (!i_5_) & (!sk[66]) & (i_3_)) + ((!i_4_) & (i_5_) & (!sk[66]) & (i_3_)));
	assign g7 = (((!sk[67]) & (g2) & (!g6)) + ((sk[67]) & (!g2) & (!g6)) + ((!sk[67]) & (g2) & (!g6)));
	assign g8 = (((!i_4_) & (i_5_) & (!sk[68]) & (!i_3_)) + ((!i_4_) & (!i_5_) & (!sk[68]) & (i_3_)) + ((!i_4_) & (!i_5_) & (!sk[68]) & (i_3_)));
	assign g9 = (((!sk[69]) & (i_6_) & (!i_7_)) + ((!sk[69]) & (i_6_) & (!i_7_)));
	assign g10 = (((!g8) & (sk[70]) & (!g9)) + ((g8) & (!sk[70]) & (!g9)) + ((!g8) & (sk[70]) & (!g9)));
	assign o_5_ = (((!i_4_) & (!sk[71]) & (i_5_) & (!g9)) + ((!i_4_) & (!sk[71]) & (!i_5_) & (g9)) + ((!i_4_) & (!sk[71]) & (i_5_) & (g9)));
	assign g12 = (((i_6_) & (!sk[72]) & (!g8)) + ((!i_6_) & (sk[72]) & (g8)));
	assign g13 = (((!i_1_) & (i_0_) & (!sk[73]) & (!i_2_)) + ((!i_1_) & (!i_0_) & (!sk[73]) & (i_2_)) + ((!i_1_) & (!i_0_) & (!sk[73]) & (i_2_)));
	assign g14 = (((!sk[74]) & (g12) & (!g13)) + ((sk[74]) & (!g12) & (!g13)) + ((!sk[74]) & (g12) & (!g13)));
	assign g15 = (((!sk[75]) & (i_6_) & (!i_7_)) + ((!sk[75]) & (i_6_) & (i_7_)));
	assign g16 = (((!sk[76]) & (g4) & (!g15)) + ((!sk[76]) & (g4) & (g15)));
	assign g17 = (((!i_1_) & (i_0_) & (!sk[77]) & (!i_2_)) + ((!i_1_) & (!i_0_) & (!sk[77]) & (i_2_)) + ((i_1_) & (!i_0_) & (sk[77]) & (!i_2_)));
	assign g18 = (((!sk[78]) & (g16) & (!g17)) + ((sk[78]) & (!g16) & (!g17)) + ((!sk[78]) & (g16) & (!g17)));
	assign g19 = (((!sk[79]) & (!i_1_) & (i_0_) & (!i_2_)) + ((!sk[79]) & (!i_1_) & (!i_0_) & (i_2_)) + ((!sk[79]) & (i_1_) & (i_0_) & (i_2_)));
	assign g20 = (((!g16) & (sk[80]) & (!g19)) + ((g16) & (!sk[80]) & (!g19)) + ((!g16) & (sk[80]) & (!g19)));
	assign g21 = (((!sk[81]) & (!i_4_) & (i_5_) & (!i_3_)) + ((!sk[81]) & (!i_4_) & (!i_5_) & (i_3_)) + ((sk[81]) & (!i_4_) & (!i_5_) & (!i_3_)));
	assign g22 = (((!g13) & (!g15) & (sk[82]) & (!g21)) + ((!g13) & (!g15) & (!sk[82]) & (g21)) + ((!g13) & (!g15) & (!sk[82]) & (g21)) + ((!g13) & (g15) & (!sk[82]) & (!g21)));
	assign g23 = (((!i_1_) & (i_0_) & (!sk[83]) & (!i_2_)) + ((!i_1_) & (!i_0_) & (!sk[83]) & (i_2_)) + ((!i_1_) & (!i_0_) & (sk[83]) & (!i_2_)) + ((!i_1_) & (!i_0_) & (!sk[83]) & (i_2_)));
	assign g24 = (((i_4_) & (!i_5_) & (!g15) & (!sk[84]) & (!g23)) + ((!i_4_) & (!i_5_) & (g15) & (!sk[84]) & (!g23)) + ((!i_4_) & (i_5_) & (g15) & (!sk[84]) & (!g23)));
	assign g25 = (((!i_1_) & (sk[85]) & (!i_0_) & (!i_2_)) + ((!i_1_) & (!sk[85]) & (i_0_) & (!i_2_)) + ((i_1_) & (!sk[85]) & (!i_0_) & (!i_2_)) + ((!i_1_) & (!sk[85]) & (i_0_) & (i_2_)));
	assign g26 = (((!g16) & (!sk[86]) & (g25)) + ((!g16) & (sk[86]) & (!g25)));
	assign g27 = (((i_1_) & (!sk[87]) & (!i_0_) & (!i_2_)) + ((!i_1_) & (!sk[87]) & (i_0_) & (!i_2_)) + ((!i_1_) & (sk[87]) & (!i_0_) & (!i_2_)) + ((!i_1_) & (!sk[87]) & (i_0_) & (!i_2_)));
	assign g28 = (((!g16) & (!sk[88]) & (g27)) + ((!g16) & (sk[88]) & (!g27)));
	assign g29 = (((!sk[89]) & (!g6) & (g15)) + ((!sk[89]) & (g6) & (g15)));
	assign g30 = (((!sk[90]) & (!g17) & (g29)) + ((sk[90]) & (!g17) & (!g29)) + ((!sk[90]) & (!g17) & (g29)));
	assign g31 = (((i_1_) & (!i_0_) & (!sk[91]) & (!i_2_)) + ((!i_1_) & (!i_0_) & (sk[91]) & (!i_2_)) + ((!i_1_) & (i_0_) & (!sk[91]) & (!i_2_)) + ((!i_1_) & (!i_0_) & (sk[91]) & (i_2_)));
	assign g32 = (((!g29) & (!sk[92]) & (g31)) + ((!g29) & (sk[92]) & (!g31)));
	assign g33 = (((!sk[93]) & (!g23) & (g29)) + ((sk[93]) & (!g23) & (!g29)) + ((!sk[93]) & (g23) & (g29)));
	assign g34 = (((!sk[94]) & (!g25) & (g29)) + ((sk[94]) & (!g25) & (!g29)) + ((!sk[94]) & (g25) & (g29)));
	assign g35 = (((i_4_) & (!i_5_) & (!sk[95]) & (!g31)) + ((!i_4_) & (i_5_) & (!sk[95]) & (!g31)) + ((i_4_) & (!i_5_) & (!sk[95]) & (!g31)));
	assign g36 = (((i_4_) & (!sk[96]) & (i_3_)) + ((!i_4_) & (!sk[96]) & (i_3_)));
	assign g37 = (((i_5_) & (!g13) & (!sk[97]) & (!g36)) + ((!i_5_) & (!g13) & (sk[97]) & (!g36)) + ((!i_5_) & (g13) & (!sk[97]) & (!g36)) + ((!i_5_) & (!g13) & (sk[97]) & (!g36)));
	assign g38 = (((!i_4_) & (!sk[98]) & (i_3_)) + ((i_4_) & (sk[98]) & (!i_3_)));
	assign g39 = (((!sk[99]) & (i_1_) & (!i_0_) & (!i_2_)) + ((!sk[99]) & (!i_1_) & (i_0_) & (!i_2_)) + ((sk[99]) & (!i_1_) & (!i_0_) & (!i_2_)));
	assign g40 = (((!g38) & (!sk[100]) & (g39)) + ((!g38) & (sk[100]) & (!g39)) + ((!g38) & (!sk[100]) & (g39)));
	assign g41 = (((i_6_) & (!sk[101]) & (!g21) & (!g31)) + ((!i_6_) & (!sk[101]) & (g21) & (!g31)) + ((!i_6_) & (sk[101]) & (!g21) & (!g31)) + ((!i_6_) & (!sk[101]) & (g21) & (g31)));
	assign g42 = (((!sk[102]) & (!g12) & (g31)) + ((sk[102]) & (!g12) & (!g31)));
	assign o_22_ = (((!sk[103]) & (i_4_) & (!i_5_) & (!g15) & (!g31)) + ((!sk[103]) & (!i_4_) & (i_5_) & (!g15) & (!g31)) + ((sk[103]) & (!i_4_) & (!i_5_) & (g15) & (!g31)));
	assign g44 = (((i_4_) & (!i_5_) & (!sk[104]) & (!i_3_)) + ((!i_4_) & (i_5_) & (!sk[104]) & (!i_3_)) + ((i_4_) & (i_5_) & (!sk[104]) & (i_3_)));
	assign g45 = (((!g6) & (!g39) & (sk[105]) & (!g44)) + ((!g6) & (g39) & (!sk[105]) & (!g44)) + ((g6) & (!g39) & (!sk[105]) & (!g44)) + ((!g6) & (!g39) & (sk[105]) & (!g44)));
	assign g46 = (((!sk[106]) & (g9) & (!g21) & (!g39)) + ((!sk[106]) & (!g9) & (g21) & (!g39)) + ((sk[106]) & (!g9) & (!g21) & (!g39)) + ((!sk[106]) & (!g9) & (g21) & (!g39)));
	assign g47 = (((!g9) & (g17) & (!sk[107]) & (!g21)) + ((!g9) & (!g17) & (sk[107]) & (!g21)) + ((g9) & (!g17) & (!sk[107]) & (!g21)) + ((!g9) & (!g17) & (sk[107]) & (!g21)));
	assign g48 = (((i_0_) & (!i_2_) & (!sk[108]) & (!g15) & (!g21)) + ((!i_0_) & (i_2_) & (!sk[108]) & (!g15) & (!g21)) + ((i_0_) & (i_2_) & (!sk[108]) & (g15) & (g21)));
	assign g49 = (((!g9) & (sk[109]) & (!g21) & (!g23)) + ((!g9) & (!sk[109]) & (g21) & (!g23)) + ((g9) & (!sk[109]) & (!g21) & (!g23)) + ((!g9) & (!sk[109]) & (g21) & (g23)));
	assign g50 = (((g8) & (!sk[110]) & (g15)) + ((!g8) & (!sk[110]) & (g15)));
	assign g51 = (((!sk[111]) & (!g27) & (g50)) + ((sk[111]) & (!g27) & (!g50)) + ((!sk[111]) & (g27) & (g50)));
	assign g52 = (((i_6_) & (!sk[112]) & (!i_7_) & (!g21) & (!g39)) + ((!i_6_) & (!sk[112]) & (i_7_) & (!g21) & (!g39)) + ((!i_6_) & (sk[112]) & (!i_7_) & (!g21) & (!g39)) + ((!i_6_) & (!sk[112]) & (i_7_) & (!g21) & (!g39)) + ((!i_6_) & (!sk[112]) & (i_7_) & (!g21) & (!g39)));
	assign g53 = (((!sk[113]) & (g15) & (!g19) & (!g21)) + ((!sk[113]) & (!g15) & (g19) & (!g21)) + ((sk[113]) & (!g15) & (!g19) & (!g21)) + ((!sk[113]) & (!g15) & (g19) & (!g21)));
	assign g54 = (((!i_6_) & (!i_7_) & (!sk[114]) & (g6) & (!g21) & (!g27)) + ((!i_6_) & (!i_7_) & (!sk[114]) & (g6) & (!g21) & (!g27)) + ((!i_6_) & (!i_7_) & (!sk[114]) & (g6) & (!g21) & (!g27)) + ((!i_6_) & (!i_7_) & (!sk[114]) & (!g6) & (g21) & (!g27)) + ((!i_6_) & (!i_7_) & (!sk[114]) & (!g6) & (g21) & (!g27)) + ((!i_6_) & (!i_7_) & (!sk[114]) & (!g6) & (g21) & (!g27)));
	assign g55 = (((i_6_) & (!g6) & (!g36) & (!sk[115]) & (!g39)) + ((!i_6_) & (g6) & (!g36) & (!sk[115]) & (!g39)) + ((i_6_) & (g6) & (!g36) & (!sk[115]) & (g39)) + ((!i_6_) & (!g6) & (g36) & (sk[115]) & (g39)));
	assign g56 = (((i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (g13)) + ((!i_4_) & (i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (g13)) + ((!i_4_) & (!i_5_) & (i_6_) & (!i_7_) & (!i_3_) & (g13)) + ((!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (i_3_) & (g13)) + ((!i_4_) & (!i_5_) & (!i_6_) & (i_7_) & (i_3_) & (g13)));
	assign g57 = (((i_6_) & (!sk[117]) & (!g13) & (!g21) & (!g56)) + ((!i_6_) & (!sk[117]) & (g13) & (!g21) & (!g56)) + ((i_6_) & (!sk[117]) & (!g13) & (!g21) & (!g56)) + ((!i_6_) & (sk[117]) & (!g13) & (!g21) & (!g56)) + ((!i_6_) & (!sk[117]) & (g13) & (!g21) & (!g56)));
	assign g58 = (((!sk[118]) & (!g55) & (g57)) + ((!sk[118]) & (!g55) & (g57)));
	assign g59 = (((!g27) & (g29) & (!sk[119]) & (!g36)) + ((g27) & (!g29) & (!sk[119]) & (!g36)) + ((!g27) & (!g29) & (sk[119]) & (g36)));
	assign g60 = (((i_5_) & (!sk[120]) & (!g12) & (!g38)) + ((!i_5_) & (!sk[120]) & (g12) & (!g38)) + ((!i_5_) & (sk[120]) & (!g12) & (!g38)) + ((!i_5_) & (sk[120]) & (!g12) & (!g38)));
	assign g61 = (((!i_6_) & (!i_7_) & (g4) & (!g21) & (!sk[121]) & (!g25)) + ((!i_6_) & (!i_7_) & (!g4) & (g21) & (!sk[121]) & (!g25)) + ((!i_6_) & (i_7_) & (g4) & (!g21) & (!sk[121]) & (!g25)) + ((i_6_) & (!i_7_) & (g4) & (!g21) & (!sk[121]) & (!g25)) + ((i_6_) & (!i_7_) & (!g4) & (g21) & (!sk[121]) & (!g25)));
	assign g62 = (((!sk[122]) & (!g5) & (g61)) + ((sk[122]) & (g5) & (!g61)));
	assign g63 = (((i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (g19)) + ((!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (i_3_) & (g19)) + ((!i_4_) & (!i_5_) & (i_6_) & (!i_7_) & (i_3_) & (!g19)) + ((!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (g19)) + ((!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (g19)));
	assign g64 = (((g27) & (!g50) & (g53) & (!g60) & (g62) & (!g63)) + ((!g27) & (!g50) & (g53) & (g60) & (g62) & (!g63)));
	assign g65 = (((i_6_) & (!sk[125]) & (!i_7_) & (!g6) & (!g27)) + ((!i_6_) & (!sk[125]) & (i_7_) & (!g6) & (!g27)) + ((!i_6_) & (!sk[125]) & (i_7_) & (g6) & (!g27)) + ((i_6_) & (!sk[125]) & (!i_7_) & (g6) & (!g27)));
	assign g66 = (((i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (!g25)) + ((!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (!g25)) + ((i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (!g25)) + ((!i_4_) & (i_5_) & (!i_6_) & (!i_7_) & (i_3_) & (!g25)) + ((!i_4_) & (!i_5_) & (!i_6_) & (i_7_) & (i_3_) & (!g25)) + ((!i_4_) & (i_5_) & (i_6_) & (i_7_) & (!i_3_) & (!g25)));
	assign g67 = (((!g15) & (!g21) & (g25) & (!g27) & (!sk[127]) & (!g44)) + ((!g15) & (!g21) & (!g25) & (g27) & (!sk[127]) & (!g44)) + ((!g15) & (!g21) & (!g25) & (!g27) & (sk[127]) & (g44)) + ((g15) & (g21) & (!g25) & (!g27) & (sk[127]) & (!g44)));
	assign g68 = (((i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (i_3_) & (g19)) + ((!i_4_) & (i_5_) & (!i_6_) & (!i_7_) & (i_3_) & (g19)) + ((!i_4_) & (i_5_) & (i_6_) & (i_7_) & (!i_3_) & (g19)));
	assign g69 = (((!i_5_) & (g16) & (!sk[1]) & (!g27) & (!g38) & (!g68)) + ((!i_5_) & (!g16) & (!sk[1]) & (!g27) & (g38) & (!g68)) + ((!i_5_) & (!g16) & (!sk[1]) & (!g27) & (!g38) & (g68)) + ((!i_5_) & (!g16) & (sk[1]) & (!g27) & (!g38) & (!g68)) + ((!i_5_) & (!g16) & (sk[1]) & (g27) & (!g38) & (!g68)) + ((i_5_) & (!g16) & (!sk[1]) & (!g27) & (g38) & (!g68)));
	assign g70 = (((!g59) & (g64) & (!g65) & (!g66) & (!g67) & (g69)));
	assign g71 = (((!sk[3]) & (!i_6_) & (i_7_) & (!g4) & (!g21) & (!g31)) + ((!sk[3]) & (!i_6_) & (!i_7_) & (!g4) & (g21) & (!g31)) + ((!sk[3]) & (!i_6_) & (!i_7_) & (!g4) & (!g21) & (g31)) + ((!sk[3]) & (i_6_) & (!i_7_) & (!g4) & (g21) & (!g31)) + ((!sk[3]) & (!i_6_) & (i_7_) & (g4) & (!g21) & (!g31)) + ((sk[3]) & (i_6_) & (!i_7_) & (g4) & (!g21) & (!g31)));
	assign g72 = (((!g5) & (!g31) & (!sk[4]) & (g71)) + ((g5) & (!g31) & (sk[4]) & (!g71)) + ((!g5) & (g31) & (sk[4]) & (!g71)));
	assign g73 = (((!sk[5]) & (!g15) & (!g21) & (g23)) + ((sk[5]) & (g15) & (g21) & (!g23)));
	assign g74 = (((i_6_) & (!g21) & (!sk[6]) & (!g23) & (!g30)) + ((!i_6_) & (!g21) & (!sk[6]) & (g23) & (!g30)) + ((i_6_) & (!g21) & (!sk[6]) & (!g23) & (g30)) + ((!i_6_) & (!g21) & (!sk[6]) & (g23) & (g30)) + ((!i_6_) & (!g21) & (sk[6]) & (!g23) & (g30)));
	assign g75 = (((!sk[7]) & (!g17) & (!g36) & (g49)) + ((!sk[7]) & (!g17) & (!g36) & (g49)) + ((!sk[7]) & (!g17) & (!g36) & (g49)));
	assign g76 = (((!i_6_) & (!i_7_) & (!g6) & (g21) & (!g23) & (!g31)) + ((!i_6_) & (i_7_) & (g6) & (!g21) & (!g23) & (!g31)));
	assign g77 = (((i_4_) & (!sk[9]) & (!i_5_) & (!i_3_) & (!g15)) + ((!i_4_) & (!sk[9]) & (i_5_) & (!i_3_) & (!g15)) + ((i_4_) & (!sk[9]) & (!i_5_) & (!i_3_) & (!g15)) + ((!i_4_) & (!sk[9]) & (i_5_) & (!i_3_) & (g15)));
	assign g78 = (((!sk[10]) & (g31) & (!g77)) + ((sk[10]) & (!g31) & (g77)));
	assign g79 = (((!sk[11]) & (g2) & (!g8)) + ((sk[11]) & (!g2) & (!g8)) + ((!sk[11]) & (g2) & (!g8)));
	assign g80 = (((i_7_) & (!sk[12]) & (!g8)) + ((i_7_) & (!sk[12]) & (g8)));
	assign g81 = (((g17) & (!sk[13]) & (!g38) & (!g79) & (!g80)) + ((g17) & (!sk[13]) & (g38) & (!g79) & (!g80)) + ((!g17) & (!sk[13]) & (g38) & (!g79) & (!g80)) + ((g17) & (!sk[13]) & (!g38) & (!g79) & (!g80)) + ((g17) & (!sk[13]) & (!g38) & (!g79) & (g80)));
	assign g82 = (((g12) & (!g16) & (!g23) & (!sk[14]) & (!g38)) + ((!g12) & (g16) & (!g23) & (!sk[14]) & (!g38)) + ((g12) & (!g16) & (!g23) & (!sk[14]) & (!g38)) + ((!g12) & (g16) & (!g23) & (!sk[14]) & (!g38)) + ((!g12) & (!g16) & (!g23) & (sk[14]) & (g38)));
	assign g83 = (((g78) & (!g81) & (!sk[15]) & (!g82)) + ((!g78) & (!g81) & (!sk[15]) & (g82)) + ((!g78) & (!g81) & (sk[15]) & (!g82)));
	assign g84 = (((g72) & (!g73) & (g74) & (g75) & (g354) & (g83)));
	assign g85 = (((i_6_) & (!i_7_) & (!sk[17]) & (!g4) & (!g39)) + ((!i_6_) & (i_7_) & (!sk[17]) & (!g4) & (!g39)) + ((i_6_) & (!i_7_) & (!sk[17]) & (g4) & (g39)) + ((!i_6_) & (i_7_) & (!sk[17]) & (g4) & (g39)));
	assign g86 = (((!sk[18]) & (g5) & (!g39) & (!g85)) + ((!sk[18]) & (g5) & (!g39) & (!g85)) + ((sk[18]) & (!g5) & (!g39) & (!g85)));
	assign g87 = (((g12) & (!g38) & (!g39) & (!sk[19]) & (!g86)) + ((!g12) & (!g38) & (!g39) & (!sk[19]) & (g86)) + ((!g12) & (!g38) & (!g39) & (!sk[19]) & (g86)) + ((!g12) & (!g38) & (!g39) & (!sk[19]) & (g86)));
	assign g88 = (((!sk[20]) & (i_6_) & (!i_7_) & (!g6) & (!g8) & (!g39)) + ((!sk[20]) & (!i_6_) & (!i_7_) & (!g6) & (g8) & (!g39)) + ((sk[20]) & (!i_6_) & (!i_7_) & (g6) & (!g8) & (g39)) + ((!sk[20]) & (i_6_) & (i_7_) & (!g6) & (g8) & (g39)));
	assign g89 = (((!i_6_) & (!i_7_) & (g17) & (g21) & (!sk[21]) & (!g39)) + ((i_6_) & (!i_7_) & (!g17) & (!g21) & (!sk[21]) & (!g39)) + ((!i_6_) & (!i_7_) & (!g17) & (g21) & (!sk[21]) & (!g39)) + ((!i_6_) & (!i_7_) & (!g17) & (g21) & (!sk[21]) & (g39)) + ((!i_6_) & (i_7_) & (!g17) & (g21) & (!sk[21]) & (g39)));
	assign g90 = (((!sk[22]) & (g13) & (!g29) & (!g31) & (!g50) & (!g89)) + ((!sk[22]) & (!g13) & (!g29) & (!g31) & (g50) & (!g89)) + ((sk[22]) & (!g13) & (!g29) & (!g31) & (!g50) & (!g89)) + ((!sk[22]) & (g13) & (!g29) & (g31) & (!g50) & (!g89)) + ((!sk[22]) & (!g13) & (!g29) & (g31) & (g50) & (!g89)) + ((!sk[22]) & (g13) & (!g29) & (!g31) & (!g50) & (!g89)));
	assign g91 = (((g18) & (!sk[23]) & (!g35) & (!g87) & (!g88) & (!g90)) + ((!g18) & (!sk[23]) & (!g35) & (!g87) & (g88) & (!g90)) + ((g18) & (!sk[23]) & (!g35) & (g87) & (!g88) & (g90)));
	assign g92 = (((g32) & (!g54) & (g58) & (g70) & (g84) & (g91)));
	assign g93 = (((!sk[25]) & (i_5_) & (!i_3_) & (!i_1_)) + ((!sk[25]) & (i_5_) & (!i_3_) & (!i_1_)) + ((sk[25]) & (!i_5_) & (i_3_) & (i_1_)));
	assign g94 = (((i_4_) & (!i_0_) & (!sk[26]) & (!i_2_) & (!g15) & (!g93)) + ((!i_4_) & (!i_0_) & (!sk[26]) & (!i_2_) & (g15) & (!g93)) + ((!i_4_) & (i_0_) & (!sk[26]) & (i_2_) & (g15) & (!g93)));
	assign g95 = (((!sk[27]) & (g17) & (!g21)) + ((!sk[27]) & (g17) & (g21)));
	assign g96 = (((g13) & (!g29) & (!sk[28]) & (!g36) & (!g95)) + ((!g13) & (!g29) & (!sk[28]) & (!g36) & (g95)) + ((!g13) & (!g29) & (sk[28]) & (!g36) & (!g95)) + ((!g13) & (!g29) & (sk[28]) & (!g36) & (!g95)));
	assign g97 = (((g18) & (!sk[29]) & (!g96)) + ((g18) & (!sk[29]) & (g96)));
	assign g98 = (((g12) & (!g16) & (!sk[30]) & (!g25) & (!g31) & (!g44)) + ((!g12) & (!g16) & (!sk[30]) & (!g25) & (g31) & (!g44)) + ((!g12) & (!g16) & (!sk[30]) & (g25) & (g31) & (!g44)) + ((!g12) & (!g16) & (!sk[30]) & (!g25) & (g31) & (!g44)) + ((!g12) & (!g16) & (sk[30]) & (g25) & (!g31) & (!g44)) + ((!g12) & (!g16) & (sk[30]) & (!g25) & (!g31) & (!g44)));
	assign g99 = (((i_6_) & (!sk[31]) & (!i_7_) & (!g13) & (!g21) & (!g39)) + ((!i_6_) & (!sk[31]) & (i_7_) & (!g13) & (!g21) & (!g39)) + ((!i_6_) & (sk[31]) & (!i_7_) & (g13) & (g21) & (!g39)) + ((!i_6_) & (sk[31]) & (!i_7_) & (!g13) & (g21) & (g39)) + ((!i_6_) & (sk[31]) & (!i_7_) & (!g13) & (g21) & (g39)));
	assign g100 = (((!g55) & (!g98) & (!sk[32]) & (g99)) + ((!g55) & (g98) & (sk[32]) & (!g99)));
	assign g101 = (((!sk[33]) & (!i_6_) & (!g21) & (g25)) + ((sk[33]) & (!i_6_) & (g21) & (!g25)));
	assign g102 = (((!sk[34]) & (i_1_) & (!i_0_) & (!i_2_) & (!g50) & (!g101)) + ((!sk[34]) & (!i_1_) & (i_0_) & (!i_2_) & (!g50) & (!g101)) + ((!sk[34]) & (!i_1_) & (i_0_) & (!i_2_) & (!g50) & (!g101)) + ((!sk[34]) & (!i_1_) & (i_0_) & (i_2_) & (!g50) & (!g101)) + ((sk[34]) & (!i_1_) & (!i_0_) & (!i_2_) & (!g50) & (!g101)) + ((sk[34]) & (!i_1_) & (!i_0_) & (i_2_) & (!g50) & (!g101)) + ((!sk[34]) & (i_1_) & (!i_0_) & (!i_2_) & (!g50) & (!g101)));
	assign g103 = (((!sk[35]) & (g16) & (!g19) & (!g29) & (!g36) & (!g102)) + ((!sk[35]) & (!g16) & (g19) & (!g29) & (!g36) & (!g102)) + ((sk[35]) & (!g16) & (!g19) & (!g29) & (!g36) & (g102)) + ((!sk[35]) & (!g16) & (g19) & (!g29) & (!g36) & (g102)));
	assign g104 = (((i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (g39)) + ((!i_4_) & (i_5_) & (i_6_) & (!i_7_) & (!i_3_) & (g39)) + ((!i_4_) & (i_5_) & (!i_6_) & (i_7_) & (!i_3_) & (g39)) + ((!i_4_) & (!i_5_) & (i_6_) & (i_7_) & (!i_3_) & (g39)) + ((!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (i_3_) & (g39)));
	assign g105 = (((i_4_) & (!sk[37]) & (!i_5_) & (!i_3_) & (!g15) & (!g27)) + ((!i_4_) & (!sk[37]) & (i_5_) & (!i_3_) & (!g15) & (!g27)) + ((i_4_) & (!sk[37]) & (!i_5_) & (!i_3_) & (!g15) & (!g27)) + ((!i_4_) & (sk[37]) & (!i_5_) & (!i_3_) & (g15) & (!g27)));
	assign g106 = (((i_4_) & (!sk[38]) & (!i_5_) & (!g2) & (!i_3_) & (!g25)) + ((!i_4_) & (!sk[38]) & (i_5_) & (!g2) & (!i_3_) & (!g25)) + ((i_4_) & (!sk[38]) & (!i_5_) & (!g2) & (!i_3_) & (!g25)) + ((i_4_) & (!sk[38]) & (i_5_) & (!g2) & (!i_3_) & (!g25)) + ((!i_4_) & (!sk[38]) & (i_5_) & (!g2) & (i_3_) & (!g25)));
	assign g107 = (((g27) & (!sk[39]) & (!g29) & (!g36) & (!g105) & (!g106)) + ((!g27) & (!sk[39]) & (g29) & (!g36) & (!g105) & (!g106)) + ((g27) & (!sk[39]) & (!g29) & (!g36) & (!g105) & (!g106)) + ((!g27) & (sk[39]) & (!g29) & (!g36) & (!g105) & (!g106)));
	assign g108 = (((g64) & (!g100) & (!g103) & (!sk[40]) & (!g104) & (!g107)) + ((!g64) & (!g100) & (g103) & (!sk[40]) & (!g104) & (!g107)) + ((!g64) & (g100) & (!g103) & (!sk[40]) & (!g104) & (g107)) + ((g64) & (g100) & (g103) & (!sk[40]) & (!g104) & (g107)));
	assign g109 = (((i_6_) & (!g17) & (!g21) & (!sk[41]) & (!g23) & (!g44)) + ((!i_6_) & (!g17) & (g21) & (!sk[41]) & (!g23) & (!g44)) + ((!i_6_) & (g17) & (!g21) & (!sk[41]) & (!g23) & (g44)) + ((!i_6_) & (!g17) & (g21) & (!sk[41]) & (!g23) & (!g44)));
	assign g110 = (((!sk[42]) & (!i_5_) & (g17) & (!g36) & (!g109)) + ((!sk[42]) & (!i_5_) & (!g17) & (!g36) & (g109)) + ((!sk[42]) & (i_5_) & (!g17) & (!g36) & (!g109)) + ((sk[42]) & (!i_5_) & (!g17) & (!g36) & (!g109)) + ((!sk[42]) & (!i_5_) & (g17) & (!g36) & (!g109)));
	assign g111 = (((!sk[43]) & (i_6_) & (!i_7_) & (!g6) & (!g17)) + ((!sk[43]) & (!i_6_) & (i_7_) & (!g6) & (!g17)) + ((!sk[43]) & (!i_6_) & (!i_7_) & (!g6) & (g17)) + ((!sk[43]) & (i_6_) & (!i_7_) & (g6) & (g17)) + ((!sk[43]) & (!i_6_) & (i_7_) & (g6) & (g17)));
	assign g112 = (((i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (!g23)) + ((!i_4_) & (!i_5_) & (i_6_) & (!i_7_) & (!i_3_) & (!g23)) + ((!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (i_3_) & (!g23)) + ((!i_4_) & (!i_5_) & (i_6_) & (i_7_) & (!i_3_) & (!g23)));
	assign g113 = (((!i_4_) & (i_5_) & (!i_6_) & (i_7_) & (i_3_) & (!g31)) + ((!i_4_) & (i_5_) & (i_6_) & (!i_7_) & (i_3_) & (!g31)) + ((!i_4_) & (!i_5_) & (!i_6_) & (i_7_) & (i_3_) & (!g31)) + ((!i_4_) & (i_5_) & (i_6_) & (i_7_) & (!i_3_) & (!g31)));
	assign g114 = (((!sk[46]) & (g110) & (!g111) & (!g112) & (!g113)) + ((!sk[46]) & (!g110) & (g111) & (!g112) & (!g113)) + ((!sk[46]) & (!g110) & (!g111) & (!g112) & (g113)) + ((!sk[46]) & (g110) & (!g111) & (!g112) & (!g113)));
	assign g115 = (((!sk[47]) & (!g15) & (g21)) + ((!sk[47]) & (!g15) & (g21)));
	assign g116 = (((!sk[48]) & (i_4_) & (!g23) & (!g29) & (!g31) & (!g115)) + ((!sk[48]) & (!i_4_) & (!g23) & (g29) & (!g31) & (!g115)) + ((!sk[48]) & (!i_4_) & (g23) & (!g29) & (!g31) & (g115)) + ((sk[48]) & (!i_4_) & (!g23) & (!g29) & (g31) & (!g115)) + ((sk[48]) & (!i_4_) & (!g23) & (!g29) & (!g31) & (!g115)) + ((sk[48]) & (!i_4_) & (g23) & (!g29) & (g31) & (!g115)) + ((sk[48]) & (!i_4_) & (g23) & (!g29) & (!g31) & (!g115)));
	assign g117 = (((!g27) & (!sk[49]) & (g115)) + ((!g27) & (!sk[49]) & (g115)));
	assign g118 = (((!sk[50]) & (g12) & (!g13) & (!g38) & (!g50)) + ((!sk[50]) & (!g12) & (g13) & (!g38) & (!g50)) + ((!sk[50]) & (g12) & (g13) & (!g38) & (!g50)) + ((!sk[50]) & (!g12) & (g13) & (g38) & (!g50)) + ((!sk[50]) & (!g12) & (!g13) & (!g38) & (g50)) + ((!sk[50]) & (!g12) & (g13) & (!g38) & (g50)));
	assign g119 = (((g13) & (!sk[51]) & (!g16) & (!g29) & (!g31) & (!g79)) + ((!g13) & (!sk[51]) & (!g16) & (g29) & (!g31) & (!g79)) + ((!g13) & (sk[51]) & (!g16) & (!g29) & (g31) & (!g79)) + ((!g13) & (sk[51]) & (!g16) & (!g29) & (g31) & (!g79)) + ((!g13) & (!sk[51]) & (g16) & (!g29) & (!g31) & (g79)) + ((!g13) & (sk[51]) & (!g16) & (!g29) & (!g31) & (g79)));
	assign g120 = (((g22) & (!g117) & (!g118) & (!sk[52]) & (!g81) & (!g119)) + ((!g22) & (!g117) & (g118) & (!sk[52]) & (!g81) & (!g119)) + ((!g22) & (g117) & (!g118) & (!sk[52]) & (!g81) & (g119)) + ((g22) & (!g117) & (!g118) & (!sk[52]) & (!g81) & (g119)));
	assign g121 = (((g97) & (!g108) & (!sk[53]) & (!g114) & (!g116) & (!g120)) + ((!g97) & (!g108) & (!sk[53]) & (g114) & (!g116) & (!g120)) + ((!g97) & (g108) & (!sk[53]) & (!g114) & (!g116) & (g120)) + ((g97) & (g108) & (!sk[53]) & (g114) & (g116) & (g120)));
	assign g122 = (((i_4_) & (i_5_) & (!i_3_) & (!i_1_) & (i_0_) & (!i_2_)) + ((i_4_) & (!i_5_) & (!i_3_) & (!i_1_) & (!i_0_) & (!i_2_)) + ((i_4_) & (i_5_) & (i_3_) & (!i_1_) & (!i_0_) & (i_2_)));
	assign g123 = (((i_4_) & (!i_3_) & (!g9) & (!sk[55]) & (!i_0_) & (!i_2_)) + ((!i_4_) & (!i_3_) & (g9) & (!sk[55]) & (!i_0_) & (!i_2_)) + ((!i_4_) & (i_3_) & (!g9) & (!sk[55]) & (!i_0_) & (i_2_)) + ((i_4_) & (!i_3_) & (!g9) & (!sk[55]) & (i_0_) & (!i_2_)) + ((!i_4_) & (!i_3_) & (g9) & (!sk[55]) & (!i_0_) & (i_2_)));
	assign g124 = (((i_5_) & (!i_1_) & (!sk[56]) & (!g123)) + ((!i_5_) & (i_1_) & (!sk[56]) & (!g123)) + ((!i_5_) & (!i_1_) & (sk[56]) & (g123)));
	assign g125 = (((!sk[57]) & (i_6_) & (!g5) & (!g21) & (!g23) & (!g38)) + ((!sk[57]) & (!i_6_) & (!g5) & (!g21) & (g23) & (!g38)) + ((!sk[57]) & (!i_6_) & (!g5) & (!g21) & (!g23) & (g38)) + ((sk[57]) & (!i_6_) & (!g5) & (!g21) & (!g23) & (!g38)) + ((!sk[57]) & (i_6_) & (!g5) & (g21) & (!g23) & (!g38)));
	assign g126 = (((!sk[58]) & (i_6_) & (!i_7_) & (!g4) & (!g23) & (!g109)) + ((!sk[58]) & (!i_6_) & (!i_7_) & (!g4) & (!g23) & (g109)) + ((!sk[58]) & (!i_6_) & (!i_7_) & (!g4) & (g23) & (!g109)) + ((!sk[58]) & (i_6_) & (i_7_) & (!g4) & (!g23) & (!g109)) + ((sk[58]) & (!i_6_) & (!i_7_) & (!g4) & (!g23) & (!g109)) + ((sk[58]) & (!i_6_) & (!i_7_) & (!g4) & (!g23) & (!g109)));
	assign g127 = (((!g16) & (!sk[59]) & (g23) & (!g125) & (!g126)) + ((!g16) & (!sk[59]) & (!g23) & (g125) & (!g126)) + ((!g16) & (!sk[59]) & (g23) & (!g125) & (g126)) + ((!g16) & (sk[59]) & (!g23) & (!g125) & (g126)));
	assign g128 = (((!sk[60]) & (g23) & (!g79) & (!g127)) + ((!sk[60]) & (!g23) & (g79) & (!g127)) + ((!sk[60]) & (g23) & (!g79) & (g127)) + ((!sk[60]) & (!g23) & (g79) & (g127)));
	assign g129 = (((!i_6_) & (!sk[61]) & (i_7_) & (!g19) & (!g21)) + ((!i_6_) & (!sk[61]) & (!i_7_) & (g19) & (!g21)) + ((!i_6_) & (!sk[61]) & (!i_7_) & (g19) & (g21)) + ((!i_6_) & (!sk[61]) & (!i_7_) & (g19) & (g21)));
	assign g130 = (((!sk[62]) & (!g53) & (g129)) + ((sk[62]) & (g53) & (!g129)));
	assign g131 = (((!g27) & (g31) & (!sk[63]) & (!g50) & (!g59)) + ((!g27) & (!g31) & (!sk[63]) & (g50) & (!g59)) + ((g27) & (g31) & (!sk[63]) & (!g50) & (!g59)) + ((!g27) & (!g31) & (sk[63]) & (!g50) & (!g59)));
	assign g132 = (((!g19) & (!g38) & (g72) & (g130) & (g354) & (g131)) + ((!g19) & (!g38) & (g72) & (g130) & (g354) & (g131)));
	assign g133 = (((!i_6_) & (i_7_) & (!g6) & (!sk[65]) & (!g13)) + ((!i_6_) & (!i_7_) & (g6) & (!sk[65]) & (!g13)) + ((!i_6_) & (!i_7_) & (g6) & (!sk[65]) & (g13)) + ((!i_6_) & (!i_7_) & (g6) & (!sk[65]) & (g13)));
	assign g134 = (((!i_6_) & (g4) & (!sk[66]) & (!g17) & (!g38)) + ((!i_6_) & (!g4) & (!sk[66]) & (g17) & (!g38)) + ((!i_6_) & (!g4) & (!sk[66]) & (!g17) & (g38)) + ((!i_6_) & (!g4) & (!sk[66]) & (g17) & (g38)) + ((i_6_) & (g4) & (!sk[66]) & (g17) & (!g38)));
	assign g135 = (((!sk[67]) & (!i_6_) & (g8) & (!g17)) + ((!sk[67]) & (!i_6_) & (g8) & (g17)));
	assign g136 = (((!sk[68]) & (!g133) & (g310)) + ((sk[68]) & (!g133) & (!g310)));
	assign g137 = (((!sk[69]) & (!g13) & (g29) & (!g36)) + ((!sk[69]) & (g13) & (g29) & (!g36)) + ((sk[69]) & (g13) & (!g29) & (g36)));
	assign g138 = (((!i_6_) & (i_7_) & (!g4) & (!g21) & (!sk[70]) & (!g27)) + ((!i_6_) & (!i_7_) & (g4) & (!g21) & (!sk[70]) & (!g27)) + ((!i_6_) & (!i_7_) & (!g4) & (g21) & (!sk[70]) & (!g27)) + ((!i_6_) & (!i_7_) & (!g4) & (!g21) & (!sk[70]) & (g27)) + ((i_6_) & (!i_7_) & (!g4) & (g21) & (!sk[70]) & (!g27)) + ((!i_6_) & (!i_7_) & (g4) & (!g21) & (!sk[70]) & (!g27)));
	assign g139 = (((!i_5_) & (!g31) & (g36) & (!sk[71]) & (!g137) & (!g138)) + ((!i_5_) & (!g31) & (!g36) & (!sk[71]) & (g137) & (!g138)) + ((!i_5_) & (!g31) & (!g36) & (!sk[71]) & (!g137) & (g138)) + ((!i_5_) & (g31) & (!g36) & (!sk[71]) & (!g137) & (!g138)) + ((!i_5_) & (!g31) & (!g36) & (sk[71]) & (!g137) & (!g138)) + ((i_5_) & (!g31) & (!g36) & (sk[71]) & (!g137) & (!g138)));
	assign g140 = (((!sk[72]) & (!i_6_) & (i_7_) & (!g6) & (!g8) & (!g27)) + ((!sk[72]) & (!i_6_) & (!i_7_) & (g6) & (!g8) & (!g27)) + ((!sk[72]) & (!i_6_) & (!i_7_) & (!g6) & (g8) & (!g27)) + ((!sk[72]) & (!i_6_) & (!i_7_) & (!g6) & (!g8) & (g27)) + ((!sk[72]) & (!i_6_) & (!i_7_) & (!g6) & (g8) & (!g27)) + ((!sk[72]) & (!i_6_) & (!i_7_) & (g6) & (!g8) & (!g27)));
	assign g141 = (((i_1_) & (!i_0_) & (!g50) & (g136) & (g139) & (!g140)) + ((!i_1_) & (i_0_) & (!g50) & (g136) & (g139) & (!g140)) + ((!i_1_) & (!i_0_) & (!g50) & (g136) & (g139) & (!g140)));
	assign g142 = (((!g2) & (!sk[74]) & (g6) & (!g25) & (!g50)) + ((!g2) & (!sk[74]) & (!g6) & (g25) & (!g50)) + ((!g2) & (!sk[74]) & (!g6) & (!g25) & (g50)) + ((!g2) & (!sk[74]) & (g6) & (!g25) & (!g50)));
	assign g143 = (((!g7) & (!g23) & (g78) & (!sk[75]) & (!g65) & (!g142)) + ((!g7) & (!g23) & (!g78) & (!sk[75]) & (g65) & (!g142)) + ((!g7) & (!g23) & (!g78) & (!sk[75]) & (!g65) & (g142)) + ((!g7) & (g23) & (!g78) & (!sk[75]) & (!g65) & (!g142)) + ((g7) & (!g23) & (!g78) & (sk[75]) & (!g65) & (!g142)));
	assign g144 = (((!sk[76]) & (!g2) & (g4) & (!g27) & (!g38)) + ((!sk[76]) & (!g2) & (!g4) & (g27) & (!g38)) + ((!sk[76]) & (!g2) & (!g4) & (!g27) & (g38)) + ((!sk[76]) & (!g2) & (g4) & (!g27) & (!g38)));
	assign g145 = (((!i_5_) & (g12) & (!g31) & (!sk[77]) & (!g38) & (!g144)) + ((!i_5_) & (!g12) & (!g31) & (!sk[77]) & (g38) & (!g144)) + ((!i_5_) & (!g12) & (!g31) & (!sk[77]) & (!g38) & (g144)) + ((!i_5_) & (!g12) & (g31) & (!sk[77]) & (!g38) & (!g144)) + ((!i_5_) & (!g12) & (!g31) & (sk[77]) & (!g38) & (!g144)) + ((!i_5_) & (!g12) & (!g31) & (!sk[77]) & (g38) & (!g144)));
	assign g146 = (((!i_6_) & (!i_7_) & (g8) & (i_1_) & (i_0_) & (!i_2_)) + ((!i_6_) & (i_7_) & (g8) & (!i_1_) & (!i_0_) & (!i_2_)) + ((!i_6_) & (!i_7_) & (g8) & (!i_1_) & (!i_0_) & (i_2_)) + ((!i_6_) & (i_7_) & (g8) & (!i_1_) & (!i_0_) & (i_2_)));
	assign g147 = (((!i_4_) & (i_5_) & (!i_6_) & (!i_7_) & (i_3_) & (g17)) + ((i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (i_3_) & (g17)) + ((!i_4_) & (!i_5_) & (i_6_) & (i_7_) & (i_3_) & (g17)));
	assign g148 = (((!i_6_) & (g21) & (!g27) & (!sk[80]) & (!g147)) + ((!i_6_) & (!g21) & (!g27) & (!sk[80]) & (g147)) + ((!i_6_) & (!g21) & (g27) & (!sk[80]) & (!g147)) + ((!i_6_) & (!g21) & (!g27) & (sk[80]) & (!g147)) + ((i_6_) & (!g21) & (!g27) & (sk[80]) & (!g147)));
	assign g149 = (((!i_4_) & (!i_5_) & (!i_3_) & (!i_1_) & (!i_0_) & (i_2_)) + ((!i_4_) & (!i_5_) & (!i_3_) & (i_1_) & (!i_0_) & (!i_2_)) + ((!i_4_) & (!i_5_) & (!i_3_) & (!i_1_) & (i_0_) & (!i_2_)) + ((!i_4_) & (!i_5_) & (i_3_) & (!i_1_) & (!i_0_) & (!i_2_)) + ((!i_4_) & (!i_5_) & (!i_3_) & (!i_1_) & (i_0_) & (i_2_)) + ((i_4_) & (!i_5_) & (!i_3_) & (!i_1_) & (!i_0_) & (!i_2_)) + ((i_4_) & (!i_5_) & (!i_3_) & (!i_1_) & (!i_0_) & (!i_2_)));
	assign g150 = (((!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (!g19)) + ((i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (!g19)) + ((!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (!g19)) + ((!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (!g19)) + ((!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (!g19)));
	assign g151 = (((!g343) & (g145) & (!g146) & (!g148) & (!sk[83]) & (!g333)) + ((!g343) & (!g145) & (g146) & (!g148) & (!sk[83]) & (!g333)) + ((!g343) & (!g145) & (!g146) & (g148) & (!sk[83]) & (!g333)) + ((!g343) & (!g145) & (!g146) & (!g148) & (!sk[83]) & (g333)) + ((g343) & (g145) & (!g146) & (g148) & (!sk[83]) & (g333)));
	assign g152 = (((!g128) & (!sk[84]) & (g132) & (!g141) & (!g143) & (!g151)) + ((!g128) & (!sk[84]) & (!g132) & (g141) & (!g143) & (!g151)) + ((!g128) & (!sk[84]) & (!g132) & (!g141) & (g143) & (!g151)) + ((!g128) & (!sk[84]) & (!g132) & (!g141) & (!g143) & (g151)) + ((g128) & (!sk[84]) & (g132) & (g141) & (g143) & (g151)));
	assign g153 = (((!g5) & (g16) & (!sk[85]) & (!g31) & (!g71)) + ((!g5) & (!g16) & (!sk[85]) & (!g31) & (g71)) + ((!g5) & (!g16) & (!sk[85]) & (g31) & (!g71)) + ((g5) & (!g16) & (sk[85]) & (!g31) & (!g71)));
	assign g154 = (((!sk[86]) & (!g7) & (g17) & (!g36) & (!g50) & (!g111)) + ((!sk[86]) & (!g7) & (!g17) & (!g36) & (!g50) & (g111)) + ((sk[86]) & (!g7) & (!g17) & (!g36) & (!g50) & (!g111)) + ((!sk[86]) & (!g7) & (!g17) & (g36) & (!g50) & (!g111)) + ((!sk[86]) & (!g7) & (!g17) & (!g36) & (g50) & (!g111)) + ((!sk[86]) & (g7) & (g17) & (!g36) & (!g50) & (!g111)));
	assign g155 = (((!i_4_) & (i_5_) & (!i_6_) & (!sk[87]) & (!i_3_) & (!g23)) + ((!i_4_) & (!i_5_) & (i_6_) & (!sk[87]) & (!i_3_) & (!g23)) + ((!i_4_) & (!i_5_) & (!i_6_) & (!sk[87]) & (i_3_) & (!g23)) + ((!i_4_) & (!i_5_) & (!i_6_) & (!sk[87]) & (!i_3_) & (g23)) + ((i_4_) & (i_5_) & (!i_6_) & (!sk[87]) & (!i_3_) & (!g23)) + ((i_4_) & (!i_5_) & (!i_6_) & (!sk[87]) & (i_3_) & (!g23)) + ((!i_4_) & (i_5_) & (i_6_) & (!sk[87]) & (i_3_) & (!g23)));
	assign g156 = (((!g31) & (!g41) & (!sk[88]) & (g50) & (!g155)) + ((!g31) & (!g41) & (!sk[88]) & (!g50) & (g155)) + ((g31) & (g41) & (!sk[88]) & (!g50) & (!g155)) + ((!g31) & (g41) & (!sk[88]) & (!g50) & (!g155)));
	assign g157 = (((!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (i_3_) & (!g23)) + ((i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (!g23)) + ((!i_4_) & (!i_5_) & (i_6_) & (!i_7_) & (!i_3_) & (!g23)) + ((!i_4_) & (i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (!g23)) + ((!i_4_) & (!i_5_) & (i_6_) & (i_7_) & (!i_3_) & (!g23)) + ((!i_4_) & (!i_5_) & (!i_6_) & (i_7_) & (i_3_) & (!g23)));
	assign g158 = (((g126) & (!g310) & (g153) & (g154) & (g156) & (!g157)));
	assign g159 = (((!sk[91]) & (!g15) & (g21) & (!g39) & (!g86)) + ((!sk[91]) & (!g15) & (!g21) & (g39) & (!g86)) + ((!sk[91]) & (!g15) & (!g21) & (!g39) & (g86)) + ((!sk[91]) & (!g15) & (!g21) & (!g39) & (g86)) + ((!sk[91]) & (!g15) & (!g21) & (!g39) & (g86)));
	assign g160 = (((!i_4_) & (!sk[92]) & (i_3_) & (!g13) & (!g15)) + ((!i_4_) & (!sk[92]) & (!i_3_) & (g13) & (!g15)) + ((!i_4_) & (!sk[92]) & (!i_3_) & (!g13) & (g15)) + ((!i_4_) & (!sk[92]) & (i_3_) & (g13) & (g15)));
	assign g161 = (((g38) & (!sk[93]) & (g39) & (!g79) & (!g80)) + ((!g38) & (!sk[93]) & (!g39) & (g79) & (!g80)) + ((!g38) & (!sk[93]) & (g39) & (!g79) & (!g80)) + ((!g38) & (!sk[93]) & (!g39) & (!g79) & (g80)) + ((!g38) & (!sk[93]) & (g39) & (!g79) & (g80)));
	assign g162 = (((i_4_) & (!i_5_) & (i_3_) & (!g13) & (!g15) & (g39)) + ((!i_4_) & (!i_5_) & (!i_3_) & (g13) & (!g15) & (!g39)) + ((!i_4_) & (!i_5_) & (!i_3_) & (g13) & (g15) & (!g39)) + ((!i_4_) & (i_5_) & (i_3_) & (!g13) & (g15) & (g39)));
	assign g163 = (((!sk[95]) & (!g12) & (g13) & (!g38) & (!g161) & (!g162)) + ((!sk[95]) & (!g12) & (!g13) & (!g38) & (g161) & (!g162)) + ((!sk[95]) & (!g12) & (!g13) & (!g38) & (!g161) & (g162)) + ((sk[95]) & (!g12) & (!g13) & (!g38) & (!g161) & (!g162)) + ((!sk[95]) & (!g12) & (!g13) & (g38) & (!g161) & (!g162)) + ((!sk[95]) & (!g12) & (g13) & (!g38) & (!g161) & (!g162)));
	assign g164 = (((i_6_) & (!g21) & (!g39) & (g159) & (!g160) & (g163)) + ((!i_6_) & (!g21) & (!g39) & (g159) & (!g160) & (g163)) + ((!i_6_) & (!g21) & (!g39) & (g159) & (!g160) & (g163)));
	assign g165 = (((!g32) & (g54) & (!g70) & (!g158) & (!sk[97]) & (!g164)) + ((!g32) & (!g54) & (g70) & (!g158) & (!sk[97]) & (!g164)) + ((!g32) & (!g54) & (!g70) & (g158) & (!sk[97]) & (!g164)) + ((!g32) & (!g54) & (!g70) & (!g158) & (!sk[97]) & (g164)) + ((g32) & (!g54) & (g70) & (g158) & (!sk[97]) & (g164)));
	assign g166 = (((!g17) & (!sk[98]) & (g74) & (!g75) & (!g60)) + ((!g17) & (!sk[98]) & (!g74) & (g75) & (!g60)) + ((!g17) & (!sk[98]) & (!g74) & (!g75) & (g60)) + ((!g17) & (!sk[98]) & (g74) & (g75) & (!g60)) + ((!g17) & (!sk[98]) & (g74) & (g75) & (g60)));
	assign g167 = (((!i_6_) & (i_7_) & (!g6) & (!sk[99]) & (!g21) & (!g31)) + ((!i_6_) & (!i_7_) & (g6) & (!sk[99]) & (!g21) & (!g31)) + ((!i_6_) & (!i_7_) & (!g6) & (!sk[99]) & (g21) & (!g31)) + ((!i_6_) & (!i_7_) & (!g6) & (!sk[99]) & (!g21) & (g31)) + ((!i_6_) & (i_7_) & (g6) & (!sk[99]) & (!g21) & (!g31)) + ((i_6_) & (!i_7_) & (g6) & (!sk[99]) & (!g21) & (!g31)) + ((i_6_) & (!i_7_) & (!g6) & (!sk[99]) & (g21) & (!g31)));
	assign g168 = (((!i_6_) & (g6) & (!sk[100]) & (!g23) & (!g36) & (!g117)) + ((!i_6_) & (!g6) & (!sk[100]) & (!g23) & (g36) & (!g117)) + ((!i_6_) & (!g6) & (!sk[100]) & (!g23) & (!g36) & (g117)) + ((!i_6_) & (!g6) & (!sk[100]) & (g23) & (!g36) & (!g117)) + ((!i_6_) & (!g6) & (sk[100]) & (!g23) & (!g36) & (!g117)) + ((!i_6_) & (!g6) & (sk[100]) & (!g23) & (!g36) & (!g117)));
	assign g169 = (((!g13) & (g29) & (!g82) & (!sk[101]) & (!g167) & (!g168)) + ((!g13) & (!g29) & (g82) & (!sk[101]) & (!g167) & (!g168)) + ((!g13) & (!g29) & (!g82) & (!sk[101]) & (g167) & (!g168)) + ((!g13) & (!g29) & (!g82) & (!sk[101]) & (!g167) & (g168)) + ((!g13) & (!g29) & (!g82) & (!sk[101]) & (!g167) & (g168)));
	assign g170 = (((!g13) & (g36) & (!sk[102]) & (!g95)) + ((!g13) & (!g36) & (sk[102]) & (!g95)) + ((!g13) & (!g36) & (sk[102]) & (!g95)));
	assign g171 = (((!g17) & (!sk[103]) & (g77) & (!g170)) + ((!g17) & (sk[103]) & (!g77) & (g170)) + ((!g17) & (!sk[103]) & (g77) & (g170)));
	assign g172 = (((!sk[104]) & (!g17) & (g50) & (!g73)) + ((sk[104]) & (!g17) & (!g50) & (!g73)) + ((!sk[104]) & (!g17) & (g50) & (!g73)));
	assign g173 = (((!sk[105]) & (i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!g31)) + ((!sk[105]) & (!i_4_) & (!i_5_) & (i_6_) & (!i_7_) & (!g31)) + ((!sk[105]) & (i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!g31)) + ((sk[105]) & (!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!g31)) + ((!sk[105]) & (!i_4_) & (i_5_) & (i_6_) & (i_7_) & (!g31)));
	assign g174 = (((!sk[106]) & (!g56) & (!g171) & (g172) & (!g173)) + ((!sk[106]) & (g56) & (!g171) & (!g172) & (g173)) + ((!sk[106]) & (!g56) & (g171) & (g172) & (!g173)));
	assign g175 = (((!g166) & (!sk[107]) & (!g108) & (g169) & (!g174)) + ((g166) & (!sk[107]) & (!g108) & (!g169) & (g174)) + ((g166) & (!sk[107]) & (g108) & (g169) & (g174)));
	assign g176 = (((i_5_) & (!g29) & (!g31) & (!g36) & (!sk[108]) & (!g54)) + ((!i_5_) & (!g29) & (g31) & (!g36) & (!sk[108]) & (!g54)) + ((!i_5_) & (!g29) & (g31) & (!g36) & (!sk[108]) & (!g54)) + ((i_5_) & (!g29) & (!g31) & (!g36) & (!sk[108]) & (!g54)) + ((!i_5_) & (!g29) & (!g31) & (!g36) & (sk[108]) & (!g54)));
	assign g177 = (((!sk[109]) & (!g39) & (g50) & (!g343)) + ((sk[109]) & (!g39) & (!g50) & (g343)) + ((!sk[109]) & (g39) & (!g50) & (g343)));
	assign g178 = (((i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (g19)) + ((!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (i_3_) & (g19)) + ((!i_4_) & (i_5_) & (!i_6_) & (i_7_) & (!i_3_) & (g19)) + ((!i_4_) & (i_5_) & (i_6_) & (!i_7_) & (!i_3_) & (g19)) + ((!i_4_) & (!i_5_) & (i_6_) & (!i_7_) & (i_3_) & (!g19)));
	assign g179 = (((!g20) & (!g62) & (g177) & (!sk[111]) & (!g178)) + ((g20) & (!g62) & (!g177) & (!sk[111]) & (g178)) + ((g20) & (g62) & (g177) & (!sk[111]) & (!g178)));
	assign g180 = (((g12) & (!g13) & (!g38) & (!sk[112]) & (!g39) & (!g50)) + ((!g12) & (!g13) & (g38) & (!sk[112]) & (!g39) & (!g50)) + ((!g12) & (!g13) & (!g38) & (sk[112]) & (!g39) & (!g50)) + ((!g12) & (!g13) & (!g38) & (sk[112]) & (!g39) & (!g50)) + ((!g12) & (!g13) & (!g38) & (sk[112]) & (!g39) & (!g50)));
	assign g181 = (((!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (i_3_) & (!g27)) + ((!i_4_) & (!i_5_) & (i_6_) & (!i_7_) & (i_3_) & (!g27)));
	assign g182 = (((g144) & (!sk[114]) & (!g181)) + ((!g144) & (sk[114]) & (!g181)));
	assign g183 = (((i_6_) & (!sk[115]) & (!i_7_) & (!g6) & (!g8) & (!g17)) + ((!i_6_) & (!sk[115]) & (!i_7_) & (g6) & (!g8) & (!g17)) + ((!i_6_) & (!sk[115]) & (!i_7_) & (g6) & (!g8) & (g17)) + ((i_6_) & (!sk[115]) & (i_7_) & (!g6) & (g8) & (g17)));
	assign g184 = (((g16) & (!sk[116]) & (!g17) & (g39) & (!g77)) + ((!g16) & (!sk[116]) & (!g17) & (g39) & (!g77)) + ((g16) & (!sk[116]) & (!g17) & (!g39) & (g77)) + ((!g16) & (sk[116]) & (g17) & (!g39) & (g77)));
	assign g185 = (((!i_4_) & (!i_5_) & (!i_3_) & (i_1_) & (!i_0_) & (i_2_)) + ((!i_4_) & (!i_5_) & (!i_3_) & (i_1_) & (i_0_) & (!i_2_)) + ((i_4_) & (!i_5_) & (!i_3_) & (!i_1_) & (i_0_) & (!i_2_)) + ((i_4_) & (!i_5_) & (i_3_) & (i_1_) & (!i_0_) & (!i_2_)));
	assign g186 = (((g17) & (!g60) & (!g183) & (!sk[118]) & (!g184) & (!g185)) + ((!g17) & (!g60) & (g183) & (!sk[118]) & (!g184) & (!g185)) + ((!g17) & (!g60) & (!g183) & (sk[118]) & (!g184) & (!g185)) + ((!g17) & (g60) & (!g183) & (sk[118]) & (!g184) & (!g185)));
	assign g187 = (((g129) & (!g153) & (!g180) & (!g182) & (!sk[119]) & (!g186)) + ((!g129) & (!g153) & (g180) & (!g182) & (!sk[119]) & (!g186)) + ((!g129) & (g153) & (g180) & (g182) & (!sk[119]) & (g186)));
	assign g188 = (((g128) & (!g176) & (!sk[120]) & (!g90) & (!g179) & (!g187)) + ((!g128) & (!g176) & (!sk[120]) & (g90) & (!g179) & (!g187)) + ((g128) & (g176) & (!sk[120]) & (g90) & (g179) & (g187)));
	assign g189 = (((!i_6_) & (!g8) & (!sk[121]) & (g31) & (!g38)) + ((!i_6_) & (!g8) & (sk[121]) & (!g31) & (g38)) + ((!i_6_) & (g8) & (sk[121]) & (!g31) & (!g38)) + ((i_6_) & (!g8) & (!sk[121]) & (!g31) & (g38)));
	assign g190 = (((!g57) & (!g189) & (g88) & (!sk[122]) & (!g158)) + ((g57) & (!g189) & (!g88) & (!sk[122]) & (g158)) + ((g57) & (!g189) & (!g88) & (!sk[122]) & (g158)));
	assign g191 = (((!sk[123]) & (!g21) & (!g39) & (g87) & (!g178)) + ((!sk[123]) & (g21) & (!g39) & (!g87) & (g178)) + ((!sk[123]) & (!g21) & (!g39) & (g87) & (!g178)) + ((!sk[123]) & (!g21) & (!g39) & (g87) & (!g178)));
	assign g192 = (((g5) & (!g19) & (!g25) & (!g44) & (!sk[124]) & (!g130)) + ((!g5) & (!g19) & (g25) & (!g44) & (!sk[124]) & (!g130)) + ((g5) & (!g19) & (g25) & (!g44) & (!sk[124]) & (g130)) + ((!g5) & (!g19) & (g25) & (!g44) & (!sk[124]) & (g130)) + ((g5) & (!g19) & (!g25) & (!g44) & (!sk[124]) & (g130)) + ((!g5) & (!g19) & (!g25) & (!g44) & (sk[124]) & (g130)));
	assign g193 = (((g20) & (!g55) & (!g133) & (!sk[125]) & (!g182) & (!g192)) + ((!g20) & (!g55) & (g133) & (!sk[125]) & (!g182) & (!g192)) + ((g20) & (!g55) & (!g133) & (!sk[125]) & (g182) & (g192)));
	assign g194 = (((g139) & (!sk[126]) & (!g190) & (!g191) & (!g322) & (!g193)) + ((!g139) & (!sk[126]) & (!g190) & (g191) & (!g322) & (!g193)) + ((g139) & (!sk[126]) & (g190) & (g191) & (g322) & (g193)));
	assign g195 = (((i_4_) & (!i_5_) & (!sk[127]) & (!i_3_) & (!g13) & (!g39)) + ((!i_4_) & (!i_5_) & (!sk[127]) & (i_3_) & (!g13) & (!g39)) + ((i_4_) & (!i_5_) & (!sk[127]) & (i_3_) & (!g13) & (g39)) + ((!i_4_) & (!i_5_) & (sk[127]) & (!i_3_) & (g13) & (!g39)));
	assign g196 = (((g16) & (!g29) & (!sk[0]) & (!g31) & (!g39) & (!g195)) + ((!g16) & (!g29) & (!sk[0]) & (g31) & (!g39) & (!g195)) + ((!g16) & (!g29) & (!sk[0]) & (g31) & (!g39) & (!g195)) + ((!g16) & (!g29) & (!sk[0]) & (g31) & (!g39) & (!g195)) + ((!g16) & (!g29) & (sk[0]) & (!g31) & (!g39) & (!g195)) + ((!g16) & (!g29) & (sk[0]) & (!g31) & (!g39) & (!g195)));
	assign g197 = (((!i_6_) & (!i_7_) & (!sk[1]) & (g4) & (!g31)) + ((i_6_) & (!i_7_) & (!sk[1]) & (!g4) & (g31)) + ((!i_6_) & (i_7_) & (!sk[1]) & (g4) & (!g31)) + ((i_6_) & (!i_7_) & (!sk[1]) & (g4) & (!g31)));
	assign g198 = (((g13) & (!g77) & (!g197) & (!g63) & (!sk[2]) & (!g180)) + ((!g13) & (!g77) & (g197) & (!g63) & (!sk[2]) & (!g180)) + ((!g13) & (!g77) & (!g197) & (!g63) & (sk[2]) & (g180)) + ((!g13) & (!g77) & (!g197) & (!g63) & (sk[2]) & (g180)));
	assign g199 = (((g61) & (!sk[3]) & (!g172) & (!g103) & (!g196) & (!g198)) + ((!g61) & (!sk[3]) & (!g172) & (g103) & (!g196) & (!g198)) + ((!g61) & (!sk[3]) & (g172) & (g103) & (g196) & (g198)));
	assign g200 = (((!g12) & (!g23) & (!sk[4]) & (g27) & (!g60)) + ((g12) & (!g23) & (!sk[4]) & (!g27) & (g60)) + ((!g12) & (!g23) & (sk[4]) & (!g27) & (!g60)) + ((g12) & (!g23) & (sk[4]) & (!g27) & (!g60)));
	assign g201 = (((g16) & (!g25) & (!g38) & (!sk[5]) & (!g189) & (!g200)) + ((!g16) & (!g25) & (g38) & (!sk[5]) & (!g189) & (!g200)) + ((!g16) & (!g25) & (!g38) & (sk[5]) & (!g189) & (!g200)) + ((!g16) & (g25) & (!g38) & (sk[5]) & (!g189) & (!g200)));
	assign g202 = (((i_6_) & (i_7_) & (!g6) & (!g21) & (!g27) & (!g137)) + ((!i_6_) & (!i_7_) & (!g6) & (!g21) & (!g27) & (!g137)) + ((!i_6_) & (i_7_) & (!g6) & (!g21) & (!g27) & (!g137)) + ((!i_6_) & (!i_7_) & (!g6) & (!g21) & (!g27) & (!g137)) + ((!i_6_) & (!i_7_) & (!g6) & (!g21) & (g27) & (!g137)));
	assign g203 = (((!sk[7]) & (!g21) & (g38) & (!g39)) + ((!sk[7]) & (g21) & (!g38) & (g39)) + ((!sk[7]) & (!g21) & (g38) & (g39)));
	assign g204 = (((i_5_) & (!g16) & (!g23) & (!g27) & (!g38) & (!g203)) + ((!i_5_) & (!g16) & (g23) & (g27) & (!g38) & (!g203)) + ((!i_5_) & (!g16) & (!g23) & (!g27) & (!g38) & (!g203)));
	assign g205 = (((!g12) & (g25) & (g27) & (!g29) & (!g36) & (g204)) + ((!g12) & (!g25) & (!g27) & (!g29) & (!g36) & (g204)) + ((!g12) & (g25) & (!g27) & (!g29) & (!g36) & (g204)));
	assign g206 = (((!sk[10]) & (g48) & (!g95) & (!g184) & (!g116) & (!g205)) + ((!sk[10]) & (!g48) & (!g95) & (g184) & (!g116) & (!g205)) + ((sk[10]) & (!g48) & (!g95) & (!g184) & (g116) & (g205)));
	assign g207 = (((g166) & (g199) & (g311) & (g201) & (g202) & (g206)));
	assign g208 = (((!g12) & (!sk[12]) & (g25) & (!g38)) + ((g12) & (sk[12]) & (!g25) & (!g38)) + ((!g12) & (sk[12]) & (!g25) & (g38)) + ((g12) & (!sk[12]) & (!g25) & (g38)));
	assign g209 = (((!g110) & (!sk[13]) & (g135) & (!g208)) + ((g110) & (!sk[13]) & (!g135) & (g208)) + ((g110) & (sk[13]) & (!g135) & (!g208)));
	assign g210 = (((!sk[14]) & (!g49) & (g144) & (!g111)) + ((!sk[14]) & (g49) & (!g144) & (g111)) + ((sk[14]) & (g49) & (!g144) & (!g111)));
	assign g211 = (((!sk[15]) & (!g12) & (!g27) & (g29) & (!g36)) + ((!sk[15]) & (!g12) & (!g27) & (g29) & (!g36)) + ((sk[15]) & (g12) & (!g27) & (!g29) & (!g36)) + ((!sk[15]) & (g12) & (!g27) & (!g29) & (g36)) + ((sk[15]) & (!g12) & (!g27) & (!g29) & (g36)));
	assign g212 = (((!i_4_) & (!i_5_) & (!i_6_) & (!i_3_) & (!g25) & (g32)) + ((!i_4_) & (!i_5_) & (!i_6_) & (!i_3_) & (g25) & (g32)) + ((!i_4_) & (!i_5_) & (!i_6_) & (!i_3_) & (!g25) & (g32)) + ((!i_4_) & (!i_5_) & (!i_6_) & (!i_3_) & (!g25) & (g32)));
	assign g213 = (((g26) & (!g85) & (!g134) & (!g211) & (!g89) & (g212)));
	assign g214 = (((g169) & (!g199) & (!g209) & (!sk[18]) & (!g210) & (!g213)) + ((!g169) & (!g199) & (g209) & (!sk[18]) & (!g210) & (!g213)) + ((g169) & (g199) & (g209) & (!sk[18]) & (g210) & (g213)));
	assign g215 = (((i_4_) & (!i_3_) & (!i_1_) & (!i_0_) & (!i_2_) & (!g1)) + ((!i_4_) & (!i_3_) & (!i_1_) & (i_0_) & (!i_2_) & (g1)));
	assign g216 = (((i_4_) & (!i_3_) & (!g12) & (!sk[20]) & (!g13) & (!g15)) + ((!i_4_) & (!i_3_) & (g12) & (!sk[20]) & (!g13) & (!g15)) + ((!i_4_) & (!i_3_) & (g12) & (!sk[20]) & (g13) & (!g15)) + ((!i_4_) & (i_3_) & (!g12) & (sk[20]) & (g13) & (g15)));
	assign g217 = (((!sk[21]) & (!g13) & (g38) & (!g216)) + ((!sk[21]) & (g13) & (!g38) & (g216)) + ((sk[21]) & (!g13) & (!g38) & (!g216)) + ((!sk[21]) & (!g13) & (g38) & (!g216)));
	assign g218 = (((!g171) & (!sk[22]) & (!g87) & (g162) & (!g217)) + ((g171) & (!sk[22]) & (!g87) & (!g162) & (g217)) + ((g171) & (!sk[22]) & (g87) & (!g162) & (g217)));
	assign g219 = (((!sk[23]) & (!g31) & (g44) & (!g176)) + ((!sk[23]) & (g31) & (!g44) & (g176)) + ((sk[23]) & (!g31) & (!g44) & (g176)));
	assign g220 = (((!g23) & (!g31) & (g41) & (!sk[24]) & (!g50)) + ((!g23) & (!g31) & (g41) & (!sk[24]) & (!g50)) + ((g23) & (g31) & (g41) & (!sk[24]) & (!g50)) + ((g23) & (!g31) & (!g41) & (!sk[24]) & (g50)));
	assign g221 = (((!g39) & (!sk[25]) & (!g115) & (g189) & (!g220)) + ((g39) & (!sk[25]) & (!g115) & (!g189) & (g220)) + ((!g39) & (sk[25]) & (!g115) & (!g189) & (g220)) + ((!g39) & (sk[25]) & (!g115) & (!g189) & (g220)));
	assign g222 = (((i_6_) & (!g21) & (!g23) & (!sk[26]) & (!g153) & (!g24)) + ((!i_6_) & (!g21) & (g23) & (!sk[26]) & (!g153) & (!g24)) + ((!i_6_) & (!g21) & (g23) & (!sk[26]) & (g153) & (!g24)) + ((!i_6_) & (!g21) & (!g23) & (sk[26]) & (g153) & (!g24)) + ((!i_6_) & (!g21) & (!g23) & (sk[26]) & (g153) & (!g24)));
	assign g223 = (((!g17) & (g218) & (g219) & (g70) & (g221) & (g222)));
	assign g224 = (((i_4_) & (!i_5_) & (!sk[28]) & (!i_3_) & (!g9) & (!g17)) + ((!i_4_) & (!i_5_) & (!sk[28]) & (i_3_) & (!g9) & (!g17)) + ((i_4_) & (!i_5_) & (!sk[28]) & (!i_3_) & (!g9) & (g17)) + ((!i_4_) & (!i_5_) & (sk[28]) & (!i_3_) & (!g9) & (g17)));
	assign g225 = (((g51) & (!sk[29]) & (!g53)) + ((g51) & (!sk[29]) & (g53)));
	assign g226 = (((!sk[30]) & (g62) & (!g101)) + ((!sk[30]) & (g62) & (!g101)));
	assign g227 = (((g20) & (!g23) & (!g25) & (!g36) & (!sk[31]) & (!g50)) + ((!g20) & (!g23) & (g25) & (!g36) & (!sk[31]) & (!g50)) + ((g20) & (g23) & (g25) & (!g36) & (!sk[31]) & (!g50)) + ((g20) & (g23) & (!g25) & (!g36) & (!sk[31]) & (!g50)) + ((g20) & (!g23) & (g25) & (!g36) & (!sk[31]) & (!g50)) + ((g20) & (!g23) & (!g25) & (!g36) & (!sk[31]) & (!g50)));
	assign g228 = (((!g7) & (!g19) & (!sk[32]) & (g27) & (!g36)) + ((!g7) & (!g19) & (sk[32]) & (!g27) & (!g36)) + ((g7) & (!g19) & (!sk[32]) & (!g27) & (g36)) + ((!g7) & (g19) & (sk[32]) & (!g27) & (g36)));
	assign g229 = (((g26) & (!g63) & (!g211) & (!g208) & (!g76) & (!g228)));
	assign g230 = (((!g71) & (g225) & (g226) & (g143) & (g227) & (g229)));
	assign g231 = (((i_6_) & (!sk[35]) & (!i_7_) & (!g6) & (!g8) & (!g31)) + ((!i_6_) & (!sk[35]) & (!i_7_) & (g6) & (!g8) & (!g31)) + ((i_6_) & (!sk[35]) & (i_7_) & (!g6) & (g8) & (!g31)));
	assign g232 = (((g12) & (!sk[36]) & (!g38) & (g39) & (!g115)) + ((!g12) & (!sk[36]) & (!g38) & (g39) & (!g115)) + ((!g12) & (!sk[36]) & (g38) & (g39) & (!g115)) + ((!g12) & (!sk[36]) & (!g38) & (g39) & (g115)) + ((g12) & (!sk[36]) & (!g38) & (!g39) & (g115)));
	assign g233 = (((g138) & (!g145) & (!sk[37]) & (!g311) & (!g231) & (!g232)) + ((!g138) & (!g145) & (!sk[37]) & (g311) & (!g231) & (!g232)) + ((!g138) & (g145) & (!sk[37]) & (g311) & (!g231) & (!g232)));
	assign g234 = (((g49) & (g86) & (!g73) & (!g137) & (!g24) & (g154)));
	assign g235 = (((g58) & (!g136) & (!sk[39]) & (!g230) & (!g233) & (!g234)) + ((!g58) & (!g136) & (!sk[39]) & (g230) & (!g233) & (!g234)) + ((g58) & (g136) & (!sk[39]) & (g230) & (g233) & (g234)));
	assign g236 = (((i_3_) & (!g39) & (!g137) & (g219) & (g70) & (g190)) + ((!i_3_) & (!g39) & (!g137) & (g219) & (g70) & (g190)));
	assign g237 = (((g13) & (g38) & (!sk[41]) & (!g1)) + ((!g13) & (g38) & (!sk[41]) & (!g1)) + ((g13) & (!g38) & (!sk[41]) & (g1)));
	assign g238 = (((!i_3_) & (!sk[42]) & (i_1_) & (!i_0_)) + ((!i_3_) & (sk[42]) & (!i_1_) & (i_0_)) + ((i_3_) & (!sk[42]) & (!i_1_) & (i_0_)));
	assign g239 = (((i_4_) & (!i_5_) & (!i_2_) & (!g15) & (!sk[43]) & (!g238)) + ((!i_4_) & (!i_5_) & (i_2_) & (!g15) & (!sk[43]) & (!g238)) + ((!i_4_) & (!i_5_) & (!i_2_) & (g15) & (sk[43]) & (!g238)));
	assign g240 = (((!g138) & (!g145) & (!sk[44]) & (g311) & (!g231)) + ((g138) & (!g145) & (!sk[44]) & (!g311) & (g231)) + ((!g138) & (g145) & (!sk[44]) & (g311) & (!g231)));
	assign g241 = (((!sk[45]) & (!i_6_) & (!g19) & (g21) & (!g62)) + ((sk[45]) & (!i_6_) & (!g19) & (!g21) & (g62)) + ((!sk[45]) & (i_6_) & (!g19) & (!g21) & (g62)) + ((!sk[45]) & (i_6_) & (!g19) & (!g21) & (g62)));
	assign g242 = (((g12) & (!g25) & (!g29) & (!sk[46]) & (!g36) & (!g50)) + ((!g12) & (!g25) & (g29) & (!sk[46]) & (!g36) & (!g50)) + ((g12) & (!g25) & (!g29) & (!sk[46]) & (!g36) & (!g50)) + ((!g12) & (!g25) & (g29) & (!sk[46]) & (!g36) & (!g50)) + ((!g12) & (!g25) & (!g29) & (sk[46]) & (g36) & (!g50)) + ((!g12) & (!g25) & (!g29) & (sk[46]) & (!g36) & (g50)));
	assign g243 = (((!g181) & (!sk[47]) & (g241) & (!g242)) + ((g181) & (!sk[47]) & (!g241) & (g242)) + ((!g181) & (!sk[47]) & (g241) & (!g242)));
	assign g244 = (((!sk[48]) & (!g16) & (g21) & (!g38)) + ((!sk[48]) & (g16) & (!g21) & (g38)) + ((sk[48]) & (!g16) & (!g21) & (!g38)));
	assign g245 = (((!sk[49]) & (i_4_) & (!i_5_) & (!i_3_) & (!g15) & (!g19)) + ((!sk[49]) & (!i_4_) & (!i_5_) & (i_3_) & (!g15) & (!g19)) + ((!sk[49]) & (!i_4_) & (!i_5_) & (i_3_) & (g15) & (g19)) + ((sk[49]) & (!i_4_) & (i_5_) & (!i_3_) & (g15) & (g19)));
	assign g246 = (((g19) & (!sk[50]) & (!g29) & (!g39) & (!g244) & (!g245)) + ((!g19) & (!sk[50]) & (!g29) & (g39) & (!g244) & (!g245)) + ((!g19) & (sk[50]) & (!g29) & (!g39) & (!g244) & (!g245)) + ((!g19) & (sk[50]) & (!g29) & (!g39) & (!g244) & (!g245)) + ((!g19) & (!sk[50]) & (!g29) & (g39) & (g244) & (!g245)));
	assign g247 = (((g97) & (!g84) & (!sk[51]) & (!g240) & (!g243) & (!g309)) + ((!g97) & (!g84) & (!sk[51]) & (g240) & (!g243) & (!g309)) + ((g97) & (g84) & (!sk[51]) & (g240) & (g243) & (g309)));
	assign g248 = (((!i_4_) & (!i_3_) & (g13) & (!sk[52]) & (!g15)) + ((i_4_) & (!i_3_) & (!g13) & (!sk[52]) & (g15)) + ((!i_4_) & (!i_3_) & (g13) & (!sk[52]) & (g15)));
	assign g249 = (((i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (i_3_) & (g19)) + ((!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (i_3_) & (g19)) + ((!i_4_) & (!i_5_) & (i_6_) & (i_7_) & (i_3_) & (g19)) + ((!i_4_) & (!i_5_) & (i_6_) & (!i_7_) & (i_3_) & (!g19)));
	assign g250 = (((i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (!g31)) + ((i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (!g31)) + ((!i_4_) & (i_5_) & (!i_6_) & (!i_7_) & (i_3_) & (!g31)) + ((!i_4_) & (i_5_) & (i_6_) & (i_7_) & (i_3_) & (!g31)) + ((!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (i_3_) & (!g31)) + ((!i_4_) & (i_5_) & (!i_6_) & (!i_7_) & (!i_3_) & (!g31)));
	assign g251 = (((!g9) & (!g13) & (!sk[55]) & (g19) & (!g21)) + ((g9) & (g13) & (!sk[55]) & (!g19) & (g21)) + ((g9) & (!g13) & (!sk[55]) & (!g19) & (g21)) + ((g9) & (!g13) & (!sk[55]) & (g19) & (g21)));
	assign g252 = (((!g249) & (!sk[56]) & (!g156) & (g250) & (!g251)) + ((g249) & (!sk[56]) & (!g156) & (!g250) & (g251)) + ((!g249) & (sk[56]) & (g156) & (!g250) & (!g251)));
	assign g253 = (((!sk[57]) & (g71) & (!g225) & (!g114) & (!g227) & (!g252)) + ((!sk[57]) & (!g71) & (!g225) & (g114) & (!g227) & (!g252)) + ((!sk[57]) & (!g71) & (g225) & (g114) & (g227) & (g252)));
	assign g254 = (((!sk[58]) & (g7) & (!g17) & (!g50) & (!g62) & (!g142)) + ((!sk[58]) & (!g7) & (!g17) & (g50) & (!g62) & (!g142)) + ((sk[58]) & (!g7) & (!g17) & (!g50) & (g62) & (!g142)) + ((!sk[58]) & (g7) & (!g17) & (!g50) & (g62) & (!g142)));
	assign g255 = (((g2) & (!g4) & (!sk[59]) & (!g27) & (!g29) & (!g36)) + ((!g2) & (!g4) & (!sk[59]) & (g27) & (!g29) & (!g36)) + ((!g2) & (!g4) & (sk[59]) & (!g27) & (g29) & (!g36)) + ((!g2) & (!g4) & (sk[59]) & (!g27) & (!g29) & (g36)) + ((!g2) & (g4) & (sk[59]) & (!g27) & (!g29) & (!g36)));
	assign g256 = (((!sk[60]) & (!g29) & (!g39) & (g244) & (!g255)) + ((!sk[60]) & (g29) & (!g39) & (!g244) & (g255)) + ((sk[60]) & (!g29) & (!g39) & (!g244) & (!g255)) + ((!sk[60]) & (!g29) & (!g39) & (g244) & (!g255)));
	assign g257 = (((!g248) & (g98) & (g141) & (g253) & (g254) & (g256)));
	assign g258 = (((!g13) & (!g21) & (!g39) & (!g50) & (g170) & (g163)) + ((!g13) & (!g21) & (!g39) & (!g50) & (g170) & (g163)) + ((!g13) & (!g21) & (!g39) & (!g50) & (g170) & (g163)) + ((!g13) & (!g21) & (!g39) & (!g50) & (g170) & (g163)));
	assign g259 = (((g10) & (!g17) & (!g38) & (!g183) & (!sk[63]) & (!g142)) + ((!g10) & (!g17) & (g38) & (!g183) & (!sk[63]) & (!g142)) + ((g10) & (!g17) & (!g38) & (!g183) & (!sk[63]) & (!g142)) + ((g10) & (!g17) & (!g38) & (!g183) & (!sk[63]) & (!g142)));
	assign g260 = (((!i_6_) & (!g16) & (!sk[64]) & (g21) & (!g23)) + ((i_6_) & (!g16) & (!sk[64]) & (!g21) & (g23)) + ((!i_6_) & (g16) & (sk[64]) & (!g21) & (!g23)) + ((i_6_) & (!g16) & (!sk[64]) & (g21) & (!g23)));
	assign g261 = (((g219) & (!g226) & (!sk[65]) & (!g245) & (!g259) & (!g260)) + ((!g219) & (!g226) & (!sk[65]) & (g245) & (!g259) & (!g260)) + ((g219) & (g226) & (!sk[65]) & (!g245) & (g259) & (!g260)));
	assign g262 = (((g105) & (!g132) & (!g201) & (!sk[66]) & (!g258) & (!g261)) + ((!g105) & (!g132) & (g201) & (!sk[66]) & (!g258) & (!g261)) + ((!g105) & (g132) & (g201) & (!sk[66]) & (g258) & (g261)));
	assign g263 = (((!sk[67]) & (i_6_) & (!i_7_) & (!g6) & (!g27) & (!g31)) + ((!sk[67]) & (!i_6_) & (!i_7_) & (g6) & (!g27) & (!g31)) + ((!sk[67]) & (i_6_) & (i_7_) & (!g6) & (g27) & (g31)) + ((sk[67]) & (!i_6_) & (!i_7_) & (!g6) & (g27) & (g31)));
	assign g264 = (((!i_6_) & (!i_7_) & (!g8) & (!g21) & (g27) & (g263)) + ((i_6_) & (i_7_) & (!g8) & (!g21) & (!g27) & (g263)) + ((i_6_) & (!i_7_) & (!g8) & (!g21) & (!g27) & (g263)) + ((!i_6_) & (!i_7_) & (!g8) & (!g21) & (!g27) & (g263)));
	assign g265 = (((!g25) & (!sk[69]) & (g36) & (!g264)) + ((g25) & (!sk[69]) & (!g36) & (g264)) + ((!g25) & (sk[69]) & (!g36) & (g264)));
	assign g266 = (((!g18) & (!sk[70]) & (g47) & (!g118)) + ((g18) & (!sk[70]) & (!g47) & (g118)) + ((g18) & (!sk[70]) & (g47) & (!g118)));
	assign g267 = (((g23) & (!g50) & (!g101) & (!g130) & (!sk[71]) & (!g266)) + ((!g23) & (!g50) & (g101) & (!g130) & (!sk[71]) & (!g266)) + ((g23) & (!g50) & (!g101) & (g130) & (!sk[71]) & (g266)) + ((!g23) & (!g50) & (!g101) & (g130) & (sk[71]) & (g266)));
	assign g268 = (((i_4_) & (!i_5_) & (i_3_) & (g13) & (!g15) & (!g17)) + ((!i_4_) & (i_5_) & (i_3_) & (g13) & (g15) & (!g17)) + ((!i_4_) & (!i_5_) & (!i_3_) & (!g13) & (g15) & (g17)));
	assign g269 = (((g125) & (!g88) & (!g195) & (!sk[73]) & (!g209) & (!g268)) + ((!g125) & (!g88) & (g195) & (!sk[73]) & (!g209) & (!g268)) + ((!g125) & (!g88) & (!g195) & (sk[73]) & (g209) & (!g268)));
	assign g270 = (((g265) & (!sk[74]) & (!g191) & (!g254) & (!g267) & (!g269)) + ((!g265) & (!sk[74]) & (!g191) & (g254) & (!g267) & (!g269)) + ((g265) & (!sk[74]) & (g191) & (g254) & (g267) & (g269)));
	assign g271 = (((!g15) & (!g21) & (g39) & (!sk[75]) & (!g268)) + ((g15) & (!g21) & (!g39) & (!sk[75]) & (g268)) + ((!g15) & (!g21) & (!g39) & (sk[75]) & (!g268)) + ((!g15) & (!g21) & (!g39) & (sk[75]) & (!g268)) + ((!g15) & (!g21) & (!g39) & (sk[75]) & (!g268)));
	assign g272 = (((!g219) & (!g221) & (!sk[76]) & (g266) & (!g271)) + ((g219) & (!g221) & (!sk[76]) & (!g266) & (g271)) + ((g219) & (g221) & (!sk[76]) & (g266) & (g271)));
	assign g273 = (((!g16) & (!g38) & (!g39) & (!g60) & (!g105) & (!g101)) + ((!g16) & (!g38) & (!g39) & (g60) & (!g105) & (!g101)));
	assign g274 = (((!sk[78]) & (i_4_) & (!i_3_) & (!g16) & (!g19) & (!g25)) + ((!sk[78]) & (!i_4_) & (!i_3_) & (g16) & (!g19) & (!g25)) + ((!sk[78]) & (!i_4_) & (!i_3_) & (g16) & (!g19) & (!g25)) + ((!sk[78]) & (i_4_) & (i_3_) & (!g16) & (g19) & (!g25)) + ((!sk[78]) & (i_4_) & (!i_3_) & (!g16) & (!g19) & (!g25)));
	assign g275 = (((!sk[79]) & (g142) & (!g183) & (!g222) & (!g273) & (!g274)) + ((!sk[79]) & (!g142) & (!g183) & (g222) & (!g273) & (!g274)) + ((!sk[79]) & (!g142) & (!g183) & (g222) & (g273) & (!g274)));
	assign g276 = (((g59) & (!g64) & (!g177) & (!g272) & (!sk[80]) & (!g275)) + ((!g59) & (!g64) & (g177) & (!g272) & (!sk[80]) & (!g275)) + ((!g59) & (g64) & (g177) & (g272) & (!sk[80]) & (g275)));
	assign g277 = (((!i_6_) & (!sk[81]) & (g17) & (!g21)) + ((i_6_) & (!sk[81]) & (!g17) & (g21)) + ((!i_6_) & (!sk[81]) & (g17) & (g21)));
	assign g278 = (((i_4_) & (!i_3_) & (!i_1_) & (!i_0_) & (!i_2_) & (!g79)) + ((!i_4_) & (!i_3_) & (!i_1_) & (!i_0_) & (!i_2_) & (!g79)) + ((i_4_) & (i_3_) & (i_1_) & (!i_0_) & (i_2_) & (!g79)));
	assign g279 = (((g12) & (!g23) & (!g39) & (!g80) & (!sk[83]) & (!g278)) + ((!g12) & (!g23) & (g39) & (!g80) & (!sk[83]) & (!g278)) + ((!g12) & (!g23) & (!g39) & (!g80) & (sk[83]) & (!g278)) + ((!g12) & (g23) & (!g39) & (!g80) & (sk[83]) & (!g278)) + ((!g12) & (!g23) & (!g39) & (!g80) & (sk[83]) & (!g278)) + ((!g12) & (g23) & (!g39) & (!g80) & (sk[83]) & (!g278)));
	assign g280 = (((g85) & (!g71) & (!g277) & (!sk[84]) & (!g125) & (!g279)) + ((!g85) & (!g71) & (g277) & (!sk[84]) & (!g125) & (!g279)) + ((!g85) & (!g71) & (!g277) & (sk[84]) & (!g125) & (g279)));
	assign g281 = (((g74) & (!sk[85]) & (!g70) & (!g196) & (!g272) & (!g280)) + ((!g74) & (!sk[85]) & (!g70) & (g196) & (!g272) & (!g280)) + ((g74) & (!sk[85]) & (g70) & (g196) & (g272) & (g280)));
	assign g282 = (((!g73) & (!sk[86]) & (g74) & (!g75)) + ((g73) & (!sk[86]) & (!g74) & (g75)) + ((!g73) & (!sk[86]) & (g74) & (g75)));
	assign g283 = (((!g2) & (!g6) & (!sk[87]) & (g25) & (!g38)) + ((!g2) & (!g6) & (sk[87]) & (!g25) & (g38)) + ((!g2) & (g6) & (sk[87]) & (!g25) & (!g38)) + ((g2) & (!g6) & (!sk[87]) & (!g25) & (g38)));
	assign g284 = (((!i_4_) & (!i_3_) & (g13) & (!sk[88]) & (!g23)) + ((i_4_) & (i_3_) & (g13) & (!sk[88]) & (!g23)) + ((i_4_) & (!i_3_) & (!g13) & (!sk[88]) & (g23)) + ((i_4_) & (!i_3_) & (!g13) & (sk[88]) & (!g23)));
	assign g285 = (((!g26) & (!sk[89]) & (g283) & (!g284)) + ((g26) & (!sk[89]) & (!g283) & (g284)) + ((g26) & (sk[89]) & (!g283) & (!g284)));
	assign g286 = (((!i_6_) & (!i_7_) & (!g6) & (g8) & (g17) & (!g23)) + ((!i_6_) & (i_7_) & (!g6) & (g8) & (g17) & (!g23)) + ((!i_6_) & (!i_7_) & (g6) & (!g8) & (!g17) & (!g23)) + ((!i_6_) & (!i_7_) & (!g6) & (g8) & (!g17) & (!g23)));
	assign g287 = (((!sk[91]) & (g39) & (!g60) & (!g244) & (!g285) & (!g286)) + ((!sk[91]) & (!g39) & (!g60) & (g244) & (!g285) & (!g286)) + ((sk[91]) & (!g39) & (!g60) & (!g244) & (g285) & (!g286)) + ((!sk[91]) & (!g39) & (g60) & (g244) & (g285) & (!g286)));
	assign g288 = (((g282) & (!sk[92]) & (!g264) & (!g179) & (!g267) & (!g287)) + ((!g282) & (!sk[92]) & (!g264) & (g179) & (!g267) & (!g287)) + ((g282) & (!sk[92]) & (g264) & (g179) & (g267) & (g287)));
	assign g289 = (((!g17) & (!g60) & (!sk[93]) & (g127) & (!g147)) + ((g17) & (!g60) & (!sk[93]) & (!g127) & (g147)) + ((!g17) & (!g60) & (!sk[93]) & (g127) & (!g147)) + ((!g17) & (g60) & (!sk[93]) & (g127) & (!g147)));
	assign g290 = (((!g21) & (g33) & (!sk[94]) & (!g39)) + ((!g21) & (g33) & (!sk[94]) & (!g39)) + ((g21) & (!g33) & (!sk[94]) & (g39)));
	assign g291 = (((g218) & (!g230) & (!g240) & (!g289) & (!sk[95]) & (!g290)) + ((!g218) & (!g230) & (g240) & (!g289) & (!sk[95]) & (!g290)) + ((g218) & (g230) & (g240) & (g289) & (!sk[95]) & (g290)));
	assign g292 = (((i_6_) & (!i_7_) & (!g8) & (!g17) & (!sk[96]) & (!g21)) + ((!i_6_) & (!i_7_) & (g8) & (!g17) & (!sk[96]) & (!g21)) + ((!i_6_) & (i_7_) & (g8) & (g17) & (!sk[96]) & (!g21)) + ((!i_6_) & (!i_7_) & (!g8) & (g17) & (sk[96]) & (g21)) + ((!i_6_) & (!i_7_) & (!g8) & (g17) & (sk[96]) & (g21)));
	assign g293 = (((!i_5_) & (!sk[97]) & (!g17) & (g38) & (!g79)) + ((i_5_) & (!sk[97]) & (g17) & (g38) & (!g79)) + ((i_5_) & (!sk[97]) & (!g17) & (!g38) & (g79)) + ((!i_5_) & (sk[97]) & (g17) & (!g38) & (!g79)));
	assign g294 = (((i_4_) & (i_5_) & (!i_3_) & (!g15) & (!g17) & (!g27)) + ((!i_4_) & (i_5_) & (!i_3_) & (g15) & (g17) & (!g27)) + ((!i_4_) & (i_5_) & (i_3_) & (g15) & (!g17) & (!g27)));
	assign g295 = (((i_4_) & (!i_5_) & (!i_3_) & (g13) & (!g15) & (!g17)) + ((i_4_) & (!i_5_) & (!i_3_) & (!g13) & (!g15) & (g17)) + ((!i_4_) & (i_5_) & (!i_3_) & (g13) & (g15) & (!g17)));
	assign g296 = (((!g293) & (!sk[100]) & (!g216) & (g294) & (!g295)) + ((g293) & (!sk[100]) & (!g216) & (!g294) & (g295)) + ((!g293) & (sk[100]) & (!g216) & (!g294) & (!g295)));
	assign g297 = (((g117) & (!g62) & (!g283) & (!g292) & (!sk[101]) & (!g296)) + ((!g117) & (!g62) & (g283) & (!g292) & (!sk[101]) & (!g296)) + ((!g117) & (g62) & (!g283) & (!g292) & (sk[101]) & (g296)));
	assign g298 = (((!sk[102]) & (!g100) & (!g253) & (g273) & (!g297)) + ((!sk[102]) & (g100) & (!g253) & (!g273) & (g297)) + ((!sk[102]) & (g100) & (g253) & (g273) & (g297)));
	assign g299 = (((!sk[103]) & (!g20) & (g26) & (!g249)) + ((!sk[103]) & (g20) & (!g26) & (g249)) + ((!sk[103]) & (g20) & (g26) & (!g249)));
	assign g300 = (((g84) & (!g240) & (!sk[104]) & (!g243) & (!g258) & (!g308)) + ((!g84) & (!g240) & (!sk[104]) & (g243) & (!g258) & (!g308)) + ((g84) & (g240) & (!sk[104]) & (g243) & (g258) & (g308)));
	assign g301 = (((!g10) & (g51) & (!sk[105]) & (!g118)) + ((g10) & (!g51) & (!sk[105]) & (g118)) + ((g10) & (g51) & (!sk[105]) & (!g118)));
	assign g302 = (((g159) & (!g66) & (!g192) & (!g294) & (!sk[106]) & (!g301)) + ((!g159) & (!g66) & (g192) & (!g294) & (!sk[106]) & (!g301)) + ((g159) & (!g66) & (g192) & (!g294) & (!sk[106]) & (g301)));
	assign g303 = (((g96) & (!g84) & (!g179) & (!g233) & (!sk[107]) & (!g302)) + ((!g96) & (!g84) & (g179) & (!g233) & (!sk[107]) & (!g302)) + ((g96) & (g84) & (g179) & (g233) & (!sk[107]) & (g302)));
	assign g304 = (((!g171) & (!sk[108]) & (g162) & (!g217)) + ((g171) & (!sk[108]) & (!g162) & (g217)));
	assign g305 = (((!i_3_) & (!g12) & (!i_1_) & (i_0_) & (!i_2_) & (!g142)) + ((!i_3_) & (!g12) & (!i_1_) & (!i_0_) & (i_2_) & (!g142)) + ((!i_3_) & (!g12) & (!i_1_) & (i_0_) & (i_2_) & (!g142)) + ((!i_3_) & (!g12) & (i_1_) & (!i_0_) & (!i_2_) & (!g142)) + ((!i_3_) & (!g12) & (i_1_) & (!i_0_) & (!i_2_) & (!g142)) + ((i_3_) & (!g12) & (!i_1_) & (!i_0_) & (!i_2_) & (!g142)));
	assign g306 = (((g39) & (!g79) & (!sk[110]) & (!g80) & (!g241) & (!g305)) + ((!g39) & (!g79) & (!sk[110]) & (g80) & (!g241) & (!g305)) + ((!g39) & (!g79) & (sk[110]) & (!g80) & (g241) & (g305)) + ((!g39) & (g79) & (sk[110]) & (!g80) & (g241) & (g305)));
	assign g307 = (((!sk[111]) & (g304) & (!g265) & (!g289) & (!g299) & (!g306)) + ((!sk[111]) & (!g304) & (!g265) & (g289) & (!g299) & (!g306)) + ((!sk[111]) & (g304) & (g265) & (g289) & (g299) & (g306)));
	assign g308 = (((!g25) & (!g21) & (!g19) & (!i_6_) & (g299) & (g18)) + ((!g25) & (!g21) & (!g19) & (i_6_) & (g299) & (g18)) + ((g25) & (!g21) & (!g19) & (!i_6_) & (g299) & (g18)));
	assign g309 = (((!i_2_) & (!i_3_) & (g246) & (!g50) & (i_0_) & (!i_1_)) + ((!i_2_) & (!i_3_) & (g246) & (!g50) & (!i_0_) & (i_1_)) + ((!i_2_) & (!i_3_) & (g246) & (!g50) & (!i_0_) & (!i_1_)) + ((!i_2_) & (i_3_) & (g246) & (!g50) & (!i_0_) & (!i_1_)));
	assign g310 = (((!sk[114]) & (i_3_) & (!i_5_) & (!i_4_) & (!i_6_) & (!g17)) + ((!sk[114]) & (!i_3_) & (!i_5_) & (i_4_) & (!i_6_) & (!g17)) + ((sk[114]) & (!i_3_) & (!i_5_) & (!i_4_) & (!i_6_) & (g17)) + ((!sk[114]) & (i_3_) & (!i_5_) & (!i_4_) & (!i_6_) & (g17)));
	assign g311 = (((!sk[115]) & (g312) & (!g313)) + ((sk[115]) & (!g312) & (!g313)));
	assign g312 = (((!sk[116]) & (i_6_) & (!g314)) + ((sk[116]) & (!i_6_) & (g314)));
	assign g313 = (((!sk[117]) & (i_6_) & (!g317)) + ((!sk[117]) & (i_6_) & (g317)));
	assign g314 = (((!sk[118]) & (g315) & (!g316)) + ((sk[118]) & (!g315) & (!g316)));
	assign g315 = (((!sk[119]) & (i_3_) & (!g319)) + ((sk[119]) & (!i_3_) & (g319)));
	assign g316 = (((!sk[120]) & (i_3_) & (!g320)) + ((!sk[120]) & (i_3_) & (g320)));
	assign g317 = (((i_3_) & (!sk[121]) & (!g318)) + ((i_3_) & (!sk[121]) & (!g318)));
	assign g318 = (((i_3_) & (!sk[122]) & (!g321)) + ((i_3_) & (!sk[122]) & (g321)));
	assign g319 = (((!i_5_) & (!sk[123]) & (g27) & (!i_4_)) + ((i_5_) & (sk[123]) & (!g27) & (!i_4_)) + ((i_5_) & (!sk[123]) & (!g27) & (i_4_)) + ((!i_5_) & (sk[123]) & (!g27) & (i_4_)));
	assign g320 = (((!sk[124]) & (g31) & (!i_4_)) + ((sk[124]) & (!g31) & (!i_4_)));
	assign g321 = (((i_7_) & (!i_5_) & (g31) & (!sk[125]) & (!i_4_)) + ((!i_7_) & (!i_5_) & (g31) & (!sk[125]) & (!i_4_)) + ((!i_7_) & (!i_5_) & (g31) & (!sk[125]) & (i_4_)) + ((i_7_) & (!i_5_) & (!g31) & (!sk[125]) & (i_4_)) + ((!i_7_) & (!i_5_) & (!g31) & (sk[125]) & (!i_4_)));
	assign g322 = (((!sk[126]) & (g323) & (!g324)) + ((sk[126]) & (!g323) & (!g324)));
	assign g323 = (((i_6_) & (!sk[127]) & (!g325)) + ((!i_6_) & (sk[127]) & (g325)));
	assign g324 = (((!sk[0]) & (i_6_) & (!g328)) + ((!sk[0]) & (i_6_) & (g328)));
	assign g325 = (((g326) & (!sk[1]) & (!g327)) + ((!g326) & (sk[1]) & (!g327)));
	assign g326 = (((!sk[2]) & (i_3_) & (!g330)) + ((sk[2]) & (!i_3_) & (g330)));
	assign g327 = (((i_3_) & (!sk[3]) & (!g331)) + ((i_3_) & (!sk[3]) & (g331)));
	assign g328 = (((!sk[4]) & (i_3_) & (!g329)) + ((!sk[4]) & (i_3_) & (!g329)));
	assign g329 = (((i_3_) & (!sk[5]) & (!g332)) + ((i_3_) & (!sk[5]) & (g332)));
	assign g330 = (((!i_5_) & (!sk[6]) & (i_4_) & (!g27)) + ((i_5_) & (sk[6]) & (!i_4_) & (!g27)) + ((i_5_) & (!sk[6]) & (!i_4_) & (g27)) + ((!i_5_) & (sk[6]) & (!i_4_) & (g27)));
	assign g331 = (((!sk[7]) & (!i_5_) & (i_4_) & (!g25)) + ((!sk[7]) & (i_5_) & (i_4_) & (!g25)) + ((sk[7]) & (!i_5_) & (!i_4_) & (g25)) + ((!sk[7]) & (i_5_) & (!i_4_) & (g25)));
	assign g332 = (((!i_5_) & (!sk[8]) & (!i_4_) & (i_7_) & (!g25)) + ((i_5_) & (!sk[8]) & (!i_4_) & (!i_7_) & (g25)) + ((!i_5_) & (sk[8]) & (!i_4_) & (!i_7_) & (g25)) + ((i_5_) & (sk[8]) & (i_4_) & (!i_7_) & (!g25)) + ((!i_5_) & (sk[8]) & (!i_4_) & (!i_7_) & (!g25)));
	assign g333 = (((g334) & (!sk[9]) & (!g335)) + ((!g334) & (sk[9]) & (!g335)));
	assign g334 = (((!sk[10]) & (g39) & (!g336)) + ((sk[10]) & (!g39) & (g336)));
	assign g335 = (((g39) & (!sk[11]) & (!g339)) + ((g39) & (!sk[11]) & (g339)));
	assign g336 = (((!sk[12]) & (g337) & (!g338)) + ((sk[12]) & (!g337) & (!g338)));
	assign g337 = (((g7) & (!sk[13]) & (!g340)) + ((!g7) & (sk[13]) & (g340)));
	assign g338 = (((g7) & (!sk[14]) & (!g341)) + ((g7) & (!sk[14]) & (g341)));
	assign g339 = (((g7) & (!sk[15]) & (!g342)) + ((g7) & (!sk[15]) & (g342)));
	assign g340 = (((!g149) & (g150) & (!sk[16]) & (!g25)) + ((g149) & (g150) & (!sk[16]) & (g25)) + ((g149) & (!g150) & (!sk[16]) & (g25)));
	assign g341 = (((!sk[17]) & (g149) & (!g150)) + ((!sk[17]) & (g149) & (g150)));
	assign g342 = (((!g149) & (!g150) & (!sk[18]) & (g38) & (!g79)) + ((g149) & (!g150) & (!sk[18]) & (!g38) & (g79)) + ((g149) & (g150) & (!sk[18]) & (!g38) & (g79)));
	assign g343 = (((!sk[19]) & (g344) & (!g345)) + ((sk[19]) & (!g344) & (!g345)));
	assign g344 = (((!sk[20]) & (i_4_) & (!g346)) + ((sk[20]) & (!i_4_) & (g346)));
	assign g345 = (((i_4_) & (!sk[21]) & (!g349)) + ((i_4_) & (!sk[21]) & (g349)));
	assign g346 = (((!sk[22]) & (g347) & (!g348)) + ((sk[22]) & (!g347) & (!g348)));
	assign g347 = (((i_3_) & (!sk[23]) & (!g13)) + ((!i_3_) & (sk[23]) & (!g13)));
	assign g348 = (((i_3_) & (!sk[24]) & (!g352)) + ((i_3_) & (!sk[24]) & (g352)));
	assign g349 = (((!sk[25]) & (g350) & (!g351)) + ((sk[25]) & (!g350) & (!g351)));
	assign g350 = (((!sk[26]) & (i_3_) & (!g353)) + ((sk[26]) & (!i_3_) & (g353)));
	assign g351 = (((i_3_) & (!sk[27]) & (!g39)) + ((i_3_) & (!sk[27]) & (!g39)));
	assign g352 = (((!g39) & (!i_7_) & (!i_6_) & (sk[28]) & (!i_5_)) + ((!g39) & (!i_7_) & (!i_6_) & (sk[28]) & (!i_5_)) + ((g39) & (!i_7_) & (!i_6_) & (!sk[28]) & (i_5_)) + ((!g39) & (!i_7_) & (i_6_) & (!sk[28]) & (!i_5_)) + ((g39) & (!i_7_) & (!i_6_) & (!sk[28]) & (i_5_)));
	assign g353 = (((!g13) & (sk[29]) & (!i_5_)) + ((g13) & (!sk[29]) & (!i_5_)) + ((!g13) & (sk[29]) & (i_5_)));
	assign g354 = (((!sk[30]) & (g355) & (!g356)) + ((sk[30]) & (!g355) & (!g356)));
	assign g355 = (((g23) & (!sk[31]) & (!g357)) + ((!g23) & (sk[31]) & (g357)));
	assign g356 = (((g23) & (!sk[32]) & (!g360)) + ((g23) & (!sk[32]) & (g360)));
	assign g357 = (((g358) & (!sk[33]) & (!g359)) + ((!g358) & (sk[33]) & (!g359)));
	assign g358 = (((!sk[34]) & (i_3_) & (!g362)) + ((sk[34]) & (!i_3_) & (g362)));
	assign g359 = (((i_3_) & (!sk[35]) & (!g363)) + ((i_3_) & (!sk[35]) & (g363)));
	assign g360 = (((i_3_) & (!sk[36]) & (!g361)) + ((!i_3_) & (sk[36]) & (!g361)));
	assign g361 = (((!sk[37]) & (i_3_) & (!g364)) + ((sk[37]) & (!i_3_) & (g364)));
	assign g362 = (((!sk[38]) & (!i_5_) & (!i_6_) & (g31) & (!i_4_)) + ((sk[38]) & (i_5_) & (!i_6_) & (!g31) & (!i_4_)) + ((sk[38]) & (!i_5_) & (i_6_) & (!g31) & (!i_4_)) + ((sk[38]) & (!i_5_) & (!i_6_) & (!g31) & (i_4_)) + ((!sk[38]) & (i_5_) & (!i_6_) & (!g31) & (i_4_)));
	assign g363 = (((!i_5_) & (!i_6_) & (i_7_) & (!sk[39]) & (!i_4_)) + ((i_5_) & (!i_6_) & (!i_7_) & (!sk[39]) & (i_4_)) + ((!i_5_) & (!i_6_) & (!i_7_) & (sk[39]) & (!i_4_)) + ((!i_5_) & (!i_6_) & (!i_7_) & (sk[39]) & (!i_4_)) + ((!i_5_) & (!i_6_) & (!i_7_) & (sk[39]) & (!i_4_)));
	assign g364 = (((!i_5_) & (!sk[40]) & (!i_6_) & (g31) & (!i_4_)) + ((i_5_) & (sk[40]) & (!i_6_) & (!g31) & (!i_4_)) + ((!i_5_) & (sk[40]) & (i_6_) & (!g31) & (!i_4_)) + ((i_5_) & (!sk[40]) & (!i_6_) & (!g31) & (i_4_)) + ((!i_5_) & (sk[40]) & (!i_6_) & (!g31) & (i_4_)));
	assign g365 = (((!sk[41]) & (i_1_) & (!g366)) + ((sk[41]) & (!i_1_) & (g366)));
	assign g366 = (((g367) & (!sk[42]) & (!g368)) + ((!g367) & (sk[42]) & (!g368)));
	assign g367 = (((!sk[43]) & (i_5_) & (!g369)) + ((sk[43]) & (!i_5_) & (g369)));
	assign g368 = (((!sk[44]) & (i_5_) & (!g370)) + ((!sk[44]) & (i_5_) & (g370)));
	assign g369 = (((!i_4_) & (!i_2_) & (i_6_) & (!sk[45]) & (!i_0_)) + ((i_4_) & (!i_2_) & (!i_6_) & (!sk[45]) & (i_0_)) + ((!i_4_) & (!i_2_) & (!i_6_) & (sk[45]) & (i_0_)));
	assign g370 = (((!sk[46]) & (!i_4_) & (!i_2_) & (i_3_) & (!i_0_)) + ((!sk[46]) & (i_4_) & (!i_2_) & (!i_3_) & (i_0_)) + ((!sk[46]) & (i_4_) & (!i_2_) & (!i_3_) & (i_0_)) + ((sk[46]) & (i_4_) & (!i_2_) & (!i_3_) & (!i_0_)) + ((!sk[46]) & (i_4_) & (i_2_) & (i_3_) & (!i_0_)));

endmodule